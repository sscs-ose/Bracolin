* NGSPICE file created from PR_pfets.ext - technology: gf180mcuD

.subckt PR_pfets VS2_A VG VS2_B VC_A VC_B VS1 VD1 VB
X0 VB.t71 VB.t70 VB.t71 VB.t4 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1 VB.t69 VB.t68 VB.t69 VB.t1 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2 VS2_A VG.t0 a_1844_3098# VB.t4 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3 VD1 VG.t1 a_1844_1166# VB.t4 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4 VB.t67 VB.t66 VB.t67 VB.t7 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5 VB.t65 VB.t64 VB.t65 VB.t26 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6 a_438_3098# VG.t2 VS2_B.t0 VB.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X7 VD1 VG.t3 a_1844_1932# VB.t4 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X8 a_438_1166# VG.t4 VD1.t2 VB.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X9 VC_A VG.t5 a_438_0# VB.t56 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X10 VB.t63 VB.t62 VB.t63 VB.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X11 VB.t61 VB.t60 VB.t61 VB.t29 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X12 VB.t59 VB.t58 VB.t59 VB.t26 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X13 a_438_1932# VG.t6 VD1.t3 VB.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X14 VB.t57 VB.t55 VB.t57 VB.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X15 VB.t54 VB.t53 VB.t54 VB.t29 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X16 VB.t52 VB.t51 VB.t52 VB.t26 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X17 VB.t50 VB.t49 VB.t50 VB.t10 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X18 VB.t48 VB.t47 VB.t48 VB.t7 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X19 VB.t46 VB.t45 VB.t46 VB.t29 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X20 VC_B VG.t7 a_438_3098# VB.t56 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X21 VB.t44 VB.t43 VB.t44 VB.t29 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X22 VS1 VG.t8 a_438_1166# VB.t56 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X23 VB.t42 VB.t41 VB.t42 VB.t29 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X24 VB.t40 VB.t39 VB.t40 VB.t26 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X25 VB.t38 VB.t37 VB.t38 VB.t26 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X26 VB.t36 VB.t35 VB.t36 VB.t7 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X27 VB.t34 VB.t33 VB.t34 VB.t10 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X28 VS2_B VG.t9 a_1844_0# VB.t4 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X29 VB.t32 VB.t31 VB.t32 VB.t21 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X30 VS1 VG.t10 a_438_1932# VB.t56 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X31 VB.t30 VB.t28 VB.t30 VB.t29 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X32 VB.t27 VB.t25 VB.t27 VB.t26 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X33 VB.t24 VB.t23 VB.t24 VB.t10 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X34 VB.t22 VB.t20 VB.t22 VB.t21 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X35 VB.t19 VB.t18 VB.t19 VB.t7 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X36 VB.t17 VB.t16 VB.t17 VB.t10 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X37 VB.t15 VB.t14 VB.t15 VB.t10 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X38 VB.t13 VB.t12 VB.t13 VB.t7 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X39 VB.t11 VB.t9 VB.t11 VB.t10 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X40 VB.t8 VB.t6 VB.t8 VB.t7 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X41 a_1844_0# VG.t11 VC_B.t1 VB.t21 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X42 a_1844_3098# VG.t12 VC_A.t1 VB.t21 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X43 a_1844_1166# VG.t13 VS1.t0 VB.t21 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X44 VB.t5 VB.t3 VB.t5 VB.t4 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X45 a_438_0# VG.t14 VS2_A.t0 VB.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X46 a_1844_1932# VG.t15 VS1.t1 VB.t21 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X47 VB.t2 VB.t0 VB.t2 VB.t1 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
R0 VB.n61 VB.n5 477.971
R1 VB.n58 VB.n6 470.842
R2 VB.n61 VB.n6 470.842
R3 VB.n58 VB.n5 469.683
R4 VB.t4 VB.t29 142.035
R5 VB.t1 VB.t10 142.035
R6 VB.t29 VB.t26 96.2717
R7 VB.t21 VB.t4 96.2717
R8 VB.t56 VB.t1 96.2717
R9 VB.t10 VB.t7 96.2717
R10 VB.t26 VB.n5 80.6158
R11 VB.t7 VB.n6 80.6158
R12 VB.n59 VB.t21 69.831
R13 VB.n60 VB.t56 63.7293
R14 VB.n60 VB.n59 8.47508
R15 VB.n20 VB.t53 8.10567
R16 VB.n20 VB.t51 8.10567
R17 VB.n18 VB.t43 8.10567
R18 VB.n18 VB.t39 8.10567
R19 VB.n17 VB.t28 8.10567
R20 VB.n17 VB.t25 8.10567
R21 VB.n13 VB.t41 8.10567
R22 VB.n13 VB.t37 8.10567
R23 VB.n12 VB.t45 8.10567
R24 VB.n12 VB.t64 8.10567
R25 VB.n69 VB.t60 8.10567
R26 VB.n69 VB.t58 8.10567
R27 VB.n53 VB.t68 8.10567
R28 VB.n27 VB.t55 8.10567
R29 VB.n7 VB.t20 8.10567
R30 VB.n23 VB.t70 8.10567
R31 VB.n50 VB.t35 8.10567
R32 VB.n50 VB.t33 8.10567
R33 VB.n48 VB.t18 8.10567
R34 VB.n48 VB.t16 8.10567
R35 VB.n47 VB.t6 8.10567
R36 VB.n47 VB.t9 8.10567
R37 VB.n43 VB.t12 8.10567
R38 VB.n43 VB.t14 8.10567
R39 VB.n42 VB.t66 8.10567
R40 VB.n42 VB.t23 8.10567
R41 VB.n40 VB.t47 8.10567
R42 VB.n40 VB.t49 8.10567
R43 VB.n34 VB.t0 8.10567
R44 VB.n35 VB.t62 8.10567
R45 VB.n64 VB.t31 8.10567
R46 VB.n3 VB.t3 8.10567
R47 VB.n52 VB.t69 3.20383
R48 VB.n56 VB.t57 3.20383
R49 VB.n26 VB.t22 3.20383
R50 VB.n22 VB.t71 3.20383
R51 VB.n38 VB.t2 3.20383
R52 VB.t63 VB.n4 3.20383
R53 VB.n63 VB.t32 3.20383
R54 VB.n67 VB.t5 3.20383
R55 VB.n66 VB.n65 1.73383
R56 VB.n37 VB.n36 1.73383
R57 VB.n25 VB.n24 1.73383
R58 VB.n55 VB.n54 1.73383
R59 VB.t57 VB.n55 1.4705
R60 VB.n55 VB.t69 1.4705
R61 VB.n25 VB.t71 1.4705
R62 VB.t22 VB.n25 1.4705
R63 VB.n37 VB.t63 1.4705
R64 VB.t2 VB.n37 1.4705
R65 VB.t5 VB.n66 1.4705
R66 VB.n66 VB.t32 1.4705
R67 VB.n8 VB.t52 1.00929
R68 VB.n9 VB.t40 1.00929
R69 VB.n10 VB.t27 1.00929
R70 VB.n11 VB.t38 1.00929
R71 VB.n0 VB.t65 1.00929
R72 VB.n2 VB.t59 1.00929
R73 VB.n28 VB.t34 1.00929
R74 VB.n29 VB.t17 1.00929
R75 VB.n30 VB.t11 1.00929
R76 VB.n31 VB.t15 1.00929
R77 VB.n32 VB.t24 1.00929
R78 VB.n33 VB.t50 1.00929
R79 VB.n8 VB.t54 1.00871
R80 VB.n9 VB.t44 1.00871
R81 VB.n10 VB.t30 1.00871
R82 VB.n11 VB.t42 1.00871
R83 VB.n0 VB.t46 1.00871
R84 VB.n2 VB.t61 1.00871
R85 VB.n28 VB.t36 1.00871
R86 VB.n29 VB.t19 1.00871
R87 VB.n30 VB.t8 1.00871
R88 VB.n31 VB.t13 1.00871
R89 VB.n32 VB.t67 1.00871
R90 VB.n33 VB.t48 1.00871
R91 VB.n51 VB.n28 0.470768
R92 VB.n21 VB.n8 0.470735
R93 VB.n39 VB.n33 0.468749
R94 VB.n41 VB.n32 0.468749
R95 VB.n44 VB.n31 0.468749
R96 VB.n46 VB.n30 0.468749
R97 VB.n49 VB.n29 0.468749
R98 VB.n68 VB.n2 0.468749
R99 VB.n1 VB.n0 0.468749
R100 VB.n14 VB.n11 0.468749
R101 VB.n16 VB.n10 0.468749
R102 VB.n19 VB.n9 0.468749
R103 VB.n45 VB.n6 0.10728
R104 VB.n58 VB.n57 0.10728
R105 VB.n59 VB.n58 0.10728
R106 VB.n15 VB.n5 0.10728
R107 VB.n62 VB.n61 0.1055
R108 VB.n61 VB.n60 0.1055
R109 VB.n50 VB.n49 0.0382419
R110 VB.n41 VB.n40 0.0382419
R111 VB.n20 VB.n19 0.0376172
R112 VB.n48 VB.n47 0.0364748
R113 VB.n43 VB.n42 0.0364748
R114 VB.n18 VB.n17 0.0358793
R115 VB.n13 VB.n12 0.0358793
R116 VB.n39 VB.n38 0.0308563
R117 VB.n68 VB.n67 0.0307435
R118 VB.n67 VB.n3 0.0293162
R119 VB.n65 VB.n3 0.0293162
R120 VB.n65 VB.n64 0.0293162
R121 VB.n64 VB.n63 0.0293162
R122 VB.n35 VB.n4 0.0293162
R123 VB.n36 VB.n35 0.0293162
R124 VB.n36 VB.n34 0.0293162
R125 VB.n38 VB.n34 0.0293162
R126 VB.n23 VB.n22 0.0293162
R127 VB.n24 VB.n23 0.0293162
R128 VB.n24 VB.n7 0.0293162
R129 VB.n26 VB.n7 0.0293162
R130 VB.n56 VB.n27 0.0293162
R131 VB.n54 VB.n27 0.0293162
R132 VB.n54 VB.n53 0.0293162
R133 VB.n53 VB.n52 0.0293162
R134 VB.n46 VB.n45 0.0270708
R135 VB.n16 VB.n15 0.026631
R136 VB.n22 VB.n21 0.02404
R137 VB.n52 VB.n51 0.02404
R138 VB VB.n1 0.0233414
R139 VB.n45 VB.n44 0.0222742
R140 VB.n15 VB.n14 0.0219138
R141 VB.n49 VB.n48 0.0193079
R142 VB.n47 VB.n46 0.0193079
R143 VB.n44 VB.n43 0.0193079
R144 VB.n42 VB.n41 0.0193079
R145 VB.n40 VB.n39 0.0193079
R146 VB.n19 VB.n18 0.0189966
R147 VB.n17 VB.n16 0.0189966
R148 VB.n14 VB.n13 0.0189966
R149 VB.n12 VB.n1 0.0189966
R150 VB.n69 VB.n68 0.0189966
R151 VB.n63 VB.n62 0.0185609
R152 VB.n51 VB.n50 0.0172882
R153 VB.n21 VB.n20 0.0170103
R154 VB.n57 VB.n56 0.0149081
R155 VB VB.n69 0.0147759
R156 VB.n57 VB.n26 0.0134876
R157 VB.n62 VB.n4 0.00983484
R158 VG.n28 VG.t6 8.17385
R159 VG.n38 VG.t4 8.17299
R160 VG.n60 VG.t14 8.17134
R161 VG.n2 VG.t2 8.16754
R162 VG.n18 VG.t3 8.15339
R163 VG.n35 VG.t1 8.15277
R164 VG.n50 VG.t9 8.15161
R165 VG.n5 VG.t0 8.14892
R166 VG.n57 VG.t5 8.10567
R167 VG.n43 VG.t13 8.10567
R168 VG.n11 VG.t12 8.10567
R169 VG.n22 VG.t15 8.10567
R170 VG.n25 VG.t10 8.10567
R171 VG.n9 VG.t7 8.10567
R172 VG.n54 VG.t11 8.10567
R173 VG.n37 VG.t8 8.10567
R174 VG.n23 VG.n22 4.62603
R175 VG.n44 VG.n43 4.6244
R176 VG.n55 VG.n54 4.62126
R177 VG.n12 VG.n11 4.61407
R178 VG.n26 VG.n1 4.5005
R179 VG.n21 VG.n4 4.5005
R180 VG.n20 VG.n19 4.5005
R181 VG.n13 VG.n6 4.5005
R182 VG.n15 VG.n14 4.5005
R183 VG.n8 VG.n7 4.5005
R184 VG.n53 VG.n34 4.5005
R185 VG.n52 VG.n51 4.5005
R186 VG.n47 VG.n46 4.5005
R187 VG.n45 VG.n36 4.5005
R188 VG.n41 VG.n40 4.5005
R189 VG.n58 VG.n32 4.5005
R190 VG.n25 VG.n24 2.26271
R191 VG.n42 VG.n37 2.26206
R192 VG.n57 VG.n56 2.26082
R193 VG.n10 VG.n9 2.25797
R194 VG.n14 VG.n5 1.97162
R195 VG.n51 VG.n50 1.97099
R196 VG.n19 VG.n18 1.97058
R197 VG.n46 VG.n35 1.97031
R198 VG.n2 VG.n0 1.9364
R199 VG.n61 VG.n60 1.93496
R200 VG.n39 VG.n38 1.93434
R201 VG.n29 VG.n28 1.93401
R202 VG.n30 VG.n0 1.67564
R203 VG.n30 VG.n29 1.5005
R204 VG.n62 VG.n61 1.5005
R205 VG.n39 VG.n31 1.5005
R206 VG.n24 VG.n23 0.834997
R207 VG.n44 VG.n42 0.834981
R208 VG.n56 VG.n55 0.83495
R209 VG.n12 VG.n10 0.834879
R210 VG.n27 VG.n3 0.618
R211 VG.n17 VG.n16 0.618
R212 VG.n49 VG.n48 0.613
R213 VG.n59 VG.n33 0.613
R214 VG.n31 VG.n30 0.415534
R215 VG.n18 VG.n17 0.291089
R216 VG.n48 VG.n35 0.263985
R217 VG.n16 VG.n5 0.263649
R218 VG.n50 VG.n49 0.257367
R219 VG.n40 VG.n33 0.249461
R220 VG.n28 VG.n27 0.248085
R221 VG.n59 VG.n58 0.243158
R222 VG VG.n62 0.23827
R223 VG.n10 VG.n7 0.234321
R224 VG.n56 VG.n32 0.234252
R225 VG.n42 VG.n41 0.234222
R226 VG.n24 VG.n1 0.234207
R227 VG.n3 VG.n2 0.224813
R228 VG.n27 VG.n26 0.223132
R229 VG.n38 VG.n33 0.215694
R230 VG.n8 VG.n3 0.201929
R231 VG.n48 VG.n47 0.186344
R232 VG.n60 VG 0.184128
R233 VG.n52 VG.n49 0.181639
R234 VG.n62 VG.n31 0.171986
R235 VG.n20 VG.n17 0.165105
R236 VG.n19 VG.n4 0.157683
R237 VG.n23 VG.n4 0.157683
R238 VG.n14 VG.n13 0.157683
R239 VG.n13 VG.n12 0.157683
R240 VG.n51 VG.n34 0.157683
R241 VG.n55 VG.n34 0.157683
R242 VG.n46 VG.n45 0.157683
R243 VG.n45 VG.n44 0.157683
R244 VG.n16 VG.n15 0.149429
R245 VG.n21 VG.n20 0.147342
R246 VG.n47 VG.n36 0.145435
R247 VG.n53 VG.n52 0.141766
R248 VG.n15 VG.n6 0.133357
R249 VG.n26 VG.n25 0.133132
R250 VG.n40 VG.n37 0.131409
R251 VG.n58 VG.n57 0.128095
R252 VG.n9 VG.n8 0.1205
R253 VG VG.n59 0.0267025
R254 VG.n29 VG.n1 0.0220493
R255 VG.n7 VG.n0 0.0220493
R256 VG.n61 VG.n32 0.0220493
R257 VG.n41 VG.n39 0.0220493
R258 VG.n22 VG.n21 0.0218158
R259 VG.n43 VG.n36 0.021539
R260 VG.n54 VG.n53 0.0210063
R261 VG.n11 VG.n6 0.0197857
R262 VS2_A.n1 VS2_A.n0 11.7531
R263 VS2_A.n1 VS2_A 4.90596
R264 VS2_A VS2_A.t0 3.61831
R265 VS2_A VS2_A.n1 0.3335
R266 VD1.n4 VD1.n3 4.84877
R267 VD1.n3 VD1.t3 3.65383
R268 VD1.n2 VD1.n0 3.65146
R269 VD1.n3 VD1.t2 3.57094
R270 VD1 VD1.n1 3.51291
R271 VD1 VD1.n4 2.98263
R272 VD1.n4 VD1.n2 2.71171
R273 VD1.n2 VD1 0.0608947
R274 VS2_B.n1 VS2_B.t0 12.1613
R275 VS2_B.n1 VS2_B 4.97994
R276 VS2_B VS2_B.n0 3.61831
R277 VS2_B VS2_B.n1 0.42663
R278 VC_A.n1 VC_A.t1 10.1798
R279 VC_A.n1 VC_A 4.63333
R280 VC_A VC_A.n0 3.51291
R281 VC_A VC_A.n1 0.0734
R282 VC_B.n1 VC_B.n0 9.63183
R283 VC_B.n1 VC_B 4.98908
R284 VC_B VC_B.t1 3.47265
R285 VC_B VC_B.n1 0.47975
R286 VS1 VS1.n4 4.36237
R287 VS1.n0 VS1.t0 3.73318
R288 VS1.n3 VS1.n2 3.73318
R289 VS1.n3 VS1.n1 3.4916
R290 VS1 VS1.t1 3.47383
R291 VS1.n4 VS1.n3 0.174974
R292 VS1.n4 VS1.n0 0.130788
R293 VS1.n0 VS1 0.0182632
C0 a_1844_1166# VD1 0.062843f
C1 a_438_1932# VG 0.15726f
C2 VB a_438_3098# 0.025718f
C3 VC_B a_1844_0# 0.029601f
C4 VC_A a_1844_0# 0.014894f
C5 VC_B VC_A 2.30852f
C6 VC_A a_1844_3098# 0.042568f
C7 VS2_B a_1844_0# 0.031455f
C8 VG a_1844_0# 0.130094f
C9 VS2_B VC_B 2.11591f
C10 VC_B VG 1.21933f
C11 VG a_1844_3098# 0.132974f
C12 VB VS2_A 1.303f
C13 VS2_B VC_A 0.219687f
C14 VG VC_A 2.59073f
C15 VB VS1 1.12283f
C16 VS2_B VG 2.86536f
C17 VB VD1 1.11211f
C18 VB a_438_0# 0.021515f
C19 a_438_1932# VS2_A 0.01182f
C20 a_438_1932# VS1 0.04473f
C21 VC_B a_438_3098# 0.02829f
C22 a_438_3098# VC_A 0.016091f
C23 a_438_1932# VD1 0.029183f
C24 VS2_B a_438_3098# 0.02829f
C25 a_438_3098# VG 0.158238f
C26 VG a_438_1166# 0.157264f
C27 VS1 a_1844_0# 0.013613f
C28 VC_B VS2_A 2.19085f
C29 a_1844_3098# VS2_A 0.02829f
C30 VC_A VS2_A 0.29118f
C31 VS1 VC_B 1.72732f
C32 VS1 a_1844_3098# 0.013613f
C33 VS1 VC_A 0.39497f
C34 VS2_B VS2_A 0.357159f
C35 VG VS2_A 4.61911f
C36 VD1 a_1844_0# 0.021476f
C37 VS2_B VS1 0.182793f
C38 VC_B VD1 0.191679f
C39 VS1 VG 1.46282f
C40 VD1 a_1844_3098# 0.02151f
C41 VD1 VC_A 0.241135f
C42 a_438_0# VC_A 0.043765f
C43 a_1844_1932# VG 0.1317f
C44 a_1844_1166# VG 0.131658f
C45 VS2_B VD1 1.70058f
C46 VD1 VG 1.30476f
C47 a_438_0# VG 0.15567f
C48 a_438_3098# VS2_A 0.01182f
C49 a_438_1166# VS2_A 0.01182f
C50 VS1 a_438_1166# 0.028915f
C51 VD1 a_438_1166# 0.041194f
C52 VS1 VS2_A 0.204565f
C53 VB a_1844_0# 0.021515f
C54 VB VC_B 0.895169f
C55 VB a_1844_3098# 0.025718f
C56 VB VC_A 1.76889f
C57 a_1844_1932# VS1 0.058343f
C58 a_1844_1166# VS1 0.042528f
C59 VD1 VS2_A 0.281431f
C60 a_438_0# VS2_A 0.040109f
C61 VS1 VD1 2.62467f
C62 VS2_B VB 1.73079f
C63 VB VG 10.4278f
C64 a_1844_1932# VD1 0.050814f
C65 VS1 a_1426_n1526# 2.286416f
C66 VD1 a_1426_n1526# 1.408236f
C67 VS2_A a_1426_n1526# 1.407576f
C68 VC_A a_1426_n1526# 1.310399f
C69 VC_B a_1426_n1526# 1.746819f
C70 VS2_B a_1426_n1526# 1.229475f
C71 VG a_1426_n1526# 3.806466f
C72 VB a_1426_n1526# 0.115827p
C73 VS1.t0 a_1426_n1526# 0.058936f
C74 VS1.t1 a_1426_n1526# 0.054098f
C75 VS1.n0 a_1426_n1526# 0.106711f
C76 VS1.n1 a_1426_n1526# 0.054397f
C77 VS1.n2 a_1426_n1526# 0.058936f
C78 VS1.n3 a_1426_n1526# 0.183843f
C79 VS1.n4 a_1426_n1526# 0.341766f
C80 VC_B.n0 a_1426_n1526# 0.800726f
C81 VC_B.t1 a_1426_n1526# 0.167323f
C82 VC_B.n1 a_1426_n1526# 3.93205f
C83 VC_A.t1 a_1426_n1526# 0.71089f
C84 VC_A.n0 a_1426_n1526# 0.129424f
C85 VC_A.n1 a_1426_n1526# 3.11041f
C86 VS2_B.t0 a_1426_n1526# 0.63032f
C87 VS2_B.n0 a_1426_n1526# 0.131883f
C88 VS2_B.n1 a_1426_n1526# 3.27009f
C89 VD1.n0 a_1426_n1526# 0.071501f
C90 VD1.n1 a_1426_n1526# 0.068326f
C91 VD1.n2 a_1426_n1526# 0.125926f
C92 VD1.t2 a_1426_n1526# 0.069612f
C93 VD1.t3 a_1426_n1526# 0.071558f
C94 VD1.n3 a_1426_n1526# 0.271735f
C95 VD1.n4 a_1426_n1526# 0.542154f
C96 VS2_A.n0 a_1426_n1526# 0.856096f
C97 VS2_A.t0 a_1426_n1526# 0.184022f
C98 VS2_A.n1 a_1426_n1526# 4.61084f
C99 VG.n0 a_1426_n1526# 0.259422f
C100 VG.n1 a_1426_n1526# 0.028667f
C101 VG.t6 a_1426_n1526# 0.511623f
C102 VG.t2 a_1426_n1526# 0.511482f
C103 VG.n2 a_1426_n1526# 0.300291f
C104 VG.n3 a_1426_n1526# 0.128374f
C105 VG.n4 a_1426_n1526# 0.031998f
C106 VG.t0 a_1426_n1526# 0.510946f
C107 VG.n5 a_1426_n1526# 0.309035f
C108 VG.n6 a_1426_n1526# 0.021676f
C109 VG.n7 a_1426_n1526# 0.028678f
C110 VG.n8 a_1426_n1526# 0.045794f
C111 VG.t7 a_1426_n1526# 0.509584f
C112 VG.n9 a_1426_n1526# 0.252058f
C113 VG.n10 a_1426_n1526# 0.106722f
C114 VG.t12 a_1426_n1526# 0.509584f
C115 VG.n11 a_1426_n1526# 0.229035f
C116 VG.n12 a_1426_n1526# 0.102462f
C117 VG.n13 a_1426_n1526# 0.031998f
C118 VG.n14 a_1426_n1526# 0.147319f
C119 VG.n15 a_1426_n1526# 0.040146f
C120 VG.n16 a_1426_n1526# 0.125211f
C121 VG.n17 a_1426_n1526# 0.119417f
C122 VG.t3 a_1426_n1526# 0.511047f
C123 VG.n18 a_1426_n1526# 0.299311f
C124 VG.n19 a_1426_n1526# 0.147312f
C125 VG.n20 a_1426_n1526# 0.036323f
C126 VG.n21 a_1426_n1526# 0.019611f
C127 VG.t15 a_1426_n1526# 0.509584f
C128 VG.n22 a_1426_n1526# 0.22453f
C129 VG.n23 a_1426_n1526# 0.102472f
C130 VG.n24 a_1426_n1526# 0.106717f
C131 VG.t10 a_1426_n1526# 0.509584f
C132 VG.n25 a_1426_n1526# 0.245316f
C133 VG.n26 a_1426_n1526# 0.041433f
C134 VG.n27 a_1426_n1526# 0.122271f
C135 VG.n28 a_1426_n1526# 0.291564f
C136 VG.n29 a_1426_n1526# 0.13905f
C137 VG.n30 a_1426_n1526# 2.07481f
C138 VG.n31 a_1426_n1526# 1.0376f
C139 VG.n32 a_1426_n1526# 0.028672f
C140 VG.t14 a_1426_n1526# 0.511567f
C141 VG.n33 a_1426_n1526# 0.12289f
C142 VG.n34 a_1426_n1526# 0.031998f
C143 VG.t1 a_1426_n1526# 0.511033f
C144 VG.n35 a_1426_n1526# 0.297585f
C145 VG.n36 a_1426_n1526# 0.019869f
C146 VG.t8 a_1426_n1526# 0.509584f
C147 VG.n37 a_1426_n1526# 0.246158f
C148 VG.t4 a_1426_n1526# 0.511604f
C149 VG.n38 a_1426_n1526# 0.288773f
C150 VG.n39 a_1426_n1526# 0.139054f
C151 VG.n40 a_1426_n1526# 0.045474f
C152 VG.n41 a_1426_n1526# 0.028669f
C153 VG.n42 a_1426_n1526# 0.106718f
C154 VG.t13 a_1426_n1526# 0.509584f
C155 VG.n43 a_1426_n1526# 0.225093f
C156 VG.n44 a_1426_n1526# 0.102471f
C157 VG.n45 a_1426_n1526# 0.031998f
C158 VG.n46 a_1426_n1526# 0.147303f
C159 VG.n47 a_1426_n1526# 0.039597f
C160 VG.n48 a_1426_n1526# 0.119767f
C161 VG.n49 a_1426_n1526# 0.121218f
C162 VG.t9 a_1426_n1526# 0.511007f
C163 VG.n50 a_1426_n1526# 0.299931f
C164 VG.n51 a_1426_n1526# 0.147315f
C165 VG.n52 a_1426_n1526# 0.040626f
C166 VG.n53 a_1426_n1526# 0.020386f
C167 VG.t11 a_1426_n1526# 0.509584f
C168 VG.n54 a_1426_n1526# 0.226219f
C169 VG.n55 a_1426_n1526# 0.102468f
C170 VG.n56 a_1426_n1526# 0.106719f
C171 VG.t5 a_1426_n1526# 0.509584f
C172 VG.n57 a_1426_n1526# 0.247844f
C173 VG.n58 a_1426_n1526# 0.046655f
C174 VG.n59 a_1426_n1526# 0.097988f
C175 VG.n60 a_1426_n1526# 0.287084f
C176 VG.n61 a_1426_n1526# 0.13906f
C177 VG.n62 a_1426_n1526# 0.724009f
C178 VB.n1 a_1426_n1526# 0.079215f
C179 VB.t58 a_1426_n1526# 0.02156f
C180 VB.t3 a_1426_n1526# 0.02156f
C181 VB.n3 a_1426_n1526# 0.046453f
C182 VB.n4 a_1426_n1526# 0.028126f
C183 VB.n5 a_1426_n1526# 0.367597f
C184 VB.n6 a_1426_n1526# 0.358113f
C185 VB.t26 a_1426_n1526# 0.47352f
C186 VB.t29 a_1426_n1526# 0.637785f
C187 VB.t4 a_1426_n1526# 0.637785f
C188 VB.t21 a_1426_n1526# 0.444544f
C189 VB.t20 a_1426_n1526# 0.02156f
C190 VB.n7 a_1426_n1526# 0.046453f
C191 VB.t51 a_1426_n1526# 0.02156f
C192 VB.t39 a_1426_n1526# 0.02156f
C193 VB.t25 a_1426_n1526# 0.02156f
C194 VB.t37 a_1426_n1526# 0.02156f
C195 VB.t64 a_1426_n1526# 0.02156f
C196 VB.t45 a_1426_n1526# 0.02156f
C197 VB.n12 a_1426_n1526# 0.112202f
C198 VB.t41 a_1426_n1526# 0.02156f
C199 VB.n13 a_1426_n1526# 0.112202f
C200 VB.n14 a_1426_n1526# 0.076651f
C201 VB.n15 a_1426_n1526# 0.085395f
C202 VB.n16 a_1426_n1526# 0.085123f
C203 VB.t28 a_1426_n1526# 0.02156f
C204 VB.n17 a_1426_n1526# 0.112202f
C205 VB.t43 a_1426_n1526# 0.02156f
C206 VB.n18 a_1426_n1526# 0.112202f
C207 VB.n19 a_1426_n1526# 0.104856f
C208 VB.t53 a_1426_n1526# 0.02156f
C209 VB.n20 a_1426_n1526# 0.111756f
C210 VB.n21 a_1426_n1526# 0.149015f
C211 VB.n22 a_1426_n1526# 0.037673f
C212 VB.t70 a_1426_n1526# 0.02156f
C213 VB.n23 a_1426_n1526# 0.046453f
C214 VB.n24 a_1426_n1526# 0.038736f
C215 VB.n26 a_1426_n1526# 0.030581f
C216 VB.t55 a_1426_n1526# 0.02156f
C217 VB.n27 a_1426_n1526# 0.046453f
C218 VB.t33 a_1426_n1526# 0.02156f
C219 VB.t16 a_1426_n1526# 0.02156f
C220 VB.t9 a_1426_n1526# 0.02156f
C221 VB.t14 a_1426_n1526# 0.02156f
C222 VB.t23 a_1426_n1526# 0.02156f
C223 VB.t49 a_1426_n1526# 0.02156f
C224 VB.t0 a_1426_n1526# 0.02156f
C225 VB.n34 a_1426_n1526# 0.046453f
C226 VB.t62 a_1426_n1526# 0.02156f
C227 VB.n35 a_1426_n1526# 0.046453f
C228 VB.n36 a_1426_n1526# 0.038736f
C229 VB.n38 a_1426_n1526# 0.065696f
C230 VB.n39 a_1426_n1526# 0.146258f
C231 VB.t47 a_1426_n1526# 0.02156f
C232 VB.n40 a_1426_n1526# 0.11367f
C233 VB.n41 a_1426_n1526# 0.103202f
C234 VB.t66 a_1426_n1526# 0.02156f
C235 VB.n42 a_1426_n1526# 0.1106f
C236 VB.t12 a_1426_n1526# 0.02156f
C237 VB.n43 a_1426_n1526# 0.1106f
C238 VB.n44 a_1426_n1526# 0.075464f
C239 VB.n45 a_1426_n1526# 0.083982f
C240 VB.n46 a_1426_n1526# 0.083797f
C241 VB.t6 a_1426_n1526# 0.02156f
C242 VB.n47 a_1426_n1526# 0.1106f
C243 VB.t18 a_1426_n1526# 0.02156f
C244 VB.n48 a_1426_n1526# 0.1106f
C245 VB.n49 a_1426_n1526# 0.103202f
C246 VB.t35 a_1426_n1526# 0.02156f
C247 VB.n50 a_1426_n1526# 0.110162f
C248 VB.n51 a_1426_n1526# 0.146886f
C249 VB.n52 a_1426_n1526# 0.037673f
C250 VB.t68 a_1426_n1526# 0.02156f
C251 VB.n53 a_1426_n1526# 0.046453f
C252 VB.n54 a_1426_n1526# 0.038736f
C253 VB.n56 a_1426_n1526# 0.031535f
C254 VB.n57 a_1426_n1526# 0.018413f
C255 VB.n58 a_1426_n1526# 0.066736f
C256 VB.n59 a_1426_n1526# 0.209571f
C257 VB.t7 a_1426_n1526# 0.473508f
C258 VB.t10 a_1426_n1526# 0.637785f
C259 VB.t1 a_1426_n1526# 0.637785f
C260 VB.t56 a_1426_n1526# 0.428214f
C261 VB.n60 a_1426_n1526# 0.193241f
C262 VB.n61 a_1426_n1526# 0.067324f
C263 VB.n62 a_1426_n1526# 0.018413f
C264 VB.n63 a_1426_n1526# 0.033991f
C265 VB.t31 a_1426_n1526# 0.02156f
C266 VB.n64 a_1426_n1526# 0.046453f
C267 VB.n65 a_1426_n1526# 0.038736f
C268 VB.n67 a_1426_n1526# 0.065742f
C269 VB.n68 a_1426_n1526# 0.148796f
C270 VB.t60 a_1426_n1526# 0.02156f
C271 VB.n69 a_1426_n1526# 0.074298f
.ends

