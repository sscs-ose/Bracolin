* Extracted by KLayout with GF180MCU LVS runset on : 24/04/2024 20:08

.SUBCKT inverter_PAD DVDD DVSS Y A
M$1 Y A DVDD DVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2 DVDD \$84 \$82 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$3 \$82 \$84 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$4 \$20 \$135 \$82 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$5 \$82 \$135 \$20 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$6 \$84 \$136 \$83 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$7 DVDD \$138 \$84 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$8 \$84 \$139 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$9 \$85 \$83 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$10 DVDD \$83 \$85 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$11 \$49 \$83 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$12 DVDD \$83 \$49 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$13 \$51 \$87 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$14 DVDD \$87 \$51 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$15 \$50 \$87 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$16 DVDD \$87 \$50 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$17 DVDD \$139 \$86 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$18 \$86 \$140 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$19 \$87 \$142 \$86 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$20 \$15 \$135 \$16 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$21 \$16 \$135 \$15 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$22 DVDD \$86 \$16 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$23 \$16 \$86 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$24 DVDD \$90 \$88 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$25 \$88 \$90 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$26 \$17 \$135 \$88 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$27 \$88 \$135 \$17 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$28 \$90 \$142 \$89 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$29 DVDD \$140 \$90 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$30 \$90 \$139 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$31 \$53 \$89 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$32 DVDD \$89 \$53 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$33 \$52 \$89 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$34 DVDD \$89 \$52 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$35 \$55 \$92 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$36 DVDD \$92 \$55 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$37 \$54 \$92 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$38 DVDD \$92 \$54 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$39 DVDD \$139 \$91 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$40 \$91 \$144 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$41 \$92 \$146 \$91 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$42 \$18 \$135 \$19 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$43 \$19 \$135 \$18 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$44 DVDD \$91 \$19 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$45 \$19 \$91 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$46 \$251 \$215 \$266 \$266 pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$47 \$266 \$216 \$251 \$266 pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$48 \$82 DVSS \$20 DVDD pfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P PS=3.28U
+ PD=3.28U
M$49 DVDD \$251 \$138 DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$50 \$136 \$138 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$51 DVDD \$140 \$142 DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$52 \$140 \$253 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$53 \$253 \$216 \$266 \$266 pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$54 \$266 \$217 \$253 \$266 pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$55 \$256 \$266 \$266 \$266 pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$56 \$266 \$216 \$256 \$266 pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$57 \$15 DVSS \$16 DVDD pfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P PS=3.28U
+ PD=3.28U
M$58 DVDD \$256 \$144 DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$59 \$146 \$144 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$60 \$88 DVSS \$17 DVDD pfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P PS=3.28U
+ PD=3.28U
M$61 DVDD \$257 \$139 DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$62 \$257 \$258 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$63 \$258 Y \$266 \$266 pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$64 \$266 \$216 \$258 \$266 pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$65 \$395 \$401 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$66 \$260 \$280 \$266 \$266 pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$67 \$359 \$371 \$266 \$266 pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$68 \$266 \$397 \$359 \$266 pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$69 A \$451 \$266 \$266 pfet_06v0 L=0.7U W=3.5U AS=1.54P AD=0.91P PS=7.88U
+ PD=4.02U
M$70 \$266 \$451 A \$266 pfet_06v0 L=0.7U W=3.5U AS=0.91P AD=0.91P PS=4.02U
+ PD=4.02U
M$71 A \$451 \$266 \$266 pfet_06v0 L=0.7U W=3.5U AS=0.91P AD=0.91P PS=4.02U
+ PD=4.02U
M$72 \$266 \$451 A \$266 pfet_06v0 L=0.7U W=3.5U AS=0.91P AD=0.91P PS=4.02U
+ PD=4.02U
M$73 A \$451 \$266 \$266 pfet_06v0 L=0.7U W=3.5U AS=0.91P AD=0.91P PS=4.02U
+ PD=4.02U
M$74 \$266 \$451 A \$266 pfet_06v0 L=0.7U W=3.5U AS=0.91P AD=1.54P PS=4.02U
+ PD=7.88U
M$75 \$396 \$371 \$266 \$266 pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$76 \$135 \$260 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$77 DVDD \$260 \$135 DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$78 \$175 \$135 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$79 DVDD \$135 \$175 DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$80 \$397 \$396 \$393 \$266 pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$81 \$361 \$397 \$266 \$266 pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$82 \$266 \$372 \$361 \$266 pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$83 \$372 \$371 \$397 \$266 pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$84 \$18 DVSS \$19 DVDD pfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P PS=3.28U
+ PD=3.28U
M$85 \$266 \$372 \$393 \$266 pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$86 \$448 \$458 DVDD DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.52P PS=4.88U
+ PD=2.52U
M$87 DVDD \$458 \$448 DVDD pfet_06v0 L=0.7U W=2U AS=0.52P AD=0.52P PS=2.52U
+ PD=2.52U
M$88 \$448 \$458 DVDD DVDD pfet_06v0 L=0.7U W=2U AS=0.52P AD=0.88P PS=2.52U
+ PD=4.88U
M$89 \$448 \$347 \$446 DVDD pfet_06v0 L=0.7U W=2.15U AS=0.946P AD=0.559P
+ PS=5.18U PD=2.67U
M$90 \$446 \$347 \$448 DVDD pfet_06v0 L=0.7U W=2.15U AS=0.559P AD=0.946P
+ PS=2.67U PD=5.18U
M$91 \$449 \$448 DVDD DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$92 \$456 \$457 DVDD DVDD pfet_06v0 L=0.7U W=4U AS=1.76P AD=1.04P PS=8.88U
+ PD=4.52U
M$93 DVDD \$457 \$456 DVDD pfet_06v0 L=0.7U W=4U AS=1.04P AD=1.76P PS=4.52U
+ PD=8.88U
M$94 \$459 \$457 DVDD DVDD pfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.39P PS=3.88U
+ PD=2.02U
M$95 DVDD \$457 \$459 DVDD pfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.66P PS=2.02U
+ PD=3.88U
M$96 DVDD \$347 \$446 DVDD pfet_06v0 L=0.7U W=1.9U AS=0.836P AD=0.494P PS=4.68U
+ PD=2.42U
M$97 \$446 \$347 DVDD DVDD pfet_06v0 L=0.7U W=1.9U AS=0.494P AD=0.836P PS=2.42U
+ PD=4.68U
M$98 DVSS \$459 \$446 DVDD pfet_06v0 L=0.7U W=1.9U AS=0.836P AD=0.494P PS=4.68U
+ PD=2.42U
M$99 \$446 \$459 DVSS DVDD pfet_06v0 L=0.7U W=1.9U AS=0.494P AD=0.836P PS=2.42U
+ PD=4.68U
M$100 \$448 \$456 \$459 DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$101 \$450 \$456 \$448 DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$102 \$451 \$449 \$266 \$266 pfet_06v0 L=0.7U W=2.5U AS=1.1P AD=0.65P PS=5.88U
+ PD=3.02U
M$103 \$266 \$449 \$451 \$266 pfet_06v0 L=0.7U W=2.5U AS=0.65P AD=0.65P
+ PS=3.02U PD=3.02U
M$104 \$451 \$449 \$266 \$266 pfet_06v0 L=0.7U W=2.5U AS=0.65P AD=0.65P
+ PS=3.02U PD=3.02U
M$105 \$266 \$449 \$451 \$266 pfet_06v0 L=0.7U W=2.5U AS=0.65P AD=1.1P PS=3.02U
+ PD=5.88U
M$106 \$528 \$553 \$266 \$266 pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$107 \$458 \$528 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$108 DVDD \$528 \$458 DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$109 \$529 \$458 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$110 DVDD \$458 \$529 DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$111 \$530 \$457 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$112 DVDD \$457 \$530 DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$113 \$457 \$531 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$114 DVDD \$531 \$457 DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$115 \$266 \$518 \$531 \$266 pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$116 \$532 \$359 \$266 \$266 pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$117 \$533 \$532 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$118 DVDD \$532 \$533 DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$119 \$414 \$533 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$120 DVDD \$533 \$414 DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$121 \$534 \$401 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$122 DVDD \$401 \$534 DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$123 \$401 \$535 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$124 DVDD \$535 \$401 DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$125 \$266 \$361 \$535 \$266 pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$126 Y A DVSS DVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$127 \$49 DVDD \$85 DVSS nfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P PS=3.28U
+ PD=3.28U
M$128 \$50 DVDD \$51 DVSS nfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P PS=3.28U
+ PD=3.28U
M$129 \$52 DVDD \$53 DVSS nfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P PS=3.28U
+ PD=3.28U
M$130 \$54 DVDD \$55 DVSS nfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P PS=3.28U
+ PD=3.28U
M$131 \$20 \$84 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$132 DVSS \$84 \$20 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$133 \$82 \$84 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$134 DVSS \$84 \$82 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$135 \$83 \$136 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$136 \$84 \$138 \$83 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$137 DVSS \$139 \$83 DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$138 \$85 \$83 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$139 DVSS \$83 \$85 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$140 \$85 \$175 \$49 DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$141 \$49 \$175 \$85 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$142 \$50 \$175 \$51 DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$143 \$51 \$175 \$50 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$144 \$50 \$87 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$145 DVSS \$87 \$50 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$146 \$87 \$139 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$147 \$87 \$140 \$86 DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$148 DVSS \$142 \$87 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$149 \$16 \$86 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$150 DVSS \$86 \$16 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$151 \$15 \$86 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$152 DVSS \$86 \$15 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$153 \$17 \$90 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$154 DVSS \$90 \$17 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$155 \$88 \$90 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$156 DVSS \$90 \$88 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$157 \$89 \$142 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$158 \$90 \$140 \$89 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$159 DVSS \$139 \$89 DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$160 \$53 \$89 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$161 DVSS \$89 \$53 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$162 \$53 \$175 \$52 DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$163 \$52 \$175 \$53 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$164 \$54 \$175 \$55 DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$165 \$55 \$175 \$54 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$166 \$54 \$92 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$167 DVSS \$92 \$54 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$168 \$92 \$139 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$169 \$92 \$144 \$91 DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$170 DVSS \$146 \$92 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$171 \$19 \$91 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$172 DVSS \$91 \$19 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$173 \$18 \$91 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$174 DVSS \$91 \$18 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$175 \$250 \$215 \$5 DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$176 \$251 \$216 \$250 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$177 DVSS \$251 \$138 DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$178 \$136 \$138 DVSS DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$179 DVSS \$456 \$450 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$180 DVSS \$140 \$142 DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$181 \$140 \$253 DVSS DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$182 \$480 \$458 DVSS DVSS nfet_06v0 L=0.7U W=3.2U AS=1.408P AD=0.832P
+ PS=7.28U PD=3.72U
M$183 DVSS \$458 \$480 DVSS nfet_06v0 L=0.7U W=3.2U AS=0.832P AD=0.832P
+ PS=3.72U PD=3.72U
M$184 \$480 \$458 DVSS DVSS nfet_06v0 L=0.7U W=3.2U AS=0.832P AD=0.832P
+ PS=3.72U PD=3.72U
M$185 DVSS \$458 \$480 DVSS nfet_06v0 L=0.7U W=3.2U AS=0.832P AD=0.832P
+ PS=3.72U PD=3.72U
M$186 \$480 \$458 DVSS DVSS nfet_06v0 L=0.7U W=3.2U AS=0.832P AD=1.408P
+ PS=3.72U PD=7.28U
M$187 \$254 \$216 \$253 DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$188 \$5 \$217 \$254 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$189 \$255 \$266 \$5 DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$190 \$256 \$216 \$255 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$191 DVSS \$256 \$144 DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$192 \$146 \$144 DVSS DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$193 \$448 \$457 \$459 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$194 \$450 \$457 \$448 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$195 DVSS \$257 \$139 DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$196 \$257 \$258 DVSS DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$197 DVSS \$448 \$449 DVSS nfet_06v0 L=0.7U W=4U AS=1.76P AD=1.04P PS=8.88U
+ PD=4.52U
M$198 \$449 \$448 DVSS DVSS nfet_06v0 L=0.7U W=4U AS=1.04P AD=1.76P PS=4.52U
+ PD=8.88U
M$199 \$259 Y \$258 DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$200 \$5 \$216 \$259 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$201 \$395 \$414 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$202 \$260 \$280 \$5 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$203 \$360 \$371 \$359 DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$204 \$5 \$397 \$360 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$205 \$396 \$371 \$5 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$206 \$135 \$260 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.39P PS=3.88U
+ PD=2.02U
M$207 DVSS \$260 \$135 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$208 \$175 \$135 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$209 DVSS \$135 \$175 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.66P PS=2.02U
+ PD=3.88U
M$210 \$397 \$371 \$393 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$211 \$362 \$397 \$361 DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$212 \$5 \$372 \$362 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$213 \$372 \$396 \$397 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$214 \$5 \$372 \$393 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$215 \$456 \$457 DVSS DVSS nfet_06v0 L=0.7U W=2U AS=0.88P AD=0.52P PS=4.88U
+ PD=2.52U
M$216 DVSS \$457 \$456 DVSS nfet_06v0 L=0.7U W=2U AS=0.52P AD=0.88P PS=2.52U
+ PD=4.88U
M$217 \$480 \$347 \$483 DVSS nfet_06v0 L=0.7U W=2.65U AS=1.166P AD=0.689P
+ PS=6.18U PD=3.17U
M$218 \$483 \$347 \$480 DVSS nfet_06v0 L=0.7U W=2.65U AS=0.689P AD=0.689P
+ PS=3.17U PD=3.17U
M$219 \$480 \$347 \$483 DVSS nfet_06v0 L=0.7U W=2.65U AS=0.689P AD=0.689P
+ PS=3.17U PD=3.17U
M$220 \$483 \$347 \$480 DVSS nfet_06v0 L=0.7U W=2.65U AS=0.689P AD=1.166P
+ PS=3.17U PD=6.18U
M$221 \$448 \$347 \$483 DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$222 \$483 \$347 \$448 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$223 \$448 \$347 \$483 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$224 \$483 \$347 \$448 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$225 \$483 \$450 DVDD DVSS nfet_06v0 L=0.7U W=1.3U AS=0.572P AD=0.572P
+ PS=3.48U PD=3.48U
M$226 \$528 \$553 \$5 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$227 \$458 \$528 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.39P PS=3.88U
+ PD=2.02U
M$228 DVSS \$528 \$458 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$229 \$529 \$458 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$230 DVSS \$458 \$529 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.66P PS=2.02U
+ PD=3.88U
M$231 \$530 \$457 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.39P PS=3.88U
+ PD=2.02U
M$232 DVSS \$457 \$530 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$233 \$457 \$531 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$234 DVSS \$531 \$457 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.66P PS=2.02U
+ PD=3.88U
M$235 \$5 \$518 \$531 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$236 \$532 \$359 \$5 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$237 \$533 \$532 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.39P PS=3.88U
+ PD=2.02U
M$238 DVSS \$532 \$533 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$239 \$414 \$533 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$240 DVSS \$533 \$414 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.66P PS=2.02U
+ PD=3.88U
M$241 \$451 \$449 \$5 DVSS nfet_06v0 L=0.7U W=1.25U AS=0.55P AD=0.325P PS=3.38U
+ PD=1.77U
M$242 \$5 \$449 \$451 DVSS nfet_06v0 L=0.7U W=1.25U AS=0.325P AD=0.55P PS=1.77U
+ PD=3.38U
M$243 \$534 \$401 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.39P PS=3.88U
+ PD=2.02U
M$244 DVSS \$401 \$534 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$245 \$401 \$535 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$246 DVSS \$535 \$401 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.66P PS=2.02U
+ PD=3.88U
M$247 A \$451 \$5 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.39P PS=3.88U
+ PD=2.02U
M$248 \$5 \$451 A DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$249 A \$451 \$5 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$250 \$5 \$451 A DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$251 A \$451 \$5 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$252 \$5 \$451 A DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.66P PS=2.02U
+ PD=3.88U
M$253 \$5 \$361 \$535 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
D$254 \$5 \$215 diode_pd2nw_06v0 A=0.2304P P=1.92U
D$255 \$5 \$216 diode_pd2nw_06v0 A=0.2304P P=1.92U
D$256 \$5 \$216 diode_pd2nw_06v0 A=0.2304P P=1.92U
D$257 \$5 \$217 diode_pd2nw_06v0 A=0.2304P P=1.92U
D$258 \$5 \$266 diode_pd2nw_06v0 A=0.2304P P=1.92U
D$259 \$5 \$216 diode_pd2nw_06v0 A=0.2304P P=1.92U
D$260 Y \$266 diode_pd2nw_06v0 A=1P P=4U
D$261 \$280 \$266 diode_pd2nw_06v0 A=1P P=4U
D$262 \$372 \$266 diode_pd2nw_06v0 A=1P P=4U
D$263 \$371 \$266 diode_pd2nw_06v0 A=1P P=4U
D$264 \$518 \$266 diode_pd2nw_06v0 A=1P P=4U
D$265 \$553 \$266 diode_pd2nw_06v0 A=1P P=4U
R$266 \$332 \$395 DVSS 15618.75 ppolyf_u L=35.7U W=0.8U
R$267 \$332 \$416 DVSS 15618.75 ppolyf_u L=35.7U W=0.8U
R$268 \$333 \$416 DVSS 15618.75 ppolyf_u L=35.7U W=0.8U
R$269 \$333 \$417 DVSS 15618.75 ppolyf_u L=35.7U W=0.8U
R$270 \$334 \$417 DVSS 15618.75 ppolyf_u L=35.7U W=0.8U
R$271 \$334 \$418 DVSS 15618.75 ppolyf_u L=35.7U W=0.8U
R$272 \$335 \$418 DVSS 15618.75 ppolyf_u L=35.7U W=0.8U
R$273 \$335 \$347 DVSS 10062.5 ppolyf_u L=23U W=0.8U
R$274 \$1 \$347 DVSS 392 ppolyf_u L=2.8U W=2.5U
R$275 \$1 \$347 DVSS 392 ppolyf_u L=2.8U W=2.5U
R$276 \$1 \$347 DVSS 392 ppolyf_u L=2.8U W=2.5U
R$277 \$1 \$347 DVSS 392 ppolyf_u L=2.8U W=2.5U
C$278 DVDD DVSS 2.07e-14 cap_nmos_06v0 A=9P P=12U
C$279 DVDD DVSS 2.07e-14 cap_nmos_06v0 A=9P P=12U
C$280 DVDD DVSS 2.07e-14 cap_nmos_06v0 A=9P P=12U
C$281 DVDD DVSS 2.07e-14 cap_nmos_06v0 A=9P P=12U
C$282 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$283 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$284 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$285 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$286 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$287 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$288 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$289 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$290 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$291 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
M$292 \$1 \$49 DVDD DVDD pfet_06v0_dss L=0.7U W=40U AS=31.6P AD=124.4P
+ PS=81.58U PD=46.22U
M$293 DVDD \$49 \$1 DVDD pfet_06v0_dss L=0.7U W=40U AS=124.4P AD=24.4P
+ PS=46.22U PD=41.22U
M$294 \$1 \$85 DVDD DVDD pfet_06v0_dss L=0.7U W=40U AS=24.4P AD=124.4P
+ PS=41.22U PD=46.22U
M$295 DVDD \$50 \$1 DVDD pfet_06v0_dss L=0.7U W=40U AS=124.4P AD=24.4P
+ PS=46.22U PD=41.22U
M$296 \$1 \$51 DVDD DVDD pfet_06v0_dss L=0.7U W=40U AS=24.4P AD=124.4P
+ PS=41.22U PD=46.22U
M$297 DVDD \$51 \$1 DVDD pfet_06v0_dss L=0.7U W=40U AS=124.4P AD=24.4P
+ PS=46.22U PD=41.22U
M$298 \$1 \$52 DVDD DVDD pfet_06v0_dss L=0.7U W=40U AS=24.4P AD=124.4P
+ PS=41.22U PD=46.22U
M$299 DVDD \$52 \$1 DVDD pfet_06v0_dss L=0.7U W=40U AS=124.4P AD=24.4P
+ PS=46.22U PD=41.22U
M$300 \$1 \$53 DVDD DVDD pfet_06v0_dss L=0.7U W=40U AS=24.4P AD=124.4P
+ PS=41.22U PD=46.22U
M$301 DVDD \$54 \$1 DVDD pfet_06v0_dss L=0.7U W=40U AS=124.4P AD=24.4P
+ PS=46.22U PD=41.22U
M$302 \$1 \$55 DVDD DVDD pfet_06v0_dss L=0.7U W=40U AS=24.4P AD=124.4P
+ PS=41.22U PD=46.22U
M$303 DVDD \$55 \$1 DVDD pfet_06v0_dss L=0.7U W=40U AS=124.4P AD=31.6P
+ PS=46.22U PD=81.58U
M$304 \$1 \$20 DVSS DVSS nfet_06v0_dss L=1.15U W=38U AS=30.02P AD=156.18P
+ PS=77.58U PD=46.22U
M$305 DVSS \$82 \$1 DVSS nfet_06v0_dss L=1.15U W=38U AS=156.18P AD=23.18P
+ PS=46.22U PD=39.22U
M$306 \$1 \$15 DVSS DVSS nfet_06v0_dss L=1.15U W=38U AS=23.18P AD=156.18P
+ PS=39.22U PD=46.22U
M$307 DVSS \$16 \$1 DVSS nfet_06v0_dss L=1.15U W=38U AS=156.18P AD=23.18P
+ PS=46.22U PD=39.22U
M$308 \$1 \$17 DVSS DVSS nfet_06v0_dss L=1.15U W=38U AS=23.18P AD=156.18P
+ PS=39.22U PD=46.22U
M$309 DVSS \$88 \$1 DVSS nfet_06v0_dss L=1.15U W=38U AS=156.18P AD=23.18P
+ PS=46.22U PD=39.22U
M$310 \$1 \$18 DVSS DVSS nfet_06v0_dss L=1.15U W=38U AS=23.18P AD=156.18P
+ PS=39.22U PD=46.22U
M$311 DVSS \$19 \$1 DVSS nfet_06v0_dss L=1.15U W=38U AS=156.18P AD=30.02P
+ PS=46.22U PD=77.58U
.ENDS inverter_PAD
