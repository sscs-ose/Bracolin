* Extracted by KLayout with GF180MCU LVS runset on : 16/03/2024 13:19

.SUBCKT inverter_PAD VSS DVDD DVSS NDRIVE_X NDRIVE_Y PDRIVE_X PDRIVE_Y Z ENB EN
+ A|AB ZB PDRV OE PDRV|VDD A A|PDB_OUT|Z A|PUB_OUT|Z B A|B PU_B|Z PD|ZB A|Z
M$1 A \$656 DVDD DVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2 DVDD \$91 NDRIVE_Y DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$3 NDRIVE_Y \$91 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$4 NDRIVE_X Z NDRIVE_Y DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$5 NDRIVE_Y Z NDRIVE_X DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$6 \$91 ENB \$90 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$7 DVDD EN \$91 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$8 \$91 A|AB DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$9 PDRIVE_Y \$90 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$10 DVDD \$90 PDRIVE_Y DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$11 PDRIVE_X \$90 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$12 DVDD \$90 PDRIVE_X DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$13 PDRIVE_X \$94 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$14 DVDD \$94 PDRIVE_X DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$15 PDRIVE_Y \$94 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$16 DVDD \$94 PDRIVE_Y DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$17 DVDD A|AB \$93 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$18 \$93 EN DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$19 \$94 ENB \$93 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$20 NDRIVE_X Z NDRIVE_Y DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P
+ PS=24.88U PD=12.52U
M$21 NDRIVE_Y Z NDRIVE_X DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P
+ PS=12.52U PD=12.52U
M$22 DVDD \$93 NDRIVE_Y DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$23 NDRIVE_Y \$93 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$24 DVDD \$97 NDRIVE_Y DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$25 NDRIVE_Y \$97 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$26 NDRIVE_X Z NDRIVE_Y DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P
+ PS=12.52U PD=12.52U
M$27 NDRIVE_Y Z NDRIVE_X DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P
+ PS=12.52U PD=24.88U
M$28 \$97 ENB \$96 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$29 DVDD EN \$97 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$30 \$97 A|AB DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$31 PDRIVE_Y \$96 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$32 DVDD \$96 PDRIVE_Y DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$33 PDRIVE_X \$96 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$34 DVDD \$96 PDRIVE_X DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$35 PDRIVE_X \$100 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P
+ PS=24.88U PD=12.52U
M$36 DVDD \$100 PDRIVE_X DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P
+ PS=12.52U PD=12.52U
M$37 PDRIVE_Y \$100 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P
+ PS=12.52U PD=12.52U
M$38 DVDD \$100 PDRIVE_Y DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P
+ PS=12.52U PD=24.88U
M$39 DVDD A|AB \$99 DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P PS=24.88U
+ PD=12.52U
M$40 \$99 EN DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$41 \$100 ENB \$99 DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$42 NDRIVE_X Z NDRIVE_Y DVDD pfet_06v0 L=0.7U W=12U AS=5.28P AD=3.12P
+ PS=24.88U PD=12.52U
M$43 NDRIVE_Y Z NDRIVE_X DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P
+ PS=12.52U PD=12.52U
M$44 DVDD \$99 NDRIVE_Y DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=3.12P PS=12.52U
+ PD=12.52U
M$45 NDRIVE_Y \$99 DVDD DVDD pfet_06v0 L=0.7U W=12U AS=3.12P AD=5.28P PS=12.52U
+ PD=24.88U
M$46 \$251 PDRV PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$47 PDRV|VDD OE \$251 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$48 NDRIVE_Y DVSS NDRIVE_X DVDD pfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P
+ PS=3.28U PD=3.28U
M$49 DVDD \$251 EN DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$50 ENB EN DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U PD=12.88U
M$51 DVDD EN ENB DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U PD=6.52U
M$52 EN \$253 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$53 \$253 OE PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$54 PDRV|VDD PDRV \$253 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$55 \$256 PDRV|VDD PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$56 PDRV|VDD OE \$256 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$57 NDRIVE_X DVSS NDRIVE_Y DVDD pfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P
+ PS=3.28U PD=3.28U
M$58 DVDD \$256 EN DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$59 ENB EN DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U PD=12.88U
M$60 NDRIVE_Y DVSS NDRIVE_X DVDD pfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P
+ PS=3.28U PD=3.28U
M$61 DVDD \$257 A|AB DVDD pfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$62 \$257 \$258 DVDD DVDD pfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$63 \$258 A PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$64 PDRV|VDD OE \$258 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$65 \$396 PU_B|Z DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$66 \$260 A PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$67 A|PDB_OUT|Z B PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$68 PDRV|VDD A|B A|PDB_OUT|Z PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$69 \$447 Z PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3.5U AS=1.54P AD=0.91P
+ PS=7.88U PD=4.02U
M$70 PDRV|VDD Z \$447 PDRV|VDD pfet_06v0 L=0.7U W=3.5U AS=0.91P AD=0.91P
+ PS=4.02U PD=4.02U
M$71 \$447 Z PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3.5U AS=0.91P AD=0.91P
+ PS=4.02U PD=4.02U
M$72 PDRV|VDD Z \$447 PDRV|VDD pfet_06v0 L=0.7U W=3.5U AS=0.91P AD=0.91P
+ PS=4.02U PD=4.02U
M$73 \$447 Z PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3.5U AS=0.91P AD=0.91P
+ PS=4.02U PD=4.02U
M$74 PDRV|VDD Z \$447 PDRV|VDD pfet_06v0 L=0.7U W=3.5U AS=0.91P AD=1.54P
+ PS=4.02U PD=7.88U
M$75 \$397 B PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$76 Z \$260 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U PD=3.52U
M$77 DVDD \$260 Z DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U PD=3.52U
M$78 ZB Z DVDD DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U PD=3.52U
M$79 DVDD Z ZB DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U PD=6.88U
M$80 A|B \$397 \$394 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$81 A|PUB_OUT|Z A|B PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$82 PDRV|VDD A A|PUB_OUT|Z PDRV|VDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P
+ PS=3.52U PD=6.88U
M$83 A B A|B PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U PD=6.88U
M$84 NDRIVE_X DVSS NDRIVE_Y DVDD pfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P
+ PS=3.28U PD=3.28U
M$85 PDRV|VDD A \$394 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P PS=6.88U
+ PD=6.88U
M$86 A|Z Z DVDD DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.52P PS=4.88U PD=2.52U
M$87 DVDD Z A|Z DVDD pfet_06v0 L=0.7U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$88 A|Z Z DVDD DVDD pfet_06v0 L=0.7U W=2U AS=0.52P AD=0.88P PS=2.52U PD=4.88U
M$89 A|Z A \$446 DVDD pfet_06v0 L=0.7U W=2.15U AS=0.946P AD=0.559P PS=5.18U
+ PD=2.67U
M$90 \$446 A A|Z DVDD pfet_06v0 L=0.7U W=2.15U AS=0.559P AD=0.946P PS=2.67U
+ PD=5.18U
M$91 \$449 A|Z DVDD DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$92 \$456 Z DVDD DVDD pfet_06v0 L=0.7U W=4U AS=1.76P AD=1.04P PS=8.88U PD=4.52U
M$93 DVDD Z \$456 DVDD pfet_06v0 L=0.7U W=4U AS=1.04P AD=1.76P PS=4.52U PD=8.88U
M$94 \$459 Z DVDD DVDD pfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.39P PS=3.88U
+ PD=2.02U
M$95 DVDD Z \$459 DVDD pfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.66P PS=2.02U
+ PD=3.88U
M$96 DVDD A \$446 DVDD pfet_06v0 L=0.7U W=1.9U AS=0.836P AD=0.494P PS=4.68U
+ PD=2.42U
M$97 \$446 A DVDD DVDD pfet_06v0 L=0.7U W=1.9U AS=0.494P AD=0.836P PS=2.42U
+ PD=4.68U
M$98 DVSS \$459 \$446 DVDD pfet_06v0 L=0.7U W=1.9U AS=0.836P AD=0.494P PS=4.68U
+ PD=2.42U
M$99 \$446 \$459 DVSS DVDD pfet_06v0 L=0.7U W=1.9U AS=0.494P AD=0.836P PS=2.42U
+ PD=4.68U
M$100 A|Z \$456 \$459 DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$101 \$450 \$456 A|Z DVDD pfet_06v0 L=0.7U W=2U AS=0.88P AD=0.88P PS=4.88U
+ PD=4.88U
M$102 Z \$449 PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=2.5U AS=1.1P AD=0.65P
+ PS=5.88U PD=3.02U
M$103 PDRV|VDD \$449 Z PDRV|VDD pfet_06v0 L=0.7U W=2.5U AS=0.65P AD=0.65P
+ PS=3.02U PD=3.02U
M$104 Z \$449 PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=2.5U AS=0.65P AD=0.65P
+ PS=3.02U PD=3.02U
M$105 PDRV|VDD \$449 Z PDRV|VDD pfet_06v0 L=0.7U W=2.5U AS=0.65P AD=1.1P
+ PS=3.02U PD=5.88U
M$106 \$528 A PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$107 Z \$528 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$108 DVDD \$528 Z DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$109 ZB Z DVDD DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U PD=3.52U
M$110 DVDD Z ZB DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U PD=6.88U
M$111 ZB Z DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U PD=3.52U
M$112 DVDD Z ZB DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U PD=3.52U
M$113 Z \$531 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$114 DVDD \$531 Z DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$115 PDRV|VDD A \$531 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=1.32P
+ PS=6.88U PD=6.88U
M$116 \$532 A|PDB_OUT|Z PDRV|VDD PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$117 Z \$532 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$118 DVDD \$532 Z DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$119 PD|ZB Z DVDD DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$120 DVDD Z PD|ZB DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$121 ZB PU_B|Z DVDD DVDD pfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$122 DVDD PU_B|Z ZB DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$123 PU_B|Z \$535 DVDD DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U
+ PD=3.52U
M$124 DVDD \$535 PU_B|Z DVDD pfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$125 PDRV|VDD A|PUB_OUT|Z \$535 PDRV|VDD pfet_06v0 L=0.7U W=3U AS=1.32P
+ AD=1.32P PS=6.88U PD=6.88U
M$126 A \$656 DVSS DVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$127 PDRIVE_X DVDD PDRIVE_Y DVSS nfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P
+ PS=3.28U PD=3.28U
M$128 PDRIVE_Y DVDD PDRIVE_X DVSS nfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P
+ PS=3.28U PD=3.28U
M$129 PDRIVE_X DVDD PDRIVE_Y DVSS nfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P
+ PS=3.28U PD=3.28U
M$130 PDRIVE_Y DVDD PDRIVE_X DVSS nfet_06v0 L=0.7U W=1.2U AS=0.528P AD=0.528P
+ PS=3.28U PD=3.28U
M$131 NDRIVE_X \$91 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$132 DVSS \$91 NDRIVE_X DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$133 NDRIVE_Y \$91 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$134 DVSS \$91 NDRIVE_Y DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$135 \$90 ENB DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$136 \$91 EN \$90 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$137 DVSS A|AB \$90 DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$138 PDRIVE_Y \$90 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$139 DVSS \$90 PDRIVE_Y DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$140 PDRIVE_Y ZB PDRIVE_X DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P
+ PS=12.88U PD=6.52U
M$141 PDRIVE_X ZB PDRIVE_Y DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P
+ PS=6.52U PD=12.88U
M$142 PDRIVE_Y ZB PDRIVE_X DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P
+ PS=12.88U PD=6.52U
M$143 PDRIVE_X ZB PDRIVE_Y DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P
+ PS=6.52U PD=12.88U
M$144 PDRIVE_Y \$94 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$145 DVSS \$94 PDRIVE_Y DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$146 \$94 A|AB DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$147 \$94 EN \$93 DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$148 DVSS ENB \$94 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$149 NDRIVE_Y \$93 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$150 DVSS \$93 NDRIVE_Y DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$151 NDRIVE_X \$93 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$152 DVSS \$93 NDRIVE_X DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$153 NDRIVE_X \$97 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$154 DVSS \$97 NDRIVE_X DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$155 NDRIVE_Y \$97 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$156 DVSS \$97 NDRIVE_Y DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$157 \$96 ENB DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$158 \$97 EN \$96 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$159 DVSS A|AB \$96 DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$160 PDRIVE_Y \$96 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$161 DVSS \$96 PDRIVE_Y DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$162 PDRIVE_Y ZB PDRIVE_X DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P
+ PS=12.88U PD=6.52U
M$163 PDRIVE_X ZB PDRIVE_Y DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P
+ PS=6.52U PD=12.88U
M$164 PDRIVE_Y ZB PDRIVE_X DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P
+ PS=12.88U PD=6.52U
M$165 PDRIVE_X ZB PDRIVE_Y DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P
+ PS=6.52U PD=12.88U
M$166 PDRIVE_Y \$100 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P
+ PS=12.88U PD=6.52U
M$167 DVSS \$100 PDRIVE_Y DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$168 \$100 A|AB DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$169 \$100 EN \$99 DVSS nfet_06v0 L=0.7U W=6U AS=2.64P AD=1.56P PS=12.88U
+ PD=6.52U
M$170 DVSS ENB \$100 DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$171 NDRIVE_Y \$99 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$172 DVSS \$99 NDRIVE_Y DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$173 NDRIVE_X \$99 DVSS DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=1.56P PS=6.52U
+ PD=6.52U
M$174 DVSS \$99 NDRIVE_X DVSS nfet_06v0 L=0.7U W=6U AS=1.56P AD=2.64P PS=6.52U
+ PD=12.88U
M$175 \$250 PDRV VSS DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$176 \$251 OE \$250 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$177 DVSS \$251 EN DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$178 ENB EN DVSS DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U PD=6.88U
M$179 DVSS \$456 \$450 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$180 DVSS EN ENB DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U PD=3.52U
M$181 EN \$253 DVSS DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$182 \$481 Z DVSS DVSS nfet_06v0 L=0.7U W=3.2U AS=1.408P AD=0.832P PS=7.28U
+ PD=3.72U
M$183 DVSS Z \$481 DVSS nfet_06v0 L=0.7U W=3.2U AS=0.832P AD=0.832P PS=3.72U
+ PD=3.72U
M$184 \$481 Z DVSS DVSS nfet_06v0 L=0.7U W=3.2U AS=0.832P AD=0.832P PS=3.72U
+ PD=3.72U
M$185 DVSS Z \$481 DVSS nfet_06v0 L=0.7U W=3.2U AS=0.832P AD=0.832P PS=3.72U
+ PD=3.72U
M$186 \$481 Z DVSS DVSS nfet_06v0 L=0.7U W=3.2U AS=0.832P AD=1.408P PS=3.72U
+ PD=7.28U
M$187 \$254 OE \$253 DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$188 VSS PDRV \$254 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$189 \$255 PDRV|VDD VSS DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$190 \$256 OE \$255 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$191 DVSS \$256 EN DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$192 ENB EN DVSS DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U PD=6.88U
M$193 A|Z Z \$459 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$194 \$450 Z A|Z DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$195 DVSS \$257 A|AB DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$196 \$257 \$258 DVSS DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$197 DVSS A|Z \$449 DVSS nfet_06v0 L=0.7U W=4U AS=1.76P AD=1.04P PS=8.88U
+ PD=4.52U
M$198 \$449 A|Z DVSS DVSS nfet_06v0 L=0.7U W=4U AS=1.04P AD=1.76P PS=4.52U
+ PD=8.88U
M$199 \$259 A \$258 DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$200 VSS OE \$259 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$201 \$396 PD|ZB DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$202 \$260 A VSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$203 \$361 B A|PDB_OUT|Z DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U
+ PD=3.52U
M$204 VSS A|B \$361 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U
+ PD=6.88U
M$205 \$397 B VSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$206 Z \$260 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.39P PS=3.88U
+ PD=2.02U
M$207 DVSS \$260 Z DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$208 ZB Z DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U PD=2.02U
M$209 DVSS Z ZB DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.66P PS=2.02U PD=3.88U
M$210 A|B B \$394 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$211 \$363 A|B A|PUB_OUT|Z DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P
+ PS=6.88U PD=3.52U
M$212 VSS A \$363 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U PD=6.88U
M$213 A \$397 A|B DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$214 VSS A \$394 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$215 \$456 Z DVSS DVSS nfet_06v0 L=0.7U W=2U AS=0.88P AD=0.52P PS=4.88U
+ PD=2.52U
M$216 DVSS Z \$456 DVSS nfet_06v0 L=0.7U W=2U AS=0.52P AD=0.88P PS=2.52U
+ PD=4.88U
M$217 \$481 A \$483 DVSS nfet_06v0 L=0.7U W=2.65U AS=1.166P AD=0.689P PS=6.18U
+ PD=3.17U
M$218 \$483 A \$481 DVSS nfet_06v0 L=0.7U W=2.65U AS=0.689P AD=0.689P PS=3.17U
+ PD=3.17U
M$219 \$481 A \$483 DVSS nfet_06v0 L=0.7U W=2.65U AS=0.689P AD=0.689P PS=3.17U
+ PD=3.17U
M$220 \$483 A \$481 DVSS nfet_06v0 L=0.7U W=2.65U AS=0.689P AD=1.166P PS=3.17U
+ PD=6.18U
M$221 A|Z A \$483 DVSS nfet_06v0 L=0.7U W=3U AS=1.32P AD=0.78P PS=6.88U PD=3.52U
M$222 \$483 A A|Z DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U PD=3.52U
M$223 A|Z A \$483 DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=0.78P PS=3.52U PD=3.52U
M$224 \$483 A A|Z DVSS nfet_06v0 L=0.7U W=3U AS=0.78P AD=1.32P PS=3.52U PD=6.88U
M$225 \$483 \$450 DVDD DVSS nfet_06v0 L=0.7U W=1.3U AS=0.572P AD=0.572P
+ PS=3.48U PD=3.48U
M$226 \$528 A VSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$227 Z \$528 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.39P PS=3.88U
+ PD=2.02U
M$228 DVSS \$528 Z DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$229 ZB Z DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U PD=2.02U
M$230 DVSS Z ZB DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.66P PS=2.02U PD=3.88U
M$231 ZB Z DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.39P PS=3.88U PD=2.02U
M$232 DVSS Z ZB DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U PD=2.02U
M$233 Z \$531 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$234 DVSS \$531 Z DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.66P PS=2.02U
+ PD=3.88U
M$235 VSS A \$531 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P PS=3.88U
+ PD=3.88U
M$236 \$532 A|PDB_OUT|Z VSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
M$237 Z \$532 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.39P PS=3.88U
+ PD=2.02U
M$238 DVSS \$532 Z DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$239 PD|ZB Z DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$240 DVSS Z PD|ZB DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.66P PS=2.02U
+ PD=3.88U
M$241 Z \$449 VSS DVSS nfet_06v0 L=0.7U W=1.25U AS=0.55P AD=0.325P PS=3.38U
+ PD=1.77U
M$242 VSS \$449 Z DVSS nfet_06v0 L=0.7U W=1.25U AS=0.325P AD=0.55P PS=1.77U
+ PD=3.38U
M$243 ZB PU_B|Z DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.39P PS=3.88U
+ PD=2.02U
M$244 DVSS PU_B|Z ZB DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$245 PU_B|Z \$535 DVSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$246 DVSS \$535 PU_B|Z DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.66P PS=2.02U
+ PD=3.88U
M$247 \$447 Z VSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.39P PS=3.88U
+ PD=2.02U
M$248 VSS Z \$447 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$249 \$447 Z VSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$250 VSS Z \$447 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$251 \$447 Z VSS DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.39P PS=2.02U
+ PD=2.02U
M$252 VSS Z \$447 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.39P AD=0.66P PS=2.02U
+ PD=3.88U
M$253 VSS A|PUB_OUT|Z \$535 DVSS nfet_06v0 L=0.7U W=1.5U AS=0.66P AD=0.66P
+ PS=3.88U PD=3.88U
D$254 VSS PDRV diode_pd2nw_06v0 A=0.2304P P=1.92U
D$255 VSS OE diode_pd2nw_06v0 A=0.2304P P=1.92U
D$256 VSS OE diode_pd2nw_06v0 A=0.2304P P=1.92U
D$257 VSS PDRV diode_pd2nw_06v0 A=0.2304P P=1.92U
D$258 VSS PDRV|VDD diode_pd2nw_06v0 A=0.2304P P=1.92U
D$259 VSS OE diode_pd2nw_06v0 A=0.2304P P=1.92U
D$260 A PDRV|VDD diode_pd2nw_06v0 A=1P P=4U
D$261 A PDRV|VDD diode_pd2nw_06v0 A=1P P=4U
D$262 A PDRV|VDD diode_pd2nw_06v0 A=1P P=4U
D$263 B PDRV|VDD diode_pd2nw_06v0 A=1P P=4U
D$264 A PDRV|VDD diode_pd2nw_06v0 A=1P P=4U
D$265 A PDRV|VDD diode_pd2nw_06v0 A=1P P=4U
R$266 \$332 \$396 DVSS 15618.75 ppolyf_u L=35.7U W=0.8U
R$267 \$332 \$416 DVSS 15618.75 ppolyf_u L=35.7U W=0.8U
R$268 \$333 \$416 DVSS 15618.75 ppolyf_u L=35.7U W=0.8U
R$269 \$333 \$417 DVSS 15618.75 ppolyf_u L=35.7U W=0.8U
R$270 \$334 \$417 DVSS 15618.75 ppolyf_u L=35.7U W=0.8U
R$271 \$334 \$418 DVSS 15618.75 ppolyf_u L=35.7U W=0.8U
R$272 \$335 \$418 DVSS 15618.75 ppolyf_u L=35.7U W=0.8U
R$273 \$335 A DVSS 10062.5 ppolyf_u L=23U W=0.8U
R$274 \$1 A DVSS 392 ppolyf_u L=2.8U W=2.5U
R$275 \$1 A DVSS 392 ppolyf_u L=2.8U W=2.5U
R$276 \$1 A DVSS 392 ppolyf_u L=2.8U W=2.5U
R$277 \$1 A DVSS 392 ppolyf_u L=2.8U W=2.5U
C$278 DVDD DVSS 2.07e-14 cap_nmos_06v0 A=9P P=12U
C$279 DVDD DVSS 2.07e-14 cap_nmos_06v0 A=9P P=12U
C$280 DVDD DVSS 2.07e-14 cap_nmos_06v0 A=9P P=12U
C$281 DVDD DVSS 2.07e-14 cap_nmos_06v0 A=9P P=12U
C$282 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$283 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$284 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$285 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$286 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$287 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$288 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$289 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$290 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
C$291 DVDD DVSS 1.725e-14 cap_nmos_06v0 A=7.5P P=13U
M$292 \$1 PDRIVE_X DVDD DVDD pfet_06v0_dss L=0.7U W=40U AS=31.6P AD=124.4P
+ PS=81.58U PD=46.22U
M$293 DVDD PDRIVE_X \$1 DVDD pfet_06v0_dss L=0.7U W=40U AS=124.4P AD=24.4P
+ PS=46.22U PD=41.22U
M$294 \$1 PDRIVE_Y DVDD DVDD pfet_06v0_dss L=0.7U W=40U AS=24.4P AD=124.4P
+ PS=41.22U PD=46.22U
M$295 DVDD PDRIVE_Y \$1 DVDD pfet_06v0_dss L=0.7U W=40U AS=124.4P AD=24.4P
+ PS=46.22U PD=41.22U
M$296 \$1 PDRIVE_X DVDD DVDD pfet_06v0_dss L=0.7U W=40U AS=24.4P AD=124.4P
+ PS=41.22U PD=46.22U
M$297 DVDD PDRIVE_X \$1 DVDD pfet_06v0_dss L=0.7U W=40U AS=124.4P AD=24.4P
+ PS=46.22U PD=41.22U
M$298 \$1 PDRIVE_X DVDD DVDD pfet_06v0_dss L=0.7U W=40U AS=24.4P AD=124.4P
+ PS=41.22U PD=46.22U
M$299 DVDD PDRIVE_X \$1 DVDD pfet_06v0_dss L=0.7U W=40U AS=124.4P AD=24.4P
+ PS=46.22U PD=41.22U
M$300 \$1 PDRIVE_Y DVDD DVDD pfet_06v0_dss L=0.7U W=40U AS=24.4P AD=124.4P
+ PS=41.22U PD=46.22U
M$301 DVDD PDRIVE_Y \$1 DVDD pfet_06v0_dss L=0.7U W=40U AS=124.4P AD=24.4P
+ PS=46.22U PD=41.22U
M$302 \$1 PDRIVE_X DVDD DVDD pfet_06v0_dss L=0.7U W=40U AS=24.4P AD=124.4P
+ PS=41.22U PD=46.22U
M$303 DVDD PDRIVE_X \$1 DVDD pfet_06v0_dss L=0.7U W=40U AS=124.4P AD=31.6P
+ PS=46.22U PD=81.58U
M$304 \$1 NDRIVE_X DVSS DVSS nfet_06v0_dss L=1.15U W=38U AS=30.02P AD=156.18P
+ PS=77.58U PD=46.22U
M$305 DVSS NDRIVE_Y \$1 DVSS nfet_06v0_dss L=1.15U W=38U AS=156.18P AD=23.18P
+ PS=46.22U PD=39.22U
M$306 \$1 NDRIVE_X DVSS DVSS nfet_06v0_dss L=1.15U W=38U AS=23.18P AD=156.18P
+ PS=39.22U PD=46.22U
M$307 DVSS NDRIVE_Y \$1 DVSS nfet_06v0_dss L=1.15U W=38U AS=156.18P AD=23.18P
+ PS=46.22U PD=39.22U
M$308 \$1 NDRIVE_X DVSS DVSS nfet_06v0_dss L=1.15U W=38U AS=23.18P AD=156.18P
+ PS=39.22U PD=46.22U
M$309 DVSS NDRIVE_Y \$1 DVSS nfet_06v0_dss L=1.15U W=38U AS=156.18P AD=23.18P
+ PS=46.22U PD=39.22U
M$310 \$1 NDRIVE_X DVSS DVSS nfet_06v0_dss L=1.15U W=38U AS=23.18P AD=156.18P
+ PS=39.22U PD=46.22U
M$311 DVSS NDRIVE_Y \$1 DVSS nfet_06v0_dss L=1.15U W=38U AS=156.18P AD=30.02P
+ PS=46.22U PD=77.58U
.ENDS inverter_PAD
