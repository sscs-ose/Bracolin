* Extracted by KLayout with GF180MCU LVS runset on : 09/01/2024 11:45

.SUBCKT inv_1x VDDD IN OUT VSSD
M$1 OUT IN VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$2 OUT IN VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
.ENDS inv_1x
