* NGSPICE file created from CM_nfets.ext - technology: gf180mcuD

.subckt CM_nfets VSS OUT1 OUT2 IN
X0 a_n522_n1809# IN.t12 a_n1082_n1809# VSS.t40 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1 a_352_1779# IN.t13 a_n170_882# VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2 a_2346_n15# IN.t14 a_1786_882# VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3 a_1786_n15# IN.t15 a_1264_n1809# VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4 VSS.t75 VSS.t74 VSS.t75 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5 a_1786_n3603# IN.t16 a_1264_n3603# VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6 a_912_n4500# IN.t17 a_352_n4500# VSS.t24 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X7 VSS.t73 VSS.t72 VSS.t73 VSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X8 a_n1082_n1809# IN.t18 a_n1604_n2706# VSS.t33 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X9 VSS.t71 VSS.t70 VSS.t71 VSS.t33 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X10 VSS.t69 VSS.t68 VSS.t69 VSS.t1 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X11 a_352_n2706# IN.t19 a_n170_n3603# VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X12 VSS.t67 VSS.t66 VSS.t67 VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X13 VSS.t65 VSS.t64 VSS.t65 VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X14 VSS.t63 VSS.t62 VSS.t63 VSS.t24 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X15 a_2346_1779# IN.t20 a_1786_2676# VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X16 a_n522_882# IN.t21 a_n1082_1779# VSS.t40 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X17 VSS.t61 VSS.t60 VSS.t61 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X18 a_n1082_1779# IN.t22 a_n1604_1779# VSS.t33 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X19 a_1786_1779# IN.t23 a_1264_882# VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X20 a_912_882# IN.t24 a_352_882# VSS.t24 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X21 VSS.t59 VSS.t58 VSS.t59 VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X22 a_2346_n2706# IN.t25 a_1786_n2706# VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X23 VSS.t57 VSS.t56 VSS.t57 VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X24 a_1786_n4500# IN.t26 a_n522_n4500# VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X25 VSS.t55 VSS.t54 VSS.t55 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X26 a_912_1779# IN.t27 a_352_1779# VSS.t24 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X27 a_2346_n15# IN.t28 a_1786_n15# VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X28 a_n522_n3603# IN.t29 a_n1082_n2706# VSS.t40 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X29 a_352_2676# IN.t30 a_n522_n912.t0 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X30 VSS.t53 VSS.t52 VSS.t53 VSS.t7 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X31 IN IN.t0 VSS.t86 VSS.t24 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X32 a_n1082_n2706# IN.t32 a_n1604_n2706# VSS.t33 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X33 VSS.t51 VSS.t50 VSS.t51 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X34 a_352_n3603# IN.t33 a_n170_n3603# VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X35 VSS.t49 VSS.t48 VSS.t49 VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X36 VSS.t47 VSS.t46 VSS.t47 VSS.t19 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X37 OUT1 IN.t34 a_n1082_2676# VSS.t40 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X38 IN IN.t10 VSS.t85 VSS.t24 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X39 a_1786_2676# IN.t36 VSS.t84 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X40 VSS.t45 VSS.t44 VSS.t45 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X41 VSS.t43 VSS.t42 VSS.t43 VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X42 a_2346_n4500# IN.t37 a_1786_n3603# VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X43 VSS.t41 VSS.t39 VSS.t41 VSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X44 VSS.t38 VSS.t37 VSS.t38 VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X45 a_n1082_2676# IN.t38 a_n1604_1779# VSS.t33 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X46 a_1786_n1809# IN.t39 a_1264_n1809# VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X47 VSS.t36 VSS.t35 VSS.t36 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X48 VSS.t34 VSS.t32 VSS.t34 VSS.t33 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X49 a_912_1779# IN.t40 a_352_2676# VSS.t24 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X50 a_n1082_882# IN.t41 a_n1604_n15# VSS.t33 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X51 a_n522_n3603# IN.t42 a_n1082_n3603# VSS.t40 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X52 a_352_n4500# IN.t43 VSS.t83 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X53 a_912_n2706# IN.t44 a_1786_n912# VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X54 VSS.t31 VSS.t30 VSS.t31 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X55 a_912_n2706# IN.t45 a_352_n2706# VSS.t24 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X56 a_n1082_n3603# IN.t46 a_n1604_n4500# VSS.t33 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X57 a_n522_882# IN.t47 a_n1082_882# VSS.t40 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X58 VSS.t29 VSS.t28 VSS.t29 VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X59 VSS.t27 VSS.t26 VSS.t27 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X60 a_2346_n4500# IN.t48 a_1786_n4500# VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X61 VSS IN.t8 IN.t9 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X62 a_352_882# IN.t49 a_n170_882# VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X63 a_n522_n4500# IN.t50 a_n1082_n4500# VSS.t40 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X64 a_n1082_n15# IN.t51 a_n1604_n15# VSS.t33 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X65 a_1786_n2706# IN.t52 a_1264_n3603# VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X66 VSS.t25 VSS.t23 VSS.t25 VSS.t24 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X67 VSS.t22 VSS.t21 VSS.t22 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X68 a_n1082_n4500# IN.t53 a_n1604_n4500# VSS.t33 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X69 VSS.t20 VSS.t18 VSS.t20 VSS.t19 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X70 VSS.t17 VSS.t16 VSS.t17 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X71 a_1786_882# IN.t54 a_1264_882# VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X72 a_1786_n912# IN.t56 a_912_882# VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X73 VSS IN.t6 IN.t7 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X74 a_n522_n1809# IN.t57 a_n1082_n15# VSS.t40 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X75 VSS.t15 VSS.t14 VSS.t15 VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X76 a_n1082_n912# IN.t58 OUT2.t0 VSS.t33 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X77 a_912_n4500# IN.t59 a_352_n3603# VSS.t24 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X78 a_2346_1779# IN.t60 a_1786_1779# VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X79 VSS.t13 VSS.t11 VSS.t13 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X80 VSS.t10 VSS.t9 VSS.t10 VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X81 IN IN.t2 VSS.t78 VSS.t24 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X82 VSS.t8 VSS.t6 VSS.t8 VSS.t7 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X83 VSS IN.t4 IN.t5 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X84 VSS.t5 VSS.t3 VSS.t5 VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X85 a_2346_n2706# IN.t62 a_1786_n1809# VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X86 VSS.t2 VSS.t0 VSS.t2 VSS.t1 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
R0 IN.n119 IN.t38 10.1674
R1 IN.n120 IN.t38 10.1674
R2 IN.n107 IN.t22 10.1674
R3 IN.t22 IN.n106 10.1674
R4 IN.n95 IN.t41 10.1674
R5 IN.t41 IN.n94 10.1674
R6 IN.t51 IN.n18 10.1674
R7 IN.n19 IN.t51 10.1674
R8 IN.t18 IN.n42 10.1674
R9 IN.n43 IN.t18 10.1674
R10 IN.n64 IN.t46 10.1674
R11 IN.t46 IN.n63 10.1674
R12 IN.n54 IN.t53 10.1674
R13 IN.n31 IN.t58 10.1674
R14 IN.t58 IN.n30 10.1674
R15 IN.t32 IN.n75 10.1674
R16 IN.n76 IN.t32 10.1674
R17 IN.t20 IN.n3 10.1674
R18 IN.n4 IN.t20 10.1674
R19 IN.n109 IN.t60 10.1674
R20 IN.t60 IN.n108 10.1674
R21 IN.n97 IN.t14 10.1674
R22 IN.t14 IN.n96 10.1674
R23 IN.t28 IN.n20 10.1674
R24 IN.n21 IN.t28 10.1674
R25 IN.t62 IN.n44 10.1674
R26 IN.n45 IN.t62 10.1674
R27 IN.n66 IN.t37 10.1674
R28 IN.t37 IN.n65 10.1674
R29 IN.n56 IN.t48 10.1674
R30 IN.n33 IN.t44 10.1674
R31 IN.t44 IN.n32 10.1674
R32 IN.t25 IN.n77 10.1674
R33 IN.n78 IN.t25 10.1674
R34 IN.t53 IN.n53 10.1409
R35 IN.t48 IN.n55 10.1409
R36 IN.t50 IN.n53 9.54631
R37 IN.n59 IN.t43 9.54631
R38 IN.t17 IN.n52 9.54631
R39 IN.n55 IN.t26 9.54631
R40 IN.n120 IN.t34 9.54355
R41 IN.t34 IN.n119 9.54355
R42 IN.n118 IN.t30 9.54355
R43 IN.n5 IN.t40 9.54355
R44 IN.t40 IN.n2 9.54355
R45 IN.n4 IN.t36 9.54355
R46 IN.n3 IN.t36 9.54355
R47 IN.t21 IN.n106 9.54355
R48 IN.n107 IN.t21 9.54355
R49 IN.n113 IN.t13 9.54355
R50 IN.t13 IN.n112 9.54355
R51 IN.t27 IN.n105 9.54355
R52 IN.n110 IN.t27 9.54355
R53 IN.n108 IN.t23 9.54355
R54 IN.n109 IN.t23 9.54355
R55 IN.t47 IN.n94 9.54355
R56 IN.n95 IN.t47 9.54355
R57 IN.n101 IN.t49 9.54355
R58 IN.t49 IN.n100 9.54355
R59 IN.t24 IN.n93 9.54355
R60 IN.n98 IN.t24 9.54355
R61 IN.n96 IN.t54 9.54355
R62 IN.n97 IN.t54 9.54355
R63 IN.n19 IN.t57 9.54355
R64 IN.t57 IN.n18 9.54355
R65 IN.t4 IN.n24 9.54355
R66 IN.n25 IN.t4 9.54355
R67 IN.n22 IN.t10 9.54355
R68 IN.t10 IN.n17 9.54355
R69 IN.n21 IN.t15 9.54355
R70 IN.n20 IN.t15 9.54355
R71 IN.n43 IN.t12 9.54355
R72 IN.t12 IN.n42 9.54355
R73 IN.t6 IN.n48 9.54355
R74 IN.n49 IN.t6 9.54355
R75 IN.n46 IN.t0 9.54355
R76 IN.t0 IN.n41 9.54355
R77 IN.n45 IN.t39 9.54355
R78 IN.n44 IN.t39 9.54355
R79 IN.t42 IN.n63 9.54355
R80 IN.n64 IN.t42 9.54355
R81 IN.n70 IN.t33 9.54355
R82 IN.t33 IN.n69 9.54355
R83 IN.t59 IN.n62 9.54355
R84 IN.n67 IN.t59 9.54355
R85 IN.n65 IN.t16 9.54355
R86 IN.n66 IN.t16 9.54355
R87 IN.n54 IN.t50 9.54355
R88 IN.t43 IN.n58 9.54355
R89 IN.n57 IN.t17 9.54355
R90 IN.n56 IN.t26 9.54355
R91 IN.t55 IN.n30 9.54355
R92 IN.n31 IN.t55 9.54355
R93 IN.n37 IN.t8 9.54355
R94 IN.t8 IN.n36 9.54355
R95 IN.t2 IN.n29 9.54355
R96 IN.n34 IN.t2 9.54355
R97 IN.n32 IN.t56 9.54355
R98 IN.n33 IN.t56 9.54355
R99 IN.n76 IN.t29 9.54355
R100 IN.t29 IN.n75 9.54355
R101 IN.t19 IN.n81 9.54355
R102 IN.n82 IN.t19 9.54355
R103 IN.n79 IN.t45 9.54355
R104 IN.t45 IN.n74 9.54355
R105 IN.n78 IN.t52 9.54355
R106 IN.n77 IN.t52 9.54355
R107 IN.n6 IN.t30 8.06917
R108 IN.n7 IN.n6 4.64379
R109 IN.n1 IN.n0 4.5005
R110 IN.n122 IN.n121 4.5005
R111 IN.n12 IN.n11 3.3605
R112 IN.n14 IN.n13 3.3605
R113 IN.n16 IN.n15 3.3605
R114 IN.n89 IN.t5 3.3605
R115 IN.n88 IN.t9 3.3605
R116 IN.n87 IN.t7 3.3605
R117 IN.n86 IN.n16 2.59662
R118 IN.n90 IN.n12 2.59544
R119 IN.n87 IN.n86 2.58354
R120 IN.n90 IN.n89 2.58235
R121 IN.n61 IN.n60 1.59324
R122 IN.n80 IN.n73 1.5005
R123 IN.n86 IN.n85 1.5005
R124 IN.n39 IN.n38 1.5005
R125 IN.n91 IN.n90 1.5005
R126 IN.n72 IN.n71 1.5005
R127 IN.n68 IN.n61 1.5005
R128 IN.n84 IN.n83 1.5005
R129 IN.n47 IN.n40 1.5005
R130 IN.n51 IN.n50 1.5005
R131 IN.n35 IN.n28 1.5005
R132 IN.n23 IN.n10 1.5005
R133 IN.n27 IN.n26 1.5005
R134 IN.n103 IN.n102 1.5005
R135 IN.n99 IN.n92 1.5005
R136 IN.n115 IN.n114 1.5005
R137 IN.n111 IN.n104 1.5005
R138 IN.n9 IN.n8 1.5005
R139 IN.n117 IN.n116 1.5005
R140 IN.n89 IN.n88 1.06274
R141 IN.n88 IN.n87 1.06274
R142 IN.n14 IN.n12 1.06274
R143 IN.n16 IN.n14 1.06274
R144 IN.n3 IN.n2 0.97759
R145 IN.n119 IN.n118 0.97759
R146 IN.n5 IN.n4 0.97759
R147 IN.n110 IN.n109 0.97759
R148 IN.n112 IN.n107 0.97759
R149 IN.n108 IN.n105 0.97759
R150 IN.n113 IN.n106 0.97759
R151 IN.n98 IN.n97 0.97759
R152 IN.n100 IN.n95 0.97759
R153 IN.n96 IN.n93 0.97759
R154 IN.n101 IN.n94 0.97759
R155 IN.n20 IN.n17 0.97759
R156 IN.n25 IN.n18 0.97759
R157 IN.n22 IN.n21 0.97759
R158 IN.n24 IN.n19 0.97759
R159 IN.n44 IN.n41 0.97759
R160 IN.n49 IN.n42 0.97759
R161 IN.n46 IN.n45 0.97759
R162 IN.n48 IN.n43 0.97759
R163 IN.n67 IN.n66 0.97759
R164 IN.n69 IN.n64 0.97759
R165 IN.n65 IN.n62 0.97759
R166 IN.n70 IN.n63 0.97759
R167 IN.n57 IN.n56 0.97759
R168 IN.n58 IN.n54 0.97759
R169 IN.n34 IN.n33 0.97759
R170 IN.n36 IN.n31 0.97759
R171 IN.n32 IN.n29 0.97759
R172 IN.n37 IN.n30 0.97759
R173 IN.n77 IN.n74 0.97759
R174 IN.n82 IN.n75 0.97759
R175 IN.n79 IN.n78 0.97759
R176 IN.n81 IN.n76 0.97759
R177 IN.n55 IN.n52 0.931516
R178 IN.n59 IN.n53 0.931516
R179 IN.n121 IN.n120 0.840888
R180 IN.n58 IN.n57 0.62434
R181 IN.n117 IN.n2 0.314952
R182 IN.n8 IN.n5 0.314952
R183 IN.n111 IN.n110 0.314952
R184 IN.n114 IN.n105 0.314952
R185 IN.n99 IN.n98 0.314952
R186 IN.n102 IN.n93 0.314952
R187 IN.n26 IN.n17 0.314952
R188 IN.n23 IN.n22 0.314952
R189 IN.n50 IN.n41 0.314952
R190 IN.n47 IN.n46 0.314952
R191 IN.n68 IN.n67 0.314952
R192 IN.n71 IN.n62 0.314952
R193 IN.n35 IN.n34 0.314952
R194 IN.n38 IN.n29 0.314952
R195 IN.n83 IN.n74 0.314952
R196 IN.n80 IN.n79 0.314952
R197 IN.n118 IN.n117 0.309888
R198 IN.n112 IN.n111 0.309888
R199 IN.n114 IN.n113 0.309888
R200 IN.n100 IN.n99 0.309888
R201 IN.n102 IN.n101 0.309888
R202 IN.n26 IN.n25 0.309888
R203 IN.n24 IN.n23 0.309888
R204 IN.n50 IN.n49 0.309888
R205 IN.n48 IN.n47 0.309888
R206 IN.n69 IN.n68 0.309888
R207 IN.n71 IN.n70 0.309888
R208 IN.n36 IN.n35 0.309888
R209 IN.n38 IN.n37 0.309888
R210 IN.n83 IN.n82 0.309888
R211 IN.n81 IN.n80 0.309888
R212 IN.n60 IN.n52 0.300213
R213 IN.n60 IN.n59 0.295374
R214 IN.n115 IN.n104 0.180804
R215 IN.n116 IN.n9 0.1805
R216 IN.n72 IN.n61 0.1805
R217 IN.n51 IN.n40 0.179588
R218 IN.n103 IN.n92 0.179284
R219 IN.n27 IN.n10 0.179284
R220 IN.n84 IN.n73 0.179284
R221 IN.n39 IN.n28 0.178676
R222 IN.n8 IN.n7 0.17375
R223 IN.n122 IN.n0 0.147342
R224 IN.n7 IN.n1 0.14
R225 IN.n121 IN.n1 0.14
R226 IN.n40 IN.n39 0.0947568
R227 IN.n28 IN.n27 0.0944527
R228 IN.n73 IN.n72 0.0944527
R229 IN.n116 IN.n115 0.0938446
R230 IN.n104 IN.n103 0.0932365
R231 IN.n9 IN 0.0798581
R232 IN.n91 IN.n10 0.0482365
R233 IN.n85 IN.n51 0.0482365
R234 IN IN.n122 0.0478684
R235 IN.n92 IN.n91 0.0467162
R236 IN.n85 IN.n84 0.0464122
R237 IN.n6 IN.n0 0.00405263
R238 VSS.n89 VSS.n40 752.225
R239 VSS.n91 VSS.n40 750.567
R240 VSS.n89 VSS.n39 750.383
R241 VSS.n91 VSS.n39 748.725
R242 VSS.t19 VSS.t12 275.589
R243 VSS.t33 VSS.t4 275.589
R244 VSS.t24 VSS.t1 274.022
R245 VSS.t7 VSS.t40 274.022
R246 VSS.t1 VSS.t19 175.575
R247 VSS.t40 VSS.t33 175.575
R248 VSS.t12 VSS.n39 146.779
R249 VSS.t4 VSS.n40 146.779
R250 VSS.n90 VSS.t7 90.9227
R251 VSS.n90 VSS.t24 84.6522
R252 VSS.t60 VSS.n54 8.06917
R253 VSS.n55 VSS.t60 8.06917
R254 VSS.t11 VSS.n52 8.06917
R255 VSS.n53 VSS.t11 8.06917
R256 VSS.t44 VSS.n50 8.06917
R257 VSS.n51 VSS.t44 8.06917
R258 VSS.t26 VSS.n2 8.06917
R259 VSS.n49 VSS.t26 8.06917
R260 VSS.n127 VSS.t30 8.06917
R261 VSS.t30 VSS.n126 8.06917
R262 VSS.n23 VSS.t21 8.06917
R263 VSS.t21 VSS.n22 8.06917
R264 VSS.n25 VSS.t74 8.06917
R265 VSS.t74 VSS.n24 8.06917
R266 VSS.n27 VSS.t50 8.06917
R267 VSS.t50 VSS.n26 8.06917
R268 VSS.n29 VSS.t35 8.06917
R269 VSS.t35 VSS.n28 8.06917
R270 VSS.t37 VSS.n76 8.06917
R271 VSS.n77 VSS.t37 8.06917
R272 VSS.t56 VSS.n74 8.06917
R273 VSS.n75 VSS.t56 8.06917
R274 VSS.t9 VSS.n72 8.06917
R275 VSS.n73 VSS.t9 8.06917
R276 VSS.t64 VSS.n6 8.06917
R277 VSS.n71 VSS.t64 8.06917
R278 VSS.t14 VSS.n120 8.06917
R279 VSS.n121 VSS.t14 8.06917
R280 VSS.t3 VSS.n110 8.06917
R281 VSS.n111 VSS.t3 8.06917
R282 VSS.t58 VSS.n108 8.06917
R283 VSS.n109 VSS.t58 8.06917
R284 VSS.t42 VSS.n106 8.06917
R285 VSS.n107 VSS.t42 8.06917
R286 VSS.t28 VSS.n104 8.06917
R287 VSS.n105 VSS.t28 8.06917
R288 VSS.n124 VSS.n123 4.21074
R289 VSS.n118 VSS.n1 4.21074
R290 VSS.n119 VSS.n118 4.19794
R291 VSS.n123 VSS.n122 4.19794
R292 VSS.n44 VSS.t16 4.03583
R293 VSS.n59 VSS.t18 4.03583
R294 VSS.n43 VSS.t68 4.03583
R295 VSS.n41 VSS.t62 4.03583
R296 VSS.n42 VSS.t6 4.03583
R297 VSS.n65 VSS.t72 4.03583
R298 VSS.n81 VSS.t70 4.03583
R299 VSS.n66 VSS.t66 4.03583
R300 VSS.n17 VSS.t54 4.03583
R301 VSS.n33 VSS.t46 4.03583
R302 VSS.n16 VSS.t0 4.03583
R303 VSS.n38 VSS.t23 4.03583
R304 VSS.n15 VSS.t52 4.03583
R305 VSS.n98 VSS.t39 4.03583
R306 VSS.n14 VSS.t32 4.03583
R307 VSS.n13 VSS.t48 4.03583
R308 VSS.n96 VSS.t83 3.9481
R309 VSS.n63 VSS.t84 3.78612
R310 VSS.n103 VSS.t49 3.37771
R311 VSS.t55 VSS.n30 3.37771
R312 VSS.t67 VSS.n78 3.37771
R313 VSS.t17 VSS.n56 3.37771
R314 VSS.t49 VSS.n102 3.3605
R315 VSS.n101 VSS.t34 3.3605
R316 VSS.n97 VSS.t41 3.3605
R317 VSS.n95 VSS.t53 3.3605
R318 VSS.n37 VSS.t25 3.3605
R319 VSS.n36 VSS.t2 3.3605
R320 VSS.n32 VSS.t47 3.3605
R321 VSS.n31 VSS.t55 3.3605
R322 VSS.n79 VSS.t67 3.3605
R323 VSS.n80 VSS.t71 3.3605
R324 VSS.n84 VSS.t73 3.3605
R325 VSS.t8 VSS.n85 3.3605
R326 VSS.t63 VSS.n64 3.3605
R327 VSS.n62 VSS.t69 3.3605
R328 VSS.n58 VSS.t20 3.3605
R329 VSS.n57 VSS.t17 3.3605
R330 VSS.n117 VSS.n116 2.58721
R331 VSS.n5 VSS.n4 2.58366
R332 VSS.n114 VSS.n113 2.1005
R333 VSS.n61 VSS.n60 2.1005
R334 VSS.n87 VSS.n86 2.1005
R335 VSS.n83 VSS.n82 2.1005
R336 VSS.n35 VSS.n34 2.1005
R337 VSS.n94 VSS.n93 2.1005
R338 VSS.n100 VSS.n99 2.1005
R339 VSS.n45 VSS.t61 1.6805
R340 VSS.n46 VSS.t13 1.6805
R341 VSS.n47 VSS.t45 1.6805
R342 VSS.n48 VSS.t27 1.6805
R343 VSS.n125 VSS.t31 1.6805
R344 VSS.n21 VSS.t22 1.6805
R345 VSS.n20 VSS.t75 1.6805
R346 VSS.n19 VSS.t51 1.6805
R347 VSS.n18 VSS.t36 1.6805
R348 VSS.n67 VSS.t38 1.6805
R349 VSS.n68 VSS.t57 1.6805
R350 VSS.n69 VSS.t10 1.6805
R351 VSS.n70 VSS.t65 1.6805
R352 VSS.n7 VSS.t15 1.6805
R353 VSS.n9 VSS.t5 1.6805
R354 VSS.n10 VSS.t59 1.6805
R355 VSS.n11 VSS.t43 1.6805
R356 VSS.n12 VSS.t29 1.6805
R357 VSS.n123 VSS.n5 1.47409
R358 VSS.n118 VSS.n117 1.47409
R359 VSS.n100 VSS.t41 1.2605
R360 VSS.t34 VSS.n100 1.2605
R361 VSS.n94 VSS.t25 1.2605
R362 VSS.t53 VSS.n94 1.2605
R363 VSS.n35 VSS.t47 1.2605
R364 VSS.t2 VSS.n35 1.2605
R365 VSS.n116 VSS.t86 1.2605
R366 VSS.n116 VSS.n115 1.2605
R367 VSS.n113 VSS.t78 1.2605
R368 VSS.n113 VSS.n112 1.2605
R369 VSS.n4 VSS.t85 1.2605
R370 VSS.n4 VSS.n3 1.2605
R371 VSS.t73 VSS.n83 1.2605
R372 VSS.n83 VSS.t71 1.2605
R373 VSS.n86 VSS.t63 1.2605
R374 VSS.n86 VSS.t8 1.2605
R375 VSS.n61 VSS.t20 1.2605
R376 VSS.t69 VSS.n61 1.2605
R377 VSS.n114 VSS.n5 0.489579
R378 VSS.n117 VSS.n114 0.486026
R379 VSS.n89 VSS.n88 0.08175
R380 VSS.n90 VSS.n89 0.08175
R381 VSS.n92 VSS.n91 0.08175
R382 VSS.n91 VSS.n90 0.08175
R383 VSS.n40 VSS.n8 0.0490981
R384 VSS.n39 VSS.n0 0.0490981
R385 VSS.n78 VSS.n77 0.0414574
R386 VSS.n56 VSS.n55 0.0414574
R387 VSS.n104 VSS.n103 0.0412447
R388 VSS.n30 VSS.n29 0.0412447
R389 VSS.n76 VSS.n75 0.0329468
R390 VSS.n74 VSS.n73 0.0329468
R391 VSS.n72 VSS.n71 0.0329468
R392 VSS.n110 VSS.n109 0.0329468
R393 VSS.n108 VSS.n107 0.0329468
R394 VSS.n106 VSS.n105 0.0329468
R395 VSS.n54 VSS.n53 0.0329468
R396 VSS.n52 VSS.n51 0.0329468
R397 VSS.n50 VSS.n49 0.0329468
R398 VSS.n24 VSS.n23 0.0329468
R399 VSS.n26 VSS.n25 0.0329468
R400 VSS.n28 VSS.n27 0.0329468
R401 VSS.n77 VSS.n67 0.0319894
R402 VSS.n76 VSS.n67 0.0319894
R403 VSS.n75 VSS.n68 0.0319894
R404 VSS.n74 VSS.n68 0.0319894
R405 VSS.n73 VSS.n69 0.0319894
R406 VSS.n72 VSS.n69 0.0319894
R407 VSS.n71 VSS.n70 0.0319894
R408 VSS.n70 VSS.n6 0.0319894
R409 VSS.n121 VSS.n7 0.0319894
R410 VSS.n111 VSS.n9 0.0319894
R411 VSS.n110 VSS.n9 0.0319894
R412 VSS.n109 VSS.n10 0.0319894
R413 VSS.n108 VSS.n10 0.0319894
R414 VSS.n107 VSS.n11 0.0319894
R415 VSS.n106 VSS.n11 0.0319894
R416 VSS.n105 VSS.n12 0.0319894
R417 VSS.n104 VSS.n12 0.0319894
R418 VSS.n55 VSS.n45 0.0319894
R419 VSS.n54 VSS.n45 0.0319894
R420 VSS.n53 VSS.n46 0.0319894
R421 VSS.n52 VSS.n46 0.0319894
R422 VSS.n51 VSS.n47 0.0319894
R423 VSS.n50 VSS.n47 0.0319894
R424 VSS.n49 VSS.n48 0.0319894
R425 VSS.n48 VSS.n2 0.0319894
R426 VSS.n126 VSS.n125 0.0319894
R427 VSS.n22 VSS.n21 0.0319894
R428 VSS.n23 VSS.n21 0.0319894
R429 VSS.n24 VSS.n20 0.0319894
R430 VSS.n25 VSS.n20 0.0319894
R431 VSS.n26 VSS.n19 0.0319894
R432 VSS.n27 VSS.n19 0.0319894
R433 VSS.n28 VSS.n18 0.0319894
R434 VSS.n29 VSS.n18 0.0319894
R435 VSS.n58 VSS.n57 0.031877
R436 VSS.n80 VSS.n79 0.031877
R437 VSS.n32 VSS.n31 0.031877
R438 VSS.n102 VSS.n101 0.031877
R439 VSS.n85 VSS.n84 0.0313852
R440 VSS.n37 VSS.n36 0.0313852
R441 VSS.n120 VSS.n8 0.0311383
R442 VSS.n97 VSS.n96 0.0300082
R443 VSS VSS.n127 0.0280532
R444 VSS.n57 VSS.n44 0.028041
R445 VSS.n59 VSS.n58 0.028041
R446 VSS.n60 VSS.n59 0.028041
R447 VSS.n60 VSS.n43 0.028041
R448 VSS.n62 VSS.n43 0.028041
R449 VSS.n64 VSS.n63 0.028041
R450 VSS.n64 VSS.n41 0.028041
R451 VSS.n87 VSS.n42 0.028041
R452 VSS.n85 VSS.n42 0.028041
R453 VSS.n84 VSS.n65 0.028041
R454 VSS.n82 VSS.n65 0.028041
R455 VSS.n82 VSS.n81 0.028041
R456 VSS.n81 VSS.n80 0.028041
R457 VSS.n79 VSS.n66 0.028041
R458 VSS.n31 VSS.n17 0.028041
R459 VSS.n33 VSS.n32 0.028041
R460 VSS.n34 VSS.n33 0.028041
R461 VSS.n34 VSS.n16 0.028041
R462 VSS.n36 VSS.n16 0.028041
R463 VSS.n38 VSS.n37 0.028041
R464 VSS.n93 VSS.n15 0.028041
R465 VSS.n95 VSS.n15 0.028041
R466 VSS.n98 VSS.n97 0.028041
R467 VSS.n99 VSS.n98 0.028041
R468 VSS.n99 VSS.n14 0.028041
R469 VSS.n101 VSS.n14 0.028041
R470 VSS.n102 VSS.n13 0.028041
R471 VSS.n88 VSS.n41 0.0270574
R472 VSS.n92 VSS.n38 0.0270574
R473 VSS.n122 VSS.n121 0.0169894
R474 VSS.n126 VSS.n124 0.0169894
R475 VSS.n119 VSS.n111 0.0167766
R476 VSS.n22 VSS.n1 0.0167766
R477 VSS.n120 VSS.n119 0.0166702
R478 VSS.n127 VSS.n1 0.0166702
R479 VSS.n122 VSS.n6 0.0164574
R480 VSS.n124 VSS.n2 0.0164574
R481 VSS.n56 VSS.n44 0.0108279
R482 VSS.n78 VSS.n66 0.0108279
R483 VSS.n30 VSS.n17 0.0108279
R484 VSS.n103 VSS.n13 0.0108279
R485 VSS.n63 VSS.n62 0.00384426
R486 VSS VSS.n0 0.00358511
R487 VSS.n96 VSS.n95 0.00187705
R488 VSS.n88 VSS.n87 0.00148361
R489 VSS.n93 VSS.n92 0.00148361
R490 VSS.n8 VSS.n7 0.00135106
R491 VSS.n125 VSS.n0 0.00135106
R492 a_n522_n912.t0 a_n522_n912.n0 13.2434
R493 OUT1.n6 OUT1.n5 4.5005
R494 OUT1.n5 OUT1.n4 4.5005
R495 OUT1.n4 OUT1.n0 4.5005
R496 OUT1.n6 OUT1.n0 4.5005
R497 OUT1.n2 OUT1.n1 3.3605
R498 OUT1.n3 OUT1 1.41787
R499 OUT1 OUT1.n6 0.0365963
R500 OUT1.n3 OUT1.n0 0.0309545
R501 OUT1.n6 OUT1.n2 0.0269706
R502 OUT1.n4 OUT1.n2 0.0269706
R503 OUT1.n5 OUT1.n3 0.0264091
R504 OUT2.n5 OUT2.n4 4.5005
R505 OUT2.n4 OUT2.n3 4.5005
R506 OUT2.n3 OUT2.n0 4.5005
R507 OUT2.n5 OUT2.n0 4.5005
R508 OUT2.n1 OUT2.t0 3.3605
R509 OUT2.n2 OUT2 3.25949
R510 OUT2 OUT2.n5 0.0351524
R511 OUT2.n2 OUT2.n0 0.0309545
R512 OUT2.n5 OUT2.n1 0.0269706
R513 OUT2.n3 OUT2.n1 0.0269706
R514 OUT2.n4 OUT2.n2 0.0264091
C0 a_n1082_n4500# a_n1604_n4500# 0.0284f
C1 a_352_1779# a_n170_882# 0.0284f
C2 IN a_1786_n1809# 0.111984f
C3 a_n1082_n3603# a_n522_n3603# 0.0284f
C4 IN a_2346_1779# 0.234631f
C5 IN a_1786_n3603# 0.112519f
C6 a_n170_n3603# a_352_n2706# 0.0284f
C7 a_n1082_n15# a_n1604_n15# 0.0284f
C8 a_1786_n3603# a_1264_n3603# 0.0284f
C9 a_2346_1779# a_1786_2676# 0.0284f
C10 IN a_n1082_n15# 0.111376f
C11 a_n1082_882# a_n522_882# 0.0284f
C12 a_n1082_n15# a_n522_n1809# 0.035468f
C13 IN a_n170_882# 0.403137f
C14 a_n522_n3603# a_n170_n3603# 0.210644f
C15 IN a_n522_n4500# 1.43426f
C16 IN a_n1082_n912# 0.111058f
C17 a_912_882# a_352_882# 0.037577f
C18 a_n522_n4500# a_912_n4500# 0.054819f
C19 IN a_n1082_n3603# 0.112534f
C20 a_352_n3603# a_n170_n3603# 0.0284f
C21 IN a_1786_1779# 0.112493f
C22 a_1786_n2706# a_2346_n2706# 0.0284f
C23 IN a_n1082_2676# 0.10943f
C24 a_n170_882# a_n522_882# 0.210644f
C25 IN a_n1604_n2706# 0.274115f
C26 a_n522_n4500# a_n1082_n4500# 0.0284f
C27 IN a_n170_n3603# 0.418388f
C28 a_912_882# a_1264_n1809# 0.534125f
C29 IN a_352_882# 0.143422f
C30 OUT2 a_n1604_n15# 0.085733f
C31 a_n1082_n1809# a_n1604_n2706# 0.0284f
C32 OUT2 IN 0.545908f
C33 IN a_352_n2706# 0.14613f
C34 IN a_1786_882# 0.110898f
C35 OUT2 a_n522_n1809# 0.075896f
C36 IN a_2346_n2706# 0.243632f
C37 IN a_n1082_1779# 0.11029f
C38 a_1786_n4500# a_n522_n4500# 0.0284f
C39 IN a_2346_n4500# 0.235347f
C40 IN a_n522_n3603# 0.355772f
C41 a_912_882# a_1786_n912# 0.030444f
C42 a_n1082_n2706# a_n1604_n2706# 0.0284f
C43 a_n1082_n3603# a_n1604_n4500# 0.0284f
C44 IN a_1264_n1809# 1.17554f
C45 a_2346_n15# a_1786_882# 0.0284f
C46 IN a_912_882# 1.71798f
C47 IN a_1786_n2706# 0.112493f
C48 a_1786_1779# a_1264_882# 0.0284f
C49 a_912_1779# a_352_1779# 0.0284f
C50 IN a_352_1779# 0.145777f
C51 IN a_352_n4500# 0.144763f
C52 IN a_352_n3603# 0.145782f
C53 a_1786_n2706# a_1264_n3603# 0.0284f
C54 a_n1082_2676# a_n1604_1779# 0.0284f
C55 a_n522_882# a_n1082_1779# 0.0284f
C56 IN a_1786_n912# 0.111376f
C57 a_n522_n3603# a_n1082_n2706# 0.0284f
C58 a_352_n4500# a_912_n4500# 0.0284f
C59 a_912_n4500# a_352_n3603# 0.0284f
C60 IN a_n1604_n15# 0.274083f
C61 IN a_912_1779# 0.405199f
C62 OUT2 a_n1604_1779# 0.078566f
C63 a_1786_882# a_1264_882# 0.0284f
C64 OUT1 a_n1082_2676# 0.037438f
C65 IN a_n522_n1809# 1.15854f
C66 IN a_1264_n3603# 0.388639f
C67 a_1786_1779# a_2346_1779# 0.0284f
C68 IN a_n1082_n1809# 0.111988f
C69 a_912_n2706# a_352_n2706# 0.0284f
C70 a_n1082_1779# a_n1604_1779# 0.0284f
C71 IN a_1786_2676# 0.112059f
C72 a_1786_n15# a_1264_n1809# 0.035574f
C73 IN a_912_n4500# 0.406067f
C74 a_1786_n4500# a_2346_n4500# 0.0284f
C75 a_n1082_n1809# a_n522_n1809# 0.034628f
C76 a_2346_n2706# a_912_n2706# 0.08885f
C77 OUT2 OUT1 0.111964f
C78 a_912_n4500# a_1264_n3603# 0.053799f
C79 IN a_2346_n15# 0.24359f
C80 a_912_882# a_1264_882# 0.062551f
C81 IN a_n1082_n2706# 0.112508f
C82 IN a_n522_882# 0.346971f
C83 a_912_n2706# a_1264_n1809# 0.070243f
C84 IN a_n1082_n4500# 0.112152f
C85 a_2346_n2706# a_1786_n1809# 0.0284f
C86 IN a_1786_n15# 0.111376f
C87 a_352_2676# a_912_1779# 0.0284f
C88 IN a_352_2676# 0.143307f
C89 IN a_n1604_n4500# 0.266274f
C90 a_2346_n4500# a_1786_n3603# 0.0284f
C91 a_352_882# a_n170_882# 0.0284f
C92 a_912_1779# a_1264_882# 0.053799f
C93 IN a_1264_882# 0.416734f
C94 IN a_n1604_1779# 0.265528f
C95 a_1786_n1809# a_1264_n1809# 0.034714f
C96 a_912_n2706# a_1786_n912# 0.034652f
C97 IN a_1786_n4500# 0.112137f
C98 IN a_912_n2706# 1.81086f
C99 OUT2 a_n1082_n912# 0.037147f
C100 a_1786_n15# a_2346_n15# 0.0284f
C101 a_n1082_882# a_n1604_n15# 0.0284f
C102 IN a_n1082_882# 0.11029f
C103 a_1264_n3603# a_912_n2706# 0.16936f
C104 OUT1 IN 0.460317f
.ends

