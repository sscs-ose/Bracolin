* Extracted by KLayout with GF180MCU LVS runset on : 14/04/2024 15:38

.SUBCKT SAR_Asynchronous_top D_C_11 Valid Bit_0 D_C_10 Bit_1 D_C_9 Bit_2 D_C_8
+ Bit_3 D_C_7 Bit_4 D_C_6 VSSD Set D CK11 CK9 CK8 CK7 CK6 CK5 CK4 CK3 CK2 CK1
+ clks VDDD Reset D_C_1 D_C_2 D_C_3 D_C_4 D_C_5 VCM Bit_10 Bit_9 Bit_8 Bit_7
+ Bit_6 Bit_5
M$1 \$151 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$2 \$152 \$151 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$3 \$153 CK11 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$4 \$154 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$5 \$155 \$154 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$6 \$156 \$96 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$7 \$157 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$8 \$158 \$157 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$9 \$159 CK9 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$10 \$160 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$11 \$161 \$160 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$12 \$162 CK8 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$13 \$163 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$14 \$164 \$163 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$15 \$165 CK7 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$16 \$166 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$17 \$167 \$166 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$18 \$168 CK6 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$19 \$169 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$20 \$170 \$169 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$21 \$171 CK5 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$22 \$172 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$23 \$173 \$172 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$24 \$174 CK4 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$25 \$175 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$26 \$176 \$175 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$27 \$177 CK3 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$28 \$178 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$29 \$179 \$178 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$30 \$180 CK2 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$31 \$181 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$32 \$182 \$181 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$33 \$183 CK1 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$34 \$85 \$152 D VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$35 \$971 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$36 \$86 \$85 \$971 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$37 \$972 \$86 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$38 \$87 clks \$972 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$39 \$85 \$151 \$87 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$40 \$89 \$151 \$86 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$41 \$973 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$42 CK11 \$89 \$973 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$43 \$974 CK11 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$44 \$88 Set \$974 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$45 \$89 \$152 \$88 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$46 \$91 \$155 CK11 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$47 \$975 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$48 \$92 \$91 \$975 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$49 \$976 \$92 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$50 \$93 clks \$976 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$51 \$91 \$154 \$93 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$52 \$95 \$154 \$92 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$53 \$977 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$54 \$96 \$95 \$977 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$55 \$978 \$96 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$56 \$94 Set \$978 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$57 \$95 \$155 \$94 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$58 \$97 \$158 \$96 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$59 \$979 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$60 \$98 \$97 \$979 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$61 \$980 \$98 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$62 \$99 clks \$980 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$63 \$97 \$157 \$99 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$64 \$101 \$157 \$98 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$65 \$981 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$66 CK9 \$101 \$981 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$67 \$982 CK9 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$68 \$100 Set \$982 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$69 \$101 \$158 \$100 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$70 \$103 \$161 CK9 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$71 \$983 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$72 \$104 \$103 \$983 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$73 \$984 \$104 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$74 \$105 clks \$984 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$75 \$103 \$160 \$105 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$76 \$107 \$160 \$104 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$77 \$985 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$78 CK8 \$107 \$985 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$79 \$986 CK8 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$80 \$106 Set \$986 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$81 \$107 \$161 \$106 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$82 \$109 \$164 CK8 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$83 \$987 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$84 \$110 \$109 \$987 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$85 \$988 \$110 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$86 \$111 clks \$988 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$87 \$109 \$163 \$111 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$88 \$113 \$163 \$110 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$89 \$989 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$90 CK7 \$113 \$989 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$91 \$990 CK7 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$92 \$112 Set \$990 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$93 \$113 \$164 \$112 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$94 \$115 \$167 CK7 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$95 \$991 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$96 \$116 \$115 \$991 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$97 \$992 \$116 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$98 \$117 clks \$992 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$99 \$115 \$166 \$117 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$100 \$119 \$166 \$116 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$101 \$993 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$102 CK6 \$119 \$993 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$103 \$994 CK6 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$104 \$118 Set \$994 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$105 \$119 \$167 \$118 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$106 \$121 \$170 CK6 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$107 \$995 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$108 \$122 \$121 \$995 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$109 \$996 \$122 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$110 \$123 clks \$996 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$111 \$121 \$169 \$123 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$112 \$125 \$169 \$122 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$113 \$997 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$114 CK5 \$125 \$997 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$115 \$998 CK5 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$116 \$124 Set \$998 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$117 \$125 \$170 \$124 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$118 \$127 \$173 CK5 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$119 \$999 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$120 \$128 \$127 \$999 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$121 \$1000 \$128 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$122 \$129 clks \$1000 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$123 \$127 \$172 \$129 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$124 \$131 \$172 \$128 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$125 \$1001 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$126 CK4 \$131 \$1001 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$127 \$1002 CK4 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$128 \$130 Set \$1002 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$129 \$131 \$173 \$130 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$130 \$133 \$176 CK4 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$131 \$1003 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$132 \$134 \$133 \$1003 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$133 \$1004 \$134 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$134 \$135 clks \$1004 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$135 \$133 \$175 \$135 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$136 \$137 \$175 \$134 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$137 \$1005 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$138 CK3 \$137 \$1005 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$139 \$1006 CK3 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$140 \$136 Set \$1006 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$141 \$137 \$176 \$136 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$142 \$139 \$179 CK3 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$143 \$1007 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$144 \$140 \$139 \$1007 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$145 \$1008 \$140 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$146 \$141 clks \$1008 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$147 \$139 \$178 \$141 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$148 \$143 \$178 \$140 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$149 \$1009 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$150 CK2 \$143 \$1009 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$151 \$1010 CK2 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$152 \$142 Set \$1010 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$153 \$143 \$179 \$142 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$154 \$145 \$182 CK2 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$155 \$1011 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$156 \$146 \$145 \$1011 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$157 \$1012 \$146 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$158 \$147 clks \$1012 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$159 \$145 \$181 \$147 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$160 \$150 \$181 \$146 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$161 \$1013 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$162 CK1 \$150 \$1013 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$163 \$1014 CK1 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$164 \$149 Set \$1014 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$165 \$150 \$182 \$149 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$166 \$1632 \$1806 \$1635 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$167 VDDD \$1635 \$2443 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$168 \$1633 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$169 \$1634 \$1633 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$170 \$2421 \$2558 \$2376 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$171 \$2957 Set \$2421 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$172 \$1600 \$1634 \$1635 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$173 VDDD \$1635 \$2957 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$174 \$2016 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$175 \$1601 \$1600 \$2016 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$176 \$2958 \$2376 \$1635 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$177 VDDD Reset \$2958 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$178 \$2017 \$1601 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$179 \$1602 Reset \$2017 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$180 \$2422 \$2557 \$2376 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$181 \$1600 \$1633 \$1602 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$182 \$2423 \$2557 \$2411 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$183 \$1605 \$1633 \$1601 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$184 \$2959 Reset \$2423 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$185 VDDD \$2422 \$2959 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$186 \$2018 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$187 \$1603 \$1605 \$2018 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$188 \$2960 \$2411 \$2422 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$189 VDDD Set \$2960 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$190 \$2019 \$1603 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$191 D_C_1 \$2558 \$2411 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$192 \$1604 Set \$2019 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$193 \$1605 \$1634 \$1604 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$194 VDDD \$2557 \$2558 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$195 VDDD \$1631 \$2557 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$196 \$1636 \$1603 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$197 VDDD \$1806 \$1631 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$198 VDDD CK1 \$1806 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$199 \$1606 \$1820 \$1640 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$200 VDDD \$1640 \$2445 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$201 \$1638 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$202 \$1639 \$1638 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$203 \$2425 \$2560 \$2377 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$204 \$2961 Set \$2425 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$205 \$1607 \$1639 \$1640 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$206 VDDD \$1640 \$2961 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$207 \$2020 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$208 \$1608 \$1607 \$2020 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$209 \$2962 \$2377 \$1640 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$210 VDDD Reset \$2962 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$211 \$2021 \$1608 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$212 \$1609 Reset \$2021 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$213 \$2426 \$2559 \$2377 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$214 \$1607 \$1638 \$1609 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$215 \$2427 \$2559 \$2412 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$216 \$1612 \$1638 \$1608 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$217 \$2963 Reset \$2427 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$218 VDDD \$2426 \$2963 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$219 \$2022 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$220 \$1610 \$1612 \$2022 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$221 \$2964 \$2412 \$2426 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$222 VDDD Set \$2964 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$223 \$2023 \$1610 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$224 D_C_2 \$2560 \$2412 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$225 \$1611 Set \$2023 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$226 \$1612 \$1639 \$1611 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$227 VDDD \$2559 \$2560 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$228 VDDD \$1637 \$2559 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$229 \$1641 \$1610 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$230 VDDD \$1820 \$1637 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$231 VDDD CK2 \$1820 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$232 \$1643 \$1833 \$1646 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$233 VDDD \$1646 \$2447 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$234 \$1644 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$235 \$1645 \$1644 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$236 \$2429 \$2562 \$2378 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$237 \$2965 Set \$2429 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$238 \$1613 \$1645 \$1646 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$239 VDDD \$1646 \$2965 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$240 \$2024 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$241 \$1614 \$1613 \$2024 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$242 \$2966 \$2378 \$1646 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$243 VDDD Reset \$2966 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$244 \$2025 \$1614 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$245 \$1615 Reset \$2025 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$246 \$2430 \$2561 \$2378 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$247 \$1613 \$1644 \$1615 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$248 \$2431 \$2561 \$2413 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$249 \$1618 \$1644 \$1614 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$250 \$2967 Reset \$2431 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$251 VDDD \$2430 \$2967 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$252 \$2026 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$253 \$1616 \$1618 \$2026 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$254 \$2968 \$2413 \$2430 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$255 VDDD Set \$2968 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$256 \$2027 \$1616 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$257 D_C_3 \$2562 \$2413 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$258 \$1617 Set \$2027 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$259 \$1618 \$1645 \$1617 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$260 VDDD \$2561 \$2562 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$261 VDDD \$1642 \$2561 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$262 \$1647 \$1616 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$263 VDDD \$1833 \$1642 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$264 VDDD CK3 \$1833 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$265 \$1619 \$1846 \$1651 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$266 VDDD \$1651 \$2449 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$267 \$1649 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$268 \$1650 \$1649 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$269 \$2433 \$2564 \$2379 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$270 \$2969 Set \$2433 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$271 \$1620 \$1650 \$1651 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$272 VDDD \$1651 \$2969 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$273 \$2028 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$274 \$1621 \$1620 \$2028 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$275 \$2970 \$2379 \$1651 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$276 VDDD Reset \$2970 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$277 \$2029 \$1621 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$278 \$1622 Reset \$2029 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$279 \$2434 \$2563 \$2379 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$280 \$1620 \$1649 \$1622 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$281 \$2435 \$2563 \$2414 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$282 \$1652 \$1649 \$1621 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$283 \$2971 Reset \$2435 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$284 VDDD \$2434 \$2971 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$285 \$2030 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$286 \$1623 \$1652 \$2030 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$287 \$2972 \$2414 \$2434 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$288 VDDD Set \$2972 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$289 \$2031 \$1623 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$290 D_C_4 \$2564 \$2414 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$291 \$1624 Set \$2031 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$292 \$1652 \$1650 \$1624 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$293 VDDD \$2563 \$2564 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$294 VDDD \$1648 \$2563 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$295 \$1653 \$1623 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$296 VDDD \$1846 \$1648 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$297 VDDD CK4 \$1846 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$298 \$1625 \$1859 \$1657 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$299 VDDD \$1657 \$2451 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$300 \$1655 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$301 \$1656 \$1655 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$302 \$2437 \$2566 \$2380 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$303 \$2973 Set \$2437 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$304 \$1626 \$1656 \$1657 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$305 VDDD \$1657 \$2973 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$306 \$2032 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$307 \$1627 \$1626 \$2032 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$308 \$2974 \$2380 \$1657 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$309 VDDD Reset \$2974 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$310 \$2033 \$1627 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$311 \$1628 Reset \$2033 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$312 \$2438 \$2565 \$2380 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$313 \$1626 \$1655 \$1628 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$314 \$2439 \$2565 \$2415 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$315 \$1658 \$1655 \$1627 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$316 \$2975 Reset \$2439 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$317 VDDD \$2438 \$2975 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$318 \$2034 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$319 \$1629 \$1658 \$2034 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$320 \$2976 \$2415 \$2438 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$321 VDDD Set \$2976 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$322 \$2035 \$1629 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$323 D_C_5 \$2566 \$2415 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$324 \$1630 Set \$2035 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$325 \$1658 \$1656 \$1630 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$326 VDDD \$2565 \$2566 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$327 VDDD \$1654 \$2565 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$328 \$1659 \$1629 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$329 VDDD \$1859 \$1654 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$330 VDDD CK5 \$1859 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$331 VDDD \$3580 \$3397 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$332 \$3398 \$3605 \$3331 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$333 \$3861 Set \$3398 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$334 VDDD \$3580 \$3861 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$335 \$3862 \$3331 \$3580 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$336 VDDD Reset \$3862 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$337 \$3399 \$3579 \$3331 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$338 \$3369 \$3579 \$3362 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$339 \$3863 Reset \$3369 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$340 VDDD \$3399 \$3863 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$341 \$3864 \$3362 \$3399 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$342 VDDD Set \$3864 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$343 \$3370 \$3605 \$3362 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$344 VDDD \$3579 \$3605 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$345 VDDD clks \$3579 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$346 \$3370 \$3400 \$3371 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$347 Bit_0 \$1631 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$348 VDDD \$2442 Bit_0 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$349 \$2442 \$1806 \$1635 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$350 VDDD \$3582 \$3401 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$351 VDDD \$1631 \$2442 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$352 \$3373 \$3627 \$3332 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$353 \$3865 Set \$3373 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$354 VDDD \$3582 \$3865 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$355 \$3866 \$3332 \$3582 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$356 VDDD Reset \$3866 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$357 \$3402 \$3581 \$3332 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$358 \$3374 \$3581 \$3363 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$359 \$3867 Reset \$3374 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$360 VDDD \$3402 \$3867 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$361 \$3868 \$3363 \$3402 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$362 VDDD Set \$3868 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$363 \$3375 \$3627 \$3363 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$364 VDDD \$3581 \$3627 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$365 VDDD clks \$3581 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$366 \$3375 \$3403 \$3376 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$367 Bit_1 \$1637 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$368 VDDD \$2444 Bit_1 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$369 \$2444 \$1820 \$1640 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$370 VDDD \$3584 \$3404 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$371 VDDD \$1637 \$2444 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$372 \$3378 \$3641 \$3333 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$373 \$3869 Set \$3378 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$374 VDDD \$3584 \$3869 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$375 \$3870 \$3333 \$3584 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$376 VDDD Reset \$3870 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$377 \$3379 \$3583 \$3333 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$378 \$3380 \$3583 \$3364 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$379 \$3871 Reset \$3380 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$380 VDDD \$3379 \$3871 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$381 \$3872 \$3364 \$3379 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$382 VDDD Set \$3872 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$383 \$3405 \$3641 \$3364 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$384 VDDD \$3583 \$3641 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$385 VDDD clks \$3583 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$386 \$3405 \$3406 \$3407 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$387 Bit_2 \$1642 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$388 VDDD \$2446 Bit_2 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$389 \$2446 \$1833 \$1646 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$390 VDDD \$3586 \$3408 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$391 VDDD \$1642 \$2446 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$392 \$3382 \$3655 \$3334 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$393 \$3873 Set \$3382 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$394 VDDD \$3586 \$3873 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$395 \$3874 \$3334 \$3586 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$396 VDDD Reset \$3874 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$397 \$3409 \$3585 \$3334 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$398 \$3383 \$3585 \$3365 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$399 \$3875 Reset \$3383 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$400 VDDD \$3409 \$3875 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$401 \$3876 \$3365 \$3409 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$402 VDDD Set \$3876 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$403 \$3384 \$3655 \$3365 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$404 VDDD \$3585 \$3655 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$405 VDDD clks \$3585 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$406 \$3384 \$3410 \$3385 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$407 Bit_3 \$1648 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$408 VDDD \$2448 Bit_3 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$409 \$2448 \$1846 \$1651 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$410 VDDD \$3588 \$3411 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$411 VDDD \$1648 \$2448 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$412 \$3387 \$3669 \$3335 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$413 \$3877 Set \$3387 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$414 VDDD \$3588 \$3877 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$415 \$3878 \$3335 \$3588 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$416 VDDD Reset \$3878 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$417 \$3388 \$3587 \$3335 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$418 \$3389 \$3587 \$3366 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$419 \$3879 Reset \$3389 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$420 VDDD \$3388 \$3879 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$421 \$3880 \$3366 \$3388 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$422 VDDD Set \$3880 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$423 \$3412 \$3669 \$3366 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$424 VDDD \$3587 \$3669 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$425 VDDD clks \$3587 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$426 \$3412 \$3413 \$3390 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$427 Bit_4 \$1654 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$428 VDDD \$2450 Bit_4 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$429 \$2450 \$1859 \$1657 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$430 VDDD \$3590 \$3414 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$431 VDDD \$1654 \$2450 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$432 \$3392 \$3683 \$3336 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$433 \$3881 Set \$3392 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$434 VDDD \$3590 \$3881 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$435 \$3882 \$3336 \$3590 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$436 VDDD Reset \$3882 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$437 \$3415 \$3589 \$3336 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$438 \$3393 \$3589 \$3367 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$439 \$3883 Reset \$3393 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$440 VDDD \$3415 \$3883 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$441 \$3884 \$3367 \$3415 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$442 VDDD Set \$3884 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$443 \$3394 \$3683 \$3367 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$444 VDDD \$3589 \$3683 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$445 VDDD clks \$3589 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$446 \$3394 \$3416 \$3395 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$447 \$3400 CK11 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$448 \$3614 \$3400 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$449 \$4383 \$3614 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$450 \$4384 \$4383 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$451 \$4341 \$4384 D_C_11 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$452 \$4995 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$453 \$4342 \$4341 \$4995 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$454 \$4996 \$4342 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$455 \$4343 Reset \$4996 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$456 \$4341 \$4383 \$4343 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$457 \$4345 \$4383 \$4342 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$458 \$4997 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$459 \$3370 \$4345 \$4997 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$460 \$4998 \$3370 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$461 \$4344 Set \$4998 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$462 \$4345 \$4384 \$4344 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$463 \$4385 \$3370 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$464 \$3403 \$96 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$465 \$3628 \$3403 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$466 \$4386 \$3628 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$467 \$4387 \$4386 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$468 \$4347 \$4387 D_C_10 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$469 \$4999 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$470 \$4348 \$4347 \$4999 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$471 \$5000 \$4348 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$472 \$4349 Reset \$5000 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$473 \$4347 \$4386 \$4349 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$474 \$4351 \$4386 \$4348 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$475 \$5001 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$476 \$3375 \$4351 \$5001 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$477 \$5002 \$3375 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$478 \$4350 Set \$5002 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$479 \$4351 \$4387 \$4350 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$480 \$4388 \$3375 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$481 \$3406 CK9 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$482 \$3642 \$3406 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$483 \$4389 \$3642 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$484 \$4390 \$4389 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$485 \$4353 \$4390 D_C_9 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$486 \$5003 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$487 \$4354 \$4353 \$5003 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$488 \$5004 \$4354 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$489 \$4355 Reset \$5004 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$490 \$4353 \$4389 \$4355 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$491 \$4357 \$4389 \$4354 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$492 \$5005 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$493 \$3405 \$4357 \$5005 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$494 \$5006 \$3405 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$495 \$4356 Set \$5006 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$496 \$4357 \$4390 \$4356 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$497 \$4391 \$3405 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$498 \$3410 CK8 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$499 \$3656 \$3410 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$500 \$4392 \$3656 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$501 \$4393 \$4392 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$502 \$4359 \$4393 D_C_8 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$503 \$5007 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$504 \$4360 \$4359 \$5007 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$505 \$5008 \$4360 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$506 \$4361 Reset \$5008 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$507 \$4359 \$4392 \$4361 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$508 \$4363 \$4392 \$4360 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$509 \$5009 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$510 \$3384 \$4363 \$5009 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$511 \$5010 \$3384 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$512 \$4362 Set \$5010 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$513 \$4363 \$4393 \$4362 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$514 \$4394 \$3384 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$515 \$3413 CK7 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$516 \$3670 \$3413 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$517 \$4395 \$3670 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$518 \$4396 \$4395 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$519 \$4365 \$4396 D_C_7 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$520 \$5011 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$521 \$4366 \$4365 \$5011 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$522 \$5012 \$4366 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$523 \$4367 Reset \$5012 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$524 \$4365 \$4395 \$4367 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$525 \$4369 \$4395 \$4366 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$526 \$5013 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$527 \$3412 \$4369 \$5013 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$528 \$5014 \$3412 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$529 \$4368 Set \$5014 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$530 \$4369 \$4396 \$4368 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$531 \$4397 \$3412 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$532 \$3416 CK6 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$533 \$3684 \$3416 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$534 \$4398 \$3684 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$535 \$4399 \$4398 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$536 \$4371 \$4399 D_C_6 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$537 \$5015 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$538 \$4372 \$4371 \$5015 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$539 \$5016 \$4372 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$540 \$4373 Reset \$5016 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$541 \$4371 \$4398 \$4373 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$542 \$4375 \$4398 \$4372 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$543 \$5017 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$544 \$3394 \$4375 \$5017 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$545 \$5018 \$3394 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$546 \$4374 Set \$5018 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$547 \$4375 \$4399 \$4374 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$548 \$4400 \$3394 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$549 \$4346 \$3614 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$550 \$3370 \$3400 \$4346 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$551 Bit_10 \$4346 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$552 VCM \$3614 Bit_10 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$553 \$4352 \$3628 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$554 \$3375 \$3403 \$4352 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$555 Bit_9 \$4352 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$556 VCM \$3628 Bit_9 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$557 \$4358 \$3642 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$558 \$3405 \$3406 \$4358 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$559 Bit_8 \$4358 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$560 VCM \$3642 Bit_8 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$561 \$4364 \$3656 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$562 \$3384 \$3410 \$4364 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$563 Bit_7 \$4364 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$564 VCM \$3656 Bit_7 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$565 \$4370 \$3670 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$566 \$3412 \$3413 \$4370 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$567 Bit_6 \$4370 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$568 VCM \$3670 Bit_6 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$569 \$4376 \$3684 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$570 \$3394 \$3416 \$4376 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$571 Bit_5 \$4376 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$572 VCM \$3684 Bit_5 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$573 \$85 \$151 D VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$574 \$86 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$575 VSSD \$85 \$86 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$576 \$87 \$86 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$577 VSSD clks \$87 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$578 \$85 \$152 \$87 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$579 \$89 \$152 \$86 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$580 CK11 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$581 VSSD \$89 CK11 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$582 \$88 CK11 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$583 VSSD Set \$88 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$584 \$89 \$151 \$88 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$585 \$91 \$154 CK11 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$586 \$92 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$587 VSSD \$91 \$92 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$588 \$93 \$92 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$589 VSSD clks \$93 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$590 \$91 \$155 \$93 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$591 \$95 \$155 \$92 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$592 \$96 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$593 VSSD \$95 \$96 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$594 \$94 \$96 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$595 VSSD Set \$94 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$596 \$95 \$154 \$94 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$597 \$97 \$157 \$96 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$598 \$98 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$599 VSSD \$97 \$98 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$600 \$99 \$98 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$601 VSSD clks \$99 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$602 \$97 \$158 \$99 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$603 \$101 \$158 \$98 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$604 CK9 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$605 VSSD \$101 CK9 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$606 \$100 CK9 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$607 VSSD Set \$100 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$608 \$101 \$157 \$100 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$609 \$103 \$160 CK9 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$610 \$104 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$611 VSSD \$103 \$104 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$612 \$105 \$104 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$613 VSSD clks \$105 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$614 \$103 \$161 \$105 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$615 \$107 \$161 \$104 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$616 CK8 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$617 VSSD \$107 CK8 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$618 \$106 CK8 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$619 VSSD Set \$106 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$620 \$107 \$160 \$106 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$621 \$109 \$163 CK8 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$622 \$110 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$623 VSSD \$109 \$110 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$624 \$111 \$110 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$625 VSSD clks \$111 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$626 \$109 \$164 \$111 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$627 \$113 \$164 \$110 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$628 CK7 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$629 VSSD \$113 CK7 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$630 \$112 CK7 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$631 VSSD Set \$112 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$632 \$113 \$163 \$112 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$633 \$115 \$166 CK7 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$634 \$116 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$635 VSSD \$115 \$116 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$636 \$117 \$116 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$637 VSSD clks \$117 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$638 \$115 \$167 \$117 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$639 \$119 \$167 \$116 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$640 CK6 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$641 VSSD \$119 CK6 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$642 \$118 CK6 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$643 VSSD Set \$118 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$644 \$119 \$166 \$118 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$645 \$121 \$169 CK6 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$646 \$122 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$647 VSSD \$121 \$122 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$648 \$123 \$122 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$649 VSSD clks \$123 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$650 \$121 \$170 \$123 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$651 \$125 \$170 \$122 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$652 CK5 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$653 VSSD \$125 CK5 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$654 \$124 CK5 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$655 VSSD Set \$124 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$656 \$125 \$169 \$124 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$657 \$127 \$172 CK5 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$658 \$128 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$659 VSSD \$127 \$128 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$660 \$129 \$128 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$661 VSSD clks \$129 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$662 \$127 \$173 \$129 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$663 \$131 \$173 \$128 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$664 CK4 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$665 VSSD \$131 CK4 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$666 \$130 CK4 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$667 VSSD Set \$130 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$668 \$131 \$172 \$130 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$669 \$133 \$175 CK4 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$670 \$134 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$671 VSSD \$133 \$134 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$672 \$135 \$134 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$673 VSSD clks \$135 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$674 \$133 \$176 \$135 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$675 \$137 \$176 \$134 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$676 CK3 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$677 VSSD \$137 CK3 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$678 \$136 CK3 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$679 VSSD Set \$136 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$680 \$137 \$175 \$136 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$681 \$139 \$178 CK3 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$682 \$140 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$683 VSSD \$139 \$140 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$684 \$141 \$140 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$685 VSSD clks \$141 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$686 \$139 \$179 \$141 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$687 \$143 \$179 \$140 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$688 CK2 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$689 VSSD \$143 CK2 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$690 \$142 CK2 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$691 VSSD Set \$142 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$692 \$143 \$178 \$142 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$693 \$145 \$181 CK2 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$694 \$146 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$695 VSSD \$145 \$146 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$696 \$147 \$146 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$697 VSSD clks \$147 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$698 \$145 \$182 \$147 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$699 \$150 \$182 \$146 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$700 CK1 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$701 VSSD \$150 CK1 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$702 \$149 CK1 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$703 VSSD Set \$149 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$704 \$150 \$181 \$149 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$705 \$151 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$706 \$152 \$151 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$707 \$153 CK11 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$708 \$154 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$709 \$155 \$154 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$710 Bit_0 \$1632 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$711 \$1632 \$1631 \$1635 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$712 VSSD \$1806 \$1632 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$713 \$1633 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$714 \$1634 \$1633 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$715 \$2421 \$2557 \$2376 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$716 \$156 \$96 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$717 \$2421 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$718 \$1600 \$1633 \$1635 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$719 \$157 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$720 VSSD \$1635 \$2421 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$721 \$1601 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$722 \$158 \$157 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$723 VSSD \$1600 \$1601 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$724 \$1635 \$2376 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$725 VSSD Reset \$1635 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$726 \$1602 \$1601 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$727 VSSD Reset \$1602 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$728 \$2422 \$2558 \$2376 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$729 \$1600 \$1634 \$1602 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$730 \$2423 \$2558 \$2411 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$731 \$1605 \$1634 \$1601 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$732 \$2423 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$733 VSSD \$2422 \$2423 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$734 \$1603 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$735 VSSD \$1605 \$1603 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$736 \$2422 \$2411 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$737 VSSD Set \$2422 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$738 \$1604 \$1603 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$739 D_C_1 \$2557 \$2411 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$740 VSSD Set \$1604 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$741 \$1605 \$1633 \$1604 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$742 \$1636 \$1603 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$743 \$159 CK9 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$744 \$160 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$745 \$161 \$160 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$746 Bit_1 \$1606 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$747 \$1606 \$1637 \$1640 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$748 VSSD \$1820 \$1606 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$749 \$162 CK8 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$750 \$1638 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$751 \$163 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$752 \$1639 \$1638 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$753 \$2425 \$2559 \$2377 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$754 \$164 \$163 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$755 \$2425 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$756 \$1607 \$1638 \$1640 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$757 VSSD \$1640 \$2425 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$758 \$1608 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$759 VSSD \$1607 \$1608 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$760 \$1640 \$2377 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$761 VSSD Reset \$1640 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$762 \$1609 \$1608 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$763 VSSD Reset \$1609 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$764 \$2426 \$2560 \$2377 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$765 \$1607 \$1639 \$1609 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$766 \$2427 \$2560 \$2412 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$767 \$1612 \$1639 \$1608 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$768 \$2427 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$769 VSSD \$2426 \$2427 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$770 \$1610 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$771 VSSD \$1612 \$1610 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$772 \$2426 \$2412 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$773 VSSD Set \$2426 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$774 \$1611 \$1610 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$775 D_C_2 \$2559 \$2412 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$776 VSSD Set \$1611 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$777 \$1612 \$1638 \$1611 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$778 \$1641 \$1610 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$779 \$165 CK7 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$780 \$166 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$781 \$167 \$166 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$782 Bit_2 \$1643 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$783 \$168 CK6 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$784 \$1643 \$1642 \$1646 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$785 VSSD \$1833 \$1643 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$786 \$169 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$787 \$170 \$169 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$788 \$1644 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$789 \$1645 \$1644 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$790 \$2429 \$2561 \$2378 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$791 \$2429 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$792 \$1613 \$1644 \$1646 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$793 VSSD \$1646 \$2429 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$794 \$1614 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$795 VSSD \$1613 \$1614 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$796 \$1646 \$2378 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$797 VSSD Reset \$1646 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$798 \$1615 \$1614 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$799 VSSD Reset \$1615 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$800 \$2430 \$2562 \$2378 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$801 \$1613 \$1645 \$1615 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$802 \$2431 \$2562 \$2413 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$803 \$1618 \$1645 \$1614 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$804 \$2431 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$805 VSSD \$2430 \$2431 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$806 \$1616 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$807 VSSD \$1618 \$1616 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$808 \$2430 \$2413 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$809 VSSD Set \$2430 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$810 \$1617 \$1616 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$811 D_C_3 \$2561 \$2413 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$812 VSSD Set \$1617 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$813 \$171 CK5 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$814 \$1618 \$1644 \$1617 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$815 \$172 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$816 \$1647 \$1616 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$817 \$173 \$172 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$818 \$174 CK4 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$819 Bit_3 \$1619 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$820 \$175 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$821 \$176 \$175 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$822 \$1619 \$1648 \$1651 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$823 VSSD \$1846 \$1619 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$824 \$1649 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$825 \$1650 \$1649 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$826 \$2433 \$2563 \$2379 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$827 \$2433 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$828 \$1620 \$1649 \$1651 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$829 VSSD \$1651 \$2433 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$830 \$1621 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$831 VSSD \$1620 \$1621 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$832 \$1651 \$2379 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$833 VSSD Reset \$1651 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$834 \$1622 \$1621 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$835 VSSD Reset \$1622 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$836 \$2434 \$2564 \$2379 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$837 \$1620 \$1650 \$1622 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$838 \$2435 \$2564 \$2414 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$839 \$1652 \$1650 \$1621 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$840 \$2435 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$841 VSSD \$2434 \$2435 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$842 \$1623 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$843 VSSD \$1652 \$1623 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$844 \$2434 \$2414 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$845 \$177 CK3 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$846 VSSD Set \$2434 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$847 \$1624 \$1623 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$848 D_C_4 \$2563 \$2414 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$849 VSSD Set \$1624 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$850 \$178 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$851 \$179 \$178 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$852 \$1652 \$1649 \$1624 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$853 \$1653 \$1623 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$854 \$180 CK2 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$855 \$181 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$856 \$182 \$181 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$857 Bit_4 \$1625 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$858 \$1625 \$1654 \$1657 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$859 VSSD \$1859 \$1625 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$860 \$1655 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$861 \$1656 \$1655 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$862 \$2437 \$2565 \$2380 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$863 \$2437 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$864 \$1626 \$1655 \$1657 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$865 VSSD \$1657 \$2437 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$866 \$1627 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$867 VSSD \$1626 \$1627 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$868 \$1657 \$2380 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$869 VSSD Reset \$1657 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$870 \$1628 \$1627 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$871 VSSD Reset \$1628 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$872 \$2438 \$2566 \$2380 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$873 \$1626 \$1656 \$1628 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$874 \$2439 \$2566 \$2415 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$875 \$1658 \$1656 \$1627 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$876 \$183 CK1 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$877 \$2439 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$878 VSSD \$2438 \$2439 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$879 \$1629 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$880 VSSD \$1658 \$1629 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$881 \$2438 \$2415 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$882 VSSD Set \$2438 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$883 \$1630 \$1629 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$884 D_C_5 \$2565 \$2415 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$885 VSSD Set \$1630 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$886 \$1658 \$1655 \$1630 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$887 \$1659 \$1629 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$888 \$3398 \$3579 \$3331 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$889 \$3398 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$890 VSSD \$3580 \$3398 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$891 \$3580 \$3331 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$892 VSSD Reset \$3580 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$893 \$3399 \$3605 \$3331 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$894 \$3369 \$3605 \$3362 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$895 \$3369 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$896 VSSD \$3399 \$3369 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$897 \$3399 \$3362 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$898 VSSD Set \$3399 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$899 \$3370 \$3579 \$3362 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$900 \$3371 \$3400 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$901 \$3370 \$3614 \$3371 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$902 VSSD \$3371 Bit_10 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$903 Bit_0 \$1806 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$904 \$2442 \$1631 \$1635 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$905 \$3373 \$3581 \$3332 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$906 VSSD \$1635 \$2443 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$907 \$3373 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$908 VSSD \$3582 \$3373 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$909 \$3582 \$3332 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$910 VSSD Reset \$3582 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$911 \$3402 \$3627 \$3332 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$912 \$3374 \$3627 \$3363 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$913 \$3374 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$914 VSSD \$3402 \$3374 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$915 \$3402 \$3363 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$916 VSSD Set \$3402 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$917 \$3375 \$3581 \$3363 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$918 VSSD \$2557 \$2558 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$919 \$3376 \$3403 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$920 VSSD \$1631 \$2557 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$921 \$3375 \$3628 \$3376 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$922 VSSD \$1806 \$1631 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$923 VSSD \$3376 Bit_9 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$924 VSSD CK1 \$1806 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$925 Bit_1 \$1820 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$926 \$2444 \$1637 \$1640 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$927 \$3378 \$3583 \$3333 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$928 VSSD \$1640 \$2445 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$929 \$3378 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$930 VSSD \$3584 \$3378 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$931 \$3584 \$3333 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$932 VSSD Reset \$3584 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$933 \$3379 \$3641 \$3333 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$934 \$3380 \$3641 \$3364 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$935 \$3380 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$936 VSSD \$3379 \$3380 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$937 \$3379 \$3364 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$938 VSSD Set \$3379 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$939 \$3405 \$3583 \$3364 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$940 VSSD \$2559 \$2560 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$941 \$3407 \$3406 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$942 VSSD \$1637 \$2559 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$943 \$3405 \$3642 \$3407 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$944 VSSD \$1820 \$1637 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$945 VSSD \$3407 Bit_8 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$946 VSSD CK2 \$1820 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$947 Bit_2 \$1833 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$948 \$2446 \$1642 \$1646 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$949 \$3382 \$3585 \$3334 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$950 VSSD \$1646 \$2447 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$951 \$3382 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$952 VSSD \$3586 \$3382 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$953 \$3586 \$3334 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$954 VSSD Reset \$3586 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$955 \$3409 \$3655 \$3334 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$956 \$3383 \$3655 \$3365 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$957 \$3383 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$958 VSSD \$3409 \$3383 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$959 \$3409 \$3365 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$960 VSSD Set \$3409 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$961 \$3384 \$3585 \$3365 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$962 VSSD \$2561 \$2562 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$963 \$3385 \$3410 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$964 VSSD \$1642 \$2561 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$965 \$3384 \$3656 \$3385 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$966 VSSD \$1833 \$1642 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$967 VSSD \$3385 Bit_7 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$968 VSSD CK3 \$1833 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$969 Bit_3 \$1846 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$970 \$2448 \$1648 \$1651 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$971 \$3387 \$3587 \$3335 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$972 VSSD \$1651 \$2449 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$973 \$3387 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$974 VSSD \$3588 \$3387 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$975 \$3588 \$3335 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$976 VSSD Reset \$3588 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$977 \$3388 \$3669 \$3335 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$978 \$3389 \$3669 \$3366 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$979 \$3389 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$980 VSSD \$3388 \$3389 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$981 \$3388 \$3366 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$982 VSSD Set \$3388 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$983 \$3412 \$3587 \$3366 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$984 VSSD \$2563 \$2564 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$985 \$3390 \$3413 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$986 VSSD \$1648 \$2563 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$987 \$3412 \$3670 \$3390 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$988 VSSD \$1846 \$1648 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$989 VSSD \$3390 Bit_6 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$990 VSSD CK4 \$1846 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$991 Bit_4 \$1859 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$992 \$2450 \$1654 \$1657 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$993 \$3392 \$3589 \$3336 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$994 VSSD \$1657 \$2451 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$995 \$3392 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$996 VSSD \$3590 \$3392 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$997 \$3590 \$3336 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$998 VSSD Reset \$3590 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$999 \$3415 \$3683 \$3336 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1000 \$3393 \$3683 \$3367 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1001 \$3393 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1002 VSSD \$3415 \$3393 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1003 \$3415 \$3367 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1004 VSSD Set \$3415 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1005 \$3394 \$3589 \$3367 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1006 VSSD \$2565 \$2566 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1007 \$3395 \$3416 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1008 VSSD \$1654 \$2565 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1009 \$3394 \$3684 \$3395 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1010 VSSD \$1859 \$1654 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1011 VSSD \$3395 Bit_5 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1012 VSSD CK5 \$1859 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1013 VSSD \$3580 \$3397 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1014 \$4341 \$4383 D_C_11 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1015 \$4342 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1016 VSSD \$4341 \$4342 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1017 \$4343 \$4342 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1018 VSSD Reset \$4343 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1019 \$4341 \$4384 \$4343 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1020 \$4345 \$4384 \$4342 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1021 \$3370 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1022 VSSD \$4345 \$3370 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1023 \$4344 \$3370 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1024 VSSD Set \$4344 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1025 \$4345 \$4383 \$4344 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1026 VSSD \$3579 \$3605 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1027 VSSD clks \$3579 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1028 VSSD \$3582 \$3401 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1029 \$4347 \$4386 D_C_10 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1030 \$4348 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1031 VSSD \$4347 \$4348 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1032 \$4349 \$4348 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1033 VSSD Reset \$4349 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1034 \$4347 \$4387 \$4349 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1035 \$4351 \$4387 \$4348 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1036 \$3375 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1037 VSSD \$4351 \$3375 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1038 \$4350 \$3375 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1039 VSSD Set \$4350 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1040 \$4351 \$4386 \$4350 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1041 VSSD \$3581 \$3627 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1042 VSSD clks \$3581 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1043 VSSD \$3584 \$3404 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1044 \$4353 \$4389 D_C_9 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1045 \$4354 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1046 VSSD \$4353 \$4354 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1047 \$4355 \$4354 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1048 VSSD Reset \$4355 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1049 \$4353 \$4390 \$4355 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1050 \$4357 \$4390 \$4354 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1051 \$3405 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1052 VSSD \$4357 \$3405 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1053 \$4356 \$3405 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1054 VSSD Set \$4356 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1055 \$4357 \$4389 \$4356 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1056 VSSD \$3583 \$3641 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1057 VSSD clks \$3583 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1058 VSSD \$3586 \$3408 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1059 \$4359 \$4392 D_C_8 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1060 \$4360 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1061 VSSD \$4359 \$4360 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1062 \$4361 \$4360 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1063 VSSD Reset \$4361 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1064 \$4359 \$4393 \$4361 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1065 \$4363 \$4393 \$4360 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1066 \$3384 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1067 VSSD \$4363 \$3384 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1068 \$4362 \$3384 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1069 VSSD Set \$4362 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1070 \$4363 \$4392 \$4362 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1071 VSSD \$3585 \$3655 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1072 VSSD clks \$3585 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1073 VSSD \$3588 \$3411 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1074 \$4365 \$4395 D_C_7 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1075 \$4366 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1076 VSSD \$4365 \$4366 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1077 \$4367 \$4366 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1078 VSSD Reset \$4367 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1079 \$4365 \$4396 \$4367 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1080 \$4369 \$4396 \$4366 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1081 \$3412 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1082 VSSD \$4369 \$3412 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1083 \$4368 \$3412 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1084 VSSD Set \$4368 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1085 \$4369 \$4395 \$4368 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1086 VSSD \$3587 \$3669 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1087 VSSD clks \$3587 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1088 VSSD \$3590 \$3414 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1089 \$4371 \$4398 D_C_6 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1090 \$4372 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1091 VSSD \$4371 \$4372 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1092 \$4373 \$4372 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1093 VSSD Reset \$4373 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1094 \$4371 \$4399 \$4373 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1095 \$4375 \$4399 \$4372 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1096 \$3394 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1097 VSSD \$4375 \$3394 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1098 \$4374 \$3394 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1099 VSSD Set \$4374 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1100 \$4375 \$4398 \$4374 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1101 VSSD \$3589 \$3683 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1102 VSSD clks \$3589 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1103 \$3400 CK11 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1104 \$3614 \$3400 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1105 \$4383 \$3614 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1106 \$4384 \$4383 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1107 \$4385 \$3370 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1108 \$3370 \$3614 \$4346 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1109 VCM \$3400 Bit_10 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1110 \$3403 \$96 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1111 \$3628 \$3403 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1112 \$4386 \$3628 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1113 \$4387 \$4386 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1114 \$4388 \$3375 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1115 \$3375 \$3628 \$4352 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1116 VCM \$3403 Bit_9 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1117 \$3406 CK9 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1118 \$3642 \$3406 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1119 \$4389 \$3642 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1120 \$4390 \$4389 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1121 \$4391 \$3405 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1122 \$3405 \$3642 \$4358 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1123 VCM \$3406 Bit_8 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1124 \$3410 CK8 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1125 \$3656 \$3410 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1126 \$4392 \$3656 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1127 \$4393 \$4392 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1128 \$4394 \$3384 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1129 \$3384 \$3656 \$4364 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1130 VCM \$3410 Bit_7 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1131 \$3413 CK7 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1132 \$3670 \$3413 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1133 \$4395 \$3670 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1134 \$4396 \$4395 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1135 \$4397 \$3412 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1136 \$3412 \$3670 \$4370 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1137 VCM \$3413 Bit_6 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1138 \$3416 CK6 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1139 \$3684 \$3416 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1140 \$4398 \$3684 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1141 \$4399 \$4398 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1142 \$4400 \$3394 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1143 \$3394 \$3684 \$4376 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1144 VCM \$3416 Bit_5 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
.ENDS SAR_Asynchronous_top
