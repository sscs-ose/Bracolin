* Extracted by KLayout with GF180MCU LVS runset on : 21/12/2023 23:00

.SUBCKT PRbiased_net_x5 ITP5 ITP4 ITP3 ITP2 ITP1 ITN1 ITN2 ITN3 ITN4 ITN5 IBN1
+ IBN2 IBN3 IBN4 IBN5 VDD VA VB IBP1 IBP2 IBP3 IBP4 IBP5 VSS
M$1 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$4 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$5 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$6 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$7 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$8 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$9 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$10 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$11 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$12 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$13 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$14 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$15 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$16 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$17 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$18 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$19 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$20 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$21 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$22 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$23 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$24 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$25 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$26 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$27 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$28 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$29 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$30 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$31 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$32 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$33 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$34 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$35 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$36 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$37 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$38 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$39 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$40 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$41 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$42 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$43 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$44 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$45 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$46 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$47 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$48 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$49 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$50 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$51 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$52 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$53 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$54 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$55 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$56 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$57 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$58 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$59 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$60 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$61 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$62 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$63 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$64 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$65 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$66 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$67 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$68 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$69 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$70 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$71 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$72 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$73 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$74 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$75 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$76 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$77 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$78 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$79 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$80 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$81 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$82 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$83 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$84 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$85 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$86 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$87 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$88 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$89 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$90 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$91 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$92 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$93 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$94 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$95 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$96 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$97 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$98 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$99 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$100 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$101 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$102 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$103 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$104 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$105 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$106 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$107 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$108 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$109 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$110 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$111 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$112 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$113 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$114 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$115 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$116 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$117 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$118 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$119 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$120 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$121 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$122 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$123 \$893 \$147 \$147 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$124 VDD \$147 \$893 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$125 \$894 \$147 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$126 \$47 \$147 \$894 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$127 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$128 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$129 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$130 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$131 \$896 \$929 VA VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$132 \$150 \$929 \$896 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$133 \$897 \$929 \$258 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$134 \$898 \$929 \$897 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$135 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$136 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$137 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$138 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$139 \$899 \$187 \$188 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$140 ITP1 \$187 \$899 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$141 \$900 IBP1 ITP1 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$142 \$929 IBP1 \$900 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$143 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$144 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$145 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$146 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$147 \$901 \$155 \$155 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$148 VDD \$155 \$901 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$149 \$902 \$155 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$150 \$48 \$155 \$902 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$151 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$152 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$153 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$154 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$155 \$903 \$930 \$898 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$156 \$158 \$930 \$903 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$157 \$904 \$930 \$260 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$158 \$905 \$930 \$904 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$159 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$160 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$161 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$162 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$163 \$906 \$189 \$190 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$164 ITP2 \$189 \$906 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$165 \$907 IBP2 ITP2 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$166 \$930 IBP2 \$907 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$167 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$168 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$169 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$170 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$171 \$908 \$163 \$163 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$172 VDD \$163 \$908 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$173 \$909 \$163 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$174 \$49 \$163 \$909 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$175 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$176 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$177 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$178 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$179 \$910 \$931 \$905 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$180 \$166 \$931 \$910 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$181 \$911 \$931 \$262 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$182 \$912 \$931 \$911 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$183 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$184 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$185 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$186 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$187 \$913 \$191 \$192 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$188 ITP3 \$191 \$913 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$189 \$914 IBP3 ITP3 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$190 \$931 IBP3 \$914 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$191 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$192 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$193 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$194 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$195 \$915 \$171 \$171 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$196 VDD \$171 \$915 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$197 \$916 \$171 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$198 \$50 \$171 \$916 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$199 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$200 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$201 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$202 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$203 \$917 \$932 \$912 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$204 \$174 \$932 \$917 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$205 \$918 \$932 \$264 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$206 \$919 \$932 \$918 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$207 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$208 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$209 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$210 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$211 \$920 \$193 \$194 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$212 ITP4 \$193 \$920 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$213 \$921 IBP4 ITP4 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$214 \$932 IBP4 \$921 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$215 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$216 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$217 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$218 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$219 \$922 \$179 \$179 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$220 VDD \$179 \$922 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$221 \$923 \$179 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$222 \$51 \$179 \$923 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$223 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$224 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$225 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$226 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$227 \$924 \$933 \$919 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$228 \$182 \$933 \$924 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$229 \$925 \$933 \$266 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$230 VB \$933 \$925 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$231 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$232 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$233 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$234 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$235 \$927 \$195 \$196 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$236 ITP5 \$195 \$927 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$237 \$928 IBP5 ITP5 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$238 \$933 IBP5 \$928 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$239 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$240 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$241 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$242 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$243 \$1054 \$147 \$47 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$244 VDD \$147 \$1054 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$245 \$1055 \$147 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$246 \$147 \$147 \$1055 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$247 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$248 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$249 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$250 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$251 \$1056 \$929 IBP1 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$252 VSS \$929 \$1056 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$253 \$1057 \$929 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$254 IBP1 \$929 \$1057 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$255 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$256 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$257 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$258 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$259 \$1058 IBP1 \$929 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$260 ITP1 IBP1 \$1058 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$261 \$1059 \$187 ITP1 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$262 \$188 \$187 \$1059 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$263 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$264 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$265 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$266 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$267 \$1060 \$155 \$48 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$268 VDD \$155 \$1060 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$269 \$1061 \$155 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$270 \$155 \$155 \$1061 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$271 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$272 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$273 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$274 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$275 \$1062 \$930 IBP2 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$276 VSS \$930 \$1062 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$277 \$1063 \$930 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$278 IBP2 \$930 \$1063 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$279 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$280 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$281 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$282 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$283 \$1064 IBP2 \$930 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$284 ITP2 IBP2 \$1064 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$285 \$1065 \$189 ITP2 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$286 \$190 \$189 \$1065 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$287 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$288 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$289 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$290 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$291 \$1066 \$163 \$49 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$292 VDD \$163 \$1066 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$293 \$1067 \$163 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$294 \$163 \$163 \$1067 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$295 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$296 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$297 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$298 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$299 \$1068 \$931 IBP3 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$300 VSS \$931 \$1068 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$301 \$1069 \$931 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$302 IBP3 \$931 \$1069 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$303 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$304 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$305 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$306 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$307 \$1070 IBP3 \$931 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$308 ITP3 IBP3 \$1070 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$309 \$1071 \$191 ITP3 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$310 \$192 \$191 \$1071 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$311 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$312 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$313 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$314 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$315 \$1072 \$171 \$50 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$316 VDD \$171 \$1072 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$317 \$1073 \$171 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$318 \$171 \$171 \$1073 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$319 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$320 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$321 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$322 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$323 \$1074 \$932 IBP4 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$324 VSS \$932 \$1074 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$325 \$1075 \$932 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$326 IBP4 \$932 \$1075 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$327 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$328 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$329 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$330 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$331 \$1076 IBP4 \$932 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$332 ITP4 IBP4 \$1076 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$333 \$1077 \$193 ITP4 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$334 \$194 \$193 \$1077 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$335 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$336 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$337 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$338 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$339 \$1078 \$179 \$51 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$340 VDD \$179 \$1078 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$341 \$1079 \$179 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$342 \$179 \$179 \$1079 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$343 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$344 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$345 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$346 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$347 \$1080 \$933 IBP5 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$348 VSS \$933 \$1080 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$349 \$1081 \$933 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$350 IBP5 \$933 \$1081 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$351 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$352 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$353 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$354 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$355 \$1082 IBP5 \$933 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$356 ITP5 IBP5 \$1082 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$357 \$1083 \$195 ITP5 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$358 \$196 \$195 \$1083 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$359 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$360 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$361 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$362 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$363 \$1189 \$147 \$147 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$364 VDD \$147 \$1189 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$365 \$1190 \$147 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$366 \$47 \$147 \$1190 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$367 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$368 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$369 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$370 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$371 \$1191 \$929 IBP1 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$372 VSS \$929 \$1191 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$373 \$1192 \$929 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$374 IBP1 \$929 \$1192 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$375 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$376 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$377 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$378 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$379 \$1193 \$187 \$188 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$380 ITP1 \$187 \$1193 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$381 \$1194 IBP1 ITP1 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$382 \$929 IBP1 \$1194 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$383 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$384 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$385 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$386 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$387 \$1195 \$155 \$155 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$388 VDD \$155 \$1195 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$389 \$1196 \$155 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$390 \$48 \$155 \$1196 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$391 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$392 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$393 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$394 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$395 \$1197 \$930 IBP2 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$396 VSS \$930 \$1197 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$397 \$1198 \$930 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$398 IBP2 \$930 \$1198 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$399 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$400 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$401 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$402 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$403 \$1199 \$189 \$190 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$404 ITP2 \$189 \$1199 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$405 \$1200 IBP2 ITP2 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$406 \$930 IBP2 \$1200 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$407 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$408 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$409 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$410 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$411 \$1201 \$163 \$163 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$412 VDD \$163 \$1201 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$413 \$1202 \$163 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$414 \$49 \$163 \$1202 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$415 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$416 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$417 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$418 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$419 \$1203 \$931 IBP3 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$420 VSS \$931 \$1203 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$421 \$1204 \$931 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$422 IBP3 \$931 \$1204 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$423 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$424 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$425 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$426 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$427 \$1205 \$191 \$192 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$428 ITP3 \$191 \$1205 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$429 \$1206 IBP3 ITP3 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$430 \$931 IBP3 \$1206 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$431 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$432 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$433 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$434 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$435 \$1207 \$171 \$171 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$436 VDD \$171 \$1207 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$437 \$1208 \$171 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$438 \$50 \$171 \$1208 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$439 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$440 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$441 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$442 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$443 \$1209 \$932 IBP4 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$444 VSS \$932 \$1209 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$445 \$1210 \$932 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$446 IBP4 \$932 \$1210 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$447 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$448 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$449 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$450 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$451 \$1211 \$193 \$194 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$452 ITP4 \$193 \$1211 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$453 \$1212 IBP4 ITP4 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$454 \$932 IBP4 \$1212 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$455 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$456 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$457 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$458 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$459 \$1213 \$179 \$179 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$460 VDD \$179 \$1213 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$461 \$1214 \$179 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$462 \$51 \$179 \$1214 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$463 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$464 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$465 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$466 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$467 \$1215 \$933 IBP5 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$468 VSS \$933 \$1215 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$469 \$1216 \$933 VSS VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$470 IBP5 \$933 \$1216 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$471 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$472 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$473 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$474 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$475 \$1217 \$195 \$196 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$476 ITP5 \$195 \$1217 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$477 \$1218 IBP5 ITP5 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$478 \$933 IBP5 \$1218 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$479 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$480 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$481 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$482 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$483 \$1349 \$147 \$47 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$484 VDD \$147 \$1349 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$485 \$1350 \$147 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$486 \$147 \$147 \$1350 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$487 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$488 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$489 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$490 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$491 \$1351 \$929 \$898 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$492 \$258 \$929 \$1351 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$493 \$1352 \$929 \$150 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$494 VA \$929 \$1352 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$495 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$496 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$497 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$498 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$499 \$1353 IBP1 \$929 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$500 ITP1 IBP1 \$1353 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$501 \$1354 \$187 ITP1 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$502 \$188 \$187 \$1354 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$503 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$504 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$505 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$506 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$507 \$1355 \$155 \$48 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$508 VDD \$155 \$1355 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$509 \$1356 \$155 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$510 \$155 \$155 \$1356 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$511 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$512 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$513 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$514 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$515 \$1357 \$930 \$905 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$516 \$260 \$930 \$1357 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$517 \$1358 \$930 \$158 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$518 \$898 \$930 \$1358 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$519 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$520 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$521 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$522 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$523 \$1359 IBP2 \$930 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$524 ITP2 IBP2 \$1359 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$525 \$1360 \$189 ITP2 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$526 \$190 \$189 \$1360 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$527 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$528 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$529 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$530 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$531 \$1361 \$163 \$49 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$532 VDD \$163 \$1361 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$533 \$1362 \$163 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$534 \$163 \$163 \$1362 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$535 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$536 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$537 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$538 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$539 \$1363 \$931 \$912 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$540 \$262 \$931 \$1363 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$541 \$1364 \$931 \$166 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$542 \$905 \$931 \$1364 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$543 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$544 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$545 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$546 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$547 \$1365 IBP3 \$931 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$548 ITP3 IBP3 \$1365 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$549 \$1366 \$191 ITP3 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$550 \$192 \$191 \$1366 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$551 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$552 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$553 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$554 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$555 \$1367 \$171 \$50 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$556 VDD \$171 \$1367 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$557 \$1368 \$171 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$558 \$171 \$171 \$1368 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$559 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$560 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$561 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$562 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$563 \$1369 \$932 \$919 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$564 \$264 \$932 \$1369 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$565 \$1370 \$932 \$174 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$566 \$912 \$932 \$1370 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$567 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$568 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$569 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$570 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$571 \$1371 IBP4 \$932 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$572 ITP4 IBP4 \$1371 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$573 \$1372 \$193 ITP4 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$574 \$194 \$193 \$1372 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$575 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$576 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$577 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$578 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$579 \$1373 \$179 \$51 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$580 VDD \$179 \$1373 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$581 \$1374 \$179 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$582 \$179 \$179 \$1374 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$583 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$584 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$585 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$586 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$587 \$1375 \$933 VB VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$588 \$266 \$933 \$1375 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$589 \$1376 \$933 \$182 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$590 \$919 \$933 \$1376 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$591 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$592 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$593 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$594 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$595 \$1377 IBP5 \$933 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$596 ITP5 IBP5 \$1377 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$597 \$1378 \$195 ITP5 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$598 \$196 \$195 \$1378 VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$599 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$600 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$601 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$602 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$603 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$604 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$605 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$606 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$607 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$608 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$609 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$610 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$611 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$612 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$613 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$614 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$615 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$616 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$617 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$618 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$619 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$620 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$621 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$622 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$623 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$624 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$625 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$626 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$627 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$628 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$629 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$630 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$631 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$632 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$633 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$634 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$635 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$636 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$637 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$638 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$639 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$640 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$641 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$642 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$643 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$644 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$645 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$646 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$647 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$648 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$649 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$650 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$651 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$652 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$653 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$654 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$655 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$656 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$657 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$658 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$659 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$660 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$661 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$662 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$663 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$664 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$665 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$666 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$667 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$668 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$669 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$670 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$671 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$672 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$673 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$674 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$675 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$676 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$677 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$678 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$679 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$680 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$681 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$682 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$683 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$684 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$685 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$686 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$687 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$688 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$689 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$690 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$691 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$692 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$693 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$694 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$695 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$696 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$697 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$698 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$699 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$700 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$701 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$702 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$703 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$704 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$705 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$706 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$707 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$708 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$709 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$710 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$711 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$712 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$713 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$714 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$715 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$716 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$717 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$718 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$719 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$720 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$721 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$722 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$723 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$724 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$725 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$726 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$727 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$728 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$729 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$730 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$731 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$732 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$733 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$734 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$735 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$736 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$737 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$738 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$739 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$740 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$741 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$742 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$743 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$744 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$745 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$746 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$747 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$748 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$749 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$750 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$751 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$752 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$753 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$754 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$755 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$756 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$757 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$758 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$759 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$760 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$761 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$762 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$763 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$764 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$765 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$766 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$767 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$768 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$769 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$770 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$771 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$772 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$773 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$774 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$775 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$776 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$777 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$778 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$779 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$780 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$781 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$782 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$783 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$784 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$785 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$786 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$787 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$788 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$789 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$790 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$791 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$792 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$793 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$794 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$795 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$796 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$797 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$798 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$799 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$800 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$801 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$802 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$803 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$804 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$805 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$806 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$807 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$808 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$809 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$810 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$811 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$812 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$813 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$814 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$815 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$816 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$817 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$818 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$819 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$820 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$821 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$822 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$823 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$824 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$825 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$826 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$827 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$828 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$829 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$830 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$831 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$832 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$833 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$834 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$835 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$836 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$837 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$838 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$839 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$840 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$841 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$842 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$843 \$148 \$187 \$147 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$844 ITN1 \$187 \$148 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$845 \$149 IBN1 ITN1 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$846 \$47 IBN1 \$149 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$847 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$848 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$849 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$850 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$851 \$151 \$47 \$150 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$852 \$187 \$47 \$151 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$853 \$152 \$47 \$187 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$854 \$258 \$47 \$152 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$855 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$856 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$857 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$858 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$859 \$153 \$188 \$188 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$860 VSS \$188 \$153 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$861 \$154 \$188 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$862 \$929 \$188 \$154 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$863 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$864 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$865 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$866 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$867 \$156 \$189 \$155 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$868 ITN2 \$189 \$156 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$869 \$157 IBN2 ITN2 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$870 \$48 IBN2 \$157 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$871 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$872 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$873 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$874 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$875 \$159 \$48 \$158 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$876 \$189 \$48 \$159 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$877 \$160 \$48 \$189 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$878 \$260 \$48 \$160 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$879 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$880 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$881 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$882 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$883 \$161 \$190 \$190 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$884 VSS \$190 \$161 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$885 \$162 \$190 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$886 \$930 \$190 \$162 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$887 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$888 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$889 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$890 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$891 \$164 \$191 \$163 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$892 ITN3 \$191 \$164 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$893 \$165 IBN3 ITN3 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$894 \$49 IBN3 \$165 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$895 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$896 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$897 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$898 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$899 \$167 \$49 \$166 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$900 \$191 \$49 \$167 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$901 \$168 \$49 \$191 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$902 \$262 \$49 \$168 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$903 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$904 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$905 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$906 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$907 \$169 \$192 \$192 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$908 VSS \$192 \$169 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$909 \$170 \$192 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$910 \$931 \$192 \$170 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$911 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$912 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$913 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$914 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$915 \$172 \$193 \$171 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$916 ITN4 \$193 \$172 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$917 \$173 IBN4 ITN4 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$918 \$50 IBN4 \$173 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$919 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$920 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$921 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$922 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$923 \$175 \$50 \$174 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$924 \$193 \$50 \$175 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$925 \$176 \$50 \$193 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$926 \$264 \$50 \$176 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$927 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$928 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$929 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$930 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$931 \$177 \$194 \$194 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$932 VSS \$194 \$177 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$933 \$178 \$194 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$934 \$932 \$194 \$178 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$935 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$936 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$937 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$938 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$939 \$180 \$195 \$179 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$940 ITN5 \$195 \$180 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$941 \$181 IBN5 ITN5 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$942 \$51 IBN5 \$181 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$943 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$944 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$945 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$946 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$947 \$183 \$51 \$182 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$948 \$195 \$51 \$183 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$949 \$184 \$51 \$195 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$950 \$266 \$51 \$184 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$951 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$952 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$953 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$954 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$955 \$185 \$196 \$196 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$956 VSS \$196 \$185 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$957 \$186 \$196 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$958 \$933 \$196 \$186 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$959 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$960 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$961 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$962 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$963 \$337 IBN1 \$47 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$964 ITN1 IBN1 \$337 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$965 \$338 \$187 ITN1 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$966 \$147 \$187 \$338 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$967 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$968 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$969 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$970 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$971 \$339 \$47 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$972 IBN1 \$47 \$339 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$973 \$340 \$47 IBN1 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$974 VDD \$47 \$340 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$975 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$976 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$977 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$978 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$979 \$341 \$188 \$929 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$980 VSS \$188 \$341 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$981 \$342 \$188 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$982 \$188 \$188 \$342 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$983 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$984 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$985 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$986 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$987 \$343 IBN2 \$48 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$988 ITN2 IBN2 \$343 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$989 \$344 \$189 ITN2 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$990 \$155 \$189 \$344 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$991 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$992 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$993 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$994 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$995 \$345 \$48 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$996 IBN2 \$48 \$345 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$997 \$346 \$48 IBN2 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$998 VDD \$48 \$346 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$999 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1000 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1001 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1002 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1003 \$347 \$190 \$930 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1004 VSS \$190 \$347 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1005 \$348 \$190 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1006 \$190 \$190 \$348 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1007 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1008 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1009 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1010 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1011 \$349 IBN3 \$49 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1012 ITN3 IBN3 \$349 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1013 \$350 \$191 ITN3 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1014 \$163 \$191 \$350 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1015 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1016 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1017 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1018 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1019 \$351 \$49 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1020 IBN3 \$49 \$351 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1021 \$352 \$49 IBN3 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1022 VDD \$49 \$352 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1023 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1024 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1025 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1026 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1027 \$353 \$192 \$931 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1028 VSS \$192 \$353 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1029 \$354 \$192 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1030 \$192 \$192 \$354 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1031 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1032 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1033 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1034 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1035 \$355 IBN4 \$50 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1036 ITN4 IBN4 \$355 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1037 \$356 \$193 ITN4 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1038 \$171 \$193 \$356 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1039 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1040 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1041 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1042 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1043 \$357 \$50 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1044 IBN4 \$50 \$357 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1045 \$358 \$50 IBN4 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1046 VDD \$50 \$358 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1047 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1048 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1049 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1050 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1051 \$359 \$194 \$932 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1052 VSS \$194 \$359 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1053 \$360 \$194 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1054 \$194 \$194 \$360 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1055 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1056 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1057 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1058 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1059 \$361 IBN5 \$51 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1060 ITN5 IBN5 \$361 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1061 \$362 \$195 ITN5 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1062 \$179 \$195 \$362 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1063 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1064 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1065 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1066 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1067 \$363 \$51 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1068 IBN5 \$51 \$363 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1069 \$364 \$51 IBN5 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1070 VDD \$51 \$364 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1071 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1072 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1073 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1074 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1075 \$365 \$196 \$933 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1076 VSS \$196 \$365 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1077 \$366 \$196 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1078 \$196 \$196 \$366 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1079 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1080 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1081 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1082 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1083 \$457 \$187 \$147 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1084 ITN1 \$187 \$457 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1085 \$458 IBN1 ITN1 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1086 \$47 IBN1 \$458 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1087 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1088 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1089 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1090 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1091 \$459 \$47 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1092 IBN1 \$47 \$459 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1093 \$460 \$47 IBN1 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1094 VDD \$47 \$460 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1095 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1096 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1097 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1098 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1099 \$461 \$188 \$188 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1100 VSS \$188 \$461 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1101 \$462 \$188 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1102 \$929 \$188 \$462 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1103 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1104 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1105 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1106 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1107 \$463 \$189 \$155 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1108 ITN2 \$189 \$463 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1109 \$464 IBN2 ITN2 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1110 \$48 IBN2 \$464 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1111 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1112 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1113 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1114 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1115 \$465 \$48 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1116 IBN2 \$48 \$465 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1117 \$466 \$48 IBN2 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1118 VDD \$48 \$466 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1119 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1120 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1121 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1122 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1123 \$467 \$190 \$190 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1124 VSS \$190 \$467 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1125 \$468 \$190 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1126 \$930 \$190 \$468 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1127 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1128 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1129 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1130 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1131 \$469 \$191 \$163 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1132 ITN3 \$191 \$469 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1133 \$470 IBN3 ITN3 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1134 \$49 IBN3 \$470 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1135 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1136 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1137 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1138 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1139 \$471 \$49 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1140 IBN3 \$49 \$471 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1141 \$472 \$49 IBN3 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1142 VDD \$49 \$472 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1143 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1144 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1145 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1146 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1147 \$473 \$192 \$192 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1148 VSS \$192 \$473 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1149 \$474 \$192 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1150 \$931 \$192 \$474 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1151 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1152 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1153 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1154 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1155 \$475 \$193 \$171 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1156 ITN4 \$193 \$475 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1157 \$476 IBN4 ITN4 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1158 \$50 IBN4 \$476 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1159 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1160 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1161 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1162 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1163 \$477 \$50 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1164 IBN4 \$50 \$477 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1165 \$478 \$50 IBN4 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1166 VDD \$50 \$478 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1167 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1168 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1169 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1170 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1171 \$479 \$194 \$194 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1172 VSS \$194 \$479 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1173 \$480 \$194 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1174 \$932 \$194 \$480 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1175 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1176 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1177 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1178 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1179 \$481 \$195 \$179 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1180 ITN5 \$195 \$481 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1181 \$482 IBN5 ITN5 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1182 \$51 IBN5 \$482 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1183 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1184 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1185 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1186 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1187 \$483 \$51 VDD VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1188 IBN5 \$51 \$483 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1189 \$484 \$51 IBN5 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1190 VDD \$51 \$484 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1191 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1192 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1193 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1194 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1195 \$485 \$196 \$196 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1196 VSS \$196 \$485 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1197 \$486 \$196 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1198 \$933 \$196 \$486 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1199 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1200 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1201 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1202 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1203 \$602 IBN1 \$47 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1204 ITN1 IBN1 \$602 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1205 \$603 \$187 ITN1 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1206 \$147 \$187 \$603 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1207 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1208 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1209 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1210 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1211 \$604 \$47 \$258 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1212 \$187 \$47 \$604 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1213 \$605 \$47 \$187 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1214 \$150 \$47 \$605 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1215 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1216 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1217 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1218 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1219 \$606 \$188 \$929 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1220 VSS \$188 \$606 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1221 \$607 \$188 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1222 \$188 \$188 \$607 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1223 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1224 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1225 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1226 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1227 \$608 IBN2 \$48 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1228 ITN2 IBN2 \$608 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1229 \$609 \$189 ITN2 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1230 \$155 \$189 \$609 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1231 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1232 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1233 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1234 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1235 \$610 \$48 \$260 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1236 \$189 \$48 \$610 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1237 \$611 \$48 \$189 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1238 \$158 \$48 \$611 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1239 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1240 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1241 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1242 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1243 \$612 \$190 \$930 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1244 VSS \$190 \$612 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1245 \$613 \$190 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1246 \$190 \$190 \$613 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1247 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1248 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1249 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1250 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1251 \$614 IBN3 \$49 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1252 ITN3 IBN3 \$614 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1253 \$615 \$191 ITN3 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1254 \$163 \$191 \$615 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1255 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1256 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1257 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1258 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1259 \$616 \$49 \$262 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1260 \$191 \$49 \$616 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1261 \$617 \$49 \$191 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1262 \$166 \$49 \$617 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1263 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1264 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1265 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1266 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1267 \$618 \$192 \$931 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1268 VSS \$192 \$618 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1269 \$619 \$192 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1270 \$192 \$192 \$619 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1271 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1272 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1273 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1274 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1275 \$620 IBN4 \$50 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1276 ITN4 IBN4 \$620 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1277 \$621 \$193 ITN4 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1278 \$171 \$193 \$621 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1279 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1280 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1281 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1282 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1283 \$622 \$50 \$264 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1284 \$193 \$50 \$622 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1285 \$623 \$50 \$193 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1286 \$174 \$50 \$623 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1287 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1288 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1289 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1290 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1291 \$624 \$194 \$932 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1292 VSS \$194 \$624 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1293 \$625 \$194 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1294 \$194 \$194 \$625 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1295 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1296 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1297 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1298 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1299 \$626 IBN5 \$51 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1300 ITN5 IBN5 \$626 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1301 \$627 \$195 ITN5 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1302 \$179 \$195 \$627 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1303 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1304 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1305 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1306 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1307 \$628 \$51 \$266 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1308 \$195 \$51 \$628 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1309 \$629 \$51 \$195 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1310 \$182 \$51 \$629 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1311 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1312 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1313 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1314 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1315 \$630 \$196 \$933 VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1316 VSS \$196 \$630 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1317 \$631 \$196 VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1318 \$196 \$196 \$631 VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1319 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1320 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1321 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1322 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1323 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1324 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1325 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1326 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1327 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1328 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1329 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1330 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1331 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1332 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1333 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1334 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1335 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1336 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1337 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1338 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1339 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1340 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1341 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1342 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1343 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1344 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1345 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1346 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1347 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1348 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1349 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1350 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1351 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1352 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1353 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1354 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1355 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1356 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1357 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1358 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1359 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1360 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1361 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1362 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1363 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1364 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1365 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1366 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1367 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1368 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1369 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1370 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1371 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1372 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1373 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1374 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1375 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1376 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1377 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1378 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1379 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1380 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1381 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1382 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1383 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1384 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1385 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1386 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1387 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1388 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1389 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1390 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1391 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1392 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1393 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1394 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1395 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1396 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1397 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1398 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1399 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1400 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1401 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1402 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1403 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1404 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1405 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1406 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1407 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1408 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1409 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1410 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1411 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1412 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1413 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1414 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1415 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1416 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1417 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1418 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1419 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1420 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1421 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1422 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1423 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1424 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1425 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1426 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1427 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1428 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1429 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1430 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1431 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1432 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1433 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1434 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1435 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1436 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1437 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1438 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1439 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1440 VSS VSS VSS VSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
.ENDS PRbiased_net_x5
