* NGSPICE file created from Filter_TOP.ext - technology: gf180mcuD

.subckt Filter_TOP VCM IN_POS IN_NEG VSS I1U VDD I1N IBNOUT OUT IBPOUT
X0 VSS.t3632 VSS.t3631 VSS.t3632 VSS.t1104 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1 a_52635_49681.t175 a_52635_34067.t65 VDD.t4975 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2 VDD.t4744 VDD.t4743 VDD.t4744 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3 VDD.t4742 VDD.t4741 VDD.t4742 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4 VDD.t4740 VDD.t4739 VDD.t4740 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5 VDD.t4738 VDD.t4737 VDD.t4738 VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6 a_100820_11614.t4 a_57977_n12421.t0 a_102796_6405# VSS.t171 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X7 a_31284_4481.t2 a_30324_4421.t0 a_30724_6405# VSS.t151 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X8 VDD.t4736 VDD.t4735 VDD.t4736 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X9 a_102756_12380# a_100820_10448.t11 VDD.t325 VDD.t298 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X10 a_36032_n36322.t0 a_53829_n36382.t8 a_55635_n36322# VDD.t297 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X11 a_33249_35053.t141 a_35502_25545.t28 VSS.t280 VSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X12 VSS.t3630 VSS.t3629 VSS.t3630 VSS.t571 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X13 VSS.t3628 VSS.t3627 VSS.t3628 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X14 a_101350_10448# a_100820_10448.t9 a_100820_10448.t10 VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X15 a_52635_49681.t174 a_52635_34067.t66 VDD.t4974 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X16 a_38619_n2651# a_31953_n19727.t74 a_38097_n2651# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X17 VDD.t4734 VDD.t4733 VDD.t4734 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X18 VSS.t3626 VSS.t3625 VSS.t3626 VSS.t905 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X19 VSS.t3624 VSS.t3623 VSS.t3624 VSS.t166 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X20 VDD.t45 a_31699_20742.t45 a_35502_24538.t23 VDD.t14 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X21 VSS.t3622 VSS.t3621 VSS.t3622 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X22 a_43817_6405# a_41891_4481.t11 VSS.t169 VSS.t158 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X23 VSS.t3620 VSS.t3619 VSS.t3620 VSS.t453 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X24 VSS.t3618 VSS.t3617 VSS.t3618 VSS.t979 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X25 VDD.t4732 VDD.t4731 VDD.t4732 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X26 a_105365_n7865# a_71281_n8397.t74 a_104527_n7865# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X27 VDD.t46 a_31699_20742.t46 a_35502_25545.t0 VDD.t38 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X28 a_52635_34067.t0 a_35922_19591.t6 a_52635_48695.t87 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X29 a_58851_n7138# a_50751_n19729.t74 a_58329_n8035# VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X30 a_53145_n19597# a_50751_n19729.t75 a_52585_n19597# VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X31 a_71864_n30339# a_65486_n36322.t8 a_71342_n30339.t2 VSS.t156 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X32 VDD.t4730 VDD.t4729 VDD.t4730 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X33 VSS.t3616 VSS.t3615 VSS.t3616 VSS.t558 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X34 a_106809_n17715.t1 a_71281_n8397.t75 a_106501_n21335# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X35 VSS.t3614 VSS.t3613 VSS.t3614 VSS.t98 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X36 VSS.t3612 VSS.t3611 VSS.t3612 VSS.t421 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X37 VDD.t4728 VDD.t4727 VDD.t4728 VDD.t18 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X38 VDD.t4726 VDD.t4725 VDD.t4726 VDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X39 a_105933_n2435# a_71281_n8397.t76 a_105365_n2435# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X40 VSS.t3610 VSS.t3609 VSS.t3610 VSS.t401 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X41 VDD.t4724 VDD.t4723 VDD.t4724 VDD.t3678 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X42 a_52635_34067.t1 a_35922_19591.t7 a_52635_48695.t86 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X43 VDD.t4722 VDD.t4721 VDD.t4722 VDD.t976 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X44 a_33249_48695.t334 a_31699_20742.t47 VDD.t48 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X45 VSS.t3608 VSS.t3607 VSS.t3608 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X46 a_52635_48695.t175 a_52635_34067.t67 VDD.t4973 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X47 VSS.t3606 VSS.t3605 VSS.t3606 VSS.t308 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X48 OUT.t107 a_35922_19591.t8 a_52635_49681.t0 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X49 VDD.t4720 VDD.t4719 VDD.t4720 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X50 VDD.t4718 VDD.t4717 VDD.t4718 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X51 VSS.t3604 VSS.t3603 VSS.t3604 VSS.t947 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X52 VSS.t3602 VSS.t3601 VSS.t3602 VSS.t908 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X53 VSS.t3600 VSS.t3599 VSS.t3600 VSS.t190 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X54 a_33249_48695.t333 a_31699_20742.t48 VDD.t50 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X55 VDD.t52 a_31699_20742.t49 a_33249_48695.t332 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X56 VDD.t4716 VDD.t4715 VDD.t4716 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X57 VSS.t3598 VSS.t3597 VSS.t3598 VSS.t1821 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X58 a_31284_n30339.t1 a_30324_n30399.t1 a_30724_n30339# VSS.t151 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X59 VSS.t3596 VSS.t3595 VSS.t3596 VSS.t339 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X60 VDD.t4714 VDD.t4713 VDD.t4714 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X61 OUT.t106 a_35922_19591.t9 a_52635_49681.t1 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X62 a_33249_35053.t88 a_35502_24538.t24 OUT.t19 VSS.t165 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X63 VDD.t4712 VDD.t4711 VDD.t4712 VDD.t944 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X64 a_38097_n5342.t1 a_100992_n29313.t0 a_101392_n29181# VSS.t332 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X65 VDD.t467 a_71281_n8397.t70 a_71281_n8397.t71 VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X66 a_101392_6405# a_100992_4421.t0 a_100820_10448.t0 VSS.t163 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X67 VDD.t4710 VDD.t4709 VDD.t4710 VDD.t875 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X68 a_52635_48695.t85 a_35922_19591.t10 a_52635_34067.t2 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X69 VDD.t54 a_31699_20742.t50 a_33249_48695.t331 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X70 VSS.t3594 VSS.t3593 VSS.t3594 VSS.t638 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X71 VDD.t4708 VDD.t4707 VDD.t4708 VDD.t2464 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X72 a_100235_n15000# a_71281_n8397.t77 a_99667_n15000# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X73 VDD.t4706 VDD.t4705 VDD.t4706 VDD.t1419 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X74 VSS.t3592 VSS.t3591 VSS.t3592 VSS.t896 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X75 a_73302_13546# a_71496_10388.t8 a_71342_4481.t2 VDD.t363 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X76 a_30724_6405# a_30324_4421.t0 a_30152_10448.t3 VSS.t150 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X77 VDD.t4704 VDD.t4703 VDD.t4704 VDD.t976 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X78 VSS.t3590 VSS.t3589 VSS.t3590 VSS.t195 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X79 VDD.t4702 VDD.t4701 VDD.t4702 VDD.t1747 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X80 VDD.t4700 VDD.t4699 VDD.t4700 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X81 VSS.t3588 VSS.t3587 VSS.t3588 VSS.t650 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X82 a_31831_n5342.t1 a_32913_n8930.t1 a_83725_n28415# VSS.t288 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X83 a_45445_n18698# a_31953_n19727.t75 a_44885_n17801# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X84 VSS.t3586 VSS.t3585 VSS.t3586 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X85 VDD.t56 a_31699_20742.t51 a_33249_48695.t330 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X86 OUT.t105 a_35922_19591.t11 a_52635_49681.t2 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X87 VDD.t4698 VDD.t4697 VDD.t4698 VDD.t944 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X88 VSS.t3584 VSS.t3583 VSS.t3584 VSS.t522 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X89 VDD.t4696 VDD.t4695 VDD.t4696 VDD.t309 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X90 VDD.t4694 VDD.t4693 VDD.t4694 VDD.t2447 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X91 VSS.t3582 VSS.t3581 VSS.t3582 VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X92 a_51711_n5344.t1 a_50751_n19729.t76 a_51151_n5344# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X93 a_66551_n17803# a_50751_n19729.t77 a_66029_n18700# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X94 a_33249_35053.t0 a_33379_34917.t3 a_33249_48695.t14 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X95 VSS.t3580 VSS.t3579 VSS.t3580 VSS.t687 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X96 a_33249_35053.t1 a_33379_34917.t4 a_33249_48695.t15 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X97 a_98829_n17715# a_71281_n8397.t78 a_98299_n16810# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X98 OUT.t104 a_35922_19591.t12 a_52635_49681.t3 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X99 VSS.t3578 VSS.t3577 VSS.t3578 VSS.t1537 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X100 a_73302_11614# a_71496_10388.t9 VSS.t3649 VDD.t363 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X101 a_73268_n29181# a_65486_n36322.t9 a_45445_n19595.t1 VSS.t154 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X102 a_90245_n6055# a_71281_n10073.t74 a_60677_10448.t0 VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X103 VDD.t4692 VDD.t4691 VDD.t4692 VDD.t544 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X104 VSS.t3576 VSS.t3575 VSS.t3576 VSS.t884 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X105 a_98829_n15000# a_71281_n8397.t79 a_98299_n15905# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X106 a_51711_n14215# a_50751_n19729.t78 a_51151_n14215# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X107 VDD.t4690 VDD.t4689 VDD.t4690 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X108 VDD.t4688 VDD.t4687 VDD.t4688 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X109 VSS.t3574 VSS.t3573 VSS.t3574 VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X110 VSS.t3572 VSS.t3571 VSS.t3572 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X111 a_33249_48695.t350 a_33379_34007.t4 a_33249_34067.t105 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X112 VDD.t4686 VDD.t4685 VDD.t4686 VDD.t568 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X113 VDD.t4684 VDD.t4683 VDD.t4684 VDD.t930 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X114 a_65486_n35156.t5 a_65486_n35156.t4 a_67422_n36322# VDD.t1 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X115 a_60285_n2653# a_50751_n19729.t79 a_59763_n3550# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X116 a_71281_n8397.t69 a_71281_n8397.t68 VDD.t466 VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X117 VDD.t4682 VDD.t4681 VDD.t4682 VDD.t1494 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X118 a_105365_n15000# a_71281_n8397.t80 a_104527_n15000# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X119 VDD.t4680 VDD.t4679 VDD.t4680 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X120 a_106676_n30339.t0 a_100820_n36322.t8 a_108602_n27257# VSS.t333 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X121 VDD.t4678 VDD.t4677 VDD.t4678 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X122 VSS.t3570 VSS.t3569 VSS.t3570 VSS.t681 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X123 a_40613_n8930# a_31953_n19727.t76 a_40053_n8930# VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X124 a_33249_48695.t351 a_33379_34007.t5 a_33249_34067.t104 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X125 VDD.t4676 VDD.t4675 VDD.t4676 VDD.t351 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X126 VDD.t4674 VDD.t4673 VDD.t4674 VDD.t341 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X127 OUT.t103 a_35922_19591.t13 a_52635_49681.t4 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X128 VSS.t3568 VSS.t3567 VSS.t3568 VSS.t834 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X129 VSS.t3566 VSS.t3565 VSS.t3566 VSS.t817 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X130 a_110225_n1530# a_71281_n8397.t81 a_109695_n5150# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X131 a_52635_48695.t84 a_35922_19591.t14 a_52635_34067.t3 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X132 a_88271_n3340# a_71281_n10073.t75 a_87433_n3340# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X133 VDD.t4762 a_83153_11614.t8 a_90935_5639# VSS.t392 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X134 VDD.t4672 VDD.t4671 VDD.t4672 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X135 VDD.t4670 VDD.t4669 VDD.t4670 VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X136 VSS.t3564 VSS.t3563 VSS.t3564 VSS.t220 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X137 a_114516_10448# a_86903_n14095.t3 a_89715_n17715.t2 VDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X138 VDD.t4668 VDD.t4667 VDD.t4668 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X139 a_39179_n8033# a_31953_n19727.t77 a_38619_n8033# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X140 VDD.t57 a_31699_20742.t52 a_35502_25545.t1 VDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X141 VSS.t3562 VSS.t3561 VSS.t3562 VSS.t653 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X142 VDD.t4666 VDD.t4665 VDD.t4666 VDD.t1714 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X143 VSS.t254 a_50751_n19729.t70 a_50751_n19729.t71 VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X144 VDD.t4664 VDD.t4663 VDD.t4664 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X145 a_84547_n15000# a_71281_n10073.t76 a_83709_n14095# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X146 VDD.t4662 VDD.t4661 VDD.t4662 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X147 a_100235_n20430# a_71281_n8397.t82 a_99667_n20430# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X148 VDD.t4660 VDD.t4659 VDD.t4660 VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X149 a_52635_49681.t5 a_35922_19591.t15 OUT.t102 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X150 VDD.t3 a_65486_n35156.t12 a_66016_n36322# VDD.t2 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X151 a_67111_n2653# a_50751_n19729.t80 a_66551_n1756# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X152 VDD.t4658 VDD.t4657 VDD.t4658 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X153 VDD.t4656 VDD.t4655 VDD.t4656 VDD.t1867 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X154 VDD.t4654 VDD.t4653 VDD.t4654 VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X155 VDD.t4652 VDD.t4651 VDD.t4652 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X156 a_54579_n4447# a_50751_n19729.t81 a_54019_n4447# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X157 a_32353_n7136# a_31953_n19727.t78 a_31831_n7136# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X158 VSS.t3560 VSS.t3559 VSS.t3560 VSS.t107 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X159 VSS.t295 a_112559_4481.t11 a_113081_5639# VSS.t294 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X160 a_30324_n30399.t1 a_30152_n36322.t8 a_36530_n29181# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X161 VDD.t4650 VDD.t4649 VDD.t4650 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X162 VDD.t4648 VDD.t4647 VDD.t4648 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X163 VSS.t3558 VSS.t3557 VSS.t3558 VSS.t868 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X164 a_34347_n7136# a_31953_n19727.t79 a_33787_n7136# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X165 VDD.t4646 VDD.t4645 VDD.t4646 VDD.t2399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X166 a_48349_n35156# a_47819_n35156.t7 a_47819_n35156.t8 VDD.t2559 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X167 VSS.t3556 VSS.t3555 VSS.t3556 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X168 a_51711_n12421.t0 a_83153_11614.t9 a_89531_6405# VSS.t393 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X169 a_101350_n34390# a_100820_n35156.t12 a_100820_n36322.t0 VDD.t523 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X170 VSS.t3554 VSS.t3553 VSS.t3554 VSS.t25 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X171 VSS.t3552 VSS.t3551 VSS.t3552 VSS.t1360 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X172 a_77225_4481.t7 a_77225_4481.t6 a_79151_5639# VSS.t318 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X173 a_106676_4481.t0 a_106830_10388.t8 a_107230_10448# VDD.t519 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X174 VDD.t4644 VDD.t4643 VDD.t4644 VDD.t898 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X175 VSS.t3550 VSS.t3549 VSS.t3550 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X176 a_33249_48695.t346 a_33379_34007.t6 a_33249_34067.t103 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X177 VSS.t3548 VSS.t3547 VSS.t3548 VSS.t65 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X178 VSS.t3546 VSS.t3545 VSS.t3546 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X179 a_57417_n8932# a_50751_n19729.t82 a_56895_n8932# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X180 VDD.t4642 VDD.t4641 VDD.t4642 VDD.t2777 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X181 a_98829_n20430# a_71281_n8397.t83 a_36032_n35156.t0 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X182 VDD.t4640 VDD.t4639 VDD.t4640 VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X183 VDD.t4638 VDD.t4637 VDD.t4638 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X184 VSS.t3544 VSS.t3543 VSS.t3544 VSS.t129 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X185 VDD.t4636 VDD.t4635 VDD.t4636 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X186 VDD.t4634 VDD.t4633 VDD.t4634 VDD.t496 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X187 a_30152_n35156.t5 a_30152_n35156.t4 a_32088_n34390# VDD.t551 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X188 VSS.t3542 VSS.t3541 VSS.t3542 VSS.t537 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X189 VDD.t4632 VDD.t4631 VDD.t4632 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X190 a_89563_13546# a_89163_10388.t8 a_89033_13546.t3 VDD.t552 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X191 a_67422_13546# a_65486_10448.t11 VDD.t4745 VDD.t866 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X192 VDD.t4630 VDD.t4629 VDD.t4630 VDD.t2382 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X193 a_51151_n17803# a_50751_n19729.t83 a_50629_n17803# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X194 VSS.t3540 VSS.t3539 VSS.t3540 VSS.t853 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X195 VDD.t4628 VDD.t4627 VDD.t4628 VDD.t1658 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X196 a_43010_10448.t4 a_36032_11614.t3 a_42442_13546# VDD.t289 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X197 VSS.t3538 VSS.t3537 VSS.t3538 VSS.t842 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X198 a_52635_34067.t4 a_35922_19591.t16 a_52635_48695.t83 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X199 a_48349_n33224# a_47819_n35156.t3 a_47819_n35156.t4 VDD.t2559 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X200 a_42047_n19595# a_31953_n19727.t80 a_41487_n19595# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X201 a_30682_10448# a_30152_10448.t4 a_30152_10448.t5 VDD.t302 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X202 VDD.t4626 VDD.t4625 VDD.t4626 VDD.t571 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X203 VDD.t4624 VDD.t4623 VDD.t4624 VDD.t955 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X204 a_32088_n36322# a_30152_n35156.t12 VDD.t4977 VDD.t2088 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X205 VDD.t4622 VDD.t4621 VDD.t4622 VDD.t855 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X206 a_105365_n20430# a_71281_n8397.t84 a_104527_n20430# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X207 VDD.t4620 VDD.t4619 VDD.t4620 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X208 VSS.t3536 VSS.t3535 VSS.t3536 VSS.t18 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X209 VDD.t4972 a_52635_34067.t68 a_52635_48695.t174 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X210 OUT.t101 a_35922_19591.t17 a_52635_49681.t6 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X211 VDD.t4618 VDD.t4617 VDD.t4618 VDD.t898 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X212 VDD.t4616 VDD.t4615 VDD.t4616 VDD.t302 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X213 a_52635_34067.t5 a_35922_19591.t18 a_52635_48695.t82 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X214 VDD.t4614 VDD.t4613 VDD.t4614 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X215 VDD.t44 a_31699_20742.t43 a_31699_20742.t44 VDD.t38 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X216 a_33249_48695.t329 a_31699_20742.t53 VDD.t59 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X217 VSS.t3534 VSS.t3533 VSS.t3534 VSS.t379 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X218 VSS.t3532 VSS.t3531 VSS.t3532 VSS.t837 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X219 OUT.t100 a_35922_19591.t19 a_52635_49681.t7 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X220 a_52635_34067.t6 a_35922_19591.t20 a_52635_48695.t81 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X221 VDD.t4612 VDD.t4611 VDD.t4612 VDD.t1818 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X222 a_89563_11614# a_89163_10388.t9 a_81205_n14095.t2 VDD.t552 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X223 a_67422_11614# a_65486_10448.t12 VDD.t4746 VDD.t866 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X224 VDD.t4610 VDD.t4609 VDD.t4610 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X225 a_44885_n6239# a_31953_n19727.t81 a_44363_n7136# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X226 a_52635_49681.t8 a_35922_19591.t21 OUT.t99 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X227 VDD.t4608 VDD.t4607 VDD.t4608 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X228 a_31953_n19727.t71 a_31953_n19727.t70 VSS.t95 VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X229 a_43010_10448.t0 a_36032_11614.t4 a_42442_11614# VDD.t289 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X230 VSS.t3530 VSS.t3529 VSS.t3530 VSS.t558 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X231 VDD.t4606 VDD.t4605 VDD.t4606 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X232 VSS.t341 a_89163_n36382.t8 a_89563_n35156# VDD.t547 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X233 VSS.t3528 VSS.t3527 VSS.t3528 VSS.t1426 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X234 VDD.t4604 VDD.t4603 VDD.t4604 VDD.t2344 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X235 VDD.t4602 VDD.t4601 VDD.t4602 VDD.t855 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X236 a_31953_n19727.t69 a_31953_n19727.t68 VSS.t94 VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X237 a_47753_n15110# a_31953_n19727.t82 a_47231_n16904# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X238 VDD.t4600 VDD.t4599 VDD.t4600 VDD.t813 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X239 VDD.t4598 VDD.t4597 VDD.t4598 VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X240 VDD.t4596 VDD.t4595 VDD.t4596 VDD.t401 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X241 VSS.t3526 VSS.t3525 VSS.t3526 VSS.t337 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X242 a_89531_6405# a_83153_11614.t10 VDD.t4763 VSS.t394 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X243 a_107339_n6055# a_71281_n8397.t85 a_106809_n5150.t2 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X244 VSS.t3524 VSS.t3523 VSS.t3524 VSS.t763 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X245 VDD.t4594 VDD.t4593 VDD.t4594 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X246 VDD.t4592 VDD.t4591 VDD.t4592 VDD.t434 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X247 a_52635_34067.t61 a_35502_24538.t25 a_33249_34067.t17 VSS.t165 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X248 VSS.t368 a_41891_n29181.t11 a_42413_n27257# VSS.t166 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X249 VDD.t4590 VDD.t4589 VDD.t4590 VDD.t667 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X250 VDD.t4588 VDD.t4587 VDD.t4588 VDD.t920 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X251 VDD.t4586 VDD.t4585 VDD.t4586 VDD.t1787 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X252 VDD.t4584 VDD.t4583 VDD.t4584 VDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X253 VDD.t4582 VDD.t4581 VDD.t4582 VDD.t423 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X254 VSS.t3522 VSS.t3521 VSS.t3522 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X255 a_33249_48695.t347 a_33379_34007.t7 a_33249_34067.t102 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X256 a_89407_n6960# a_71281_n10073.t77 a_88839_n6960# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X257 VSS.t3520 VSS.t3519 VSS.t3520 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X258 VSS.t3518 VSS.t3517 VSS.t3518 VSS.t531 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X259 VDD.t4580 VDD.t4579 VDD.t4580 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X260 a_89009_n27257.t2 a_89163_n36382.t9 a_89563_n33224# VDD.t547 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X261 a_89033_13546.t2 a_89163_10388.t10 a_90969_10448# VDD.t553 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X262 a_31699_20742.t42 a_31699_20742.t41 VDD.t43 VDD.t20 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X263 VDD.t4578 VDD.t4577 VDD.t4578 VDD.t47 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X264 a_53699_n36322.t3 a_71496_n36382.t8 a_73302_n36322# VDD.t2058 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X265 VDD.t4576 VDD.t4575 VDD.t4576 VDD.t813 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X266 VSS.t3516 VSS.t3515 VSS.t3516 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X267 VDD.t4574 VDD.t4573 VDD.t4574 VDD.t828 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X268 a_100235_n15905# a_71281_n8397.t86 a_99667_n15905# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X269 VSS.t3514 VSS.t3513 VSS.t3514 VSS.t1794 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X270 VDD.t4572 VDD.t4571 VDD.t4572 VDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X271 VDD.t4570 VDD.t4569 VDD.t4570 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X272 a_33249_48695.t16 a_33379_34917.t5 a_33249_35053.t2 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X273 VDD.t61 a_31699_20742.t54 a_33249_48695.t328 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X274 a_40613_n14213# a_31953_n19727.t83 a_40053_n14213# VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X275 VSS.t3512 VSS.t3511 VSS.t3512 VSS.t340 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X276 a_67462_n29181# a_45445_n19595.t2 a_44363_n16007.t1 VSS.t289 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X277 a_31699_20742.t40 a_31699_20742.t39 VDD.t42 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X278 VDD.t4568 VDD.t4567 VDD.t4568 VDD.t2302 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X279 VDD.t4566 VDD.t4565 VDD.t4566 VDD.t439 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X280 a_94537_n9675# a_71281_n10073.t78 a_93969_n9675# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X281 VDD.t4564 VDD.t4563 VDD.t4564 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X282 a_78344_n36322.t3 a_71366_n35156.t5 a_77776_n36322# VDD.t502 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X283 a_33249_34067.t101 a_33379_34007.t8 a_33249_48695.t348 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X284 a_52635_34067.t7 a_35922_19591.t22 a_52635_48695.t80 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X285 VDD.t4562 VDD.t4561 VDD.t4562 VDD.t351 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X286 VSS.t3510 VSS.t3509 VSS.t3510 VSS.t331 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X287 VDD.t4560 VDD.t4559 VDD.t4560 VDD.t1642 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X288 VSS.t3508 VSS.t3507 VSS.t3508 VSS.t1466 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X289 VSS.t3506 VSS.t3505 VSS.t3506 VSS.t811 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X290 VDD.t4558 VDD.t4557 VDD.t4558 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X291 VDD.t4556 VDD.t4555 VDD.t4556 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X292 a_39179_n19595.t1 a_31953_n19727.t84 a_38619_n19595# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X293 VSS.t3504 VSS.t3503 VSS.t3504 VSS.t397 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X294 VDD.t4554 VDD.t4553 VDD.t4554 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X295 VSS.t3502 VSS.t3501 VSS.t3502 VSS.t638 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X296 VSS.t3500 VSS.t3499 VSS.t3500 VSS.t808 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X297 a_60845_n19597# a_50751_n19729.t84 a_60285_n18700# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X298 VDD.t4552 VDD.t4551 VDD.t4552 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X299 VDD.t4550 VDD.t4549 VDD.t4550 VDD.t635 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X300 VDD.t4548 VDD.t4547 VDD.t4548 VDD.t828 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X301 VDD.t4546 VDD.t4545 VDD.t4546 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X302 VSS.t3498 VSS.t3497 VSS.t3498 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X303 a_71342_n30339.t0 a_71496_n36382.t9 a_71896_n36322# VDD.t2021 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X304 VDD.t4544 VDD.t4543 VDD.t4544 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X305 VSS.t3496 VSS.t3495 VSS.t3496 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X306 VDD.t4542 VDD.t4541 VDD.t4542 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X307 VSS.t3494 VSS.t3493 VSS.t3494 VSS.t1385 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X308 VSS.t3492 VSS.t3491 VSS.t3492 VSS.t297 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X309 a_60285_n19597# a_50751_n19729.t85 a_57977_n19597# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X310 a_98829_n15905# a_71281_n8397.t87 a_98299_n15905# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X311 VSS.t3490 VSS.t3489 VSS.t3490 VSS.t266 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X312 VSS.t3488 VSS.t3487 VSS.t3488 VSS.t859 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X313 VSS.t3486 VSS.t3485 VSS.t3486 VSS.t1104 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X314 a_61484_4481# a_59558_4481.t11 VSS.t400 VSS.t399 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X315 VDD.t4540 VDD.t4539 VDD.t4540 VDD.t2254 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X316 a_54229_n35156# a_53829_n36382.t9 a_53699_n35156.t1 VDD.t417 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X317 a_82573_n13190# a_71281_n10073.t79 a_81735_n13190# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X318 VDD.t4538 VDD.t4537 VDD.t4538 VDD.t2680 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X319 VDD.t4536 VDD.t4535 VDD.t4536 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X320 VDD.t4534 VDD.t4533 VDD.t4534 VDD.t610 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X321 VSS.t3484 VSS.t3483 VSS.t3484 VSS.t687 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X322 VSS.t3482 VSS.t3481 VSS.t3482 VSS.t792 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X323 a_105365_n15905# a_71281_n8397.t88 a_104527_n15905# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X324 VSS.t3480 VSS.t3479 VSS.t3480 VSS.t817 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X325 VSS.t3478 VSS.t3477 VSS.t3478 VSS.t261 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X326 VSS.t152 a_35502_25545.t29 a_33249_35053.t140 VSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X327 VDD.t4532 VDD.t4531 VDD.t4532 VDD.t792 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X328 VSS.t3476 VSS.t3475 VSS.t3476 VSS.t553 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X329 a_39179_n3548# a_31953_n19727.t85 a_38619_n3548# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X330 a_94892_n29181.t2 a_83325_n29313.t1 a_96849_n36322# VDD.t1996 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X331 VDD.t4530 VDD.t4529 VDD.t4530 VDD.t789 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X332 VDD.t4528 VDD.t4527 VDD.t4528 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X333 a_54579_n19597# a_50751_n19729.t86 a_54019_n18700# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X334 a_32353_n15110# a_31953_n19727.t86 a_31831_n15110# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X335 VSS.t3474 VSS.t3473 VSS.t3474 VSS.t220 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X336 VDD.t4526 VDD.t4525 VDD.t4526 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X337 a_64243_n18700# a_50751_n19729.t87 a_63683_n18700# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X338 a_54019_n4447# a_50751_n19729.t88 a_53497_n6241# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X339 VSS.t253 a_50751_n19729.t68 a_50751_n19729.t69 VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X340 VSS.t3472 VSS.t3471 VSS.t3472 VSS.t413 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X341 a_54229_n33224# a_53829_n36382.t10 a_36032_n36322.t1 VDD.t417 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X342 VSS.t3470 VSS.t3469 VSS.t3470 VSS.t265 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X343 a_88271_n2435# a_71281_n10073.t80 a_87433_n2435# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X344 a_31699_19142# I1U.t2 a_30377_18342# VSS.t349 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X345 VSS.t3468 VSS.t3467 VSS.t3468 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X346 a_79151_n29181# a_77225_n29181.t11 VSS.t382 VSS.t381 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X347 a_52635_34067.t8 a_35922_19591.t23 a_52635_48695.t79 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X348 VDD.t4524 VDD.t4523 VDD.t4524 VDD.t792 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X349 VSS.t3466 VSS.t3465 VSS.t3466 VSS.t775 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X350 a_52635_34067.t9 a_35922_19591.t24 a_52635_48695.t78 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X351 VSS.t3464 VSS.t3463 VSS.t3464 VSS.t409 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X352 VDD.t4522 VDD.t4521 VDD.t4522 VDD.t920 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X353 VDD.t4520 VDD.t4519 VDD.t4520 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X354 VDD.t4518 VDD.t4517 VDD.t4518 VDD.t755 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X355 a_81735_n8770# a_71281_n10073.t81 VDD.t370 VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X356 VSS.t3462 VSS.t3461 VSS.t3462 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X357 VSS.t3460 VSS.t3459 VSS.t3460 VSS.t323 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X358 a_48313_n13316# a_31953_n19727.t87 a_47753_n13316# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X359 OUT.t98 a_35922_19591.t25 a_52635_49681.t9 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X360 VDD.t4516 VDD.t4515 VDD.t4516 VDD.t2812 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X361 a_63161_n5344.t1 a_64243_n1756.t1 a_66058_7563# VSS.t377 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X362 VSS.t3458 VSS.t3457 VSS.t3458 VSS.t653 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X363 VDD.t4514 VDD.t4513 VDD.t4514 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X364 VSS.t3456 VSS.t3455 VSS.t3456 VSS.t289 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X365 VDD.t4512 VDD.t4511 VDD.t4512 VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X366 OUT.t97 a_35922_19591.t26 a_52635_49681.t10 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X367 a_33249_35053.t3 a_33379_34917.t6 a_33249_48695.t17 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X368 VSS.t3454 VSS.t3453 VSS.t3454 VSS.t1431 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X369 VDD.t4510 VDD.t4509 VDD.t4510 VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X370 VSS.t3452 VSS.t3451 VSS.t3452 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X371 VSS.t3450 VSS.t3449 VSS.t3450 VSS.t795 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X372 VDD.t63 a_31699_20742.t55 a_33249_48695.t327 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X373 a_36008_4481.t0 a_30152_11614.t8 a_37934_7563# VSS.t281 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X374 a_33249_48695.t349 a_33379_34007.t9 a_33249_34067.t100 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X375 a_58851_n14215# a_50751_n19729.t89 a_58329_n14215# VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X376 a_102796_n30339# a_100992_n29313.t0 a_38097_n5342.t2 VSS.t330 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X377 a_96011_n36322.t0 a_83325_n29313.t1 a_95443_n35156# VDD.t2422 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X378 a_98829_n8770# a_71281_n8397.t89 a_89033_n35156.t0 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X379 a_83725_n29181# a_83325_n29313.t0 a_83153_n35156.t8 VSS.t287 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X380 VSS.t3448 VSS.t3447 VSS.t3448 VSS.t281 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X381 VDD.t4508 VDD.t4507 VDD.t4508 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X382 a_52635_34067.t10 a_35922_19591.t27 a_52635_48695.t77 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X383 a_77747_7563# a_77225_4481.t11 a_71496_10388.t0 VSS.t317 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X384 a_57977_n18700# a_50751_n19729.t90 a_57417_n18700# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X385 VSS.t3446 VSS.t3445 VSS.t3446 VSS.t29 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X386 VSS.t3444 VSS.t3443 VSS.t3444 VSS.t396 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X387 VDD.t65 a_31699_20742.t56 a_33249_48695.t326 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X388 VSS.t3442 VSS.t3441 VSS.t3442 VSS.t1253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X389 VDD.t4506 VDD.t4505 VDD.t4506 VDD.t78 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X390 VDD.t4971 a_52635_34067.t69 a_52635_48695.t173 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X391 VSS.t3440 VSS.t3439 VSS.t3440 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X392 VDD.t4504 VDD.t4503 VDD.t4504 VDD.t755 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X393 VSS.t3438 VSS.t3437 VSS.t3438 VSS.t733 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X394 a_108636_13546# a_106830_10388.t9 a_106676_4481.t1 VDD.t520 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X395 VSS.t3436 VSS.t3435 VSS.t3436 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X396 VDD.t4502 VDD.t4501 VDD.t4502 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X397 VSS.t3434 VSS.t3433 VSS.t3434 VSS.t591 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X398 a_57417_n16009# a_50751_n19729.t91 a_56895_n16009.t0 VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X399 VDD.t4500 VDD.t4499 VDD.t4500 VDD.t404 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X400 a_87433_n9675# a_71281_n10073.t82 a_86903_n9675# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X401 a_33787_n17801# a_31953_n19727.t88 a_33265_n18698# VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X402 a_96011_n36322.t1 a_83325_n29313.t1 a_95443_n33224# VDD.t2422 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X403 VDD.t4498 VDD.t4497 VDD.t4498 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X404 VDD.t4496 VDD.t4495 VDD.t4496 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X405 VSS.t3432 VSS.t3431 VSS.t3432 VSS.t498 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X406 VSS.t3430 VSS.t3429 VSS.t3430 VSS.t1064 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X407 VSS.t3428 VSS.t3427 VSS.t3428 VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X408 VDD.t4494 VDD.t4493 VDD.t4494 VDD.t1370 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X409 VDD.t4492 VDD.t4491 VDD.t4492 VDD.t78 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X410 VDD.t4490 VDD.t4489 VDD.t4490 VDD.t748 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X411 VSS.t93 a_31953_n19727.t66 a_31953_n19727.t67 VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X412 VSS.t3426 VSS.t3425 VSS.t3426 VSS.t260 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X413 VSS.t3424 VSS.t3423 VSS.t3424 VSS.t748 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X414 a_33249_34067.t99 a_33379_34007.t10 a_33249_48695.t8 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X415 VSS.t3422 VSS.t3421 VSS.t3422 VSS.t0 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X416 VSS.t3420 VSS.t3419 VSS.t3420 VSS.t283 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X417 VDD.t4488 VDD.t4487 VDD.t4488 VDD.t1549 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X418 a_108636_11614# a_106830_10388.t10 VSS.t313 VDD.t520 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X419 a_64243_n8932# a_50751_n19729.t92 a_63683_n8932# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X420 a_32128_7563# a_30324_4421.t0 a_31284_4481.t2 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X421 VDD.t4486 VDD.t4485 VDD.t4486 VDD.t2189 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X422 a_66551_n4447# a_50751_n19729.t93 a_66029_n6241# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X423 a_52635_48695.t172 a_52635_34067.t70 VDD.t4970 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X424 VSS.t3418 VSS.t3417 VSS.t3418 VSS.t763 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X425 VDD.t67 a_31699_20742.t57 a_33249_48695.t325 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X426 VSS.t3416 VSS.t3415 VSS.t3416 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X427 VSS.t3414 VSS.t3413 VSS.t3414 VSS.t311 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X428 a_30152_n35156.t1 a_30324_n29313.t0 a_32128_n28415# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X429 VDD.t4484 VDD.t4483 VDD.t4484 VDD.t725 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X430 a_33249_48695.t324 a_31699_20742.t58 VDD.t69 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X431 VSS.t3412 VSS.t3411 VSS.t3412 VSS.t740 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X432 a_52635_48695.t171 a_52635_34067.t71 VDD.t4969 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X433 VDD.t71 a_31699_20742.t59 a_33249_48695.t323 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X434 VDD.t4968 a_52635_34067.t72 a_52635_49681.t173 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X435 VDD.t4482 VDD.t4481 VDD.t4482 VDD.t748 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X436 VSS.t3410 VSS.t3409 VSS.t3410 VSS.t760 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X437 VDD.t4480 VDD.t4479 VDD.t4480 VDD.t34 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X438 VSS.t3408 VSS.t3407 VSS.t3408 VSS.t1222 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X439 VSS.t3406 VSS.t3405 VSS.t3406 VSS.t1253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X440 a_33249_35053.t4 a_33379_34917.t7 a_33249_48695.t18 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X441 OUT.t96 a_35922_19591.t28 a_52635_49681.t11 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X442 a_48313_n7136# a_31953_n19727.t89 a_47753_n7136# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X443 a_45706_22884# a_35922_19591.t29 a_45138_22884# VDD.t402 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X444 VSS.t412 a_112559_n29181.t11 a_113081_n28415# VSS.t411 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X445 a_107339_n6960# a_71281_n8397.t90 a_106501_n4245# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X446 VSS.t3404 VSS.t3403 VSS.t3404 VSS.t684 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X447 VDD.t4478 VDD.t4477 VDD.t4478 VDD.t120 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X448 VDD.t4476 VDD.t4475 VDD.t4476 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X449 a_49755_12380# a_47819_10448.t11 VDD.t509 VDD.t508 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X450 VDD.t4967 a_52635_34067.t73 a_52635_48695.t170 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X451 VSS.t3402 VSS.t3401 VSS.t3402 VSS.t1306 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X452 VSS.t3400 VSS.t3399 VSS.t3400 VSS.t1303 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X453 VSS.t3398 VSS.t3397 VSS.t3398 VSS.t576 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X454 a_43848_13546# a_30324_4421.t1 a_43010_10448.t0 VDD.t290 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X455 VDD.t4474 VDD.t4473 VDD.t4474 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X456 VDD.t4472 VDD.t4471 VDD.t4472 VDD.t2160 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X457 VDD.t4470 VDD.t4469 VDD.t4470 VDD.t725 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X458 a_47819_n36322.t7 a_39179_n19595.t0 a_49795_n27257# VSS.t337 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X459 VSS.t3396 VSS.t3395 VSS.t3396 VSS.t615 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X460 a_93131_n8770# a_71281_n10073.t83 VDD.t308 VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X461 VDD.t4468 VDD.t4467 VDD.t4468 VDD.t2155 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X462 VSS.t194 a_53829_n36382.t11 a_54229_n34390# VDD.t301 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X463 a_35502_25545.t2 a_31699_20742.t60 VDD.t72 VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X464 VSS.t3394 VSS.t3393 VSS.t3394 VSS.t671 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X465 VSS.t3392 VSS.t3391 VSS.t3392 VSS.t1294 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X466 a_33249_35053.t139 a_35502_25545.t30 VSS.t176 VSS.t145 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X467 a_84017_n17715.t2 a_83325_4421.t1 a_95443_12380# VDD.t498 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X468 VDD.t4466 VDD.t4465 VDD.t4466 VDD.t55 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X469 OUT.t95 a_35922_19591.t30 a_52635_49681.t12 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X470 VSS.t3390 VSS.t3389 VSS.t3390 VSS.t107 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X471 VSS.t3388 VSS.t3387 VSS.t3388 VSS.t1287 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X472 VSS.t3386 VSS.t3385 VSS.t3386 VSS.t398 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X473 VDD.t4464 VDD.t4463 VDD.t4464 VDD.t2142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X474 VSS.t3384 VSS.t3383 VSS.t3384 VSS.t609 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X475 VSS.t3382 VSS.t3381 VSS.t3382 VSS.t304 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X476 VDD.t465 a_71281_n8397.t66 a_71281_n8397.t67 VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X477 a_105365_n1530# a_71281_n8397.t91 a_104527_n1530# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X478 OUT.t94 a_35922_19591.t31 a_52635_49681.t13 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X479 VDD.t74 a_31699_20742.t61 a_33249_48695.t322 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X480 a_43848_11614# a_30324_4421.t1 a_43010_10448.t2 VDD.t290 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X481 a_35502_25545.t3 a_31699_20742.t62 VDD.t75 VDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X482 a_38619_n12419# a_31953_n19727.t90 a_38097_n13316# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X483 VDD.t4966 a_52635_34067.t74 a_52635_48695.t169 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X484 VSS.t3380 VSS.t3379 VSS.t3380 VSS.t147 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X485 a_105933_n15000# a_71281_n8397.t92 a_105365_n15000# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X486 VSS.t3378 VSS.t3377 VSS.t3378 VSS.t284 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X487 VSS.t3376 VSS.t3375 VSS.t3376 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X488 a_90935_n30339# a_83153_n36322.t8 a_83325_n29313.t0 VSS.t452 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X489 VDD.t4965 a_52635_34067.t75 a_52635_48695.t168 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X490 VSS.t252 a_50751_n19729.t66 a_50751_n19729.t67 VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X491 VDD.t4462 VDD.t4461 VDD.t4462 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X492 a_47819_n36322.t0 a_47819_n35156.t12 a_49755_n35156# VDD.t2325 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X493 VDD.t4460 VDD.t4459 VDD.t4460 VDD.t2127 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X494 a_52635_49681.t172 a_52635_34067.t76 VDD.t4964 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X495 VDD.t4458 VDD.t4457 VDD.t4458 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X496 VSS.t3374 VSS.t3373 VSS.t3374 VSS.t310 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X497 VDD.t4456 VDD.t4455 VDD.t4456 VDD.t648 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X498 VDD.t4963 a_52635_34067.t77 a_52635_49681.t171 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X499 a_101392_n27257# a_100992_n29313.t1 a_100820_n35156.t2 VSS.t331 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X500 VDD.t4454 VDD.t4453 VDD.t4454 VDD.t2729 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X501 a_41891_n29181.t8 a_41891_n29181.t7 a_43817_n28415# VSS.t168 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X502 a_83153_10448.t11 a_83153_10448.t10 a_85089_13546# VDD.t643 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X503 a_47991_4421.t0 a_47819_11614.t8 a_54197_7563# VSS.t304 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X504 VDD.t4452 VDD.t4451 VDD.t4452 VDD.t522 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X505 VDD.t4450 VDD.t4449 VDD.t4450 VDD.t3613 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X506 VDD.t4448 VDD.t4447 VDD.t4448 VDD.t2573 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X507 VDD.t4446 VDD.t4445 VDD.t4446 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X508 a_63683_n19597# a_50751_n19729.t94 a_63161_n19597# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X509 VSS.t3372 VSS.t3371 VSS.t3372 VSS.t638 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X510 a_52635_48695.t76 a_35922_19591.t32 a_52635_34067.t11 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X511 VDD.t4444 VDD.t4443 VDD.t4444 VDD.t2570 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X512 a_106501_n6960# a_71281_n8397.t93 a_105933_n6960# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X513 a_104527_n17715# a_71281_n8397.t94 a_103997_n16810# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X514 a_71281_n8397.t65 a_71281_n8397.t64 VDD.t464 VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X515 a_58851_n1756# a_50751_n19729.t95 a_57977_n5344.t0 VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X516 VDD.t4442 VDD.t4441 VDD.t4442 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X517 OUT.t93 a_35922_19591.t33 a_52635_49681.t14 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X518 a_104527_n15000# a_71281_n8397.t95 a_103997_n15905# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X519 a_47819_n36322.t3 a_47819_n35156.t13 a_49755_n33224# VDD.t2325 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X520 VDD.t4440 VDD.t4439 VDD.t4440 VDD.t619 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X521 a_44885_n5342# a_31953_n19727.t91 VSS.t104 VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X522 VDD.t4438 VDD.t4437 VDD.t4438 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X523 VDD.t4436 VDD.t4435 VDD.t4436 VDD.t507 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X524 a_112199_n18620# a_71281_n8397.t96 a_111631_n18620# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X525 VDD.t4434 VDD.t4433 VDD.t4434 VDD.t1867 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X526 VDD.t4432 VDD.t4431 VDD.t4432 VDD.t508 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X527 VDD.t4430 VDD.t4429 VDD.t4430 VDD.t648 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X528 VSS.t3370 VSS.t3369 VSS.t3370 VSS.t528 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X529 OUT.t18 a_35502_24538.t26 a_33249_35053.t98 VSS.t190 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X530 VDD.t4792 a_47819_n35156.t14 a_48349_n35156# VDD.t2288 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X531 a_33249_48695.t9 a_33379_34007.t11 a_33249_34067.t98 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X532 VSS.t3368 VSS.t3367 VSS.t3368 VSS.t103 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X533 a_104527_n8770# a_71281_n8397.t97 a_103997_n8770.t0 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X534 VDD.t4428 VDD.t4427 VDD.t4428 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X535 a_83153_10448.t9 a_83153_10448.t8 a_85089_11614# VDD.t643 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X536 a_31953_n19727.t65 a_31953_n19727.t64 VSS.t92 VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X537 a_52635_49681.t15 a_35922_19591.t34 OUT.t92 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X538 VDD.t4426 VDD.t4425 VDD.t4426 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X539 VDD.t4424 VDD.t4423 VDD.t4424 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X540 VSS.t3366 VSS.t3365 VSS.t3366 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X541 a_111631_n9675# a_71281_n8397.t98 a_111063_n9675# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X542 a_47753_n14213# a_31953_n19727.t92 a_47231_n14213# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X543 VSS.t3364 VSS.t3363 VSS.t3364 VSS.t979 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X544 VSS.t3362 VSS.t3361 VSS.t3362 VSS.t681 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X545 VDD.t4422 VDD.t4421 VDD.t4422 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X546 a_46879_n19595# a_31953_n19727.t93 a_46319_n18698# VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X547 VDD.t77 a_31699_20742.t63 a_33249_48695.t321 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X548 VDD.t4420 VDD.t4419 VDD.t4420 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X549 a_49795_4481# a_47991_5507.t1 a_48951_4481.t2 VSS.t338 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X550 VDD.t4962 a_52635_34067.t78 a_52635_48695.t167 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X551 a_83709_n19525# a_71281_n10073.t84 a_83141_n19525# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X552 VDD.t4418 VDD.t4417 VDD.t4418 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X553 a_101350_n36322# a_100820_n35156.t13 a_100820_n36322.t1 VDD.t523 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X554 VSS.t3360 VSS.t3359 VSS.t3360 VSS.t553 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X555 VDD.t4416 VDD.t4415 VDD.t4416 VDD.t2099 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X556 VDD.t4414 VDD.t4413 VDD.t4414 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X557 VDD.t4412 VDD.t4411 VDD.t4412 VDD.t638 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X558 a_52635_34067.t12 a_35922_19591.t35 a_52635_48695.t75 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X559 VSS.t3358 VSS.t3357 VSS.t3358 VSS.t868 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X560 VDD.t4410 VDD.t4409 VDD.t4410 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X561 VSS.t3356 VSS.t3355 VSS.t3356 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X562 a_33249_48695.t320 a_31699_20742.t64 VDD.t79 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X563 VDD.t4408 VDD.t4407 VDD.t4408 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X564 VDD.t4961 a_52635_34067.t79 a_52635_49681.t170 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X565 VDD.t4406 VDD.t4405 VDD.t4406 VDD.t501 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X566 a_42047_n4445# a_31953_n19727.t94 a_41487_n4445# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X567 VDD.t4404 VDD.t4403 VDD.t4404 VDD.t625 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X568 VSS.t3354 VSS.t3353 VSS.t3354 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X569 a_106830_10388.t2 a_112559_4481.t12 a_114485_6405# VSS.t292 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X570 VDD.t4793 a_47819_n35156.t15 a_48349_n33224# VDD.t2288 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X571 VSS.t188 a_41891_4481.t12 a_42413_6405# VSS.t166 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X572 a_114485_n27257# a_112559_n29181.t12 VSS.t414 VSS.t413 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X573 a_30152_n35156.t7 a_30152_n35156.t6 a_32088_n36322# VDD.t551 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X574 a_54019_n17803# a_50751_n19729.t96 a_53497_n18700# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X575 a_71896_n35156# a_71496_n36382.t10 a_71366_n35156.t4 VDD.t2251 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X576 a_81735_n7865# a_71281_n10073.t85 a_81205_n7865# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X577 a_105933_n20430# a_71281_n8397.t99 a_105365_n20430# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X578 VDD.t4402 VDD.t4401 VDD.t4402 VDD.t643 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X579 VSS.t3352 VSS.t3351 VSS.t3352 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X580 a_59558_n29181.t1 a_47991_n29313.t1 a_61515_n34390# VDD.t546 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X581 a_32913_n6239# a_31953_n19727.t95 a_32353_n6239# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X582 VDD.t4400 VDD.t4399 VDD.t4400 VDD.t1611 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X583 a_33249_34067.t97 a_33379_34007.t12 a_33249_48695.t109 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X584 a_54197_n30339# a_47819_n36322.t8 a_53675_n30339.t3 VSS.t306 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X585 VDD.t4398 VDD.t4397 VDD.t4398 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X586 a_98829_n7865# a_71281_n8397.t100 a_98299_n7865# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X587 VSS.t3350 VSS.t3349 VSS.t3350 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X588 VDD.t4396 VDD.t4395 VDD.t4396 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X589 VDD.t4394 VDD.t4393 VDD.t4394 VDD.t598 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X590 VSS.t3348 VSS.t3347 VSS.t3348 VSS.t422 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X591 a_33249_34067.t96 a_33379_34007.t13 a_33249_48695.t110 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X592 VDD.t4392 VDD.t4391 VDD.t4392 VDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X593 VSS.t3346 VSS.t3345 VSS.t3346 VSS.t699 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X594 VDD.t4390 VDD.t4389 VDD.t4390 VDD.t625 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X595 a_33249_48695.t319 a_31699_20742.t65 VDD.t80 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X596 VSS.t3344 VSS.t3343 VSS.t3344 VSS.t288 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X597 VSS.t3342 VSS.t3341 VSS.t3342 VSS.t1594 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X598 a_71896_n33224# a_71496_n36382.t11 a_53699_n36322.t2 VDD.t2251 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X599 VSS.t3340 VSS.t3339 VSS.t3340 VSS.t1244 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X600 VSS.t3338 VSS.t3337 VSS.t3338 VSS.t690 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X601 VDD.t4388 VDD.t4387 VDD.t4388 VDD.t1818 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X602 a_96849_n35156# a_89033_n35156.t5 a_96011_n36322.t0 VDD.t2240 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X603 VDD.t4386 VDD.t4385 VDD.t4386 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X604 VSS.t3336 VSS.t3335 VSS.t3336 VSS.t644 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X605 VSS.t3334 VSS.t3333 VSS.t3334 VSS.t1315 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X606 a_33249_35053.t5 a_33379_34917.t8 a_33249_48695.t19 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X607 a_84547_n6960# a_71281_n10073.t86 a_83709_n6960# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X608 VSS.t3332 VSS.t3331 VSS.t3332 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X609 a_104527_n20430# a_71281_n8397.t101 a_53699_n35156.t2 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X610 a_93131_n19525# a_71281_n10073.t87 a_92601_n19525# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X611 a_52635_48695.t166 a_52635_34067.t80 VDD.t4960 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X612 VDD.t4384 VDD.t4383 VDD.t4384 VDD.t2079 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X613 a_60677_n36322.t1 a_53699_n35156.t3 a_60109_n34390# VDD.t545 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X614 a_56895_n16009.t1 a_100992_4421.t0 a_101392_6405# VSS.t162 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X615 VSS.t3330 VSS.t3329 VSS.t3330 VSS.t676 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X616 a_88271_n19525# a_71281_n10073.t88 a_87433_n19525# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X617 VDD.t4382 VDD.t4381 VDD.t4382 VDD.t2076 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X618 VSS.t3328 VSS.t3327 VSS.t3328 VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X619 VDD.t4380 VDD.t4379 VDD.t4380 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X620 VDD.t4978 a_30152_n35156.t13 a_30682_n35156# VDD.t2228 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X621 VDD.t518 a_47819_n36322.t9 a_55601_n29181# VSS.t307 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X622 a_108602_n30339# a_100820_n36322.t9 a_100992_n29313.t0 VSS.t334 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X623 a_45445_n14213# a_31953_n19727.t96 a_44885_n13316# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X624 VSS.t3326 VSS.t3325 VSS.t3326 VSS.t266 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X625 VSS.t3324 VSS.t3323 VSS.t3324 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X626 VDD.t4378 VDD.t4377 VDD.t4378 VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X627 a_113081_6405# a_112559_4481.t6 a_112559_4481.t7 VSS.t293 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X628 a_52635_34067.t13 a_35922_19591.t36 a_52635_48695.t74 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X629 a_96849_n33224# a_89033_n35156.t6 a_96011_n36322.t1 VDD.t2240 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X630 VSS.t3322 VSS.t3321 VSS.t3322 VSS.t721 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X631 a_100235_n14095# a_71281_n8397.t102 a_99667_n14095# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X632 a_65486_11614.t5 a_64243_n1756.t1 a_67462_6405# VSS.t378 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X633 VDD.t4376 VDD.t4375 VDD.t4376 VDD.t1787 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X634 VSS.t3320 VSS.t3319 VSS.t3320 VSS.t498 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X635 a_66551_n13318# a_50751_n19729.t97 a_66029_n14215# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X636 a_39179_n3548# a_31953_n19727.t97 a_38619_n2651# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X637 a_42413_6405# a_41891_4481.t5 a_41891_4481.t6 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X638 VDD.t4374 VDD.t4373 VDD.t4374 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X639 VSS.t3318 VSS.t3317 VSS.t3318 VSS.t681 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X640 a_32353_n14213# a_31953_n19727.t98 a_31831_n15110# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X641 VDD.t4372 VDD.t4371 VDD.t4372 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X642 a_79151_6405# a_77225_4481.t12 VSS.t320 VSS.t319 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X643 VDD.t4370 VDD.t4369 VDD.t4370 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X644 VDD.t4979 a_30152_n35156.t14 a_30682_n33224# VDD.t2228 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X645 a_54229_13546# a_53829_10388.t8 a_53699_13546.t1 VDD.t3678 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X646 OUT.t91 a_35922_19591.t37 a_52635_49681.t16 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X647 a_53699_n35156.t0 a_53829_n36382.t12 a_55635_n35156# VDD.t297 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X648 VDD.t4368 VDD.t4367 VDD.t4368 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X649 VDD.t4366 VDD.t4365 VDD.t4366 VDD.t2061 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X650 a_32353_n1754# a_31953_n19727.t99 a_31831_n2651# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X651 VSS.t3316 VSS.t3315 VSS.t3316 VSS.t423 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X652 VDD.t4364 VDD.t4363 VDD.t4364 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X653 VSS.t3314 VSS.t3313 VSS.t3314 VSS.t609 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X654 VSS.t3312 VSS.t3311 VSS.t3312 VSS.t12 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X655 VSS.t3310 VSS.t3309 VSS.t3310 VSS.t183 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X656 VDD.t4362 VDD.t4361 VDD.t4362 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X657 a_34347_n2651# a_31953_n19727.t100 a_33787_n1754# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X658 a_90935_4481# a_83153_11614.t11 a_83325_4421.t0 VSS.t395 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X659 a_41487_n16904# a_31953_n19727.t101 a_40965_n16904# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X660 a_35781_n7136# a_31953_n19727.t102 a_35221_n6239# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X661 a_33249_48695.t318 a_31699_20742.t66 VDD.t81 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X662 VSS.t3308 VSS.t3307 VSS.t3308 VSS.t908 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X663 a_52635_49681.t169 a_52635_34067.t81 VDD.t4959 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X664 a_52635_34067.t14 a_35922_19591.t38 a_52635_48695.t73 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X665 a_113037_n17715# a_71281_n8397.t103 a_78344_n36322.t0 VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X666 VDD.t4360 VDD.t4359 VDD.t4360 VDD.t32 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X667 a_98829_n14095# a_71281_n8397.t104 VDD.t473 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X668 a_93131_n7865# a_71281_n10073.t89 a_92601_n7865# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X669 a_50751_n19729.t65 a_50751_n19729.t64 VSS.t251 VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X670 VSS.t3306 VSS.t3305 VSS.t3306 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X671 VDD.t4358 VDD.t4357 VDD.t4358 VDD.t1419 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X672 a_52635_34067.t15 a_35922_19591.t39 a_52635_48695.t72 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X673 a_113037_n15000# a_71281_n8397.t105 a_112199_n15000# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X674 a_33249_48695.t317 a_31699_20742.t67 VDD.t83 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X675 VDD.t4356 VDD.t4355 VDD.t4356 VDD.t2485 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X676 a_54229_11614# a_53829_10388.t9 a_53699_11614.t2 VDD.t3678 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X677 VSS.t3304 VSS.t3303 VSS.t3304 VSS.t354 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X678 a_52635_48695.t165 a_52635_34067.t82 VDD.t4958 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X679 a_53699_n36322.t1 a_53829_n36382.t13 a_55635_n33224# VDD.t297 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X680 VDD.t4354 VDD.t4353 VDD.t4354 VDD.t976 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X681 VSS.t3302 VSS.t3301 VSS.t3302 VSS.t1157 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X682 VDD.t84 a_31699_20742.t68 a_33249_48695.t316 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X683 a_83141_n18620# a_71281_n10073.t90 a_82573_n18620# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X684 VSS.t3300 VSS.t3299 VSS.t3300 VSS.t553 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X685 a_105365_n14095# a_71281_n8397.t106 a_104527_n14095# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X686 a_66058_4481# a_65658_4421.t1 a_65486_10448.t10 VSS.t376 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X687 VDD.t4352 VDD.t4351 VDD.t4352 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X688 VDD.t4350 VDD.t4349 VDD.t4350 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X689 a_83153_n35156.t10 a_83325_n29313.t0 a_85129_n30339# VSS.t285 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X690 a_105933_n15905# a_71281_n8397.t107 a_105365_n15905# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X691 a_72603_n10073# I1N.t4 a_71281_n10073.t72 VSS.t429 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X692 a_95105_n13190# a_71281_n10073.t91 a_94537_n13190# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X693 VDD.t85 a_31699_20742.t69 a_33249_48695.t315 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X694 VDD.t4348 VDD.t4347 VDD.t4348 VDD.t1419 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X695 a_52635_34067.t16 a_35922_19591.t40 a_52635_48695.t71 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X696 a_89715_n16810.t1 a_71281_n10073.t92 a_89407_n13190# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X697 VDD.t4346 VDD.t4345 VDD.t4346 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X698 VDD.t4344 VDD.t4343 VDD.t4344 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X699 a_57417_n15112# a_50751_n19729.t98 a_56895_n15112# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X700 a_53829_n36382.t0 a_59558_n29181.t11 a_61484_n27257# VSS.t398 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X701 a_95943_n6960# a_71281_n10073.t93 a_95105_n6960# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X702 VDD.t4342 VDD.t4341 VDD.t4342 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X703 VSS.t3298 VSS.t3297 VSS.t3298 VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X704 a_44885_n16904# a_31953_n19727.t103 a_44363_n17801# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X705 VDD.t41 a_31699_20742.t37 a_31699_20742.t38 VDD.t16 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X706 VDD.t4340 VDD.t4339 VDD.t4340 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X707 VDD.t86 a_31699_20742.t70 a_33249_48695.t314 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X708 VDD.t4338 VDD.t4337 VDD.t4338 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X709 a_52635_34067.t17 a_35922_19591.t41 a_52635_48695.t70 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X710 OUT.t90 a_35922_19591.t42 a_52635_49681.t17 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X711 VSS.t3296 VSS.t3295 VSS.t3296 VSS.t65 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X712 a_81735_n18620# a_71281_n10073.t94 a_81205_n19525# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X713 VDD.t4336 VDD.t4335 VDD.t4336 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X714 VSS.t91 a_31953_n19727.t62 a_31953_n19727.t63 VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X715 VSS.t3294 VSS.t3293 VSS.t3294 VSS.t615 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X716 VDD.t4334 VDD.t4333 VDD.t4334 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X717 a_57417_n4447# a_50751_n19729.t99 a_56895_n4447# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X718 VDD.t4332 VDD.t4331 VDD.t4332 VDD.t638 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X719 a_33249_35053.t6 a_33379_34917.t9 a_33249_48695.t20 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X720 a_93969_n8770# a_71281_n10073.t95 a_93131_n8770# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X721 VDD.t4330 VDD.t4329 VDD.t4330 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X722 VDD.t4328 VDD.t4327 VDD.t4328 VDD.t1515 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X723 a_104527_n15905# a_71281_n8397.t108 a_103997_n15905# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X724 a_112199_n4245# a_71281_n8397.t109 a_111631_n4245# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X725 VSS.t3292 VSS.t3291 VSS.t3292 VSS.t1256 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X726 VDD.t4326 VDD.t4325 VDD.t4326 VDD.t944 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X727 VDD.t4324 VDD.t4323 VDD.t4324 VDD.t1373 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X728 VDD.t327 a_30152_10448.t12 a_30682_12380# VDD.t326 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X729 VDD.t4322 VDD.t4321 VDD.t4322 VDD.t1370 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X730 a_51151_n13318# a_50751_n19729.t100 a_50629_n13318# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X731 a_71896_13546# a_71496_10388.t10 a_71366_13546.t3 VDD.t351 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X732 VDD.t4320 VDD.t4319 VDD.t4320 VDD.t1365 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X733 VSS.t3290 VSS.t3289 VSS.t3290 VSS.t795 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X734 a_94537_n3340# a_71281_n10073.t96 a_93969_n3340# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X735 a_96849_12380# a_81205_n14095.t3 a_84017_n17715.t4 VDD.t499 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X736 VDD.t4318 VDD.t4317 VDD.t4318 VDD.t78 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X737 a_42413_n30339# a_41891_n29181.t12 a_36162_n36382.t2 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X738 a_88839_n13190# a_71281_n10073.t97 a_88271_n13190# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X739 a_73302_10448# a_71496_10388.t11 a_71342_7563.t2 VDD.t363 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X740 VDD.t4316 VDD.t4315 VDD.t4316 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X741 VDD.t463 a_71281_n8397.t62 a_71281_n8397.t63 VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X742 VDD.t4314 VDD.t4313 VDD.t4314 VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X743 VSS.t3288 VSS.t3287 VSS.t3288 VSS.t604 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X744 a_104527_n7865# a_71281_n8397.t110 a_103997_n7865# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X745 a_52635_34067.t18 a_35922_19591.t43 a_52635_48695.t69 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X746 a_82573_n9675# a_71281_n10073.t98 a_81735_n9675# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X747 OUT.t89 a_35922_19591.t44 a_52635_49681.t18 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X748 a_75585_n9297# I1N.t5 VSS.t431 VSS.t430 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X749 VSS.t3286 VSS.t3285 VSS.t3286 VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X750 a_113037_n20430# a_71281_n8397.t111 a_112199_n20430# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X751 a_65486_n36322.t0 a_65486_n35156.t13 a_67422_n35156# VDD.t1 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X752 VDD.t4312 VDD.t4311 VDD.t4312 VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X753 VDD.t4310 VDD.t4309 VDD.t4310 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X754 VDD.t4308 VDD.t4307 VDD.t4308 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X755 a_50751_n19729.t63 a_50751_n19729.t62 VSS.t250 VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X756 OUT.t88 a_35922_19591.t45 a_52635_49681.t19 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X757 VDD.t4306 VDD.t4305 VDD.t4306 VDD.t1354 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X758 a_99667_n9675# a_71281_n8397.t112 a_98829_n9675# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X759 a_71896_11614# a_71496_10388.t12 a_71366_11614.t2 VDD.t351 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X760 a_102756_n34390# a_100820_n35156.t14 VDD.t525 VDD.t524 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X761 a_34347_n13316# a_31953_n19727.t104 a_33787_n12419# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X762 a_52635_48695.t68 a_35922_19591.t46 a_52635_34067.t19 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X763 a_33249_35053.t7 a_33379_34917.t10 a_33249_48695.t21 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X764 a_95414_n28415# a_94892_n29181.t11 a_89163_n36382.t0 VSS.t353 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X765 VDD.t4304 VDD.t4303 VDD.t4304 VDD.t1349 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X766 a_94892_n29181.t4 a_94892_n29181.t3 a_96818_n30339# VSS.t352 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X767 a_33249_34067.t95 a_33379_34007.t14 a_33249_48695.t157 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X768 VSS.t3284 VSS.t3283 VSS.t3284 VSS.t979 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X769 VSS.t3282 VSS.t3281 VSS.t3282 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X770 VDD.t4302 VDD.t4301 VDD.t4302 VDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X771 VDD.t4300 VDD.t4299 VDD.t4300 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X772 a_30152_10448.t0 a_30324_4421.t0 a_32128_5639# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X773 a_35502_25545.t4 a_31699_20742.t71 VDD.t87 VDD.t20 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X774 a_33249_35053.t8 a_33379_34917.t11 a_33249_48695.t22 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X775 VDD.t503 a_47819_11614.t9 a_55601_6405# VSS.t307 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X776 VDD.t4298 VDD.t4297 VDD.t4298 VDD.t1711 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X777 VDD.t4296 VDD.t4295 VDD.t4296 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X778 VDD.t4294 VDD.t4293 VDD.t4294 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X779 VSS.t3280 VSS.t3279 VSS.t3280 VSS.t550 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X780 VDD.t375 a_71281_n10073.t70 a_71281_n10073.t71 VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X781 a_46319_n17801# a_31953_n19727.t105 a_45797_n18698# VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X782 a_65486_n36322.t1 a_65486_n35156.t14 a_67422_n33224# VDD.t1 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X783 a_40613_n8930# a_31953_n19727.t106 a_40053_n8033# VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X784 VDD.t4292 VDD.t4291 VDD.t4292 VDD.t2777 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X785 VSS.t3278 VSS.t3277 VSS.t3278 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X786 VDD.t4 a_65486_n35156.t15 a_66016_n35156# VDD.t2 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X787 VSS.t3276 VSS.t3275 VSS.t3276 VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X788 VSS.t3274 VSS.t3273 VSS.t3274 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X789 a_33249_35053.t9 a_33379_34917.t12 a_33249_48695.t23 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X790 VDD.t4290 VDD.t4289 VDD.t4290 VDD.t2559 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X791 a_57977_n8932# a_50751_n19729.t101 a_57417_n8932# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X792 a_79182_13546# a_65658_4421.t2 a_78344_10448.t5 VDD.t571 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X793 VDD.t4288 VDD.t4287 VDD.t4288 VDD.t955 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X794 VSS.t3272 VSS.t3271 VSS.t3272 VSS.t1126 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X795 VSS.t3270 VSS.t3269 VSS.t3270 VSS.t1034 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X796 VSS.t3268 VSS.t3267 VSS.t3268 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X797 a_43817_n29181# a_41891_n29181.t13 VSS.t369 VSS.t158 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X798 VDD.t4286 VDD.t4285 VDD.t4286 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X799 VDD.t4284 VDD.t4283 VDD.t4284 VDD.t49 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X800 VDD.t4282 VDD.t4281 VDD.t4282 VDD.t898 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X801 a_33249_48695.t158 a_33379_34007.t15 a_33249_34067.t94 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X802 VDD.t88 a_31699_20742.t72 a_35502_24538.t22 VDD.t25 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X803 VSS.t3266 VSS.t3265 VSS.t3266 VSS.t182 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X804 VDD.t4280 VDD.t4279 VDD.t4280 VDD.t2777 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X805 VDD.t4278 VDD.t4277 VDD.t4278 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X806 a_40053_n7136# a_31953_n19727.t107 a_39531_n8033# VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X807 a_49795_n29181# a_39179_n19595.t2 a_38097_n16007.t1 VSS.t338 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X808 VDD.t5 a_65486_n35156.t16 a_66016_n33224# VDD.t2 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X809 a_71281_n10073.t69 a_71281_n10073.t68 VDD.t362 VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X810 VDD.t4957 a_52635_34067.t83 a_52635_49681.t168 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X811 a_31831_n5342.t2 a_83325_n29313.t2 a_83725_n27257# VSS.t288 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X812 VSS.t3264 VSS.t3263 VSS.t3264 VSS.t14 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X813 VDD.t4956 a_52635_34067.t84 a_52635_48695.t164 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X814 OUT.t87 a_35922_19591.t47 a_52635_49681.t20 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X815 VDD.t4276 VDD.t4275 VDD.t4276 VDD.t12 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X816 VDD.t4274 VDD.t4273 VDD.t4274 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X817 VDD.t89 a_31699_20742.t73 a_33249_48695.t313 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X818 VSS.t3262 VSS.t3261 VSS.t3262 VSS.t1111 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X819 VSS.t3260 VSS.t3259 VSS.t3260 VSS.t464 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X820 a_60080_n30339# a_59558_n29181.t12 a_53829_n36382.t1 VSS.t397 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X821 a_54197_4481# a_47819_11614.t10 a_53675_4481.t2 VSS.t306 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X822 a_112199_n21335# a_71281_n8397.t113 a_111631_n21335# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X823 a_102796_5639# a_100992_4421.t0 a_56895_n16009.t1 VSS.t172 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X824 VSS.t3258 VSS.t3257 VSS.t3258 VSS.t37 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X825 VSS.t3256 VSS.t3255 VSS.t3256 VSS.t185 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X826 a_93969_n19525# a_71281_n10073.t99 a_93131_n19525# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X827 VDD.t4272 VDD.t4271 VDD.t4272 VDD.t955 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X828 VDD.t4270 VDD.t4269 VDD.t4270 VDD.t1917 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X829 a_79182_11614# a_65658_4421.t2 a_78344_10448.t2 VDD.t571 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X830 a_52635_34067.t20 a_35922_19591.t48 a_52635_48695.t67 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X831 OUT.t86 a_35922_19591.t49 a_52635_49681.t21 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X832 a_40613_n14213# a_31953_n19727.t108 a_41487_n16007# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X833 VDD.t4268 VDD.t4267 VDD.t4268 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X834 a_41487_n7136# a_31953_n19727.t109 a_40965_n8033# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X835 a_35781_n19595# a_31953_n19727.t110 a_35221_n18698# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X836 VSS.t3254 VSS.t3253 VSS.t3254 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X837 a_32088_n35156# a_30152_n35156.t15 VDD.t4980 VDD.t2088 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X838 a_35221_n6239# a_31953_n19727.t111 a_34699_n6239# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X839 a_53675_n30339.t0 a_53829_n36382.t14 a_54229_n36322# VDD.t301 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X840 a_55601_6405# a_47819_11614.t11 a_47991_5507.t1 VSS.t305 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X841 VDD.t4266 VDD.t4265 VDD.t4266 VDD.t1904 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X842 VDD.t4264 VDD.t4263 VDD.t4264 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X843 a_71281_n8397.t61 a_71281_n8397.t60 VDD.t462 VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X844 VSS.t3252 VSS.t3251 VSS.t3252 VSS.t591 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X845 VSS.t3250 VSS.t3249 VSS.t3250 VSS.t475 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X846 a_87433_n3340# a_71281_n10073.t100 a_86903_n4245# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X847 VSS.t3248 VSS.t3247 VSS.t3248 VSS.t103 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X848 VDD.t4262 VDD.t4261 VDD.t4262 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X849 a_106501_n15000# a_71281_n8397.t114 a_105933_n15000# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X850 a_89563_10448# a_89163_10388.t11 a_71366_13546.t1 VDD.t552 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X851 a_67422_10448# a_65486_10448.t13 VDD.t4747 VDD.t866 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X852 VSS.t3246 VSS.t3245 VSS.t3246 VSS.t588 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X853 a_36162_10388.t5 a_36032_11614.t5 a_43848_12380# VDD.t287 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X854 VDD.t4260 VDD.t4259 VDD.t4260 VDD.t547 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X855 VDD.t4258 VDD.t4257 VDD.t4258 VDD.t2349 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X856 VSS.t3244 VSS.t3243 VSS.t3244 VSS.t1615 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X857 VSS.t3242 VSS.t3241 VSS.t3242 VSS.t495 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X858 VSS.t3240 VSS.t3239 VSS.t3240 VSS.t681 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X859 a_43010_10448.t1 a_30324_4421.t1 a_42442_10448# VDD.t289 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X860 a_101641_n6960# a_71281_n8397.t115 a_100803_n6960# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X861 a_32088_n33224# a_30152_n35156.t16 VDD.t4981 VDD.t2088 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X862 VSS.t3238 VSS.t3237 VSS.t3238 VSS.t1821 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X863 VDD.t4256 VDD.t4255 VDD.t4256 VDD.t1893 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X864 VDD.t4254 VDD.t4253 VDD.t4254 VDD.t855 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X865 a_113037_n18620# a_71281_n8397.t116 a_112199_n15905# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X866 VSS.t249 a_50751_n19729.t60 a_50751_n19729.t61 VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X867 OUT.t85 a_35922_19591.t50 a_52635_49681.t22 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X868 VDD.t373 a_71281_n10073.t66 a_71281_n10073.t67 VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X869 a_32913_n5342.t0 a_31953_n19727.t112 a_32353_n5342# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X870 VSS.t3236 VSS.t3235 VSS.t3236 VSS.t478 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X871 a_52635_48695.t163 a_52635_34067.t85 VDD.t4955 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X872 VSS.t3234 VSS.t3233 VSS.t3234 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X873 a_33249_48695.t0 a_33379_34007.t16 a_33249_34067.t93 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X874 a_52635_34067.t58 a_35502_24538.t27 a_33249_34067.t16 VSS.t190 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X875 VDD.t4252 VDD.t4251 VDD.t4252 VDD.t1884 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X876 VDD.t366 a_71281_n10073.t64 a_71281_n10073.t65 VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X877 a_50751_n19729.t59 a_50751_n19729.t58 VSS.t248 VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X878 VDD.t4250 VDD.t4249 VDD.t4250 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X879 VDD.t4248 VDD.t4247 VDD.t4248 VDD.t667 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X880 VSS.t3232 VSS.t3231 VSS.t3232 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X881 VSS.t3230 VSS.t3229 VSS.t3230 VSS.t60 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X882 VDD.t4246 VDD.t4245 VDD.t4246 VDD.t828 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X883 VDD.t4244 VDD.t4243 VDD.t4244 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X884 a_71366_n35156.t2 a_71496_n36382.t12 a_73302_n35156# VDD.t2058 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X885 VDD.t4242 VDD.t4241 VDD.t4242 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X886 VDD.t4240 VDD.t4239 VDD.t4240 VDD.t813 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X887 a_45138_23609# a_35922_19591.t51 a_44608_22884# VDD.t405 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X888 VDD.t4238 VDD.t4237 VDD.t4238 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X889 VSS.t3228 VSS.t3227 VSS.t3228 VSS.t501 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X890 a_41891_4481.t8 a_41891_4481.t7 a_43817_7563# VSS.t168 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X891 VSS.t3226 VSS.t3225 VSS.t3226 VSS.t1157 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X892 VDD.t4236 VDD.t4235 VDD.t4236 VDD.t667 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X893 VDD.t4234 VDD.t4233 VDD.t4234 VDD.t2680 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X894 OUT.t84 a_35922_19591.t52 a_52635_49681.t23 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X895 VDD.t4232 VDD.t4231 VDD.t4232 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X896 VSS.t3224 VSS.t3223 VSS.t3224 VSS.t976 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X897 a_78344_n36322.t2 a_65658_n29313.t1 a_77776_n35156# VDD.t502 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X898 VSS.t3222 VSS.t3221 VSS.t3222 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X899 a_66058_n29181# a_65658_n29313.t0 a_65486_n35156.t8 VSS.t376 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X900 VSS.t3220 VSS.t3219 VSS.t3220 VSS.t490 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X901 a_81735_n17715# a_71281_n10073.t101 a_81205_n21335# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X902 a_39179_n16007.t1 a_31953_n19727.t113 a_38619_n16007# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X903 a_33249_34067.t92 a_33379_34007.t17 a_33249_48695.t1 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X904 a_33249_48695.t312 a_31699_20742.t74 VDD.t90 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X905 a_71366_n36322.t0 a_71496_n36382.t13 a_73302_n33224# VDD.t2058 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X906 a_52635_49681.t167 a_52635_34067.t86 VDD.t4954 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X907 VDD.t4230 VDD.t4229 VDD.t4230 VDD.t635 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X908 a_93969_n7865# a_71281_n10073.t102 a_93131_n7865# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X909 a_33249_48695.t311 a_31699_20742.t75 VDD.t91 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X910 VSS.t3218 VSS.t3217 VSS.t3218 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X911 VSS.t90 a_31953_n19727.t60 a_31953_n19727.t61 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X912 a_33249_34067.t91 a_33379_34007.t18 a_33249_48695.t5 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X913 VSS.t3216 VSS.t3215 VSS.t3216 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X914 VSS.t364 a_71496_n36382.t14 a_71896_n35156# VDD.t2021 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X915 a_48313_n2651# a_31953_n19727.t114 a_47753_n1754# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X916 a_106501_n20430# a_71281_n8397.t117 a_105933_n20430# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X917 a_33787_n13316# a_31953_n19727.t115 a_33265_n14213# VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X918 VSS.t3214 VSS.t3213 VSS.t3214 VSS.t155 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X919 a_66551_n12421# a_50751_n19729.t102 VSS.t267 VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X920 VSS.t3212 VSS.t3211 VSS.t3212 VSS.t534 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X921 a_60285_n16009# a_50751_n19729.t103 a_59411_n14215# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X922 a_94537_n2435# a_71281_n10073.t103 a_93969_n2435# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X923 VDD.t4228 VDD.t4227 VDD.t4228 VDD.t1850 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X924 VDD.t4226 VDD.t4225 VDD.t4226 VDD.t417 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X925 VSS.t3210 VSS.t3209 VSS.t3210 VSS.t149 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X926 a_45445_n6239# a_31953_n19727.t116 a_44885_n4445# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X927 VDD.t4224 VDD.t4223 VDD.t4224 VDD.t2680 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X928 a_78344_n36322.t2 a_65658_n29313.t1 a_77776_n33224# VDD.t502 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X929 VSS.t3208 VSS.t3207 VSS.t3208 VSS.t531 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X930 VDD.t4222 VDD.t4221 VDD.t4222 VDD.t337 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X931 a_59558_n29181.t2 a_47991_n29313.t1 a_61515_n36322# VDD.t546 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X932 VDD.t4220 VDD.t4219 VDD.t4220 VDD.t1611 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X933 VDD.t4218 VDD.t4217 VDD.t4218 VDD.t792 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X934 VDD.t4216 VDD.t4215 VDD.t4216 VDD.t610 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X935 VDD.t4214 VDD.t4213 VDD.t4214 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X936 a_64243_n6241# a_50751_n19729.t104 a_63683_n4447# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X937 VDD.t4212 VDD.t4211 VDD.t4212 VDD.t635 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X938 a_51711_n19597# a_50751_n19729.t105 a_51151_n19597# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X939 a_100820_10448.t1 a_100992_4421.t0 a_102796_7563# VSS.t171 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X940 VDD.t4210 VDD.t4209 VDD.t4210 VDD.t507 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X941 a_31284_4481.t2 a_30324_5507.t1 a_30724_7563# VSS.t151 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X942 VSS.t3206 VSS.t3205 VSS.t3206 VSS.t411 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X943 VSS.t3204 VSS.t3203 VSS.t3204 VSS.t129 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X944 a_71342_n27257.t0 a_71496_n36382.t15 a_71896_n33224# VDD.t2021 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X945 a_33249_34067.t90 a_33379_34007.t19 a_33249_48695.t6 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X946 a_34347_n3548# a_31953_n19727.t117 a_35221_n5342# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X947 VSS.t3202 VSS.t3201 VSS.t3202 VSS.t148 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X948 a_89163_n36382.t4 a_89033_n35156.t7 a_96849_n35156# VDD.t1996 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X949 VSS.t3200 VSS.t3199 VSS.t3200 VSS.t478 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X950 a_40613_n3548# a_31953_n19727.t118 a_40053_n3548# VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X951 VDD.t4208 VDD.t4207 VDD.t4208 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X952 VDD.t4206 VDD.t4205 VDD.t4206 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X953 a_83141_n21335# a_71281_n10073.t104 a_82573_n21335# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X954 VDD.t4204 VDD.t4203 VDD.t4204 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X955 a_50751_n19729.t57 a_50751_n19729.t56 VSS.t247 VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X956 VDD.t4202 VDD.t4201 VDD.t4202 VDD.t1824 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X957 a_52635_34067.t12 a_35922_19591.t53 a_52635_48695.t66 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X958 VDD.t4200 VDD.t4199 VDD.t4200 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X959 VDD.t4198 VDD.t4197 VDD.t4198 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X960 VDD.t4196 VDD.t4195 VDD.t4196 VDD.t1821 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X961 VSS.t3198 VSS.t3197 VSS.t3198 VSS.t459 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X962 a_52635_34067.t21 a_35922_19591.t54 a_52635_48695.t65 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X963 a_33249_34067.t89 a_33379_34007.t20 a_33249_48695.t7 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X964 a_111063_n8770# a_71281_n8397.t118 a_110225_n8770# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X965 VSS.t3196 VSS.t3195 VSS.t3196 VSS.t229 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X966 a_85129_5639# a_83325_4421.t0 a_50629_n16009.t1 VSS.t309 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X967 VDD.t4194 VDD.t4193 VDD.t4194 VDD.t610 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X968 VDD.t4192 VDD.t4191 VDD.t4192 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X969 a_43817_7563# a_41891_4481.t13 VSS.t159 VSS.t158 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X970 VDD.t4190 VDD.t4189 VDD.t4190 VDD.t2231 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X971 VDD.t92 a_31699_20742.t76 a_33249_48695.t310 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X972 a_60677_n36322.t2 a_53699_n35156.t4 a_60109_n36322# VDD.t545 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X973 a_83709_n4245# a_71281_n10073.t105 a_83141_n4245# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X974 a_32088_12380# a_30152_10448.t13 VDD.t304 VDD.t303 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X975 OUT.t83 a_35922_19591.t55 a_52635_49681.t24 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X976 a_38097_n5342.t2 a_39179_n8930.t1 a_101392_n30339# VSS.t332 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X977 VSS.t3194 VSS.t3193 VSS.t3194 VSS.t1037 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X978 a_111631_n3340# a_71281_n8397.t119 a_111063_n3340# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X979 VDD.t4188 VDD.t4187 VDD.t4188 VDD.t535 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X980 a_89163_n36382.t5 a_89033_n35156.t8 a_96849_n33224# VDD.t1996 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X981 VSS.t3192 VSS.t3191 VSS.t3192 VSS.t487 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X982 VSS.t3190 VSS.t3189 VSS.t3190 VSS.t284 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X983 VDD.t4186 VDD.t4185 VDD.t4186 VDD.t1209 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X984 VDD.t4184 VDD.t4183 VDD.t4184 VDD.t755 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X985 VDD.t4182 VDD.t4181 VDD.t4182 VDD.t2422 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X986 VSS.t3188 VSS.t3187 VSS.t3188 VSS.t947 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X987 a_81735_n21335# a_71281_n10073.t106 a_81205_n21335# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X988 VSS.t3186 VSS.t3185 VSS.t3186 VSS.t937 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X989 VDD.t4180 VDD.t4179 VDD.t4180 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X990 VDD.t4178 VDD.t4177 VDD.t4178 VDD.t1796 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X991 a_87433_n19525# a_71281_n10073.t107 a_86903_n19525# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X992 VSS.t3184 VSS.t3183 VSS.t3184 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X993 VSS.t3182 VSS.t3181 VSS.t3182 VSS.t229 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X994 VSS.t3180 VSS.t3179 VSS.t3180 VSS.t1025 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X995 a_101392_7563# a_57977_n12421.t0 a_100820_11614.t6 VSS.t163 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X996 a_33249_34067.t141 a_35502_25545.t31 VSS.t204 VSS.t31 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X997 VSS.t3178 VSS.t3177 VSS.t3178 VSS.t168 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X998 VDD.t4176 VDD.t4175 VDD.t4176 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X999 a_81735_n1530# a_71281_n10073.t108 a_81205_n5150# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1000 a_33249_48695.t106 a_33379_34007.t21 a_33249_34067.t88 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1001 a_45445_n19595.t1 a_65486_n36322.t10 a_71864_n28415# VSS.t157 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1002 VDD.t4174 VDD.t4173 VDD.t4174 VDD.t755 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1003 VSS.t3176 VSS.t3175 VSS.t3176 VSS.t868 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1004 a_33249_35053.t10 a_33379_34917.t13 a_33249_48695.t24 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1005 a_30724_7563# a_30324_5507.t1 a_30152_11614.t3 VSS.t150 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1006 VDD.t4172 VDD.t4171 VDD.t4172 VDD.t1780 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1007 a_73268_n30339# a_65486_n36322.t11 a_65658_n29313.t0 VSS.t154 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1008 VDD.t4953 a_52635_34067.t87 a_52635_48695.t162 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1009 a_98829_n1530# a_71281_n8397.t120 a_98299_n5150# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1010 a_51151_n12421# a_50751_n19729.t106 a_50629_n13318# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1011 VDD.t4170 VDD.t4169 VDD.t4170 VDD.t1333 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1012 VDD.t4168 VDD.t4167 VDD.t4168 VDD.t1262 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1013 a_71281_n8397.t59 a_71281_n8397.t58 VDD.t461 VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1014 a_52635_49681.t166 a_52635_34067.t88 VDD.t4952 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1015 VDD.t4166 VDD.t4165 VDD.t4166 VDD.t748 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1016 VDD.t4164 VDD.t4163 VDD.t4164 VDD.t1338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1017 a_65677_n17803# a_50751_n19729.t107 a_65117_n17803# VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1018 VDD.t4162 VDD.t4161 VDD.t4162 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1019 VDD.t4160 VDD.t4159 VDD.t4160 VDD.t1183 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1020 a_33249_48695.t309 a_31699_20742.t77 VDD.t93 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1021 a_52635_49681.t165 a_52635_34067.t89 VDD.t4951 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1022 a_105933_n14095# a_71281_n8397.t121 a_105365_n14095# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1023 VSS.t3174 VSS.t3173 VSS.t3174 VSS.t596 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1024 VDD.t4158 VDD.t4157 VDD.t4158 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1025 VDD.t4156 VDD.t4155 VDD.t4156 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1026 a_52635_48695.t161 a_52635_34067.t90 VDD.t4950 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1027 a_30724_n28415# a_30324_n30399.t1 a_30152_n36322.t3 VSS.t150 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1028 VSS.t3172 VSS.t3171 VSS.t3172 VSS.t105 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1029 a_106501_n15905# a_71281_n8397.t122 a_105933_n15905# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1030 a_61484_n29181# a_59558_n29181.t13 VSS.t444 VSS.t399 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1031 a_108636_10448# a_106830_10388.t11 a_106676_7563.t0 VDD.t520 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1032 a_33249_34067.t140 a_35502_25545.t32 VSS.t179 VSS.t16 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1033 VDD.t4154 VDD.t4153 VDD.t4154 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1034 a_87433_n2435# a_71281_n10073.t109 a_53699_11614.t0 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1035 VDD.t4152 VDD.t4151 VDD.t4152 VDD.t1177 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1036 VSS.t3170 VSS.t3169 VSS.t3170 VSS.t190 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1037 VDD.t4150 VDD.t4149 VDD.t4150 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1038 a_52635_48695.t160 a_52635_34067.t91 VDD.t4949 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1039 a_100820_n36322.t5 a_39179_n8930.t1 a_102796_n29181# VSS.t329 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1040 VDD.t4148 VDD.t4147 VDD.t4148 VDD.t725 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1041 VSS.t3168 VSS.t3167 VSS.t3168 VSS.t998 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1042 VDD.t4146 VDD.t4145 VDD.t4146 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1043 VSS.t3166 VSS.t3165 VSS.t3166 VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1044 a_60285_n8932# a_50751_n19729.t108 a_57977_n8932# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1045 VDD.t4948 a_52635_34067.t92 a_52635_49681.t164 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1046 VDD.t4144 VDD.t4143 VDD.t4144 VDD.t1373 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1047 a_35221_n17801# a_31953_n19727.t119 a_34699_n18698# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1048 VDD.t4142 VDD.t4141 VDD.t4142 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1049 VDD.t460 a_71281_n8397.t56 a_71281_n8397.t57 VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1050 VSS.t3164 VSS.t3163 VSS.t3164 VSS.t837 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1051 VSS.t3162 VSS.t3161 VSS.t3162 VSS.t588 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1052 a_104527_n14095# a_71281_n8397.t123 VDD.t475 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1053 VDD.t4140 VDD.t4139 VDD.t4140 VDD.t429 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1054 VDD.t4138 VDD.t4137 VDD.t4138 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1055 a_95105_n4245# a_71281_n10073.t110 a_94537_n4245# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1056 a_33249_48695.t308 a_31699_20742.t78 VDD.t94 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1057 VDD.t4136 VDD.t4135 VDD.t4136 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1058 a_30324_n29313.t0 a_30152_n36322.t9 a_36530_n30339# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1059 VDD.t4134 VDD.t4133 VDD.t4134 VDD.t1299 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1060 VSS.t3160 VSS.t3159 VSS.t3160 VSS.t834 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1061 VSS.t3158 VSS.t3157 VSS.t3158 VSS.t1064 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1062 VDD.t95 a_31699_20742.t79 a_33249_48695.t307 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1063 VDD.t4132 VDD.t4131 VDD.t4132 VDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1064 VDD.t4130 VDD.t4129 VDD.t4130 VDD.t697 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1065 VDD.t4947 a_52635_34067.t93 a_52635_49681.t163 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1066 VDD.t4128 VDD.t4127 VDD.t4128 VDD.t1515 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1067 a_89407_n13190# a_71281_n10073.t111 a_88839_n13190# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1068 a_54019_n13318# a_50751_n19729.t109 a_53497_n14215# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1069 VSS.t3156 VSS.t3155 VSS.t3156 VSS.t1360 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1070 VSS.t3154 VSS.t3153 VSS.t3154 VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1071 VDD.t4126 VDD.t4125 VDD.t4126 VDD.t2777 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1072 VSS.t3152 VSS.t3151 VSS.t3152 VSS.t68 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1073 VDD.t97 a_31699_20742.t80 a_33249_48695.t306 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1074 a_103997_n8770.t1 a_106830_n36382.t8 a_108636_n34390# VDD.t1290 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1075 VDD.t4124 VDD.t4123 VDD.t4124 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1076 a_36008_7563.t1 a_36162_10388.t8 a_36562_13546# VDD.t3613 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1077 VDD.t4122 VDD.t4121 VDD.t4122 VDD.t2573 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1078 VDD.t4120 VDD.t4119 VDD.t4120 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1079 a_100803_n13190# a_71281_n8397.t124 a_100235_n13190# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1080 a_32913_n8930.t1 a_83153_n36322.t9 a_89531_n28415# VSS.t453 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1081 VDD.t4118 VDD.t4117 VDD.t4118 VDD.t2570 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1082 VDD.t4946 a_52635_34067.t94 a_52635_48695.t159 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1083 a_40613_n19595# a_31953_n19727.t120 a_40053_n19595# VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1084 VSS.t3150 VSS.t3149 VSS.t3150 VSS.t537 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1085 a_93131_n1530# a_71281_n10073.t112 a_92601_n5150# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1086 a_43848_10448# a_36032_11614.t6 a_43010_10448.t1 VDD.t290 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1087 VDD.t4116 VDD.t4115 VDD.t4116 VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1088 a_107198_n29181# a_100820_n36322.t10 VDD.t539 VSS.t335 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1089 a_83325_4421.t0 a_83153_11614.t12 a_89531_7563# VSS.t393 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1090 VDD.t4114 VDD.t4113 VDD.t4114 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1091 a_73268_5639# a_65486_11614.t8 a_64243_n1756.t1 VSS.t421 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1092 VDD.t4112 VDD.t4111 VDD.t4112 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1093 VDD.t4110 VDD.t4109 VDD.t4110 VDD.t2325 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1094 VDD.t4108 VDD.t4107 VDD.t4108 VDD.t20 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1095 VSS.t180 a_71496_10388.t13 a_71896_12380# VDD.t353 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1096 VSS.t3148 VSS.t3147 VSS.t3148 VSS.t1821 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1097 VDD.t98 a_31699_20742.t81 a_35502_25545.t5 VDD.t34 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1098 a_52635_34067.t59 a_35502_24538.t28 a_33249_34067.t15 VSS.t183 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1099 VDD.t4106 VDD.t4105 VDD.t4106 VDD.t288 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1100 a_102756_n36322# a_100820_n35156.t15 VDD.t526 VDD.t524 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1101 a_52635_34067.t17 a_35922_19591.t56 a_52635_48695.t64 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1102 VSS.t3146 VSS.t3145 VSS.t3146 VSS.t107 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1103 VSS.t3144 VSS.t3143 VSS.t3144 VSS.t721 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1104 VDD.t4104 VDD.t4103 VDD.t4104 VDD.t2118 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1105 VDD.t4102 VDD.t4101 VDD.t4102 VDD.t64 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1106 VDD.t4100 VDD.t4099 VDD.t4100 VDD.t2573 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1107 VSS.t425 a_36162_10388.t9 a_36562_11614# VDD.t3613 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1108 VSS.t3142 VSS.t3141 VSS.t3142 VSS.t834 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1109 a_48391_n28415# a_39179_n19595.t0 a_47819_n36322.t5 VSS.t339 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1110 a_35221_n5342# a_31953_n19727.t121 a_34347_n7136# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1111 VDD.t4098 VDD.t4097 VDD.t4098 VDD.t2570 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1112 VDD.t4096 VDD.t4095 VDD.t4096 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1113 VDD.t4094 VDD.t4093 VDD.t4094 VDD.t401 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1114 a_32913_n16904# a_31953_n19727.t122 a_32353_n16904# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1115 a_33249_35053.t11 a_33379_34917.t14 a_33249_48695.t25 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1116 a_63683_n16009# a_50751_n19729.t110 VSS.t268 VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1117 VDD.t4092 VDD.t4091 VDD.t4092 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1118 VDD.t4090 VDD.t4089 VDD.t4090 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1119 VDD.t4764 a_83153_11614.t13 a_90935_6405# VSS.t392 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1120 VSS.t3140 VSS.t3139 VSS.t3140 VSS.t808 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1121 VDD.t4088 VDD.t4087 VDD.t4088 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1122 VDD.t99 a_31699_20742.t82 a_35502_24538.t21 VDD.t25 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1123 VSS.t3138 VSS.t3137 VSS.t3138 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1124 VDD.t4086 VDD.t4085 VDD.t4086 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1125 a_95943_n20430# a_71281_n10073.t113 a_95105_n19525# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1126 VDD.t4084 VDD.t4083 VDD.t4084 VDD.t1265 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1127 a_84547_n6055# a_71281_n10073.t114 a_43010_10448.t3 VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1128 a_52635_49681.t25 a_35922_19591.t57 OUT.t82 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1129 VDD.t4082 VDD.t4081 VDD.t4082 VDD.t2288 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1130 VDD.t4080 VDD.t4079 VDD.t4080 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1131 VDD.t4078 VDD.t4077 VDD.t4078 VDD.t1708 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1132 a_51151_n8035# a_50751_n19729.t111 a_50629_n8932# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1133 a_30152_n36322.t2 a_30324_n30399.t1 a_32128_n27257# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1134 VDD.t4076 VDD.t4075 VDD.t4076 VDD.t1867 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1135 VDD.t4074 VDD.t4073 VDD.t4074 VDD.t648 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1136 VSS.t3136 VSS.t3135 VSS.t3136 VSS.t650 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1137 VDD.t100 a_31699_20742.t83 a_33249_48695.t305 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1138 VSS.t296 a_112559_4481.t13 a_113081_6405# VSS.t294 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1139 VDD.t4072 VDD.t4071 VDD.t4072 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1140 a_45706_24920# a_35922_19591.t58 a_45138_24920# VDD.t402 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X1141 VDD.t4945 a_52635_34067.t95 a_52635_48695.t158 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1142 a_83153_11614.t4 a_83153_10448.t12 a_85089_10448# VDD.t643 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1143 VDD.t4070 VDD.t4069 VDD.t4070 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1144 a_53145_n8932# a_50751_n19729.t112 a_52585_n8035# VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1145 VDD.t4068 VDD.t4067 VDD.t4068 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1146 VDD.t4066 VDD.t4065 VDD.t4066 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1147 a_31953_n19727.t59 a_31953_n19727.t58 VSS.t89 VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1148 VSS.t415 a_112559_n29181.t13 a_113081_n27257# VSS.t411 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1149 VSS.t3134 VSS.t3133 VSS.t3134 VSS.t558 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1150 a_101350_n35156# a_100820_n35156.t6 a_100820_n35156.t7 VDD.t523 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1151 VSS.t3132 VSS.t3131 VSS.t3132 VSS.t380 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1152 VSS.t3130 VSS.t3129 VSS.t3130 VSS.t1537 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1153 a_111063_n7865# a_71281_n8397.t125 a_110225_n7865# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1154 a_33249_35053.t12 a_33379_34917.t15 a_33249_48695.t26 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1155 VSS.t3128 VSS.t3127 VSS.t3128 VSS.t531 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1156 a_71496_10388.t1 a_77225_4481.t13 a_79151_6405# VSS.t318 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1157 VSS.t3126 VSS.t3125 VSS.t3126 VSS.t455 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1158 VDD.t4064 VDD.t4063 VDD.t4064 VDD.t625 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1159 a_41487_n12419# a_31953_n19727.t123 a_39179_n12419# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1160 VSS.t3124 VSS.t3123 VSS.t3124 VSS.t424 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1161 VSS.t3122 VSS.t3121 VSS.t3122 VSS.t856 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1162 VDD.t4062 VDD.t4061 VDD.t4062 VDD.t1867 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1163 a_94537_n19525# a_71281_n10073.t115 a_93969_n19525# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1164 a_89531_7563# a_83153_11614.t14 a_89009_7563.t1 VSS.t394 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1165 VDD.t4060 VDD.t4059 VDD.t4060 VDD.t2251 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1166 a_104527_n1530# a_71281_n8397.t126 a_103997_n5150# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1167 a_33249_35053.t13 a_33379_34917.t16 a_33249_48695.t27 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1168 a_111631_n2435# a_71281_n8397.t127 a_111063_n2435# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1169 a_82573_n3340# a_71281_n10073.t116 a_81735_n3340# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1170 VDD.t4058 VDD.t4057 VDD.t4058 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1171 VDD.t4056 VDD.t4055 VDD.t4056 VDD.t1112 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1172 VSS.t181 a_35502_25545.t33 a_33249_34067.t139 VSS.t27 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1173 a_71496_10388.t4 a_71366_11614.t3 a_79182_12380# VDD.t1841 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1174 VSS.t3120 VSS.t3119 VSS.t3120 VSS.t509 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1175 a_30152_n36322.t4 a_30152_n35156.t17 a_32088_n35156# VDD.t551 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1176 a_33249_34067.t138 a_35502_25545.t34 VSS.t212 VSS.t137 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1177 a_33249_48695.t304 a_31699_20742.t84 VDD.t101 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1178 a_67462_n30339# a_65658_n29313.t0 a_44363_n16007.t2 VSS.t289 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1179 VDD.t4054 VDD.t4053 VDD.t4054 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1180 VDD.t4052 VDD.t4051 VDD.t4052 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1181 a_33249_48695.t28 a_33379_34917.t17 a_33249_35053.t14 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1182 a_47753_n4445# a_31953_n19727.t124 a_47231_n6239# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1183 a_99667_n3340# a_71281_n8397.t128 a_98829_n3340# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1184 a_101350_n33224# a_100820_n35156.t4 a_100820_n35156.t5 VDD.t523 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1185 a_48313_n19595# a_31953_n19727.t125 a_47753_n18698# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1186 a_33249_34067.t87 a_33379_34007.t22 a_33249_48695.t107 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1187 VSS.t3118 VSS.t3117 VSS.t3118 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1188 VDD.t102 a_31699_20742.t85 a_35502_25545.t6 VDD.t16 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1189 VSS.t3116 VSS.t3115 VSS.t3116 VSS.t775 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1190 VSS.t3114 VSS.t3113 VSS.t3114 VSS.t842 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1191 a_52635_48695.t157 a_52635_34067.t96 VDD.t4944 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1192 VDD.t103 a_31699_20742.t86 a_33249_48695.t303 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1193 a_35502_25545.t27 a_35502_25545.t26 VSS.t211 VSS.t41 nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X1194 VDD.t4050 VDD.t4049 VDD.t4050 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1195 a_58851_n19597# a_50751_n19729.t113 VSS.t269 VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1196 VSS.t3112 VSS.t3111 VSS.t3112 VSS.t687 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1197 VDD.t4048 VDD.t4047 VDD.t4048 VDD.t2240 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1198 a_113037_n15000# a_71281_n8397.t129 a_112199_n14095# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1199 a_90245_n8770# a_71281_n10073.t117 a_89407_n8770# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1200 a_63161_n5344.t2 a_65658_4421.t1 a_66058_4481# VSS.t377 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1201 a_60845_n15112# a_50751_n19729.t114 a_60285_n14215# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1202 a_63683_n7138# a_50751_n19729.t115 a_63161_n7138# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1203 a_30152_n36322.t5 a_30152_n35156.t18 a_32088_n33224# VDD.t551 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1204 VDD.t4046 VDD.t4045 VDD.t4046 VDD.t1818 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1205 VSS.t3110 VSS.t3109 VSS.t3110 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1206 a_52635_49681.t26 a_35922_19591.t59 OUT.t81 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1207 VDD.t4044 VDD.t4043 VDD.t4044 VDD.t1218 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1208 a_36008_7563.t2 a_30152_11614.t9 a_37934_4481# VSS.t281 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1209 a_65677_n7138# a_50751_n19729.t116 a_65117_n7138# VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1210 a_44885_n12419# a_31953_n19727.t126 a_44363_n13316# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1211 a_77747_4481# a_77225_4481.t0 a_77225_4481.t1 VSS.t317 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1212 VDD.t4042 VDD.t4041 VDD.t4042 VDD.t2228 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1213 a_60285_n15112# a_50751_n19729.t117 a_59763_n16906# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1214 a_36162_n36382.t3 a_41891_n29181.t14 a_43817_n27257# VSS.t168 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1215 a_100803_n4245# a_71281_n8397.t130 a_100235_n4245# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1216 VDD.t4040 VDD.t4039 VDD.t4040 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1217 VDD.t4038 VDD.t4037 VDD.t4038 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1218 a_52635_34067.t22 a_35922_19591.t60 a_52635_48695.t63 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1219 VDD.t4036 VDD.t4035 VDD.t4036 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1220 VSS.t3108 VSS.t3107 VSS.t3108 VSS.t671 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1221 VDD.t104 a_31699_20742.t87 a_33249_48695.t302 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1222 a_71281_n10073.t63 a_71281_n10073.t62 VDD.t364 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1223 VDD.t4034 VDD.t4033 VDD.t4034 VDD.t2485 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1224 a_95943_n6055# a_71281_n10073.t118 a_78344_10448.t0 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1225 VSS.t3106 VSS.t3105 VSS.t3106 VSS.t102 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1226 VDD.t4032 VDD.t4031 VDD.t4032 VDD.t1818 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1227 VDD.t4030 VDD.t4029 VDD.t4030 VDD.t1787 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1228 VDD.t4028 VDD.t4027 VDD.t4028 VDD.t1081 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1229 VDD.t4026 VDD.t4025 VDD.t4026 VDD.t60 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1230 a_84547_n18620# a_71281_n10073.t119 a_83709_n18620# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1231 VDD.t4024 VDD.t4023 VDD.t4024 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1232 VDD.t4022 VDD.t4021 VDD.t4022 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1233 a_40613_n2651# a_31953_n19727.t127 a_40053_n2651# VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1234 VSS.t3104 VSS.t3103 VSS.t3104 VSS.t399 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1235 VDD.t4020 VDD.t4019 VDD.t4020 VDD.t2485 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1236 a_54579_n15112# a_50751_n19729.t118 a_54019_n14215# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1237 VDD.t4018 VDD.t4017 VDD.t4018 VDD.t297 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1238 VSS.t3102 VSS.t3101 VSS.t3102 VSS.t353 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1239 VSS.t3100 VSS.t3099 VSS.t3100 VSS.t196 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1240 VDD.t4016 VDD.t4015 VDD.t4016 VDD.t1653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1241 a_64243_n14215# a_50751_n19729.t119 a_63683_n14215# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1242 a_79151_n30339# a_77225_n29181.t12 VSS.t383 VSS.t381 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1243 VDD.t4014 VDD.t4013 VDD.t4014 VDD.t406 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1244 VSS.t202 a_35502_25545.t35 a_33249_34067.t137 VSS.t21 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1245 a_33249_48695.t301 a_31699_20742.t88 VDD.t105 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1246 a_32128_4481# a_30324_5507.t1 a_31284_4481.t1 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1247 a_52635_49681.t162 a_52635_34067.t97 VDD.t4943 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1248 a_32353_n8930# a_31953_n19727.t128 a_31831_n8930# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1249 VDD.t4012 VDD.t4011 VDD.t4012 VDD.t60 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1250 VDD.t4010 VDD.t4009 VDD.t4010 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1251 VDD.t4008 VDD.t4007 VDD.t4008 VDD.t1787 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1252 VSS.t3098 VSS.t3097 VSS.t3098 VSS.t740 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1253 VDD.t4006 VDD.t4005 VDD.t4006 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1254 a_34347_n8930# a_31953_n19727.t129 a_33787_n8930# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1255 VDD.t4004 VDD.t4003 VDD.t4004 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1256 VDD.t4002 VDD.t4001 VDD.t4002 VDD.t2485 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1257 a_45706_24195# a_35922_19591.t61 a_45138_24195# VDD.t402 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X1258 a_33249_35053.t15 a_33379_34917.t18 a_33249_48695.t29 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1259 a_77747_n28415# a_77225_n29181.t13 a_71496_n36382.t2 VSS.t379 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1260 VDD.t4000 VDD.t3999 VDD.t4000 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1261 a_40053_n1754# a_31953_n19727.t130 VSS.t109 VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1262 a_35502_24538.t20 a_31699_20742.t89 VDD.t106 VDD.t14 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1263 a_83725_n30339# a_32913_n8930.t1 a_83153_n36322.t3 VSS.t287 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1264 VDD.t3998 VDD.t3997 VDD.t3998 VDD.t404 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1265 a_54229_10448# a_53829_10388.t10 a_36032_13546.t0 VDD.t3678 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1266 a_33249_34067.t86 a_33379_34007.t23 a_33249_48695.t108 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1267 VDD.t3996 VDD.t3995 VDD.t3996 VDD.t549 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1268 VDD.t40 a_31699_20742.t35 a_31699_20742.t36 VDD.t34 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1269 a_52635_49681.t161 a_52635_34067.t98 VDD.t4942 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1270 a_33249_34067.t14 a_35502_24538.t29 a_52635_34067.t56 VSS.t185 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1271 VDD.t3994 VDD.t3993 VDD.t3994 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1272 a_46319_n13316# a_31953_n19727.t131 a_45797_n14213# VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1273 VSS.t3096 VSS.t3095 VSS.t3096 VSS.t1253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1274 VSS.t3094 VSS.t3093 VSS.t3094 VSS.t1426 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1275 VDD.t3992 VDD.t3991 VDD.t3992 VDD.t1049 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1276 a_33249_48695.t300 a_31699_20742.t90 VDD.t107 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1277 VDD.t3990 VDD.t3989 VDD.t3990 VDD.t47 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1278 VSS.t3092 VSS.t3091 VSS.t3092 VSS.t108 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1279 a_57977_n14215# a_50751_n19729.t120 a_57417_n14215# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1280 VSS.t3090 VSS.t3089 VSS.t3090 VSS.t859 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1281 VSS.t3088 VSS.t3087 VSS.t3088 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1282 VDD.t3988 VDD.t3987 VDD.t3988 VDD.t1180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1283 VSS.t3086 VSS.t3085 VSS.t3086 VSS.t2036 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X1284 VDD.t108 a_31699_20742.t91 a_33249_48695.t299 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1285 a_52635_49681.t27 a_35922_19591.t62 OUT.t80 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1286 a_52635_34067.t22 a_35922_19591.t63 a_52635_48695.t62 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1287 a_41487_n1754# a_31953_n19727.t132 a_39179_n1754# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1288 VDD.t3986 VDD.t3985 VDD.t3986 VDD.t925 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1289 VDD.t3984 VDD.t3983 VDD.t3984 VDD.t555 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1290 VSS.t3084 VSS.t3083 VSS.t3084 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1291 VSS.t3082 VSS.t3081 VSS.t3082 VSS.t795 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1292 a_89715_n17715.t3 a_100992_4421.t1 a_113110_12380# VDD.t336 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1293 VSS.t3080 VSS.t3079 VSS.t3080 VSS.t229 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1294 VDD.t3982 VDD.t3981 VDD.t3982 VDD.t1419 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1295 a_57977_n6241# a_50751_n19729.t121 a_57417_n4447# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1296 VDD.t3980 VDD.t3979 VDD.t3980 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1297 VSS.t3078 VSS.t3077 VSS.t3078 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1298 VSS.t3076 VSS.t3075 VSS.t3076 VSS.t1615 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1299 a_71281_n10073.t61 a_71281_n10073.t60 VDD.t361 VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1300 VDD.t3978 VDD.t3977 VDD.t3978 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1301 a_51151_n3550# a_50751_n19729.t122 a_50629_n4447# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1302 VSS.t3074 VSS.t3073 VSS.t3074 VSS.t877 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1303 VDD.t3976 VDD.t3975 VDD.t3976 VDD.t1365 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1304 a_35502_25545.t7 a_31699_20742.t92 VDD.t109 VDD.t32 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1305 VSS.t3072 VSS.t3071 VSS.t3072 VSS.t591 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1306 VDD.t3974 VDD.t3973 VDD.t3974 VDD.t1155 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1307 VSS.t3070 VSS.t3069 VSS.t3070 VSS.t944 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1308 VDD.t459 a_71281_n8397.t54 a_71281_n8397.t55 VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1309 a_53145_n3550# a_50751_n19729.t123 a_52585_n3550# VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1310 VDD.t3972 VDD.t3971 VDD.t3972 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1311 a_52635_34067.t23 a_35922_19591.t64 a_52635_48695.t61 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1312 VDD.t3970 VDD.t3969 VDD.t3970 VDD.t120 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1313 VSS.t3068 VSS.t3067 VSS.t3068 VSS.t153 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1314 VSS.t3066 VSS.t3065 VSS.t3066 VSS.t591 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1315 VSS.t3064 VSS.t3063 VSS.t3064 VSS.t721 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1316 VDD.t3968 VDD.t3967 VDD.t3968 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1317 VSS.t3062 VSS.t3061 VSS.t3062 VSS.t596 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1318 VDD.t3966 VDD.t3965 VDD.t3966 VDD.t910 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1319 a_110225_n9675# a_71281_n8397.t131 a_109695_n9675# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1320 a_52635_34067.t24 a_35922_19591.t65 a_52635_48695.t60 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1321 VDD.t3964 VDD.t3963 VDD.t3964 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1322 a_33249_48695.t2 a_33379_34007.t24 a_33249_34067.t85 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1323 VSS.t3060 VSS.t3059 VSS.t3060 VSS.t588 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1324 VDD.t3962 VDD.t3961 VDD.t3962 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1325 VSS.t3058 VSS.t3057 VSS.t3058 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1326 VSS.t3056 VSS.t3055 VSS.t3056 VSS.t3 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1327 VSS.t3054 VSS.t3053 VSS.t3054 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1328 a_37968_13546# a_36162_10388.t10 a_36008_4481.t2 VDD.t1711 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1329 a_47991_4421.t0 a_47819_11614.t12 a_54197_4481# VSS.t304 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1330 VDD.t4941 a_52635_34067.t99 a_52635_49681.t160 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1331 VSS.t3052 VSS.t3051 VSS.t3052 VSS.t1222 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1332 VSS.t3050 VSS.t3049 VSS.t3050 VSS.t1466 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1333 a_33249_34067.t84 a_33379_34007.t25 a_33249_48695.t3 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1334 a_33249_35053.t16 a_33379_34917.t19 a_33249_48695.t30 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1335 a_85129_n29181# a_32913_n8930.t2 a_31831_n5342.t1 VSS.t286 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1336 VDD.t3960 VDD.t3959 VDD.t3960 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1337 VDD.t3958 VDD.t3957 VDD.t3958 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1338 VDD.t3956 VDD.t3955 VDD.t3956 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1339 a_93969_n1530# a_71281_n10073.t120 a_93131_n1530# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1340 VSS.t3048 VSS.t3047 VSS.t3048 VSS.t495 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1341 a_99667_n13190# a_71281_n8397.t132 a_98829_n13190# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1342 a_33249_34067.t83 a_33379_34007.t26 a_33249_48695.t4 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1343 VDD.t3954 VDD.t3953 VDD.t3954 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1344 VDD.t3952 VDD.t3951 VDD.t3952 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1345 VSS.t345 a_89163_10388.t12 a_89563_12380# VDD.t554 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1346 VSS.t3046 VSS.t3045 VSS.t3046 VSS.t1385 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1347 a_114485_5639# a_112559_4481.t14 VSS.t298 VSS.t297 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1348 a_47753_n19595# a_31953_n19727.t133 VSS.t110 VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1349 VSS.t3044 VSS.t3043 VSS.t3044 VSS.t615 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1350 a_111063_n13190# a_71281_n8397.t133 a_110225_n13190# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1351 a_71896_10448# a_71496_10388.t14 a_53699_13546.t3 VDD.t351 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1352 VDD.t3950 VDD.t3949 VDD.t3950 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1353 VDD.t3948 VDD.t3947 VDD.t3948 VDD.t917 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1354 a_113037_n6055# a_71281_n8397.t134 VDD.t476 VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1355 VSS.t3042 VSS.t3041 VSS.t3042 VSS.t760 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1356 VDD.t3946 VDD.t3945 VDD.t3946 VDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1357 VDD.t3944 VDD.t3943 VDD.t3944 VDD.t1570 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1358 VDD.t3942 VDD.t3941 VDD.t3942 VDD.t965 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1359 a_37968_11614# a_36162_10388.t11 VSS.t426 VDD.t1711 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1360 VSS.t3040 VSS.t3039 VSS.t3040 VSS.t757 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1361 VSS.t3038 VSS.t3037 VSS.t3038 VSS.t681 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1362 a_82573_n2435# a_71281_n10073.t121 a_81735_n2435# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1363 VSS.t3036 VSS.t3035 VSS.t3036 VSS.t1594 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1364 a_54019_n12421# a_50751_n19729.t124 VSS.t270 VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1365 VDD.t3940 VDD.t3939 VDD.t3940 VDD.t1957 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1366 VSS.t3034 VSS.t3033 VSS.t3034 VSS.t684 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1367 a_52635_34067.t25 a_35922_19591.t66 a_52635_48695.t59 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1368 a_52635_48695.t58 a_35922_19591.t67 a_52635_34067.t26 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1369 VDD.t3938 VDD.t3937 VDD.t3938 VDD.t287 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1370 a_89531_n29181# a_83153_n36322.t10 VDD.t4780 VSS.t454 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1371 VDD.t3936 VDD.t3935 VDD.t3936 VDD.t1333 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1372 a_106501_n14095# a_71281_n8397.t135 a_105933_n14095# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1373 VDD.t3934 VDD.t3933 VDD.t3934 VDD.t2 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1374 VSS.t88 a_31953_n19727.t56 a_31953_n19727.t57 VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1375 a_99667_n2435# a_71281_n8397.t136 a_98829_n2435# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1376 VSS.t3032 VSS.t3031 VSS.t3032 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1377 VDD.t3932 VDD.t3931 VDD.t3932 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1378 a_33249_35053.t17 a_33379_34917.t20 a_33249_48695.t31 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1379 a_65117_n7138# a_50751_n19729.t125 a_64595_n8035# VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1380 VDD.t3930 VDD.t3929 VDD.t3930 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1381 VDD.t3928 VDD.t3927 VDD.t3928 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1382 a_101641_n6055# a_71281_n8397.t137 a_101111_n6055.t0 VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1383 VDD.t3926 VDD.t3925 VDD.t3926 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1384 VSS.t3030 VSS.t3029 VSS.t3030 VSS.t68 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1385 VSS.t3028 VSS.t3027 VSS.t3028 VSS.t671 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1386 VSS.t3026 VSS.t3025 VSS.t3026 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1387 VDD.t3924 VDD.t3923 VDD.t3924 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1388 a_52635_49681.t159 a_52635_34067.t100 VDD.t4940 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1389 VDD.t3922 VDD.t3921 VDD.t3922 VDD.t1936 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1390 a_38097_n16007.t1 a_47991_n29313.t0 a_48391_n29181# VSS.t340 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1391 VSS.t3024 VSS.t3023 VSS.t3024 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1392 a_90245_n8770# a_71281_n10073.t122 a_89407_n7865# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1393 VDD.t3920 VDD.t3919 VDD.t3920 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1394 VDD.t3918 VDD.t3917 VDD.t3918 VDD.t398 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1395 VDD.t3916 VDD.t3915 VDD.t3916 VDD.t1540 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1396 VDD.t3914 VDD.t3913 VDD.t3914 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1397 VDD.t110 a_31699_20742.t93 a_33249_48695.t298 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1398 VSS.t3022 VSS.t3021 VSS.t3022 VSS.t609 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1399 VDD.t3912 VDD.t3911 VDD.t3912 VDD.t1209 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1400 VDD.t4939 a_52635_34067.t101 a_52635_48695.t156 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1401 a_112559_n29181.t10 a_112559_n29181.t9 a_114485_n28415# VSS.t409 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1402 a_33379_34007.t27 IN_POS.t1 cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
X1403 VDD.t3910 VDD.t3909 VDD.t3910 VDD.t2777 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1404 VSS.t3020 VSS.t3019 VSS.t3020 VSS.t534 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1405 VDD.t3908 VDD.t3907 VDD.t3908 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1406 VDD.t3906 VDD.t3905 VDD.t3906 VDD.t664 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1407 a_67111_n8932# a_50751_n19729.t126 a_66551_n8035# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1408 a_67462_5639# a_65658_4421.t0 a_63161_n5344.t1 VSS.t289 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1409 VDD.t3904 VDD.t3903 VDD.t3904 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1410 a_63683_n15112# a_50751_n19729.t127 a_63161_n15112# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1411 VSS.t3018 VSS.t3017 VSS.t3018 VSS.t305 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1412 VSS.t3016 VSS.t3015 VSS.t3016 VSS.t1431 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1413 VDD.t3902 VDD.t3901 VDD.t3902 VDD.t2349 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1414 a_33249_35053.t18 a_33379_34917.t21 a_33249_48695.t32 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1415 a_33249_34067.t13 a_35502_24538.t30 a_52635_34067.t57 VSS.t184 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1416 VDD.t3900 VDD.t3899 VDD.t3900 VDD.t398 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1417 VSS.t3014 VSS.t3013 VSS.t3014 VSS.t644 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1418 a_88839_n4245# a_71281_n10073.t123 a_88271_n4245# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1419 VDD.t4766 a_30152_n36322.t10 a_37934_n28415# VSS.t281 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1420 VDD.t3898 VDD.t3897 VDD.t3898 VDD.t2088 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1421 a_79182_10448# a_71366_11614.t4 a_78344_10448.t3 VDD.t571 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1422 VDD.t3896 VDD.t3895 VDD.t3896 VDD.t955 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1423 VDD.t3894 VDD.t3893 VDD.t3894 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1424 VDD.t3892 VDD.t3891 VDD.t3892 VDD.t1299 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1425 a_45445_n18698# a_31953_n19727.t134 a_44885_n18698# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1426 VDD.t3890 VDD.t3889 VDD.t3890 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1427 a_33249_35053.t19 a_33379_34917.t22 a_33249_48695.t33 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1428 VSS.t3012 VSS.t3011 VSS.t3012 VSS.t817 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1429 VSS.t3010 VSS.t3009 VSS.t3010 VSS.t891 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1430 a_35781_n15110# a_31953_n19727.t135 a_35221_n15110# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1431 a_94892_4481.t1 a_94892_4481.t0 a_96818_5639# VSS.t396 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1432 a_84547_n17715# a_71281_n10073.t124 a_84017_n17715.t0 VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1433 VSS.t3008 VSS.t3007 VSS.t3008 VSS.t2475 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X1434 VSS.t3006 VSS.t3005 VSS.t3006 VSS.t638 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1435 VSS.t290 a_53829_n36382.t15 a_54229_n35156# VDD.t301 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1436 VDD.t3888 VDD.t3887 VDD.t3888 VDD.t3747 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1437 a_33249_48695.t297 a_31699_20742.t94 VDD.t111 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1438 VSS.t3004 VSS.t3003 VSS.t3004 VSS.t478 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1439 VSS.t3002 VSS.t3001 VSS.t3002 VSS.t733 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1440 OUT.t17 a_35502_24538.t31 a_33249_35053.t89 VSS.t183 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1441 a_66551_n18700# a_50751_n19729.t128 a_66029_n18700# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1442 VSS.t3000 VSS.t2999 VSS.t3000 VSS.t484 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1443 VSS.t2998 VSS.t2997 VSS.t2998 VSS.t1244 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1444 a_52635_34067.t25 a_35922_19591.t68 a_52635_48695.t57 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1445 VDD.t3886 VDD.t3885 VDD.t3886 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1446 a_46879_n14213# a_31953_n19727.t136 a_46319_n14213# VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1447 VDD.t3884 VDD.t3883 VDD.t3884 VDD.t1936 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1448 a_89033_n36322.t1 a_106830_n36382.t9 a_108636_n36322# VDD.t1290 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1449 VDD.t3882 VDD.t3881 VDD.t3882 VDD.t965 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1450 VDD.t3880 VDD.t3879 VDD.t3880 VDD.t2349 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1451 VSS.t2996 VSS.t2995 VSS.t2996 VSS.t60 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1452 a_32353_n19595# a_31953_n19727.t137 a_31831_n19595# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1453 VDD.t39 a_31699_20742.t33 a_31699_20742.t34 VDD.t38 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1454 VDD.t4938 a_52635_34067.t102 a_52635_49681.t158 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1455 VDD.t3878 VDD.t3877 VDD.t3878 VDD.t1505 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1456 VDD.t3876 VDD.t3875 VDD.t3876 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1457 VSS.t2994 VSS.t2993 VSS.t2994 VSS.t1064 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1458 a_95414_n27257# a_94892_n29181.t9 a_94892_n29181.t10 VSS.t353 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1459 VDD.t3874 VDD.t3873 VDD.t3874 VDD.t920 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X1460 VSS.t2992 VSS.t2991 VSS.t2992 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1461 VDD.t3872 VDD.t3871 VDD.t3872 VDD.t1086 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1462 a_38619_n4445# a_31953_n19727.t138 a_38097_n4445# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1463 a_53675_n27257.t1 a_53829_n36382.t16 a_54229_n33224# VDD.t301 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1464 VSS.t2990 VSS.t2989 VSS.t2990 VSS.t338 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1465 a_33249_34067.t136 a_35502_25545.t36 VSS.t201 VSS.t31 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1466 VDD.t3870 VDD.t3869 VDD.t3870 VDD.t962 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1467 VDD.t3868 VDD.t3867 VDD.t3868 VDD.t667 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1468 VDD.t324 a_100820_10448.t12 a_101350_12380# VDD.t293 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1469 VSS.t2988 VSS.t2987 VSS.t2988 VSS.t509 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1470 VDD.t458 a_71281_n8397.t52 a_71281_n8397.t53 VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1471 a_33249_34067.t135 a_35502_25545.t37 VSS.t177 VSS.t137 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1472 a_112559_4481.t5 a_112559_4481.t4 a_114485_7563# VSS.t292 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1473 a_50629_n16009.t1 a_51711_n12421.t0 a_83725_5639# VSS.t311 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1474 VSS.t197 a_41891_4481.t14 a_42413_7563# VSS.t166 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1475 VDD.t3866 VDD.t3865 VDD.t3866 VDD.t1489 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1476 VDD.t3864 VDD.t3863 VDD.t3864 VDD.t1164 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1477 VDD.t3862 VDD.t3861 VDD.t3862 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1478 VDD.t3860 VDD.t3859 VDD.t3860 VDD.t2058 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1479 VSS.t2986 VSS.t2985 VSS.t2986 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1480 a_52635_34067.t27 a_35922_19591.t69 a_52635_48695.t56 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1481 VSS.t2984 VSS.t2983 VSS.t2984 VSS.t1253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1482 VDD.t3858 VDD.t3857 VDD.t3858 VDD.t1486 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1483 a_31699_20742.t32 a_31699_20742.t31 VDD.t37 VDD.t32 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1484 a_71281_n8397.t72 I1N.t6 a_75585_n10973# VSS.t312 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X1485 a_33249_35053.t20 a_33379_34917.t23 a_33249_48695.t34 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1486 VDD.t3856 VDD.t3855 VDD.t3856 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1487 a_63683_n6241# a_50751_n19729.t129 a_63161_n7138# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1488 a_33249_48695.t296 a_31699_20742.t95 VDD.t112 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1489 VDD.t3854 VDD.t3853 VDD.t3854 VDD.t1265 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1490 a_52635_48695.t155 a_52635_34067.t103 VDD.t4937 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1491 VSS.t2982 VSS.t2981 VSS.t2982 VSS.t157 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1492 a_33249_48695.t295 a_31699_20742.t96 VDD.t113 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1493 VSS.t2980 VSS.t2979 VSS.t2980 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1494 VSS.t2978 VSS.t2977 VSS.t2978 VSS.t1306 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1495 a_96818_5639# a_94892_4481.t11 VSS.t3637 VSS.t1303 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1496 VSS.t2976 VSS.t2975 VSS.t2976 VSS.t576 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1497 a_33249_35053.t21 a_33379_34917.t24 a_33249_48695.t35 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1498 VDD.t3852 VDD.t3851 VDD.t3852 VDD.t1481 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1499 VDD.t3850 VDD.t3849 VDD.t3850 VDD.t502 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1500 a_50751_n19729.t55 a_50751_n19729.t54 VSS.t246 VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1501 a_53675_n27257.t2 a_47819_n36322.t10 a_55601_n30339# VSS.t307 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1502 a_113110_13546# a_86903_n14095.t4 a_106830_10388.t4 VDD.t337 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1503 a_33249_34067.t134 a_35502_25545.t38 VSS.t200 VSS.t16 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1504 a_83141_n4245# a_71281_n10073.t125 a_82573_n4245# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1505 VSS.t2974 VSS.t2973 VSS.t2974 VSS.t690 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1506 a_52635_49681.t157 a_52635_34067.t104 VDD.t4936 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1507 VDD.t3848 VDD.t3847 VDD.t3848 VDD.t309 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1508 VDD.t3846 VDD.t3845 VDD.t3846 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1509 VDD.t3844 VDD.t3843 VDD.t3844 VDD.t789 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1510 VDD.t3842 VDD.t3841 VDD.t3842 VDD.t635 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1511 VSS.t2972 VSS.t2971 VSS.t2972 VSS.t1294 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1512 a_48349_13546# a_47819_10448.t12 a_47819_11614.t0 VDD.t507 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1513 VDD.t377 a_71281_n10073.t126 a_83709_n21335# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1514 VDD.t3840 VDD.t3839 VDD.t3840 VDD.t2021 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1515 a_100235_n4245# a_71281_n8397.t138 a_99667_n4245# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1516 VDD.t3838 VDD.t3837 VDD.t3838 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1517 a_56895_n16009.t1 a_57977_n12421.t0 a_101392_7563# VSS.t162 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1518 VSS.t2970 VSS.t2969 VSS.t2970 VSS.t676 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1519 VSS.t2968 VSS.t2967 VSS.t2968 VSS.t150 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1520 VSS.t2966 VSS.t2965 VSS.t2966 VSS.t1287 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1521 VSS.t2964 VSS.t2963 VSS.t2964 VSS.t490 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1522 a_39179_n19595.t0 a_47819_n36322.t11 a_54197_n28415# VSS.t304 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1523 VSS.t2962 VSS.t2961 VSS.t2962 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1524 a_59411_n7138# a_50751_n19729.t130 a_60285_n5344# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1525 VSS.t2960 VSS.t2959 VSS.t2960 VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1526 a_107339_n6960# a_71281_n8397.t139 a_106501_n6960# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1527 a_33249_35053.t22 a_33379_34917.t25 a_33249_48695.t36 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1528 VDD.t3836 VDD.t3835 VDD.t3836 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1529 VDD.t3834 VDD.t3833 VDD.t3834 VDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1530 VSS.t2958 VSS.t2957 VSS.t2958 VSS.t763 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1531 a_65677_n13318# a_50751_n19729.t131 a_65117_n13318# VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1532 a_113110_11614# a_86903_n14095.t5 a_106830_10388.t5 VDD.t337 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1533 VDD.t3832 VDD.t3831 VDD.t3832 VDD.t1042 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1534 a_101641_n20430# a_71281_n8397.t140 a_100803_n19525# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1535 a_48313_n8930# a_31953_n19727.t139 a_47753_n8930# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1536 a_113081_7563# a_112559_4481.t15 a_106830_10388.t0 VSS.t293 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1537 a_51151_n18700# a_50751_n19729.t132 a_50629_n19597# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1538 a_51711_n8035# a_50751_n19729.t133 a_51151_n7138# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1539 VDD.t3830 VDD.t3829 VDD.t3830 VDD.t2680 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1540 VDD.t3828 VDD.t3827 VDD.t3828 VDD.t536 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1541 VDD.t3826 VDD.t3825 VDD.t3826 VDD.t610 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1542 a_65486_10448.t8 a_65658_4421.t0 a_67462_7563# VSS.t378 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1543 VDD.t3824 VDD.t3823 VDD.t3824 VDD.t2231 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1544 VSS.t2956 VSS.t2955 VSS.t2956 VSS.t591 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1545 VSS.t2954 VSS.t2953 VSS.t2954 VSS.t668 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1546 VDD.t3822 VDD.t3821 VDD.t3822 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1547 a_53829_n36382.t4 a_53699_n35156.t5 a_61515_n35156# VDD.t546 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1548 a_86903_n14095.t0 a_106830_10388.t12 a_108636_12380# VDD.t521 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1549 a_48349_11614# a_47819_10448.t13 a_47819_11614.t1 VDD.t507 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1550 VDD.t3820 VDD.t3819 VDD.t3820 VDD.t1611 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1551 a_67422_n34390# a_65486_n35156.t17 VDD.t7 VDD.t6 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1552 a_83725_5639# a_51711_n12421.t0 a_83153_11614.t3 VSS.t310 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1553 a_42413_7563# a_41891_4481.t15 a_36162_10388.t3 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1554 a_51711_n16009.t1 a_50751_n19729.t134 a_51151_n16009# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1555 VSS.t2952 VSS.t2951 VSS.t2952 VSS.t588 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1556 VDD.t3818 VDD.t3817 VDD.t3818 VDD.t1996 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1557 VDD.t3816 VDD.t3815 VDD.t3816 VDD.t427 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1558 VSS.t2950 VSS.t2949 VSS.t2950 VSS.t398 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1559 a_52635_49681.t28 a_35922_19591.t70 OUT.t79 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1560 VDD.t114 a_31699_20742.t97 a_33249_48695.t294 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1561 a_79151_7563# a_77225_4481.t14 VSS.t321 VSS.t319 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1562 a_33249_34067.t133 a_35502_25545.t39 VSS.t22 VSS.t21 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1563 VSS.t44 a_35502_25545.t40 a_33249_35053.t138 VSS.t25 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1564 a_60285_n4447# a_50751_n19729.t135 a_59763_n6241# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1565 a_33249_48695.t293 a_31699_20742.t98 VDD.t116 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1566 a_113037_n6960# a_71281_n8397.t141 a_112199_n4245# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1567 VSS.t2948 VSS.t2947 VSS.t2948 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1568 a_35221_n13316# a_31953_n19727.t140 a_34699_n14213# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1569 VDD.t4935 a_52635_34067.t105 a_52635_49681.t156 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1570 VDD.t3814 VDD.t3813 VDD.t3814 VDD.t905 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1571 VDD.t3812 VDD.t3811 VDD.t3812 VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1572 VDD.t3810 VDD.t3809 VDD.t3810 VDD.t2231 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1573 VDD.t3808 VDD.t3807 VDD.t3808 VDD.t60 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1574 VDD.t3806 VDD.t3805 VDD.t3806 VDD.t1218 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1575 VDD.t3804 VDD.t3803 VDD.t3804 VDD.t893 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1576 VDD.t3802 VDD.t3801 VDD.t3802 VDD.t390 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1577 a_53829_n36382.t5 a_53699_n35156.t6 a_61515_n33224# VDD.t546 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1578 VDD.t3800 VDD.t3799 VDD.t3800 VDD.t1611 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1579 VSS.t2946 VSS.t2945 VSS.t2946 VSS.t395 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1580 VDD.t3798 VDD.t3797 VDD.t3798 VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1581 VSS.t2944 VSS.t2943 VSS.t2944 VSS.t528 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1582 a_60677_n36322.t1 a_47991_n29313.t1 a_60109_n35156# VDD.t545 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1583 VSS.t2942 VSS.t2941 VSS.t2942 VSS.t453 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1584 VSS.t24 a_35502_25545.t41 a_33249_35053.t137 VSS.t18 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1585 a_107339_n20430# a_71281_n8397.t142 a_106501_n19525# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1586 a_110225_n13190# a_71281_n8397.t143 a_109695_n16810# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1587 a_33249_48695.t37 a_33379_34917.t26 a_33249_35053.t23 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1588 a_67111_n4447# a_50751_n19729.t136 a_66551_n3550# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1589 VSS.t2940 VSS.t2939 VSS.t2940 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1590 VDD.t3796 VDD.t3795 VDD.t3796 VDD.t1799 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1591 VSS.t2938 VSS.t2937 VSS.t2938 VSS.t868 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1592 VDD.t374 a_71281_n10073.t58 a_71281_n10073.t59 VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1593 VSS.t2936 VSS.t2935 VSS.t2936 VSS.t553 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1594 VDD.t3794 VDD.t3793 VDD.t3794 VDD.t1424 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1595 a_111063_n1530# a_71281_n8397.t144 a_110225_n1530# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1596 VSS.t2934 VSS.t2933 VSS.t2934 VSS.t550 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1597 VSS.t2932 VSS.t2931 VSS.t2932 VSS.t376 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1598 VSS.t2930 VSS.t2929 VSS.t2930 VSS.t814 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1599 VDD.t3792 VDD.t3791 VDD.t3792 VDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1600 VDD.t4934 a_52635_34067.t106 a_52635_49681.t155 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1601 VDD.t3790 VDD.t3789 VDD.t3790 VDD.t875 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1602 OUT.t16 a_35502_24538.t32 a_33249_35053.t90 VSS.t184 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1603 VDD.t3788 VDD.t3787 VDD.t3788 VDD.t401 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1604 a_82573_n15000# a_71281_n10073.t127 a_81735_n15000# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1605 a_60677_n36322.t1 a_47991_n29313.t1 a_60109_n33224# VDD.t545 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1606 a_51151_n2653# a_50751_n19729.t137 a_50629_n2653# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1607 VSS.t2928 VSS.t2927 VSS.t2928 VSS.t339 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1608 VDD.t3786 VDD.t3785 VDD.t3786 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1609 VSS.t2926 VSS.t2925 VSS.t2926 VSS.t12 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1610 VSS.t2924 VSS.t2923 VSS.t2924 VSS.t183 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1611 VDD.t4933 a_52635_34067.t107 a_52635_48695.t154 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1612 a_33249_35053.t91 a_35502_24538.t33 OUT.t15 VSS.t185 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1613 VDD.t3784 VDD.t3783 VDD.t3784 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1614 a_52635_49681.t154 a_52635_34067.t108 VDD.t4932 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1615 VSS.t2922 VSS.t2921 VSS.t2922 VSS.t795 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1616 a_53145_n2653# a_50751_n19729.t138 a_52585_n2653# VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1617 a_52635_49681.t153 a_52635_34067.t109 VDD.t4931 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1618 VDD.t3782 VDD.t3781 VDD.t3782 VDD.t1408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1619 VSS.t2920 VSS.t2919 VSS.t2920 VSS.t618 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1620 VDD.t3780 VDD.t3779 VDD.t3780 VDD.t925 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1621 VSS.t2918 VSS.t2917 VSS.t2918 VSS.t1594 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1622 a_52635_49681.t152 a_52635_34067.t110 VDD.t4930 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1623 VSS.t445 a_59558_n29181.t14 a_60080_n29181# VSS.t401 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1624 VDD.t3778 VDD.t3777 VDD.t3778 VDD.t852 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1625 VSS.t2916 VSS.t2915 VSS.t2916 VSS.t534 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1626 VDD.t4776 a_65486_11614.t9 a_73268_5639# VSS.t422 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1627 VSS.t2914 VSS.t2913 VSS.t2914 VSS.t733 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1628 VDD.t3776 VDD.t3775 VDD.t3776 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1629 VSS.t2912 VSS.t2911 VSS.t2912 VSS.t615 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1630 VDD.t3774 VDD.t3773 VDD.t3774 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1631 VDD.t3772 VDD.t3771 VDD.t3772 VDD.t550 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1632 VSS.t2910 VSS.t2909 VSS.t2910 VSS.t650 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1633 VDD.t3770 VDD.t3769 VDD.t3770 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1634 a_32913_n12419# a_31953_n19727.t141 a_32353_n12419# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1635 VDD.t3768 VDD.t3767 VDD.t3768 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1636 a_46274_23609# a_35922_19591.t71 a_45706_23609# VDD.t407 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X1637 VSS.t2908 VSS.t2907 VSS.t2908 VSS.t1315 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1638 VDD.t3766 VDD.t3765 VDD.t3766 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1639 VSS.t2906 VSS.t2905 VSS.t2906 VSS.t1615 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1640 VSS.t291 a_35502_25545.t42 a_33249_34067.t132 VSS.t27 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1641 VSS.t187 a_35502_24538.t34 a_41100_19075# VSS.t186 nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X1642 VSS.t2904 VSS.t2903 VSS.t2904 VSS.t604 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1643 VSS.t2902 VSS.t2901 VSS.t2902 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1644 VDD.t3764 VDD.t3763 VDD.t3764 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1645 a_33249_48695.t292 a_31699_20742.t99 VDD.t117 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1646 VDD.t3762 VDD.t3761 VDD.t3762 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1647 VDD.t3760 VDD.t3759 VDD.t3760 VDD.t697 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1648 VDD.t3758 VDD.t3757 VDD.t3758 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1649 VDD.t3756 VDD.t3755 VDD.t3756 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1650 VSS.t2900 VSS.t2899 VSS.t2900 VSS.t1537 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1651 VSS.t2898 VSS.t2897 VSS.t2898 VSS.t478 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1652 VDD.t3754 VDD.t3753 VDD.t3754 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1653 VDD.t3752 VDD.t3751 VDD.t3752 VDD.t910 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1654 VDD.t3750 VDD.t3749 VDD.t3750 VDD.t3570 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1655 VDD.t3748 VDD.t3746 VDD.t3748 VDD.t3747 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1656 a_33249_48695.t291 a_31699_20742.t100 VDD.t118 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1657 a_67111_n17803# a_50751_n19729.t139 a_66551_n17803# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1658 a_52635_49681.t151 a_52635_34067.t111 VDD.t4929 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1659 a_105365_n9675# a_71281_n8397.t145 a_104527_n9675# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1660 a_63683_n1756# a_50751_n19729.t140 a_63161_n2653# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1661 VSS.t2896 VSS.t2895 VSS.t2896 VSS.t772 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1662 VDD.t119 a_31699_20742.t101 a_33249_48695.t290 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1663 VDD.t3745 VDD.t3744 VDD.t3745 VDD.t979 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1664 a_105933_n4245# a_71281_n8397.t146 a_105365_n4245# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1665 VSS.t245 a_50751_n19729.t52 a_50751_n19729.t53 VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1666 a_82573_n20430# a_71281_n10073.t128 a_81735_n20430# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1667 a_53675_4481.t3 a_47819_11614.t13 a_55601_7563# VSS.t307 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1668 VDD.t3743 VDD.t3742 VDD.t3743 VDD.t697 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1669 VDD.t3741 VDD.t3740 VDD.t3741 VDD.t1155 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1670 VDD.t3739 VDD.t3738 VDD.t3739 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1671 a_65677_n2653# a_50751_n19729.t141 a_65117_n1756# VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1672 VSS.t2894 VSS.t2893 VSS.t2894 VSS.t704 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1673 VSS.t2892 VSS.t2891 VSS.t2892 VSS.t1034 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1674 a_71864_5639# a_65486_11614.t10 VDD.t4777 VSS.t423 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1675 VDD.t3737 VDD.t3736 VDD.t3737 VDD.t801 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1676 a_43817_n30339# a_41891_n29181.t15 VSS.t370 VSS.t158 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1677 a_42442_13546# a_36032_11614.t7 a_36162_10388.t6 VDD.t288 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1678 VDD.t3735 VDD.t3734 VDD.t3735 VDD.t1515 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1679 VDD.t3733 VDD.t3732 VDD.t3733 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1680 VSS.t2890 VSS.t2889 VSS.t2890 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1681 VDD.t3731 VDD.t3730 VDD.t3731 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1682 a_53829_10388.t0 a_53699_11614.t3 a_61515_12380# VDD.t1512 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1683 VDD.t3729 VDD.t3728 VDD.t3729 VDD.t2118 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1684 VDD.t3727 VDD.t3726 VDD.t3727 VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1685 a_38619_n17801# a_31953_n19727.t142 a_38097_n17801# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1686 VSS.t2888 VSS.t2887 VSS.t2888 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1687 a_100235_n18620# a_71281_n8397.t147 a_99667_n18620# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1688 VSS.t2886 VSS.t2885 VSS.t2886 VSS.t568 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1689 VDD.t3725 VDD.t3724 VDD.t3725 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1690 VSS.t2884 VSS.t2883 VSS.t2884 VSS.t908 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1691 a_49795_n30339# a_47991_n29313.t0 a_38097_n16007.t2 VSS.t338 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1692 VDD.t3723 VDD.t3722 VDD.t3723 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1693 VSS.t2882 VSS.t2881 VSS.t2882 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1694 VSS.t2880 VSS.t2879 VSS.t2880 VSS.t377 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1695 a_31953_n19727.t55 a_31953_n19727.t54 VSS.t87 VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1696 a_52635_48695.t55 a_35922_19591.t72 a_52635_34067.t28 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1697 a_52635_34067.t62 a_35502_24538.t35 a_33249_34067.t12 VSS.t196 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1698 VDD.t3721 VDD.t3720 VDD.t3721 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1699 a_33249_34067.t82 a_33379_34007.t28 a_33249_48695.t111 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1700 a_96818_n28415# a_94892_n29181.t12 VSS.t355 VSS.t354 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1701 a_111631_n13190# a_71281_n8397.t148 a_111063_n13190# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1702 a_65658_n29313.t0 a_65486_n36322.t12 a_71864_n27257# VSS.t157 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1703 a_33249_48695.t289 a_31699_20742.t102 VDD.t121 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1704 a_42442_11614# a_36032_11614.t8 a_36162_10388.t7 VDD.t288 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1705 VDD.t3719 VDD.t3718 VDD.t3719 VDD.t1515 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1706 VSS.t2878 VSS.t2877 VSS.t2878 VSS.t1157 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1707 VDD.t3717 VDD.t3716 VDD.t3717 VDD.t2118 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1708 VDD.t3715 VDD.t3714 VDD.t3715 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1709 VDD.t3713 VDD.t3712 VDD.t3713 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1710 a_36032_11614.t1 a_36162_10388.t12 a_37968_12380# VDD.t1494 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1711 VDD.t3711 VDD.t3710 VDD.t3711 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1712 a_33249_48695.t288 a_31699_20742.t103 VDD.t123 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1713 a_102756_n35156# a_100820_n35156.t16 VDD.t527 VDD.t524 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1714 VSS.t2876 VSS.t2875 VSS.t2876 VSS.t568 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1715 VSS.t2874 VSS.t2873 VSS.t2874 VSS.t410 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1716 a_36162_10388.t2 a_41891_4481.t16 a_43817_4481# VSS.t168 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1717 a_35781_n15110# a_31953_n19727.t143 a_35221_n14213# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1718 VDD.t3709 VDD.t3708 VDD.t3709 VDD.t2573 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1719 a_36008_4481.t3 a_36162_10388.t13 a_36562_10448# VDD.t3613 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1720 VDD.t3707 VDD.t3706 VDD.t3707 VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1721 VDD.t3705 VDD.t3704 VDD.t3705 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1722 VSS.t2872 VSS.t2871 VSS.t2872 VSS.t108 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1723 a_98829_n18620# a_71281_n8397.t149 a_98299_n19525# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1724 a_30152_11614.t0 a_30324_5507.t1 a_32128_6405# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1725 VDD.t3703 VDD.t3702 VDD.t3703 VDD.t2570 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1726 VDD.t3701 VDD.t3700 VDD.t3701 VDD.t398 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1727 VDD.t3699 VDD.t3698 VDD.t3699 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1728 VSS.t2870 VSS.t2869 VSS.t2870 VSS.t464 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1729 VSS.t2868 VSS.t2867 VSS.t2868 VSS.t306 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1730 a_33249_34067.t131 a_35502_25545.t43 VSS.t208 VSS.t145 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1731 a_33787_n18698# a_31953_n19727.t144 a_33265_n18698# VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1732 a_30724_n27257# a_30324_n29313.t1 a_30152_n35156.t3 VSS.t150 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1733 VSS.t2866 VSS.t2865 VSS.t2866 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1734 VDD.t3697 VDD.t3696 VDD.t3697 VDD.t352 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1735 VDD.t3695 VDD.t3694 VDD.t3695 VDD.t1867 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1736 VSS.t2864 VSS.t2863 VSS.t2864 VSS.t650 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1737 VDD.t3693 VDD.t3692 VDD.t3693 VDD.t337 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1738 a_105365_n18620# a_71281_n8397.t150 a_104527_n18620# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1739 a_55601_7563# a_47819_11614.t14 a_47991_4421.t0 VSS.t305 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1740 VSS.t2862 VSS.t2861 VSS.t2862 VSS.t56 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1741 a_102756_n33224# a_100820_n35156.t17 VDD.t528 VDD.t524 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1742 VSS.t2860 VSS.t2859 VSS.t2860 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1743 VSS.t2858 VSS.t2857 VSS.t2858 VSS.t60 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1744 VDD.t3691 VDD.t3690 VDD.t3691 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1745 VDD.t3689 VDD.t3688 VDD.t3689 VDD.t404 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1746 a_33249_35053.t136 a_35502_25545.t44 VSS.t206 VSS.t29 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1747 VDD.t3687 VDD.t3686 VDD.t3687 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1748 a_33249_48695.t287 a_31699_20742.t104 VDD.t124 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1749 VSS.t2856 VSS.t2855 VSS.t2856 VSS.t641 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1750 VDD.t3685 VDD.t3684 VDD.t3685 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1751 a_52635_48695.t54 a_35922_19591.t73 a_52635_34067.t29 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1752 VDD.t3683 VDD.t3682 VDD.t3683 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1753 VDD.t3681 VDD.t3680 VDD.t3681 VDD.t523 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1754 VSS.t2854 VSS.t2853 VSS.t2854 VSS.t1256 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1755 VDD.t36 a_31699_20742.t29 a_31699_20742.t30 VDD.t14 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1756 VSS.t2852 VSS.t2851 VSS.t2852 VSS.t379 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1757 VDD.t3679 VDD.t3677 VDD.t3679 VDD.t3678 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1758 VDD.t3676 VDD.t3675 VDD.t3676 VDD.t2921 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1759 a_110225_n3340# a_71281_n8397.t151 a_109695_n4245# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1760 a_100820_11614.t5 a_57977_n12421.t0 a_102796_4481# VSS.t171 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1761 a_33249_48695.t112 a_33379_34007.t29 a_33249_34067.t81 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1762 a_31284_4481.t1 a_30324_4421.t2 a_30724_4481# VSS.t151 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1763 VDD.t331 a_71281_n10073.t56 a_71281_n10073.t57 VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1764 a_58851_n8035# a_50751_n19729.t142 a_58329_n8035# VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1765 a_52635_49681.t150 a_52635_34067.t112 VDD.t4928 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1766 VSS.t2850 VSS.t2849 VSS.t2850 VSS.t337 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1767 VSS.t2848 VSS.t2847 VSS.t2848 VSS.t384 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1768 VDD.t125 a_31699_20742.t105 a_33249_48695.t286 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1769 a_52635_49681.t149 a_52635_34067.t113 VDD.t4927 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1770 VDD.t3674 VDD.t3673 VDD.t3674 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1771 VDD.t3672 VDD.t3671 VDD.t3672 VDD.t551 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1772 VDD.t3670 VDD.t3669 VDD.t3670 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1773 VDD.t3668 VDD.t3667 VDD.t3668 VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1774 VDD.t3666 VDD.t3665 VDD.t3666 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1775 a_57417_n16906# a_50751_n19729.t143 a_56895_n17803# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1776 VSS.t2846 VSS.t2845 VSS.t2846 VSS.t37 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1777 VSS.t2844 VSS.t2843 VSS.t2844 VSS.t185 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1778 VDD.t3664 VDD.t3663 VDD.t3664 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1779 VDD.t3662 VDD.t3661 VDD.t3662 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1780 a_102796_6405# a_57977_n12421.t2 a_56895_n16009.t1 VSS.t172 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1781 VDD.t3660 VDD.t3659 VDD.t3660 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1782 VDD.t3658 VDD.t3657 VDD.t3658 VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1783 VDD.t126 a_31699_20742.t106 a_33249_48695.t285 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1784 VDD.t3656 VDD.t3655 VDD.t3656 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1785 a_82573_n15905# a_71281_n10073.t129 a_81735_n15905# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1786 a_43817_4481# a_41891_4481.t17 VSS.t189 VSS.t158 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1787 a_33249_35053.t24 a_33379_34917.t27 a_33249_48695.t38 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1788 VSS.t2842 VSS.t2841 VSS.t2842 VSS.t976 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1789 a_66058_n30339# a_45445_n19595.t1 a_65486_n36322.t5 VSS.t376 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1790 a_48313_n15110# a_31953_n19727.t145 a_47753_n15110# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1791 a_112199_n6960# a_71281_n8397.t152 a_111631_n6960# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1792 a_83325_n29313.t0 a_83153_n36322.t11 a_89531_n27257# VSS.t453 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1793 VDD.t3654 VDD.t3653 VDD.t3654 VDD.t553 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1794 VDD.t3652 VDD.t3651 VDD.t3652 VDD.t120 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1795 VSS.t244 a_50751_n19729.t50 a_50751_n19729.t51 VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1796 a_89563_n34390# a_89163_n36382.t10 a_89033_n35156.t2 VDD.t548 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1797 a_52635_49681.t29 a_35922_19591.t74 OUT.t78 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1798 VDD.t3650 VDD.t3649 VDD.t3650 VDD.t1818 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1799 VDD.t3648 VDD.t3647 VDD.t3648 VDD.t522 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1800 VSS.t2840 VSS.t2839 VSS.t2840 VSS.t501 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1801 VDD.t3646 VDD.t3645 VDD.t3646 VDD.t49 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1802 VSS.t2838 VSS.t2837 VSS.t2838 VSS.t947 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1803 VSS.t2836 VSS.t2835 VSS.t2836 VSS.t1615 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1804 VDD.t3644 VDD.t3643 VDD.t3644 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1805 VDD.t3642 VDD.t3641 VDD.t3642 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1806 VDD.t127 a_31699_20742.t107 a_33249_48695.t284 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1807 VSS.t2834 VSS.t2833 VSS.t2834 VSS.t262 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1808 VSS.t2832 VSS.t2831 VSS.t2832 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1809 VDD.t3640 VDD.t3639 VDD.t3640 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1810 VSS.t2830 VSS.t2829 VSS.t2830 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1811 VDD.t3638 VDD.t3637 VDD.t3638 VDD.t1086 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1812 a_41100_19075# a_35502_24538.t36 a_40578_19075# VSS.t191 nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X1813 VDD.t3636 VDD.t3635 VDD.t3636 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1814 VSS.t2828 VSS.t2827 VSS.t2828 VSS.t490 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1815 a_35502_24538.t19 a_31699_20742.t108 VDD.t128 VDD.t18 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1816 a_48391_n27257# a_47991_n29313.t2 a_47819_n35156.t11 VSS.t339 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1817 a_101392_4481# a_100992_4421.t2 a_100820_10448.t0 VSS.t163 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1818 VDD.t3634 VDD.t3633 VDD.t3634 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1819 a_65677_n13318# a_50751_n19729.t144 a_65117_n12421# VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1820 VSS.t2826 VSS.t2825 VSS.t2826 VSS.t1466 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1821 VDD.t3632 VDD.t3631 VDD.t3632 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1822 a_51711_n6241# a_50751_n19729.t145 a_51151_n6241# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1823 a_89715_n5150.t1 a_71281_n10073.t130 a_89407_n1530# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1824 VSS.t2824 VSS.t2823 VSS.t2824 VSS.t1126 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1825 VSS.t2822 VSS.t2821 VSS.t2822 VSS.t339 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1826 a_65486_n36322.t6 a_45445_n19595.t1 a_67462_n29181# VSS.t378 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1827 VSS.t2820 VSS.t2819 VSS.t2820 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1828 a_30724_4481# a_30324_4421.t2 a_30152_10448.t1 VSS.t150 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1829 VDD.t3630 VDD.t3629 VDD.t3630 VDD.t1787 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1830 VDD.t3628 VDD.t3627 VDD.t3628 VDD.t499 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1831 a_51711_n16906# a_50751_n19729.t146 a_51151_n15112# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1832 a_107198_5639# a_100820_11614.t8 VDD.t422 VSS.t182 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1833 VSS.t2818 VSS.t2817 VSS.t2818 VSS.t650 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1834 a_33249_48695.t39 a_33379_34917.t28 a_33249_35053.t25 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1835 VDD.t3626 VDD.t3625 VDD.t3626 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1836 VSS.t2816 VSS.t2815 VSS.t2816 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1837 a_65117_n1756# a_50751_n19729.t147 a_64243_n5344.t0 VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1838 VSS.t2814 VSS.t2813 VSS.t2814 VSS.t1111 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1839 a_33249_34067.t80 a_33379_34007.t30 a_33249_48695.t113 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1840 VSS.t2812 VSS.t2811 VSS.t2812 VSS.t259 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1841 VSS.t2810 VSS.t2809 VSS.t2810 VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1842 VDD.t4926 a_52635_34067.t114 a_52635_49681.t148 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1843 VSS.t2808 VSS.t2807 VSS.t2808 VSS.t263 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1844 VDD.t3624 VDD.t3623 VDD.t3624 VDD.t1180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1845 a_33249_35053.t26 a_33379_34917.t29 a_33249_48695.t40 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1846 VSS.t2806 VSS.t2805 VSS.t2806 VSS.t1537 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1847 a_52635_48695.t153 a_52635_34067.t115 VDD.t4925 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1848 VDD.t3622 VDD.t3621 VDD.t3622 VDD.t78 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1849 a_90969_13546# a_89163_10388.t13 a_89009_4481.t2 VDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1850 a_33249_48695.t283 a_31699_20742.t109 VDD.t129 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1851 VSS.t2804 VSS.t2803 VSS.t2804 VSS.t459 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1852 VDD.t3620 VDD.t3619 VDD.t3620 VDD.t2485 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1853 VSS.t243 a_50751_n19729.t48 a_50751_n19729.t49 VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1854 VSS.t448 a_106830_n36382.t10 a_107230_n34390# VDD.t845 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1855 VSS.t2802 VSS.t2801 VSS.t2802 VSS.t498 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1856 a_89407_n8770# a_71281_n10073.t131 a_88839_n8770# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1857 VSS.t2800 VSS.t2799 VSS.t2800 VSS.t937 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1858 a_67111_n2653# a_50751_n19729.t148 a_66551_n2653# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1859 VDD.t3618 VDD.t3617 VDD.t3618 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1860 VDD.t3616 VDD.t3615 VDD.t3616 VDD.t836 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1861 VDD.t3614 VDD.t3612 VDD.t3614 VDD.t3613 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1862 VDD.t3611 VDD.t3610 VDD.t3611 VDD.t1251 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1863 a_32353_n8033# a_31953_n19727.t146 a_31831_n8930# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1864 a_53145_n7138# a_50751_n19729.t149 a_54019_n5344# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1865 a_40053_n8930# a_31953_n19727.t147 a_39179_n5342.t0 VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1866 VDD.t3609 VDD.t3608 VDD.t3609 VDD.t1180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1867 a_71281_n8397.t51 a_71281_n8397.t50 VDD.t457 VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1868 a_54019_n18700# a_50751_n19729.t150 a_53497_n18700# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1869 a_40053_n12419# a_31953_n19727.t148 VSS.t111 VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1870 VSS.t2798 VSS.t2797 VSS.t2798 VSS.t647 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1871 VDD.t3607 VDD.t3606 VDD.t3607 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1872 a_90969_11614# a_89163_10388.t14 VSS.t346 VDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1873 VDD.t3605 VDD.t3604 VDD.t3605 VDD.t1042 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1874 VDD.t3603 VDD.t3602 VDD.t3603 VDD.t2299 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X1875 a_34347_n8930# a_31953_n19727.t149 a_33787_n8033# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1876 VSS.t2796 VSS.t2795 VSS.t2796 VSS.t409 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1877 VSS.t2794 VSS.t2793 VSS.t2794 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1878 VSS.t2792 VSS.t2791 VSS.t2792 VSS.t336 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1879 VDD.t511 a_47819_10448.t14 a_48349_12380# VDD.t510 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1880 VSS.t2790 VSS.t2789 VSS.t2790 VSS.t349 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1881 VDD.t3601 VDD.t3600 VDD.t3601 VDD.t823 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1882 VSS.t2788 VSS.t2787 VSS.t2788 VSS.t265 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1883 VSS.t2786 VSS.t2785 VSS.t2786 VSS.t531 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1884 VDD.t3599 VDD.t3598 VDD.t3599 VDD.t427 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1885 a_67422_n36322# a_65486_n35156.t18 VDD.t8 VDD.t6 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1886 VDD.t3597 VDD.t3596 VDD.t3597 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1887 a_41487_n8930# a_31953_n19727.t150 VSS.t112 VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1888 a_33249_48695.t282 a_31699_20742.t110 VDD.t130 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1889 VSS.t2784 VSS.t2783 VSS.t2784 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1890 VSS.t2782 VSS.t2781 VSS.t2782 VSS.t1431 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1891 VSS.t2780 VSS.t2779 VSS.t2780 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1892 VDD.t3595 VDD.t3594 VDD.t3595 VDD.t810 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1893 VSS.t2778 VSS.t2777 VSS.t2778 VSS.t281 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1894 VSS.t2776 VSS.t2775 VSS.t2776 VSS.t571 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1895 VDD.t3593 VDD.t3592 VDD.t3593 VDD.t3354 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1896 a_33249_48695.t41 a_33379_34917.t30 a_33249_35053.t27 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1897 VDD.t4924 a_52635_34067.t116 a_52635_49681.t147 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1898 VSS.t2774 VSS.t2773 VSS.t2774 VSS.t633 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1899 VDD.t4923 a_52635_34067.t117 a_52635_48695.t152 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1900 a_61484_n30339# a_59558_n29181.t15 VSS.t446 VSS.t399 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1901 a_83325_4421.t0 a_83153_11614.t15 a_89531_4481# VSS.t393 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1902 VSS.t2772 VSS.t2771 VSS.t2772 VSS.t868 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1903 a_98829_n17715# a_71281_n8397.t153 a_98299_n21335# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1904 VSS.t2770 VSS.t2769 VSS.t2770 VSS.t842 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1905 a_100820_n35156.t3 a_100992_n29313.t0 a_102796_n30339# VSS.t329 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1906 VSS.t2768 VSS.t2767 VSS.t2768 VSS.t733 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1907 VSS.t2766 VSS.t2765 VSS.t2766 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1908 VDD.t3591 VDD.t3590 VDD.t3591 VDD.t338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1909 a_85129_6405# a_51711_n12421.t2 a_50629_n16009.t1 VSS.t309 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1910 VDD.t3589 VDD.t3588 VDD.t3589 VDD.t55 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1911 VDD.t3587 VDD.t3586 VDD.t3587 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1912 VDD.t3585 VDD.t3584 VDD.t3585 VDD.t917 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1913 a_52635_49681.t30 a_35922_19591.t75 OUT.t77 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1914 VSS.t2764 VSS.t2763 VSS.t2764 VSS.t282 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1915 VSS.t2762 VSS.t2761 VSS.t2762 VSS.t1157 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1916 VDD.t131 a_31699_20742.t111 a_35502_25545.t8 VDD.t38 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1917 VDD.t3583 VDD.t3582 VDD.t3583 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1918 VSS.t2760 VSS.t2759 VSS.t2760 VSS.t558 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1919 VDD.t456 a_71281_n8397.t48 a_71281_n8397.t49 VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1920 VDD.t3581 VDD.t3580 VDD.t3581 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1921 a_58851_n3550# a_50751_n19729.t151 a_58329_n3550# VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1922 VSS.t2758 VSS.t2757 VSS.t2758 VSS.t487 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1923 VDD.t3579 VDD.t3578 VDD.t3579 VDD.t1957 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1924 a_95443_n34390# a_89033_n35156.t9 a_89163_n36382.t6 VDD.t795 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1925 VDD.t3577 VDD.t3576 VDD.t3577 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1926 a_95443_12380# a_83325_4421.t1 a_94892_4481.t8 VDD.t497 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1927 VSS.t2756 VSS.t2755 VSS.t2756 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1928 VSS.t2754 VSS.t2753 VSS.t2754 VSS.t537 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1929 a_44885_n7136# a_31953_n19727.t151 a_44363_n7136# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1930 VSS.t2752 VSS.t2751 VSS.t2752 VSS.t699 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1931 VSS.t2750 VSS.t2749 VSS.t2750 VSS.t33 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1932 a_34347_n17801# a_31953_n19727.t152 a_33787_n17801# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1933 VDD.t340 a_71281_n10073.t54 a_71281_n10073.t55 VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1934 VDD.t3575 VDD.t3574 VDD.t3575 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1935 VDD.t3573 VDD.t3572 VDD.t3573 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1936 a_52635_49681.t31 a_35922_19591.t76 OUT.t76 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1937 a_52635_49681.t32 a_35922_19591.t77 OUT.t75 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1938 a_90245_n17715# a_71281_n10073.t132 a_89715_n16810.t0 VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1939 a_46879_n7136# a_31953_n19727.t153 a_46319_n7136# VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1940 VDD.t3571 VDD.t3569 VDD.t3571 VDD.t3570 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1941 VSS.t2748 VSS.t2747 VSS.t2748 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1942 VDD.t3568 VDD.t3567 VDD.t3568 VDD.t1841 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1943 VDD.t295 a_65486_n36322.t13 a_73268_n28415# VSS.t155 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1944 VDD.t3566 VDD.t3565 VDD.t3566 VDD.t917 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1945 a_95105_n15000# a_71281_n10073.t133 a_94537_n15000# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1946 a_47753_n16007# a_31953_n19727.t154 a_46879_n17801# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1947 a_110225_n2435# a_71281_n8397.t154 VDD.t477 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1948 a_88271_n4245# a_71281_n10073.t134 a_87433_n4245# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1949 VSS.t2746 VSS.t2745 VSS.t2746 VSS.t612 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1950 a_90245_n15000# a_71281_n10073.t135 a_89407_n15000# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1951 VDD.t3564 VDD.t3563 VDD.t3564 VDD.t1936 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1952 VDD.t3562 VDD.t3561 VDD.t3562 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1953 VDD.t3560 VDD.t3559 VDD.t3560 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1954 a_37968_10448# a_36162_10388.t14 a_36008_7563.t0 VDD.t1711 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1955 VDD.t3558 VDD.t3557 VDD.t3558 VDD.t1195 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1956 VDD.t3556 VDD.t3555 VDD.t3556 VDD.t1957 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1957 VSS.t2744 VSS.t2743 VSS.t2744 VSS.t99 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1958 a_77747_n27257# a_77225_n29181.t3 a_77225_n29181.t4 VSS.t379 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1959 a_100235_n21335# a_71281_n8397.t155 a_99667_n21335# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1960 VSS.t2742 VSS.t2741 VSS.t2742 VSS.t837 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1961 VDD.t3554 VDD.t3553 VDD.t3554 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1962 VDD.t3552 VDD.t3551 VDD.t3552 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1963 VSS.t2740 VSS.t2739 VSS.t2740 VSS.t282 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1964 a_42047_n7136# a_31953_n19727.t155 a_41487_n6239# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1965 VDD.t4748 a_65486_10448.t14 a_66016_12380# VDD.t1338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1966 VSS.t2738 VSS.t2737 VSS.t2738 VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1967 VSS.t2736 VSS.t2735 VSS.t2736 VSS.t558 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1968 VDD.t132 a_31699_20742.t112 a_33249_48695.t281 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1969 VDD.t3550 VDD.t3549 VDD.t3550 VDD.t3423 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1970 VDD.t3548 VDD.t3547 VDD.t3548 VDD.t1333 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1971 a_112559_n29181.t2 a_100992_n29313.t2 a_114516_n34390# VDD.t538 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1972 a_60677_10448.t1 a_53699_11614.t4 a_60109_13546# VDD.t664 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1973 a_32128_n28415# a_30324_n29313.t0 a_31284_n30339.t2 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1974 VSS.t2734 VSS.t2733 VSS.t2734 VSS.t39 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1975 VSS.t2732 VSS.t2731 VSS.t2732 VSS.t192 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1976 a_107198_n30339# a_100820_n36322.t11 a_106676_n30339.t1 VSS.t335 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1977 a_52635_49681.t146 a_52635_34067.t118 VDD.t4922 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1978 VSS.t2730 VSS.t2729 VSS.t2730 VSS.t522 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1979 a_89531_4481# a_83153_11614.t16 a_89009_4481.t0 VSS.t394 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1980 a_71281_n10073.t53 a_71281_n10073.t52 VDD.t368 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1981 VDD.t3546 VDD.t3545 VDD.t3546 VDD.t1936 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1982 VDD.t3544 VDD.t3543 VDD.t3544 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1983 VDD.t3542 VDD.t3541 VDD.t3542 VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1984 a_88839_n15000# a_71281_n10073.t136 a_88271_n15000# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1985 VDD.t3540 VDD.t3539 VDD.t3540 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1986 a_30324_5507.t0 a_50751_n19729.t152 a_51151_n1756# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1987 a_33249_34067.t79 a_33379_34007.t31 a_33249_48695.t102 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1988 a_98829_n21335# a_71281_n8397.t156 a_98299_n21335# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1989 VDD.t3538 VDD.t3537 VDD.t3538 VDD.t1333 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1990 VDD.t3536 VDD.t3535 VDD.t3536 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1991 VSS.t3638 a_94892_4481.t12 a_95414_5639# VSS.t1037 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1992 a_60677_10448.t2 a_53699_11614.t5 a_60109_11614# VDD.t664 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1993 VSS.t2728 VSS.t2727 VSS.t2728 VSS.t304 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1994 a_60845_n19597# a_50751_n19729.t153 a_60285_n19597# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1995 a_101350_12380# a_100820_10448.t3 a_100820_10448.t4 VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1996 a_33249_34067.t78 a_33379_34007.t32 a_33249_48695.t103 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1997 VSS.t2726 VSS.t2725 VSS.t2726 VSS.t357 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1998 VDD.t3534 VDD.t3533 VDD.t3534 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1999 a_36530_n28415# a_30152_n36322.t11 VDD.t4767 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2000 a_106809_n5150.t1 a_103997_n8770.t5 a_113110_n34390# VDD.t537 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2001 a_33249_48695.t280 a_31699_20742.t113 VDD.t133 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2002 VSS.t207 a_35502_25545.t45 a_33249_35053.t135 VSS.t25 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2003 VDD.t3532 VDD.t3531 VDD.t3532 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2004 a_105365_n21335# a_71281_n8397.t157 a_104527_n21335# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2005 VDD.t540 a_100820_n36322.t12 a_108602_n29181# VSS.t333 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2006 VSS.t2724 VSS.t2723 VSS.t2724 VSS.t108 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2007 VSS.t2722 VSS.t2721 VSS.t2722 VSS.t576 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2008 a_33249_34067.t130 a_35502_25545.t46 VSS.t178 VSS.t145 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2009 VDD.t3530 VDD.t3529 VDD.t3530 VDD.t979 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2010 a_45445_n16904# a_31953_n19727.t156 a_44885_n15110# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2011 VDD.t3528 VDD.t3527 VDD.t3528 VDD.t1299 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2012 VSS.t2720 VSS.t2719 VSS.t2720 VSS.t1025 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2013 VDD.t3526 VDD.t3525 VDD.t3526 VDD.t301 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2014 a_95105_n20430# a_71281_n10073.t137 a_94537_n20430# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2015 a_50751_n19729.t47 a_50751_n19729.t46 VSS.t242 VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2016 OUT.t14 a_35502_24538.t37 a_33249_35053.t96 VSS.t196 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2017 a_89009_4481.t1 a_83153_11614.t17 a_90935_7563# VSS.t392 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2018 VSS.t2718 VSS.t2717 VSS.t2718 VSS.t1466 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2019 VDD.t3524 VDD.t3523 VDD.t3524 VDD.t500 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2020 a_90245_n20430# a_71281_n10073.t138 a_89407_n20430# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2021 VDD.t3522 VDD.t3521 VDD.t3522 VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2022 a_83709_n6960# a_71281_n10073.t139 a_83141_n6960# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2023 VSS.t2716 VSS.t2715 VSS.t2716 VSS.t808 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2024 a_39179_n6239# a_31953_n19727.t157 a_38619_n4445# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2025 VDD.t3520 VDD.t3519 VDD.t3520 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2026 VDD.t3518 VDD.t3517 VDD.t3518 VDD.t720 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2027 VDD.t3516 VDD.t3515 VDD.t3516 VDD.t1164 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2028 VDD.t3514 VDD.t3513 VDD.t3514 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2029 a_103997_n8770.t2 a_106830_n36382.t11 a_108636_n35156# VDD.t1290 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2030 a_54579_n19597# a_50751_n19729.t154 a_54019_n19597# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2031 VDD.t3512 VDD.t3511 VDD.t3512 VDD.t2349 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2032 a_32353_n16007# a_31953_n19727.t158 a_31284_n30339.t0 VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2033 VSS.t19 a_35502_25545.t47 a_33249_35053.t134 VSS.t18 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2034 a_33249_48695.t104 a_33379_34007.t33 a_33249_34067.t77 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2035 VSS.t2714 VSS.t2713 VSS.t2714 VSS.t856 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2036 VSS.t299 a_112559_4481.t16 a_113081_7563# VSS.t294 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2037 VDD.t3510 VDD.t3509 VDD.t3510 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2038 a_54019_n5344# a_50751_n19729.t155 a_53145_n3550# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2039 a_64243_n19597# a_50751_n19729.t156 a_63683_n19597# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2040 a_49755_n34390# a_47819_n35156.t16 VDD.t4794 VDD.t707 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2041 a_107339_n6055# a_71281_n8397.t158 a_106809_n6055.t1 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2042 a_32353_n3548# a_31953_n19727.t159 a_31831_n4445# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2043 VDD.t3508 VDD.t3507 VDD.t3508 VDD.t1299 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2044 a_73268_6405# a_65486_11614.t11 a_64243_n1756.t1 VSS.t421 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2045 VSS.t2712 VSS.t2711 VSS.t2712 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2046 a_34347_n3548# a_31953_n19727.t160 a_33787_n3548# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2047 a_77225_4481.t5 a_77225_4481.t4 a_79151_7563# VSS.t318 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2048 I1U.t1 I1U.t0 VSS.t350 VSS.t349 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X2049 a_88839_n20430# a_71281_n10073.t140 a_88271_n20430# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2050 VDD.t3506 VDD.t3505 VDD.t3506 VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2051 a_89407_n7865# a_71281_n10073.t141 a_88839_n7865# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2052 a_33249_48695.t279 a_31699_20742.t114 VDD.t135 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2053 VDD.t3504 VDD.t3503 VDD.t3504 VDD.t1164 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2054 a_95414_5639# a_94892_4481.t13 a_89163_10388.t0 VSS.t998 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2055 VSS.t2710 VSS.t2709 VSS.t2710 VSS.t868 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2056 VCM.t1 a_106830_n36382.t12 a_108636_n33224# VDD.t1290 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2057 VDD.t3502 VDD.t3501 VDD.t3502 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2058 VSS.t2708 VSS.t2707 VSS.t2708 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2059 a_48313_n15110# a_31953_n19727.t161 a_47753_n14213# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2060 a_52635_48695.t53 a_35922_19591.t78 a_52635_34067.t30 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2061 VDD.t3500 VDD.t3499 VDD.t3500 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2062 VDD.t3498 VDD.t3497 VDD.t3498 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2063 a_52635_48695.t151 a_52635_34067.t119 VDD.t4921 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2064 a_46319_n18698# a_31953_n19727.t162 a_45797_n18698# VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2065 a_105933_n18620# a_71281_n8397.t159 a_105365_n18620# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2066 a_105365_n3340# a_71281_n8397.t160 a_104527_n3340# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2067 VSS.t2706 VSS.t2705 VSS.t2706 VSS.t1244 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X2068 VSS.t241 a_50751_n19729.t44 a_50751_n19729.t45 VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2069 a_35922_19591.t5 a_35502_25545.t48 VSS.t42 VSS.t41 nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X2070 VSS.t2704 VSS.t2703 VSS.t2704 VSS.t588 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2071 a_57977_n19597# a_50751_n19729.t157 a_57417_n19597# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2072 VDD.t3496 VDD.t3495 VDD.t3496 VDD.t1265 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2073 VDD.t3494 VDD.t3493 VDD.t3494 VDD.t14 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2074 VSS.t2702 VSS.t2701 VSS.t2702 VSS.t775 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2075 VSS.t2700 VSS.t2699 VSS.t2700 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2076 VDD.t3492 VDD.t3491 VDD.t3492 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2077 VDD.t3490 VDD.t3489 VDD.t3490 VDD.t322 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2078 VDD.t3488 VDD.t3487 VDD.t3488 VDD.t930 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2079 a_106830_n36382.t7 a_112559_n29181.t14 a_114485_n27257# VSS.t409 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2080 VSS.t2698 VSS.t2697 VSS.t2698 VSS.t266 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2081 VSS.t2696 VSS.t2695 VSS.t2696 VSS.t1064 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2082 VDD.t3486 VDD.t3485 VDD.t3486 VDD.t1127 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2083 VSS.t2694 VSS.t2693 VSS.t2694 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2084 VSS.t2692 VSS.t2691 VSS.t2692 VSS.t671 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2085 VSS.t2690 VSS.t2689 VSS.t2690 VSS.t528 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2086 VDD.t3484 VDD.t3483 VDD.t3484 VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2087 VSS.t2688 VSS.t2687 VSS.t2688 VSS.t262 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2088 VSS.t2686 VSS.t2685 VSS.t2686 VSS.t377 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2089 VSS.t2684 VSS.t2683 VSS.t2684 VSS.t215 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2090 VSS.t2682 VSS.t2681 VSS.t2682 VSS.t795 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2091 VDD.t3482 VDD.t3481 VDD.t3482 VDD.t406 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2092 VSS.t2680 VSS.t2679 VSS.t2680 VSS.t1431 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2093 VSS.t2678 VSS.t2677 VSS.t2678 VSS.t281 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2094 VDD.t3480 VDD.t3479 VDD.t3480 VDD.t64 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2095 VDD.t3478 VDD.t3477 VDD.t3478 VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2096 a_36008_n30339.t0 a_30152_n36322.t12 a_37934_n27257# VSS.t281 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2097 a_106501_n8770# a_71281_n8397.t161 a_105933_n8770# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2098 VSS.t2676 VSS.t2675 VSS.t2676 VSS.t1315 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2099 a_104527_n18620# a_71281_n8397.t162 a_103997_n19525# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2100 VSS.t2674 VSS.t2673 VSS.t2674 VSS.t317 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2101 VDD.t3476 VDD.t3475 VDD.t3476 VDD.t1265 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2102 a_46319_n7136# a_31953_n19727.t163 a_45797_n8033# VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2103 VSS.t2672 VSS.t2671 VSS.t2672 VSS.t401 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2104 VDD.t3474 VDD.t3473 VDD.t3474 VDD.t568 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X2105 VDD.t3472 VDD.t3471 VDD.t3472 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2106 a_82573_n14095# a_71281_n10073.t142 a_81735_n14095# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2107 a_52635_48695.t52 a_35922_19591.t79 a_52635_34067.t31 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2108 VDD.t136 a_31699_20742.t115 a_33249_48695.t278 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2109 VDD.t138 a_31699_20742.t116 a_33249_48695.t277 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2110 VSS.t2670 VSS.t2669 VSS.t2670 VSS.t308 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2111 a_114516_12380# a_86903_n14095.t6 a_89715_n17715.t4 VDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2112 a_95105_n6960# a_71281_n10073.t143 a_94537_n6960# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2113 VSS.t2668 VSS.t2667 VSS.t2668 VSS.t908 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2114 a_52635_49681.t145 a_52635_34067.t120 VDD.t4920 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2115 a_113110_10448# a_100992_4421.t1 a_112559_4481.t9 VDD.t337 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2116 VSS.t2666 VSS.t2665 VSS.t2666 VSS.t733 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2117 VSS.t371 a_41891_n29181.t16 a_42413_n29181# VSS.t166 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2118 VDD.t3470 VDD.t3469 VDD.t3470 VDD.t546 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2119 VSS.t2664 VSS.t2663 VSS.t2664 VSS.t591 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2120 a_33249_48695.t276 a_31699_20742.t117 VDD.t139 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2121 VDD.t3468 VDD.t3467 VDD.t3468 VDD.t1611 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2122 a_66551_n5344# a_50751_n19729.t158 a_65677_n3550# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2123 VDD.t4919 a_52635_34067.t121 a_52635_48695.t150 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2124 VSS.t2662 VSS.t2661 VSS.t2662 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2125 a_35502_24538.t18 a_31699_20742.t118 VDD.t140 VDD.t18 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2126 VSS.t2660 VSS.t2659 VSS.t2660 VSS.t262 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2127 a_48349_10448# a_47819_10448.t4 a_47819_10448.t5 VDD.t507 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2128 a_95105_n15905# a_71281_n10073.t144 a_94537_n15905# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2129 VSS.t2658 VSS.t2657 VSS.t2658 VSS.t834 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2130 a_90245_n18620# a_71281_n10073.t145 a_89407_n15905# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2131 VSS.t2656 VSS.t2655 VSS.t2656 VSS.t259 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2132 VDD.t4918 a_52635_34067.t122 a_52635_49681.t144 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2133 VDD.t3466 VDD.t3465 VDD.t3466 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2134 VDD.t3464 VDD.t3463 VDD.t3464 VDD.t1439 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2135 VSS.t2654 VSS.t2653 VSS.t2654 VSS.t263 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2136 a_48313_n8930# a_31953_n19727.t164 a_47753_n8033# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2137 VDD.t3462 VDD.t3461 VDD.t3462 VDD.t1799 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2138 a_89563_n36322# a_89163_n36382.t11 a_89033_n36322.t3 VDD.t548 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2139 OUT.t13 a_35502_24538.t38 a_33249_35053.t97 VSS.t193 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2140 a_59411_n7138# a_50751_n19729.t159 a_58851_n7138# VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2141 VDD.t3460 VDD.t3459 VDD.t3460 VDD.t630 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2142 VDD.t3458 VDD.t3457 VDD.t3458 VDD.t1442 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2143 VDD.t3456 VDD.t3455 VDD.t3456 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2144 VSS.t2652 VSS.t2651 VSS.t2652 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2145 VSS.t314 a_106830_10388.t13 a_107230_12380# VDD.t519 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2146 a_33249_35053.t133 a_35502_25545.t49 VSS.t15 VSS.t14 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2147 VDD.t3454 VDD.t3453 VDD.t3454 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2148 VSS.t2650 VSS.t2649 VSS.t2650 VSS.t148 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2149 a_30682_n34390# a_30152_n35156.t19 a_30152_n36322.t6 VDD.t622 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2150 a_67111_n13318# a_50751_n19729.t160 a_66551_n13318# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2151 VDD.t3452 VDD.t3451 VDD.t3452 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2152 VDD.t3450 VDD.t3449 VDD.t3450 VDD.t2231 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2153 VDD.t3448 VDD.t3447 VDD.t3448 VDD.t1218 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2154 a_33249_35053.t28 a_33379_34917.t31 a_33249_48695.t42 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2155 VDD.t3446 VDD.t3445 VDD.t3446 VDD.t545 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2156 VSS.t2648 VSS.t2647 VSS.t2648 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2157 a_81735_n9675# a_71281_n10073.t146 a_81205_n9675# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2158 VDD.t3444 VDD.t3443 VDD.t3444 VDD.t2299 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X2159 VSS.t2646 VSS.t2645 VSS.t2646 VSS.t740 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2160 VSS.t2644 VSS.t2643 VSS.t2644 VSS.t638 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2161 VSS.t2642 VSS.t2641 VSS.t2642 VSS.t908 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2162 a_72603_n10973# I1N.t2 I1N.t3 VSS.t429 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X2163 VSS.t2640 VSS.t2639 VSS.t2640 VSS.t760 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2164 VDD.t141 a_31699_20742.t119 a_33249_48695.t275 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2165 a_98829_n9675# a_71281_n8397.t163 a_98299_n9675# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2166 a_88839_n15905# a_71281_n10073.t147 a_88271_n15905# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2167 VSS.t2638 VSS.t2637 VSS.t2638 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2168 VDD.t3442 VDD.t3441 VDD.t3442 VDD.t1799 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2169 a_30682_12380# a_30152_10448.t10 a_30152_10448.t11 VDD.t302 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2170 VDD.t3440 VDD.t3439 VDD.t3440 VDD.t603 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2171 VDD.t4917 a_52635_34067.t123 a_52635_49681.t143 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2172 VSS.t2636 VSS.t2635 VSS.t2636 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2173 a_42047_n17801# a_31953_n19727.t165 a_41487_n16904# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2174 VSS.t2634 VSS.t2633 VSS.t2634 VSS.t354 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2175 a_77225_n29181.t8 a_77225_n29181.t7 a_79151_n28415# VSS.t380 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2176 VSS.t2632 VSS.t2631 VSS.t2632 VSS.t859 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2177 VDD.t4781 a_83153_n36322.t12 a_90935_n28415# VSS.t455 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2178 a_55635_n34390# a_53829_n36382.t17 VSS.t175 VDD.t367 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2179 VDD.t3438 VDD.t3437 VDD.t3438 VDD.t1218 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2180 VSS.t2630 VSS.t2629 VSS.t2630 VSS.t265 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2181 a_52635_48695.t149 a_52635_34067.t124 VDD.t4916 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2182 VDD.t3436 VDD.t3435 VDD.t3436 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2183 VDD.t3434 VDD.t3433 VDD.t3434 VDD.t309 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2184 a_38619_n13316# a_31953_n19727.t166 a_38097_n13316# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2185 VSS.t2628 VSS.t2627 VSS.t2628 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2186 VDD.t3432 VDD.t3431 VDD.t3432 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2187 VDD.t3430 VDD.t3429 VDD.t3430 VDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2188 a_64243_n1756.t1 a_65486_11614.t12 a_71864_5639# VSS.t424 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2189 a_52585_n17803# a_50751_n19729.t161 a_52063_n18700# VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2190 VSS.t2626 VSS.t2625 VSS.t2626 VSS.t196 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2191 VCM.t2 a_33379_34007.t0 cap_mim_2f0_m4m5_noshield c_width=9.8u c_length=9.8u
X2192 VSS.t2624 VSS.t2623 VSS.t2624 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2193 VDD.t3428 VDD.t3427 VDD.t3428 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2194 a_84547_n8770# a_71281_n10073.t148 a_83709_n8770# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2195 VDD.t3426 VDD.t3425 VDD.t3426 VDD.t930 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2196 VSS.t2622 VSS.t2621 VSS.t2622 VSS.t687 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2197 VDD.t3424 VDD.t3422 VDD.t3424 VDD.t3423 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2198 a_52635_49681.t33 a_35922_19591.t80 OUT.t74 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2199 VDD.t3421 VDD.t3420 VDD.t3421 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2200 a_60109_n34390# a_53699_n35156.t7 a_53829_n36382.t6 VDD.t543 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2201 VDD.t3419 VDD.t3418 VDD.t3419 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2202 a_33249_35053.t132 a_35502_25545.t50 VSS.t47 VSS.t29 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2203 a_47991_n29313.t0 a_47819_n36322.t12 a_54197_n27257# VSS.t304 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2204 VDD.t3417 VDD.t3416 VDD.t3417 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2205 VDD.t3415 VDD.t3414 VDD.t3415 VDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2206 a_85129_n30339# a_83325_n29313.t0 a_31831_n5342.t2 VSS.t286 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2207 VDD.t3413 VDD.t3412 VDD.t3413 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2208 VDD.t3411 VDD.t3410 VDD.t3411 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2209 a_78344_10448.t4 a_71366_11614.t5 a_77776_13546# VDD.t3570 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2210 a_36032_13546.t1 a_53829_10388.t11 a_55635_13546# VDD.t3747 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2211 a_33249_48695.t43 a_33379_34917.t32 a_33249_35053.t29 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2212 VSS.t2620 VSS.t2619 VSS.t2620 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2213 a_58851_n2653# a_50751_n19729.t162 a_58329_n3550# VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2214 VSS.t2618 VSS.t2617 VSS.t2618 VSS.t687 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2215 a_106676_n30339.t2 a_106830_n36382.t13 a_107230_n36322# VDD.t845 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2216 VDD.t3409 VDD.t3408 VDD.t3409 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2217 VDD.t3407 VDD.t3406 VDD.t3407 VDD.t836 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2218 a_33249_48695.t274 a_31699_20742.t120 VDD.t142 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2219 VDD.t3405 VDD.t3404 VDD.t3405 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2220 a_52635_48695.t148 a_52635_34067.t125 VDD.t4915 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2221 VSS.t2616 VSS.t2615 VSS.t2616 VSS.t1256 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2222 a_81205_n14095.t1 a_89163_10388.t15 a_90969_12380# VDD.t553 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2223 VDD.t3403 VDD.t3402 VDD.t3403 VDD.t1799 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2224 VDD.t3401 VDD.t3400 VDD.t3401 VDD.t27 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2225 VSS.t2614 VSS.t2613 VSS.t2614 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2226 VDD.t3399 VDD.t3398 VDD.t3399 VDD.t353 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2227 VDD.t3397 VDD.t3396 VDD.t3397 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2228 VDD.t3395 VDD.t3394 VDD.t3395 VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2229 VSS.t2612 VSS.t2611 VSS.t2612 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2230 VDD.t3393 VDD.t3392 VDD.t3393 VDD.t1052 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2231 VSS.t2610 VSS.t2609 VSS.t2610 VSS.t1426 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2232 VDD.t3391 VDD.t3390 VDD.t3391 VDD.t3013 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2233 VSS.t2608 VSS.t2607 VSS.t2608 VSS.t757 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2234 VDD.t3389 VDD.t3388 VDD.t3389 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2235 VSS.t2606 VSS.t2605 VSS.t2606 VSS.t304 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2236 VDD.t3387 VDD.t3386 VDD.t3387 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2237 VSS.t2604 VSS.t2603 VSS.t2604 VSS.t653 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2238 a_46879_n19595# a_31953_n19727.t167 a_46319_n19595# VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2239 a_78344_10448.t1 a_71366_11614.t6 a_77776_11614# VDD.t3570 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2240 a_53699_11614.t1 a_53829_10388.t12 a_55635_11614# VDD.t3747 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2241 VDD.t3385 VDD.t3384 VDD.t3385 VDD.t823 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2242 a_35922_19591.t1 a_35922_19591.t0 a_46274_24920# VDD.t390 pfet_03v3 ad=0.78p pd=3.7u as=0.78p ps=3.7u w=1.2u l=2u
X2243 VSS.t2602 VSS.t2601 VSS.t2602 VSS.t905 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2244 a_89531_n30339# a_83153_n36322.t13 a_89009_n30339.t0 VSS.t454 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2245 a_113037_n18620# a_71281_n8397.t164 a_112199_n18620# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2246 VSS.t2600 VSS.t2599 VSS.t2600 VSS.t261 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2247 a_40613_n3548# a_31953_n19727.t168 a_41487_n5342# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2248 a_93131_n9675# a_71281_n10073.t149 a_92601_n9675# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2249 VSS.t2598 VSS.t2597 VSS.t2598 VSS.t156 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2250 VDD.t3383 VDD.t3382 VDD.t3383 VDD.t810 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2251 VSS.t2596 VSS.t2595 VSS.t2596 VSS.t229 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2252 VDD.t3381 VDD.t3380 VDD.t3381 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2253 VDD.t3379 VDD.t3378 VDD.t3379 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2254 VSS.t2594 VSS.t2593 VSS.t2594 VSS.t853 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2255 VDD.t3377 VDD.t3376 VDD.t3377 VDD.t38 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2256 a_39179_n16904# a_31953_n19727.t169 a_38619_n16904# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2257 a_38097_n16007.t2 a_39179_n19595.t0 a_48391_n30339# VSS.t340 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2258 a_32913_n8033# a_31953_n19727.t170 a_32353_n7136# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2259 VSS.t2592 VSS.t2591 VSS.t2592 VSS.t681 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2260 VDD.t3375 VDD.t3374 VDD.t3375 VDD.t697 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2261 VDD.t3373 VDD.t3372 VDD.t3373 VDD.t1155 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2262 VDD.t3371 VDD.t3370 VDD.t3371 VDD.t1515 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2263 VDD.t3369 VDD.t3368 VDD.t3369 VDD.t2924 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2264 VDD.t3367 VDD.t3366 VDD.t3367 VDD.t305 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2265 VDD.t3365 VDD.t3364 VDD.t3365 VDD.t1405 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2266 VDD.t3363 VDD.t3362 VDD.t3363 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2267 VSS.t2590 VSS.t2589 VSS.t2590 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2268 a_52635_49681.t34 a_35922_19591.t81 OUT.t73 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2269 VSS.t2588 VSS.t2587 VSS.t2588 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2270 VSS.t2586 VSS.t2585 VSS.t2586 VSS.t213 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2271 a_100803_n6960# a_71281_n8397.t165 a_100235_n6960# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2272 a_71281_n8397.t47 a_71281_n8397.t46 VDD.t455 VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2273 VDD.t143 a_31699_20742.t121 a_33249_48695.t273 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2274 a_105365_n2435# a_71281_n8397.t166 a_104527_n2435# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2275 VSS.t2584 VSS.t2583 VSS.t2584 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2276 VSS.t2582 VSS.t2581 VSS.t2582 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2277 VSS.t2580 VSS.t2579 VSS.t2580 VSS.t151 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2278 VSS.t2578 VSS.t2577 VSS.t2578 VSS.t868 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2279 a_33249_48695.t272 a_31699_20742.t122 VDD.t144 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2280 a_60285_n16906# a_50751_n19729.t163 a_59763_n16906# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2281 VSS.t2576 VSS.t2575 VSS.t2576 VSS.t3 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2282 a_106830_10388.t1 a_112559_4481.t17 a_114485_4481# VSS.t292 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2283 VSS.t167 a_41891_4481.t18 a_42413_4481# VSS.t166 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2284 a_33249_48695.t271 a_31699_20742.t123 VDD.t145 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2285 a_95443_n36322# a_89033_n35156.t10 a_89163_n36382.t7 VDD.t795 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2286 a_95943_n8770# a_71281_n10073.t150 a_95105_n8770# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2287 VDD.t3361 VDD.t3360 VDD.t3361 VDD.t2464 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2288 VDD.t3359 VDD.t3358 VDD.t3359 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2289 VSS.t2574 VSS.t2573 VSS.t2574 VSS.t896 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2290 VDD.t3357 VDD.t3356 VDD.t3357 VDD.t1155 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2291 VDD.t3355 VDD.t3353 VDD.t3355 VDD.t3354 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2292 a_53699_13546.t2 a_71496_10388.t15 a_73302_13546# VDD.t352 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2293 VDD.t3352 VDD.t3351 VDD.t3352 VDD.t789 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2294 VDD.t3350 VDD.t3349 VDD.t3350 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2295 a_42442_10448# a_30324_4421.t1 a_41891_4481.t0 VDD.t288 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2296 VDD.t3348 VDD.t3347 VDD.t3348 VDD.t1015 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2297 VDD.t3346 VDD.t3345 VDD.t3346 VDD.t524 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2298 a_114485_6405# a_112559_4481.t18 VSS.t300 VSS.t297 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2299 VSS.t2572 VSS.t2571 VSS.t2572 VSS.t1385 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2300 VDD.t3344 VDD.t3343 VDD.t3344 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2301 VDD.t3342 VDD.t3341 VDD.t3342 VDD.t320 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2302 VSS.t2570 VSS.t2569 VSS.t2570 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2303 VDD.t3340 VDD.t3339 VDD.t3340 VDD.t2118 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2304 VDD.t3338 VDD.t3337 VDD.t3338 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2305 a_106501_n7865# a_71281_n8397.t167 a_105933_n7865# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2306 a_45445_n14213# a_31953_n19727.t171 a_44885_n14213# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2307 a_104527_n17715# a_71281_n8397.t168 a_103997_n21335# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2308 VDD.t454 a_71281_n8397.t44 a_71281_n8397.t45 VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2309 VDD.t3336 VDD.t3335 VDD.t3336 VDD.t2447 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2310 VSS.t2568 VSS.t2567 VSS.t2568 VSS.t690 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2311 a_71281_n10073.t51 a_71281_n10073.t50 VDD.t334 VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2312 VSS.t86 a_31953_n19727.t52 a_31953_n19727.t53 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2313 a_48313_n4445# a_31953_n19727.t172 a_47753_n3548# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2314 a_112199_n19525# a_71281_n8397.t169 a_111631_n19525# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2315 VSS.t85 a_31953_n19727.t50 a_31953_n19727.t51 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2316 VDD.t146 a_31699_20742.t124 a_33249_48695.t270 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2317 a_66551_n14215# a_50751_n19729.t164 a_66029_n14215# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2318 a_71366_11614.t1 a_71496_10388.t16 a_73302_11614# VDD.t352 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2319 a_61515_n34390# a_47991_n29313.t1 a_60677_n36322.t1 VDD.t544 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2320 VSS.t2566 VSS.t2565 VSS.t2566 VSS.t644 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2321 VSS.t2564 VSS.t2563 VSS.t2564 VSS.t1315 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2322 a_52635_34067.t64 a_35502_24538.t39 a_33249_34067.t11 VSS.t193 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2323 a_52635_49681.t35 a_35922_19591.t82 OUT.t72 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2324 VSS.t2562 VSS.t2561 VSS.t2562 VSS.t884 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2325 VDD.t342 a_71281_n10073.t48 a_71281_n10073.t49 VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2326 a_104527_n9675# a_71281_n8397.t170 a_103997_n9675# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2327 a_65677_n19597# a_50751_n19729.t165 a_65117_n18700# VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2328 a_112559_n29181.t0 a_100992_n29313.t2 a_114516_n36322# VDD.t538 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2329 a_56895_n16009.t2 a_100992_4421.t2 a_101392_4481# VSS.t162 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2330 VSS.t2560 VSS.t2559 VSS.t2560 VSS.t676 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2331 a_45445_n6239# a_31953_n19727.t173 a_44885_n6239# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2332 a_47819_n36322.t6 a_39179_n19595.t0 a_49795_n29181# VSS.t337 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2333 a_89407_n15000# a_71281_n10073.t151 a_88839_n15000# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2334 VDD.t3334 VDD.t3333 VDD.t3334 VDD.t1322 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2335 a_33249_34067.t76 a_33379_34007.t34 a_33249_48695.t105 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2336 a_32353_n2651# a_31953_n19727.t174 a_31831_n2651# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2337 VSS.t2558 VSS.t2557 VSS.t2558 VSS.t877 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2338 VSS.t2556 VSS.t2555 VSS.t2556 VSS.t340 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2339 a_71281_n8397.t43 a_71281_n8397.t42 VDD.t453 VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2340 a_52635_48695.t147 a_52635_34067.t126 VDD.t4914 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2341 VDD.t3332 VDD.t3331 VDD.t3332 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2342 a_113081_4481# a_112559_4481.t2 a_112559_4481.t3 VSS.t293 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2343 VDD.t3330 VDD.t3329 VDD.t3330 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2344 VSS.t2554 VSS.t2553 VSS.t2554 VSS.t944 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2345 VSS.t2552 VSS.t2551 VSS.t2552 VSS.t484 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X2346 a_100803_n15000# a_71281_n8397.t171 a_100235_n15000# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2347 a_34347_n2651# a_31953_n19727.t175 a_33787_n2651# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2348 a_65486_11614.t7 a_64243_n1756.t1 a_67462_4481# VSS.t378 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2349 VDD.t3328 VDD.t3327 VDD.t3328 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2350 a_41487_n17801# a_31953_n19727.t176 a_40965_n18698# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2351 a_35781_n7136# a_31953_n19727.t177 a_35221_n7136# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2352 VSS.t2550 VSS.t2549 VSS.t2550 VSS.t811 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2353 a_57977_n12421.t0 a_100820_11614.t9 a_107198_5639# VSS.t153 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2354 VSS.t2548 VSS.t2547 VSS.t2548 VSS.t397 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2355 a_33249_48695.t269 a_31699_20742.t125 VDD.t147 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2356 a_52635_49681.t142 a_52635_34067.t127 VDD.t4913 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2357 VSS.t2546 VSS.t2545 VSS.t2546 VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2358 a_42413_4481# a_41891_4481.t3 a_41891_4481.t4 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2359 a_35221_n18698# a_31953_n19727.t178 a_34699_n18698# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2360 VDD.t148 a_31699_20742.t126 a_33249_48695.t268 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2361 a_33249_34067.t75 a_33379_34007.t35 a_33249_48695.t10 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2362 a_105933_n21335# a_71281_n8397.t172 a_105365_n21335# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2363 a_79151_4481# a_77225_4481.t15 VSS.t322 VSS.t319 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2364 a_107230_13546# a_106830_10388.t14 OUT.t0 VDD.t522 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2365 a_106809_n5150.t0 a_103997_n8770.t6 a_113110_n36322# VDD.t537 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2366 a_67462_6405# a_64243_n1756.t2 a_63161_n5344.t1 VSS.t289 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2367 VSS.t2544 VSS.t2543 VSS.t2544 VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2368 VDD.t3326 VDD.t3325 VDD.t3326 VDD.t390 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X2369 VSS.t2542 VSS.t2541 VSS.t2542 VSS.t495 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2370 a_33249_48695.t11 a_33379_34007.t36 a_33249_34067.t74 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2371 VSS.t2540 VSS.t2539 VSS.t2540 VSS.t525 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2372 a_35502_25545.t9 a_31699_20742.t127 VDD.t149 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2373 a_101392_n29181# a_100992_n29313.t0 a_100820_n35156.t0 VSS.t331 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2374 a_72603_n8397# I1N.t7 a_71281_n8397.t73 VSS.t429 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X2375 VSS.t2538 VSS.t2537 VSS.t2538 VSS.t908 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2376 VSS.t2536 VSS.t2535 VSS.t2536 VSS.t792 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2377 a_89163_10388.t1 a_94892_4481.t14 a_96818_6405# VSS.t396 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2378 VDD.t3324 VDD.t3323 VDD.t3324 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2379 VDD.t3322 VDD.t3321 VDD.t3322 VDD.t2399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2380 a_107230_11614# a_106830_10388.t15 a_86903_n14095.t1 VDD.t522 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2381 VDD.t3320 VDD.t3319 VDD.t3320 VDD.t2573 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2382 a_84547_n8770# a_71281_n10073.t152 a_83709_n7865# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2383 VDD.t3318 VDD.t3317 VDD.t3318 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2384 a_96818_n27257# a_94892_n29181.t13 VSS.t356 VSS.t354 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2385 VDD.t3316 VDD.t3315 VDD.t3316 VDD.t519 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2386 VDD.t3314 VDD.t3313 VDD.t3314 VDD.t720 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2387 a_104527_n21335# a_71281_n8397.t173 a_103997_n21335# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2388 VDD.t3312 VDD.t3311 VDD.t3312 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2389 a_44885_n17801# a_31953_n19727.t179 a_44363_n17801# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2390 VDD.t3310 VDD.t3309 VDD.t3310 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2391 a_44885_n1754# a_31953_n19727.t180 a_44363_n2651# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2392 a_49755_n36322# a_47819_n35156.t17 VDD.t4795 VDD.t707 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2393 VSS.t2534 VSS.t2533 VSS.t2534 VSS.t699 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2394 VSS.t2532 VSS.t2531 VSS.t2532 VSS.t1064 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2395 VSS.t2530 VSS.t2529 VSS.t2530 VSS.t1157 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2396 VDD.t3308 VDD.t3307 VDD.t3308 VDD.t1086 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2397 a_57417_n5344# a_50751_n19729.t166 a_48951_4481.t0 VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2398 a_46879_n2651# a_31953_n19727.t181 a_46319_n1754# VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2399 a_79182_n34390# a_65658_n29313.t1 a_78344_n36322.t2 VDD.t2382 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2400 VSS.t2528 VSS.t2527 VSS.t2528 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2401 a_89407_n20430# a_71281_n10073.t153 a_88839_n20430# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2402 VSS.t2526 VSS.t2525 VSS.t2526 VSS.t668 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2403 VDD.t3306 VDD.t3305 VDD.t3306 VDD.t1142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2404 VDD.t3304 VDD.t3303 VDD.t3304 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2405 VSS.t2524 VSS.t2523 VSS.t2524 VSS.t553 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2406 a_33249_48695.t12 a_33379_34007.t37 a_33249_34067.t73 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2407 a_51151_n14215# a_50751_n19729.t167 a_50629_n15112# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2408 VSS.t2522 VSS.t2521 VSS.t2522 VSS.t323 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2409 a_100803_n20430# a_71281_n8397.t174 a_100235_n20430# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2410 VSS.t2520 VSS.t2519 VSS.t2520 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2411 VSS.t2518 VSS.t2517 VSS.t2518 VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2412 VSS.t2516 VSS.t2515 VSS.t2516 VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2413 a_50629_n16009.t1 a_83325_4421.t0 a_83725_6405# VSS.t311 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2414 VDD.t4912 a_52635_34067.t128 a_52635_48695.t146 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2415 a_106501_n18620# a_71281_n8397.t175 a_105933_n18620# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2416 VDD.t3302 VDD.t3301 VDD.t3302 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2417 a_114485_n29181# a_112559_n29181.t15 VSS.t416 VSS.t413 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2418 VDD.t3300 VDD.t3299 VDD.t3300 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2419 a_87433_n6055# a_71281_n10073.t154 a_86903_n5150# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2420 OUT.t12 a_35502_24538.t40 a_33249_35053.t103 VSS.t192 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2421 VSS.t2514 VSS.t2513 VSS.t2514 VSS.t615 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2422 VSS.t2512 VSS.t2511 VSS.t2512 VSS.t155 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2423 VDD.t3298 VDD.t3297 VDD.t3298 VDD.t1086 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2424 VSS.t2510 VSS.t2509 VSS.t2510 VSS.t1253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2425 VDD.t4911 a_52635_34067.t129 a_52635_49681.t141 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2426 a_55601_n28415# a_47819_n36322.t13 a_39179_n19595.t0 VSS.t305 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2427 a_50751_n19729.t43 a_50751_n19729.t42 VSS.t240 VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2428 VDD.t3296 VDD.t3295 VDD.t3296 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2429 a_101641_n8770# a_71281_n8397.t176 a_100803_n8770# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2430 VSS.t2508 VSS.t2507 VSS.t2508 VSS.t1256 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2431 a_77776_n34390# a_71366_n35156.t6 a_71496_n36382.t6 VDD.t2344 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2432 a_34347_n13316# a_31953_n19727.t182 a_33787_n13316# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2433 a_67111_n13318# a_50751_n19729.t168 a_66551_n12421# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2434 VDD.t3294 VDD.t3293 VDD.t3294 VDD.t1262 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2435 a_113037_n17715# a_71281_n8397.t177 a_112507_n17715.t1 VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2436 VSS.t2506 VSS.t2505 VSS.t2506 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2437 VSS.t2504 VSS.t2503 VSS.t2504 VSS.t1306 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2438 a_96818_6405# a_94892_4481.t15 VSS.t3639 VSS.t1303 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2439 VSS.t2502 VSS.t2501 VSS.t2502 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2440 VSS.t2500 VSS.t2499 VSS.t2500 VSS.t576 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2441 VSS.t2498 VSS.t2497 VSS.t2498 VSS.t891 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2442 VSS.t2496 VSS.t2495 VSS.t2496 VSS.t604 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2443 VDD.t3292 VDD.t3291 VDD.t3292 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2444 VSS.t2494 VSS.t2493 VSS.t2494 VSS.t148 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2445 a_83141_n19525# a_71281_n10073.t155 a_82573_n19525# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2446 VSS.t2492 VSS.t2491 VSS.t2492 VSS.t1294 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2447 VDD.t3290 VDD.t3289 VDD.t3290 VDD.t510 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2448 VSS.t2490 VSS.t2489 VSS.t2490 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2449 VSS.t2488 VSS.t2487 VSS.t2488 VSS.t0 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2450 VSS.t2486 VSS.t2485 VSS.t2486 VSS.t748 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2451 VSS.t2484 VSS.t2483 VSS.t2484 VSS.t1287 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2452 VSS.t2482 VSS.t2481 VSS.t2482 VSS.t283 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2453 VDD.t4784 a_83153_10448.t13 a_83683_13546# VDD.t3354 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2454 VDD.t3288 VDD.t3287 VDD.t3288 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2455 VDD.t150 a_31699_20742.t128 a_33249_48695.t267 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2456 a_95105_n14095# a_71281_n10073.t156 a_94537_n14095# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2457 VDD.t3286 VDD.t3285 VDD.t3286 VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2458 VSS.t2480 VSS.t2479 VSS.t2480 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2459 VSS.t2478 VSS.t2477 VSS.t2478 VSS.t105 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2460 VDD.t3284 VDD.t3283 VDD.t3284 VDD.t1180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2461 VSS.t2476 VSS.t2474 VSS.t2476 VSS.t2475 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X2462 VDD.t3282 VDD.t3281 VDD.t3282 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2463 a_63683_n16906# a_50751_n19729.t169 a_63161_n17803# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2464 a_90245_n15000# a_71281_n10073.t157 a_89407_n14095# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2465 a_88839_n6960# a_71281_n10073.t158 a_88271_n6960# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2466 VDD.t151 a_31699_20742.t129 a_33249_48695.t266 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2467 a_53675_7563.t2 a_47819_11614.t15 a_55601_4481# VSS.t307 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2468 a_90969_10448# a_89163_10388.t16 a_89009_7563.t2 VDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2469 VDD.t3280 VDD.t3279 VDD.t3280 VDD.t1042 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2470 VDD.t35 a_31699_20742.t27 a_31699_20742.t28 VDD.t34 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2471 a_95943_n8770# a_71281_n10073.t159 a_95105_n7865# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2472 a_112559_4481.t8 a_100992_4421.t1 a_114516_13546# VDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2473 a_33249_48695.t265 a_31699_20742.t130 VDD.t152 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2474 VDD.t4910 a_52635_34067.t130 a_52635_48695.t145 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2475 VDD.t3278 VDD.t3277 VDD.t3278 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2476 a_33249_35053.t30 a_33379_34917.t33 a_33249_48695.t44 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2477 VSS.t440 a_36162_n36382.t8 a_36562_n34390# VDD.t2302 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2478 VDD.t4909 a_52635_34067.t131 a_52635_48695.t144 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2479 VSS.t2473 VSS.t2472 VSS.t2473 VSS.t284 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2480 VSS.t2471 VSS.t2470 VSS.t2471 VSS.t498 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2481 VSS.t2469 VSS.t2468 VSS.t2469 VSS.t618 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2482 a_89407_n1530# a_71281_n10073.t160 a_88839_n1530# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2483 VSS.t2467 VSS.t2466 VSS.t2467 VSS.t550 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2484 a_67422_n35156# a_65486_n35156.t19 VDD.t9 VDD.t6 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2485 a_83725_6405# a_83325_4421.t0 a_83153_10448.t0 VSS.t310 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2486 VSS.t447 a_59558_n29181.t16 a_60080_n30339# VSS.t401 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2487 a_81735_n19525# a_71281_n10073.t161 a_81205_n19525# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2488 a_51151_n8932# a_50751_n19729.t170 a_50629_n8932# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2489 a_40053_n8033# a_31953_n19727.t183 a_39531_n8033# VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2490 VDD.t4785 a_83153_10448.t14 a_83683_11614# VDD.t3354 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2491 a_52635_48695.t51 a_35922_19591.t83 a_52635_34067.t32 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2492 a_93969_n9675# a_71281_n10073.t162 a_93131_n9675# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2493 a_53145_n8932# a_50751_n19729.t171 a_52585_n8932# VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2494 VDD.t3276 VDD.t3275 VDD.t3276 VDD.t630 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2495 VDD.t3274 VDD.t3273 VDD.t3274 VDD.t638 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2496 VSS.t2465 VSS.t2464 VSS.t2465 VSS.t817 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X2497 VDD.t3272 VDD.t3271 VDD.t3272 VDD.t1042 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2498 VDD.t3270 VDD.t3269 VDD.t3270 VDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2499 VDD.t3268 VDD.t3267 VDD.t3268 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2500 a_112559_4481.t10 a_100992_4421.t1 a_114516_11614# VDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2501 VDD.t3266 VDD.t3265 VDD.t3266 VDD.t496 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2502 a_94537_n4245# a_71281_n10073.t163 a_93969_n4245# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2503 a_30682_n36322# a_30152_n35156.t20 a_30152_n36322.t7 VDD.t622 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2504 a_88839_n14095# a_71281_n10073.t164 a_88271_n14095# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2505 a_35781_n19595# a_31953_n19727.t184 a_35221_n19595# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2506 a_41487_n8033# a_31953_n19727.t185 a_40965_n8033# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2507 VDD.t3264 VDD.t3263 VDD.t3264 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2508 VDD.t3262 VDD.t3261 VDD.t3262 VDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2509 VSS.t2463 VSS.t2462 VSS.t2463 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2510 a_35221_n7136# a_31953_n19727.t186 a_34699_n8033# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2511 a_67422_n33224# a_65486_n35156.t20 VDD.t10 VDD.t6 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2512 a_89407_n15905# a_71281_n10073.t165 a_88839_n15905# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2513 VDD.t3260 VDD.t3259 VDD.t3260 VDD.t2254 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2514 VSS.t2461 VSS.t2460 VSS.t2461 VSS.t528 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2515 VDD.t3258 VDD.t3257 VDD.t3258 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2516 a_112507_n17715.t0 a_71281_n8397.t178 a_112199_n21335# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2517 VDD.t3256 VDD.t3255 VDD.t3256 VDD.t1206 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2518 VDD.t3254 VDD.t3253 VDD.t3254 VDD.t603 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2519 a_100803_n15905# a_71281_n8397.t179 a_100235_n15905# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2520 a_36562_13546# a_36162_10388.t15 a_36032_13546.t3 VDD.t3423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2521 VSS.t2459 VSS.t2458 VSS.t2459 VSS.t147 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2522 VSS.t2457 VSS.t2456 VSS.t2457 VSS.t284 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2523 VDD.t3252 VDD.t3251 VDD.t3252 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2524 VDD.t3250 VDD.t3249 VDD.t3250 VDD.t598 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2525 a_55635_n36322# a_53829_n36382.t18 a_53675_n27257.t0 VDD.t367 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2526 VSS.t2455 VSS.t2454 VSS.t2455 VSS.t490 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2527 VDD.t3248 VDD.t3247 VDD.t3248 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2528 VDD.t3246 VDD.t3245 VDD.t3246 VDD.t917 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2529 a_41660_19698# a_35502_24538.t41 a_41100_20251# VSS.t186 nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X2530 VSS.t2453 VSS.t2452 VSS.t2453 VSS.t525 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2531 a_65117_n17803# a_50751_n19729.t172 a_64595_n18700# VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2532 a_55601_4481# a_47819_11614.t16 a_47991_4421.t0 VSS.t305 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2533 a_35502_24538.t17 a_31699_20742.t131 VDD.t153 VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2534 VDD.t3244 VDD.t3243 VDD.t3244 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2535 VDD.t3242 VDD.t3241 VDD.t3242 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2536 a_71281_n10073.t47 a_71281_n10073.t46 VDD.t354 VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2537 a_53829_n36382.t2 a_59558_n29181.t17 a_61484_n29181# VSS.t398 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2538 VSS.t2451 VSS.t2450 VSS.t2451 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2539 VDD.t3240 VDD.t3239 VDD.t3240 VDD.t1957 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2540 a_60109_n36322# a_53699_n35156.t8 a_53829_n36382.t7 VDD.t543 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2541 a_59411_n17803# a_50751_n19729.t173 a_58851_n17803# VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2542 VDD.t452 a_71281_n8397.t40 a_71281_n8397.t41 VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2543 a_83141_n6960# a_71281_n10073.t166 a_82573_n6960# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2544 a_36562_11614# a_36162_10388.t16 a_36032_11614.t2 VDD.t3423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2545 VDD.t3238 VDD.t3237 VDD.t3238 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2546 VDD.t3236 VDD.t3235 VDD.t3236 VDD.t1333 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2547 a_33379_34007.t27 IN_POS.t0 cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
X2548 a_59558_4481.t7 a_59558_4481.t6 a_61484_5639# VSS.t398 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2549 VDD.t3234 VDD.t3233 VDD.t3234 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2550 a_33249_35053.t100 a_35502_24538.t42 OUT.t11 VSS.t195 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2551 VDD.t4778 a_65486_11614.t13 a_73268_6405# VSS.t422 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2552 VDD.t3232 VDD.t3231 VDD.t3232 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2553 a_100235_n6960# a_71281_n8397.t180 a_99667_n6960# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2554 a_83709_n13190# a_71281_n10073.t167 a_83141_n13190# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2555 a_46319_n1754# a_31953_n19727.t187 VSS.t113 VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2556 VDD.t3230 VDD.t3229 VDD.t3230 VDD.t406 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2557 VDD.t3228 VDD.t3227 VDD.t3228 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2558 VSS.t2449 VSS.t2448 VSS.t2449 VSS.t1064 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2559 a_47753_n6239# a_31953_n19727.t188 a_47231_n6239# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2560 VSS.t2447 VSS.t2446 VSS.t2447 VSS.t330 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2561 VDD.t3226 VDD.t3225 VDD.t3226 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2562 VDD.t3224 VDD.t3223 VDD.t3224 VDD.t1936 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2563 a_52635_49681.t36 a_35922_19591.t84 OUT.t71 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2564 VDD.t3222 VDD.t3221 VDD.t3222 VDD.t598 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2565 VSS.t2445 VSS.t2444 VSS.t2445 VSS.t63 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2566 VDD.t3220 VDD.t3219 VDD.t3220 VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2567 VSS.t2443 VSS.t2442 VSS.t2443 VSS.t568 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2568 a_81735_n3340# a_71281_n10073.t168 a_81205_n4245# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2569 a_52635_48695.t143 a_52635_34067.t132 VDD.t4908 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2570 VDD.t3218 VDD.t3217 VDD.t3218 VDD.t833 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2571 a_71281_n8397.t39 a_71281_n8397.t38 VDD.t451 VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2572 VDD.t3216 VDD.t3215 VDD.t3216 VDD.t798 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2573 VSS.t2441 VSS.t2440 VSS.t2441 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2574 a_94892_4481.t9 a_83325_4421.t1 a_96849_13546# VDD.t500 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2575 VDD.t3214 VDD.t3213 VDD.t3214 VDD.t1378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2576 a_99667_n15000# a_71281_n8397.t181 a_98829_n15000# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2577 a_59411_n17803# a_50751_n19729.t174 a_60285_n16009# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2578 a_60677_10448.t3 a_47991_4421.t1 a_60109_10448# VDD.t664 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2579 a_71281_n8397.t37 a_71281_n8397.t36 VDD.t450 VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2580 a_98829_n3340# a_71281_n8397.t182 a_98299_n4245# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2581 VDD.t3212 VDD.t3211 VDD.t3212 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2582 VSS.t84 a_31953_n19727.t48 a_31953_n19727.t49 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2583 VSS.t2439 VSS.t2438 VSS.t2439 VSS.t63 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2584 VSS.t2437 VSS.t2436 VSS.t2437 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2585 VSS.t2435 VSS.t2434 VSS.t2435 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2586 VSS.t2433 VSS.t2432 VSS.t2433 VSS.t763 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X2587 a_48313_n2651# a_31953_n19727.t189 a_47753_n2651# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2588 a_111063_n15000# a_71281_n8397.t183 a_110225_n15000# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2589 a_33787_n14213# a_31953_n19727.t190 a_33265_n14213# VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2590 VSS.t2431 VSS.t2430 VSS.t2431 VSS.t501 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2591 a_59411_n2653# a_50751_n19729.t175 a_58851_n1756# VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2592 VDD.t3210 VDD.t3209 VDD.t3210 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2593 a_113037_n6960# a_71281_n8397.t184 a_112199_n6960# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2594 VSS.t2429 VSS.t2428 VSS.t2429 VSS.t814 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2595 VSS.t2427 VSS.t2426 VSS.t2427 VSS.t979 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2596 VDD.t3208 VDD.t3207 VDD.t3208 VDD.t1299 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2597 VSS.t2425 VSS.t2424 VSS.t2425 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2598 VSS.t2423 VSS.t2422 VSS.t2423 VSS.t168 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2599 VDD.t3206 VDD.t3205 VDD.t3206 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2600 VSS.t2421 VSS.t2420 VSS.t2421 VSS.t1157 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2601 a_45445_n5342.t1 a_31953_n19727.t191 a_44885_n5342# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2602 VDD.t3204 VDD.t3203 VDD.t3204 VDD.t1177 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2603 VDD.t3202 VDD.t3201 VDD.t3202 VDD.t2680 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2604 a_33249_48695.t45 a_33379_34917.t34 a_33249_35053.t31 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2605 a_30152_10448.t2 a_30324_4421.t0 a_32128_7563# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2606 VDD.t3200 VDD.t3199 VDD.t3200 VDD.t2774 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2607 a_94892_4481.t10 a_83325_4421.t1 a_96849_11614# VDD.t500 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2608 VDD.t3198 VDD.t3197 VDD.t3198 VDD.t979 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2609 VDD.t449 a_71281_n8397.t34 a_71281_n8397.t35 VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2610 VDD.t3196 VDD.t3195 VDD.t3196 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2611 a_33249_35053.t131 a_35502_25545.t51 VSS.t164 VSS.t14 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2612 VSS.t2419 VSS.t2418 VSS.t2419 VSS.t490 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2613 VSS.t2417 VSS.t2416 VSS.t2417 VSS.t834 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2614 a_87433_n4245# a_71281_n10073.t169 a_86903_n4245# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2615 VDD.t3194 VDD.t3193 VDD.t3194 VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2616 a_43010_n36322.t3 a_36032_n35156.t5 a_42442_n34390# VDD.t2189 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2617 VDD.t3192 VDD.t3191 VDD.t3192 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2618 a_64243_n5344.t1 a_50751_n19729.t176 a_63683_n5344# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2619 a_71864_6405# a_65486_11614.t14 VDD.t4779 VSS.t423 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2620 a_33249_48695.t13 a_33379_34007.t38 a_33249_34067.t72 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2621 VDD.t154 a_31699_20742.t132 a_33249_48695.t264 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2622 a_93131_n13190# a_71281_n10073.t170 a_92601_n16810# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2623 VDD.t3190 VDD.t3189 VDD.t3190 VDD.t1290 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2624 a_101641_n8770# a_71281_n8397.t185 a_100803_n7865# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2625 a_88271_n13190# a_71281_n10073.t171 a_87433_n13190# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2626 a_31953_n19727.t47 a_31953_n19727.t46 VSS.t83 VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2627 a_53145_n17803# a_50751_n19729.t177 a_54019_n16009# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2628 VSS.t2415 VSS.t2414 VSS.t2415 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2629 VDD.t4907 a_52635_34067.t133 a_52635_48695.t142 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2630 a_71342_n30339.t3 a_65486_n36322.t14 a_73268_n27257# VSS.t155 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2631 VDD.t3188 VDD.t3187 VDD.t3188 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2632 a_33249_48695.t263 a_31699_20742.t133 VDD.t155 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2633 VSS.t2413 VSS.t2412 VSS.t2413 VSS.t733 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2634 VDD.t3186 VDD.t3185 VDD.t3186 VDD.t2464 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2635 a_64243_n16009.t1 a_50751_n19729.t178 a_63683_n16009# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2636 VDD.t3184 VDD.t3183 VDD.t3184 VDD.t979 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2637 a_71281_n10073.t45 a_71281_n10073.t44 VDD.t356 VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2638 VSS.t2411 VSS.t2410 VSS.t2411 VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2639 a_52635_49681.t37 a_35922_19591.t85 OUT.t70 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2640 VDD.t3182 VDD.t3181 VDD.t3182 VDD.t2570 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2641 VDD.t3180 VDD.t3179 VDD.t3180 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2642 VSS.t2409 VSS.t2408 VSS.t2409 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2643 VSS.t2407 VSS.t2406 VSS.t2407 VSS.t1157 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2644 a_45138_22884# a_35922_19591.t86 a_44608_22884# VDD.t405 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X2645 a_100820_10448.t8 a_100820_10448.t7 a_102756_13546# VDD.t322 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2646 VDD.t3178 VDD.t3177 VDD.t3178 VDD.t2160 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2647 VSS.t2405 VSS.t2404 VSS.t2405 VSS.t171 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2648 VSS.t2403 VSS.t2402 VSS.t2403 VSS.t151 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2649 VDD.t3176 VDD.t3175 VDD.t3176 VDD.t2155 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2650 a_31831_n5342.t1 a_83325_n29313.t0 a_83725_n29181# VSS.t288 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2651 VSS.t2401 VSS.t2400 VSS.t2401 VSS.t380 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2652 VDD.t3174 VDD.t3173 VDD.t3174 VDD.t1164 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2653 a_32128_n27257# a_30324_n30399.t1 a_31284_n30339.t1 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2654 VSS.t2399 VSS.t2398 VSS.t2399 VSS.t1104 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2655 VDD.t3172 VDD.t3171 VDD.t3172 VDD.t2447 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2656 a_40053_n3548# a_31953_n19727.t192 a_39531_n3548# VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2657 VDD.t3170 VDD.t3169 VDD.t3170 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2658 VSS.t2397 VSS.t2396 VSS.t2397 VSS.t455 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2659 VDD.t3168 VDD.t3167 VDD.t3168 VDD.t944 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2660 a_99667_n20430# a_71281_n8397.t186 a_98829_n20430# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2661 a_102796_7563# a_100992_4421.t0 a_56895_n16009.t1 VSS.t172 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2662 VSS.t2395 VSS.t2394 VSS.t2395 VSS.t459 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2663 VDD.t3166 VDD.t3165 VDD.t3166 VDD.t2142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2664 a_61515_n36322# a_47991_n29313.t1 a_60677_n36322.t2 VDD.t544 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2665 VSS.t82 a_31953_n19727.t44 a_31953_n19727.t45 VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2666 VDD.t3164 VDD.t3163 VDD.t3164 VDD.t1265 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2667 VSS.t2393 VSS.t2392 VSS.t2393 VSS.t10 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2668 VDD.t3162 VDD.t3161 VDD.t3162 VDD.t60 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2669 a_93131_n3340# a_71281_n10073.t172 a_92601_n4245# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2670 a_73302_12380# a_71496_10388.t17 VSS.t173 VDD.t363 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2671 a_57977_n16009.t1 a_50751_n19729.t179 a_57417_n16009# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2672 VSS.t2391 VSS.t2390 VSS.t2391 VSS.t158 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2673 VSS.t2389 VSS.t2388 VSS.t2389 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2674 VDD.t3160 VDD.t3159 VDD.t3160 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2675 a_111063_n20430# a_71281_n8397.t187 a_110225_n20430# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2676 VSS.t2387 VSS.t2386 VSS.t2387 VSS.t772 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2677 VDD.t3158 VDD.t3157 VDD.t3158 VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2678 a_42047_n13316# a_31953_n19727.t193 a_41487_n12419# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2679 a_100820_10448.t6 a_100820_10448.t5 a_102756_11614# VDD.t322 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2680 a_41487_n3548# a_31953_n19727.t194 a_40965_n3548# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2681 VSS.t2385 VSS.t2384 VSS.t2385 VSS.t452 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2682 a_31699_20742.t26 a_31699_20742.t25 VDD.t33 VDD.t32 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2683 VSS.t2383 VSS.t2382 VSS.t2383 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2684 a_37968_n34390# a_36162_n36382.t9 VSS.t441 VDD.t2127 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2685 a_52585_n13318# a_50751_n19729.t180 a_52063_n14215# VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2686 VSS.t2381 VSS.t2380 VSS.t2381 VSS.t704 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2687 VDD.t156 a_31699_20742.t134 a_35502_25545.t10 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2688 a_65486_n35156.t9 a_65658_n29313.t0 a_67462_n30339# VSS.t378 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2689 a_52635_48695.t141 a_52635_34067.t134 VDD.t4906 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2690 VDD.t157 a_31699_20742.t135 a_33249_48695.t262 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2691 a_36530_n27257# a_30152_n36322.t13 a_36008_n27257.t1 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2692 a_52635_48695.t140 a_52635_34067.t135 VDD.t4905 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2693 a_106501_n21335# a_71281_n8397.t188 a_105933_n21335# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2694 VDD.t3156 VDD.t3155 VDD.t3156 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2695 VSS.t2379 VSS.t2378 VSS.t2379 VSS.t947 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2696 a_52635_49681.t140 a_52635_34067.t136 VDD.t4904 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2697 VSS.t2377 VSS.t2376 VSS.t2377 VSS.t681 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2698 a_33249_35053.t130 a_35502_25545.t52 VSS.t161 VSS.t31 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2699 VSS.t2375 VSS.t2374 VSS.t2375 VSS.t568 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2700 VDD.t3154 VDD.t3153 VDD.t3154 VDD.t1439 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2701 VDD.t3152 VDD.t3151 VDD.t3152 VDD.t532 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2702 a_52635_49681.t139 a_52635_34067.t137 VDD.t4903 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2703 a_44363_n16007.t1 a_45445_n19595.t1 a_66058_n28415# VSS.t377 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2704 VSS.t2373 VSS.t2372 VSS.t2373 VSS.t163 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2705 a_85089_13546# a_83153_10448.t15 VDD.t4786 VDD.t1442 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2706 a_41100_20251# a_35502_24538.t0 a_35502_24538.t1 VSS.t191 nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X2707 VDD.t3150 VDD.t3149 VDD.t3150 VDD.t47 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2708 VDD.t4902 a_52635_34067.t138 a_52635_48695.t139 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2709 VDD.t3148 VDD.t3147 VDD.t3148 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2710 VDD.t3146 VDD.t3145 VDD.t3146 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2711 VDD.t3144 VDD.t3143 VDD.t3144 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2712 a_105933_n6960# a_71281_n8397.t189 a_105365_n6960# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2713 a_32913_n1754# a_31953_n19727.t195 a_32353_n1754# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2714 VSS.t2371 VSS.t2370 VSS.t2371 VSS.t150 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2715 VDD.t3142 VDD.t3141 VDD.t3142 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2716 VSS.t2369 VSS.t2368 VSS.t2369 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2717 a_52635_49681.t38 a_35922_19591.t87 OUT.t69 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2718 VDD.t3140 VDD.t3139 VDD.t3140 VDD.t944 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2719 VDD.t3138 VDD.t3137 VDD.t3138 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2720 a_106501_n1530# a_71281_n8397.t190 a_105933_n1530# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2721 a_113081_n28415# a_112559_n29181.t16 a_106830_n36382.t6 VSS.t410 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2722 VDD.t3136 VDD.t3135 VDD.t3136 VDD.t429 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2723 a_33249_34067.t71 a_33379_34007.t39 a_33249_48695.t335 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2724 VDD.t3134 VDD.t3133 VDD.t3134 VDD.t2399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2725 VDD.t3132 VDD.t3131 VDD.t3132 VDD.t1439 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2726 a_33249_35053.t129 a_35502_25545.t53 VSS.t199 VSS.t16 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2727 a_85089_11614# a_83153_10448.t16 VDD.t4787 VDD.t1442 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2728 VDD.t3130 VDD.t3129 VDD.t3130 VDD.t2099 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2729 a_52635_34067.t60 a_35502_24538.t43 a_33249_34067.t10 VSS.t195 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2730 a_111063_n9675# a_71281_n8397.t191 a_110225_n9675# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2731 VDD.t3128 VDD.t3127 VDD.t3128 VDD.t529 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2732 VDD.t3126 VDD.t3125 VDD.t3126 VDD.t1099 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2733 a_89563_n35156# a_89163_n36382.t12 a_89033_n35156.t1 VDD.t548 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2734 a_33249_48695.t261 a_31699_20742.t136 VDD.t158 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2735 VDD.t3124 VDD.t3123 VDD.t3124 VDD.t1218 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2736 a_104527_n3340# a_71281_n8397.t192 a_103997_n4245# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2737 a_77225_n29181.t0 a_65658_n29313.t1 a_79182_n34390# VDD.t501 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2738 VDD.t3122 VDD.t3121 VDD.t3122 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2739 VDD.t3120 VDD.t3119 VDD.t3120 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2740 VDD.t339 a_71281_n10073.t42 a_71281_n10073.t43 VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2741 VSS.t2367 VSS.t2366 VSS.t2367 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2742 a_111631_n4245# a_71281_n8397.t193 a_111063_n4245# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2743 VSS.t2365 VSS.t2364 VSS.t2365 VSS.t650 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2744 a_52635_34067.t57 a_35502_24538.t44 a_33249_34067.t9 VSS.t192 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2745 VDD.t159 a_31699_20742.t137 a_33249_48695.t260 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2746 a_79182_n36322# a_65658_n29313.t1 a_78344_n36322.t3 VDD.t2382 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2747 VDD.t3118 VDD.t3117 VDD.t3118 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2748 a_67111_n8932# a_50751_n19729.t181 a_66551_n8932# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2749 VSS.t2363 VSS.t2362 VSS.t2363 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2750 a_54019_n14215# a_50751_n19729.t182 a_53497_n14215# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2751 VDD.t3116 VDD.t3115 VDD.t3116 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2752 VSS.t2361 VSS.t2360 VSS.t2361 VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2753 a_71281_n8397.t33 a_71281_n8397.t32 VDD.t448 VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2754 VSS.t2359 VSS.t2358 VSS.t2359 VSS.t306 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2755 VDD.t3114 VDD.t3113 VDD.t3114 VDD.t1112 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2756 VSS.t2357 VSS.t2356 VSS.t2357 VSS.t68 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2757 a_39179_n12419# a_31953_n19727.t196 a_38619_n12419# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2758 VSS.t2355 VSS.t2354 VSS.t2355 VSS.t641 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2759 VSS.t2353 VSS.t2352 VSS.t2353 VSS.t1126 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2760 VDD.t3112 VDD.t3111 VDD.t3112 VDD.t1799 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2761 a_89563_n33224# a_89163_n36382.t13 a_71366_n36322.t2 VDD.t548 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2762 VSS.t2351 VSS.t2350 VSS.t2351 VSS.t217 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2763 VSS.t2349 VSS.t2348 VSS.t2349 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2764 VDD.t3110 VDD.t3109 VDD.t3110 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2765 a_52635_48695.t50 a_35922_19591.t88 a_52635_34067.t33 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2766 VDD.t3108 VDD.t3107 VDD.t3108 VDD.t55 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2767 VSS.t2347 VSS.t2346 VSS.t2347 VSS.t571 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2768 VSS.t2345 VSS.t2344 VSS.t2345 VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2769 a_81735_n2435# a_71281_n10073.t173 a_36032_11614.t0 VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2770 a_99667_n15905# a_71281_n8397.t194 a_98829_n15905# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2771 a_107198_6405# a_100820_11614.t10 VDD.t418 VSS.t182 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2772 VSS.t2343 VSS.t2342 VSS.t2343 VSS.t1064 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2773 a_47819_10448.t10 a_47991_4421.t0 a_49795_5639# VSS.t337 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2774 VDD.t3106 VDD.t3105 VDD.t3106 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2775 OUT.t68 a_35922_19591.t89 a_52635_49681.t39 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2776 VSS.t385 a_77225_n29181.t14 a_77747_n28415# VSS.t384 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2777 VSS.t2341 VSS.t2340 VSS.t2341 VSS.t531 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2778 VDD.t3104 VDD.t3103 VDD.t3104 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2779 a_33249_48695.t336 a_33379_34007.t40 a_33249_34067.t70 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2780 VDD.t3102 VDD.t3101 VDD.t3102 VDD.t680 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2781 a_98829_n2435# a_71281_n8397.t195 VDD.t478 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2782 VSS.t2339 VSS.t2338 VSS.t2339 VSS.t1111 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2783 a_89563_12380# a_89163_10388.t17 a_81205_n14095.t2 VDD.t552 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2784 a_67422_12380# a_65486_10448.t15 VDD.t4749 VDD.t866 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2785 a_111063_n15905# a_71281_n8397.t196 a_110225_n15905# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2786 a_71266_n4019.t2 a_71266_n4019.t0 a_75602_n4019# VDD.t1665 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X2787 a_77776_n36322# a_71366_n35156.t7 a_71496_n36382.t7 VDD.t2344 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2788 VDD.t3100 VDD.t3099 VDD.t3100 VDD.t2079 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2789 VDD.t447 a_71281_n8397.t30 a_71281_n8397.t31 VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2790 a_43010_10448.t0 a_30324_4421.t1 a_42442_12380# VDD.t289 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2791 a_61515_13546# a_47991_4421.t1 a_60677_10448.t5 VDD.t3013 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2792 VDD.t3098 VDD.t3097 VDD.t3098 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2793 VDD.t3096 VDD.t3095 VDD.t3096 VDD.t2076 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2794 a_33249_48695.t46 a_33379_34917.t35 a_33249_35053.t32 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2795 VSS.t2337 VSS.t2336 VSS.t2337 VSS.t334 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2796 VDD.t3094 VDD.t3093 VDD.t3094 VDD.t855 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2797 VDD.t3092 VDD.t3091 VDD.t3092 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2798 VSS.t2335 VSS.t2334 VSS.t2335 VSS.t558 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2799 a_35781_n2651# a_31953_n19727.t197 a_35221_n1754# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2800 a_32913_n18698# a_31953_n19727.t198 a_32353_n17801# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2801 VDD.t3090 VDD.t3089 VDD.t3090 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2802 a_84017_n5150.t0 a_71281_n10073.t174 a_83709_n1530# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2803 VSS.t2333 VSS.t2332 VSS.t2333 VSS.t393 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2804 VDD.t3088 VDD.t3087 VDD.t3088 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2805 VSS.t2331 VSS.t2330 VSS.t2331 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2806 I1N.t1 I1N.t0 a_75585_n8397# VSS.t312 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X2807 a_85129_7563# a_83325_4421.t0 a_50629_n16009.t1 VSS.t309 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2808 VSS.t449 a_106830_n36382.t14 a_107230_n35156# VDD.t845 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2809 VDD.t3086 VDD.t3085 VDD.t3086 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2810 VSS.t2329 VSS.t2328 VSS.t2329 VSS.t944 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2811 VDD.t3084 VDD.t3083 VDD.t3084 VDD.t836 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2812 a_110225_n17715# a_71281_n8397.t197 a_109695_n16810# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2813 a_61515_11614# a_47991_4421.t1 a_60677_10448.t4 VDD.t3013 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2814 VSS.t2327 VSS.t2326 VSS.t2327 VSS.t487 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2815 VDD.t3082 VDD.t3081 VDD.t3082 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2816 VSS.t2325 VSS.t2324 VSS.t2325 VSS.t834 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2817 a_43848_n34390# a_30324_n29313.t2 a_43010_n36322.t3 VDD.t2061 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2818 a_30152_10448.t7 a_30152_10448.t6 a_32088_13546# VDD.t305 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2819 a_110225_n15000# a_71281_n8397.t198 a_109695_n15905# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2820 a_53675_7563.t1 a_53829_10388.t13 a_54229_13546# VDD.t1405 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2821 VSS.t2323 VSS.t2322 VSS.t2323 VSS.t609 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2822 VDD.t3080 VDD.t3079 VDD.t3080 VDD.t813 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2823 a_35502_24538.t16 a_31699_20742.t138 VDD.t160 VDD.t20 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2824 a_33249_34067.t69 a_33379_34007.t41 a_33249_48695.t337 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2825 a_31953_n19727.t43 a_31953_n19727.t42 VSS.t81 VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2826 a_89009_7563.t0 a_83153_11614.t18 a_90935_4481# VSS.t392 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2827 a_93969_n13190# a_71281_n10073.t175 a_93131_n13190# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2828 a_78344_10448.t3 a_65658_4421.t2 a_77776_10448# VDD.t3570 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2829 a_53699_13546.t0 a_53829_10388.t14 a_55635_10448# VDD.t3747 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2830 a_36008_n30339.t2 a_36162_n36382.t10 a_36562_n36322# VDD.t2302 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2831 VSS.t2321 VSS.t2320 VSS.t2321 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2832 VDD.t3078 VDD.t3077 VDD.t3078 VDD.t398 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2833 VDD.t3076 VDD.t3075 VDD.t3076 VDD.t823 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2834 a_48391_5639# a_47991_5507.t1 a_47819_11614.t7 VSS.t339 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2835 VDD.t3074 VDD.t3073 VDD.t3074 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2836 a_52635_48695.t138 a_52635_34067.t139 VDD.t4901 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2837 a_106676_n27257.t2 a_106830_n36382.t15 a_107230_n33224# VDD.t845 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2838 VDD.t3072 VDD.t3071 VDD.t3072 VDD.t78 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2839 VSS.t2319 VSS.t2318 VSS.t2319 VSS.t495 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2840 a_41487_n13316# a_31953_n19727.t199 a_40965_n14213# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2841 VDD.t161 a_31699_20742.t139 a_33249_48695.t259 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2842 VDD.t3070 VDD.t3069 VDD.t3070 VDD.t836 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2843 VSS.t2317 VSS.t2316 VSS.t2317 VSS.t522 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2844 a_38619_n6239# a_31953_n19727.t200 a_38097_n7136# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2845 VSS.t301 a_112559_4481.t19 a_113081_4481# VSS.t294 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2846 VSS.t2315 VSS.t2314 VSS.t2315 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2847 VDD.t3068 VDD.t3067 VDD.t3068 VDD.t935 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2848 VDD.t3066 VDD.t3065 VDD.t3066 VDD.t810 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2849 a_89407_n14095# a_71281_n10073.t176 a_88839_n14095# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2850 VDD.t3064 VDD.t3063 VDD.t3064 VDD.t1155 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2851 VSS.t417 a_53829_10388.t15 a_54229_11614# VDD.t1405 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2852 a_30152_10448.t9 a_30152_10448.t8 a_32088_11614# VDD.t305 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2853 VDD.t3062 VDD.t3061 VDD.t3062 VDD.t25 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2854 VDD.t3060 VDD.t3059 VDD.t3060 VDD.t2299 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X2855 a_52635_49681.t138 a_52635_34067.t140 VDD.t4900 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2856 VDD.t162 a_31699_20742.t140 a_33249_48695.t258 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2857 VDD.t4899 a_52635_34067.t141 a_52635_48695.t137 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2858 a_47753_n5342# a_31953_n19727.t201 a_46879_n7136# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2859 VDD.t3058 VDD.t3057 VDD.t3058 VDD.t823 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2860 a_100803_n14095# a_71281_n8397.t199 a_100235_n14095# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2861 VDD.t3056 VDD.t3055 VDD.t3056 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2862 VSS.t2313 VSS.t2312 VSS.t2313 VSS.t285 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2863 a_48313_n19595# a_31953_n19727.t202 a_47753_n19595# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2864 a_35502_24538.t15 a_31699_20742.t141 VDD.t163 VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2865 VSS.t2311 VSS.t2310 VSS.t2311 VSS.t220 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2866 VSS.t2309 VSS.t2308 VSS.t2309 VSS.t558 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2867 a_33249_48695.t47 a_33379_34917.t36 a_33249_35053.t33 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2868 a_71496_10388.t2 a_77225_4481.t16 a_79151_4481# VSS.t318 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2869 a_71496_n36382.t3 a_77225_n29181.t15 a_79151_n27257# VSS.t380 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2870 VDD.t3054 VDD.t3053 VDD.t3054 VDD.t2254 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2871 VSS.t51 a_35502_25545.t54 a_33249_35053.t128 VSS.t27 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2872 a_93131_n2435# a_71281_n10073.t177 a_71366_11614.t0 VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2873 a_89009_n30339.t1 a_83153_n36322.t14 a_90935_n27257# VSS.t455 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2874 VDD.t3052 VDD.t3051 VDD.t3052 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2875 VSS.t2307 VSS.t2306 VSS.t2307 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2876 VDD.t31 a_31699_20742.t23 a_31699_20742.t24 VDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2877 VDD.t3050 VDD.t3049 VDD.t3050 VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2878 VSS.t2305 VSS.t2304 VSS.t2305 VSS.t394 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2879 VDD.t3048 VDD.t3047 VDD.t3048 VDD.t810 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2880 a_95443_n35156# a_83325_n29313.t1 a_94892_n29181.t1 VDD.t795 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2881 a_60845_n15112# a_50751_n19729.t183 a_60285_n15112# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2882 VSS.t2303 VSS.t2302 VSS.t2303 VSS.t495 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2883 a_63683_n8035# a_50751_n19729.t184 a_63161_n8932# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2884 VSS.t2301 VSS.t2300 VSS.t2301 VSS.t33 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2885 a_106676_n27257.t1 a_100820_n36322.t13 a_108602_n30339# VSS.t333 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2886 VSS.t2299 VSS.t2298 VSS.t2299 VSS.t498 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2887 a_51711_n16906# a_50751_n19729.t185 a_51151_n16906# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2888 a_44885_n13316# a_31953_n19727.t203 a_44363_n13316# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2889 a_65677_n8932# a_50751_n19729.t186 a_65117_n8035# VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2890 VDD.t3046 VDD.t3045 VDD.t3046 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2891 VDD.t3044 VDD.t3043 VDD.t3044 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2892 VDD.t3042 VDD.t3041 VDD.t3042 VDD.t1322 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2893 VDD.t3040 VDD.t3039 VDD.t3040 VDD.t303 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2894 VDD.t3038 VDD.t3037 VDD.t3038 VDD.t2349 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2895 VSS.t2297 VSS.t2296 VSS.t2297 VSS.t63 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2896 VSS.t2295 VSS.t2294 VSS.t2295 VSS.t478 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2897 VSS.t2293 VSS.t2292 VSS.t2293 VSS.t647 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2898 a_52635_48695.t49 a_35922_19591.t90 a_52635_34067.t34 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2899 VSS.t2291 VSS.t2290 VSS.t2291 VSS.t1077 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X2900 a_95413_n5150.t0 a_71281_n10073.t178 a_95105_n1530# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2901 VDD.t3036 VDD.t3035 VDD.t3036 VDD.t1349 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2902 a_39179_n8930.t1 a_100820_n36322.t14 a_107198_n28415# VSS.t336 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2903 a_110225_n20430# a_71281_n8397.t200 a_71366_n35156.t0 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2904 a_33249_48695.t48 a_33379_34917.t37 a_33249_35053.t34 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2905 a_95443_n33224# a_83325_n29313.t1 a_94892_n29181.t1 VDD.t795 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2906 VDD.t3034 VDD.t3033 VDD.t3034 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2907 a_60845_n7138# a_50751_n19729.t187 a_60285_n7138# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2908 VSS.t2289 VSS.t2288 VSS.t2289 VSS.t160 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2909 VSS.t2287 VSS.t2286 VSS.t2287 VSS.t305 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2910 a_71366_13546.t2 a_71496_10388.t18 a_73302_10448# VDD.t352 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2911 VDD.t3032 VDD.t3031 VDD.t3032 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2912 VSS.t2285 VSS.t2284 VSS.t2285 VSS.t39 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2913 VSS.t2283 VSS.t2282 VSS.t2283 VSS.t192 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2914 a_33249_48695.t257 a_31699_20742.t142 VDD.t164 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2915 a_54579_n15112# a_50751_n19729.t188 a_54019_n15112# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2916 a_52635_48695.t136 a_52635_34067.t142 VDD.t4898 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2917 a_106830_n36382.t0 a_103997_n8770.t7 a_114516_n35156# VDD.t538 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2918 VDD.t3030 VDD.t3029 VDD.t3030 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2919 VSS.t2281 VSS.t2280 VSS.t2281 VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2920 VDD.t3028 VDD.t3027 VDD.t3028 VDD.t1322 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2921 a_93969_n3340# a_71281_n10073.t179 a_93131_n3340# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2922 VDD.t3026 VDD.t3025 VDD.t3026 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2923 VDD.t3024 VDD.t3023 VDD.t3024 VDD.t560 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2924 a_64243_n16906# a_50751_n19729.t189 a_63683_n15112# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2925 VSS.t2279 VSS.t2278 VSS.t2279 VSS.t891 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2926 VSS.t2277 VSS.t2276 VSS.t2277 VSS.t633 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2927 VDD.t3022 VDD.t3021 VDD.t3022 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2928 VSS.t2275 VSS.t2274 VSS.t2275 VSS.t352 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2929 a_33249_48695.t49 a_33379_34917.t38 a_33249_35053.t35 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2930 a_33249_34067.t129 a_35502_25545.t55 VSS.t23 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2931 VDD.t446 a_71281_n8397.t28 a_71281_n8397.t29 VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2932 a_37934_n28415# a_30152_n36322.t14 a_30324_n30399.t1 VSS.t282 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2933 a_104527_n2435# a_71281_n8397.t201 VDD.t479 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2934 a_82573_n4245# a_71281_n10073.t180 a_81735_n4245# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2935 a_35221_n15110# a_31953_n19727.t204 a_34699_n16904# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2936 a_106830_n36382.t3 a_103997_n8770.t8 a_114516_n33224# VDD.t538 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2937 VSS.t3640 a_94892_4481.t16 a_95414_6405# VSS.t1037 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2938 a_111631_n15000# a_71281_n8397.t202 a_111063_n15000# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2939 a_73268_7563# a_65486_11614.t15 a_65658_4421.t0 VSS.t421 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2940 VDD.t3020 VDD.t3019 VDD.t3020 VDD.t755 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2941 VDD.t3018 VDD.t3017 VDD.t3018 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2942 a_40053_n2651# a_31953_n19727.t205 a_39531_n3548# VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2943 a_33249_48695.t338 a_33379_34007.t42 a_33249_34067.t68 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2944 VSS.t2273 VSS.t2272 VSS.t2273 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2945 a_67111_n19597# a_50751_n19729.t190 a_66551_n18700# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2946 VSS.t2271 VSS.t2270 VSS.t2271 VSS.t537 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2947 a_106809_n5150.t1 a_100992_n29313.t2 a_113110_n35156# VDD.t537 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2948 a_99667_n4245# a_71281_n8397.t203 a_98829_n4245# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2949 VDD.t165 a_31699_20742.t143 a_35502_25545.t11 VDD.t34 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2950 a_52635_34067.t35 a_35922_19591.t91 a_52635_48695.t48 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2951 VDD.t3016 VDD.t3015 VDD.t3016 VDD.t2299 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X2952 a_46319_n14213# a_31953_n19727.t206 a_45797_n14213# VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2953 VDD.t3014 VDD.t3012 VDD.t3014 VDD.t3013 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2954 a_57977_n16906# a_50751_n19729.t191 a_57417_n15112# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2955 VDD.t3011 VDD.t3010 VDD.t3011 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2956 VDD.t3009 VDD.t3008 VDD.t3009 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2957 a_41487_n2651# a_31953_n19727.t207 a_40965_n3548# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2958 VSS.t2269 VSS.t2268 VSS.t2269 VSS.t612 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2959 VSS.t2267 VSS.t2266 VSS.t2267 VSS.t1025 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2960 VDD.t3007 VDD.t3006 VDD.t3007 VDD.t1142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2961 VDD.t378 a_71281_n10073.t181 a_89407_n9675# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2962 a_35221_n1754# a_31953_n19727.t208 a_32913_n1754# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2963 VDD.t3005 VDD.t3004 VDD.t3005 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2964 VSS.t2265 VSS.t2264 VSS.t2265 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2965 a_43010_n36322.t2 a_36032_n35156.t6 a_42442_n36322# VDD.t2189 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2966 a_108636_12380# a_106830_10388.t16 VSS.t315 VDD.t520 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2967 a_52585_n12421# a_50751_n19729.t192 a_51711_n16009.t0 VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2968 a_57977_n5344.t1 a_50751_n19729.t193 a_57417_n5344# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2969 a_107230_10448# a_106830_10388.t17 a_89033_13546.t0 VDD.t522 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2970 VDD.t3003 VDD.t3002 VDD.t3003 VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2971 a_106809_n5150.t1 a_100992_n29313.t2 a_113110_n33224# VDD.t537 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2972 a_38619_n18698# a_31953_n19727.t209 a_38097_n19595# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2973 VDD.t3001 VDD.t3000 VDD.t3001 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2974 a_37934_5639# a_30152_11614.t10 a_30324_5507.t1 VSS.t282 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2975 VDD.t2999 VDD.t2998 VDD.t2999 VDD.t720 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2976 a_33249_34067.t67 a_33379_34007.t43 a_33249_48695.t339 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2977 a_30152_n36322.t1 a_30324_n30399.t1 a_32128_n29181# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2978 VDD.t4897 a_52635_34067.t143 a_52635_48695.t135 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2979 VDD.t2997 VDD.t2996 VDD.t2997 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2980 VSS.t2263 VSS.t2262 VSS.t2263 VSS.t859 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2981 a_51151_n4447# a_50751_n19729.t194 a_50629_n4447# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2982 VDD.t2995 VDD.t2994 VDD.t2995 VDD.t1086 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2983 VDD.t2993 VDD.t2992 VDD.t2993 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2984 VSS.t2261 VSS.t2260 VSS.t2261 VSS.t397 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2985 a_49755_n35156# a_47819_n35156.t18 VDD.t4796 VDD.t707 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2986 VSS.t372 a_41891_n29181.t17 a_42413_n30339# VSS.t166 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2987 VSS.t32 a_35502_25545.t56 a_33249_35053.t127 VSS.t31 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2988 VDD.t2991 VDD.t2990 VDD.t2991 VDD.t1142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2989 a_44885_n8930# a_31953_n19727.t210 a_44363_n8930# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2990 VDD.t343 a_71281_n10073.t40 a_71281_n10073.t41 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2991 VDD.t2989 VDD.t2988 VDD.t2989 VDD.t1917 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2992 a_50751_n19729.t41 a_50751_n19729.t40 VSS.t239 VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2993 VSS.t3645 a_112559_n29181.t17 a_113081_n29181# VSS.t411 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2994 VSS.t2259 VSS.t2258 VSS.t2259 VSS.t795 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2995 VDD.t2987 VDD.t2986 VDD.t2987 VDD.t1262 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2996 a_88271_n6960# a_71281_n10073.t182 a_87433_n6960# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2997 a_33249_35053.t36 a_33379_34917.t39 a_33249_48695.t50 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2998 a_84547_n20430# a_71281_n10073.t183 a_83709_n19525# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2999 VSS.t2257 VSS.t2256 VSS.t2257 VSS.t106 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3000 a_46879_n8930# a_31953_n19727.t211 a_46319_n8930# VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3001 VDD.t4896 a_52635_34067.t144 a_52635_48695.t134 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3002 VDD.t2985 VDD.t2984 VDD.t2985 VDD.t2160 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3003 a_87433_n13190# a_71281_n10073.t184 a_86903_n16810# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3004 VDD.t2983 VDD.t2982 VDD.t2983 VDD.t2542 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3005 VDD.t2981 VDD.t2980 VDD.t2981 VDD.t2155 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3006 VDD.t2979 VDD.t2978 VDD.t2979 VDD.t401 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3007 VSS.t2255 VSS.t2254 VSS.t2255 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3008 VDD.t2977 VDD.t2976 VDD.t2977 VDD.t720 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3009 VSS.t2253 VSS.t2252 VSS.t2253 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3010 VSS.t2251 VSS.t2250 VSS.t2251 VSS.t261 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3011 a_95414_6405# a_94892_4481.t6 a_94892_4481.t7 VSS.t998 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3012 a_110225_n15905# a_71281_n8397.t204 a_109695_n15905# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3013 a_107230_n34390# a_106830_n36382.t16 a_103997_n8770.t3 VDD.t1904 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3014 VDD.t2975 VDD.t2974 VDD.t2975 VDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3015 VSS.t2249 VSS.t2248 VSS.t2249 VSS.t490 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3016 VSS.t2247 VSS.t2246 VSS.t2247 VSS.t475 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3017 VSS.t358 a_94892_n29181.t14 a_95414_n28415# VSS.t357 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3018 a_49755_n33224# a_47819_n35156.t19 VDD.t4797 VDD.t707 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3019 VDD.t2973 VDD.t2972 VDD.t2973 VDD.t363 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3020 a_111631_n20430# a_71281_n8397.t205 a_111063_n20430# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3021 VDD.t2971 VDD.t2970 VDD.t2971 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3022 VSS.t2245 VSS.t2244 VSS.t2245 VSS.t591 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3023 VDD.t2969 VDD.t2968 VDD.t2969 VDD.t2142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3024 VSS.t2243 VSS.t2242 VSS.t2243 VSS.t102 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3025 VSS.t2241 VSS.t2240 VSS.t2241 VSS.t944 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3026 VDD.t2967 VDD.t2966 VDD.t2967 VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3027 VDD.t2965 VDD.t2964 VDD.t2965 VDD.t1262 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3028 VSS.t17 a_35502_25545.t57 a_33249_35053.t126 VSS.t16 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3029 VSS.t2239 VSS.t2238 VSS.t2239 VSS.t588 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3030 VSS.t2237 VSS.t2236 VSS.t2237 VSS.t576 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3031 a_36032_n35156.t1 a_36162_n36382.t11 a_37968_n34390# VDD.t1893 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3032 VDD.t2963 VDD.t2962 VDD.t2963 VDD.t401 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3033 VSS.t2235 VSS.t2234 VSS.t2235 VSS.t638 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3034 VSS.t2233 VSS.t2232 VSS.t2233 VSS.t41 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X3035 VSS.t2231 VSS.t2230 VSS.t2231 VSS.t217 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3036 a_43848_12380# a_36032_11614.t9 a_43010_10448.t2 VDD.t290 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3037 VSS.t2229 VSS.t2228 VSS.t2229 VSS.t264 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3038 VDD.t2961 VDD.t2960 VDD.t2961 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3039 a_31953_n19727.t41 a_31953_n19727.t40 VSS.t80 VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3040 a_37968_n36322# a_36162_n36382.t12 a_36008_n27257.t3 VDD.t2127 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3041 VDD.t166 a_31699_20742.t144 a_35502_24538.t14 VDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3042 a_65117_n13318# a_50751_n19729.t195 a_64595_n14215# VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3043 VSS.t2227 VSS.t2226 VSS.t2227 VSS.t1821 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X3044 VDD.t167 a_31699_20742.t145 a_33249_48695.t256 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3045 VDD.t2959 VDD.t2958 VDD.t2959 VDD.t1884 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3046 a_52635_49681.t40 a_35922_19591.t92 OUT.t67 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3047 VSS.t2225 VSS.t2224 VSS.t2225 VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3048 a_63683_n3550# a_50751_n19729.t196 a_63161_n4447# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3049 VSS.t2223 VSS.t2222 VSS.t2223 VSS.t495 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3050 VDD.t480 a_71281_n8397.t206 a_100803_n1530# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3051 VDD.t168 a_31699_20742.t146 a_33249_48695.t255 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3052 a_40053_n17801# a_31953_n19727.t212 a_39531_n18698# VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3053 a_33249_34067.t66 a_33379_34007.t44 a_33249_48695.t340 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3054 VDD.t4895 a_52635_34067.t145 a_52635_49681.t137 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3055 VSS.t2221 VSS.t2220 VSS.t2221 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3056 a_59411_n13318# a_50751_n19729.t197 a_58851_n13318# VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3057 a_65117_n8035# a_50751_n19729.t198 a_64595_n8035# VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3058 VDD.t2957 VDD.t2956 VDD.t2957 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3059 VDD.t2955 VDD.t2954 VDD.t2955 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3060 a_36162_n36382.t0 a_41891_n29181.t18 a_43817_n29181# VSS.t168 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3061 VDD.t2953 VDD.t2952 VDD.t2953 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3062 a_65677_n3550# a_50751_n19729.t199 a_65117_n3550# VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3063 VDD.t2951 VDD.t2950 VDD.t2951 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3064 VSS.t2219 VSS.t2218 VSS.t2219 VSS.t687 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3065 VDD.t2949 VDD.t2948 VDD.t2949 VDD.t1042 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3066 VSS.t2217 VSS.t2216 VSS.t2217 VSS.t760 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3067 a_47819_10448.t1 a_47819_10448.t0 a_49755_13546# VDD.t496 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3068 VDD.t2947 VDD.t2946 VDD.t2947 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3069 VSS.t2215 VSS.t2214 VSS.t2215 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3070 a_50751_n19729.t72 a_71266_n4019.t0 a_75602_n4978# VDD.t1665 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3071 VDD.t2945 VDD.t2944 VDD.t2945 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3072 VDD.t2943 VDD.t2942 VDD.t2943 VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3073 VDD.t2941 VDD.t2940 VDD.t2941 VDD.t6 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3074 VDD.t2939 VDD.t2938 VDD.t2939 VDD.t429 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3075 VDD.t355 a_71281_n10073.t38 a_71281_n10073.t39 VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3076 VDD.t2937 VDD.t2936 VDD.t2937 VDD.t289 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3077 VDD.t2935 VDD.t2934 VDD.t2935 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3078 VDD.t2933 VDD.t2932 VDD.t2933 VDD.t648 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3079 VDD.t2931 VDD.t2930 VDD.t2931 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3080 VDD.t2929 VDD.t2928 VDD.t2929 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3081 a_83153_11614.t5 a_83153_10448.t17 a_85089_12380# VDD.t643 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3082 VDD.t2927 VDD.t2926 VDD.t2927 VDD.t1206 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3083 VSS.t2213 VSS.t2212 VSS.t2213 VSS.t814 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3084 VDD.t4788 a_83153_10448.t18 a_83683_10448# VDD.t3354 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3085 VDD.t2925 VDD.t2923 VDD.t2925 VDD.t2924 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3086 VDD.t2922 VDD.t2920 VDD.t2922 VDD.t2921 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3087 VDD.t2919 VDD.t2918 VDD.t2919 VDD.t2099 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3088 a_71281_n8397.t27 a_71281_n8397.t26 VDD.t445 VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3089 VDD.t2917 VDD.t2916 VDD.t2917 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3090 a_47819_10448.t3 a_47819_10448.t2 a_49755_11614# VDD.t496 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3091 VDD.t2915 VDD.t2914 VDD.t2915 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3092 VDD.t2913 VDD.t2912 VDD.t2913 VDD.t630 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3093 VSS.t2211 VSS.t2210 VSS.t2211 VSS.t834 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3094 a_107339_n8770# a_71281_n8397.t207 a_106501_n8770# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3095 a_77225_n29181.t1 a_65658_n29313.t1 a_79182_n36322# VDD.t501 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3096 VDD.t169 a_31699_20742.t147 a_33249_48695.t254 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3097 a_45445_n19595.t0 a_31953_n19727.t213 a_44885_n19595# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3098 a_106830_10388.t6 a_86903_n14095.t7 a_114516_10448# VDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3099 a_30682_n35156# a_30152_n35156.t10 a_30152_n35156.t11 VDD.t622 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3100 a_34347_n14213# a_31953_n19727.t214 a_35221_n16007# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3101 VDD.t4753 a_83153_n35156.t11 a_83683_n34390# VDD.t1850 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3102 a_58851_n8932# a_50751_n19729.t200 VSS.t271 VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3103 VSS.t38 a_35502_25545.t58 a_33249_34067.t128 VSS.t37 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3104 OUT.t66 a_35922_19591.t93 a_52635_49681.t41 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3105 VDD.t2911 VDD.t2910 VDD.t2911 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3106 VSS.t2209 VSS.t2208 VSS.t2209 VSS.t653 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3107 VDD.t2909 VDD.t2908 VDD.t2909 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3108 VDD.t2907 VDD.t2906 VDD.t2907 VDD.t1206 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3109 a_93969_n2435# a_71281_n10073.t185 a_93131_n2435# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3110 VSS.t2207 VSS.t2206 VSS.t2207 VSS.t528 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3111 a_99667_n14095# a_71281_n8397.t208 a_98829_n14095# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3112 a_66551_n19597# a_50751_n19729.t201 a_64243_n19597# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3113 VDD.t2905 VDD.t2904 VDD.t2905 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3114 a_55601_n27257# a_47819_n36322.t14 a_47991_n29313.t0 VSS.t305 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3115 VDD.t2903 VDD.t2902 VDD.t2903 VDD.t603 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3116 VDD.t2901 VDD.t2900 VDD.t2901 VDD.t630 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3117 VDD.t2899 VDD.t2898 VDD.t2899 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3118 a_111063_n14095# a_71281_n8397.t209 a_110225_n14095# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3119 VSS.t2205 VSS.t2204 VSS.t2205 VSS.t1426 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3120 VSS.t2203 VSS.t2202 VSS.t2203 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3121 a_30682_n33224# a_30152_n35156.t8 a_30152_n35156.t9 VDD.t622 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3122 a_113037_n6055# a_71281_n8397.t210 a_112507_n6055.t1 VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3123 a_55635_n35156# a_53829_n36382.t19 VSS.t391 VDD.t367 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3124 VDD.t2897 VDD.t2896 VDD.t2897 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3125 VSS.t402 a_59558_4481.t12 a_60080_5639# VSS.t401 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3126 a_111631_n15905# a_71281_n8397.t211 a_111063_n15905# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3127 a_31699_17542# I1U.t3 a_30377_18342# VSS.t349 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X3128 VSS.t2201 VSS.t2200 VSS.t2201 VSS.t891 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3129 a_38619_n5342# a_31953_n19727.t215 a_38097_n5342.t0 VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3130 a_64243_n1756.t1 a_65486_11614.t16 a_71864_6405# VSS.t424 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3131 a_33249_48695.t341 a_33379_34007.t45 a_33249_34067.t65 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3132 VDD.t2895 VDD.t2894 VDD.t2895 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3133 VDD.t2893 VDD.t2892 VDD.t2893 VDD.t1824 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3134 VSS.t2199 VSS.t2198 VSS.t2199 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3135 a_83153_10448.t3 a_83325_4421.t0 a_85129_5639# VSS.t308 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3136 VSS.t2197 VSS.t2196 VSS.t2197 VSS.t908 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3137 VDD.t2891 VDD.t2890 VDD.t2891 VDD.t1821 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3138 VSS.t238 a_50751_n19729.t38 a_50751_n19729.t39 VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3139 VDD.t2889 VDD.t2888 VDD.t2889 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3140 a_95413_n16810.t0 a_71281_n10073.t186 a_95105_n13190# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3141 VDD.t2887 VDD.t2886 VDD.t2887 VDD.t322 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3142 VCM.t3 a_33379_34007.t1 cap_mim_2f0_m4m5_noshield c_width=9.8u c_length=9.8u
X3143 VDD.t2885 VDD.t2884 VDD.t2885 VDD.t852 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3144 VDD.t2883 VDD.t2882 VDD.t2883 VDD.t2079 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3145 VDD.t2881 VDD.t2880 VDD.t2881 VDD.t603 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3146 a_52635_48695.t47 a_35922_19591.t94 a_52635_34067.t36 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3147 VDD.t2879 VDD.t2878 VDD.t2879 VDD.t2076 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3148 a_65486_10448.t5 a_65486_10448.t4 a_67422_13546# VDD.t1378 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3149 a_60109_n35156# a_47991_n29313.t1 a_59558_n29181.t0 VDD.t543 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3150 VDD.t170 a_31699_20742.t148 a_33249_48695.t253 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3151 VSS.t2195 VSS.t2194 VSS.t2195 VSS.t332 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3152 a_35502_24538.t13 a_31699_20742.t149 VDD.t171 VDD.t20 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3153 a_113110_n34390# a_103997_n8770.t9 a_106830_n36382.t2 VDD.t535 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3154 a_36562_10448# a_36162_10388.t17 a_33379_34917.t1 VDD.t3423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3155 a_33249_34067.t64 a_33379_34007.t46 a_33249_48695.t342 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3156 VDD.t4894 a_52635_34067.t146 a_52635_49681.t136 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3157 a_55635_n33224# a_53829_n36382.t20 a_53675_n30339.t1 VDD.t367 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3158 VDD.t2877 VDD.t2876 VDD.t2877 VDD.t404 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3159 VSS.t2193 VSS.t2192 VSS.t2193 VSS.t772 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3160 a_35502_25545.t12 a_31699_20742.t150 VDD.t172 VDD.t32 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3161 a_82573_n18620# a_71281_n10073.t187 a_81735_n18620# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3162 a_111063_n3340# a_71281_n8397.t212 a_110225_n3340# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3163 a_33249_35053.t125 a_35502_25545.t59 VSS.t28 VSS.t27 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3164 VDD.t2875 VDD.t2874 VDD.t2875 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3165 VSS.t2191 VSS.t2190 VSS.t2191 VSS.t687 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3166 a_52635_48695.t133 a_52635_34067.t147 VDD.t4893 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3167 VSS.t2189 VSS.t2188 VSS.t2189 VSS.t721 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3168 VSS.t2187 VSS.t2186 VSS.t2187 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3169 a_41891_n29181.t2 a_30324_n29313.t2 a_43848_n34390# VDD.t1796 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3170 VDD.t2873 VDD.t2872 VDD.t2873 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3171 VDD.t2871 VDD.t2870 VDD.t2871 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3172 VDD.t2869 VDD.t2868 VDD.t2869 VDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3173 a_46319_n8930# a_31953_n19727.t216 a_45445_n5342.t0 VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3174 a_65486_10448.t3 a_65486_10448.t2 a_67422_11614# VDD.t1378 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3175 a_60109_n33224# a_47991_n29313.t1 a_59558_n29181.t0 VDD.t543 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3176 a_94537_n13190# a_71281_n10073.t188 a_93969_n13190# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3177 VSS.t2185 VSS.t2184 VSS.t2185 VSS.t292 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3178 VSS.t2183 VSS.t2182 VSS.t2183 VSS.t166 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3179 a_43848_n36322# a_30324_n29313.t2 a_43010_n36322.t2 VDD.t2061 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3180 VDD.t2867 VDD.t2866 VDD.t2867 VDD.t1747 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3181 VDD.t2865 VDD.t2864 VDD.t2865 VDD.t404 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3182 VDD.t2863 VDD.t2862 VDD.t2863 VDD.t1780 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3183 a_52635_34067.t29 a_35922_19591.t95 a_52635_48695.t46 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3184 VDD.t2861 VDD.t2860 VDD.t2861 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3185 VSS.t2181 VSS.t2180 VSS.t2181 VSS.t154 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3186 VSS.t2179 VSS.t2178 VSS.t2179 VSS.t377 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3187 VSS.t2177 VSS.t2176 VSS.t2177 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3188 a_33249_34067.t63 a_33379_34007.t47 a_33249_48695.t343 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3189 VDD.t2859 VDD.t2858 VDD.t2859 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3190 VDD.t2857 VDD.t2856 VDD.t2857 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3191 a_114485_7563# a_112559_4481.t20 VSS.t302 VSS.t297 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3192 VSS.t2175 VSS.t2174 VSS.t2175 VSS.t1385 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3193 VSS.t2173 VSS.t2172 VSS.t2173 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3194 a_60845_n7138# a_50751_n19729.t202 a_60285_n6241# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3195 a_33249_48695.t51 a_33379_34917.t40 a_33249_35053.t37 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3196 a_47819_n35156.t1 a_47991_n29313.t0 a_49795_n30339# VSS.t337 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3197 VDD.t173 a_31699_20742.t151 a_33249_48695.t252 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3198 a_52635_48695.t132 a_52635_34067.t148 VDD.t4892 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3199 VDD.t2855 VDD.t2854 VDD.t2855 VDD.t979 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3200 a_65677_n14215# a_50751_n19729.t203 a_65117_n14215# VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3201 a_51151_n19597# a_50751_n19729.t204 a_50629_n19597# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3202 VDD.t2853 VDD.t2852 VDD.t2853 VDD.t120 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3203 a_51711_n8035# a_50751_n19729.t205 a_51151_n8035# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3204 VDD.t4891 a_52635_34067.t149 a_52635_49681.t135 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3205 VSS.t2171 VSS.t2170 VSS.t2171 VSS.t410 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3206 VDD.t2851 VDD.t2850 VDD.t2851 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3207 a_89163_10388.t4 a_81205_n14095.t4 a_96849_10448# VDD.t500 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3208 VSS.t2169 VSS.t2168 VSS.t2169 VSS.t690 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3209 VDD.t2849 VDD.t2848 VDD.t2849 VDD.t798 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3210 a_54229_12380# a_53829_10388.t16 a_53699_11614.t2 VDD.t3678 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3211 VSS.t2167 VSS.t2166 VSS.t2167 VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3212 VDD.t2847 VDD.t2846 VDD.t2847 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3213 a_33249_48695.t251 a_31699_20742.t152 VDD.t174 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3214 VSS.t2165 VSS.t2164 VSS.t2165 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3215 VDD.t4890 a_52635_34067.t150 a_52635_48695.t131 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3216 VDD.t2845 VDD.t2844 VDD.t2845 VDD.t962 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X3217 VDD.t2843 VDD.t2842 VDD.t2843 VDD.t49 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3218 VSS.t2163 VSS.t2162 VSS.t2163 VSS.t162 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3219 VSS.t2161 VSS.t2160 VSS.t2161 VSS.t676 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3220 VSS.t2159 VSS.t2158 VSS.t2159 VSS.t490 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3221 a_60285_n5344# a_50751_n19729.t206 a_59411_n3550# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3222 VDD.t2841 VDD.t2840 VDD.t2841 VDD.t402 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X3223 VSS.t2157 VSS.t2156 VSS.t2157 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3224 a_65117_n3550# a_50751_n19729.t207 a_64595_n3550# VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3225 VDD.t2839 VDD.t2838 VDD.t2839 VDD.t120 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3226 a_35221_n14213# a_31953_n19727.t217 a_34699_n14213# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3227 VDD.t2837 VDD.t2836 VDD.t2837 VDD.t2464 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3228 VSS.t2155 VSS.t2154 VSS.t2155 VSS.t293 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3229 a_34347_n19595# a_31953_n19727.t218 a_33787_n18698# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3230 VDD.t2835 VDD.t2834 VDD.t2835 VDD.t1419 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3231 VSS.t2153 VSS.t2152 VSS.t2153 VSS.t1244 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X3232 VDD.t2833 VDD.t2832 VDD.t2833 VDD.t55 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3233 VDD.t2831 VDD.t2830 VDD.t2831 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3234 a_101392_n30339# a_39179_n8930.t1 a_100820_n36322.t4 VSS.t331 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3235 VSS.t2151 VSS.t2150 VSS.t2151 VSS.t378 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3236 a_71281_n8397.t25 a_71281_n8397.t24 VDD.t443 VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3237 VSS.t2149 VSS.t2148 VSS.t2149 VSS.t283 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3238 VDD.t2829 VDD.t2828 VDD.t2829 VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3239 VSS.t49 a_35502_25545.t60 a_33249_34067.t127 VSS.t25 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3240 a_52635_48695.t45 a_35922_19591.t96 a_52635_34067.t37 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3241 VSS.t2147 VSS.t2146 VSS.t2147 VSS.t160 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3242 VSS.t2145 VSS.t2144 VSS.t2145 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3243 VDD.t175 a_31699_20742.t153 a_35502_24538.t12 VDD.t16 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3244 VDD.t176 a_31699_20742.t154 a_33249_48695.t250 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3245 VSS.t2143 VSS.t2142 VSS.t2143 VSS.t319 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3246 VSS.t2141 VSS.t2140 VSS.t2141 VSS.t1360 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3247 a_67462_7563# a_65658_4421.t0 a_63161_n5344.t1 VSS.t289 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3248 VDD.t2827 VDD.t2826 VDD.t2827 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3249 a_52585_n7138# a_50751_n19729.t208 a_52063_n8035# VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3250 VDD.t2825 VDD.t2824 VDD.t2825 VDD.t427 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3251 VDD.t2823 VDD.t2822 VDD.t2823 VDD.t2447 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3252 a_67111_n4447# a_50751_n19729.t209 a_66551_n4447# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3253 VSS.t2139 VSS.t2138 VSS.t2139 VSS.t905 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3254 VDD.t2821 VDD.t2820 VDD.t2821 VDD.t2464 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3255 VDD.t2819 VDD.t2818 VDD.t2819 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3256 VSS.t2137 VSS.t2136 VSS.t2137 VSS.t384 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3257 VDD.t2817 VDD.t2816 VDD.t2817 VDD.t2261 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3258 VDD.t2815 VDD.t2814 VDD.t2815 VDD.t780 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3259 a_52635_49681.t134 a_52635_34067.t151 VDD.t4889 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3260 a_54579_n7138# a_50751_n19729.t210 a_54019_n7138# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3261 VSS.t2135 VSS.t2134 VSS.t2135 VSS.t399 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3262 a_33249_48695.t249 a_31699_20742.t155 VDD.t177 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3263 a_61515_n35156# a_53699_n35156.t9 a_60677_n36322.t3 VDD.t544 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3264 a_52635_48695.t130 a_52635_34067.t152 VDD.t4888 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3265 VSS.t2133 VSS.t2132 VSS.t2133 VSS.t537 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3266 a_94892_4481.t3 a_94892_4481.t2 a_96818_7563# VSS.t396 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3267 VSS.t35 a_35502_25545.t61 a_33249_34067.t126 VSS.t18 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3268 a_71864_n28415# a_65486_n36322.t15 VDD.t296 VSS.t156 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3269 a_100820_11614.t2 a_100820_10448.t13 a_102756_10448# VDD.t322 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3270 VDD.t2813 VDD.t2811 VDD.t2813 VDD.t2812 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3271 VSS.t2131 VSS.t2130 VSS.t2131 VSS.t853 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3272 VSS.t2129 VSS.t2128 VSS.t2129 VSS.t553 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3273 VSS.t2127 VSS.t2126 VSS.t2127 VSS.t877 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3274 a_52635_48695.t129 a_52635_34067.t153 VDD.t4887 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3275 VDD.t2810 VDD.t2809 VDD.t2810 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3276 VDD.t2808 VDD.t2807 VDD.t2808 VDD.t2447 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3277 VSS.t46 a_35502_25545.t62 a_35922_19591.t4 VSS.t45 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X3278 VDD.t2806 VDD.t2805 VDD.t2806 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3279 VDD.t2804 VDD.t2803 VDD.t2804 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3280 VDD.t2802 VDD.t2801 VDD.t2802 VDD.t34 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3281 a_31284_n30339.t2 a_30324_n30399.t1 a_30724_n28415# VSS.t151 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3282 a_107339_n8770# a_71281_n8397.t213 a_106501_n7865# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3283 a_57977_n12421.t0 a_100820_11614.t11 a_107198_6405# VSS.t153 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3284 a_71896_12380# a_71496_10388.t19 a_71366_11614.t2 VDD.t351 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3285 a_47753_n16904# a_31953_n19727.t219 a_47231_n16904# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3286 a_114485_n30339# a_112559_n29181.t18 VSS.t3646 VSS.t413 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3287 a_61515_n33224# a_53699_n35156.t10 a_60677_n36322.t1 VDD.t544 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3288 VSS.t2125 VSS.t2124 VSS.t2125 VSS.t1064 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3289 VSS.t2123 VSS.t2122 VSS.t2123 VSS.t814 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3290 a_95414_n29181# a_94892_n29181.t7 a_94892_n29181.t8 VSS.t353 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3291 VDD.t2800 VDD.t2799 VDD.t2800 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3292 a_52635_48695.t44 a_35922_19591.t97 a_52635_34067.t8 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3293 VSS.t2121 VSS.t2120 VSS.t2121 VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3294 VSS.t2119 VSS.t2118 VSS.t2119 VSS.t106 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3295 VDD.t2798 VDD.t2797 VDD.t2798 VDD.t1099 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3296 a_32913_n14213# a_31953_n19727.t220 a_32353_n13316# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3297 VDD.t178 a_31699_20742.t156 a_33249_48695.t248 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3298 VDD.t2796 VDD.t2795 VDD.t2796 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3299 VSS.t2117 VSS.t2116 VSS.t2117 VSS.t896 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3300 VSS.t2115 VSS.t2114 VSS.t2115 VSS.t261 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3301 a_33249_48695.t52 a_33379_34917.t41 a_33249_35053.t38 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3302 VSS.t2113 VSS.t2112 VSS.t2113 VSS.t165 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3303 a_52635_49681.t42 a_35922_19591.t98 OUT.t65 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3304 a_85089_n34390# a_83153_n35156.t12 VDD.t4754 VDD.t1708 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3305 VSS.t2111 VSS.t2110 VSS.t2111 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3306 a_50629_n16009.t1 a_51711_n12421.t0 a_83725_7563# VSS.t311 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3307 a_52635_48695.t128 a_52635_34067.t154 VDD.t4886 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3308 a_32913_n8930.t0 a_31953_n19727.t221 a_32353_n8930# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3309 VSS.t2109 VSS.t2108 VSS.t2109 VSS.t615 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3310 VDD.t2794 VDD.t2793 VDD.t2794 VDD.t2399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3311 VSS.t2107 VSS.t2106 VSS.t2107 VSS.t1253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3312 VDD.t2792 VDD.t2791 VDD.t2792 VDD.t1439 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3313 a_33249_48695.t247 a_31699_20742.t157 VDD.t179 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3314 VDD.t2790 VDD.t2789 VDD.t2790 VDD.t1099 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3315 VDD.t2788 VDD.t2787 VDD.t2788 VDD.t548 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3316 a_65117_n12421# a_50751_n19729.t211 a_64243_n16009.t0 VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3317 a_45138_24920# a_35922_19591.t99 a_44608_24195# VDD.t405 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X3318 a_110225_n6055# a_71281_n8397.t214 a_109695_n5150# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3319 a_85089_10448# a_83153_10448.t19 VDD.t4789 VDD.t1442 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3320 VDD.t2786 VDD.t2785 VDD.t2786 VDD.t401 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3321 VSS.t2105 VSS.t2104 VSS.t2105 VSS.t531 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3322 VDD.t2784 VDD.t2783 VDD.t2784 VDD.t925 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3323 a_63683_n2653# a_50751_n19729.t212 a_63161_n2653# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3324 VSS.t2103 VSS.t2102 VSS.t2103 VSS.t1306 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3325 a_96818_7563# a_94892_4481.t17 VSS.t3641 VSS.t1303 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3326 VSS.t2101 VSS.t2100 VSS.t2101 VSS.t884 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3327 VSS.t2099 VSS.t2098 VSS.t2099 VSS.t576 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3328 a_33249_34067.t62 a_33379_34007.t48 a_33249_48695.t344 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3329 VDD.t2782 VDD.t2781 VDD.t2782 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3330 a_59411_n13318# a_50751_n19729.t213 a_58851_n12421# VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3331 VDD.t2780 VDD.t2779 VDD.t2780 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3332 VDD.t2778 VDD.t2776 VDD.t2778 VDD.t2777 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3333 VDD.t2775 VDD.t2773 VDD.t2775 VDD.t2774 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3334 VSS.t2097 VSS.t2096 VSS.t2097 VSS.t604 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3335 VDD.t2772 VDD.t2771 VDD.t2772 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3336 VSS.t2095 VSS.t2094 VSS.t2095 VSS.t1244 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X3337 VSS.t2093 VSS.t2092 VSS.t2093 VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3338 a_65677_n2653# a_50751_n19729.t214 a_65117_n2653# VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3339 VDD.t2770 VDD.t2769 VDD.t2770 VDD.t402 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X3340 VSS.t2091 VSS.t2090 VSS.t2091 VSS.t289 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3341 a_48951_4481.t1 a_47991_5507.t1 a_48391_5639# VSS.t340 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3342 a_110225_n14095# a_71281_n8397.t215 VDD.t481 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3343 VSS.t2089 VSS.t2088 VSS.t2089 VSS.t1294 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3344 VDD.t2768 VDD.t2767 VDD.t2768 VDD.t1917 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3345 a_79182_n35156# a_71366_n35156.t8 a_78344_n36322.t1 VDD.t2382 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3346 VDD.t2766 VDD.t2765 VDD.t2766 VDD.t2399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3347 VDD.t2764 VDD.t2763 VDD.t2764 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3348 VSS.t2087 VSS.t2086 VSS.t2087 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3349 a_52635_34067.t35 a_35922_19591.t100 a_52635_48695.t43 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3350 a_71281_n10073.t37 a_71281_n10073.t36 VDD.t357 VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3351 VSS.t2085 VSS.t2084 VSS.t2085 VSS.t498 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3352 a_111063_n2435# a_71281_n8397.t216 a_110225_n2435# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3353 VDD.t2762 VDD.t2761 VDD.t2762 VDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3354 VDD.t2760 VDD.t2759 VDD.t2760 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3355 VDD.t2758 VDD.t2757 VDD.t2758 VDD.t955 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3356 a_79182_12380# a_71366_11614.t7 a_78344_10448.t2 VDD.t571 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3357 a_112199_n8770# a_71281_n8397.t217 a_111631_n8770# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3358 VSS.t2083 VSS.t2082 VSS.t2083 VSS.t264 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3359 VSS.t2081 VSS.t2080 VSS.t2081 VSS.t1287 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3360 OUT.t64 a_35922_19591.t101 a_52635_49681.t43 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3361 VSS.t2079 VSS.t2078 VSS.t2079 VSS.t811 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3362 a_60080_5639# a_59558_4481.t13 a_53829_10388.t4 VSS.t397 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3363 a_33249_35053.t39 a_33379_34917.t42 a_33249_48695.t53 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3364 a_33249_48695.t246 a_31699_20742.t158 VDD.t180 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3365 VSS.t2077 VSS.t2076 VSS.t2077 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3366 a_60845_n2653# a_50751_n19729.t215 a_60285_n1756# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3367 VSS.t2075 VSS.t2074 VSS.t2075 VSS.t772 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3368 a_107230_n36322# a_106830_n36382.t17 VCM.t0 VDD.t1904 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3369 VDD.t2756 VDD.t2755 VDD.t2756 VDD.t910 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3370 a_33249_48695.t345 a_33379_34007.t49 a_33249_34067.t61 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3371 VSS.t2073 VSS.t2072 VSS.t2073 VSS.t307 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3372 a_33249_48695.t245 a_31699_20742.t159 VDD.t181 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3373 VDD.t2754 VDD.t2753 VDD.t2754 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3374 VSS.t2071 VSS.t2070 VSS.t2071 VSS.t591 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3375 VSS.t2069 VSS.t2068 VSS.t2069 VSS.t647 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3376 a_79182_n33224# a_71366_n35156.t9 a_78344_n36322.t2 VDD.t2382 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3377 a_51711_n3550# a_50751_n19729.t216 a_51151_n3550# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3378 VDD.t2752 VDD.t2751 VDD.t2752 VDD.t677 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3379 VDD.t2750 VDD.t2749 VDD.t2750 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3380 a_83725_7563# a_51711_n12421.t0 a_83153_11614.t2 VSS.t310 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3381 VSS.t2067 VSS.t2066 VSS.t2067 VSS.t336 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3382 VSS.t2065 VSS.t2064 VSS.t2065 VSS.t588 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3383 VDD.t2748 VDD.t2747 VDD.t2748 VDD.t674 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3384 a_33379_34007.t2 a_36162_n36382.t13 a_37968_n36322# VDD.t1893 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3385 a_77776_n35156# a_65658_n29313.t1 a_77225_n29181.t2 VDD.t2344 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3386 a_32353_n16904# a_31953_n19727.t222 a_31831_n17801# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3387 VDD.t414 a_35922_19591.t102 a_45706_22884# VDD.t407 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X3388 VDD.t2746 VDD.t2745 VDD.t2746 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3389 VSS.t2063 VSS.t2062 VSS.t2063 VSS.t684 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3390 VSS.t2061 VSS.t2060 VSS.t2061 VSS.t792 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3391 a_90245_n3340# a_71281_n10073.t189 a_89407_n3340# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3392 VDD.t2744 VDD.t2743 VDD.t2744 VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3393 VDD.t2742 VDD.t2741 VDD.t2742 VDD.t1081 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3394 a_44363_n16007.t2 a_65658_n29313.t2 a_66058_n27257# VSS.t377 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3395 VDD.t2740 VDD.t2739 VDD.t2740 VDD.t288 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3396 a_33249_34067.t125 a_35502_25545.t63 VSS.t53 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3397 a_33787_n19595# a_31953_n19727.t223 a_32913_n16007.t1 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3398 VDD.t2738 VDD.t2737 VDD.t2738 VDD.t1884 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3399 VDD.t2736 VDD.t2735 VDD.t2736 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3400 a_33249_35053.t40 a_33379_34917.t43 a_33249_48695.t54 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3401 VDD.t2734 VDD.t2733 VDD.t2734 VDD.t845 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3402 a_35781_n8930# a_31953_n19727.t224 a_35221_n8930# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3403 VSS.t2059 VSS.t2058 VSS.t2059 VSS.t633 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3404 VDD.t2732 VDD.t2731 VDD.t2732 VDD.t836 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3405 VDD.t2730 VDD.t2728 VDD.t2730 VDD.t2729 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3406 VSS.t2057 VSS.t2056 VSS.t2057 VSS.t671 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3407 VSS.t2055 VSS.t2054 VSS.t2055 VSS.t528 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3408 VDD.t2727 VDD.t2726 VDD.t2727 VDD.t935 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3409 VDD.t2725 VDD.t2724 VDD.t2725 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3410 a_77776_n33224# a_65658_n29313.t1 a_77225_n29181.t2 VDD.t2344 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3411 a_52635_49681.t133 a_52635_34067.t155 VDD.t4885 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3412 VSS.t2053 VSS.t2052 VSS.t2053 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3413 VDD.t2723 VDD.t2722 VDD.t2723 VDD.t1653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3414 VDD.t2721 VDD.t2720 VDD.t2721 VDD.t425 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3415 a_61515_10448# a_53699_11614.t6 a_60677_10448.t3 VDD.t3013 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3416 a_52635_49681.t44 a_35922_19591.t103 OUT.t63 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3417 a_113081_n27257# a_112559_n29181.t7 a_112559_n29181.t8 VSS.t410 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3418 VSS.t2051 VSS.t2050 VSS.t2051 VSS.t282 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3419 VDD.t2719 VDD.t2718 VDD.t2719 VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3420 VDD.t2717 VDD.t2716 VDD.t2717 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3421 a_30152_11614.t1 a_30324_5507.t1 a_32128_4481# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3422 VSS.t2049 VSS.t2048 VSS.t2049 VSS.t381 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3423 VSS.t2047 VSS.t2046 VSS.t2047 VSS.t609 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3424 a_59558_n29181.t4 a_59558_n29181.t3 a_61484_n30339# VSS.t398 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3425 VDD.t2715 VDD.t2714 VDD.t2715 VDD.t823 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3426 a_39179_n6239# a_31953_n19727.t225 a_38619_n6239# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3427 a_33249_48695.t244 a_31699_20742.t160 VDD.t182 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3428 a_52635_48695.t127 a_52635_34067.t156 VDD.t4884 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3429 VDD.t2713 VDD.t2712 VDD.t2713 VDD.t619 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3430 VDD.t2711 VDD.t2710 VDD.t2711 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3431 a_52635_48695.t126 a_52635_34067.t157 VDD.t4883 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3432 VSS.t442 a_36162_n36382.t14 a_36562_n35156# VDD.t2302 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3433 VDD.t2709 VDD.t2708 VDD.t2709 VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3434 VDD.t183 a_31699_20742.t161 a_33249_48695.t243 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3435 VDD.t4882 a_52635_34067.t158 a_52635_49681.t132 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3436 a_54019_n7138# a_50751_n19729.t217 a_53497_n8035# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3437 VSS.t324 a_77225_4481.t17 a_77747_5639# VSS.t323 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3438 VDD.t2707 VDD.t2706 VDD.t2707 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3439 a_82573_n21335# a_71281_n10073.t190 a_81735_n21335# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3440 VDD.t2705 VDD.t2704 VDD.t2705 VDD.t935 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3441 VDD.t2703 VDD.t2702 VDD.t2703 VDD.t810 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3442 a_33249_34067.t124 a_35502_25545.t64 VSS.t30 VSS.t29 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3443 a_33249_48695.t114 a_33379_34007.t50 a_33249_34067.t60 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3444 VSS.t2045 VSS.t2044 VSS.t2045 VSS.t305 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3445 VSS.t2043 VSS.t2042 VSS.t2043 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3446 VSS.t2041 VSS.t2040 VSS.t2041 VSS.t287 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3447 a_57417_n17803# a_50751_n19729.t218 a_56895_n17803# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3448 VSS.t2039 VSS.t2038 VSS.t2039 VSS.t612 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3449 a_53675_4481.t0 a_53829_10388.t17 a_54229_10448# VDD.t1405 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3450 a_30152_11614.t6 a_30152_10448.t14 a_32088_10448# VDD.t305 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3451 a_90969_n34390# a_89163_n36382.t14 VSS.t342 VDD.t549 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3452 VSS.t2037 VSS.t2035 VSS.t2037 VSS.t2036 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X3453 VDD.t2701 VDD.t2700 VDD.t2701 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3454 a_45138_24195# a_35922_19591.t104 a_44608_24195# VDD.t405 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X3455 a_33249_48695.t55 a_33379_34917.t44 a_33249_35053.t41 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3456 VDD.t184 a_31699_20742.t162 a_33249_48695.t242 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3457 VSS.t2034 VSS.t2033 VSS.t2034 VSS.t1253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3458 VDD.t2699 VDD.t2698 VDD.t2699 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3459 a_100235_n19525# a_71281_n8397.t218 a_99667_n19525# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3460 VSS.t2032 VSS.t2031 VSS.t2032 VSS.t638 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3461 VDD.t2697 VDD.t2696 VDD.t2697 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3462 a_36008_n27257.t2 a_36162_n36382.t15 a_36562_n33224# VDD.t2302 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3463 VDD.t4755 a_83153_n35156.t13 a_83683_n36322# VDD.t1850 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3464 VSS.t2030 VSS.t2029 VSS.t2030 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3465 VDD.t2695 VDD.t2694 VDD.t2695 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3466 a_46879_n14213# a_31953_n19727.t226 a_47753_n16007# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3467 a_33249_48695.t115 a_33379_34007.t51 a_33249_34067.t59 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3468 a_75585_n10073# I1N.t8 VSS.t432 VSS.t430 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X3469 VSS.t2028 VSS.t2027 VSS.t2028 VSS.t534 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3470 a_71342_4481.t0 a_65486_11614.t17 a_73268_7563# VSS.t422 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3471 VDD.t4881 a_52635_34067.t159 a_52635_49681.t131 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3472 VDD.t2693 VDD.t2692 VDD.t2693 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3473 VDD.t2691 VDD.t2690 VDD.t2691 VDD.t298 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3474 VDD.t2689 VDD.t2688 VDD.t2689 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3475 VDD.t2687 VDD.t2686 VDD.t2687 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3476 VDD.t2685 VDD.t2684 VDD.t2685 VDD.t2254 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3477 VSS.t2026 VSS.t2025 VSS.t2026 VSS.t105 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3478 VDD.t2683 VDD.t2682 VDD.t2683 VDD.t795 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3479 VDD.t2681 VDD.t2679 VDD.t2681 VDD.t2680 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3480 a_111631_n14095# a_71281_n8397.t219 a_111063_n14095# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3481 VSS.t386 a_77225_n29181.t16 a_77747_n27257# VSS.t384 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3482 OUT.t62 a_35922_19591.t105 a_52635_49681.t45 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3483 a_102796_4481# a_57977_n12421.t0 a_56895_n16009.t2 VSS.t172 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3484 VSS.t2024 VSS.t2023 VSS.t2024 VSS.t979 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3485 VDD.t2678 VDD.t2677 VDD.t2678 VDD.t404 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3486 VDD.t300 a_100820_11614.t12 a_108602_5639# VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3487 VSS.t2022 VSS.t2021 VSS.t2022 VSS.t748 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3488 VSS.t2020 VSS.t2019 VSS.t2020 VSS.t338 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3489 a_30324_5507.t1 a_30152_11614.t11 a_36530_5639# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3490 a_52635_34067.t58 a_35502_24538.t45 a_33249_34067.t8 VSS.t190 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3491 a_52635_48695.t42 a_35922_19591.t106 a_52635_34067.t12 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3492 VSS.t2018 VSS.t2017 VSS.t2018 VSS.t478 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3493 a_52585_n18700# a_50751_n19729.t219 a_52063_n18700# VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3494 a_98829_n19525# a_71281_n8397.t220 a_98299_n19525# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3495 VDD.t2676 VDD.t2675 VDD.t2676 VDD.t1824 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3496 VDD.t2674 VDD.t2673 VDD.t2674 VDD.t2254 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3497 VDD.t2672 VDD.t2671 VDD.t2672 VDD.t1821 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3498 VDD.t2670 VDD.t2669 VDD.t2670 VDD.t32 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3499 VDD.t185 a_31699_20742.t163 a_35502_25545.t13 VDD.t25 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3500 VSS.t2016 VSS.t2015 VSS.t2016 VSS.t357 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3501 VSS.t2014 VSS.t2013 VSS.t2014 VSS.t501 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3502 a_105365_n19525# a_71281_n8397.t221 a_104527_n19525# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3503 a_113110_n36322# a_103997_n8770.t10 a_106830_n36382.t1 VDD.t535 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3504 VDD.t2668 VDD.t2667 VDD.t2668 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3505 VDD.t2666 VDD.t2665 VDD.t2666 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3506 VDD.t2664 VDD.t2663 VDD.t2664 VDD.t538 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3507 VSS.t2012 VSS.t2011 VSS.t2012 VSS.t1222 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3508 a_53829_10388.t3 a_59558_4481.t14 a_61484_6405# VSS.t398 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3509 a_52635_34067.t30 a_35922_19591.t107 a_52635_48695.t41 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3510 VSS.t2010 VSS.t2009 VSS.t2010 VSS.t576 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3511 VSS.t2008 VSS.t2007 VSS.t2008 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3512 VSS.t2006 VSS.t2005 VSS.t2006 VSS.t490 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3513 a_65117_n2653# a_50751_n19729.t220 a_64595_n3550# VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3514 VDD.t2662 VDD.t2661 VDD.t2662 VDD.t1322 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3515 a_33249_35053.t42 a_33379_34917.t45 a_33249_48695.t56 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3516 VDD.t2660 VDD.t2659 VDD.t2660 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3517 a_95105_n18620# a_71281_n10073.t191 a_94537_n18620# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3518 a_33249_34067.t58 a_33379_34007.t52 a_33249_48695.t116 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3519 a_71864_7563# a_65486_11614.t18 a_71342_7563.t0 VSS.t423 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3520 a_66551_n7138# a_50751_n19729.t221 a_66029_n8035# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3521 a_52635_49681.t130 a_52635_34067.t160 VDD.t4880 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3522 a_90245_n18620# a_71281_n10073.t192 a_89407_n18620# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3523 a_33249_48695.t57 a_33379_34917.t46 a_33249_35053.t43 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3524 a_41891_n29181.t1 a_30324_n29313.t2 a_43848_n36322# VDD.t1796 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3525 a_110225_n4245# a_71281_n8397.t222 a_109695_n4245# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3526 VSS.t2004 VSS.t2003 VSS.t2004 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3527 VSS.t2002 VSS.t2001 VSS.t2002 VSS.t615 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3528 a_71281_n10073.t35 a_71281_n10073.t34 VDD.t376 VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3529 a_52635_49681.t46 a_35922_19591.t108 OUT.t61 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3530 a_31831_n5342.t2 a_32913_n8930.t1 a_83725_n30339# VSS.t288 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3531 VDD.t2658 VDD.t2657 VDD.t2658 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3532 VDD.t2656 VDD.t2655 VDD.t2656 VDD.t298 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3533 VDD.t2654 VDD.t2653 VDD.t2654 VDD.t120 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3534 VDD.t2652 VDD.t2651 VDD.t2652 VDD.t1570 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3535 VDD.t2650 VDD.t2649 VDD.t2650 VDD.t64 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3536 VDD.t482 a_71281_n8397.t223 a_100803_n13190# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3537 VDD.t2648 VDD.t2647 VDD.t2648 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3538 VSS.t26 a_35502_25545.t65 a_33249_34067.t123 VSS.t25 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3539 VDD.t4775 a_71266_n4019.t0 a_72596_n4019# VDD.t1188 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3540 VDD.t2646 VDD.t2645 VDD.t2646 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3541 VDD.t2644 VDD.t2643 VDD.t2644 VDD.t1780 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3542 VDD.t2642 VDD.t2641 VDD.t2642 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3543 VDD.t2640 VDD.t2639 VDD.t2640 VDD.t537 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3544 VSS.t237 a_50751_n19729.t36 a_50751_n19729.t37 VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3545 a_45445_n19595.t1 a_65486_n36322.t16 a_71864_n29181# VSS.t157 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3546 a_40613_n13316# a_31953_n19727.t227 a_40053_n12419# VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3547 VSS.t2000 VSS.t1999 VSS.t2000 VSS.t1157 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3548 VDD.t2638 VDD.t2637 VDD.t2638 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3549 VSS.t1998 VSS.t1997 VSS.t1998 VSS.t1594 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X3550 a_54579_n7138# a_50751_n19729.t222 a_54019_n6241# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3551 a_108602_5639# a_100820_11614.t13 a_57977_n12421.t0 VSS.t147 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3552 a_36530_5639# a_30152_11614.t12 VDD.t488 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3553 a_112199_n7865# a_71281_n8397.t224 a_111631_n7865# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3554 a_52635_48695.t40 a_35922_19591.t109 a_52635_34067.t13 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3555 a_88839_n18620# a_71281_n10073.t193 a_88271_n18620# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3556 a_54019_n19597# a_50751_n19729.t223 a_51711_n19597# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3557 a_40053_n13316# a_31953_n19727.t228 a_39531_n14213# VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3558 a_33249_48695.t58 a_33379_34917.t47 a_33249_35053.t44 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3559 a_94537_n6960# a_71281_n10073.t194 a_93969_n6960# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3560 VDD.t4879 a_52635_34067.t161 a_52635_49681.t129 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3561 VDD.t2636 VDD.t2635 VDD.t2636 VDD.t47 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3562 VSS.t1996 VSS.t1995 VSS.t1996 VSS.t106 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3563 VDD.t2634 VDD.t2633 VDD.t2634 VDD.t976 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3564 a_108636_n34390# a_106830_n36382.t18 VSS.t450 VDD.t1540 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3565 a_33249_34067.t122 a_35502_25545.t66 VSS.t50 VSS.t18 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3566 a_43010_n36322.t3 a_30324_n29313.t2 a_42442_n35156# VDD.t2189 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3567 VSS.t43 a_35502_25545.t67 a_33249_34067.t121 VSS.t37 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3568 a_52635_48695.t39 a_35922_19591.t110 a_52635_34067.t38 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3569 VDD.t2632 VDD.t2631 VDD.t2632 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3570 a_30724_n29181# a_30324_n29313.t0 a_30152_n35156.t0 VSS.t150 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3571 VSS.t1994 VSS.t1993 VSS.t1994 VSS.t459 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3572 a_60109_13546# a_53699_11614.t7 a_53829_10388.t1 VDD.t2542 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3573 VDD.t186 a_31699_20742.t164 a_35502_24538.t11 VDD.t16 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3574 VSS.t1992 VSS.t1991 VSS.t1992 VSS.t681 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3575 VDD.t2630 VDD.t2629 VDD.t2630 VDD.t720 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3576 a_35221_n8930# a_31953_n19727.t229 VSS.t114 VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3577 a_38619_n15110# a_31953_n19727.t230 a_38097_n15110# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3578 VDD.t2628 VDD.t2627 VDD.t2628 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3579 a_33249_34067.t57 a_33379_34007.t53 a_33249_48695.t117 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3580 VDD.t2626 VDD.t2625 VDD.t2626 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3581 VDD.t2624 VDD.t2623 VDD.t2624 VDD.t707 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3582 VDD.t2622 VDD.t2621 VDD.t2622 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3583 VSS.t1990 VSS.t1989 VSS.t1990 VSS.t733 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3584 VSS.t1988 VSS.t1987 VSS.t1988 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3585 VDD.t483 a_71281_n8397.t225 a_106501_n13190# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3586 VSS.t1986 VSS.t1985 VSS.t1986 VSS.t647 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3587 a_90245_n3340# a_71281_n10073.t195 a_89407_n2435# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3588 VSS.t1984 VSS.t1983 VSS.t1984 VSS.t395 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3589 VDD.t2620 VDD.t2619 VDD.t2620 VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3590 VSS.t1982 VSS.t1981 VSS.t1982 VSS.t531 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3591 a_100992_n29313.t0 a_100820_n36322.t15 a_107198_n27257# VSS.t336 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3592 VDD.t2618 VDD.t2617 VDD.t2618 VDD.t1142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3593 a_102796_n28415# a_100992_n29313.t0 a_38097_n5342.t1 VSS.t330 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3594 VSS.t1980 VSS.t1979 VSS.t1980 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3595 VDD.t2616 VDD.t2615 VDD.t2616 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3596 VDD.t2614 VDD.t2613 VDD.t2614 VDD.t336 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3597 VSS.t1978 VSS.t1977 VSS.t1978 VSS.t528 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3598 a_43010_n36322.t3 a_30324_n29313.t2 a_42442_n33224# VDD.t2189 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3599 VDD.t2612 VDD.t2611 VDD.t2612 VDD.t1747 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3600 a_60109_11614# a_53699_11614.t8 a_53829_10388.t2 VDD.t2542 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3601 VDD.t2610 VDD.t2609 VDD.t2610 VDD.t2160 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3602 a_83709_n8770# a_71281_n10073.t196 a_83141_n8770# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3603 VDD.t2608 VDD.t2607 VDD.t2608 VDD.t2155 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3604 VDD.t2606 VDD.t2605 VDD.t2606 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3605 VSS.t236 a_50751_n19729.t34 a_50751_n19729.t35 VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3606 VSS.t1976 VSS.t1975 VSS.t1976 VSS.t1104 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3607 a_52635_34067.t39 a_35922_19591.t111 a_52635_48695.t38 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3608 VSS.t1974 VSS.t1973 VSS.t1974 VSS.t553 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3609 VSS.t1972 VSS.t1971 VSS.t1972 VSS.t376 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3610 a_44885_n8033# a_31953_n19727.t231 a_44363_n8930# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3611 a_33249_35053.t124 a_35502_25545.t68 VSS.t20 VSS.t3 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3612 VDD.t2604 VDD.t2603 VDD.t2604 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3613 VDD.t2602 VDD.t2601 VDD.t2602 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3614 VSS.t1970 VSS.t1969 VSS.t1970 VSS.t633 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3615 VDD.t2600 VDD.t2599 VDD.t2600 VDD.t2142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3616 a_46879_n8930# a_31953_n19727.t232 a_46319_n8033# VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3617 a_85129_4481# a_51711_n12421.t0 a_50629_n16009.t2 VSS.t309 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3618 VSS.t1968 VSS.t1967 VSS.t1968 VSS.t10 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3619 VDD.t2598 VDD.t2597 VDD.t2598 VDD.t1505 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3620 VSS.t1966 VSS.t1965 VSS.t1966 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3621 a_52635_48695.t37 a_35922_19591.t112 a_52635_34067.t16 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3622 VDD.t2596 VDD.t2595 VDD.t2596 VDD.t1262 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3623 VDD.t2594 VDD.t2593 VDD.t2594 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3624 VDD.t2592 VDD.t2591 VDD.t2592 VDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3625 VSS.t1964 VSS.t1963 VSS.t1964 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3626 VDD.t2590 VDD.t2589 VDD.t2590 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3627 a_32913_n8930.t1 a_83153_n36322.t15 a_89531_n29181# VSS.t453 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3628 a_37934_n27257# a_30152_n36322.t15 a_30324_n29313.t0 VSS.t282 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3629 VDD.t2588 VDD.t2587 VDD.t2588 VDD.t2160 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3630 VDD.t2586 VDD.t2585 VDD.t2586 VDD.t2155 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3631 VSS.t1962 VSS.t1961 VSS.t1962 VSS.t699 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3632 VSS.t1960 VSS.t1959 VSS.t1960 VSS.t487 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3633 VDD.t2584 VDD.t2583 VDD.t2584 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3634 a_52635_49681.t47 a_35922_19591.t113 OUT.t60 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3635 VDD.t2582 VDD.t2581 VDD.t2582 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3636 a_37968_n35156# a_36162_n36382.t16 VSS.t443 VDD.t2127 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3637 a_89407_n9675# a_71281_n10073.t197 a_88839_n9675# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3638 VSS.t1958 VSS.t1957 VSS.t1958 VSS.t704 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3639 a_41487_n18698# a_31953_n19727.t233 a_40965_n18698# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3640 a_42047_n7136# a_31953_n19727.t234 a_41487_n7136# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3641 VDD.t2580 VDD.t2579 VDD.t2580 VDD.t2142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3642 VDD.t2578 VDD.t2577 VDD.t2578 VDD.t1489 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3643 VDD.t2576 VDD.t2575 VDD.t2576 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3644 VSS.t1956 VSS.t1955 VSS.t1956 VSS.t596 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3645 VDD.t2574 VDD.t2572 VDD.t2574 VDD.t2573 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3646 VSS.t427 a_36162_10388.t18 a_36562_12380# VDD.t3613 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3647 VSS.t1954 VSS.t1953 VSS.t1954 VSS.t568 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3648 a_77776_13546# a_71366_11614.t8 a_71496_10388.t5 VDD.t2924 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3649 a_55635_13546# a_53829_10388.t18 a_53675_4481.t1 VDD.t2921 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3650 a_48391_n29181# a_47991_n29313.t0 a_47819_n35156.t2 VSS.t339 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3651 a_33249_35053.t45 a_33379_34917.t48 a_33249_48695.t59 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3652 VDD.t2571 VDD.t2569 VDD.t2571 VDD.t2570 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3653 a_71281_n8397.t23 a_71281_n8397.t22 VDD.t441 VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3654 a_83153_n35156.t5 a_83153_n35156.t4 a_85089_n34390# VDD.t1486 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3655 VSS.t1952 VSS.t1951 VSS.t1952 VSS.t264 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3656 VSS.t1950 VSS.t1949 VSS.t1950 VSS.t612 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3657 a_33249_35053.t46 a_33379_34917.t49 a_33249_48695.t60 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3658 VDD.t2568 VDD.t2567 VDD.t2568 VDD.t1714 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3659 a_33249_35053.t104 a_35502_24538.t46 OUT.t10 VSS.t190 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3660 VDD.t2566 VDD.t2565 VDD.t2566 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3661 VSS.t1948 VSS.t1947 VSS.t1948 VSS.t1126 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3662 VSS.t1946 VSS.t1945 VSS.t1946 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3663 a_52635_49681.t128 a_52635_34067.t162 VDD.t4878 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3664 a_37968_n33224# a_36162_n36382.t17 a_36008_n30339.t3 VDD.t2127 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3665 a_51711_n3550# a_50751_n19729.t224 a_51151_n2653# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3666 a_33249_34067.t56 a_33379_34007.t54 a_33249_48695.t118 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3667 a_85089_n36322# a_83153_n35156.t14 VDD.t4756 VDD.t1708 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3668 VDD.t2564 VDD.t2563 VDD.t2564 VDD.t60 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3669 VDD.t30 a_31699_20742.t21 a_31699_20742.t22 VDD.t25 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3670 a_52635_49681.t127 a_52635_34067.t163 VDD.t4877 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3671 VDD.t2562 VDD.t2561 VDD.t2562 VDD.t1481 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3672 VSS.t1944 VSS.t1943 VSS.t1944 VSS.t307 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3673 a_87433_n6960# a_71281_n10073.t198 a_86903_n7865# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3674 VDD.t187 a_31699_20742.t165 a_33249_48695.t241 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3675 a_107198_7563# a_100820_11614.t14 a_106676_7563.t2 VSS.t182 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3676 VSS.t1942 VSS.t1941 VSS.t1942 VSS.t650 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3677 a_77776_11614# a_71366_11614.t9 a_71496_10388.t6 VDD.t2924 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3678 a_55635_11614# a_53829_10388.t19 VSS.t418 VDD.t2921 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3679 a_52635_34067.t39 a_35922_19591.t114 a_52635_48695.t36 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3680 VDD.t2560 VDD.t2558 VDD.t2560 VDD.t2559 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3681 VDD.t2557 VDD.t2556 VDD.t2557 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3682 VDD.t2555 VDD.t2554 VDD.t2555 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3683 VSS.t1940 VSS.t1939 VSS.t1940 VSS.t1111 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3684 a_44885_n18698# a_31953_n19727.t235 a_44363_n19595# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3685 VDD.t188 a_31699_20742.t166 a_33249_48695.t240 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3686 VDD.t2553 VDD.t2552 VDD.t2553 VDD.t630 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3687 VDD.t2551 VDD.t2550 VDD.t2551 VDD.t2099 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3688 a_47819_11614.t3 a_47819_10448.t15 a_49755_10448# VDD.t496 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3689 VDD.t2549 VDD.t2548 VDD.t2549 VDD.t898 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3690 VDD.t2547 VDD.t2546 VDD.t2547 VDD.t622 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3691 VSS.t1938 VSS.t1937 VSS.t1938 VSS.t1537 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3692 a_71496_n36382.t0 a_71366_n35156.t10 a_79182_n35156# VDD.t501 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3693 a_45445_n16007.t1 a_31953_n19727.t236 a_44885_n16007# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3694 a_95105_n8770# a_71281_n10073.t199 a_94537_n8770# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3695 VDD.t2545 VDD.t2544 VDD.t2545 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3696 VSS.t1936 VSS.t1935 VSS.t1936 VSS.t650 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3697 a_90935_n28415# a_83153_n36322.t16 a_32913_n8930.t1 VSS.t452 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3698 a_53145_n17803# a_50751_n19729.t225 a_52585_n17803# VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3699 VDD.t2543 VDD.t2541 VDD.t2543 VDD.t2542 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3700 a_114516_n34390# a_100992_n29313.t2 a_106809_n5150.t1 VDD.t536 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3701 VDD.t2540 VDD.t2539 VDD.t2540 VDD.t1658 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3702 VSS.t359 a_94892_n29181.t15 a_95414_n27257# VSS.t357 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3703 a_33249_48695.t61 a_33379_34917.t50 a_33249_35053.t47 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3704 VDD.t2538 VDD.t2537 VDD.t2538 VDD.t1206 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3705 VDD.t2536 VDD.t2535 VDD.t2536 VDD.t603 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3706 a_71281_n10073.t33 a_71281_n10073.t32 VDD.t344 VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3707 a_66551_n16009# a_50751_n19729.t226 a_65677_n14215# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3708 a_39179_n5342.t1 a_31953_n19727.t237 a_38619_n5342# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3709 VDD.t2534 VDD.t2533 VDD.t2534 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3710 VSS.t1934 VSS.t1933 VSS.t1934 VSS.t641 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3711 VDD.t2532 VDD.t2531 VDD.t2532 VDD.t2099 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3712 a_90245_n17715# a_71281_n10073.t200 a_89715_n17715.t0 VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3713 a_52585_n1756# a_50751_n19729.t227 a_51711_n5344.t0 VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3714 VDD.t484 a_71281_n8397.t226 a_106501_n1530# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3715 VSS.t1932 VSS.t1931 VSS.t1932 VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3716 VDD.t2530 VDD.t2529 VDD.t2530 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3717 VDD.t2528 VDD.t2527 VDD.t2528 VDD.t367 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3718 a_54019_n6241# a_50751_n19729.t228 a_53497_n6241# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3719 VDD.t2526 VDD.t2525 VDD.t2526 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3720 VSS.t1930 VSS.t1929 VSS.t1930 VSS.t576 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3721 a_71496_n36382.t1 a_71366_n35156.t11 a_79182_n33224# VDD.t501 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3722 a_32353_n4445# a_31953_n19727.t238 a_31831_n4445# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3723 VDD.t189 a_31699_20742.t167 a_33249_48695.t239 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3724 a_54579_n2653# a_50751_n19729.t229 a_54019_n1756# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3725 VDD.t2524 VDD.t2523 VDD.t2524 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3726 a_33249_35053.t48 a_33379_34917.t51 a_33249_48695.t62 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3727 a_33249_48695.t238 a_31699_20742.t168 VDD.t190 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3728 a_47819_11614.t5 a_47991_5507.t1 a_49795_6405# VSS.t337 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3729 VSS.t1928 VSS.t1927 VSS.t1928 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3730 a_31953_n19727.t39 a_31953_n19727.t38 VSS.t79 VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3731 VSS.t1926 VSS.t1925 VSS.t1926 VSS.t392 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3732 a_33249_34067.t120 a_35502_25545.t69 VSS.t36 VSS.t29 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3733 VDD.t191 a_31699_20742.t169 a_33249_48695.t237 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3734 VDD.t2522 VDD.t2521 VDD.t2522 VDD.t547 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3735 VDD.t2520 VDD.t2519 VDD.t2520 VDD.t543 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3736 VDD.t2518 VDD.t2517 VDD.t2518 VDD.t500 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3737 VSS.t1924 VSS.t1923 VSS.t1924 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3738 VSS.t1922 VSS.t1921 VSS.t1922 VSS.t905 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3739 VDD.t2516 VDD.t2515 VDD.t2516 VDD.t2079 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3740 VDD.t4876 a_52635_34067.t164 a_52635_49681.t126 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3741 VSS.t1920 VSS.t1919 VSS.t1920 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3742 VDD.t2514 VDD.t2513 VDD.t2514 VDD.t2076 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3743 VSS.t1918 VSS.t1917 VSS.t1918 VSS.t464 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3744 VSS.t1916 VSS.t1915 VSS.t1916 VSS.t306 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3745 VDD.t349 a_71281_n10073.t30 a_71281_n10073.t31 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3746 VSS.t1914 VSS.t1913 VSS.t1914 VSS.t294 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3747 VSS.t1912 VSS.t1911 VSS.t1912 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3748 VSS.t1910 VSS.t1909 VSS.t1910 VSS.t156 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3749 a_46319_n19595# a_31953_n19727.t239 a_45445_n16007.t0 VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3750 a_52635_48695.t35 a_35922_19591.t115 a_52635_34067.t40 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3751 a_73268_4481# a_65486_11614.t19 a_65658_4421.t0 VSS.t421 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3752 VDD.t2512 VDD.t2511 VDD.t2512 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3753 VSS.t1908 VSS.t1907 VSS.t1908 VSS.t41 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X3754 VDD.t2510 VDD.t2509 VDD.t2510 VDD.t1424 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3755 VDD.t2508 VDD.t2507 VDD.t2508 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3756 OUT.t59 a_35922_19591.t116 a_52635_49681.t48 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3757 VSS.t1906 VSS.t1905 VSS.t1906 VSS.t105 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3758 a_33249_34067.t7 a_35502_24538.t47 a_52635_34067.t62 VSS.t165 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3759 VDD.t2506 VDD.t2505 VDD.t2506 VDD.t425 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3760 a_31953_n19727.t73 a_71266_n4019.t0 a_75602_n3060# VDD.t1665 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3761 a_33249_35053.t49 a_33379_34917.t52 a_33249_48695.t63 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3762 VDD.t2504 VDD.t2503 VDD.t2504 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3763 VSS.t1904 VSS.t1903 VSS.t1904 VSS.t318 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3764 VDD.t2502 VDD.t2501 VDD.t2502 VDD.t2079 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3765 VDD.t2500 VDD.t2499 VDD.t2500 VDD.t1653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3766 VDD.t2498 VDD.t2497 VDD.t2498 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3767 a_65486_11614.t1 a_65486_10448.t16 a_67422_10448# VDD.t1378 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3768 VDD.t2496 VDD.t2495 VDD.t2496 VDD.t828 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3769 VDD.t2494 VDD.t2493 VDD.t2494 VDD.t2076 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3770 VSS.t1902 VSS.t1901 VSS.t1902 VSS.t151 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3771 VDD.t2492 VDD.t2491 VDD.t2492 VDD.t798 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3772 VSS.t1900 VSS.t1899 VSS.t1900 VSS.t60 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3773 a_52635_49681.t125 a_52635_34067.t165 VDD.t4875 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3774 a_43848_n35156# a_36032_n35156.t7 a_43010_n36322.t1 VDD.t2061 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3775 a_52635_48695.t125 a_52635_34067.t166 VDD.t4874 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3776 VSS.t1898 VSS.t1897 VSS.t1898 VSS.t795 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3777 a_54197_n28415# a_47819_n36322.t15 VDD.t493 VSS.t306 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3778 VDD.t2490 VDD.t2489 VDD.t2490 VDD.t1408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3779 a_44885_n3548# a_31953_n19727.t240 a_44363_n4445# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3780 VDD.t192 a_31699_20742.t170 a_33249_48695.t236 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3781 a_48391_6405# a_47991_4421.t0 a_47819_10448.t9 VSS.t339 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3782 VSS.t1896 VSS.t1895 VSS.t1896 VSS.t896 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3783 a_52635_48695.t124 a_52635_34067.t167 VDD.t4873 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3784 VSS.t1894 VSS.t1893 VSS.t1894 VSS.t1077 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X3785 a_46319_n8033# a_31953_n19727.t241 a_45797_n8033# VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3786 VDD.t2488 VDD.t2487 VDD.t2488 VDD.t1642 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3787 a_33249_48695.t235 a_31699_20742.t171 VDD.t193 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3788 a_95105_n21335# a_71281_n10073.t201 a_94537_n21335# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3789 VSS.t1892 VSS.t1891 VSS.t1892 VSS.t509 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3790 VDD.t4872 a_52635_34067.t168 a_52635_49681.t124 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3791 a_89033_n35156.t3 a_89163_n36382.t15 a_90969_n34390# VDD.t550 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3792 a_57417_n7138# a_50751_n19729.t230 a_56895_n7138# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3793 a_46879_n3548# a_31953_n19727.t242 a_46319_n3548# VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3794 VSS.t1890 VSS.t1889 VSS.t1890 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3795 VSS.t1888 VSS.t1887 VSS.t1888 VSS.t137 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3796 a_47753_n12419# a_31953_n19727.t243 a_45445_n12419# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3797 VDD.t379 a_71281_n10073.t202 a_89407_n21335# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3798 a_83709_n7865# a_71281_n10073.t203 a_83141_n7865# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3799 VSS.t1886 VSS.t1885 VSS.t1886 VSS.t262 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3800 VDD.t2486 VDD.t2484 VDD.t2486 VDD.t2485 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3801 VDD.t2483 VDD.t2482 VDD.t2483 VDD.t798 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3802 VDD.t2481 VDD.t2480 VDD.t2481 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3803 a_51151_n16009# a_50751_n19729.t231 a_50629_n16009.t0 VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3804 a_43848_n33224# a_36032_n35156.t8 a_43010_n36322.t3 VDD.t2061 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3805 VDD.t2479 VDD.t2478 VDD.t2479 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3806 VSS.t1884 VSS.t1883 VSS.t1884 VSS.t528 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3807 a_77747_n29181# a_77225_n29181.t9 a_77225_n29181.t10 VSS.t379 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3808 a_90969_n36322# a_89163_n36382.t16 a_89009_n27257.t3 VDD.t549 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3809 a_111631_n6960# a_71281_n8397.t227 a_111063_n6960# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3810 a_33249_35053.t50 a_33379_34917.t53 a_33249_48695.t64 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3811 VSS.t1882 VSS.t1881 VSS.t1882 VSS.t215 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3812 a_66551_n6241# a_50751_n19729.t232 a_66029_n6241# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3813 VDD.t2477 VDD.t2476 VDD.t2477 VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3814 VDD.t194 a_31699_20742.t172 a_35502_25545.t14 VDD.t14 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3815 VDD.t347 a_71281_n10073.t28 a_71281_n10073.t29 VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3816 VDD.t2475 VDD.t2474 VDD.t2475 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3817 VDD.t2473 VDD.t2472 VDD.t2473 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3818 VDD.t4871 a_52635_34067.t169 a_52635_49681.t123 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3819 VDD.t2471 VDD.t2470 VDD.t2471 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3820 a_108602_n28415# a_100820_n36322.t16 a_39179_n8930.t1 VSS.t334 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3821 VSS.t1880 VSS.t1879 VSS.t1880 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3822 VDD.t2469 VDD.t2468 VDD.t2469 VDD.t1714 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3823 a_52635_49681.t49 a_35922_19591.t117 OUT.t58 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3824 a_83709_n15000# a_71281_n10073.t204 a_83141_n15000# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3825 VDD.t4774 a_71266_n4019.t0 a_72596_n4978# VDD.t1188 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3826 VDD.t2467 VDD.t2466 VDD.t2467 VDD.t417 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3827 VSS.t1878 VSS.t1877 VSS.t1878 VSS.t884 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3828 VDD.t2465 VDD.t2463 VDD.t2465 VDD.t2464 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3829 VDD.t195 a_31699_20742.t173 a_33249_48695.t234 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3830 VDD.t2462 VDD.t2461 VDD.t2462 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3831 a_59411_n8932# a_50751_n19729.t233 a_58851_n8035# VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3832 VDD.t2460 VDD.t2459 VDD.t2460 VDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3833 a_66016_13546# a_65486_10448.t17 a_65486_11614.t3 VDD.t2261 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3834 VDD.t2458 VDD.t2457 VDD.t2458 VDD.t398 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3835 VDD.t2456 VDD.t2455 VDD.t2456 VDD.t780 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3836 VSS.t1876 VSS.t1875 VSS.t1876 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3837 a_33249_34067.t55 a_33379_34007.t55 a_33249_48695.t119 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3838 VDD.t2454 VDD.t2453 VDD.t2454 VDD.t792 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3839 VDD.t2452 VDD.t2451 VDD.t2452 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3840 a_31953_n19727.t37 a_31953_n19727.t36 VSS.t78 VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3841 a_67111_n15112# a_50751_n19729.t234 a_66551_n14215# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3842 a_88839_n21335# a_71281_n10073.t205 a_88271_n21335# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3843 VSS.t1874 VSS.t1873 VSS.t1874 VSS.t498 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3844 VSS.t1872 VSS.t1871 VSS.t1872 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3845 VDD.t196 a_31699_20742.t174 a_33249_48695.t233 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3846 VDD.t4870 a_52635_34067.t170 a_52635_49681.t122 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3847 a_65117_n18700# a_50751_n19729.t235 a_64595_n18700# VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3848 VDD.t2450 VDD.t2449 VDD.t2450 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3849 VSS.t3642 a_94892_4481.t18 a_95414_7563# VSS.t1037 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3850 a_33249_48695.t232 a_31699_20742.t175 VDD.t197 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3851 VSS.t1870 VSS.t1869 VSS.t1870 VSS.t1034 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3852 VSS.t1868 VSS.t1867 VSS.t1868 VSS.t158 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3853 VSS.t1866 VSS.t1865 VSS.t1866 VSS.t609 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3854 VDD.t2448 VDD.t2446 VDD.t2448 VDD.t2447 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3855 a_100803_n8770# a_71281_n8397.t228 a_100235_n8770# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3856 a_33249_34067.t119 a_35502_25545.t70 VSS.t52 VSS.t14 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3857 a_105933_n19525# a_71281_n8397.t229 a_105365_n19525# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3858 a_105365_n4245# a_71281_n8397.t230 a_104527_n4245# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3859 VDD.t2445 VDD.t2444 VDD.t2445 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3860 VDD.t2443 VDD.t2442 VDD.t2443 VDD.t780 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3861 VDD.t2441 VDD.t2440 VDD.t2441 VDD.t855 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3862 a_66016_11614# a_65486_10448.t18 a_65486_11614.t2 VDD.t2261 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3863 VDD.t2439 VDD.t2438 VDD.t2439 VDD.t18 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3864 a_59411_n19597# a_50751_n19729.t236 a_58851_n18700# VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3865 a_42047_n17801# a_31953_n19727.t244 a_41487_n17801# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3866 VSS.t1864 VSS.t1863 VSS.t1864 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3867 VSS.t1862 VSS.t1861 VSS.t1862 VSS.t338 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3868 VDD.t2437 VDD.t2436 VDD.t2437 VDD.t544 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3869 a_30152_n35156.t2 a_30324_n29313.t0 a_32128_n30339# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3870 a_38619_n14213# a_31953_n19727.t245 a_38097_n15110# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3871 VSS.t1860 VSS.t1859 VSS.t1860 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3872 VSS.t1858 VSS.t1857 VSS.t1858 VSS.t1025 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3873 VDD.t2435 VDD.t2434 VDD.t2435 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3874 VDD.t2433 VDD.t2432 VDD.t2433 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3875 a_35922_19591.t3 a_35502_25545.t71 VSS.t6 VSS.t5 nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X3876 VDD.t2431 VDD.t2430 VDD.t2431 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3877 a_93131_n17715# a_71281_n10073.t206 a_92601_n16810# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3878 VDD.t2429 VDD.t2428 VDD.t2429 VDD.t1665 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X3879 VDD.t2427 VDD.t2426 VDD.t2427 VDD.t568 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X3880 VDD.t2425 VDD.t2424 VDD.t2425 VDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3881 VSS.t1856 VSS.t1855 VSS.t1856 VSS.t1466 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3882 VSS.t1854 VSS.t1853 VSS.t1854 VSS.t21 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3883 VDD.t360 a_71281_n10073.t26 a_71281_n10073.t27 VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3884 VSS.t3647 a_112559_n29181.t19 a_113081_n30339# VSS.t411 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3885 a_93131_n15000# a_71281_n10073.t207 a_92601_n15905# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3886 VSS.t1852 VSS.t1851 VSS.t1852 VSS.t98 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3887 VDD.t2423 VDD.t2421 VDD.t2423 VDD.t2422 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3888 VDD.t198 a_31699_20742.t176 a_33249_48695.t231 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3889 VDD.t2420 VDD.t2419 VDD.t2420 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3890 a_88271_n15000# a_71281_n10073.t208 a_87433_n15000# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3891 VDD.t2418 VDD.t2417 VDD.t2418 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3892 a_31699_19142# I1U.t4 a_30377_19942# VSS.t349 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X3893 a_106501_n9675# a_71281_n8397.t231 a_105933_n9675# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3894 a_83153_n35156.t9 a_83325_n29313.t0 a_85129_n28415# VSS.t285 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3895 a_104527_n19525# a_71281_n8397.t232 a_103997_n19525# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3896 VDD.t2416 VDD.t2415 VDD.t2416 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3897 a_33249_48695.t120 a_33379_34007.t56 a_33249_34067.t54 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3898 a_52635_48695.t34 a_35922_19591.t118 a_52635_34067.t12 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3899 VDD.t2414 VDD.t2413 VDD.t2414 VDD.t1570 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3900 a_32353_n12419# a_31953_n19727.t246 a_31831_n13316# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3901 VSS.t1850 VSS.t1849 VSS.t1850 VSS.t859 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3902 a_95105_n7865# a_71281_n10073.t209 a_94537_n7865# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3903 VSS.t1848 VSS.t1847 VSS.t1848 VSS.t263 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3904 a_54019_n1756# a_50751_n19729.t237 VSS.t272 VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3905 VDD.t4869 a_52635_34067.t171 a_52635_49681.t121 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3906 a_83709_n20430# a_71281_n10073.t210 a_83141_n20430# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3907 a_37968_12380# a_36162_10388.t19 VSS.t428 VDD.t1711 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3908 VDD.t2412 VDD.t2411 VDD.t2412 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3909 a_52635_49681.t120 a_52635_34067.t172 VDD.t4868 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3910 VSS.t1846 VSS.t1845 VSS.t1846 VSS.t495 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3911 a_89407_n18620# a_71281_n10073.t211 a_88839_n18620# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3912 VSS.t1844 VSS.t1843 VSS.t1844 VSS.t537 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3913 VDD.t2410 VDD.t2409 VDD.t2410 VDD.t962 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X3914 a_83683_13546# a_83153_10448.t20 a_83153_11614.t6 VDD.t2774 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3915 a_95414_7563# a_94892_4481.t19 a_89163_10388.t2 VSS.t998 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3916 VSS.t1842 VSS.t1841 VSS.t1842 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3917 VDD.t2408 VDD.t2407 VDD.t2408 VDD.t748 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3918 a_100803_n18620# a_71281_n8397.t233 a_100235_n18620# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3919 VDD.t2406 VDD.t2405 VDD.t2406 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3920 VDD.t2404 VDD.t2403 VDD.t2404 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3921 VDD.t2402 VDD.t2401 VDD.t2402 VDD.t1549 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3922 a_33249_35053.t51 a_33379_34917.t54 a_33249_48695.t65 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3923 VDD.t2400 VDD.t2398 VDD.t2400 VDD.t2399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3924 VSS.t1840 VSS.t1839 VSS.t1840 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3925 VSS.t1838 VSS.t1837 VSS.t1838 VSS.t478 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3926 VDD.t2397 VDD.t2396 VDD.t2397 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3927 VDD.t2395 VDD.t2394 VDD.t2395 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3928 a_108636_n36322# a_106830_n36382.t19 a_106676_n27257.t3 VDD.t1540 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3929 VDD.t2393 VDD.t2392 VDD.t2393 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3930 VSS.t1836 VSS.t1835 VSS.t1836 VSS.t588 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3931 VDD.t2391 VDD.t2390 VDD.t2391 VDD.t1099 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3932 VDD.t2389 VDD.t2388 VDD.t2389 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3933 VDD.t2387 VDD.t2386 VDD.t2387 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3934 a_72596_n4019# a_71266_n4019.t0 a_71266_n4019.t0 VDD.t994 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X3935 VDD.t2385 VDD.t2384 VDD.t2385 VDD.t725 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3936 VSS.t1834 VSS.t1833 VSS.t1834 VSS.t699 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3937 a_52635_49681.t50 a_35922_19591.t119 OUT.t57 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3938 a_42413_n28415# a_41891_n29181.t19 a_36162_n36382.t1 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3939 a_41891_n29181.t6 a_41891_n29181.t5 a_43817_n30339# VSS.t168 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3940 a_37934_6405# a_30152_11614.t13 a_30324_5507.t1 VSS.t282 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3941 a_83683_11614# a_83153_10448.t21 a_83153_11614.t7 VDD.t2774 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3942 a_52635_34067.t32 a_35922_19591.t120 a_52635_48695.t33 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3943 VSS.t1832 VSS.t1831 VSS.t1832 VSS.t1426 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3944 a_106830_n36382.t4 a_112559_n29181.t20 a_114485_n29181# VSS.t409 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3945 VSS.t1830 VSS.t1829 VSS.t1830 VSS.t868 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3946 a_52635_48695.t123 a_52635_34067.t173 VDD.t4867 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3947 a_33249_34067.t53 a_33379_34007.t57 a_33249_48695.t121 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3948 a_39179_n18698# a_31953_n19727.t247 a_38619_n17801# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3949 a_33249_48695.t230 a_31699_20742.t177 VDD.t199 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3950 VDD.t2383 VDD.t2381 VDD.t2383 VDD.t2382 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3951 a_60845_n17803# a_50751_n19729.t238 a_60285_n16906# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3952 a_32913_n8033# a_31953_n19727.t248 a_32353_n8033# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3953 a_33249_48695.t229 a_31699_20742.t178 VDD.t200 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3954 VDD.t2380 VDD.t2379 VDD.t2380 VDD.t677 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3955 VSS.t1828 VSS.t1827 VSS.t1828 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3956 VDD.t2378 VDD.t2377 VDD.t2378 VDD.t508 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3957 VSS.t1826 VSS.t1825 VSS.t1826 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3958 VSS.t1824 VSS.t1823 VSS.t1824 VSS.t1431 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3959 VDD.t2376 VDD.t2375 VDD.t2376 VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3960 a_57417_n13318# a_50751_n19729.t239 a_56895_n13318# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3961 VDD.t2374 VDD.t2373 VDD.t2374 VDD.t674 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3962 VDD.t2372 VDD.t2371 VDD.t2372 VDD.t1917 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3963 a_93131_n20430# a_71281_n10073.t212 VDD.t380 VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3964 VSS.t1822 VSS.t1820 VSS.t1822 VSS.t1821 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X3965 a_33249_48695.t228 a_31699_20742.t179 VDD.t201 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3966 VSS.t1819 VSS.t1818 VSS.t1819 VSS.t905 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3967 VSS.t1817 VSS.t1816 VSS.t1817 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3968 VDD.t2370 VDD.t2369 VDD.t2370 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3969 VSS.t1815 VSS.t1814 VSS.t1815 VSS.t976 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3970 a_88271_n20430# a_71281_n10073.t213 a_87433_n20430# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3971 a_60285_n17803# a_50751_n19729.t240 a_59763_n18700# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3972 VSS.t1813 VSS.t1812 VSS.t1813 VSS.t376 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3973 VDD.t2368 VDD.t2367 VDD.t2368 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3974 VDD.t4768 a_30152_n36322.t16 a_37934_n29181# VSS.t281 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3975 a_94892_n29181.t6 a_94892_n29181.t5 a_96818_n28415# VSS.t352 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3976 a_71864_n27257# a_65486_n36322.t17 a_71342_n27257.t2 VSS.t156 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3977 VDD.t381 a_71281_n10073.t214 a_83709_n9675# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3978 a_46319_n3548# a_31953_n19727.t249 a_45797_n3548# VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3979 VDD.t2366 VDD.t2365 VDD.t2366 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3980 a_33249_48695.t66 a_33379_34917.t55 a_33249_35053.t52 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3981 a_107230_n35156# a_106830_n36382.t20 a_103997_n8770.t4 VDD.t1904 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3982 VDD.t2364 VDD.t2363 VDD.t2364 VDD.t498 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3983 VDD.t2362 VDD.t2361 VDD.t2362 VDD.t1642 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3984 VSS.t1811 VSS.t1810 VSS.t1811 VSS.t733 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3985 VDD.t2360 VDD.t2359 VDD.t2360 VDD.t677 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3986 VDD.t2358 VDD.t2357 VDD.t2358 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3987 VDD.t2356 VDD.t2355 VDD.t2356 VDD.t905 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3988 VDD.t2354 VDD.t2353 VDD.t2354 VDD.t674 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3989 VDD.t2352 VDD.t2351 VDD.t2352 VDD.t1917 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3990 VDD.t2350 VDD.t2348 VDD.t2350 VDD.t2349 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3991 VDD.t2347 VDD.t2346 VDD.t2347 VDD.t1505 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3992 VDD.t2345 VDD.t2343 VDD.t2345 VDD.t2344 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3993 a_66551_n1756# a_50751_n19729.t241 VSS.t273 VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3994 VDD.t2342 VDD.t2341 VDD.t2342 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3995 VDD.t2340 VDD.t2339 VDD.t2340 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3996 a_112199_n1530# a_71281_n8397.t234 a_111631_n1530# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3997 a_33249_34067.t52 a_33379_34007.t58 a_33249_48695.t122 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3998 VSS.t1809 VSS.t1808 VSS.t1809 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3999 a_33249_35053.t53 a_33379_34917.t56 a_33249_48695.t67 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4000 VDD.t2338 VDD.t2337 VDD.t2338 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4001 a_54579_n17803# a_50751_n19729.t242 a_54019_n16906# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4002 VDD.t2336 VDD.t2335 VDD.t2336 VDD.t925 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4003 a_31284_n30339.t1 a_30324_n29313.t1 a_30724_n27257# VSS.t151 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4004 a_36032_n35156.t2 a_36162_n36382.t18 a_37968_n35156# VDD.t1893 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4005 VDD.t2334 VDD.t2333 VDD.t2334 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4006 VDD.t202 a_31699_20742.t180 a_35502_24538.t10 VDD.t38 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4007 a_64243_n16906# a_50751_n19729.t243 a_63683_n16906# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4008 VSS.t1807 VSS.t1806 VSS.t1807 VSS.t837 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4009 VDD.t2332 VDD.t2331 VDD.t2332 VDD.t406 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4010 VDD.t2330 VDD.t2329 VDD.t2330 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4011 a_33787_n7136# a_31953_n19727.t250 a_33265_n8033# VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4012 VDD.t2328 VDD.t2327 VDD.t2328 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4013 VDD.t2326 VDD.t2324 VDD.t2326 VDD.t2325 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4014 a_107230_n33224# a_106830_n36382.t21 a_89033_n36322.t0 VDD.t1904 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4015 a_52635_48695.t32 a_35922_19591.t121 a_52635_34067.t41 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4016 a_48313_n4445# a_31953_n19727.t251 a_47753_n4445# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4017 VDD.t2323 VDD.t2322 VDD.t2323 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4018 VSS.t1805 VSS.t1804 VSS.t1805 VSS.t896 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4019 VSS.t77 a_31953_n19727.t34 a_31953_n19727.t35 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4020 a_66551_n15112# a_50751_n19729.t244 a_66029_n16906# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4021 a_59411_n3550# a_50751_n19729.t245 a_58851_n3550# VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4022 a_82573_n6960# a_71281_n10073.t215 a_81735_n6960# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4023 VDD.t2321 VDD.t2320 VDD.t2321 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4024 VSS.t434 I1N.t9 a_72603_n8397# VSS.t433 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X4025 a_33249_48695.t227 a_31699_20742.t181 VDD.t203 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4026 VDD.t2319 VDD.t2318 VDD.t2319 VDD.t1884 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4027 a_52635_49681.t119 a_52635_34067.t174 VDD.t4866 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4028 VDD.t2317 VDD.t2316 VDD.t2317 VDD.t1489 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4029 a_65677_n19597# a_50751_n19729.t246 a_65117_n19597# VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4030 VDD.t2315 VDD.t2314 VDD.t2315 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4031 a_45445_n8033# a_31953_n19727.t252 a_44885_n7136# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4032 a_114485_4481# a_112559_4481.t21 VSS.t303 VSS.t297 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4033 VSS.t1803 VSS.t1802 VSS.t1803 VSS.t1385 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4034 VDD.t2313 VDD.t2312 VDD.t2313 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4035 a_83709_n15905# a_71281_n10073.t216 a_83141_n15905# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4036 VDD.t2311 VDD.t2310 VDD.t2311 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4037 a_99667_n6960# a_71281_n8397.t235 a_98829_n6960# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4038 a_36032_n36322.t2 a_36162_n36382.t19 a_37968_n33224# VDD.t1893 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4039 a_83153_n35156.t1 a_83153_n35156.t0 a_85089_n36322# VDD.t1486 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4040 VSS.t1801 VSS.t1800 VSS.t1801 VSS.t817 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4041 a_64243_n8035# a_50751_n19729.t247 a_63683_n7138# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4042 VDD.t2309 VDD.t2308 VDD.t2309 VDD.t406 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4043 a_60080_n28415# a_59558_n29181.t18 a_53829_n36382.t3 VSS.t397 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4044 VSS.t1799 VSS.t1798 VSS.t1799 VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4045 VDD.t2307 VDD.t2306 VDD.t2307 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4046 OUT.t56 a_35922_19591.t122 a_52635_49681.t51 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4047 VDD.t2305 VDD.t2304 VDD.t2305 VDD.t910 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4048 a_113037_n20430# a_71281_n8397.t236 a_112199_n19525# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4049 VSS.t1797 VSS.t1796 VSS.t1797 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4050 VDD.t2303 VDD.t2301 VDD.t2303 VDD.t2302 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4051 VSS.t1795 VSS.t1793 VSS.t1795 VSS.t1794 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4052 a_33249_35053.t54 a_33379_34917.t57 a_33249_48695.t68 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4053 a_35781_n8930# a_31953_n19727.t253 a_35221_n8033# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4054 VDD.t2300 VDD.t2298 VDD.t2300 VDD.t2299 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X4055 VDD.t2297 VDD.t2296 VDD.t2297 VDD.t962 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4056 VDD.t2295 VDD.t2294 VDD.t2295 VDD.t1481 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4057 a_31953_n19727.t33 a_31953_n19727.t32 VSS.t76 VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4058 VDD.t2293 VDD.t2292 VDD.t2293 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4059 VDD.t2291 VDD.t2290 VDD.t2291 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4060 VDD.t2289 VDD.t2287 VDD.t2289 VDD.t2288 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4061 a_33249_48695.t123 a_33379_34007.t59 a_33249_34067.t51 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4062 VDD.t2286 VDD.t2285 VDD.t2286 VDD.t1884 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4063 a_57977_n16906# a_50751_n19729.t248 a_57417_n16906# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4064 VDD.t204 a_31699_20742.t182 a_33249_48695.t226 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4065 VSS.t1792 VSS.t1791 VSS.t1792 VSS.t884 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4066 a_35221_n19595# a_31953_n19727.t254 VSS.t115 VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4067 a_65658_4421.t0 a_65486_11614.t20 a_71864_7563# VSS.t424 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4068 VDD.t2284 VDD.t2283 VDD.t2284 VDD.t47 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4069 a_52635_49681.t118 a_52635_34067.t175 VDD.t4865 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4070 VDD.t2282 VDD.t2281 VDD.t2282 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4071 VSS.t1790 VSS.t1789 VSS.t1790 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4072 a_33249_48695.t69 a_33379_34917.t58 a_33249_35053.t55 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4073 VDD.t2280 VDD.t2279 VDD.t2280 VDD.t935 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4074 VDD.t4864 a_52635_34067.t176 a_52635_48695.t122 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4075 VDD.t2278 VDD.t2277 VDD.t2278 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4076 VDD.t2276 VDD.t2275 VDD.t2276 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4077 VSS.t1788 VSS.t1787 VSS.t1788 VSS.t475 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4078 VDD.t2274 VDD.t2273 VDD.t2274 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4079 VDD.t2272 VDD.t2271 VDD.t2272 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4080 VSS.t1786 VSS.t1785 VSS.t1786 VSS.t721 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4081 VSS.t1784 VSS.t1783 VSS.t1784 VSS.t937 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4082 a_100803_n7865# a_71281_n8397.t237 a_100235_n7865# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4083 VDD.t2270 VDD.t2269 VDD.t2270 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4084 OUT.t9 a_35502_24538.t48 a_33249_35053.t101 VSS.t183 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4085 VDD.t2268 VDD.t2267 VDD.t2268 VDD.t1251 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4086 VDD.t2266 VDD.t2265 VDD.t2266 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4087 VDD.t4863 a_52635_34067.t177 a_52635_49681.t117 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4088 VDD.t2264 VDD.t2263 VDD.t2264 VDD.t625 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4089 VDD.t2262 VDD.t2260 VDD.t2262 VDD.t2261 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4090 a_39179_n19595.t0 a_47819_n36322.t16 a_54197_n29181# VSS.t304 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4091 VDD.t2259 VDD.t2258 VDD.t2259 VDD.t866 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4092 VDD.t2257 VDD.t2256 VDD.t2257 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4093 a_88839_n8770# a_71281_n10073.t217 a_88271_n8770# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4094 VSS.t1782 VSS.t1781 VSS.t1782 VSS.t808 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4095 VDD.t2255 VDD.t2253 VDD.t2255 VDD.t2254 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4096 VDD.t4757 a_83153_n35156.t15 a_83683_n35156# VDD.t1850 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4097 VDD.t2252 VDD.t2250 VDD.t2252 VDD.t2251 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4098 VDD.t382 a_71281_n10073.t218 a_95105_n9675# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4099 a_114516_n36322# a_100992_n29313.t2 a_106809_n5150.t0 VDD.t536 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4100 OUT.t55 a_35922_19591.t123 a_52635_49681.t52 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4101 VDD.t2249 VDD.t2248 VDD.t2249 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4102 a_93131_n15905# a_71281_n10073.t219 a_92601_n15905# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4103 a_113110_12380# a_100992_4421.t1 a_112559_4481.t9 VDD.t337 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4104 VSS.t1780 VSS.t1779 VSS.t1780 VSS.t687 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4105 a_89407_n3340# a_71281_n10073.t220 a_88839_n3340# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4106 VSS.t1778 VSS.t1777 VSS.t1778 VSS.t213 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4107 a_67462_4481# a_64243_n1756.t1 a_63161_n5344.t2 VSS.t289 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4108 a_88271_n15905# a_71281_n10073.t221 a_87433_n15905# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4109 a_46274_24920# a_35922_19591.t124 a_45706_24920# VDD.t407 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X4110 a_48349_12380# a_47819_10448.t6 a_47819_10448.t7 VDD.t507 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4111 a_44885_n2651# a_31953_n19727.t255 a_44363_n2651# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4112 VSS.t1776 VSS.t1775 VSS.t1776 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4113 a_52635_49681.t53 a_35922_19591.t125 OUT.t54 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4114 VSS.t1774 VSS.t1773 VSS.t1774 VSS.t330 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4115 VDD.t346 a_71281_n10073.t24 a_71281_n10073.t25 VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4116 VDD.t2247 VDD.t2246 VDD.t2247 VDD.t49 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4117 a_33249_35053.t123 a_35502_25545.t72 VSS.t4 VSS.t3 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4118 VDD.t205 a_31699_20742.t183 a_33249_48695.t225 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4119 VDD.t2245 VDD.t2244 VDD.t2245 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4120 a_57417_n6241# a_50751_n19729.t249 a_56895_n7138# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4121 a_46879_n2651# a_31953_n19727.t256 a_46319_n2651# VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4122 a_52635_48695.t31 a_35922_19591.t126 a_52635_34067.t42 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4123 a_93969_n15000# a_71281_n10073.t222 a_93131_n15000# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4124 VSS.t1772 VSS.t1771 VSS.t1772 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4125 a_89163_10388.t3 a_94892_4481.t20 a_96818_4481# VSS.t396 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4126 VSS.t403 a_59558_4481.t15 a_60080_6405# VSS.t401 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4127 VDD.t4758 a_83153_n35156.t16 a_83683_n33224# VDD.t1850 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4128 VSS.t1770 VSS.t1769 VSS.t1770 VSS.t399 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4129 VDD.t350 a_71281_n10073.t22 a_71281_n10073.t23 VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4130 VDD.t2243 VDD.t2242 VDD.t2243 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4131 VDD.t2241 VDD.t2239 VDD.t2241 VDD.t2240 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4132 a_33249_35053.t122 a_35502_25545.t73 VSS.t2 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4133 VDD.t2238 VDD.t2237 VDD.t2238 VDD.t1824 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4134 OUT.t53 a_35922_19591.t127 a_52635_49681.t54 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4135 VSS.t1768 VSS.t1767 VSS.t1768 VSS.t329 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4136 a_83153_11614.t0 a_51711_n12421.t0 a_85129_6405# VSS.t308 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4137 VDD.t2236 VDD.t2235 VDD.t2236 VDD.t1821 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4138 a_51151_n15112# a_50751_n19729.t250 a_50629_n15112# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4139 VSS.t1766 VSS.t1765 VSS.t1766 VSS.t908 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4140 a_33249_34067.t50 a_33379_34007.t60 a_33249_48695.t124 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4141 a_33249_35053.t94 a_35502_24538.t49 OUT.t8 VSS.t165 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4142 a_33249_35053.t56 a_33379_34917.t59 a_33249_48695.t70 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4143 a_71281_n10073.t21 a_71281_n10073.t20 VDD.t359 VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4144 VDD.t2234 VDD.t2233 VDD.t2234 VDD.t2231 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4145 a_52635_48695.t121 a_52635_34067.t178 VDD.t4862 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4146 a_102756_13546# a_100820_10448.t14 VDD.t299 VDD.t298 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4147 VSS.t1764 VSS.t1763 VSS.t1764 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4148 VDD.t2232 VDD.t2230 VDD.t2232 VDD.t2231 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4149 VDD.t2229 VDD.t2227 VDD.t2229 VDD.t2228 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4150 a_32913_n18698# a_31953_n19727.t257 a_32353_n18698# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4151 VSS.t1762 VSS.t1761 VSS.t1762 VSS.t215 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4152 a_42047_n2651# a_31953_n19727.t258 a_41487_n1754# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4153 a_113110_n35156# a_100992_n29313.t2 a_112559_n29181.t1 VDD.t535 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4154 VDD.t440 a_71281_n8397.t20 a_71281_n8397.t21 VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4155 VSS.t1760 VSS.t1759 VSS.t1760 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4156 VSS.t1758 VSS.t1757 VSS.t1758 VSS.t1064 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4157 VDD.t2226 VDD.t2225 VDD.t2226 VDD.t677 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4158 VDD.t2224 VDD.t2223 VDD.t2224 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4159 VSS.t1756 VSS.t1755 VSS.t1756 VSS.t763 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4160 VDD.t2222 VDD.t2221 VDD.t2222 VDD.t1824 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4161 VDD.t2220 VDD.t2219 VDD.t2220 VDD.t1424 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4162 a_32913_n3548# a_31953_n19727.t259 a_32353_n3548# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4163 VSS.t1754 VSS.t1753 VSS.t1754 VSS.t775 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4164 VDD.t2218 VDD.t2217 VDD.t2218 VDD.t1821 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4165 a_34347_n14213# a_31953_n19727.t260 a_33787_n14213# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4166 VSS.t1752 VSS.t1751 VSS.t1752 VSS.t834 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4167 VSS.t1750 VSS.t1749 VSS.t1750 VSS.t868 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4168 VDD.t2216 VDD.t2215 VDD.t2216 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4169 VDD.t2214 VDD.t2213 VDD.t2214 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4170 a_36162_n36382.t4 a_36032_n35156.t9 a_43848_n35156# VDD.t1796 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4171 a_102756_11614# a_100820_10448.t15 VDD.t419 VDD.t298 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4172 a_50629_n16009.t2 a_83325_4421.t2 a_83725_4481# VSS.t311 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4173 VSS.t1748 VSS.t1747 VSS.t1748 VSS.t377 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4174 OUT.t52 a_35922_19591.t128 a_52635_49681.t55 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4175 VDD.t2212 VDD.t2211 VDD.t2212 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4176 VDD.t2210 VDD.t2209 VDD.t2210 VDD.t297 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4177 a_33249_35053.t57 a_33379_34917.t60 a_33249_48695.t71 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4178 a_113110_n33224# a_100992_n29313.t2 a_112559_n29181.t1 VDD.t535 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4179 VDD.t2208 VDD.t2207 VDD.t2208 VDD.t1195 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4180 a_35502_25545.t15 a_31699_20742.t184 VDD.t206 VDD.t14 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4181 VSS.t1746 VSS.t1745 VSS.t1746 VSS.t281 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4182 a_83141_n8770# a_71281_n10073.t223 a_82573_n8770# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4183 VDD.t2206 VDD.t2205 VDD.t2206 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4184 VDD.t2204 VDD.t2203 VDD.t2204 VDD.t1780 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4185 VSS.t1744 VSS.t1743 VSS.t1744 VSS.t1253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4186 VDD.t2202 VDD.t2201 VDD.t2202 VDD.t1408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4187 VSS.t1742 VSS.t1741 VSS.t1742 VSS.t317 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4188 VDD.t2200 VDD.t2199 VDD.t2200 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4189 a_52635_48695.t30 a_35922_19591.t129 a_52635_34067.t22 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4190 VSS.t1740 VSS.t1739 VSS.t1740 VSS.t484 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4191 a_52635_49681.t56 a_35922_19591.t130 OUT.t51 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4192 VSS.t1738 VSS.t1737 VSS.t1738 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4193 VSS.t210 a_35502_25545.t74 a_33249_34067.t118 VSS.t14 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4194 VDD.t2198 VDD.t2197 VDD.t2198 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4195 a_100235_n8770# a_71281_n8397.t238 a_99667_n8770# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4196 VSS.t1736 VSS.t1735 VSS.t1736 VSS.t335 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4197 a_36162_n36382.t6 a_36032_n35156.t10 a_43848_n33224# VDD.t1796 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4198 VSS.t1734 VSS.t1733 VSS.t1734 VSS.t224 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4199 a_71366_n36322.t3 a_89163_n36382.t17 a_90969_n36322# VDD.t550 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4200 VSS.t1732 VSS.t1731 VSS.t1732 VSS.t1306 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4201 a_96818_4481# a_94892_4481.t21 VSS.t3643 VSS.t1303 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4202 VDD.t4861 a_52635_34067.t179 a_52635_49681.t116 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4203 VSS.t1730 VSS.t1729 VSS.t1730 VSS.t576 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4204 VSS.t1728 VSS.t1727 VSS.t1728 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4205 VDD.t2196 VDD.t2195 VDD.t2196 VDD.t925 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4206 a_54019_n16009# a_50751_n19729.t251 a_53145_n14215# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4207 a_63683_n17803# a_50751_n19729.t252 a_63161_n17803# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4208 VDD.t2194 VDD.t2193 VDD.t2194 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4209 VSS.t1726 VSS.t1725 VSS.t1726 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4210 VDD.t2192 VDD.t2191 VDD.t2192 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4211 VSS.t1724 VSS.t1723 VSS.t1724 VSS.t259 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4212 a_93969_n20430# a_71281_n10073.t224 a_93131_n20430# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4213 VDD.t2190 VDD.t2188 VDD.t2190 VDD.t2189 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4214 VDD.t2187 VDD.t2186 VDD.t2187 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4215 VDD.t2185 VDD.t2184 VDD.t2185 VDD.t320 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4216 VDD.t2183 VDD.t2182 VDD.t2183 VDD.t1747 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4217 VSS.t1722 VSS.t1721 VSS.t1722 VSS.t1294 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4218 a_81735_n6055# a_71281_n10073.t225 a_81205_n5150# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4219 a_99667_n18620# a_71281_n8397.t239 a_98829_n18620# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4220 VDD.t2181 VDD.t2180 VDD.t2181 VDD.t1780 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4221 VSS.t1720 VSS.t1719 VSS.t1720 VSS.t1315 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4222 VDD.t2179 VDD.t2178 VDD.t2179 VDD.t1549 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4223 VDD.t2177 VDD.t2176 VDD.t2177 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4224 a_95414_n30339# a_94892_n29181.t16 a_89163_n36382.t1 VSS.t353 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4225 VSS.t1718 VSS.t1717 VSS.t1718 VSS.t1287 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4226 a_38097_n5342.t1 a_39179_n8930.t1 a_101392_n28415# VSS.t332 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4227 a_33249_35053.t58 a_33379_34917.t61 a_33249_48695.t72 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4228 a_72603_n9297# I1N.t10 a_71281_n10073.t73 VSS.t429 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X4229 a_111063_n18620# a_71281_n8397.t240 a_110225_n18620# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4230 a_98829_n6055# a_71281_n8397.t241 a_98299_n5150# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4231 VDD.t2175 VDD.t2174 VDD.t2175 VDD.t2118 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4232 a_89407_n21335# a_71281_n10073.t226 a_88839_n21335# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4233 VSS.t1716 VSS.t1715 VSS.t1716 VSS.t877 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4234 VSS.t1714 VSS.t1713 VSS.t1714 VSS.t148 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4235 VSS.t209 a_35502_25545.t24 a_35502_25545.t25 VSS.t45 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X4236 VDD.t2173 VDD.t2172 VDD.t2173 VDD.t1183 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4237 VDD.t2171 VDD.t2170 VDD.t2171 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4238 a_31953_n19727.t31 a_31953_n19727.t30 VSS.t75 VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4239 VSS.t1712 VSS.t1711 VSS.t1712 VSS.t452 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4240 a_113037_n8770# a_71281_n8397.t242 a_112199_n8770# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4241 a_52635_49681.t57 a_35922_19591.t131 OUT.t50 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4242 VDD.t2169 VDD.t2168 VDD.t2169 VDD.t910 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4243 a_100803_n21335# a_71281_n8397.t243 a_100235_n21335# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4244 VDD.t2167 VDD.t2166 VDD.t2167 VDD.t1747 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4245 a_46274_23609# a_35922_19591.t132 a_45706_24195# VDD.t407 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X4246 VSS.t1710 VSS.t1709 VSS.t1710 VSS.t817 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4247 a_100992_4421.t0 a_100820_11614.t15 a_107198_7563# VSS.t153 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4248 VSS.t1708 VSS.t1707 VSS.t1708 VSS.t740 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4249 VDD.t2165 VDD.t2164 VDD.t2165 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4250 VDD.t2163 VDD.t2162 VDD.t2163 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4251 a_35221_n8033# a_31953_n19727.t261 a_34699_n8033# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4252 VDD.t2161 VDD.t2159 VDD.t2161 VDD.t2160 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4253 a_83725_4481# a_83325_4421.t2 a_83153_10448.t1 VSS.t310 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4254 a_106501_n19525# a_71281_n8397.t244 a_105933_n19525# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4255 VDD.t2158 VDD.t2157 VDD.t2158 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4256 a_35781_n4445# a_31953_n19727.t262 a_35221_n3548# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4257 a_60109_10448# a_47991_4421.t1 a_59558_4481.t10 VDD.t2542 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4258 VDD.t2156 VDD.t2154 VDD.t2156 VDD.t2155 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4259 a_87433_n6055# a_71281_n10073.t227 a_86903_n9675# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4260 VDD.t2153 VDD.t2152 VDD.t2153 VDD.t697 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4261 a_53145_n13318# a_50751_n19729.t253 a_52585_n13318# VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4262 VSS.t1706 VSS.t1705 VSS.t1706 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4263 VDD.t2151 VDD.t2150 VDD.t2151 VDD.t1373 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4264 a_101111_n6055.t1 a_71281_n8397.t245 a_100803_n9675# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4265 a_72596_n4978# a_71266_n4019.t0 a_31953_n19727.t72 VDD.t994 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X4266 VDD.t2149 VDD.t2148 VDD.t2149 VDD.t1370 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4267 VDD.t2147 VDD.t2146 VDD.t2147 VDD.t326 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4268 a_73268_n28415# a_65486_n36322.t18 a_45445_n19595.t1 VSS.t154 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4269 VDD.t2145 VDD.t2144 VDD.t2145 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4270 a_52635_48695.t29 a_35922_19591.t133 a_52635_34067.t22 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4271 VDD.t2143 VDD.t2141 VDD.t2143 VDD.t2142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4272 VDD.t2140 VDD.t2139 VDD.t2140 VDD.t499 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4273 VDD.t2138 VDD.t2137 VDD.t2138 VDD.t1365 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4274 VSS.t1704 VSS.t1703 VSS.t1704 VSS.t856 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4275 VDD.t2136 VDD.t2135 VDD.t2136 VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4276 a_33249_35053.t95 a_35502_24538.t50 OUT.t7 VSS.t185 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4277 VSS.t1702 VSS.t1701 VSS.t1702 VSS.t908 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4278 VSS.t34 a_35502_25545.t75 a_33249_35053.t121 VSS.t33 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4279 a_52635_34067.t63 a_35502_24538.t51 a_33249_34067.t6 VSS.t183 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4280 VSS.t1700 VSS.t1699 VSS.t1700 VSS.t528 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4281 VDD.t2134 VDD.t2133 VDD.t2134 VDD.t1714 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4282 a_83709_n1530# a_71281_n10073.t228 a_83141_n1530# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4283 VDD.t2132 VDD.t2131 VDD.t2132 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4284 VSS.t1698 VSS.t1697 VSS.t1698 VSS.t853 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4285 VDD.t2130 VDD.t2129 VDD.t2130 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4286 a_33249_34067.t49 a_33379_34007.t61 a_33249_48695.t125 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4287 VDD.t2128 VDD.t2126 VDD.t2128 VDD.t2127 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4288 a_63683_n8932# a_50751_n19729.t254 a_63161_n8932# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4289 a_33249_34067.t48 a_33379_34007.t62 a_33249_48695.t126 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4290 a_96818_n29181# a_94892_n29181.t17 VSS.t360 VSS.t354 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4291 VDD.t2125 VDD.t2124 VDD.t2125 VDD.t1354 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4292 a_57417_n12421# a_50751_n19729.t255 a_56895_n13318# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4293 a_42442_12380# a_30324_4421.t1 a_41891_4481.t0 VDD.t288 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4294 a_41487_n15110# a_31953_n19727.t263 a_40965_n16904# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4295 VDD.t2123 VDD.t2122 VDD.t2123 VDD.t893 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4296 a_65677_n8932# a_50751_n19729.t256 a_65117_n8932# VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4297 VDD.t2121 VDD.t2120 VDD.t2121 VDD.t1349 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4298 a_52635_48695.t120 a_52635_34067.t180 VDD.t4860 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4299 VDD.t2119 VDD.t2117 VDD.t2119 VDD.t2118 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4300 a_33249_35053.t59 a_33379_34917.t62 a_33249_48695.t73 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4301 a_52635_48695.t119 a_52635_34067.t181 VDD.t4859 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4302 VDD.t2116 VDD.t2115 VDD.t2116 VDD.t554 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4303 a_35502_24538.t9 a_31699_20742.t185 VDD.t207 VDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4304 VSS.t1696 VSS.t1695 VSS.t1696 VSS.t1615 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4305 a_88839_n7865# a_71281_n10073.t229 a_88271_n7865# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4306 VDD.t208 a_31699_20742.t186 a_33249_48695.t224 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4307 VDD.t2114 VDD.t2113 VDD.t2114 VDD.t1714 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4308 a_87433_n17715# a_71281_n10073.t230 a_86903_n16810# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4309 VSS.t1694 VSS.t1693 VSS.t1694 VSS.t484 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4310 a_46319_n2651# a_31953_n19727.t264 a_45797_n3548# VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4311 VSS.t1692 VSS.t1691 VSS.t1692 VSS.t591 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4312 a_52635_49681.t115 a_52635_34067.t182 VDD.t4858 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4313 a_47753_n7136# a_31953_n19727.t265 a_47231_n8033# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4314 a_57417_n1756# a_50751_n19729.t257 a_56895_n2653# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4315 a_93131_n6055# a_71281_n10073.t231 a_92601_n5150# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4316 VSS.t40 a_35502_25545.t76 a_33249_35053.t120 VSS.t39 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4317 a_33249_48695.t223 a_31699_20742.t187 VDD.t209 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4318 a_52635_49681.t114 a_52635_34067.t183 VDD.t4857 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4319 a_87433_n15000# a_71281_n10073.t232 a_86903_n15905# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4320 a_89407_n2435# a_71281_n10073.t233 a_88839_n2435# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4321 VSS.t1690 VSS.t1689 VSS.t1690 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4322 VSS.t1688 VSS.t1687 VSS.t1688 VSS.t165 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4323 VSS.t1686 VSS.t1685 VSS.t1686 VSS.t588 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4324 VDD.t210 a_31699_20742.t188 a_33249_48695.t222 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4325 VSS.t1684 VSS.t1683 VSS.t1684 VSS.t304 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4326 VDD.t2112 VDD.t2111 VDD.t2112 VDD.t1957 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4327 VDD.t2110 VDD.t2109 VDD.t2110 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4328 VSS.t1682 VSS.t1681 VSS.t1682 VSS.t306 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4329 VDD.t2108 VDD.t2107 VDD.t2108 VDD.t2 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4330 a_30324_n30399.t1 a_30152_n36322.t17 a_36530_n28415# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4331 a_85089_n35156# a_83153_n35156.t17 VDD.t4759 VDD.t1708 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4332 VDD.t2106 VDD.t2105 VDD.t2106 VDD.t1127 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4333 a_93969_n15905# a_71281_n10073.t234 a_93131_n15905# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4334 VSS.t1680 VSS.t1679 VSS.t1680 VSS.t671 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4335 VDD.t2104 VDD.t2103 VDD.t2104 VDD.t1658 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4336 VDD.t2102 VDD.t2101 VDD.t2102 VDD.t78 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4337 a_71342_7563.t1 a_65486_11614.t21 a_73268_4481# VSS.t422 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4338 a_55635_10448# a_53829_10388.t20 a_53675_7563.t0 VDD.t2921 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4339 VSS.t1678 VSS.t1677 VSS.t1678 VSS.t1360 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4340 a_77776_10448# a_65658_4421.t2 a_77225_4481.t8 VDD.t2924 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4341 VDD.t2100 VDD.t2098 VDD.t2100 VDD.t2099 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4342 a_44885_n15110# a_31953_n19727.t266 a_44363_n15110# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4343 a_102796_n27257# a_39179_n8930.t1 a_38097_n5342.t2 VSS.t330 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4344 VSS.t1676 VSS.t1675 VSS.t1676 VSS.t1256 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4345 a_59411_n2653# a_50751_n19729.t258 a_58851_n2653# VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4346 VDD.t2097 VDD.t2096 VDD.t2097 VDD.t501 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4347 a_61484_5639# a_59558_4481.t16 VSS.t404 VSS.t399 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4348 VSS.t1674 VSS.t1673 VSS.t1674 VSS.t763 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4349 a_85089_n33224# a_83153_n35156.t18 VDD.t4760 VDD.t1708 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4350 VSS.t1672 VSS.t1671 VSS.t1672 VSS.t681 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4351 VSS.t1670 VSS.t1669 VSS.t1670 VSS.t537 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4352 VSS.t1668 VSS.t1667 VSS.t1668 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4353 VDD.t2095 VDD.t2094 VDD.t2095 VDD.t1512 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4354 a_105933_n8770# a_71281_n8397.t246 a_105365_n8770# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4355 VDD.t2093 VDD.t2092 VDD.t2093 VDD.t1658 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4356 VSS.t1666 VSS.t1665 VSS.t1666 VSS.t334 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4357 a_33249_48695.t221 a_31699_20742.t189 VDD.t211 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4358 a_52635_48695.t118 a_52635_34067.t184 VDD.t4856 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4359 a_64243_n6241# a_50751_n19729.t259 a_63683_n6241# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4360 a_48951_4481.t1 a_47991_4421.t0 a_48391_6405# VSS.t340 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4361 VSS.t1664 VSS.t1663 VSS.t1664 VSS.t68 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4362 a_33249_48695.t220 a_31699_20742.t190 VDD.t212 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4363 a_33249_48695.t219 a_31699_20742.t191 VDD.t213 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4364 VDD.t2091 VDD.t2090 VDD.t2091 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4365 VDD.t214 a_31699_20742.t192 a_35502_24538.t8 VDD.t38 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4366 a_106501_n3340# a_71281_n8397.t247 a_105933_n3340# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4367 VDD.t2089 VDD.t2087 VDD.t2089 VDD.t2088 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4368 VDD.t215 a_31699_20742.t193 a_33249_48695.t218 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4369 a_31953_n19727.t29 a_31953_n19727.t28 VSS.t74 VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4370 VSS.t1662 VSS.t1661 VSS.t1662 VSS.t811 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4371 a_60080_6405# a_59558_4481.t2 a_59558_4481.t3 VSS.t397 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4372 VDD.t2086 VDD.t2085 VDD.t2086 VDD.t406 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4373 a_95105_n1530# a_71281_n10073.t235 a_94537_n1530# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4374 VSS.t1660 VSS.t1659 VSS.t1660 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4375 VSS.t1658 VSS.t1657 VSS.t1658 VSS.t149 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4376 VDD.t2084 VDD.t2083 VDD.t2084 VDD.t390 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4377 a_104527_n6055# a_71281_n8397.t248 a_103997_n5150# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4378 VSS.t1656 VSS.t1655 VSS.t1656 VSS.t264 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4379 a_112199_n13190# a_71281_n8397.t249 a_111631_n13190# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4380 a_71864_4481# a_65486_11614.t22 a_71342_4481.t1 VSS.t423 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4381 a_83141_n7865# a_71281_n10073.t236 a_82573_n7865# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4382 VSS.t1654 VSS.t1653 VSS.t1654 VSS.t609 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4383 a_71281_n8397.t19 a_71281_n8397.t18 VDD.t438 VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4384 VDD.t2082 VDD.t2081 VDD.t2082 VDD.t287 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4385 VSS.t1652 VSS.t1651 VSS.t1652 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4386 a_52635_49681.t58 a_35922_19591.t134 OUT.t49 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4387 VDD.t2080 VDD.t2078 VDD.t2080 VDD.t2079 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4388 a_87433_n20430# a_71281_n10073.t237 VDD.t383 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4389 VSS.t1650 VSS.t1649 VSS.t1650 VSS.t534 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4390 VDD.t2077 VDD.t2075 VDD.t2077 VDD.t2076 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4391 VDD.t2074 VDD.t2073 VDD.t2074 VDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4392 VDD.t2072 VDD.t2071 VDD.t2072 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4393 a_100235_n7865# a_71281_n8397.t250 a_99667_n7865# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4394 VDD.t2070 VDD.t2069 VDD.t2070 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4395 VSS.t73 a_31953_n19727.t26 a_31953_n19727.t27 VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4396 VSS.t1648 VSS.t1647 VSS.t1648 VSS.t145 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4397 a_52635_48695.t28 a_35922_19591.t135 a_52635_34067.t43 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4398 a_83709_n14095# a_71281_n10073.t238 a_83141_n14095# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4399 VSS.t1646 VSS.t1645 VSS.t1646 VSS.t792 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4400 VSS.t1644 VSS.t1643 VSS.t1644 VSS.t644 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4401 VSS.t72 a_31953_n19727.t24 a_31953_n19727.t25 VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4402 VDD.t2068 VDD.t2067 VDD.t2068 VDD.t1354 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4403 a_40053_n18698# a_31953_n19727.t267 a_39531_n18698# VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4404 a_52635_49681.t113 a_52635_34067.t185 VDD.t4855 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4405 VDD.t2066 VDD.t2065 VDD.t2066 VDD.t1642 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4406 VSS.t1642 VSS.t1641 VSS.t1642 VSS.t531 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4407 VDD.t2064 VDD.t2063 VDD.t2064 VDD.t667 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4408 a_81735_n4245# a_71281_n10073.t239 a_81205_n4245# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4409 VDD.t437 a_71281_n8397.t16 a_71281_n8397.t17 VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4410 VSS.t1640 VSS.t1639 VSS.t1640 VSS.t1157 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4411 VSS.t1638 VSS.t1637 VSS.t1638 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4412 VDD.t4854 a_52635_34067.t186 a_52635_48695.t117 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4413 a_42047_n13316# a_31953_n19727.t268 a_41487_n13316# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4414 VSS.t1636 VSS.t1635 VSS.t1636 VSS.t478 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4415 VDD.t216 a_31699_20742.t194 a_33249_48695.t217 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4416 a_41487_n4445# a_31953_n19727.t269 a_40965_n6239# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4417 a_52635_49681.t112 a_52635_34067.t187 VDD.t4853 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4418 a_35221_n3548# a_31953_n19727.t270 a_34699_n3548# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4419 VSS.t1634 VSS.t1633 VSS.t1634 VSS.t285 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4420 VDD.t2062 VDD.t2060 VDD.t2062 VDD.t2061 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4421 VDD.t2059 VDD.t2057 VDD.t2059 VDD.t2058 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4422 VDD.t2056 VDD.t2055 VDD.t2056 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4423 VDD.t2054 VDD.t2053 VDD.t2054 VDD.t1653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4424 VDD.t436 a_71281_n8397.t14 a_71281_n8397.t15 VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4425 a_98829_n4245# a_71281_n8397.t251 a_98299_n4245# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4426 VDD.t2052 VDD.t2051 VDD.t2052 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4427 a_52585_n14215# a_50751_n19729.t260 a_52063_n14215# VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4428 a_57977_n8035# a_50751_n19729.t261 a_57417_n7138# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4429 a_67462_n28415# a_65658_n29313.t0 a_44363_n16007.t1 VSS.t289 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4430 VDD.t2050 VDD.t2049 VDD.t2050 VDD.t674 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4431 VSS.t1632 VSS.t1631 VSS.t1632 VSS.t172 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4432 VDD.t2048 VDD.t2047 VDD.t2048 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4433 a_113037_n8770# a_71281_n8397.t252 a_112199_n7865# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4434 a_33249_34067.t47 a_33379_34007.t63 a_33249_48695.t127 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4435 VDD.t2046 VDD.t2045 VDD.t2046 VDD.t1642 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4436 VSS.t1630 VSS.t1629 VSS.t1630 VSS.t286 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4437 VSS.t325 a_77225_4481.t18 a_77747_6405# VSS.t323 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4438 VDD.t2044 VDD.t2043 VDD.t2044 VDD.t502 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4439 a_95943_n17715# a_71281_n10073.t240 a_95413_n16810.t1 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4440 VDD.t2042 VDD.t2041 VDD.t2042 VDD.t1099 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4441 a_84547_n3340# a_71281_n10073.t241 a_83709_n3340# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4442 VDD.t2040 VDD.t2039 VDD.t2040 VDD.t64 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4443 a_33249_34067.t5 a_35502_24538.t52 a_52635_34067.t64 VSS.t185 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4444 VDD.t2038 VDD.t2037 VDD.t2038 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4445 a_33249_35053.t60 a_33379_34917.t63 a_33249_48695.t74 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4446 a_90935_n27257# a_83153_n36322.t17 a_83325_n29313.t0 VSS.t452 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4447 VDD.t2036 VDD.t2035 VDD.t2036 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4448 VDD.t4852 a_52635_34067.t188 a_52635_48695.t116 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4449 a_95943_n15000# a_71281_n10073.t242 a_95105_n15000# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4450 VDD.t2034 VDD.t2033 VDD.t2034 VDD.t1653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4451 VDD.t2032 VDD.t2031 VDD.t2032 VDD.t635 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4452 VDD.t2030 VDD.t2029 VDD.t2030 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4453 VDD.t2028 VDD.t2027 VDD.t2028 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4454 VDD.t2026 VDD.t2025 VDD.t2026 VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4455 a_93131_n14095# a_71281_n10073.t243 IBPOUT.t0 VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4456 VDD.t2024 VDD.t2023 VDD.t2024 VDD.t798 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4457 a_110225_n18620# a_71281_n8397.t253 a_109695_n19525# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4458 VDD.t2022 VDD.t2020 VDD.t2022 VDD.t2021 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4459 a_32913_n3548# a_31953_n19727.t271 a_32353_n2651# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4460 VDD.t2019 VDD.t2018 VDD.t2019 VDD.t1251 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4461 a_90969_n35156# a_89163_n36382.t18 VSS.t343 VDD.t549 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4462 a_52635_49681.t111 a_52635_34067.t189 VDD.t4851 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4463 a_88271_n14095# a_71281_n10073.t244 a_87433_n14095# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4464 a_33249_48695.t75 a_33379_34917.t64 a_33249_35053.t61 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4465 VDD.t2017 VDD.t2016 VDD.t2017 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4466 VDD.t2015 VDD.t2014 VDD.t2015 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4467 VSS.t1628 VSS.t1627 VSS.t1628 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4468 VDD.t2013 VDD.t2012 VDD.t2013 VDD.t1052 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4469 a_65117_n8932# a_50751_n19729.t262 VSS.t274 VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4470 VSS.t1626 VSS.t1625 VSS.t1626 VSS.t757 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4471 a_59558_4481.t5 a_59558_4481.t4 a_61484_7563# VSS.t398 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4472 VSS.t1624 VSS.t1623 VSS.t1624 VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4473 VDD.t2011 VDD.t2010 VDD.t2011 VDD.t1180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4474 VDD.t217 a_31699_20742.t195 a_33249_48695.t216 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4475 VSS.t1622 VSS.t1621 VSS.t1622 VSS.t160 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4476 VDD.t4850 a_52635_34067.t190 a_52635_48695.t115 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4477 VDD.t2009 VDD.t2008 VDD.t2009 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4478 VSS.t1620 VSS.t1619 VSS.t1620 VSS.t684 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4479 a_90969_12380# a_89163_10388.t18 VSS.t347 VDD.t555 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4480 VDD.t2007 VDD.t2006 VDD.t2007 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4481 VDD.t2005 VDD.t2004 VDD.t2005 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4482 a_65658_n29313.t0 a_65486_n36322.t19 a_71864_n30339# VSS.t157 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4483 VSS.t1618 VSS.t1617 VSS.t1618 VSS.t454 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4484 VDD.t2003 VDD.t2002 VDD.t2003 VDD.t610 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4485 a_71281_n10073.t19 a_71281_n10073.t18 VDD.t371 VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4486 VSS.t1616 VSS.t1614 VSS.t1616 VSS.t1615 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4487 VDD.t2001 VDD.t2000 VDD.t2001 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4488 VDD.t4849 a_52635_34067.t191 a_52635_49681.t110 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4489 a_94537_n15000# a_71281_n10073.t245 a_93969_n15000# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4490 VDD.t1999 VDD.t1998 VDD.t1999 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4491 VDD.t1997 VDD.t1995 VDD.t1997 VDD.t1996 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4492 a_90969_n33224# a_89163_n36382.t19 a_89009_n30339.t2 VDD.t549 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4493 VSS.t1613 VSS.t1612 VSS.t1613 VSS.t671 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4494 VDD.t1994 VDD.t1993 VDD.t1994 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4495 VSS.t1611 VSS.t1610 VSS.t1611 VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4496 VSS.t1609 VSS.t1608 VSS.t1609 VSS.t748 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4497 VDD.t421 a_100820_11614.t16 a_108602_6405# VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4498 a_30324_5507.t1 a_30152_11614.t14 a_36530_6405# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4499 VSS.t1607 VSS.t1606 VSS.t1607 VSS.t340 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4500 VSS.t1605 VSS.t1604 VSS.t1605 VSS.t352 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4501 VSS.t1603 VSS.t1602 VSS.t1603 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4502 a_54019_n15112# a_50751_n19729.t263 a_53497_n16906# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4503 a_99667_n21335# a_71281_n8397.t254 a_98829_n21335# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4504 a_30724_n30339# a_30324_n30399.t1 a_30152_n36322.t0 VSS.t150 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4505 a_39179_n14213# a_31953_n19727.t272 a_38619_n13316# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4506 a_79151_n28415# a_77225_n29181.t17 VSS.t387 VSS.t381 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4507 a_87433_n15905# a_71281_n10073.t246 a_86903_n15905# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4508 VSS.t1601 VSS.t1600 VSS.t1601 VSS.t609 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4509 VDD.t1992 VDD.t1991 VDD.t1992 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4510 VDD.t1990 VDD.t1989 VDD.t1990 VDD.t390 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4511 VDD.t1988 VDD.t1987 VDD.t1988 VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4512 VDD.t1986 VDD.t1985 VDD.t1986 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4513 VDD.t1984 VDD.t1983 VDD.t1984 VDD.t429 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4514 a_93131_n4245# a_71281_n10073.t247 a_92601_n4245# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4515 a_33249_48695.t215 a_31699_20742.t196 VDD.t218 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4516 a_33787_n1754# a_31953_n19727.t273 VSS.t116 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4517 VSS.t1599 VSS.t1598 VSS.t1599 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4518 VDD.t1982 VDD.t1981 VDD.t1982 VDD.t780 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4519 a_66016_10448# a_65486_10448.t6 a_65486_10448.t7 VDD.t2261 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4520 a_111063_n21335# a_71281_n8397.t255 a_110225_n21335# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4521 VDD.t1980 VDD.t1979 VDD.t1980 VDD.t303 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4522 VDD.t1978 VDD.t1977 VDD.t1978 VDD.t401 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4523 a_35781_n17801# a_31953_n19727.t274 a_35221_n16904# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4524 a_33249_48695.t214 a_31699_20742.t197 VDD.t219 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4525 VSS.t1597 VSS.t1596 VSS.t1597 VSS.t1157 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4526 a_60285_n13318# a_50751_n19729.t264 a_59763_n14215# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4527 VSS.t1595 VSS.t1593 VSS.t1595 VSS.t1594 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X4528 VDD.t1976 VDD.t1975 VDD.t1976 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4529 a_33249_48695.t213 a_31699_20742.t198 VDD.t220 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4530 a_45445_n1754# a_31953_n19727.t275 a_44885_n1754# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4531 VSS.t1592 VSS.t1591 VSS.t1592 VSS.t108 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4532 VDD.t1974 VDD.t1973 VDD.t1974 VDD.t1209 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4533 a_83141_n13190# a_71281_n10073.t248 a_82573_n13190# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4534 a_100803_n1530# a_71281_n8397.t256 a_100235_n1530# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4535 a_83725_n28415# a_32913_n8930.t1 a_83153_n36322.t0 VSS.t287 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4536 a_95943_n20430# a_71281_n10073.t249 a_95105_n20430# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4537 a_52635_48695.t114 a_52635_34067.t192 VDD.t4848 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4538 a_54197_n27257# a_47819_n36322.t17 a_53675_n27257.t3 VSS.t306 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4539 VDD.t1972 VDD.t1971 VDD.t1972 VDD.t1015 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4540 a_64243_n1756.t0 a_50751_n19729.t265 a_63683_n1756# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4541 VSS.t1590 VSS.t1589 VSS.t1590 VSS.t1126 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4542 VSS.t1588 VSS.t1587 VSS.t1588 VSS.t1253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4543 VSS.t1586 VSS.t1585 VSS.t1586 VSS.t638 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4544 VSS.t1584 VSS.t1583 VSS.t1584 VSS.t56 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4545 VDD.t1970 VDD.t1969 VDD.t1970 VDD.t1549 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4546 VDD.t291 a_65486_n36322.t20 a_73268_n29181# VSS.t155 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4547 a_95943_n3340# a_71281_n10073.t250 a_95105_n3340# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4548 a_35781_n2651# a_31953_n19727.t276 a_35221_n2651# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4549 VDD.t1968 VDD.t1967 VDD.t1968 VDD.t917 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4550 VSS.t1582 VSS.t1581 VSS.t1582 VSS.t733 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4551 VDD.t1966 VDD.t1965 VDD.t1966 VDD.t1570 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4552 a_33249_34067.t46 a_33379_34007.t64 a_33249_48695.t128 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4553 VDD.t1964 VDD.t1963 VDD.t1964 VDD.t1195 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4554 a_107198_4481# a_100820_11614.t17 a_106676_4481.t3 VSS.t182 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4555 VDD.t1962 VDD.t1961 VDD.t1962 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4556 a_105933_n7865# a_71281_n8397.t257 a_105365_n7865# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4557 a_53145_n13318# a_50751_n19729.t266 a_52585_n12421# VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4558 VSS.t1580 VSS.t1579 VSS.t1580 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4559 VDD.t1960 VDD.t1959 VDD.t1960 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4560 VSS.t1578 VSS.t1577 VSS.t1578 VSS.t531 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4561 VSS.t1576 VSS.t1575 VSS.t1576 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4562 VDD.t1958 VDD.t1956 VDD.t1958 VDD.t1957 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4563 VDD.t1955 VDD.t1954 VDD.t1955 VDD.t1439 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4564 VDD.t1953 VDD.t1952 VDD.t1953 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4565 VDD.t1951 VDD.t1950 VDD.t1951 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4566 a_52635_48695.t113 a_52635_34067.t193 VDD.t4847 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4567 VSS.t1574 VSS.t1573 VSS.t1574 VSS.t1111 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4568 VSS.t1572 VSS.t1571 VSS.t1572 VSS.t397 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4569 a_81735_n13190# a_71281_n10073.t251 a_81205_n16810# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4570 VDD.t328 a_71281_n10073.t16 a_71281_n10073.t17 VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4571 VDD.t1949 VDD.t1948 VDD.t1949 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4572 a_35502_25545.t16 a_31699_20742.t199 VDD.t221 VDD.t18 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4573 VDD.t1947 VDD.t1946 VDD.t1947 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4574 a_83325_n29313.t0 a_83153_n36322.t18 a_89531_n30339# VSS.t453 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4575 a_106501_n2435# a_71281_n8397.t258 a_105933_n2435# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4576 a_94537_n20430# a_71281_n10073.t252 a_93969_n20430# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4577 a_108602_6405# a_100820_11614.t18 a_57977_n12421.t0 VSS.t147 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4578 a_36530_6405# a_30152_11614.t15 VDD.t489 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4579 VDD.t1945 VDD.t1944 VDD.t1945 VDD.t1183 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4580 a_52635_48695.t27 a_35922_19591.t136 a_52635_34067.t1 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4581 a_49795_5639# a_47991_4421.t0 a_48951_4481.t1 VSS.t338 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4582 VDD.t1943 VDD.t1942 VDD.t1943 VDD.t1549 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4583 a_32128_n29181# a_30324_n30399.t2 a_31284_n30339.t2 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4584 VDD.t1941 VDD.t1940 VDD.t1941 VDD.t320 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4585 a_108602_n27257# a_100820_n36322.t17 a_100992_n29313.t0 VSS.t334 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4586 a_49755_13546# a_47819_10448.t16 VDD.t512 VDD.t508 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4587 VDD.t1939 VDD.t1938 VDD.t1939 VDD.t1570 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4588 a_52635_49681.t109 a_52635_34067.t194 VDD.t4846 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4589 VSS.t1570 VSS.t1569 VSS.t1570 VSS.t550 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4590 VDD.t1937 VDD.t1935 VDD.t1937 VDD.t1936 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4591 VDD.t1934 VDD.t1933 VDD.t1934 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4592 VDD.t1932 VDD.t1931 VDD.t1932 VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4593 VDD.t4773 a_71266_n4019.t0 a_72596_n3060# VDD.t1188 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X4594 a_52635_49681.t59 a_35922_19591.t137 OUT.t48 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4595 a_33249_48695.t212 a_31699_20742.t200 VDD.t222 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4596 VDD.t1930 VDD.t1929 VDD.t1930 VDD.t1177 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4597 a_108636_n35156# a_106830_n36382.t22 VSS.t451 VDD.t1540 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4598 a_111631_n18620# a_71281_n8397.t259 a_111063_n18620# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4599 a_104527_n4245# a_71281_n8397.t260 a_103997_n4245# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4600 VDD.t1928 VDD.t1927 VDD.t1928 VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4601 VSS.t1568 VSS.t1567 VSS.t1568 VSS.t475 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4602 VSS.t1566 VSS.t1565 VSS.t1566 VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4603 a_71281_n10073.t15 a_71281_n10073.t14 VDD.t348 VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4604 VSS.t1564 VSS.t1563 VSS.t1564 VSS.t309 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4605 a_41487_n14213# a_31953_n19727.t277 a_40965_n14213# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4606 a_48391_n30339# a_39179_n19595.t0 a_47819_n36322.t4 VSS.t339 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4607 VDD.t4845 a_52635_34067.t195 a_52635_49681.t108 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4608 VDD.t1926 VDD.t1925 VDD.t1926 VDD.t1322 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4609 a_38619_n7136# a_31953_n19727.t278 a_38097_n7136# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4610 VDD.t1924 VDD.t1923 VDD.t1924 VDD.t1049 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4611 VSS.t1562 VSS.t1561 VSS.t1562 VSS.t1222 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4612 VSS.t1560 VSS.t1559 VSS.t1560 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4613 VSS.t1558 VSS.t1557 VSS.t1558 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4614 a_84017_n17715.t5 a_81205_n14095.t5 a_95443_13546# VDD.t498 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4615 a_83683_10448# a_83153_10448.t4 a_83153_10448.t5 VDD.t2774 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4616 a_60677_10448.t2 a_47991_4421.t1 a_60109_12380# VDD.t664 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4617 VDD.t435 a_71281_n8397.t12 a_71281_n8397.t13 VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4618 VSS.t1556 VSS.t1555 VSS.t1556 VSS.t487 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4619 VSS.t1554 VSS.t1553 VSS.t1554 VSS.t704 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4620 a_49755_11614# a_47819_10448.t17 VDD.t513 VDD.t508 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4621 VDD.t1922 VDD.t1921 VDD.t1922 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4622 VSS.t1552 VSS.t1551 VSS.t1552 VSS.t609 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4623 VDD.t1920 VDD.t1919 VDD.t1920 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4624 VDD.t1918 VDD.t1916 VDD.t1918 VDD.t1917 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4625 a_33249_48695.t129 a_33379_34007.t65 a_33249_34067.t45 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4626 a_36530_n29181# a_30152_n36322.t18 VDD.t4769 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4627 VSS.t1550 VSS.t1549 VSS.t1550 VSS.t484 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4628 VDD.t1915 VDD.t1914 VDD.t1915 VDD.t49 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4629 a_108636_n33224# a_106830_n36382.t23 a_106676_n30339.t3 VDD.t1540 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4630 VSS.t1548 VSS.t1547 VSS.t1548 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4631 VSS.t1546 VSS.t1545 VSS.t1546 VSS.t615 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4632 VSS.t1544 VSS.t1543 VSS.t1544 VSS.t568 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4633 a_33249_35053.t119 a_35502_25545.t77 VSS.t48 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4634 VDD.t1913 VDD.t1912 VDD.t1913 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4635 VDD.t1911 VDD.t1910 VDD.t1911 VDD.t568 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4636 VSS.t1542 VSS.t1541 VSS.t1542 VSS.t650 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4637 VDD.t1909 VDD.t1908 VDD.t1909 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4638 a_33249_48695.t76 a_33379_34917.t65 a_33249_35053.t62 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4639 VDD.t1907 VDD.t1906 VDD.t1907 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4640 a_33249_34067.t44 a_33379_34007.t66 a_33249_48695.t130 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4641 VSS.t1540 VSS.t1539 VSS.t1540 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4642 VDD.t1905 VDD.t1903 VDD.t1905 VDD.t1904 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4643 VSS.t8 a_35502_25545.t78 a_33249_35053.t118 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4644 a_84017_n17715.t2 a_81205_n14095.t6 a_95443_11614# VDD.t498 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4645 a_51711_n8932# a_50751_n19729.t267 a_51151_n8932# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4646 VDD.t1902 VDD.t1901 VDD.t1902 VDD.t780 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4647 VDD.t1900 VDD.t1899 VDD.t1900 VDD.t552 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4648 a_33249_34067.t43 a_33379_34007.t67 a_33249_48695.t131 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4649 a_51711_n18700# a_50751_n19729.t268 a_51151_n17803# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4650 VSS.t1538 VSS.t1536 VSS.t1538 VSS.t1537 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4651 VDD.t1898 VDD.t1897 VDD.t1898 VDD.t677 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4652 a_44885_n14213# a_31953_n19727.t279 a_44363_n15110# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4653 VDD.t1896 VDD.t1895 VDD.t1896 VDD.t674 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4654 VDD.t1894 VDD.t1892 VDD.t1894 VDD.t1893 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4655 a_83153_n36322.t1 a_32913_n8930.t1 a_85129_n27257# VSS.t285 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4656 VDD.t1891 VDD.t1890 VDD.t1891 VDD.t1505 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4657 VDD.t1889 VDD.t1888 VDD.t1889 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4658 a_95943_n18620# a_71281_n10073.t253 a_95105_n15905# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4659 VSS.t1535 VSS.t1534 VSS.t1535 VSS.t668 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4660 a_110225_n6960# a_71281_n8397.t261 a_109695_n7865# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4661 a_84547_n3340# a_71281_n10073.t254 a_83709_n2435# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4662 a_88271_n8770# a_71281_n10073.t255 a_87433_n8770# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4663 VDD.t1887 VDD.t1886 VDD.t1887 VDD.t353 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4664 a_52635_49681.t60 a_35922_19591.t138 OUT.t47 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4665 VDD.t1885 VDD.t1883 VDD.t1885 VDD.t1884 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4666 a_60845_n8932# a_50751_n19729.t269 a_60285_n8035# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4667 VDD.t1882 VDD.t1881 VDD.t1882 VDD.t12 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4668 VDD.t1880 VDD.t1879 VDD.t1880 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4669 VSS.t1533 VSS.t1532 VSS.t1533 VSS.t224 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4670 a_52635_34067.t36 a_35922_19591.t139 a_52635_48695.t26 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4671 VSS.t435 I1N.t11 a_72603_n10073# VSS.t433 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X4672 a_110225_n17715# a_71281_n8397.t262 a_109695_n21335# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4673 a_33249_34067.t42 a_33379_34007.t68 a_33249_48695.t132 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4674 a_50751_n19729.t33 a_50751_n19729.t32 VSS.t235 VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4675 VSS.t1531 VSS.t1530 VSS.t1531 VSS.t596 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4676 VDD.t1878 VDD.t1877 VDD.t1878 VDD.t1489 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4677 VSS.t1529 VSS.t1528 VSS.t1529 VSS.t650 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4678 VDD.t1876 VDD.t1875 VDD.t1876 VDD.t1164 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4679 VDD.t1874 VDD.t1873 VDD.t1874 VDD.t1505 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4680 VDD.t1872 VDD.t1871 VDD.t1872 VDD.t404 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4681 VSS.t1527 VSS.t1526 VSS.t1527 VSS.t98 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4682 a_93969_n14095# a_71281_n10073.t256 a_93131_n14095# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4683 a_52635_48695.t112 a_52635_34067.t196 VDD.t4844 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4684 a_83153_n36322.t4 a_83153_n35156.t19 a_85089_n35156# VDD.t1486 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4685 a_90935_5639# a_83153_11614.t19 a_51711_n12421.t0 VSS.t395 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4686 VSS.t1525 VSS.t1524 VSS.t1525 VSS.t641 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4687 a_52635_49681.t107 a_52635_34067.t197 VDD.t4843 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4688 VSS.t1523 VSS.t1522 VSS.t1523 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4689 a_94537_n15905# a_71281_n10073.t257 a_93969_n15905# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4690 a_71266_n4019.t0 I1N.t12 a_75585_n9297# VSS.t312 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X4691 VSS.t1521 VSS.t1520 VSS.t1521 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4692 VDD.t1870 VDD.t1869 VDD.t1870 VDD.t1188 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X4693 VDD.t1868 VDD.t1866 VDD.t1868 VDD.t1867 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4694 VDD.t1865 VDD.t1864 VDD.t1865 VDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4695 a_52635_49681.t106 a_52635_34067.t198 VDD.t4842 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4696 a_60285_n7138# a_50751_n19729.t270 a_59763_n8035# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4697 VDD.t1863 VDD.t1862 VDD.t1863 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4698 a_42413_n27257# a_41891_n29181.t9 a_41891_n29181.t10 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4699 VDD.t1861 VDD.t1860 VDD.t1861 VDD.t1481 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4700 VDD.t1859 VDD.t1858 VDD.t1859 VDD.t1127 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4701 VDD.t4841 a_52635_34067.t199 a_52635_48695.t111 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4702 VDD.t1857 VDD.t1856 VDD.t1857 VDD.t1489 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4703 a_35221_n16007# a_31953_n19727.t280 a_34347_n17801# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4704 VSS.t1519 VSS.t1518 VSS.t1519 VSS.t184 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4705 a_47819_10448.t8 a_47991_4421.t0 a_49795_7563# VSS.t337 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4706 VSS.t1517 VSS.t1516 VSS.t1517 VSS.t1064 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4707 a_67111_n19597# a_50751_n19729.t271 a_66551_n19597# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4708 a_101641_n3340# a_71281_n8397.t263 a_100803_n3340# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4709 a_66058_5639# a_64243_n1756.t1 a_65486_11614.t6 VSS.t376 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4710 VSS.t1515 VSS.t1514 VSS.t1515 VSS.t553 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4711 VDD.t1855 VDD.t1854 VDD.t1855 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4712 a_33249_34067.t41 a_33379_34007.t69 a_33249_48695.t133 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4713 OUT.t6 a_35502_24538.t53 a_33249_35053.t102 VSS.t196 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4714 VDD.t1853 VDD.t1852 VDD.t1853 VDD.t523 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4715 a_83153_n36322.t7 a_83153_n35156.t20 a_85089_n33224# VDD.t1486 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4716 a_33249_35053.t117 a_35502_25545.t79 VSS.t125 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4717 VSS.t1513 VSS.t1512 VSS.t1513 VSS.t168 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4718 VDD.t1851 VDD.t1849 VDD.t1851 VDD.t1850 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4719 a_89163_n36382.t2 a_94892_n29181.t18 a_96818_n27257# VSS.t352 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4720 a_31699_20742.t0 I1U.t5 a_30377_19942# VSS.t349 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X4721 a_52635_48695.t25 a_35922_19591.t140 a_52635_34067.t4 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4722 VDD.t1848 VDD.t1847 VDD.t1848 VDD.t1481 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4723 a_35221_n2651# a_31953_n19727.t281 a_34699_n3548# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4724 VDD.t1846 VDD.t1845 VDD.t1846 VDD.t1112 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4725 VDD.t1844 VDD.t1843 VDD.t1844 VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4726 VDD.t1842 VDD.t1840 VDD.t1842 VDD.t1841 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4727 VDD.t1839 VDD.t1838 VDD.t1839 VDD.t120 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4728 VSS.t1511 VSS.t1510 VSS.t1511 VSS.t332 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4729 VSS.t3644 a_94892_4481.t22 a_95414_4481# VSS.t1037 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4730 VDD.t1837 VDD.t1836 VDD.t1837 VDD.t551 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4731 a_33249_48695.t211 a_31699_20742.t201 VDD.t223 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4732 a_114516_n35156# a_103997_n8770.t11 a_106809_n5150.t3 VDD.t536 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4733 a_63683_n13318# a_50751_n19729.t272 a_63161_n13318# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4734 VSS.t1509 VSS.t1508 VSS.t1509 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4735 a_52635_49681.t61 a_35922_19591.t141 OUT.t46 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4736 a_57977_n6241# a_50751_n19729.t273 a_57417_n6241# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4737 VSS.t1507 VSS.t1506 VSS.t1507 VSS.t421 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4738 VDD.t1835 VDD.t1834 VDD.t1835 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4739 VDD.t1833 VDD.t1832 VDD.t1833 VDD.t55 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4740 VSS.t1505 VSS.t1504 VSS.t1505 VSS.t618 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4741 VDD.t1831 VDD.t1830 VDD.t1831 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4742 a_38619_n19595# a_31953_n19727.t282 a_38097_n19595# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4743 VSS.t1503 VSS.t1502 VSS.t1503 VSS.t401 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4744 VSS.t1501 VSS.t1500 VSS.t1501 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4745 VDD.t224 a_31699_20742.t202 a_33249_48695.t210 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4746 a_52635_48695.t24 a_35922_19591.t142 a_52635_34067.t6 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4747 a_31699_20742.t20 a_31699_20742.t19 VDD.t29 VDD.t18 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4748 a_51151_n5344# a_50751_n19729.t274 a_31284_4481.t0 VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4749 VDD.t1829 VDD.t1828 VDD.t1829 VDD.t568 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4750 VDD.t1827 VDD.t1826 VDD.t1827 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4751 a_88839_n1530# a_71281_n10073.t258 a_88271_n1530# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4752 VSS.t1499 VSS.t1498 VSS.t1499 VSS.t834 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4753 a_95943_n3340# a_71281_n10073.t259 a_95105_n2435# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4754 VSS.t1497 VSS.t1496 VSS.t1497 VSS.t1025 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4755 a_110225_n21335# a_71281_n8397.t264 a_109695_n21335# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4756 VDD.t1825 VDD.t1823 VDD.t1825 VDD.t1824 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4757 a_77747_n30339# a_77225_n29181.t18 a_71496_n36382.t4 VSS.t379 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4758 a_50751_n19729.t31 a_50751_n19729.t30 VSS.t234 VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4759 VDD.t1822 VDD.t1820 VDD.t1822 VDD.t1821 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4760 VDD.t1819 VDD.t1817 VDD.t1819 VDD.t1818 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4761 VSS.t1495 VSS.t1494 VSS.t1495 VSS.t171 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4762 VDD.t1816 VDD.t1815 VDD.t1816 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4763 VSS.t1493 VSS.t1492 VSS.t1493 VSS.t151 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4764 a_114516_n33224# a_103997_n8770.t12 a_106809_n5150.t1 VDD.t536 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4765 VDD.t1814 VDD.t1813 VDD.t1814 VDD.t55 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4766 a_46879_n13316# a_31953_n19727.t283 a_46319_n12419# VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4767 a_48391_7563# a_47991_5507.t1 a_47819_11614.t4 VSS.t339 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4768 VSS.t124 a_35502_25545.t80 a_33249_35053.t116 VSS.t33 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4769 VSS.t1491 VSS.t1490 VSS.t1491 VSS.t260 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4770 VDD.t1812 VDD.t1811 VDD.t1812 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4771 VSS.t1489 VSS.t1488 VSS.t1489 VSS.t154 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4772 VDD.t494 a_47819_n36322.t18 a_55601_n28415# VSS.t307 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4773 VSS.t1487 VSS.t1486 VSS.t1487 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4774 VDD.t1810 VDD.t1809 VDD.t1810 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4775 VDD.t1808 VDD.t1807 VDD.t1808 VDD.t535 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4776 a_93969_n4245# a_71281_n10073.t260 a_93131_n4245# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4777 VDD.t1806 VDD.t1805 VDD.t1806 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4778 VDD.t1804 VDD.t1803 VDD.t1804 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4779 a_32913_n16904# a_31953_n19727.t284 a_32353_n15110# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4780 VDD.t1802 VDD.t1801 VDD.t1802 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4781 a_33249_34067.t40 a_33379_34007.t70 a_33249_48695.t134 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4782 a_60080_n27257# a_59558_n29181.t7 a_59558_n29181.t8 VSS.t397 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4783 VSS.t1485 VSS.t1484 VSS.t1485 VSS.t158 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4784 a_42047_n8930# a_31953_n19727.t285 a_41487_n8930# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4785 VDD.t1800 VDD.t1798 VDD.t1800 VDD.t1799 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4786 VDD.t1797 VDD.t1795 VDD.t1797 VDD.t1796 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4787 VDD.t1794 VDD.t1793 VDD.t1794 VDD.t1081 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4788 VDD.t1792 VDD.t1791 VDD.t1792 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4789 VDD.t1790 VDD.t1789 VDD.t1790 VDD.t1424 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4790 VDD.t1788 VDD.t1786 VDD.t1788 VDD.t1787 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4791 a_47753_n1754# a_31953_n19727.t286 a_45445_n1754# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4792 a_71281_n8397.t11 a_71281_n8397.t10 VDD.t433 VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4793 a_71496_n36382.t5 a_77225_n29181.t19 a_79151_n29181# VSS.t380 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4794 OUT.t45 a_35922_19591.t143 a_52635_49681.t62 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4795 a_33249_35053.t63 a_33379_34917.t66 a_33249_48695.t77 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4796 VDD.t4782 a_83153_n36322.t19 a_90935_n29181# VSS.t455 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4797 a_102756_10448# a_100820_10448.t16 VDD.t372 VDD.t298 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4798 VSS.t123 a_35502_25545.t81 a_33249_35053.t115 VSS.t39 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4799 a_95414_4481# a_94892_4481.t4 a_94892_4481.t5 VSS.t998 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4800 VDD.t1785 VDD.t1784 VDD.t1785 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4801 a_40613_n17801# a_31953_n19727.t287 a_40053_n17801# VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4802 VDD.t28 a_31699_20742.t17 a_31699_20742.t18 VDD.t27 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4803 VDD.t4840 a_52635_34067.t200 a_52635_48695.t110 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4804 VDD.t1783 VDD.t1782 VDD.t1783 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4805 a_65117_n14215# a_50751_n19729.t275 a_64595_n14215# VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4806 VSS.t1483 VSS.t1482 VSS.t1483 VSS.t947 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4807 VDD.t1781 VDD.t1779 VDD.t1781 VDD.t1780 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4808 VSS.t1481 VSS.t1480 VSS.t1481 VSS.t475 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4809 VSS.t1479 VSS.t1478 VSS.t1479 VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4810 a_63683_n4447# a_50751_n19729.t276 a_63161_n4447# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4811 VSS.t1477 VSS.t1476 VSS.t1477 VSS.t498 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4812 VDD.t1778 VDD.t1777 VDD.t1778 VDD.t1408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4813 VSS.t1475 VSS.t1474 VSS.t1475 VSS.t588 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4814 a_59411_n14215# a_50751_n19729.t277 a_58851_n14215# VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4815 VSS.t1473 VSS.t1472 VSS.t1473 VSS.t163 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4816 VDD.t1776 VDD.t1775 VDD.t1776 VDD.t1424 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4817 a_50751_n19729.t29 a_50751_n19729.t28 VSS.t233 VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4818 VSS.t1471 VSS.t1470 VSS.t1471 VSS.t509 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4819 VDD.t1774 VDD.t1773 VDD.t1774 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4820 VSS.t1469 VSS.t1468 VSS.t1469 VSS.t137 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4821 VSS.t1467 VSS.t1465 VSS.t1467 VSS.t1466 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4822 a_71281_n8397.t9 a_71281_n8397.t8 VDD.t431 VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4823 VSS.t1464 VSS.t1463 VSS.t1464 VSS.t283 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4824 VDD.t1772 VDD.t1771 VDD.t1772 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4825 a_60285_n12421# a_50751_n19729.t278 VSS.t275 VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4826 a_89033_n35156.t4 a_89163_n36382.t20 a_90969_n35156# VDD.t550 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4827 a_33249_34067.t39 a_33379_34007.t71 a_33249_48695.t135 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4828 a_57417_n18700# a_50751_n19729.t279 a_56895_n19597# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4829 VSS.t1462 VSS.t1461 VSS.t1462 VSS.t1077 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X4830 VSS.t1460 VSS.t1459 VSS.t1460 VSS.t150 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4831 a_83141_n1530# a_71281_n10073.t261 a_82573_n1530# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4832 a_35502_25545.t23 a_35502_25545.t22 VSS.t203 VSS.t5 nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X4833 VSS.t1458 VSS.t1457 VSS.t1458 VSS.t1360 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4834 VSS.t1456 VSS.t1455 VSS.t1456 VSS.t568 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4835 VDD.t1770 VDD.t1769 VDD.t1770 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4836 VDD.t1768 VDD.t1767 VDD.t1768 VDD.t1049 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4837 VDD.t1766 VDD.t1765 VDD.t1766 VDD.t833 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4838 VDD.t1764 VDD.t1763 VDD.t1764 VDD.t1052 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4839 VSS.t1454 VSS.t1453 VSS.t1454 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4840 a_60845_n4447# a_50751_n19729.t280 a_60285_n3550# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4841 VDD.t1762 VDD.t1761 VDD.t1762 VDD.t1408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4842 a_100235_n1530# a_71281_n8397.t265 a_99667_n1530# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4843 VSS.t1452 VSS.t1451 VSS.t1452 VSS.t464 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4844 VDD.t1760 VDD.t1759 VDD.t1760 VDD.t434 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4845 a_54197_5639# a_47819_11614.t17 VDD.t504 VSS.t306 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4846 a_33249_48695.t209 a_31699_20742.t203 VDD.t225 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4847 a_52635_49681.t105 a_52635_34067.t201 VDD.t4839 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4848 VDD.t1758 VDD.t1757 VDD.t1758 VDD.t1373 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4849 VDD.t1756 VDD.t1755 VDD.t1756 VDD.t1370 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4850 VDD.t329 a_30152_10448.t15 a_30682_13546# VDD.t326 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4851 VDD.t1754 VDD.t1753 VDD.t1754 VDD.t336 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4852 a_89033_n36322.t2 a_89163_n36382.t21 a_90969_n33224# VDD.t550 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4853 a_78344_10448.t1 a_65658_4421.t2 a_77776_12380# VDD.t3570 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4854 a_53699_11614.t1 a_53829_10388.t21 a_55635_12380# VDD.t3747 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4855 VSS.t1450 VSS.t1449 VSS.t1450 VSS.t537 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4856 a_96849_13546# a_83325_4421.t1 a_84017_n17715.t3 VDD.t499 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4857 VDD.t1752 VDD.t1751 VDD.t1752 VDD.t1365 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4858 VSS.t1448 VSS.t1447 VSS.t1448 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4859 a_88271_n7865# a_71281_n10073.t262 a_87433_n7865# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4860 VDD.t1750 VDD.t1749 VDD.t1750 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4861 a_101641_n17715# a_71281_n8397.t266 a_43010_n36322.t0 VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4862 a_87433_n14095# a_71281_n10073.t263 a_86903_n14095.t2 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4863 VDD.t1748 VDD.t1746 VDD.t1748 VDD.t1747 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4864 a_101641_n15000# a_71281_n8397.t267 a_100803_n15000# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4865 VSS.t1446 VSS.t1445 VSS.t1446 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4866 VDD.t1745 VDD.t1744 VDD.t1745 VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4867 a_111631_n21335# a_71281_n8397.t268 a_111063_n21335# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4868 VDD.t1743 VDD.t1742 VDD.t1743 VDD.t1373 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4869 VDD.t1741 VDD.t1740 VDD.t1741 VDD.t1370 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4870 VDD.t330 a_30152_10448.t16 a_30682_11614# VDD.t326 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4871 VDD.t1739 VDD.t1738 VDD.t1739 VDD.t1354 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4872 VSS.t1444 VSS.t1443 VSS.t1444 VSS.t537 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4873 VDD.t1737 VDD.t1736 VDD.t1737 VDD.t1365 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4874 VSS.t1442 VSS.t1441 VSS.t1442 VSS.t795 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4875 a_96849_11614# a_83325_4421.t1 a_84017_n17715.t4 VDD.t499 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4876 VDD.t1735 VDD.t1734 VDD.t1735 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4877 VDD.t1733 VDD.t1732 VDD.t1733 VDD.t1349 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4878 VDD.t485 a_71281_n8397.t269 a_112199_n1530# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4879 VSS.t122 a_35502_25545.t82 a_33249_35053.t114 VSS.t37 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4880 VSS.t1440 VSS.t1439 VSS.t1440 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4881 a_33249_34067.t4 a_35502_24538.t54 a_52635_34067.t60 VSS.t196 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4882 a_48313_n17801# a_31953_n19727.t288 a_47753_n16904# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4883 a_112559_n29181.t4 a_112559_n29181.t3 a_114485_n30339# VSS.t409 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4884 a_33249_48695.t208 a_31699_20742.t204 VDD.t226 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4885 VDD.t1731 VDD.t1730 VDD.t1731 VDD.t305 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4886 VSS.t1438 VSS.t1437 VSS.t1438 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4887 VSS.t1436 VSS.t1435 VSS.t1436 VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4888 VSS.t1434 VSS.t1433 VSS.t1434 VSS.t21 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4889 VDD.t227 a_31699_20742.t205 a_33249_48695.t207 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4890 a_58851_n17803# a_50751_n19729.t281 a_58329_n18700# VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4891 VSS.t1432 VSS.t1430 VSS.t1432 VSS.t1431 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4892 VSS.t1429 VSS.t1428 VSS.t1429 VSS.t349 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4893 VDD.t228 a_31699_20742.t206 a_33249_48695.t206 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4894 VDD.t1729 VDD.t1728 VDD.t1729 VDD.t1354 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4895 VDD.t1727 VDD.t1726 VDD.t1727 VDD.t554 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4896 a_52635_48695.t109 a_52635_34067.t202 VDD.t4838 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4897 VDD.t1725 VDD.t1724 VDD.t1725 VDD.t1015 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4898 a_101641_n3340# a_71281_n8397.t270 a_100803_n2435# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4899 VDD.t1723 VDD.t1722 VDD.t1723 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4900 VDD.t1721 VDD.t1720 VDD.t1721 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4901 VDD.t1719 VDD.t1718 VDD.t1719 VDD.t1349 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4902 a_36008_n27257.t0 a_30152_n36322.t19 a_37934_n30339# VSS.t281 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4903 a_107339_n17715# a_71281_n8397.t271 a_60677_n36322.t0 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4904 a_47991_5507.t0 a_50751_n19729.t282 a_57417_n1756# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4905 a_37934_7563# a_30152_11614.t16 a_30324_4421.t0 VSS.t282 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4906 a_33249_48695.t205 a_31699_20742.t207 VDD.t229 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4907 a_52635_48695.t108 a_52635_34067.t203 VDD.t4837 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4908 a_107339_n15000# a_71281_n8397.t272 a_106501_n15000# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4909 VSS.t1427 VSS.t1425 VSS.t1427 VSS.t1426 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4910 VSS.t1424 VSS.t1423 VSS.t1424 VSS.t531 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4911 VSS.t1422 VSS.t1421 VSS.t1422 VSS.t393 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4912 VSS.t1420 VSS.t1419 VSS.t1420 VSS.t733 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4913 a_65658_4421.t0 a_65486_11614.t23 a_71864_4481# VSS.t424 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4914 VDD.t1717 VDD.t1716 VDD.t1717 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4915 VDD.t1715 VDD.t1713 VDD.t1715 VDD.t1714 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4916 VDD.t1712 VDD.t1710 VDD.t1712 VDD.t1711 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4917 VSS.t1418 VSS.t1417 VSS.t1418 VSS.t495 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4918 VSS.t1416 VSS.t1415 VSS.t1416 VSS.t289 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4919 VDD.t1709 VDD.t1707 VDD.t1709 VDD.t1708 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4920 a_71366_11614.t1 a_71496_10388.t20 a_73302_12380# VDD.t352 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4921 VDD.t1706 VDD.t1705 VDD.t1706 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4922 VDD.t1704 VDD.t1703 VDD.t1704 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4923 VDD.t1702 VDD.t1701 VDD.t1702 VDD.t64 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4924 VDD.t1700 VDD.t1699 VDD.t1700 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4925 a_38097_n5342.t2 a_100992_n29313.t1 a_101392_n27257# VSS.t332 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4926 a_101641_n20430# a_71281_n8397.t273 a_100803_n20430# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4927 VDD.t1698 VDD.t1697 VDD.t1698 VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4928 VSS.t1414 VSS.t1413 VSS.t1414 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4929 VDD.t1696 VDD.t1695 VDD.t1696 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4930 VSS.t1412 VSS.t1411 VSS.t1412 VSS.t378 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4931 VSS.t1410 VSS.t1409 VSS.t1410 VSS.t1034 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4932 VDD.t1694 VDD.t1693 VDD.t1694 VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4933 VSS.t1408 VSS.t1407 VSS.t1408 VSS.t478 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4934 a_43817_n28415# a_41891_n29181.t20 VSS.t373 VSS.t158 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4935 VDD.t230 a_31699_20742.t208 a_33249_48695.t204 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4936 VDD.t4836 a_52635_34067.t204 a_52635_48695.t107 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4937 VDD.t26 a_31699_20742.t15 a_31699_20742.t16 VDD.t25 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4938 a_106809_n6055.t0 a_71281_n8397.t274 a_106501_n9675# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4939 VSS.t1406 VSS.t1405 VSS.t1406 VSS.t687 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4940 VSS.t1404 VSS.t1403 VSS.t1404 VSS.t944 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4941 a_33249_48695.t203 a_31699_20742.t209 VDD.t231 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4942 a_52635_49681.t104 a_52635_34067.t205 VDD.t4835 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4943 VDD.t1692 VDD.t1691 VDD.t1692 VDD.t20 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4944 VSS.t1402 VSS.t1401 VSS.t1402 VSS.t1237 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4945 VDD.t1690 VDD.t1689 VDD.t1690 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4946 a_49795_n28415# a_47991_n29313.t0 a_38097_n16007.t1 VSS.t338 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4947 a_33249_48695.t202 a_31699_20742.t210 VDD.t232 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4948 a_100820_n35156.t11 a_100820_n35156.t10 a_102756_n34390# VDD.t532 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4949 a_50751_n19729.t27 a_50751_n19729.t26 VSS.t232 VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4950 a_41891_4481.t1 a_30324_4421.t1 a_43848_13546# VDD.t287 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4951 VDD.t1688 VDD.t1687 VDD.t1688 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4952 VSS.t1400 VSS.t1399 VSS.t1400 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4953 VSS.t1398 VSS.t1397 VSS.t1398 VSS.t558 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4954 VDD.t1686 VDD.t1685 VDD.t1686 VDD.t1658 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4955 VDD.t1684 VDD.t1683 VDD.t1684 VDD.t425 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4956 VDD.t1682 VDD.t1681 VDD.t1682 VDD.t341 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4957 VSS.t1396 VSS.t1395 VSS.t1396 VSS.t495 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4958 a_73268_n27257# a_65486_n36322.t21 a_65658_n29313.t0 VSS.t154 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4959 VDD.t1680 VDD.t1679 VDD.t1680 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4960 VSS.t1394 VSS.t1393 VSS.t1394 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4961 VSS.t1392 VSS.t1391 VSS.t1392 VSS.t98 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4962 a_72596_n3060# a_71266_n4019.t0 a_50751_n19729.t73 VDD.t994 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X4963 VSS.t1390 VSS.t1389 VSS.t1390 VSS.t297 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4964 VSS.t1388 VSS.t1387 VSS.t1388 VSS.t394 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4965 VSS.t1386 VSS.t1384 VSS.t1386 VSS.t1385 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4966 a_105365_n6960# a_71281_n8397.t275 a_104527_n6960# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4967 VSS.t1383 VSS.t1382 VSS.t1383 VSS.t263 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4968 a_60285_n6241# a_50751_n19729.t283 a_59763_n6241# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4969 VDD.t1678 VDD.t1677 VDD.t1678 VDD.t423 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4970 VSS.t1381 VSS.t1380 VSS.t1381 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4971 VDD.t1676 VDD.t1675 VDD.t1676 VDD.t301 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4972 VDD.t1674 VDD.t1673 VDD.t1674 VDD.t439 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4973 VSS.t1379 VSS.t1378 VSS.t1379 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4974 VSS.t231 a_50751_n19729.t24 a_50751_n19729.t25 VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4975 a_107339_n20430# a_71281_n8397.t276 a_106501_n20430# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4976 a_95943_n15000# a_71281_n10073.t264 a_95105_n14095# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4977 a_105933_n1530# a_71281_n8397.t277 a_105365_n1530# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4978 a_34347_n19595# a_31953_n19727.t289 a_33787_n19595# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4979 VDD.t530 a_100820_n35156.t18 a_101350_n34390# VDD.t529 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4980 a_52635_49681.t63 a_35922_19591.t144 OUT.t44 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4981 VDD.t1672 VDD.t1671 VDD.t1672 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4982 a_33249_48695.t201 a_31699_20742.t211 VDD.t233 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4983 a_41891_4481.t2 a_30324_4421.t1 a_43848_11614# VDD.t287 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4984 VDD.t1670 VDD.t1669 VDD.t1670 VDD.t965 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4985 a_107230_12380# a_106830_10388.t18 a_86903_n14095.t1 VDD.t522 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4986 VDD.t1668 VDD.t1667 VDD.t1668 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4987 VSS.t1377 VSS.t1376 VSS.t1377 VSS.t381 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4988 a_47991_n29313.t0 a_47819_n36322.t19 a_54197_n30339# VSS.t304 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4989 VSS.t1375 VSS.t1374 VSS.t1375 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4990 VSS.t1373 VSS.t1372 VSS.t1373 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4991 VSS.t13 a_35502_25545.t83 a_33249_35053.t113 VSS.t12 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4992 VDD.t4834 a_52635_34067.t206 a_52635_49681.t103 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4993 a_75585_n10973# I1N.t13 VSS.t436 VSS.t430 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X4994 VDD.t1666 VDD.t1664 VDD.t1666 VDD.t1665 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X4995 a_82573_n19525# a_71281_n10073.t265 a_81735_n19525# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4996 a_111063_n4245# a_71281_n8397.t278 a_110225_n4245# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4997 a_52585_n8035# a_50751_n19729.t284 a_52063_n8035# VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4998 a_33249_48695.t200 a_31699_20742.t212 VDD.t234 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4999 a_65677_n7138# a_50751_n19729.t285 a_66551_n5344# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5000 a_63683_n12421# a_50751_n19729.t286 a_63161_n13318# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5001 VDD.t1663 VDD.t1662 VDD.t1663 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5002 a_54579_n8932# a_50751_n19729.t287 a_54019_n8035# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5003 VDD.t1661 VDD.t1660 VDD.t1661 VDD.t293 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5004 VSS.t1371 VSS.t1370 VSS.t1371 VSS.t1104 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5005 VSS.t1369 VSS.t1368 VSS.t1369 VSS.t287 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5006 VDD.t1659 VDD.t1657 VDD.t1659 VDD.t1658 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5007 VSS.t1367 VSS.t1366 VSS.t1367 VSS.t571 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5008 VSS.t71 a_31953_n19727.t22 a_31953_n19727.t23 VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5009 a_94537_n14095# a_71281_n10073.t266 a_93969_n14095# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5010 a_30324_n29313.t0 a_30152_n36322.t20 a_36530_n27257# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5011 VDD.t1656 VDD.t1655 VDD.t1656 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5012 VSS.t1365 VSS.t1364 VSS.t1365 VSS.t1253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5013 VDD.t1654 VDD.t1652 VDD.t1654 VDD.t1653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5014 a_35781_n13316# a_31953_n19727.t290 a_35221_n12419# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5015 VSS.t1363 VSS.t1362 VSS.t1363 VSS.t868 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5016 VDD.t1651 VDD.t1650 VDD.t1651 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5017 VDD.t1649 VDD.t1648 VDD.t1649 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5018 a_33249_34067.t117 a_35502_25545.t84 VSS.t11 VSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5019 VDD.t1647 VDD.t1646 VDD.t1647 VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5020 a_36562_n34390# a_36162_n36382.t20 a_36032_n35156.t3 VDD.t680 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5021 a_33249_34067.t38 a_33379_34007.t72 a_33249_48695.t136 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5022 VSS.t1361 VSS.t1359 VSS.t1361 VSS.t1360 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5023 VSS.t1358 VSS.t1357 VSS.t1358 VSS.t289 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5024 a_55601_n29181# a_47819_n36322.t20 a_39179_n19595.t0 VSS.t305 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5025 VSS.t1356 VSS.t1355 VSS.t1356 VSS.t224 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5026 a_101641_n18620# a_71281_n8397.t279 a_100803_n15905# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5027 VSS.t1354 VSS.t1353 VSS.t1354 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5028 VDD.t1645 VDD.t1644 VDD.t1645 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5029 a_90245_n6055# a_71281_n10073.t267 a_89715_n5150.t0 VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5030 VSS.t1352 VSS.t1351 VSS.t1352 VSS.t558 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5031 VSS.t1350 VSS.t1349 VSS.t1350 VSS.t976 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5032 a_47753_n17801# a_31953_n19727.t291 a_47231_n18698# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5033 a_66058_n28415# a_45445_n19595.t1 a_65486_n36322.t7 VSS.t376 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5034 a_52635_48695.t106 a_52635_34067.t207 VDD.t4833 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5035 VDD.t1643 VDD.t1641 VDD.t1643 VDD.t1642 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5036 VDD.t1640 VDD.t1639 VDD.t1640 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5037 VDD.t1638 VDD.t1637 VDD.t1638 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5038 VSS.t405 a_59558_4481.t17 a_60080_7563# VSS.t401 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5039 VSS.t205 a_35502_25545.t20 a_35502_25545.t21 VSS.t129 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X5040 VSS.t1348 VSS.t1347 VSS.t1348 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5041 VSS.t1346 VSS.t1345 VSS.t1346 VSS.t891 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5042 VSS.t1344 VSS.t1343 VSS.t1344 VSS.t396 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5043 VDD.t1636 VDD.t1635 VDD.t1636 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5044 VSS.t1342 VSS.t1341 VSS.t1342 VSS.t537 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5045 a_32913_n14213# a_31953_n19727.t292 a_32353_n14213# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5046 VDD.t1634 VDD.t1633 VDD.t1634 VDD.t55 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5047 a_83153_10448.t2 a_83325_4421.t0 a_85129_7563# VSS.t308 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5048 VSS.t1340 VSS.t1339 VSS.t1340 VSS.t908 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5049 VSS.t1338 VSS.t1337 VSS.t1338 VSS.t877 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5050 a_38619_n1754# a_31953_n19727.t293 a_38097_n2651# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5051 VDD.t1632 VDD.t1631 VDD.t1632 VDD.t549 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5052 VSS.t1336 VSS.t1335 VSS.t1336 VSS.t868 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5053 VDD.t1630 VDD.t1629 VDD.t1630 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5054 VDD.t1628 VDD.t1627 VDD.t1628 VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5055 VDD.t1626 VDD.t1625 VDD.t1626 VDD.t1251 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5056 a_100992_4421.t0 a_100820_11614.t19 a_107198_4481# VSS.t153 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5057 VDD.t4832 a_52635_34067.t208 a_52635_48695.t105 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5058 a_53145_n19597# a_50751_n19729.t288 a_52585_n18700# VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5059 VDD.t1624 VDD.t1623 VDD.t1624 VDD.t994 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X5060 VSS.t1334 VSS.t1333 VSS.t1334 VSS.t1064 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5061 VDD.t1622 VDD.t1621 VDD.t1622 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5062 VDD.t1620 VDD.t1619 VDD.t1620 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5063 VSS.t1332 VSS.t1331 VSS.t1332 VSS.t837 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5064 VSS.t1330 VSS.t1329 VSS.t1330 VSS.t1222 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5065 VDD.t1618 VDD.t1617 VDD.t1618 VDD.t546 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5066 VDD.t1616 VDD.t1615 VDD.t1616 VDD.t521 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5067 a_33249_48695.t137 a_33379_34007.t73 a_33249_34067.t37 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5068 VDD.t1614 VDD.t1613 VDD.t1614 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5069 VDD.t1612 VDD.t1610 VDD.t1612 VDD.t1611 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5070 VSS.t1328 VSS.t1327 VSS.t1328 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5071 a_32088_13546# a_30152_10448.t17 VDD.t332 VDD.t303 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5072 VDD.t1609 VDD.t1608 VDD.t1609 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5073 a_84017_n16810.t1 a_71281_n10073.t268 a_83709_n13190# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5074 VDD.t235 a_31699_20742.t213 a_35502_24538.t7 VDD.t34 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5075 VSS.t9 a_35502_25545.t85 a_33249_35053.t112 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5076 a_107339_n18620# a_71281_n8397.t280 a_106501_n15905# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5077 a_33249_48695.t199 a_31699_20742.t214 VDD.t236 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5078 VSS.t1326 VSS.t1325 VSS.t1326 VSS.t522 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5079 VDD.t1607 VDD.t1606 VDD.t1607 VDD.t1251 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5080 VDD.t1605 VDD.t1604 VDD.t1605 VDD.t1209 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5081 VSS.t1324 VSS.t1323 VSS.t1324 VSS.t311 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5082 VSS.t1322 VSS.t1321 VSS.t1322 VSS.t615 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5083 a_33249_48695.t198 a_31699_20742.t215 VDD.t237 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5084 VSS.t1320 VSS.t1319 VSS.t1320 VSS.t795 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5085 VDD.t4790 a_83153_10448.t22 a_83683_12380# VDD.t3354 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5086 VDD.t1603 VDD.t1602 VDD.t1603 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5087 a_33249_48695.t197 a_31699_20742.t216 VDD.t238 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5088 VDD.t1601 VDD.t1600 VDD.t1601 VDD.t905 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5089 VDD.t1599 VDD.t1598 VDD.t1599 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5090 VDD.t1597 VDD.t1596 VDD.t1597 VDD.t893 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5091 VSS.t1318 VSS.t1317 VSS.t1318 VSS.t1253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5092 VSS.t1316 VSS.t1314 VSS.t1316 VSS.t1315 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5093 a_106830_10388.t7 a_86903_n14095.t8 a_114516_12380# VDD.t338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5094 a_32088_11614# a_30152_10448.t18 VDD.t333 VDD.t303 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5095 VDD.t1595 VDD.t1594 VDD.t1595 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5096 VDD.t1593 VDD.t1592 VDD.t1593 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5097 VSS.t1313 VSS.t1312 VSS.t1313 VSS.t531 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5098 VDD.t1591 VDD.t1590 VDD.t1591 VDD.t545 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5099 a_45445_n16904# a_31953_n19727.t294 a_44885_n16904# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5100 VSS.t1311 VSS.t1310 VSS.t1311 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5101 a_60845_n2653# a_50751_n19729.t289 a_60285_n2653# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5102 VSS.t1309 VSS.t1308 VSS.t1309 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5103 VSS.t1307 VSS.t1305 VSS.t1307 VSS.t1306 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5104 VSS.t1304 VSS.t1302 VSS.t1304 VSS.t1303 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5105 VSS.t1301 VSS.t1300 VSS.t1301 VSS.t576 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5106 VSS.t1299 VSS.t1298 VSS.t1299 VSS.t591 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5107 VDD.t1589 VDD.t1588 VDD.t1589 VDD.t1209 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5108 a_33787_n8930# a_31953_n19727.t295 a_32913_n5342.t1 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5109 VSS.t1297 VSS.t1296 VSS.t1297 VSS.t333 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5110 VDD.t1587 VDD.t1586 VDD.t1587 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5111 a_33249_48695.t78 a_33379_34917.t67 a_33249_35053.t64 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5112 VDD.t1585 VDD.t1584 VDD.t1585 VDD.t27 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5113 a_51711_n6241# a_50751_n19729.t290 a_51151_n4447# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5114 a_67462_n27257# a_45445_n19595.t1 a_44363_n16007.t2 VSS.t289 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5115 a_66551_n16906# a_50751_n19729.t291 a_66029_n16906# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5116 a_31699_20742.t14 a_31699_20742.t13 VDD.t24 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5117 VSS.t1295 VSS.t1293 VSS.t1295 VSS.t1294 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5118 VSS.t1292 VSS.t1291 VSS.t1292 VSS.t937 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5119 VDD.t1583 VDD.t1582 VDD.t1583 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5120 VDD.t1581 VDD.t1580 VDD.t1581 VDD.t1183 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5121 a_32353_n17801# a_31953_n19727.t296 a_31831_n17801# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5122 VSS.t117 a_31953_n19727.t297 a_44885_n8930# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5123 VDD.t1579 VDD.t1578 VDD.t1579 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5124 VDD.t4831 a_52635_34067.t209 a_52635_49681.t102 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5125 VSS.t1290 VSS.t1289 VSS.t1290 VSS.t834 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5126 VDD.t1577 VDD.t1576 VDD.t1577 VDD.t875 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5127 VDD.t1575 VDD.t1574 VDD.t1575 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5128 a_51711_n14215# a_50751_n19729.t292 a_51151_n13318# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5129 VDD.t1573 VDD.t1572 VDD.t1573 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5130 VSS.t1288 VSS.t1286 VSS.t1288 VSS.t1287 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5131 VSS.t1285 VSS.t1284 VSS.t1285 VSS.t490 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5132 VDD.t1571 VDD.t1569 VDD.t1571 VDD.t1570 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5133 VSS.t1283 VSS.t1282 VSS.t1283 VSS.t808 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5134 VDD.t1568 VDD.t1567 VDD.t1568 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5135 VDD.t1566 VDD.t1565 VDD.t1566 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5136 a_60285_n1756# a_50751_n19729.t293 VSS.t276 VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5137 VDD.t1564 VDD.t1563 VDD.t1564 VDD.t1177 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5138 a_33249_35053.t105 a_35502_24538.t55 OUT.t5 VSS.t184 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5139 VDD.t1562 VDD.t1561 VDD.t1562 VDD.t1195 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5140 a_52635_48695.t104 a_52635_34067.t210 VDD.t4830 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5141 VDD.t1560 VDD.t1559 VDD.t1560 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5142 a_52635_48695.t23 a_35922_19591.t145 a_52635_34067.t15 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5143 VSS.t1281 VSS.t1280 VSS.t1281 VSS.t908 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5144 VSS.t1279 VSS.t1278 VSS.t1279 VSS.t310 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5145 VDD.t1558 VDD.t1557 VDD.t1558 VDD.t852 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5146 VDD.t1556 VDD.t1555 VDD.t1556 VDD.t1183 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5147 a_36562_12380# a_36162_10388.t20 a_36032_11614.t2 VDD.t3423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5148 VSS.t1277 VSS.t1276 VSS.t1277 VSS.t760 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5149 VSS.t1275 VSS.t1274 VSS.t1275 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5150 VDD.t1554 VDD.t1553 VDD.t1554 VDD.t521 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5151 VDD.t1552 VDD.t1551 VDD.t1552 VDD.t60 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5152 a_33379_34917.t68 IN_NEG.t1 cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
X5153 a_42442_n34390# a_36032_n35156.t11 a_36162_n36382.t7 VDD.t560 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5154 a_33249_35053.t111 a_35502_25545.t86 VSS.t126 VSS.t37 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5155 VDD.t4829 a_52635_34067.t211 a_52635_48695.t103 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5156 VDD.t1550 VDD.t1548 VDD.t1550 VDD.t1549 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5157 VDD.t1547 VDD.t1546 VDD.t1547 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5158 a_61484_n28415# a_59558_n29181.t19 VSS.t3633 VSS.t399 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5159 a_110225_n6055# a_71281_n8397.t281 a_109695_n9675# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5160 a_39179_n8033# a_31953_n19727.t298 a_38619_n7136# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5161 a_96818_n30339# a_94892_n29181.t19 VSS.t361 VSS.t354 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5162 VDD.t1545 VDD.t1544 VDD.t1545 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5163 VDD.t1543 VDD.t1542 VDD.t1543 VDD.t1177 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5164 VDD.t1541 VDD.t1539 VDD.t1541 VDD.t1540 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5165 a_100820_n35156.t1 a_100992_n29313.t0 a_102796_n28415# VSS.t329 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5166 VDD.t1538 VDD.t1537 VDD.t1538 VDD.t1195 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5167 a_52585_n3550# a_50751_n19729.t294 a_52063_n3550# VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5168 VDD.t1536 VDD.t1535 VDD.t1536 VDD.t833 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5169 a_54019_n8035# a_50751_n19729.t295 a_53497_n8035# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5170 VDD.t1534 VDD.t1533 VDD.t1534 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5171 a_32353_n6239# a_31953_n19727.t299 a_31831_n7136# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5172 a_54579_n4447# a_50751_n19729.t296 a_54019_n3550# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5173 VSS.t1273 VSS.t1272 VSS.t1273 VSS.t528 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5174 VSS.t1271 VSS.t1270 VSS.t1271 VSS.t853 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5175 VDD.t1532 VDD.t1531 VDD.t1532 VDD.t78 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5176 VSS.t1269 VSS.t1268 VSS.t1269 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5177 a_31953_n19727.t21 a_31953_n19727.t20 VSS.t70 VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5178 VDD.t1530 VDD.t1529 VDD.t1530 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5179 VSS.t1267 VSS.t1266 VSS.t1267 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5180 a_33249_48695.t196 a_31699_20742.t217 VDD.t239 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5181 VDD.t1528 VDD.t1527 VDD.t1528 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5182 a_79151_n27257# a_77225_n29181.t20 VSS.t388 VSS.t381 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5183 OUT.t108 a_33379_34917.t0 cap_mim_2f0_m4m5_noshield c_width=9.8u c_length=9.8u
X5184 a_112199_n9675# a_71281_n8397.t282 a_111631_n9675# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5185 a_49755_10448# a_47819_10448.t18 VDD.t514 VDD.t508 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5186 VSS.t1265 VSS.t1264 VSS.t1265 VSS.t775 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5187 VDD.t1526 VDD.t1525 VDD.t1526 VDD.t425 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5188 VSS.t1263 VSS.t1262 VSS.t1263 VSS.t45 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X5189 VSS.t1261 VSS.t1260 VSS.t1261 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5190 a_33249_48695.t79 a_33379_34917.t69 a_33249_35053.t65 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5191 a_94537_n8770# a_71281_n10073.t269 a_93969_n8770# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5192 VDD.t1524 VDD.t1523 VDD.t1524 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5193 VDD.t1522 VDD.t1521 VDD.t1522 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5194 VSS.t1259 VSS.t1258 VSS.t1259 VSS.t814 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5195 a_63161_n5344.t1 a_64243_n1756.t1 a_66058_5639# VSS.t377 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5196 a_71342_7563.t3 a_71496_10388.t21 a_71896_13546# VDD.t353 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5197 a_89163_10388.t5 a_81205_n14095.t7 a_96849_12380# VDD.t500 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5198 VDD.t1520 VDD.t1519 VDD.t1520 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5199 VDD.t1518 VDD.t1517 VDD.t1518 VDD.t801 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5200 a_51151_n16906# a_50751_n19729.t297 a_50629_n17803# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5201 VDD.t1516 VDD.t1514 VDD.t1516 VDD.t1515 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5202 a_84017_n17715.t1 a_83325_4421.t1 a_95443_10448# VDD.t498 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5203 VDD.t490 a_30152_11614.t17 a_37934_5639# VSS.t281 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5204 VDD.t1513 VDD.t1511 VDD.t1513 VDD.t1512 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5205 VSS.t1257 VSS.t1255 VSS.t1257 VSS.t1256 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5206 a_42047_n19595# a_31953_n19727.t300 a_41487_n18698# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5207 a_83725_n27257# a_83325_n29313.t2 a_83153_n35156.t8 VSS.t287 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5208 VDD.t1510 VDD.t1509 VDD.t1510 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5209 a_77747_5639# a_77225_4481.t19 a_71496_10388.t3 VSS.t317 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5210 a_52635_48695.t22 a_35922_19591.t146 a_52635_34067.t18 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5211 VDD.t1508 VDD.t1507 VDD.t1508 VDD.t434 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5212 VDD.t1506 VDD.t1504 VDD.t1506 VDD.t1505 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5213 VSS.t1254 VSS.t1252 VSS.t1254 VSS.t1253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5214 a_90245_n6960# a_71281_n10073.t270 a_89407_n4245# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5215 a_52585_n19597# a_50751_n19729.t298 VSS.t277 VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5216 a_107198_n28415# a_100820_n36322.t18 VDD.t541 VSS.t335 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5217 VSS.t1251 VSS.t1250 VSS.t1251 VSS.t166 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5218 VDD.t1503 VDD.t1502 VDD.t1503 VDD.t423 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5219 VSS.t1249 VSS.t1248 VSS.t1249 VSS.t422 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5220 a_52635_49681.t64 a_35922_19591.t147 OUT.t43 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5221 VSS.t1247 VSS.t1246 VSS.t1247 VSS.t307 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5222 VSS.t170 a_71496_10388.t22 a_71896_11614# VDD.t353 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5223 a_59411_n8932# a_50751_n19729.t299 a_58851_n8932# VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5224 VDD.t1501 VDD.t1500 VDD.t1501 VDD.t321 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5225 VDD.t1499 VDD.t1498 VDD.t1499 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5226 a_52635_48695.t102 a_52635_34067.t212 VDD.t4828 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5227 VSS.t1245 VSS.t1243 VSS.t1245 VSS.t1244 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X5228 a_33249_48695.t80 a_33379_34917.t70 a_33249_35053.t66 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5229 VDD.t1497 VDD.t1496 VDD.t1497 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5230 VDD.t1495 VDD.t1493 VDD.t1495 VDD.t1494 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5231 VDD.t1492 VDD.t1491 VDD.t1492 VDD.t524 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5232 VDD.t1490 VDD.t1488 VDD.t1490 VDD.t1489 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5233 a_52635_48695.t101 a_52635_34067.t213 VDD.t4827 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5234 a_48951_4481.t1 a_47991_5507.t1 a_48391_7563# VSS.t340 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5235 VDD.t1487 VDD.t1485 VDD.t1487 VDD.t1486 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5236 a_66551_n8035# a_50751_n19729.t300 a_66029_n8035# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5237 a_32128_5639# a_30324_4421.t0 a_31284_4481.t2 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5238 a_88271_n1530# a_71281_n10073.t271 a_87433_n1530# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5239 VSS.t1242 VSS.t1241 VSS.t1242 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5240 VDD.t1484 VDD.t1483 VDD.t1484 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5241 VSS.t1240 VSS.t1239 VSS.t1240 VSS.t292 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5242 a_33249_48695.t81 a_33379_34917.t71 a_33249_35053.t67 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5243 VSS.t1238 VSS.t1236 VSS.t1238 VSS.t1237 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X5244 VSS.t1235 VSS.t1234 VSS.t1235 VSS.t166 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5245 VSS.t1233 VSS.t1232 VSS.t1233 VSS.t811 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5246 VSS.t1231 VSS.t1230 VSS.t1231 VSS.t740 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5247 a_60080_7563# a_59558_4481.t18 a_53829_10388.t5 VSS.t397 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5248 VDD.t1482 VDD.t1480 VDD.t1482 VDD.t1481 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5249 VSS.t1229 VSS.t1228 VSS.t1229 VSS.t259 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5250 VSS.t1227 VSS.t1226 VSS.t1227 VSS.t638 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5251 VDD.t1479 VDD.t1478 VDD.t1479 VDD.t1112 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5252 a_77225_4481.t10 a_65658_4421.t2 a_79182_13546# VDD.t1841 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5253 VSS.t1225 VSS.t1224 VSS.t1225 VSS.t772 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5254 a_100820_11614.t1 a_100820_10448.t17 a_102756_12380# VDD.t322 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5255 a_33249_48695.t138 a_33379_34007.t74 a_33249_34067.t36 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5256 VDD.t1477 VDD.t1476 VDD.t1477 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5257 a_53829_10388.t6 a_59558_4481.t19 a_61484_4481# VSS.t398 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5258 VSS.t1223 VSS.t1221 VSS.t1223 VSS.t1222 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5259 VDD.t1475 VDD.t1474 VDD.t1475 VDD.t1127 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5260 VSS.t1220 VSS.t1219 VSS.t1220 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5261 a_33249_34067.t35 a_33379_34007.t75 a_33249_48695.t139 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5262 VDD.t1473 VDD.t1472 VDD.t1473 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5263 a_35502_24538.t6 a_31699_20742.t218 VDD.t240 VDD.t32 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5264 a_40613_n13316# a_31953_n19727.t301 a_40053_n13316# VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5265 a_65677_n17803# a_50751_n19729.t301 a_66551_n16009# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5266 VSS.t1218 VSS.t1217 VSS.t1218 VSS.t423 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5267 a_35502_24538.t5 a_31699_20742.t219 VDD.t241 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5268 a_52635_48695.t100 a_52635_34067.t214 VDD.t4826 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5269 VDD.t4825 a_52635_34067.t215 a_52635_48695.t99 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5270 VSS.t1216 VSS.t1215 VSS.t1216 VSS.t856 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5271 a_100820_n35156.t9 a_100820_n35156.t8 a_102756_n36322# VDD.t532 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5272 a_35502_25545.t17 a_31699_20742.t220 VDD.t242 VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5273 a_40053_n14213# a_31953_n19727.t302 a_39531_n14213# VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5274 a_61484_6405# a_59558_4481.t20 VSS.t406 VSS.t399 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5275 VSS.t1214 VSS.t1213 VSS.t1214 VSS.t615 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5276 VSS.t1212 VSS.t1211 VSS.t1212 VSS.t690 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5277 VDD.t1471 VDD.t1470 VDD.t1471 VDD.t1112 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5278 VSS.t1210 VSS.t1209 VSS.t1210 VSS.t687 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5279 a_77225_4481.t9 a_65658_4421.t2 a_79182_11614# VDD.t1841 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5280 a_39179_n18698# a_31953_n19727.t303 a_38619_n18698# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5281 VSS.t1208 VSS.t1207 VSS.t1208 VSS.t792 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5282 a_33249_48695.t195 a_31699_20742.t221 VDD.t243 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5283 a_52635_49681.t65 a_35922_19591.t148 OUT.t42 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5284 VDD.t1469 VDD.t1468 VDD.t1469 VDD.t341 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5285 VDD.t1467 VDD.t1466 VDD.t1467 VDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5286 VDD.t1465 VDD.t1464 VDD.t1465 VDD.t536 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5287 VDD.t1463 VDD.t1462 VDD.t1463 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5288 VDD.t1461 VDD.t1460 VDD.t1461 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5289 a_44363_n16007.t1 a_65658_n29313.t0 a_66058_n29181# VSS.t377 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5290 VDD.t1459 VDD.t1458 VDD.t1459 VDD.t1127 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5291 VSS.t1206 VSS.t1205 VSS.t1206 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5292 VDD.t1457 VDD.t1456 VDD.t1457 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5293 VDD.t1455 VDD.t1454 VDD.t1455 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5294 VDD.t1453 VDD.t1452 VDD.t1453 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5295 a_87433_n8770# a_71281_n10073.t272 VDD.t384 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5296 VSS.t1204 VSS.t1203 VSS.t1204 VSS.t162 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5297 VSS.t1202 VSS.t1201 VSS.t1202 VSS.t676 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5298 VSS.t1200 VSS.t1199 VSS.t1200 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5299 a_60285_n18700# a_50751_n19729.t302 a_59763_n18700# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5300 VDD.t1451 VDD.t1450 VDD.t1451 VDD.t398 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5301 VDD.t1449 VDD.t1448 VDD.t1449 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5302 VDD.t1447 VDD.t1446 VDD.t1447 VDD.t439 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5303 a_38619_n16007# a_31953_n19727.t304 a_38097_n16007.t0 VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5304 VSS.t1198 VSS.t1197 VSS.t1198 VSS.t1157 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5305 VDD.t1445 VDD.t1444 VDD.t1445 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5306 VSS.t1196 VSS.t1195 VSS.t1196 VSS.t265 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5307 VSS.t1194 VSS.t1193 VSS.t1194 VSS.t293 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5308 a_113081_n29181# a_112559_n29181.t5 a_112559_n29181.t6 VSS.t410 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5309 VSS.t1192 VSS.t1191 VSS.t1192 VSS.t817 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X5310 VSS.t1190 VSS.t1189 VSS.t1190 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5311 VSS.t1188 VSS.t1187 VSS.t1188 VSS.t224 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5312 VDD.t1443 VDD.t1441 VDD.t1443 VDD.t1442 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5313 VDD.t1440 VDD.t1438 VDD.t1440 VDD.t1439 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5314 VSS.t1186 VSS.t1185 VSS.t1186 VSS.t378 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5315 VDD.t1437 VDD.t1436 VDD.t1437 VDD.t801 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5316 VDD.t1435 VDD.t1434 VDD.t1435 VDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5317 VDD.t531 a_100820_n35156.t19 a_101350_n36322# VDD.t529 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5318 a_85089_12380# a_83153_10448.t23 VDD.t4791 VDD.t1442 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5319 VDD.t1433 VDD.t1432 VDD.t1433 VDD.t1081 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5320 VSS.t1184 VSS.t1183 VSS.t1184 VSS.t160 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5321 a_33249_48695.t194 a_31699_20742.t222 VDD.t244 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5322 VDD.t1431 VDD.t1430 VDD.t1431 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5323 VSS.t1182 VSS.t1181 VSS.t1182 VSS.t319 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5324 VSS.t326 a_77225_4481.t20 a_77747_7563# VSS.t323 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5325 VSS.t1180 VSS.t1179 VSS.t1180 VSS.t795 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5326 a_47991_5507.t1 a_47819_11614.t18 a_54197_5639# VSS.t304 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5327 VSS.t1178 VSS.t1177 VSS.t1178 VSS.t653 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5328 a_54019_n3550# a_50751_n19729.t303 a_53497_n3550# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5329 VSS.t230 a_50751_n19729.t22 a_50751_n19729.t23 VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5330 a_33249_48695.t193 a_31699_20742.t223 VDD.t245 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5331 VSS.t1176 VSS.t1175 VSS.t1176 VSS.t145 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5332 a_95105_n19525# a_71281_n10073.t273 a_94537_n19525# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5333 a_33249_34067.t34 a_33379_34007.t76 a_33249_48695.t140 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5334 VSS.t1174 VSS.t1173 VSS.t1174 VSS.t671 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5335 VSS.t1172 VSS.t1171 VSS.t1172 VSS.t733 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5336 a_41660_19698# a_35502_24538.t56 a_41100_19698# VSS.t186 nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X5337 a_90245_n20430# a_71281_n10073.t274 a_89407_n19525# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5338 VSS.t1170 VSS.t1169 VSS.t1170 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5339 a_107339_n3340# a_71281_n8397.t283 a_106501_n3340# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5340 VDD.t1429 VDD.t1428 VDD.t1429 VDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5341 VDD.t1427 VDD.t1426 VDD.t1427 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5342 VDD.t1425 VDD.t1423 VDD.t1425 VDD.t1424 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5343 VDD.t1422 VDD.t1421 VDD.t1422 VDD.t1081 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5344 VDD.t1420 VDD.t1418 VDD.t1420 VDD.t1419 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5345 a_101641_n15000# a_71281_n8397.t284 a_100803_n14095# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5346 VSS.t1168 VSS.t1167 VSS.t1168 VSS.t681 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5347 a_45706_23609# a_35922_19591.t149 a_45138_23609# VDD.t402 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X5348 a_48313_n13316# a_31953_n19727.t305 a_47753_n12419# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5349 VDD.t1417 VDD.t1416 VDD.t1417 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5350 VDD.t1415 VDD.t1414 VDD.t1415 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5351 a_33249_34067.t116 a_35502_25545.t87 VSS.t134 VSS.t3 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5352 a_36562_n36322# a_36162_n36382.t21 a_36032_n36322.t3 VDD.t680 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5353 a_47753_n8930# a_31953_n19727.t306 VSS.t118 VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5354 VDD.t1413 VDD.t1412 VDD.t1413 VDD.t1206 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5355 VSS.t389 a_77225_n29181.t21 a_77747_n29181# VSS.t384 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5356 a_41487_n19595# a_31953_n19727.t307 VSS.t119 VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5357 VSS.t1166 VSS.t1165 VSS.t1166 VSS.t31 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5358 VDD.t1411 VDD.t1410 VDD.t1411 VDD.t1049 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5359 a_58851_n13318# a_50751_n19729.t304 a_58329_n14215# VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5360 a_42047_n8930# a_31953_n19727.t308 a_41487_n8033# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5361 VDD.t1409 VDD.t1407 VDD.t1409 VDD.t1408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5362 VDD.t1406 VDD.t1404 VDD.t1406 VDD.t1405 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5363 VSS.t1164 VSS.t1163 VSS.t1164 VSS.t213 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5364 VSS.t1162 VSS.t1161 VSS.t1162 VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5365 a_88839_n19525# a_71281_n10073.t275 a_88271_n19525# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5366 VSS.t1160 VSS.t1159 VSS.t1160 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5367 VSS.t1158 VSS.t1156 VSS.t1158 VSS.t1157 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5368 VSS.t1155 VSS.t1154 VSS.t1155 VSS.t748 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5369 a_106676_4481.t2 a_100820_11614.t20 a_108602_7563# VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5370 a_30324_4421.t0 a_30152_11614.t18 a_36530_7563# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5371 a_94537_n7865# a_71281_n10073.t276 a_93969_n7865# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5372 a_89715_n17715.t5 a_86903_n14095.t9 a_113110_13546# VDD.t336 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5373 VDD.t1403 VDD.t1402 VDD.t1403 VDD.t550 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5374 a_33249_48695.t141 a_33379_34007.t77 a_33249_34067.t33 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5375 VSS.t1153 VSS.t1152 VSS.t1153 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5376 VSS.t1151 VSS.t1150 VSS.t1151 VSS.t217 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5377 VDD.t246 a_31699_20742.t224 a_35502_24538.t4 VDD.t34 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5378 a_33249_48695.t192 a_31699_20742.t225 VDD.t247 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5379 a_52635_48695.t98 a_52635_34067.t216 VDD.t4824 VDD.t391 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5380 VSS.t69 a_31953_n19727.t18 a_31953_n19727.t19 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5381 VSS.t1149 VSS.t1148 VSS.t1149 VSS.t704 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5382 VDD.t1401 VDD.t1400 VDD.t1401 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5383 VSS.t1147 VSS.t1146 VSS.t1147 VSS.t1034 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5384 VSS.t1145 VSS.t1144 VSS.t1145 VSS.t158 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5385 VDD.t1399 VDD.t1398 VDD.t1399 VDD.t1049 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5386 VDD.t248 a_31699_20742.t226 a_35502_25545.t4 VDD.t25 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5387 a_66016_n34390# a_65486_n35156.t21 a_65486_n36322.t2 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5388 VDD.t1397 VDD.t1396 VDD.t1397 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5389 VDD.t1395 VDD.t1394 VDD.t1395 VDD.t925 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5390 VSS.t1143 VSS.t1142 VSS.t1143 VSS.t615 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5391 a_71342_n27257.t3 a_65486_n36322.t22 a_73268_n30339# VSS.t155 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5392 VDD.t1393 VDD.t1392 VDD.t1393 VDD.t1052 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5393 a_51711_n12421.t1 a_50751_n19729.t305 a_51151_n12421# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5394 VSS.t1141 VSS.t1140 VSS.t1141 VSS.t16 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5395 VSS.t1139 VSS.t1138 VSS.t1139 VSS.t193 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5396 a_61515_12380# a_53699_11614.t9 a_60677_10448.t4 VDD.t3013 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5397 VSS.t1137 VSS.t1136 VSS.t1137 VSS.t568 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5398 VSS.t1135 VSS.t1134 VSS.t1135 VSS.t338 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5399 a_107339_n15000# a_71281_n8397.t285 a_106501_n14095# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5400 a_89715_n17715.t3 a_86903_n14095.t10 a_113110_11614# VDD.t336 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5401 VDD.t1391 VDD.t1390 VDD.t1391 VDD.t510 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5402 VSS.t1133 VSS.t1132 VSS.t1133 VSS.t684 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5403 a_52635_34067.t57 a_35502_24538.t57 a_33249_34067.t3 VSS.t192 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5404 VSS.t1131 VSS.t1130 VSS.t1131 VSS.t763 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X5405 a_33249_48695.t142 a_33379_34007.t78 a_33249_34067.t32 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5406 a_44885_n19595# a_31953_n19727.t309 a_44363_n19595# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5407 VSS.t1129 VSS.t1128 VSS.t1129 VSS.t644 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5408 a_66551_n3550# a_50751_n19729.t306 a_66029_n3550# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5409 VDD.t1389 VDD.t1388 VDD.t1389 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5410 VSS.t1127 VSS.t1125 VSS.t1127 VSS.t1126 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5411 VSS.t1124 VSS.t1123 VSS.t1124 VSS.t337 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5412 VSS.t1122 VSS.t1121 VSS.t1122 VSS.t604 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5413 a_52635_48695.t21 a_35922_19591.t150 a_52635_34067.t44 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5414 a_83709_n9675# a_71281_n10073.t277 a_83141_n9675# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5415 a_32128_n30339# a_30324_n29313.t0 a_31284_n30339.t1 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5416 VDD.t1387 VDD.t1386 VDD.t1387 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5417 VDD.t1385 VDD.t1384 VDD.t1385 VDD.t293 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5418 a_53675_n30339.t2 a_47819_n36322.t21 a_55601_n27257# VSS.t307 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5419 VSS.t1120 VSS.t1119 VSS.t1120 VSS.t671 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5420 VDD.t1383 VDD.t1382 VDD.t1383 VDD.t1052 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5421 a_111631_n8770# a_71281_n8397.t286 a_111063_n8770# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5422 VSS.t1118 VSS.t1117 VSS.t1118 VSS.t56 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5423 VSS.t1116 VSS.t1115 VSS.t1116 VSS.t182 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5424 a_33249_48695.t191 a_31699_20742.t227 VDD.t249 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5425 a_48313_n7136# a_31953_n19727.t310 a_47753_n6239# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5426 a_89009_7563.t3 a_89163_10388.t19 a_89563_13546# VDD.t554 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5427 VDD.t1381 VDD.t1380 VDD.t1381 VDD.t910 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5428 VDD.t1379 VDD.t1377 VDD.t1379 VDD.t1378 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5429 a_33249_48695.t82 a_33379_34917.t72 a_33249_35053.t68 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5430 VSS.t419 a_53829_10388.t22 a_54229_12380# VDD.t1405 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5431 a_30152_11614.t4 a_30152_10448.t19 a_32088_12380# VDD.t305 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5432 a_83709_n18620# a_71281_n10073.t278 a_83141_n18620# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5433 VDD.t1376 VDD.t1375 VDD.t1376 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5434 VDD.t1374 VDD.t1372 VDD.t1374 VDD.t1373 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5435 VDD.t250 a_31699_20742.t228 a_33249_48695.t190 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5436 VSS.t1114 VSS.t1113 VSS.t1114 VSS.t609 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5437 VDD.t388 a_30152_10448.t20 a_30682_10448# VDD.t326 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5438 VDD.t1371 VDD.t1369 VDD.t1371 VDD.t1370 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5439 a_52585_n2653# a_50751_n19729.t307 a_52063_n3550# VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5440 VSS.t1112 VSS.t1110 VSS.t1112 VSS.t1111 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5441 VDD.t1368 VDD.t1367 VDD.t1368 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5442 a_96849_10448# a_81205_n14095.t8 a_84017_n17715.t1 VDD.t499 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5443 VDD.t1366 VDD.t1364 VDD.t1366 VDD.t1365 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5444 a_108602_7563# a_100820_11614.t21 a_100992_4421.t0 VSS.t147 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5445 a_36530_7563# a_30152_11614.t19 a_36008_7563.t3 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5446 VSS.t1109 VSS.t1108 VSS.t1109 VSS.t307 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5447 VDD.t1363 VDD.t1362 VDD.t1363 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5448 a_85129_n28415# a_83325_n29313.t0 a_31831_n5342.t1 VSS.t286 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5449 a_54579_n2653# a_50751_n19729.t308 a_54019_n2653# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5450 a_32353_n5342# a_31953_n19727.t311 a_31831_n5342.t0 VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5451 a_31699_20742.t12 a_31699_20742.t11 VDD.t22 VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5452 VDD.t251 a_31699_20742.t229 a_33249_48695.t189 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5453 VSS.t1107 VSS.t1106 VSS.t1107 VSS.t650 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5454 a_33249_34067.t2 a_35502_24538.t58 a_52635_34067.t57 VSS.t184 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5455 VDD.t1361 VDD.t1360 VDD.t1361 VDD.t497 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5456 VSS.t1105 VSS.t1103 VSS.t1105 VSS.t1104 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5457 a_81735_n6960# a_71281_n10073.t279 a_81205_n7865# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5458 a_36530_n30339# a_30152_n36322.t21 a_36008_n30339.t1 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5459 a_31953_n19727.t17 a_31953_n19727.t16 VSS.t67 VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5460 VSS.t348 a_89163_10388.t20 a_89563_11614# VDD.t554 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5461 VDD.t1359 VDD.t1358 VDD.t1359 VDD.t405 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5462 VSS.t1102 VSS.t1101 VSS.t1102 VSS.t331 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5463 a_75602_n4019# a_71266_n4019.t0 VDD.t4772 VDD.t692 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X5464 VDD.t1357 VDD.t1356 VDD.t1357 VDD.t520 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5465 VSS.t1100 VSS.t1099 VSS.t1100 VSS.t641 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5466 VDD.t1355 VDD.t1353 VDD.t1355 VDD.t1354 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5467 VDD.t1352 VDD.t1351 VDD.t1352 VDD.t1015 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5468 a_98829_n6960# a_71281_n8397.t287 a_98299_n7865# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5469 a_33249_34067.t115 a_35502_25545.t88 VSS.t133 VSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5470 VDD.t1350 VDD.t1348 VDD.t1350 VDD.t1349 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5471 VSS.t1098 VSS.t1097 VSS.t1098 VSS.t638 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5472 VSS.t1096 VSS.t1095 VSS.t1096 VSS.t757 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5473 VDD.t1347 VDD.t1346 VDD.t1347 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5474 VDD.t430 a_71281_n8397.t6 a_71281_n8397.t7 VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5475 VSS.t1094 VSS.t1093 VSS.t1094 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5476 VDD.t1345 VDD.t1344 VDD.t1345 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5477 a_52635_34067.t37 a_35922_19591.t151 a_52635_48695.t20 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5478 VDD.t1343 VDD.t1342 VDD.t1343 VDD.t406 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5479 VDD.t1341 VDD.t1340 VDD.t1341 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5480 VSS.t1092 VSS.t1091 VSS.t1092 VSS.t647 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5481 a_47819_11614.t6 a_47991_5507.t1 a_49795_4481# VSS.t337 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5482 a_89531_n28415# a_83153_n36322.t20 VDD.t4783 VSS.t454 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5483 a_39179_n8930.t1 a_100820_n36322.t19 a_107198_n29181# VSS.t336 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5484 VDD.t1339 VDD.t1337 VDD.t1339 VDD.t1338 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5485 VDD.t252 a_31699_20742.t230 a_33249_48695.t188 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5486 VDD.t4823 a_52635_34067.t217 a_52635_49681.t101 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5487 VDD.t1336 VDD.t1335 VDD.t1336 VDD.t401 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5488 a_93131_n18620# a_71281_n10073.t280 a_92601_n19525# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5489 a_87433_n7865# a_71281_n10073.t281 a_86903_n7865# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5490 VDD.t1334 VDD.t1332 VDD.t1334 VDD.t1333 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5491 VDD.t1331 VDD.t1330 VDD.t1331 VDD.t1015 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5492 a_88271_n18620# a_71281_n10073.t282 a_87433_n18620# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5493 VDD.t1329 VDD.t1328 VDD.t1329 VDD.t498 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5494 VDD.t1327 VDD.t1326 VDD.t1327 VDD.t47 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5495 VDD.t1325 VDD.t1324 VDD.t1325 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5496 a_63683_n18700# a_50751_n19729.t309 a_63161_n19597# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5497 a_42442_n36322# a_36032_n35156.t12 a_36162_n36382.t5 VDD.t560 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5498 a_73302_n34390# a_71496_n36382.t16 VSS.t365 VDD.t2812 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5499 VSS.t1090 VSS.t1089 VSS.t1090 VSS.t376 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5500 VSS.t1088 VSS.t1087 VSS.t1088 VSS.t976 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5501 a_49795_6405# a_47991_5507.t2 a_48951_4481.t1 VSS.t338 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5502 VDD.t1323 VDD.t1321 VDD.t1323 VDD.t1322 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5503 VSS.t1086 VSS.t1085 VSS.t1086 VSS.t553 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5504 a_38097_n16007.t1 a_39179_n19595.t0 a_48391_n28415# VSS.t340 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5505 VDD.t4822 a_52635_34067.t218 a_52635_48695.t97 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5506 VDD.t1320 VDD.t1319 VDD.t1320 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5507 a_41100_19698# a_35502_24538.t59 a_40578_19075# VSS.t191 nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X5508 VDD.t1318 VDD.t1317 VDD.t1318 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5509 VSS.t1084 VSS.t1083 VSS.t1084 VSS.t633 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5510 a_44885_n4445# a_31953_n19727.t312 a_44363_n4445# VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5511 a_100235_n13190# a_71281_n8397.t288 a_99667_n13190# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5512 a_95105_n9675# a_71281_n10073.t283 a_94537_n9675# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5513 VSS.t1082 VSS.t1081 VSS.t1082 VSS.t413 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5514 VSS.t1080 VSS.t1079 VSS.t1080 VSS.t305 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5515 VSS.t1078 VSS.t1076 VSS.t1078 VSS.t1077 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X5516 a_57417_n8035# a_50751_n19729.t310 a_56895_n8932# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5517 a_31953_n19727.t15 a_31953_n19727.t14 VSS.t66 VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5518 VSS.t1075 VSS.t1074 VSS.t1075 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5519 VDD.t1316 VDD.t1315 VDD.t1316 VDD.t321 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5520 VDD.t1314 VDD.t1313 VDD.t1314 VDD.t47 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5521 a_37934_n29181# a_30152_n36322.t22 a_30324_n30399.t1 VSS.t282 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5522 a_47753_n13316# a_31953_n19727.t313 a_47231_n14213# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5523 VDD.t1312 VDD.t1311 VDD.t1312 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5524 VDD.t1310 VDD.t1309 VDD.t1310 VDD.t965 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5525 VSS.t1073 VSS.t1072 VSS.t1073 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5526 VDD.t1308 VDD.t1307 VDD.t1308 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5527 a_107339_n3340# a_71281_n8397.t289 a_106501_n2435# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5528 VSS.t1071 VSS.t1070 VSS.t1071 VSS.t795 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5529 VSS.t1069 VSS.t1068 VSS.t1069 VSS.t27 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5530 VDD.t1306 VDD.t1305 VDD.t1306 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5531 a_33249_48695.t187 a_31699_20742.t231 VDD.t253 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5532 VDD.t1304 VDD.t1303 VDD.t1304 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5533 a_48391_4481# a_47991_4421.t2 a_47819_10448.t9 VSS.t339 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5534 VDD.t1302 VDD.t1301 VDD.t1302 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5535 a_42047_n4445# a_31953_n19727.t314 a_41487_n3548# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5536 VDD.t1300 VDD.t1298 VDD.t1300 VDD.t1299 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5537 VSS.t1067 VSS.t1066 VSS.t1067 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5538 VDD.t1297 VDD.t1296 VDD.t1297 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5539 VSS.t1065 VSS.t1063 VSS.t1065 VSS.t1064 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5540 a_98829_n13190# a_71281_n8397.t290 a_98299_n16810# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5541 a_54019_n16906# a_50751_n19729.t311 a_53497_n16906# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5542 a_33249_48695.t186 a_31699_20742.t232 VDD.t254 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5543 a_93131_n6960# a_71281_n10073.t284 a_92601_n7865# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5544 VSS.t1062 VSS.t1061 VSS.t1062 VSS.t612 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5545 VDD.t4821 a_52635_34067.t219 a_52635_48695.t96 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5546 VDD.t1295 VDD.t1294 VDD.t1295 VDD.t434 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5547 VDD.t1293 VDD.t1292 VDD.t1293 VDD.t965 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5548 VDD.t294 a_100820_10448.t18 a_101350_13546# VDD.t293 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5549 VSS.t1060 VSS.t1059 VSS.t1060 VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5550 a_31953_n19727.t13 a_31953_n19727.t12 VSS.t64 VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5551 VDD.t255 a_31699_20742.t233 a_33249_48695.t185 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5552 a_67111_n15112# a_50751_n19729.t312 a_66551_n15112# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5553 a_36162_10388.t4 a_36032_11614.t10 a_43848_10448# VDD.t287 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5554 VDD.t1291 VDD.t1289 VDD.t1291 VDD.t1290 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5555 VDD.t1288 VDD.t1287 VDD.t1288 VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5556 a_105365_n13190# a_71281_n8397.t291 a_104527_n13190# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5557 VSS.t1058 VSS.t1057 VSS.t1058 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5558 VDD.t1286 VDD.t1285 VDD.t1286 VDD.t423 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5559 a_65117_n19597# a_50751_n19729.t313 VSS.t278 VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5560 a_35502_25545.t18 a_31699_20742.t234 VDD.t256 VDD.t20 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5561 VDD.t1284 VDD.t1283 VDD.t1284 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5562 VSS.t1056 VSS.t1055 VSS.t1056 VSS.t501 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5563 VSS.t1054 VSS.t1053 VSS.t1054 VSS.t498 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5564 VDD.t1282 VDD.t1281 VDD.t1282 VDD.t1142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5565 VSS.t1052 VSS.t1051 VSS.t1052 VSS.t550 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5566 VDD.t1280 VDD.t1279 VDD.t1280 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5567 VDD.t1278 VDD.t1277 VDD.t1278 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5568 a_59411_n19597# a_50751_n19729.t314 a_58851_n19597# VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5569 VDD.t420 a_100820_10448.t19 a_101350_11614# VDD.t293 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5570 VDD.t1276 VDD.t1275 VDD.t1276 VDD.t405 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5571 VSS.t1050 VSS.t1049 VSS.t1050 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5572 a_33249_35053.t92 a_35502_24538.t60 OUT.t4 VSS.t192 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5573 a_33249_48695.t83 a_33379_34917.t73 a_33249_35053.t69 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5574 a_33249_48695.t143 a_33379_34007.t79 a_33249_34067.t31 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5575 VSS.t1048 VSS.t1047 VSS.t1048 VSS.t498 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5576 VSS.t1046 VSS.t1045 VSS.t1046 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5577 VSS.t1044 VSS.t1043 VSS.t1044 VSS.t490 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5578 VSS.t1042 VSS.t1041 VSS.t1042 VSS.t937 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5579 VDD.t1274 VDD.t1273 VDD.t1274 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5580 VDD.t1272 VDD.t1271 VDD.t1272 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5581 VSS.t1040 VSS.t1039 VSS.t1040 VSS.t834 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5582 a_35502_24538.t3 a_31699_20742.t235 VDD.t257 VDD.t32 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5583 VDD.t1270 VDD.t1269 VDD.t1270 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5584 a_75585_n8397# I1N.t14 VSS.t437 VSS.t430 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X5585 a_45445_n12419# a_31953_n19727.t315 a_44885_n12419# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5586 a_52635_49681.t66 a_35922_19591.t152 OUT.t41 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5587 VDD.t1268 VDD.t1267 VDD.t1268 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5588 VSS.t1038 VSS.t1036 VSS.t1038 VSS.t1037 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5589 VSS.t1035 VSS.t1033 VSS.t1035 VSS.t1034 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5590 VSS.t362 a_94892_n29181.t20 a_95414_n29181# VSS.t357 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5591 a_43817_n27257# a_41891_n29181.t21 VSS.t374 VSS.t158 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5592 a_112199_n3340# a_71281_n8397.t292 a_111631_n3340# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5593 a_90935_6405# a_83153_11614.t20 a_51711_n12421.t0 VSS.t395 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5594 a_52635_48695.t95 a_52635_34067.t220 VDD.t4820 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5595 VDD.t1266 VDD.t1264 VDD.t1266 VDD.t1265 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5596 a_39179_n1754# a_31953_n19727.t316 a_38619_n1754# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5597 VDD.t1263 VDD.t1261 VDD.t1263 VDD.t1262 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5598 a_49795_n27257# a_39179_n19595.t0 a_38097_n16007.t2 VSS.t338 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5599 VSS.t1032 VSS.t1031 VSS.t1032 VSS.t576 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5600 a_32353_n13316# a_31953_n19727.t317 a_31831_n13316# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5601 VSS.t1030 VSS.t1029 VSS.t1030 VSS.t99 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5602 VDD.t1260 VDD.t1259 VDD.t1260 VDD.t930 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5603 a_71281_n8397.t5 a_71281_n8397.t4 VDD.t428 VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5604 VDD.t1258 VDD.t1257 VDD.t1258 VDD.t70 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5605 a_54019_n2653# a_50751_n19729.t315 a_53497_n3550# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5606 VSS.t1028 VSS.t1027 VSS.t1028 VSS.t184 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5607 a_104527_n6960# a_71281_n8397.t293 a_103997_n7865# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5608 VDD.t1256 VDD.t1255 VDD.t1256 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5609 a_89033_13546.t1 a_106830_10388.t19 a_108636_13546# VDD.t521 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5610 VSS.t1026 VSS.t1024 VSS.t1026 VSS.t1025 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5611 a_112199_n15000# a_71281_n8397.t294 a_111631_n15000# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5612 a_82573_n8770# a_71281_n10073.t285 a_81735_n8770# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5613 a_111631_n7865# a_71281_n8397.t295 a_111063_n7865# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5614 VSS.t1023 VSS.t1022 VSS.t1023 VSS.t63 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5615 VSS.t1021 VSS.t1020 VSS.t1021 VSS.t525 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5616 a_52635_34067.t40 a_35922_19591.t153 a_52635_48695.t19 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5617 VSS.t1019 VSS.t1018 VSS.t1019 VSS.t553 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5618 a_66058_6405# a_65658_4421.t0 a_65486_10448.t10 VSS.t376 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5619 a_71281_n10073.t13 a_71281_n10073.t12 VDD.t358 VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5620 VSS.t1017 VSS.t1016 VSS.t1017 VSS.t399 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5621 VDD.t1254 VDD.t1253 VDD.t1254 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5622 a_33249_48695.t84 a_33379_34917.t74 a_33249_35053.t70 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5623 VDD.t1252 VDD.t1250 VDD.t1252 VDD.t1251 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5624 a_83683_n34390# a_83153_n35156.t21 a_83153_n36322.t5 VDD.t2729 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5625 a_77225_n29181.t6 a_77225_n29181.t5 a_79151_n30339# VSS.t380 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5626 VDD.t1249 VDD.t1248 VDD.t1249 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5627 VSS.t1015 VSS.t1014 VSS.t1015 VSS.t329 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5628 VDD.t1247 VDD.t1246 VDD.t1247 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5629 a_99667_n8770# a_71281_n8397.t296 a_98829_n8770# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5630 a_89009_n27257.t0 a_83153_n36322.t21 a_90935_n30339# VSS.t455 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5631 VSS.t1013 VSS.t1012 VSS.t1013 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5632 a_38619_n8930# a_31953_n19727.t318 a_38097_n8930# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5633 VDD.t1245 VDD.t1244 VDD.t1245 VDD.t78 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5634 VDD.t1243 VDD.t1242 VDD.t1243 VDD.t404 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5635 VDD.t1241 VDD.t1240 VDD.t1241 VDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5636 VDD.t1239 VDD.t1238 VDD.t1239 VDD.t905 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5637 VSS.t1011 VSS.t1010 VSS.t1011 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5638 VDD.t1237 VDD.t1236 VDD.t1237 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5639 VSS.t1009 VSS.t1008 VSS.t1009 VSS.t459 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5640 a_33249_48695.t144 a_33379_34007.t80 a_33249_34067.t30 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5641 VSS.t1007 VSS.t1006 VSS.t1007 VSS.t398 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5642 VSS.t1005 VSS.t1004 VSS.t1005 VSS.t668 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5643 VDD.t1235 VDD.t1234 VDD.t1235 VDD.t893 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5644 a_86903_n14095.t0 a_106830_10388.t20 a_108636_11614# VDD.t521 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5645 VDD.t1233 VDD.t1232 VDD.t1233 VDD.t619 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5646 OUT.t40 a_35922_19591.t154 a_52635_49681.t67 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5647 VDD.t4819 a_52635_34067.t221 a_52635_48695.t94 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5648 a_58851_n12421# a_50751_n19729.t316 a_57977_n16009.t0 VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5649 VSS.t1003 VSS.t1002 VSS.t1003 VSS.t537 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5650 a_33249_34067.t114 a_35502_25545.t89 VSS.t132 VSS.t3 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5651 VDD.t1231 VDD.t1230 VDD.t1231 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5652 a_33249_48695.t184 a_31699_20742.t236 VDD.t258 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5653 VSS.t1001 VSS.t1000 VSS.t1001 VSS.t266 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5654 VSS.t999 VSS.t997 VSS.t999 VSS.t998 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5655 a_100803_n9675# a_71281_n8397.t297 a_100235_n9675# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5656 VSS.t996 VSS.t995 VSS.t996 VSS.t213 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5657 a_60845_n17803# a_50751_n19729.t317 a_60285_n17803# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5658 VDD.t1229 VDD.t1228 VDD.t1229 VDD.t905 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5659 VSS.t994 VSS.t993 VSS.t994 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5660 VDD.t1227 VDD.t1226 VDD.t1227 VDD.t893 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5661 a_57417_n14215# a_50751_n19729.t318 a_56895_n15112# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5662 VDD.t1225 VDD.t1224 VDD.t1225 VDD.t519 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5663 a_47819_11614.t2 a_47819_10448.t19 a_49755_12380# VDD.t496 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5664 VDD.t1223 VDD.t1222 VDD.t1223 VDD.t875 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5665 VDD.t1221 VDD.t1220 VDD.t1221 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5666 VDD.t1219 VDD.t1217 VDD.t1219 VDD.t1218 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5667 VDD.t1216 VDD.t1215 VDD.t1216 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5668 VSS.t992 VSS.t991 VSS.t992 VSS.t217 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5669 VSS.t990 VSS.t989 VSS.t990 VSS.t588 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5670 a_32088_10448# a_30152_10448.t21 VDD.t389 VDD.t303 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5671 VSS.t988 VSS.t987 VSS.t988 VSS.t102 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5672 a_37934_4481# a_30152_11614.t20 a_30324_4421.t0 VSS.t282 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5673 a_93131_n17715# a_71281_n10073.t286 a_92601_n21335# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5674 a_33249_48695.t183 a_31699_20742.t237 VDD.t259 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5675 VDD.t1214 VDD.t1213 VDD.t1214 VDD.t120 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5676 VDD.t369 a_71281_n10073.t10 a_71281_n10073.t11 VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5677 VSS.t62 a_31953_n19727.t10 a_31953_n19727.t11 VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5678 a_71281_n10073.t9 a_71281_n10073.t8 VDD.t345 VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5679 VDD.t1212 VDD.t1211 VDD.t1212 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5680 a_57417_n3550# a_50751_n19729.t319 a_56895_n4447# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5681 VSS.t986 VSS.t985 VSS.t986 VSS.t335 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5682 VDD.t1210 VDD.t1208 VDD.t1210 VDD.t1209 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5683 VDD.t1207 VDD.t1205 VDD.t1207 VDD.t1206 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5684 VDD.t1204 VDD.t1203 VDD.t1204 VDD.t302 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5685 VSS.t984 VSS.t983 VSS.t984 VSS.t528 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5686 VDD.t1202 VDD.t1201 VDD.t1202 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5687 a_112199_n20430# a_71281_n8397.t298 a_111631_n20430# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5688 VSS.t982 VSS.t981 VSS.t982 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5689 a_93969_n18620# a_71281_n10073.t287 a_93131_n18620# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5690 VDD.t1200 VDD.t1199 VDD.t1200 VDD.t852 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5691 VDD.t4818 a_52635_34067.t222 a_52635_49681.t100 VDD.t401 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5692 VSS.t980 VSS.t978 VSS.t980 VSS.t979 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5693 a_66551_n2653# a_50751_n19729.t320 a_66029_n3550# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5694 a_41891_4481.t10 a_41891_4481.t9 a_43817_5639# VSS.t168 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5695 VDD.t1198 VDD.t1197 VDD.t1198 VDD.t875 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5696 a_54579_n17803# a_50751_n19729.t321 a_54019_n17803# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5697 a_66058_n27257# a_65658_n29313.t2 a_65486_n35156.t11 VSS.t376 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5698 VSS.t977 VSS.t975 VSS.t977 VSS.t976 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5699 a_83709_n21335# a_71281_n10073.t288 a_83141_n21335# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5700 a_64243_n18700# a_50751_n19729.t322 a_63683_n17803# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5701 VDD.t1196 VDD.t1194 VDD.t1196 VDD.t1195 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5702 a_33787_n8033# a_31953_n19727.t319 a_33265_n8033# VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5703 VDD.t1193 VDD.t1192 VDD.t1193 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5704 a_89407_n19525# a_71281_n10073.t289 a_88839_n19525# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5705 a_46879_n3548# a_31953_n19727.t320 a_47753_n5342# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5706 a_50751_n19729.t21 a_50751_n19729.t20 VSS.t228 VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5707 VSS.t974 VSS.t973 VSS.t974 VSS.t618 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5708 VSS.t3634 a_59558_n29181.t20 a_60080_n28415# VSS.t401 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5709 VDD.t1191 VDD.t1190 VDD.t1191 VDD.t852 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5710 VSS.t972 VSS.t971 VSS.t972 VSS.t56 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5711 VDD.t1189 VDD.t1187 VDD.t1189 VDD.t1188 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X5712 a_100803_n19525# a_71281_n8397.t299 a_100235_n19525# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5713 a_45445_n8033# a_31953_n19727.t321 a_44885_n8033# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5714 VDD.t1186 VDD.t1185 VDD.t1186 VDD.t25 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5715 VSS.t970 VSS.t969 VSS.t970 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5716 VDD.t1184 VDD.t1182 VDD.t1184 VDD.t1183 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5717 a_33249_48695.t145 a_33379_34007.t81 a_33249_34067.t29 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5718 a_31699_20742.t10 a_31699_20742.t9 VDD.t21 VDD.t20 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5719 a_64243_n8035# a_50751_n19729.t323 a_63683_n8035# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5720 a_75602_n4978# a_71266_n4019.t0 VDD.t4771 VDD.t692 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X5721 VDD.t260 a_31699_20742.t238 a_33249_48695.t182 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5722 VDD.t1181 VDD.t1179 VDD.t1181 VDD.t1180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5723 a_52635_48695.t18 a_35922_19591.t155 a_52635_34067.t45 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5724 VSS.t61 a_31953_n19727.t8 a_31953_n19727.t9 VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5725 a_100820_10448.t2 a_100992_4421.t0 a_102796_5639# VSS.t171 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5726 a_31284_4481.t2 a_30324_5507.t1 a_30724_5639# VSS.t151 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5727 a_33249_48695.t181 a_31699_20742.t239 VDD.t261 VDD.t115 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5728 a_66016_n36322# a_65486_n35156.t22 a_65486_n36322.t3 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5729 VDD.t1178 VDD.t1176 VDD.t1178 VDD.t1177 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5730 a_40613_n7136# a_31953_n19727.t322 a_40053_n7136# VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5731 VSS.t968 VSS.t967 VSS.t968 VSS.t288 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5732 a_71281_n10073.t7 a_71281_n10073.t6 VDD.t365 VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5733 a_57977_n18700# a_50751_n19729.t324 a_57417_n17803# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5734 VDD.t1175 VDD.t1174 VDD.t1175 VDD.t553 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5735 VSS.t966 VSS.t965 VSS.t966 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5736 VDD.t1173 VDD.t1172 VDD.t1173 VDD.t833 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5737 a_65486_11614.t0 a_65486_10448.t19 a_67422_12380# VDD.t1378 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5738 VDD.t1171 VDD.t1170 VDD.t1171 VDD.t801 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5739 a_83141_n15000# a_71281_n10073.t290 a_82573_n15000# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5740 VSS.t964 VSS.t963 VSS.t964 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5741 VSS.t962 VSS.t961 VSS.t962 VSS.t5 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X5742 VSS.t960 VSS.t959 VSS.t960 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5743 VSS.t958 VSS.t957 VSS.t958 VSS.t856 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5744 VSS.t956 VSS.t955 VSS.t956 VSS.t464 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5745 a_54197_6405# a_47819_11614.t19 VDD.t505 VSS.t306 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5746 a_59558_4481.t8 a_47991_4421.t1 a_61515_13546# VDD.t1512 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5747 a_93131_n21335# a_71281_n10073.t291 a_92601_n21335# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5748 VDD.t1169 VDD.t1168 VDD.t1169 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5749 VSS.t954 VSS.t953 VSS.t954 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5750 a_43817_5639# a_41891_4481.t19 VSS.t174 VSS.t158 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5751 a_88271_n21335# a_71281_n10073.t292 a_87433_n21335# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5752 VDD.t1167 VDD.t1166 VDD.t1167 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5753 a_52635_48695.t17 a_35922_19591.t156 a_52635_34067.t40 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5754 VSS.t952 VSS.t951 VSS.t952 VSS.t99 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5755 VSS.t59 a_31953_n19727.t6 a_31953_n19727.t7 VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5756 VDD.t1165 VDD.t1163 VDD.t1165 VDD.t1164 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5757 VDD.t1162 VDD.t1161 VDD.t1162 VDD.t833 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5758 VDD.t1160 VDD.t1159 VDD.t1160 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5759 VDD.t1158 VDD.t1157 VDD.t1158 VDD.t801 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5760 a_81735_n17715# a_71281_n10073.t293 a_81205_n16810# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5761 VSS.t950 VSS.t949 VSS.t950 VSS.t424 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5762 VDD.t1156 VDD.t1154 VDD.t1156 VDD.t1155 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5763 VDD.t1153 VDD.t1152 VDD.t1153 VDD.t976 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5764 VDD.t1151 VDD.t1150 VDD.t1151 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5765 a_59558_4481.t9 a_47991_4421.t1 a_61515_11614# VDD.t1512 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5766 VSS.t948 VSS.t946 VSS.t948 VSS.t947 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5767 VSS.t945 VSS.t943 VSS.t945 VSS.t944 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5768 VDD.t1149 VDD.t1148 VDD.t1149 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5769 VSS.t942 VSS.t941 VSS.t942 VSS.t495 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5770 a_52635_48695.t16 a_35922_19591.t157 a_52635_34067.t24 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5771 VDD.t1147 VDD.t1146 VDD.t1147 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5772 VSS.t940 VSS.t939 VSS.t940 VSS.t681 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5773 a_81735_n15000# a_71281_n10073.t294 a_81205_n15905# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5774 a_93969_n6960# a_71281_n10073.t295 a_93131_n6960# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5775 a_33379_34917.t2 a_36162_10388.t21 a_37968_13546# VDD.t1494 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5776 a_112199_n2435# a_71281_n8397.t300 a_111631_n2435# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5777 a_42047_n15110# a_31953_n19727.t323 a_41487_n15110# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5778 VSS.t938 VSS.t936 VSS.t938 VSS.t937 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5779 VSS.t935 VSS.t934 VSS.t935 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5780 a_41487_n6239# a_31953_n19727.t324 a_40965_n6239# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5781 OUT.t39 a_35922_19591.t158 a_52635_49681.t68 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5782 a_52635_34067.t38 a_35922_19591.t159 a_52635_48695.t15 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5783 a_101392_5639# a_57977_n12421.t0 a_100820_11614.t7 VSS.t163 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5784 VDD.t1145 VDD.t1144 VDD.t1145 VDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5785 a_94537_n1530# a_71281_n10073.t296 a_93969_n1530# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5786 a_33249_48695.t146 a_33379_34007.t82 a_33249_34067.t28 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5787 VSS.t933 VSS.t932 VSS.t933 VSS.t392 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5788 a_112199_n15905# a_71281_n8397.t301 a_111631_n15905# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5789 VSS.t227 a_50751_n19729.t18 a_50751_n19729.t19 VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5790 VSS.t931 VSS.t930 VSS.t931 VSS.t478 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5791 a_30724_5639# a_30324_5507.t1 a_30152_11614.t2 VSS.t150 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5792 a_82573_n7865# a_71281_n10073.t297 a_81735_n7865# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5793 VSS.t929 VSS.t928 VSS.t929 VSS.t671 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5794 VSS.t927 VSS.t926 VSS.t927 VSS.t687 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5795 VDD.t1143 VDD.t1141 VDD.t1143 VDD.t1142 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5796 a_71342_4481.t3 a_71496_10388.t23 a_71896_10448# VDD.t353 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5797 VSS.t925 VSS.t924 VSS.t925 VSS.t495 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5798 VDD.t1140 VDD.t1139 VDD.t1140 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5799 VDD.t1138 VDD.t1137 VDD.t1138 VDD.t789 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5800 VDD.t1136 VDD.t1135 VDD.t1136 VDD.t497 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5801 a_33249_48695.t85 a_33379_34917.t75 a_33249_35053.t71 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5802 VSS.t923 VSS.t922 VSS.t923 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5803 VSS.t921 VSS.t920 VSS.t921 VSS.t195 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5804 a_36032_11614.t1 a_36162_10388.t22 a_37968_11614# VDD.t1494 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5805 VDD.t1134 VDD.t1133 VDD.t1134 VDD.t47 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5806 VSS.t919 VSS.t918 VSS.t919 VSS.t568 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5807 VSS.t917 VSS.t916 VSS.t917 VSS.t294 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5808 VDD.t1132 VDD.t1131 VDD.t1132 VDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5809 a_30324_n30399.t0 a_31953_n19727.t325 a_32353_n19595# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5810 a_99667_n7865# a_71281_n8397.t302 a_98829_n7865# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5811 a_42047_n2651# a_31953_n19727.t326 a_41487_n2651# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5812 a_33249_34067.t113 a_35502_25545.t90 VSS.t131 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5813 VSS.t407 a_59558_4481.t21 a_60080_4481# VSS.t401 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5814 a_83141_n20430# a_71281_n10073.t298 a_82573_n20430# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5815 VSS.t915 VSS.t914 VSS.t915 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5816 a_33249_48695.t86 a_33379_34917.t76 a_33249_35053.t72 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5817 a_61484_n27257# a_59558_n29181.t21 VSS.t3635 VSS.t399 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5818 a_32913_n6239# a_31953_n19727.t327 a_32353_n4445# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5819 a_83153_11614.t1 a_51711_n12421.t0 a_85129_4481# VSS.t308 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5820 a_33249_48695.t87 a_33379_34917.t77 a_33249_35053.t73 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5821 VSS.t913 VSS.t912 VSS.t913 VSS.t318 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5822 VSS.t911 VSS.t910 VSS.t911 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5823 VSS.t909 VSS.t907 VSS.t909 VSS.t908 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5824 a_100820_n36322.t7 a_39179_n8930.t1 a_102796_n27257# VSS.t329 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5825 VSS.t906 VSS.t904 VSS.t906 VSS.t905 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5826 VDD.t1130 VDD.t1129 VDD.t1130 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5827 VSS.t438 I1N.t15 a_72603_n9297# VSS.t433 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X5828 a_83709_n3340# a_71281_n10073.t299 a_83141_n3340# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5829 VDD.t4817 a_52635_34067.t223 a_52635_49681.t99 VDD.t404 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5830 VDD.t4816 a_52635_34067.t224 a_52635_49681.t98 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5831 a_73302_n36322# a_71496_n36382.t17 a_71342_n27257.t1 VDD.t2812 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5832 VDD.t1128 VDD.t1126 VDD.t1128 VDD.t1127 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5833 VDD.t1125 VDD.t1124 VDD.t1125 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5834 a_71864_n29181# a_65486_n36322.t23 VDD.t292 VSS.t156 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5835 VDD.t1123 VDD.t1122 VDD.t1123 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5836 a_52635_34067.t56 a_35502_24538.t61 a_33249_34067.t1 VSS.t193 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5837 VDD.t1121 VDD.t1120 VDD.t1121 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5838 a_81735_n20430# a_71281_n10073.t300 VDD.t385 VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5839 VDD.t1119 VDD.t1118 VDD.t1119 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5840 a_88839_n9675# a_71281_n10073.t301 a_88271_n9675# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5841 a_31284_n30339.t2 a_30324_n29313.t0 a_30724_n29181# VSS.t151 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5842 a_87433_n18620# a_71281_n10073.t302 a_86903_n19525# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5843 VDD.t1117 VDD.t1116 VDD.t1117 VDD.t925 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5844 VSS.t903 VSS.t902 VSS.t903 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5845 a_100820_n36322.t2 a_100820_n35156.t20 a_102756_n35156# VDD.t532 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5846 VDD.t1115 VDD.t1114 VDD.t1115 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5847 VDD.t1113 VDD.t1111 VDD.t1113 VDD.t1112 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5848 a_89407_n4245# a_71281_n10073.t303 a_88839_n4245# VDD.t341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5849 a_39179_n16904# a_31953_n19727.t328 a_38619_n15110# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5850 a_71496_10388.t7 a_71366_11614.t10 a_79182_10448# VDD.t1841 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5851 VDD.t1110 VDD.t1109 VDD.t1110 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5852 VSS.t901 VSS.t900 VSS.t901 VSS.t103 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5853 a_55601_n30339# a_47819_n36322.t22 a_47991_n29313.t0 VSS.t305 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5854 VSS.t899 VSS.t898 VSS.t899 VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5855 a_33249_48695.t88 a_33379_34917.t78 a_33249_35053.t74 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5856 VDD.t1108 VDD.t1107 VDD.t1108 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5857 a_33787_n3548# a_31953_n19727.t329 a_33265_n3548# VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5858 VSS.t897 VSS.t895 VSS.t897 VSS.t896 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5859 VSS.t894 VSS.t893 VSS.t894 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5860 a_71281_n10073.t5 a_71281_n10073.t4 VDD.t492 VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5861 a_33787_n12419# a_31953_n19727.t330 VSS.t120 VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5862 a_33249_48695.t180 a_31699_20742.t240 VDD.t262 VDD.t120 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5863 VSS.t892 VSS.t890 VSS.t892 VSS.t891 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5864 a_45445_n3548# a_31953_n19727.t331 a_44885_n3548# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5865 a_107198_n27257# a_100820_n36322.t20 a_106676_n27257.t0 VSS.t335 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5866 a_51711_n12421.t0 a_83153_11614.t21 a_89531_5639# VSS.t393 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5867 VDD.t1106 VDD.t1105 VDD.t1106 VDD.t14 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5868 a_48349_n34390# a_47819_n35156.t20 a_47819_n36322.t2 VDD.t2559 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5869 a_100820_n36322.t3 a_100820_n35156.t21 a_102756_n33224# VDD.t532 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5870 a_105933_n13190# a_71281_n8397.t303 a_105365_n13190# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5871 a_46879_n17801# a_31953_n19727.t332 a_46319_n17801# VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5872 VSS.t889 VSS.t888 VSS.t889 VSS.t45 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X5873 a_33249_48695.t179 a_31699_20742.t241 VDD.t263 VDD.t122 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5874 VDD.t1104 VDD.t1103 VDD.t1104 VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5875 VSS.t887 VSS.t886 VSS.t887 VSS.t25 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5876 VDD.t1102 VDD.t1101 VDD.t1102 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5877 VDD.t533 a_100820_n35156.t22 a_101350_n35156# VDD.t529 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5878 a_64243_n3550# a_50751_n19729.t325 a_63683_n3550# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5879 VDD.t1100 VDD.t1098 VDD.t1100 VDD.t1099 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5880 VDD.t1097 VDD.t1096 VDD.t1097 VDD.t910 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5881 a_51711_n18700# a_50751_n19729.t326 a_51151_n18700# VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5882 VDD.t1095 VDD.t1094 VDD.t1095 VDD.t898 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5883 VSS.t130 a_35502_25545.t91 a_35922_19591.t2 VSS.t129 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X5884 a_87433_n1530# a_71281_n10073.t304 a_86903_n5150# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5885 a_31699_20742.t8 a_31699_20742.t7 VDD.t19 VDD.t18 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5886 VDD.t1093 VDD.t1092 VDD.t1093 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5887 a_35781_n4445# a_31953_n19727.t333 a_35221_n4445# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5888 VSS.t885 VSS.t883 VSS.t885 VSS.t884 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5889 VDD.t1091 VDD.t1090 VDD.t1091 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5890 VDD.t1089 VDD.t1088 VDD.t1089 VDD.t320 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5891 VDD.t1087 VDD.t1085 VDD.t1087 VDD.t1086 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5892 a_53145_n14215# a_50751_n19729.t327 a_52585_n14215# VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5893 VSS.t882 VSS.t881 VSS.t882 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5894 VSS.t880 VSS.t879 VSS.t880 VSS.t286 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5895 a_65486_n35156.t10 a_65658_n29313.t0 a_67462_n28415# VSS.t378 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5896 a_71281_n8397.t3 a_71281_n8397.t2 VDD.t426 VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5897 VSS.t878 VSS.t876 VSS.t878 VSS.t877 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5898 VSS.t875 VSS.t874 VSS.t875 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5899 VDD.t1084 VDD.t1083 VDD.t1084 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5900 VDD.t534 a_100820_n35156.t23 a_101350_n33224# VDD.t529 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5901 a_104527_n13190# a_71281_n8397.t304 a_103997_n16810# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5902 VSS.t873 VSS.t872 VSS.t873 VSS.t18 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5903 a_95105_n3340# a_71281_n10073.t305 a_94537_n3340# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5904 VDD.t1082 VDD.t1080 VDD.t1082 VDD.t1081 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5905 a_31699_17542# I1U.t6 VSS.t351 VSS.t349 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X5906 VSS.t871 VSS.t870 VSS.t871 VSS.t153 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5907 a_83141_n15905# a_71281_n10073.t306 a_82573_n15905# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5908 VDD.t264 a_31699_20742.t242 a_33249_48695.t178 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5909 VDD.t1079 VDD.t1078 VDD.t1079 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5910 a_52635_49681.t69 a_35922_19591.t160 OUT.t38 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5911 a_52635_34067.t46 a_35922_19591.t161 a_52635_48695.t14 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5912 a_83141_n9675# a_71281_n10073.t307 a_82573_n9675# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5913 VSS.t869 VSS.t867 VSS.t869 VSS.t868 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5914 VSS.t866 VSS.t865 VSS.t866 VSS.t757 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5915 VDD.t1077 VDD.t1076 VDD.t1077 VDD.t920 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X5916 VDD.t1075 VDD.t1074 VDD.t1075 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5917 a_33249_48695.t89 a_33379_34917.t79 a_33249_35053.t75 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5918 VDD.t1073 VDD.t1072 VDD.t1073 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5919 VDD.t1071 VDD.t1070 VDD.t1071 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5920 a_36562_n35156# a_36162_n36382.t22 a_36032_n35156.t4 VDD.t680 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5921 VSS.t864 VSS.t863 VSS.t864 VSS.t558 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5922 VSS.t344 a_89163_n36382.t22 a_89563_n34390# VDD.t547 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5923 a_41487_n16007# a_31953_n19727.t334 a_40613_n17801# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5924 VDD.t265 a_31699_20742.t243 a_33249_48695.t177 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5925 VSS.t862 VSS.t861 VSS.t862 VSS.t454 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5926 VDD.t1069 VDD.t1068 VDD.t1069 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5927 VSS.t860 VSS.t858 VSS.t860 VSS.t859 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5928 VSS.t128 a_35502_25545.t92 a_33249_34067.t112 VSS.t33 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5929 a_100235_n9675# a_71281_n8397.t305 a_99667_n9675# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5930 VDD.t1067 VDD.t1066 VDD.t1067 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5931 VDD.t515 a_47819_10448.t20 a_48349_13546# VDD.t510 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5932 a_33249_48695.t147 a_33379_34007.t83 a_33249_34067.t27 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5933 VSS.t857 VSS.t855 VSS.t857 VSS.t856 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5934 a_89531_5639# a_83153_11614.t22 VDD.t4765 VSS.t394 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5935 VDD.t1065 VDD.t1064 VDD.t1065 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5936 a_93969_n21335# a_71281_n10073.t308 a_93131_n21335# VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5937 a_47753_n8033# a_31953_n19727.t335 a_47231_n8033# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5938 a_57417_n2653# a_50751_n19729.t328 a_56895_n2653# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5939 VSS.t854 VSS.t852 VSS.t854 VSS.t853 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5940 VDD.t1063 VDD.t1062 VDD.t1063 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5941 a_81735_n15905# a_71281_n10073.t309 a_81205_n15905# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5942 VSS.t851 VSS.t850 VSS.t851 VSS.t596 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5943 a_81735_n6055# a_71281_n10073.t310 a_81205_n9675# VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5944 VSS.t849 VSS.t848 VSS.t849 VSS.t102 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5945 a_99667_n19525# a_71281_n8397.t306 a_98829_n19525# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5946 VDD.t1061 VDD.t1060 VDD.t1061 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5947 VDD.t1059 VDD.t1058 VDD.t1059 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5948 VDD.t1057 VDD.t1056 VDD.t1057 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5949 VSS.t847 VSS.t846 VSS.t847 VSS.t340 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5950 a_36562_n33224# a_36162_n36382.t23 a_33379_34007.t3 VDD.t680 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5951 a_60845_n8932# a_50751_n19729.t329 a_60285_n8932# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5952 a_33249_48695.t90 a_33379_34917.t80 a_33249_35053.t76 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5953 a_83683_n36322# a_83153_n35156.t22 a_83153_n36322.t6 VDD.t2729 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5954 VDD.t1055 VDD.t1054 VDD.t1055 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5955 VDD.t266 a_31699_20742.t244 a_35502_25545.t19 VDD.t16 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5956 a_52635_34067.t40 a_35922_19591.t162 a_52635_48695.t13 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5957 VSS.t845 VSS.t844 VSS.t845 VSS.t490 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5958 VSS.t843 VSS.t841 VSS.t843 VSS.t842 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X5959 VDD.t1053 VDD.t1051 VDD.t1053 VDD.t1052 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5960 VDD.t1050 VDD.t1048 VDD.t1050 VDD.t1049 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5961 a_50751_n19729.t17 a_50751_n19729.t16 VSS.t226 VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5962 a_111063_n19525# a_71281_n8397.t307 a_110225_n19525# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5963 a_98829_n6055# a_71281_n8397.t308 a_98299_n9675# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5964 VSS.t840 VSS.t839 VSS.t840 VSS.t65 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5965 VDD.t1047 VDD.t1046 VDD.t1047 VDD.t828 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5966 a_52635_49681.t70 a_35922_19591.t163 OUT.t37 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5967 VDD.t516 a_47819_10448.t21 a_48349_11614# VDD.t510 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5968 VDD.t1045 VDD.t1044 VDD.t1045 VDD.t60 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5969 VSS.t127 a_35502_25545.t93 a_33249_34067.t111 VSS.t39 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5970 VDD.t1043 VDD.t1041 VDD.t1043 VDD.t1042 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5971 VDD.t1040 VDD.t1039 VDD.t1040 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5972 VSS.t838 VSS.t836 VSS.t838 VSS.t837 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5973 VDD.t1038 VDD.t1037 VDD.t1038 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5974 a_112507_n6055.t0 a_71281_n8397.t309 a_112199_n9675# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5975 a_89715_n17715.t2 a_100992_4421.t1 a_113110_10448# VDD.t336 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5976 VDD.t1036 VDD.t1035 VDD.t1036 VDD.t619 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5977 a_52635_48695.t12 a_35922_19591.t164 a_52635_34067.t47 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5978 a_44885_n16007# a_31953_n19727.t336 a_44363_n16007.t0 VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5979 a_95943_n18620# a_71281_n10073.t311 a_95105_n18620# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5980 a_33249_48695.t148 a_33379_34007.t84 a_33249_34067.t26 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5981 VDD.t1034 VDD.t1033 VDD.t1034 VDD.t49 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5982 VDD.t1032 VDD.t1031 VDD.t1032 VDD.t6 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5983 VSS.t835 VSS.t833 VSS.t835 VSS.t834 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5984 a_84547_n6055# a_71281_n10073.t312 a_84017_n5150.t1 VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5985 a_52635_49681.t97 a_52635_34067.t225 VDD.t4815 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5986 VSS.t832 VSS.t831 VSS.t832 VSS.t571 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5987 a_95443_13546# a_81205_n14095.t9 a_89163_10388.t6 VDD.t497 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5988 a_33249_48695.t176 a_31699_20742.t245 VDD.t267 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5989 a_35221_n16904# a_31953_n19727.t337 a_34699_n16904# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5990 VSS.t830 VSS.t829 VSS.t830 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5991 VDD.t1030 VDD.t1029 VDD.t1030 VDD.t935 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5992 VDD.t268 a_31699_20742.t246 a_33249_48695.t175 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5993 VSS.t828 VSS.t827 VSS.t828 VSS.t671 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5994 VDD.t1028 VDD.t1027 VDD.t1028 VDD.t638 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5995 VDD.t1026 VDD.t1025 VDD.t1026 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5996 VDD.t1024 VDD.t1023 VDD.t1024 VDD.t962 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5997 VDD.t1022 VDD.t1021 VDD.t1022 VDD.t49 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5998 a_111063_n6960# a_71281_n8397.t310 a_110225_n6960# VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5999 a_33249_48695.t91 a_33379_34917.t81 a_33249_35053.t77 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6000 VSS.t826 VSS.t825 VSS.t826 VSS.t558 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6001 a_54229_n34390# a_53829_n36382.t21 a_53699_n35156.t0 VDD.t417 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6002 VSS.t824 VSS.t823 VSS.t824 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6003 a_83709_n2435# a_71281_n10073.t313 a_83141_n2435# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6004 a_94537_n18620# a_71281_n10073.t314 a_93969_n18620# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6005 a_95443_11614# a_81205_n14095.t10 a_89163_10388.t7 VDD.t497 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6006 a_111631_n1530# a_71281_n8397.t311 a_111063_n1530# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6007 VSS.t822 VSS.t821 VSS.t822 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6008 VDD.t1020 VDD.t1019 VDD.t1020 VDD.t792 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6009 VDD.t4750 a_65486_10448.t20 a_66016_13546# VDD.t1338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6010 VDD.t1018 VDD.t1017 VDD.t1018 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6011 OUT.t36 a_35922_19591.t165 a_52635_49681.t71 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6012 a_48951_4481.t2 a_47991_4421.t2 a_48391_4481# VSS.t340 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6013 VSS.t820 VSS.t819 VSS.t820 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6014 a_89009_4481.t3 a_89163_10388.t21 a_89563_10448# VDD.t554 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6015 VSS.t818 VSS.t816 VSS.t818 VSS.t817 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X6016 VDD.t1016 VDD.t1014 VDD.t1016 VDD.t1015 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6017 VDD.t1013 VDD.t1012 VDD.t1013 VDD.t598 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6018 VSS.t815 VSS.t813 VSS.t815 VSS.t814 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6019 VSS.t812 VSS.t810 VSS.t812 VSS.t811 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6020 a_60080_4481# a_59558_4481.t0 a_59558_4481.t1 VSS.t397 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6021 a_33249_48695.t174 a_31699_20742.t247 VDD.t269 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6022 a_40613_n19595# a_31953_n19727.t338 a_40053_n18698# VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6023 VSS.t58 a_31953_n19727.t4 a_31953_n19727.t5 VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6024 a_87433_n17715# a_71281_n10073.t315 a_86903_n21335# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6025 VSS.t809 VSS.t807 VSS.t809 VSS.t808 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6026 VDD.t4814 a_52635_34067.t226 a_52635_49681.t96 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6027 a_93131_n6055# a_71281_n10073.t316 a_92601_n9675# VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6028 VSS.t806 VSS.t805 VSS.t806 VSS.t99 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6029 VDD.t486 a_71281_n8397.t312 a_112199_n13190# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6030 VDD.t4813 a_52635_34067.t227 a_52635_49681.t95 VDD.t416 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6031 VSS.t804 VSS.t803 VSS.t804 VSS.t525 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6032 VDD.t4751 a_65486_10448.t21 a_66016_11614# VDD.t1338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6033 VDD.t1011 VDD.t1010 VDD.t1011 VDD.t38 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6034 a_40053_n19595# a_31953_n19727.t339 a_39179_n16007.t0 VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6035 VSS.t802 VSS.t801 VSS.t802 VSS.t149 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6036 VDD.t1009 VDD.t1008 VDD.t1009 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6037 a_101350_13546# a_100820_10448.t20 a_100820_11614.t3 VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6038 a_42047_n15110# a_31953_n19727.t340 a_41487_n14213# VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6039 a_41487_n5342# a_31953_n19727.t341 a_40613_n7136# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6040 a_35221_n4445# a_31953_n19727.t342 a_34699_n6239# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6041 VSS.t800 VSS.t799 VSS.t800 VSS.t522 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6042 a_33249_48695.t92 a_33379_34917.t82 a_33249_35053.t78 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6043 a_100803_n3340# a_71281_n8397.t313 a_100235_n3340# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6044 VDD.t1007 VDD.t1006 VDD.t1007 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6045 VDD.t1005 VDD.t1004 VDD.t1005 VDD.t82 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6046 VDD.t1003 VDD.t1002 VDD.t1003 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6047 VSS.t798 VSS.t797 VSS.t798 VSS.t411 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6048 VSS.t225 a_50751_n19729.t14 a_50751_n19729.t15 VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6049 VSS.t796 VSS.t794 VSS.t796 VSS.t795 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6050 a_42442_n35156# a_30324_n29313.t2 a_41891_n29181.t0 VDD.t560 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6051 a_57977_n8035# a_50751_n19729.t330 a_57417_n8035# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6052 VSS.t793 VSS.t791 VSS.t793 VSS.t792 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6053 a_96011_n36322.t0 a_89033_n35156.t11 a_95443_n34390# VDD.t2422 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6054 VSS.t790 VSS.t789 VSS.t790 VSS.t186 nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X6055 a_52635_48695.t11 a_35922_19591.t166 a_52635_34067.t48 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6056 VSS.t788 VSS.t787 VSS.t788 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6057 VDD.t1001 VDD.t1000 VDD.t1001 VDD.t290 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6058 a_95943_n6055# a_71281_n10073.t317 a_95413_n5150.t1 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6059 VSS.t786 VSS.t785 VSS.t786 VSS.t29 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6060 VDD.t999 VDD.t998 VDD.t999 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6061 VDD.t4812 a_52635_34067.t228 a_52635_49681.t94 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6062 a_51151_n7138# a_50751_n19729.t331 a_50629_n7138# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6063 VSS.t439 I1N.t16 a_72603_n10973# VSS.t433 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X6064 a_101350_11614# a_100820_10448.t21 a_100820_11614.t0 VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6065 VDD.t997 VDD.t996 VDD.t997 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6066 a_105933_n9675# a_71281_n8397.t314 a_105365_n9675# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6067 VSS.t784 VSS.t783 VSS.t784 VSS.t591 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6068 a_53145_n7138# a_50751_n19729.t332 a_52585_n7138# VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6069 VDD.t995 VDD.t993 VDD.t995 VDD.t994 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X6070 VDD.t992 VDD.t991 VDD.t992 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6071 VDD.t990 VDD.t989 VDD.t990 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6072 VDD.t988 VDD.t987 VDD.t988 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6073 a_42442_n33224# a_30324_n29313.t2 a_41891_n29181.t0 VDD.t560 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6074 a_33249_48695.t173 a_31699_20742.t248 VDD.t270 VDD.t78 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6075 VDD.t542 a_100820_n36322.t21 a_108602_n28415# VSS.t333 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6076 VSS.t782 VSS.t781 VSS.t782 VSS.t509 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6077 a_106501_n4245# a_71281_n8397.t315 a_105933_n4245# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6078 VSS.t135 a_35502_25545.t94 a_33249_34067.t110 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X6079 a_33249_35053.t110 a_35502_25545.t95 VSS.t143 VSS.t137 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6080 VSS.t780 VSS.t779 VSS.t780 VSS.t668 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6081 a_52635_49681.t93 a_52635_34067.t229 VDD.t4811 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6082 VDD.t986 VDD.t985 VDD.t986 VDD.t62 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6083 VSS.t778 VSS.t777 VSS.t778 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6084 VSS.t776 VSS.t774 VSS.t776 VSS.t775 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6085 VDD.t984 VDD.t983 VDD.t984 VDD.t748 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6086 VSS.t773 VSS.t771 VSS.t773 VSS.t772 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6087 a_95105_n2435# a_71281_n10073.t318 a_94537_n2435# VDD.t314 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6088 VSS.t327 a_77225_4481.t21 a_77747_4481# VSS.t323 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6089 OUT.t109 a_33379_34917.t0 cap_mim_2f0_m4m5_noshield c_width=9.8u c_length=9.8u
X6090 VDD.t982 VDD.t981 VDD.t982 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6091 VDD.t980 VDD.t978 VDD.t980 VDD.t979 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6092 VDD.t4810 a_52635_34067.t230 a_52635_48695.t93 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6093 a_85129_n27257# a_32913_n8930.t1 a_31831_n5342.t2 VSS.t286 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6094 VDD.t977 VDD.t975 VDD.t977 VDD.t976 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6095 VDD.t974 VDD.t973 VDD.t974 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6096 a_63161_n5344.t1 a_65658_4421.t0 a_66058_6405# VSS.t377 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6097 a_104527_n6055# a_71281_n8397.t316 a_103997_n9675# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6098 VDD.t972 VDD.t971 VDD.t972 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6099 a_112199_n14095# a_71281_n8397.t317 a_111631_n14095# VDD.t427 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6100 VSS.t770 VSS.t769 VSS.t770 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6101 VDD.t970 VDD.t969 VDD.t970 VDD.t55 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6102 VDD.t4761 a_30152_11614.t21 a_37934_6405# VSS.t281 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6103 VDD.t968 VDD.t967 VDD.t968 VDD.t725 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6104 a_47753_n3548# a_31953_n19727.t343 a_47231_n3548# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6105 VDD.t966 VDD.t964 VDD.t966 VDD.t965 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6106 a_87433_n21335# a_71281_n10073.t319 a_86903_n21335# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6107 VSS.t768 VSS.t767 VSS.t768 VSS.t168 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6108 VDD.t963 VDD.t961 VDD.t963 VDD.t962 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X6109 VSS.t766 VSS.t765 VSS.t766 VSS.t103 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6110 VDD.t960 VDD.t959 VDD.t960 VDD.t398 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6111 a_77747_6405# a_77225_4481.t2 a_77225_4481.t3 VSS.t317 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6112 VDD.t17 a_31699_20742.t5 a_31699_20742.t6 VDD.t16 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6113 VSS.t764 VSS.t762 VSS.t764 VSS.t763 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X6114 VDD.t958 VDD.t957 VDD.t958 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6115 a_33249_48695.t149 a_33379_34007.t85 a_33249_34067.t25 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6116 VSS.t761 VSS.t759 VSS.t761 VSS.t760 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6117 a_33249_48695.t93 a_33379_34917.t83 a_33249_35053.t79 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6118 VSS.t758 VSS.t756 VSS.t758 VSS.t757 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6119 VSS.t223 a_50751_n19729.t12 a_50751_n19729.t13 VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6120 OUT.t35 a_35922_19591.t167 a_52635_49681.t72 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6121 VSS.t755 VSS.t754 VSS.t755 VSS.t398 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6122 a_44363_n16007.t2 a_45445_n19595.t1 a_66058_n30339# VSS.t377 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6123 VDD.t956 VDD.t954 VDD.t956 VDD.t955 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6124 a_58851_n18700# a_50751_n19729.t333 a_58329_n18700# VSS.t229 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6125 a_39179_n14213# a_31953_n19727.t344 a_38619_n14213# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6126 a_52635_48695.t10 a_35922_19591.t168 a_52635_34067.t49 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6127 a_33249_48695.t172 a_31699_20742.t249 VDD.t271 VDD.t49 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6128 a_60845_n13318# a_50751_n19729.t334 a_60285_n13318# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6129 VDD.t272 a_31699_20742.t250 a_33249_48695.t171 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6130 a_89531_n27257# a_83153_n36322.t22 a_89009_n27257.t1 VSS.t454 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6131 a_102796_n29181# a_39179_n8930.t2 a_38097_n5342.t1 VSS.t330 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6132 VSS.t753 VSS.t752 VSS.t753 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6133 a_33787_n2651# a_31953_n19727.t345 a_33265_n3548# VSS.t68 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6134 a_50751_n19729.t11 a_50751_n19729.t10 VSS.t222 VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6135 VDD.t953 VDD.t952 VDD.t953 VDD.t930 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6136 VDD.t951 VDD.t950 VDD.t951 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6137 VDD.t323 a_100820_10448.t22 a_101350_10448# VDD.t293 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6138 a_61484_7563# a_59558_4481.t22 VSS.t408 VSS.t399 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6139 a_60109_12380# a_47991_4421.t1 a_59558_4481.t10 VDD.t2542 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6140 VDD.t949 VDD.t948 VDD.t949 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6141 a_35781_n17801# a_31953_n19727.t346 a_35221_n17801# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6142 a_52635_49681.t73 a_35922_19591.t169 OUT.t34 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6143 a_60285_n14215# a_50751_n19729.t335 a_59763_n14215# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6144 VDD.t4809 a_52635_34067.t231 a_52635_49681.t92 VDD.t410 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6145 OUT.t3 a_35502_24538.t62 a_33249_35053.t93 VSS.t193 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6146 a_113081_n30339# a_112559_n29181.t21 a_106830_n36382.t5 VSS.t410 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6147 VDD.t947 VDD.t946 VDD.t947 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6148 VSS.t751 VSS.t750 VSS.t751 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6149 VSS.t749 VSS.t747 VSS.t749 VSS.t748 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6150 a_106676_7563.t3 a_100820_11614.t22 a_108602_4481# VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6151 a_45445_n3548# a_31953_n19727.t347 a_44885_n2651# VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6152 a_30324_4421.t0 a_30152_11614.t22 a_36530_4481# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6153 VDD.t945 VDD.t943 VDD.t945 VDD.t944 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6154 a_38097_n16007.t2 a_47991_n29313.t2 a_48391_n27257# VSS.t340 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6155 a_32128_6405# a_30324_5507.t2 a_31284_4481.t2 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6156 VDD.t942 VDD.t941 VDD.t942 VDD.t407 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X6157 VDD.t940 VDD.t939 VDD.t940 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6158 a_64243_n3550# a_50751_n19729.t336 a_63683_n2653# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6159 VDD.t938 VDD.t937 VDD.t938 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6160 VDD.t936 VDD.t934 VDD.t936 VDD.t935 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6161 VDD.t933 VDD.t932 VDD.t933 VDD.t363 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6162 OUT.t33 a_35922_19591.t170 a_52635_49681.t74 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6163 VSS.t142 a_35502_25545.t96 a_33249_35053.t109 VSS.t21 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6164 a_95943_n17715# a_71281_n10073.t320 VDD.t386 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6165 VSS.t746 VSS.t744 VSS.t746 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6166 VDD.t931 VDD.t929 VDD.t931 VDD.t930 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6167 a_114516_13546# a_100992_4421.t1 a_89715_n17715.t1 VDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6168 VSS.t743 VSS.t742 VSS.t743 VSS.t618 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6169 VSS.t741 VSS.t739 VSS.t741 VSS.t740 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6170 a_110225_n8770# a_71281_n8397.t318 VDD.t487 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6171 a_84547_n6960# a_71281_n10073.t321 a_83709_n4245# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6172 VSS.t738 VSS.t737 VSS.t738 VSS.t401 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6173 a_54579_n13318# a_50751_n19729.t337 a_54019_n13318# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6174 a_40613_n2651# a_31953_n19727.t348 a_40053_n1754# VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6175 VDD.t928 VDD.t927 VDD.t928 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6176 a_33249_48695.t150 a_33379_34007.t86 a_33249_34067.t24 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6177 a_33249_34067.t23 a_33379_34007.t87 a_33249_48695.t151 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6178 a_47819_n35156.t10 a_47819_n35156.t9 a_49755_n34390# VDD.t2325 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6179 a_39179_n8930.t0 a_31953_n19727.t349 a_38619_n8930# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6180 a_52635_34067.t50 a_35922_19591.t171 a_52635_48695.t9 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6181 VDD.t926 VDD.t924 VDD.t926 VDD.t925 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6182 a_64243_n14215# a_50751_n19729.t338 a_63683_n13318# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6183 VDD.t923 VDD.t922 VDD.t923 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6184 a_110225_n19525# a_71281_n8397.t319 a_109695_n19525# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6185 a_33249_48695.t94 a_33379_34917.t84 a_33249_35053.t80 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6186 a_52635_34067.t41 a_35922_19591.t172 a_52635_48695.t8 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6187 VDD.t4808 a_52635_34067.t232 a_52635_49681.t91 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6188 a_33249_48695.t170 a_31699_20742.t251 VDD.t273 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6189 VSS.t736 VSS.t735 VSS.t736 VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6190 a_114516_11614# a_100992_4421.t1 a_89715_n17715.t4 VDD.t335 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6191 VSS.t375 a_41891_n29181.t22 a_42413_n28415# VSS.t166 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6192 VDD.t921 VDD.t919 VDD.t921 VDD.t920 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X6193 VDD.t918 VDD.t916 VDD.t918 VDD.t917 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6194 VDD.t915 VDD.t914 VDD.t915 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6195 VSS.t390 a_77225_n29181.t22 a_77747_n30339# VSS.t384 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6196 VDD.t491 a_71281_n10073.t2 a_71281_n10073.t3 VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6197 VSS.t734 VSS.t732 VSS.t734 VSS.t733 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6198 a_106676_7563.t1 a_106830_10388.t21 a_107230_13546# VDD.t519 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6199 a_33249_48695.t95 a_33379_34917.t85 a_33249_35053.t81 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6200 a_82573_n1530# a_71281_n10073.t322 a_81735_n1530# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6201 OUT.t1 a_106830_10388.t22 a_108636_10448# VDD.t521 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6202 VDD.t4798 a_47819_n35156.t21 a_48349_n34390# VDD.t2288 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6203 VSS.t731 VSS.t729 VSS.t731 VSS.t730 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6204 VDD.t913 VDD.t912 VDD.t913 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6205 a_46319_n12419# a_31953_n19727.t350 VSS.t121 VSS.t60 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6206 VDD.t911 VDD.t909 VDD.t911 VDD.t910 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6207 a_106501_n13190# a_71281_n8397.t320 a_105933_n13190# VDD.t425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6208 a_52635_49681.t75 a_35922_19591.t173 OUT.t32 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6209 VSS.t728 VSS.t727 VSS.t728 VSS.t106 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6210 a_99667_n1530# a_71281_n8397.t321 a_98829_n1530# VDD.t434 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6211 a_108602_4481# a_100820_11614.t23 a_100992_4421.t0 VSS.t147 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6212 a_57977_n14215# a_50751_n19729.t339 a_57417_n13318# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6213 a_38619_n8033# a_31953_n19727.t351 a_38097_n8930# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6214 a_36530_4481# a_30152_11614.t23 a_36008_4481.t1 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6215 VSS.t726 VSS.t725 VSS.t726 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6216 a_48349_n36322# a_47819_n35156.t22 a_47819_n36322.t1 VDD.t2559 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6217 a_101641_n6055# a_71281_n8397.t322 a_96011_n36322.t3 VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6218 a_30682_13546# a_30152_10448.t22 a_30152_11614.t7 VDD.t302 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6219 a_33249_34067.t109 a_35502_25545.t97 VSS.t141 VSS.t33 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6220 VDD.t908 VDD.t907 VDD.t908 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6221 a_77776_12380# a_65658_4421.t2 a_77225_4481.t8 VDD.t2924 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6222 a_55635_12380# a_53829_10388.t23 VSS.t420 VDD.t2921 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6223 a_33249_48695.t169 a_31699_20742.t252 VDD.t274 VDD.t134 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6224 VSS.t724 VSS.t723 VSS.t724 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6225 VSS.t722 VSS.t720 VSS.t722 VSS.t721 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6226 VSS.t316 a_106830_10388.t23 a_107230_11614# VDD.t519 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6227 VDD.t906 VDD.t904 VDD.t906 VDD.t905 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6228 VDD.t903 VDD.t902 VDD.t903 VDD.t548 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6229 VDD.t901 VDD.t900 VDD.t901 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6230 VDD.t899 VDD.t897 VDD.t899 VDD.t898 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6231 VSS.t719 VSS.t718 VSS.t719 VSS.t191 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X6232 VDD.t896 VDD.t895 VDD.t896 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6233 a_57977_n3550# a_50751_n19729.t340 a_57417_n3550# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6234 a_90245_n6960# a_71281_n10073.t323 a_89407_n6960# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6235 VDD.t894 VDD.t892 VDD.t894 VDD.t893 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6236 VSS.t717 VSS.t715 VSS.t717 VSS.t716 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6237 VDD.t891 VDD.t890 VDD.t891 VDD.t625 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6238 a_112559_4481.t1 a_112559_4481.t0 a_114485_5639# VSS.t292 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6239 VSS.t714 VSS.t712 VSS.t714 VSS.t713 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6240 VSS.t198 a_41891_4481.t20 a_42413_5639# VSS.t166 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6241 a_33249_34067.t0 a_35502_24538.t63 a_52635_34067.t59 VSS.t195 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6242 VSS.t711 VSS.t710 VSS.t711 VSS.t260 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6243 VSS.t709 VSS.t708 VSS.t709 VSS.t638 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6244 a_47991_5507.t1 a_47819_11614.t20 a_54197_6405# VSS.t304 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6245 a_71896_n34390# a_71496_n36382.t18 a_71366_n35156.t1 VDD.t2251 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6246 VDD.t889 VDD.t888 VDD.t889 VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6247 VSS.t707 VSS.t706 VSS.t707 VSS.t215 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6248 VDD.t887 VDD.t885 VDD.t887 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6249 VDD.t884 VDD.t882 VDD.t884 VDD.t883 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6250 VDD.t881 VDD.t880 VDD.t881 VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6251 a_83141_n14095# a_71281_n10073.t324 a_82573_n14095# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6252 a_90935_n29181# a_83153_n36322.t23 a_32913_n8930.t1 VSS.t452 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6253 a_100803_n2435# a_71281_n8397.t323 a_100235_n2435# VDD.t439 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6254 a_30682_11614# a_30152_10448.t23 a_30152_11614.t5 VDD.t302 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6255 VDD.t387 a_71281_n10073.t325 a_95105_n21335# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6256 VDD.t879 VDD.t877 VDD.t879 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6257 VSS.t705 VSS.t703 VSS.t705 VSS.t704 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6258 a_33249_34067.t108 a_35502_25545.t98 VSS.t140 VSS.t39 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6259 a_88839_n3340# a_71281_n10073.t326 a_88271_n3340# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6260 a_33379_34917.t68 IN_NEG.t0 cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
X6261 a_95943_n6960# a_71281_n10073.t327 a_95105_n4245# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6262 VDD.t876 VDD.t874 VDD.t876 VDD.t875 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6263 VSS.t139 a_35502_25545.t99 a_33249_34067.t107 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X6264 VSS.t702 VSS.t701 VSS.t702 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6265 VSS.t700 VSS.t698 VSS.t700 VSS.t699 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6266 VSS.t697 VSS.t696 VSS.t697 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6267 VSS.t695 VSS.t694 VSS.t695 VSS.t568 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6268 VDD.t873 VDD.t872 VDD.t873 VDD.t413 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6269 a_84547_n17715# a_71281_n10073.t328 a_84017_n16810.t0 VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6270 VSS.t693 VSS.t692 VSS.t693 VSS.t568 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6271 VSS.t691 VSS.t689 VSS.t691 VSS.t690 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6272 VSS.t688 VSS.t686 VSS.t688 VSS.t687 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6273 a_96849_n34390# a_83325_n29313.t1 a_96011_n36322.t0 VDD.t2240 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6274 OUT.t31 a_35922_19591.t174 a_52635_49681.t76 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6275 VSS.t685 VSS.t683 VSS.t685 VSS.t684 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6276 VSS.t682 VSS.t680 VSS.t682 VSS.t681 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6277 VDD.t871 VDD.t870 VDD.t871 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6278 a_33249_48695.t96 a_33379_34917.t86 a_33249_35053.t82 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6279 a_84547_n15000# a_71281_n10073.t329 a_83709_n15000# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6280 VDD.t869 VDD.t868 VDD.t869 VDD.t552 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6281 VDD.t867 VDD.t865 VDD.t867 VDD.t866 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6282 a_89009_n30339.t3 a_89163_n36382.t23 a_89563_n36322# VDD.t547 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6283 VSS.t679 VSS.t678 VSS.t679 VSS.t31 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6284 a_52635_34067.t42 a_35922_19591.t175 a_52635_48695.t7 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6285 a_71366_13546.t0 a_89163_10388.t22 a_90969_13546# VDD.t553 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6286 VDD.t864 VDD.t863 VDD.t864 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6287 a_81735_n14095# a_71281_n10073.t330 a_81205_n14095.t0 VDD.t310 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6288 a_71281_n10073.t1 a_71281_n10073.t0 VDD.t4976 VDD.t317 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6289 a_56895_n16009.t1 a_57977_n12421.t0 a_101392_5639# VSS.t162 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6290 VSS.t677 VSS.t675 VSS.t677 VSS.t676 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6291 VDD.t862 VDD.t861 VDD.t862 VDD.t289 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6292 VDD.t275 a_31699_20742.t253 a_33249_48695.t168 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6293 VDD.t860 VDD.t859 VDD.t860 VDD.t407 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X6294 a_94537_n21335# a_71281_n10073.t331 a_93969_n21335# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6295 a_47753_n18698# a_31953_n19727.t352 a_47231_n18698# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6296 a_52635_49681.t77 a_35922_19591.t176 OUT.t30 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6297 VDD.t858 VDD.t857 VDD.t858 VDD.t64 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6298 VDD.t4982 a_30152_n35156.t21 a_30682_n34390# VDD.t2228 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6299 VDD.t856 VDD.t854 VDD.t856 VDD.t855 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6300 VSS.t674 VSS.t673 VSS.t674 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6301 VSS.t672 VSS.t670 VSS.t672 VSS.t671 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6302 VDD.t853 VDD.t851 VDD.t853 VDD.t852 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6303 a_113081_5639# a_112559_4481.t22 a_106830_10388.t3 VSS.t293 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6304 a_52585_n8932# a_50751_n19729.t341 VSS.t279 VSS.t224 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6305 a_52635_48695.t6 a_35922_19591.t177 a_52635_34067.t51 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6306 VDD.t850 VDD.t849 VDD.t850 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6307 a_65486_10448.t9 a_65658_4421.t0 a_67462_5639# VSS.t378 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6308 VDD.t848 VDD.t847 VDD.t848 VDD.t49 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6309 VSS.t669 VSS.t667 VSS.t669 VSS.t668 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6310 VSS.t666 VSS.t665 VSS.t666 VSS.t609 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6311 a_111631_n19525# a_71281_n8397.t324 a_111063_n19525# VDD.t432 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6312 VDD.t846 VDD.t844 VDD.t846 VDD.t845 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6313 a_54579_n8932# a_50751_n19729.t342 a_54019_n8932# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6314 a_42413_5639# a_41891_4481.t21 a_36162_10388.t1 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6315 VDD.t843 VDD.t841 VDD.t843 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6316 VSS.t664 VSS.t663 VSS.t664 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6317 a_81205_n14095.t1 a_89163_10388.t23 a_90969_11614# VDD.t553 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6318 VDD.t840 VDD.t838 VDD.t840 VDD.t839 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6319 VDD.t837 VDD.t835 VDD.t837 VDD.t836 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6320 a_60285_n8035# a_50751_n19729.t343 a_59763_n8035# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6321 a_66016_n35156# a_65486_n35156.t2 a_65486_n35156.t3 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6322 VDD.t834 VDD.t832 VDD.t834 VDD.t833 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6323 VDD.t831 VDD.t830 VDD.t831 VDD.t64 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6324 VSS.t662 VSS.t661 VSS.t662 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6325 a_79151_5639# a_77225_4481.t22 VSS.t328 VSS.t319 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6326 VSS.t660 VSS.t659 VSS.t660 VSS.t186 nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X6327 VDD.t829 VDD.t827 VDD.t829 VDD.t828 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6328 a_52635_49681.t78 a_35922_19591.t178 OUT.t29 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6329 VSS.t658 VSS.t657 VSS.t658 VSS.t16 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6330 VSS.t656 VSS.t655 VSS.t656 VSS.t193 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6331 VSS.t654 VSS.t652 VSS.t654 VSS.t653 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6332 a_53699_n35156.t0 a_53829_n36382.t22 a_55635_n34390# VDD.t297 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6333 VSS.t651 VSS.t649 VSS.t651 VSS.t650 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6334 VSS.t648 VSS.t646 VSS.t648 VSS.t647 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6335 VDD.t826 VDD.t825 VDD.t826 VDD.t813 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6336 a_100992_n29313.t0 a_100820_n36322.t22 a_107198_n30339# VSS.t336 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6337 VDD.t824 VDD.t822 VDD.t824 VDD.t823 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6338 VDD.t821 VDD.t820 VDD.t821 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6339 VSS.t645 VSS.t643 VSS.t645 VSS.t644 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6340 a_33249_48695.t97 a_33379_34917.t87 a_33249_35053.t83 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6341 a_54197_n29181# a_47819_n36322.t23 VDD.t495 VSS.t306 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6342 VDD.t819 VDD.t817 VDD.t819 VDD.t818 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6343 VSS.t642 VSS.t640 VSS.t642 VSS.t641 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6344 VSS.t639 VSS.t637 VSS.t639 VSS.t638 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6345 VDD.t816 VDD.t815 VDD.t816 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6346 VDD.t814 VDD.t812 VDD.t814 VDD.t813 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6347 a_66016_n33224# a_65486_n35156.t0 a_65486_n35156.t1 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6348 VDD.t276 a_31699_20742.t254 a_33249_48695.t167 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6349 VDD.t811 VDD.t809 VDD.t811 VDD.t810 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6350 a_52635_34067.t52 a_35922_19591.t179 a_52635_48695.t5 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6351 OUT.t28 a_35922_19591.t180 a_52635_49681.t79 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6352 a_83141_n3340# a_71281_n10073.t332 a_82573_n3340# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6353 VDD.t808 VDD.t807 VDD.t808 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6354 a_67111_n7138# a_50751_n19729.t344 a_66551_n7138# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6355 VDD.t806 VDD.t805 VDD.t806 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6356 a_63683_n14215# a_50751_n19729.t345 a_63161_n15112# VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6357 VSS.t636 VSS.t635 VSS.t636 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6358 VDD.t804 VDD.t803 VDD.t804 VDD.t789 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6359 VSS.t634 VSS.t632 VSS.t634 VSS.t633 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6360 VSS.t631 VSS.t630 VSS.t631 VSS.t337 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6361 VDD.t802 VDD.t800 VDD.t802 VDD.t801 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6362 VDD.t799 VDD.t797 VDD.t799 VDD.t798 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6363 a_84547_n20430# a_71281_n10073.t333 a_83709_n20430# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6364 a_33249_35053.t84 a_33379_34917.t88 a_33249_48695.t98 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6365 a_53829_10388.t7 a_53699_11614.t10 a_61515_10448# VDD.t1512 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6366 OUT.t27 a_35922_19591.t181 a_52635_49681.t80 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6367 VSS.t629 VSS.t628 VSS.t629 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6368 a_100235_n3340# a_71281_n8397.t325 a_99667_n3340# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6369 VSS.t627 VSS.t626 VSS.t627 VSS.t353 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6370 a_33249_48695.t152 a_33379_34007.t88 a_33249_34067.t22 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6371 a_35502_25545.t8 a_31699_20742.t255 VDD.t277 VDD.t18 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6372 a_37934_n30339# a_30152_n36322.t23 a_30324_n29313.t0 VSS.t282 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6373 a_54229_n36322# a_53829_n36382.t23 a_53699_n36322.t0 VDD.t417 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6374 a_51151_n6241# a_50751_n19729.t346 a_50629_n7138# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6375 VSS.t625 VSS.t624 VSS.t625 VSS.t149 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6376 a_49795_7563# a_47991_4421.t0 a_48951_4481.t1 VSS.t338 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6377 a_110225_n7865# a_71281_n8397.t326 a_109695_n7865# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6378 a_108602_n29181# a_100820_n36322.t23 a_39179_n8930.t1 VSS.t334 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6379 a_88271_n9675# a_71281_n10073.t334 a_87433_n9675# VDD.t312 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6380 VDD.t796 VDD.t794 VDD.t796 VDD.t795 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6381 a_101641_n18620# a_71281_n8397.t327 a_100803_n18620# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6382 VDD.t793 VDD.t791 VDD.t793 VDD.t792 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6383 a_50751_n19729.t9 a_50751_n19729.t8 VSS.t221 VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6384 VSS.t623 VSS.t622 VSS.t623 VSS.t525 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6385 VDD.t790 VDD.t788 VDD.t790 VDD.t789 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6386 a_46879_n13316# a_31953_n19727.t353 a_46319_n13316# VSS.t65 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6387 VSS.t621 VSS.t620 VSS.t621 VSS.t378 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6388 a_32353_n18698# a_31953_n19727.t354 a_31831_n19595# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6389 VSS.t619 VSS.t617 VSS.t619 VSS.t618 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6390 VSS.t3636 a_59558_n29181.t22 a_60080_n27257# VSS.t401 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6391 a_36032_13546.t2 a_36162_10388.t23 a_37968_10448# VDD.t1494 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6392 VDD.t787 VDD.t786 VDD.t787 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6393 VSS.t616 VSS.t614 VSS.t616 VSS.t615 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6394 a_32913_n16007.t0 a_31953_n19727.t355 a_32353_n16007# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6395 VDD.t785 VDD.t784 VDD.t785 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6396 VSS.t613 VSS.t611 VSS.t613 VSS.t612 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6397 a_38619_n3548# a_31953_n19727.t356 a_38097_n4445# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6398 a_113037_n3340# a_71281_n8397.t328 a_112199_n3340# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6399 VSS.t610 VSS.t608 VSS.t610 VSS.t609 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6400 VDD.t783 VDD.t782 VDD.t783 VDD.t309 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6401 VDD.t781 VDD.t779 VDD.t781 VDD.t780 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6402 a_66016_12380# a_65486_10448.t0 a_65486_10448.t1 VDD.t2261 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6403 a_47753_n2651# a_31953_n19727.t357 a_47231_n3548# VSS.t102 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6404 a_47819_n35156.t0 a_47991_n29313.t0 a_49795_n28415# VSS.t337 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6405 a_75602_n3060# a_71266_n4019.t0 VDD.t4770 VDD.t692 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X6406 VSS.t607 VSS.t606 VSS.t607 VSS.t339 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6407 VSS.t605 VSS.t603 VSS.t605 VSS.t604 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6408 VSS.t602 VSS.t600 VSS.t602 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6409 VSS.t599 VSS.t598 VSS.t599 VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6410 VDD.t778 VDD.t777 VDD.t778 VDD.t538 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6411 VSS.t597 VSS.t595 VSS.t597 VSS.t596 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6412 VDD.t776 VDD.t775 VDD.t776 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6413 VDD.t774 VDD.t773 VDD.t774 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6414 a_73302_n35156# a_71496_n36382.t19 VSS.t366 VDD.t2812 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6415 VSS.t219 a_50751_n19729.t6 a_50751_n19729.t7 VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6416 a_65486_n35156.t7 a_65486_n35156.t6 a_67422_n34390# VDD.t1 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6417 a_101641_n6960# a_71281_n8397.t329 a_100803_n4245# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6418 a_96011_n36322.t2 a_89033_n35156.t12 a_95443_n36322# VDD.t2422 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6419 VSS.t594 VSS.t593 VSS.t594 VSS.t172 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6420 VDD.t772 VDD.t771 VDD.t772 VDD.t390 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X6421 OUT.t26 a_35922_19591.t182 a_52635_49681.t81 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6422 a_107339_n18620# a_71281_n8397.t330 a_106501_n18620# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6423 VDD.t770 VDD.t769 VDD.t770 VDD.t648 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6424 OUT.t25 a_35922_19591.t183 a_52635_49681.t82 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6425 VDD.t768 VDD.t767 VDD.t768 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6426 a_60845_n13318# a_50751_n19729.t347 a_60285_n12421# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6427 a_63683_n5344# a_50751_n19729.t348 a_63161_n5344.t0 VSS.t266 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6428 a_33249_48695.t153 a_33379_34007.t89 a_33249_34067.t21 VDD.t51 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6429 a_50751_n19729.t5 a_50751_n19729.t4 VSS.t218 VSS.t217 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6430 VDD.t766 VDD.t765 VDD.t766 VDD.t60 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6431 a_83153_n36322.t2 a_32913_n8930.t1 a_85129_n29181# VSS.t285 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6432 a_50751_n19729.t3 a_50751_n19729.t2 VSS.t216 VSS.t215 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6433 VDD.t764 VDD.t763 VDD.t764 VDD.t532 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6434 VDD.t506 a_47819_11614.t21 a_55601_5639# VSS.t307 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6435 VDD.t762 VDD.t761 VDD.t762 VDD.t406 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6436 VDD.t760 VDD.t759 VDD.t760 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6437 VDD.t758 VDD.t757 VDD.t758 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6438 VSS.t592 VSS.t590 VSS.t592 VSS.t591 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6439 a_57417_n19597# a_50751_n19729.t349 a_56895_n19597# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6440 VDD.t756 VDD.t754 VDD.t756 VDD.t755 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6441 a_33249_48695.t99 a_33379_34917.t89 a_33249_35053.t85 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6442 VSS.t363 a_94892_n29181.t21 a_95414_n30339# VSS.t357 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6443 a_73302_n33224# a_71496_n36382.t20 a_71342_n30339.t1 VDD.t2812 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6444 VDD.t278 a_31699_20742.t256 a_35502_24538.t2 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6445 VDD.t753 VDD.t752 VDD.t753 VDD.t537 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6446 VDD.t751 VDD.t750 VDD.t751 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6447 VSS.t589 VSS.t587 VSS.t589 VSS.t588 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6448 a_101392_n28415# a_39179_n8930.t1 a_100820_n36322.t6 VSS.t331 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6449 VSS.t586 VSS.t584 VSS.t586 VSS.t585 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6450 a_33249_48695.t166 a_31699_20742.t257 VDD.t279 VDD.t64 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6451 VSS.t583 VSS.t582 VSS.t583 VSS.t27 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6452 VSS.t581 VSS.t580 VSS.t581 VSS.t5 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X6453 VDD.t4807 a_52635_34067.t233 a_52635_49681.t90 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6454 VDD.t11 a_65486_n35156.t23 a_66016_n34390# VDD.t2 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6455 VDD.t749 VDD.t747 VDD.t749 VDD.t748 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6456 VSS.t579 VSS.t578 VSS.t579 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6457 VSS.t577 VSS.t575 VSS.t577 VSS.t576 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6458 a_60845_n4447# a_50751_n19729.t350 a_60285_n4447# VSS.t262 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6459 VSS.t574 VSS.t573 VSS.t574 VSS.t498 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6460 VDD.t746 VDD.t744 VDD.t746 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6461 VDD.t743 VDD.t741 VDD.t743 VDD.t742 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6462 VDD.t740 VDD.t739 VDD.t740 VDD.t307 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6463 a_88839_n2435# a_71281_n10073.t335 a_88271_n2435# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6464 VDD.t738 VDD.t737 VDD.t738 VDD.t427 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6465 VDD.t736 VDD.t735 VDD.t736 VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6466 VDD.t734 VDD.t733 VDD.t734 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6467 VDD.t732 VDD.t731 VDD.t732 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6468 VSS.t572 VSS.t570 VSS.t572 VSS.t571 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6469 a_54579_n13318# a_50751_n19729.t351 a_54019_n12421# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6470 a_84547_n18620# a_71281_n10073.t336 a_83709_n15905# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6471 VDD.t730 VDD.t729 VDD.t730 VDD.t520 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6472 VDD.t728 VDD.t727 VDD.t728 VDD.t529 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6473 IBNOUT.t0 a_50751_n19729.t352 a_63683_n12421# VSS.t263 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6474 a_90935_7563# a_83153_11614.t23 a_83325_4421.t0 VSS.t395 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6475 VDD.t726 VDD.t724 VDD.t726 VDD.t725 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6476 VDD.t723 VDD.t722 VDD.t723 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6477 VDD.t721 VDD.t719 VDD.t721 VDD.t720 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6478 VDD.t718 VDD.t717 VDD.t718 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6479 VDD.t716 VDD.t715 VDD.t716 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6480 VDD.t714 VDD.t713 VDD.t714 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6481 VDD.t712 VDD.t711 VDD.t712 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6482 a_54019_n8932# a_50751_n19729.t353 a_51711_n8932# VSS.t264 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6483 VSS.t569 VSS.t567 VSS.t569 VSS.t568 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6484 a_42413_n29181# a_41891_n29181.t3 a_41891_n29181.t4 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6485 VDD.t710 VDD.t709 VDD.t710 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6486 VSS.t566 VSS.t565 VSS.t566 VSS.t14 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6487 VSS.t564 VSS.t563 VSS.t564 VSS.t191 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X6488 a_60285_n3550# a_50751_n19729.t354 a_59763_n3550# VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6489 a_83683_12380# a_83153_10448.t6 a_83153_10448.t7 VDD.t2774 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6490 VDD.t708 VDD.t706 VDD.t708 VDD.t707 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6491 VDD.t705 VDD.t704 VDD.t705 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6492 VSS.t562 VSS.t560 VSS.t562 VSS.t561 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6493 VDD.t703 VDD.t702 VDD.t703 VDD.t555 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6494 VDD.t280 a_31699_20742.t258 a_33249_48695.t165 VDD.t55 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6495 VSS.t559 VSS.t557 VSS.t559 VSS.t558 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6496 VSS.t556 VSS.t555 VSS.t556 VSS.t553 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6497 a_52635_48695.t4 a_35922_19591.t184 a_52635_34067.t53 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6498 a_35221_n12419# a_31953_n19727.t358 a_32913_n12419# VSS.t108 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6499 VDD.t701 VDD.t699 VDD.t701 VDD.t700 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6500 VDD.t281 a_31699_20742.t259 a_33249_48695.t164 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6501 VSS.t554 VSS.t552 VSS.t554 VSS.t553 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6502 a_66058_7563# a_64243_n1756.t1 a_65486_11614.t4 VSS.t376 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6503 OUT.t24 a_35922_19591.t185 a_52635_49681.t83 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6504 VDD.t698 VDD.t696 VDD.t698 VDD.t697 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6505 VSS.t551 VSS.t549 VSS.t551 VSS.t550 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6506 a_32088_n34390# a_30152_n35156.t22 VDD.t4983 VDD.t2088 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6507 a_105365_n8770# a_71281_n8397.t331 a_104527_n8770# VDD.t429 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6508 VSS.t548 VSS.t547 VSS.t548 VSS.t220 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6509 VSS.t546 VSS.t544 VSS.t546 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6510 VDD.t282 a_31699_20742.t260 a_33249_48695.t163 VDD.t70 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6511 VDD.t695 VDD.t694 VDD.t695 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6512 VDD.t4806 a_52635_34067.t234 a_52635_48695.t92 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6513 a_48313_n17801# a_31953_n19727.t359 a_47753_n17801# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6514 a_114485_n28415# a_112559_n29181.t22 VSS.t3648 VSS.t413 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6515 a_55601_5639# a_47819_11614.t22 a_47991_5507.t1 VSS.t305 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6516 VDD.t283 a_31699_20742.t261 a_33249_48695.t162 VDD.t62 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6517 a_33249_34067.t20 a_33379_34007.t90 a_33249_48695.t154 VDD.t82 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6518 a_89163_n36382.t3 a_94892_n29181.t22 a_96818_n29181# VSS.t352 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6519 a_52635_34067.t54 a_35922_19591.t186 a_52635_48695.t3 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6520 a_105933_n3340# a_71281_n8397.t332 a_105365_n3340# VDD.t442 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6521 a_57977_n12421.t1 a_50751_n19729.t355 a_57417_n12421# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6522 VDD.t693 VDD.t691 VDD.t693 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X6523 a_33249_48695.t100 a_33379_34917.t90 a_33249_35053.t86 VDD.t53 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6524 VDD.t690 VDD.t688 VDD.t690 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6525 VDD.t687 VDD.t685 VDD.t687 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6526 VDD.t684 VDD.t682 VDD.t684 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6527 VDD.t681 VDD.t679 VDD.t681 VDD.t680 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6528 VSS.t543 VSS.t542 VSS.t543 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6529 VDD.t15 a_31699_20742.t3 a_31699_20742.t4 VDD.t14 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6530 VSS.t541 VSS.t539 VSS.t541 VSS.t540 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6531 VDD.t678 VDD.t676 VDD.t678 VDD.t677 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6532 a_57977_n3550# a_50751_n19729.t356 a_57417_n2653# VSS.t265 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6533 VSS.t538 VSS.t536 VSS.t538 VSS.t537 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6534 VSS.t535 VSS.t533 VSS.t535 VSS.t534 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6535 VDD.t675 VDD.t673 VDD.t675 VDD.t674 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6536 VDD.t424 a_71281_n8397.t0 a_71281_n8397.t1 VDD.t423 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6537 VDD.t672 VDD.t671 VDD.t672 VDD.t290 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6538 OUT.t23 a_35922_19591.t187 a_52635_49681.t84 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6539 VSS.t532 VSS.t530 VSS.t532 VSS.t531 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6540 a_47819_n35156.t6 a_47819_n35156.t5 a_49755_n36322# VDD.t2325 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6541 a_52635_34067.t55 a_35922_19591.t188 a_52635_48695.t2 VDD.t393 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6542 a_51151_n1756# a_50751_n19729.t357 a_50629_n2653# VSS.t261 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6543 VSS.t529 VSS.t527 VSS.t529 VSS.t528 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6544 VDD.t670 VDD.t669 VDD.t670 VDD.t326 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6545 VSS.t526 VSS.t524 VSS.t526 VSS.t525 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6546 VSS.t523 VSS.t521 VSS.t523 VSS.t522 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6547 VSS.t520 VSS.t519 VSS.t520 VSS.t65 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6548 a_83141_n2435# a_71281_n10073.t337 a_82573_n2435# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6549 VSS.t518 VSS.t517 VSS.t518 VSS.t260 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6550 a_52635_34067.t43 a_35922_19591.t189 a_52635_48695.t1 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6551 a_53145_n2653# a_50751_n19729.t358 a_52585_n1756# VSS.t220 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6552 VDD.t668 VDD.t666 VDD.t668 VDD.t667 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6553 VDD.t665 VDD.t663 VDD.t665 VDD.t664 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6554 VSS.t516 VSS.t515 VSS.t516 VSS.t478 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6555 a_52635_49681.t85 a_35922_19591.t190 OUT.t22 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6556 a_83683_n35156# a_83153_n35156.t2 a_83153_n35156.t3 VDD.t2729 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6557 a_100235_n2435# a_71281_n8397.t333 a_99667_n2435# VDD.t444 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6558 VDD.t662 VDD.t660 VDD.t662 VDD.t661 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6559 VDD.t4805 a_52635_34067.t235 a_52635_49681.t89 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6560 VSS.t514 VSS.t513 VSS.t514 VSS.t282 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6561 a_71366_n35156.t3 a_71496_n36382.t21 a_73302_n34390# VDD.t2058 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6562 VSS.t512 VSS.t511 VSS.t512 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6563 VDD.t659 VDD.t658 VDD.t659 VDD.t638 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6564 VSS.t510 VSS.t508 VSS.t510 VSS.t509 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6565 VSS.t507 VSS.t505 VSS.t507 VSS.t506 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6566 a_33249_35053.t108 a_35502_25545.t100 VSS.t138 VSS.t137 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6567 a_52635_48695.t91 a_52635_34067.t236 VDD.t4804 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6568 a_52635_48695.t90 a_52635_34067.t237 VDD.t4803 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6569 VDD.t657 VDD.t655 VDD.t657 VDD.t656 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6570 VDD.t517 a_47819_10448.t22 a_48349_10448# VDD.t510 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6571 a_33249_48695.t161 a_31699_20742.t262 VDD.t284 VDD.t68 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6572 a_66551_n8932# a_50751_n19729.t359 a_64243_n8932# VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6573 VDD.t654 VDD.t652 VDD.t654 VDD.t653 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6574 VSS.t136 a_35502_25545.t101 a_33249_34067.t106 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X6575 VSS.t504 VSS.t503 VSS.t504 VSS.t309 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6576 a_60080_n29181# a_59558_n29181.t9 a_59558_n29181.t10 VSS.t397 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6577 VSS.t502 VSS.t500 VSS.t502 VSS.t501 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6578 VSS.t499 VSS.t497 VSS.t499 VSS.t498 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6579 a_101641_n17715# a_71281_n8397.t334 a_101111_n17715.t1 VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6580 VDD.t4799 a_47819_n35156.t23 a_48349_n36322# VDD.t2288 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6581 VDD.t651 VDD.t650 VDD.t651 VDD.t619 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6582 VSS.t496 VSS.t494 VSS.t496 VSS.t495 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6583 a_33249_35053.t99 a_35502_24538.t64 OUT.t2 VSS.t195 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6584 a_52635_49681.t86 a_35922_19591.t191 OUT.t21 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6585 VSS.t493 VSS.t492 VSS.t493 VSS.t333 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6586 VDD.t649 VDD.t647 VDD.t649 VDD.t648 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6587 a_78344_n36322.t2 a_71366_n35156.t12 a_77776_n34390# VDD.t502 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6588 VDD.t646 VDD.t645 VDD.t646 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6589 VSS.t491 VSS.t489 VSS.t491 VSS.t490 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6590 a_83683_n33224# a_83153_n35156.t6 a_83153_n35156.t7 VDD.t2729 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6591 VSS.t488 VSS.t486 VSS.t488 VSS.t487 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6592 VDD.t644 VDD.t642 VDD.t644 VDD.t643 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6593 a_33249_48695.t155 a_33379_34007.t91 a_33249_34067.t19 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6594 VDD.t641 VDD.t640 VDD.t641 VDD.t66 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6595 VSS.t485 VSS.t483 VSS.t485 VSS.t484 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X6596 VDD.t639 VDD.t637 VDD.t639 VDD.t638 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6597 VDD.t636 VDD.t634 VDD.t636 VDD.t635 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6598 VSS.t482 VSS.t480 VSS.t482 VSS.t481 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6599 VSS.t479 VSS.t477 VSS.t479 VSS.t478 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6600 a_65486_n36322.t4 a_45445_n19595.t1 a_67462_n27257# VSS.t378 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6601 VSS.t476 VSS.t474 VSS.t476 VSS.t475 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6602 a_67111_n17803# a_50751_n19729.t360 a_66551_n16906# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6603 VDD.t633 VDD.t632 VDD.t633 VDD.t598 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6604 VDD.t631 VDD.t629 VDD.t631 VDD.t630 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6605 VSS.t367 a_71496_n36382.t22 a_71896_n34390# VDD.t2021 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6606 a_113037_n3340# a_71281_n8397.t335 a_112199_n2435# VDD.t472 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6607 VDD.t628 VDD.t627 VDD.t628 VDD.t398 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6608 a_33249_48695.t101 a_33379_34917.t91 a_33249_35053.t87 VDD.t96 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6609 VDD.t626 VDD.t624 VDD.t626 VDD.t625 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6610 a_52635_34067.t34 a_35922_19591.t192 a_52635_48695.t0 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6611 VDD.t623 VDD.t621 VDD.t623 VDD.t622 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6612 VDD.t620 VDD.t618 VDD.t620 VDD.t619 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6613 a_71896_n36322# a_71496_n36382.t23 a_71366_n36322.t1 VDD.t2251 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6614 VDD.t617 VDD.t615 VDD.t617 VDD.t616 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6615 a_33249_48695.t160 a_31699_20742.t263 VDD.t285 VDD.t76 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6616 VSS.t473 VSS.t471 VSS.t473 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6617 VDD.t4802 a_52635_34067.t238 a_52635_49681.t88 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6618 VSS.t214 a_50751_n19729.t0 a_50751_n19729.t1 VSS.t213 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6619 VSS.t470 VSS.t469 VSS.t470 VSS.t157 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6620 VDD.t614 VDD.t612 VDD.t614 VDD.t613 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6621 a_33249_48695.t159 a_31699_20742.t264 VDD.t286 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6622 VDD.t611 VDD.t609 VDD.t611 VDD.t610 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6623 a_95443_10448# a_83325_4421.t1 a_94892_4481.t8 VDD.t497 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6624 VDD.t608 VDD.t607 VDD.t608 VDD.t352 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6625 VDD.t606 VDD.t605 VDD.t606 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6626 VDD.t4801 a_52635_34067.t239 a_52635_48695.t89 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6627 VDD.t604 VDD.t602 VDD.t604 VDD.t603 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6628 VDD.t601 VDD.t600 VDD.t601 VDD.t64 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6629 a_107339_n17715# a_71281_n8397.t336 a_106809_n17715.t0 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6630 VDD.t599 VDD.t597 VDD.t599 VDD.t598 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6631 a_94892_n29181.t0 a_83325_n29313.t1 a_96849_n34390# VDD.t1996 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6632 a_38619_n16904# a_31953_n19727.t360 a_38097_n17801# VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6633 a_31699_20742.t2 a_31699_20742.t1 VDD.t13 VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6634 a_36162_10388.t0 a_41891_4481.t22 a_43817_6405# VSS.t168 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6635 VDD.t596 VDD.t595 VDD.t596 VDD.t367 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6636 VDD.t594 VDD.t592 VDD.t594 VDD.t593 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6637 VSS.t468 VSS.t466 VSS.t468 VSS.t467 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6638 VSS.t465 VSS.t463 VSS.t465 VSS.t464 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6639 a_96849_n36322# a_83325_n29313.t1 a_96011_n36322.t2 VDD.t2240 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6640 VDD.t591 VDD.t590 VDD.t591 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6641 a_54197_7563# a_47819_11614.t23 a_53675_7563.t3 VSS.t306 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6642 VDD.t589 VDD.t588 VDD.t589 VDD.t341 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6643 a_71266_n4019.t0 I1N.t17 a_75585_n10073# VSS.t312 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X6644 VSS.t462 VSS.t461 VSS.t462 VSS.t150 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6645 a_31953_n19727.t3 a_31953_n19727.t2 VSS.t57 VSS.t56 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6646 VSS.t460 VSS.t458 VSS.t460 VSS.t459 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6647 a_59558_n29181.t6 a_59558_n29181.t5 a_61484_n28415# VSS.t398 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6648 VSS.t144 a_35502_25545.t102 a_33249_35053.t107 VSS.t21 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6649 a_33249_48695.t156 a_33379_34007.t92 a_33249_34067.t18 VDD.t60 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6650 a_67111_n7138# a_50751_n19729.t361 a_66551_n6241# VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6651 VDD.t587 VDD.t585 VDD.t587 VDD.t586 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6652 VDD.t584 VDD.t582 VDD.t584 VDD.t583 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6653 VDD.t581 VDD.t580 VDD.t581 VDD.t335 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6654 a_33249_35053.t106 a_35502_25545.t103 VSS.t146 VSS.t145 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6655 VDD.t579 VDD.t578 VDD.t579 VDD.t439 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6656 a_52635_49681.t87 a_35922_19591.t193 OUT.t20 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6657 VDD.t577 VDD.t576 VDD.t577 VDD.t543 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6658 VDD.t4752 a_65486_10448.t22 a_66016_10448# VDD.t1338 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6659 VDD.t4984 a_30152_n35156.t23 a_30682_n36322# VDD.t2228 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6660 VDD.t575 VDD.t573 VDD.t575 VDD.t574 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6661 VSS.t55 a_31953_n19727.t0 a_31953_n19727.t1 VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6662 VDD.t572 VDD.t570 VDD.t572 VDD.t571 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6663 VDD.t569 VDD.t567 VDD.t569 VDD.t568 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X6664 VDD.t566 VDD.t565 VDD.t566 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6665 a_101111_n17715.t0 a_71281_n8397.t337 a_100803_n21335# VDD.t474 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6666 VSS.t457 VSS.t456 VSS.t457 VSS.t107 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6667 VDD.t4800 a_52635_34067.t240 a_52635_48695.t88 VDD.t406 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6668 VDD.t564 VDD.t562 VDD.t564 VDD.t563 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6669 a_35781_n13316# a_31953_n19727.t361 a_35221_n13316# VSS.t107 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6670 VDD.t561 VDD.t559 VDD.t561 VDD.t560 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6671 VDD.t558 VDD.t556 VDD.t558 VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
R0 VSS.n11299 VSS.n132 320062
R1 VSS.n10846 VSS.n10697 144034
R2 VSS.n11300 VSS.n11299 49361.9
R3 VSS.n9304 VSS.n9302 17249
R4 VSS.n10287 VSS.n132 12232.4
R5 VSS.n10697 VSS.n10287 9171.32
R6 VSS.n10861 VSS.n244 3502.89
R7 VSS.n11301 VSS.t763 757.145
R8 VSS.n11296 VSS.n11293 752.225
R9 VSS.n11285 VSS.n11280 752.225
R10 VSS.n563 VSS.n562 752.225
R11 VSS.n10065 VSS.n512 752.225
R12 VSS.n9891 VSS.n644 752.225
R13 VSS.n10116 VSS.n440 752.225
R14 VSS.n139 VSS.n135 752.225
R15 VSS.n11278 VSS.n144 752.225
R16 VSS.n568 VSS.n564 752.225
R17 VSS.n1181 VSS.n510 752.225
R18 VSS.n9765 VSS.n646 752.225
R19 VSS.n1235 VSS.n438 752.225
R20 VSS.n11296 VSS.n136 750.567
R21 VSS.n11285 VSS.n145 750.567
R22 VSS.n10033 VSS.n562 750.567
R23 VSS.n512 VSS.n508 750.567
R24 VSS.n9891 VSS.n645 750.567
R25 VSS.n440 VSS.n436 750.567
R26 VSS.n11291 VSS.n135 750.567
R27 VSS.n149 VSS.n144 750.567
R28 VSS.n10031 VSS.n568 750.567
R29 VSS.n1181 VSS.n509 750.567
R30 VSS.n9767 VSS.n646 750.567
R31 VSS.n1235 VSS.n437 750.567
R32 VSS.n11293 VSS.n137 750.383
R33 VSS.n11280 VSS.n146 750.383
R34 VSS.n563 VSS.n561 750.383
R35 VSS.n10065 VSS.n511 750.383
R36 VSS.n9522 VSS.n644 750.383
R37 VSS.n10116 VSS.n439 750.383
R38 VSS.n11290 VSS.n139 750.383
R39 VSS.n11278 VSS.n150 750.383
R40 VSS.n567 VSS.n564 750.383
R41 VSS.n9888 VSS.n510 750.383
R42 VSS.n9765 VSS.n797 750.383
R43 VSS.n1389 VSS.n438 750.383
R44 VSS.n137 VSS.n136 748.725
R45 VSS.n146 VSS.n145 748.725
R46 VSS.n10033 VSS.n561 748.725
R47 VSS.n511 VSS.n508 748.725
R48 VSS.n9522 VSS.n645 748.725
R49 VSS.n439 VSS.n436 748.725
R50 VSS.n11291 VSS.n11290 748.725
R51 VSS.n150 VSS.n149 748.725
R52 VSS.n10031 VSS.n567 748.725
R53 VSS.n9888 VSS.n509 748.725
R54 VSS.n9767 VSS.n797 748.725
R55 VSS.n1389 VSS.n437 748.725
R56 VSS.n9464 VSS.n1381 697.422
R57 VSS.n9466 VSS.n1382 693.922
R58 VSS.n9464 VSS.n1382 693.645
R59 VSS.n9466 VSS.n1381 688.856
R60 VSS.t817 VSS.n10847 684.903
R61 VSS.n10598 VSS.n10344 661.869
R62 VSS.n10695 VSS.n10289 661.869
R63 VSS.n10664 VSS.n10340 661.869
R64 VSS.n10661 VSS.n10343 656.895
R65 VSS.n10603 VSS.n10288 656.895
R66 VSS.n10342 VSS.n10341 656.895
R67 VSS.n10661 VSS.n10344 656.434
R68 VSS.n10603 VSS.n10289 656.434
R69 VSS.n10664 VSS.n10341 656.434
R70 VSS.n10598 VSS.n10343 653.672
R71 VSS.n10695 VSS.n10288 653.672
R72 VSS.n10342 VSS.n10340 653.672
R73 VSS.n10849 VSS.n10848 613.597
R74 VSS.n11302 VSS.n130 531.539
R75 VSS.n10845 VSS.n130 530.25
R76 VSS.n11302 VSS.n131 530.067
R77 VSS.n10845 VSS.n131 528.777
R78 VSS.n11346 VSS.n8 523.342
R79 VSS.n11360 VSS.n95 523.342
R80 VSS.n10983 VSS.n183 523.342
R81 VSS.n10928 VSS.n220 523.342
R82 VSS.n867 VSS.n505 523.342
R83 VSS.n9562 VSS.n835 523.342
R84 VSS.n11375 VSS.n5 523.342
R85 VSS.n11362 VSS.n92 523.342
R86 VSS.n10981 VSS.n180 523.342
R87 VSS.n10930 VSS.n216 523.342
R88 VSS.n1185 VSS.n1153 523.342
R89 VSS.n9541 VSS.n832 523.342
R90 VSS.n9528 VSS.n9527 523.342
R91 VSS.n9421 VSS.n1395 523.342
R92 VSS.n432 VSS.n431 523.342
R93 VSS.n10122 VSS.n421 523.342
R94 VSS.n420 VSS.n393 523.342
R95 VSS.n362 VSS.n361 523.342
R96 VSS.n10182 VSS.n349 523.342
R97 VSS.n348 VSS.n321 523.342
R98 VSS.n290 VSS.n289 523.342
R99 VSS.n10242 VSS.n277 523.342
R100 VSS.n276 VSS.n251 523.342
R101 VSS.n9117 VSS.n1532 523.342
R102 VSS.n9093 VSS.n1537 523.342
R103 VSS.n9009 VSS.n1563 523.342
R104 VSS.n9348 VSS.n1482 523.342
R105 VSS.n9298 VSS.n1507 523.342
R106 VSS.n9250 VSS.n1515 523.342
R107 VSS.n9176 VSS.n1525 523.342
R108 VSS.n11467 VSS.n7 521.869
R109 VSS.n11037 VSS.n94 521.869
R110 VSS.n11151 VSS.n182 521.869
R111 VSS.n547 VSS.n219 521.869
R112 VSS.n10068 VSS.n504 521.869
R113 VSS.n9563 VSS.n834 521.869
R114 VSS.n11469 VSS.n4 521.869
R115 VSS.n11263 VSS.n91 521.869
R116 VSS.n11153 VSS.n179 521.869
R117 VSS.n693 VSS.n215 521.869
R118 VSS.n9559 VSS.n507 521.869
R119 VSS.n9565 VSS.n831 521.869
R120 VSS.n1222 VSS.n435 521.869
R121 VSS.n9381 VSS.n1384 521.869
R122 VSS.n10120 VSS.n10119 521.869
R123 VSS.n10127 VSS.n422 521.869
R124 VSS.n10175 VSS.n394 521.869
R125 VSS.n10180 VSS.n10179 521.869
R126 VSS.n10187 VSS.n350 521.869
R127 VSS.n10235 VSS.n322 521.869
R128 VSS.n10240 VSS.n10239 521.869
R129 VSS.n10247 VSS.n278 521.869
R130 VSS.n10285 VSS.n252 521.869
R131 VSS.n9111 VSS.n1531 521.869
R132 VSS.n9090 VSS.n1555 521.869
R133 VSS.n9014 VSS.n1562 521.869
R134 VSS.n9345 VSS.n1497 521.869
R135 VSS.n9308 VSS.n1506 521.869
R136 VSS.n9247 VSS.n1514 521.869
R137 VSS.n9181 VSS.n1524 521.869
R138 VSS.n11346 VSS.n7 519.659
R139 VSS.n11360 VSS.n94 519.659
R140 VSS.n10983 VSS.n182 519.659
R141 VSS.n10928 VSS.n219 519.659
R142 VSS.n867 VSS.n504 519.659
R143 VSS.n835 VSS.n834 519.659
R144 VSS.n11375 VSS.n4 519.659
R145 VSS.n11362 VSS.n91 519.659
R146 VSS.n10981 VSS.n179 519.659
R147 VSS.n10930 VSS.n215 519.659
R148 VSS.n9559 VSS.n1153 519.659
R149 VSS.n9541 VSS.n831 519.659
R150 VSS.n9528 VSS.n1222 519.659
R151 VSS.n9421 VSS.n1384 519.659
R152 VSS.n10120 VSS.n431 519.659
R153 VSS.n10127 VSS.n421 519.659
R154 VSS.n10175 VSS.n393 519.659
R155 VSS.n10180 VSS.n361 519.659
R156 VSS.n10187 VSS.n349 519.659
R157 VSS.n10235 VSS.n321 519.659
R158 VSS.n10240 VSS.n289 519.659
R159 VSS.n10247 VSS.n277 519.659
R160 VSS.n10285 VSS.n251 519.659
R161 VSS.n9111 VSS.n1532 519.659
R162 VSS.n9093 VSS.n1555 519.659
R163 VSS.n9009 VSS.n1562 519.659
R164 VSS.n9348 VSS.n1497 519.659
R165 VSS.n9298 VSS.n1506 519.659
R166 VSS.n9250 VSS.n1514 519.659
R167 VSS.n9176 VSS.n1524 519.659
R168 VSS.n11467 VSS.n8 516.342
R169 VSS.n11037 VSS.n95 516.342
R170 VSS.n11151 VSS.n183 516.342
R171 VSS.n547 VSS.n220 516.342
R172 VSS.n10068 VSS.n505 516.342
R173 VSS.n9563 VSS.n9562 516.342
R174 VSS.n11469 VSS.n5 516.342
R175 VSS.n11263 VSS.n92 516.342
R176 VSS.n11153 VSS.n180 516.342
R177 VSS.n693 VSS.n216 516.342
R178 VSS.n1185 VSS.n507 516.342
R179 VSS.n9565 VSS.n832 516.342
R180 VSS.n9527 VSS.n435 516.342
R181 VSS.n9381 VSS.n1395 516.342
R182 VSS.n10119 VSS.n432 516.342
R183 VSS.n10122 VSS.n422 516.342
R184 VSS.n420 VSS.n394 516.342
R185 VSS.n10179 VSS.n362 516.342
R186 VSS.n10182 VSS.n350 516.342
R187 VSS.n348 VSS.n322 516.342
R188 VSS.n10239 VSS.n290 516.342
R189 VSS.n10242 VSS.n278 516.342
R190 VSS.n276 VSS.n252 516.342
R191 VSS.n9117 VSS.n1531 516.342
R192 VSS.n9090 VSS.n1537 516.342
R193 VSS.n9014 VSS.n1563 516.342
R194 VSS.n9345 VSS.n1482 516.342
R195 VSS.n9308 VSS.n1507 516.342
R196 VSS.n9247 VSS.n1515 516.342
R197 VSS.n9181 VSS.n1525 516.342
R198 VSS.t5 VSS.t1077 412.349
R199 VSS.t129 VSS.t842 412.349
R200 VSS.n10848 VSS.t817 407.188
R201 VSS.t763 VSS.n11300 407.188
R202 VSS.n10851 VSS.n249 383.618
R203 VSS.n10852 VSS.n10851 381.962
R204 VSS.n249 VSS.n248 381.132
R205 VSS.n10852 VSS.n248 379.474
R206 VSS.t1594 VSS.t186 362.154
R207 VSS.t191 VSS.t1821 358.87
R208 VSS.t409 VSS.t856 303.373
R209 VSS.t410 VSS.t905 303.373
R210 VSS.t896 VSS.t333 303.373
R211 VSS.t335 VSS.t1466 303.373
R212 VSS.t329 VSS.t944 303.373
R213 VSS.t757 VSS.t331 303.373
R214 VSS.t772 VSS.t352 303.373
R215 VSS.t353 VSS.t1360 303.269
R216 VSS.t891 VSS.t455 303.269
R217 VSS.t454 VSS.t571 303.269
R218 VSS.t814 VSS.t285 303.269
R219 VSS.t287 VSS.t721 303.269
R220 VSS.t1111 VSS.t998 300.337
R221 VSS.t464 VSS.t392 300.337
R222 VSS.t394 VSS.t877 300.337
R223 VSS.t308 VSS.t808 300.337
R224 VSS.t310 VSS.t690 300.337
R225 VSS.t292 VSS.t1294 300.236
R226 VSS.t704 VSS.t293 300.236
R227 VSS.t644 VSS.t0 300.236
R228 VSS.t182 VSS.t501 300.236
R229 VSS.t171 VSS.t487 300.236
R230 VSS.t163 VSS.t760 300.236
R231 VSS.t396 VSS.t811 296.584
R232 VSS.n10858 VSS.n243 267.474
R233 VSS.n10862 VSS.n243 266.829
R234 VSS.n10858 VSS.n242 266.276
R235 VSS.n10862 VSS.n242 265.632
R236 VSS.t45 VSS.t5 262.702
R237 VSS.t41 VSS.t129 262.702
R238 VSS.t317 VSS.t853 256.925
R239 VSS.t740 VSS.t422 256.925
R240 VSS.t423 VSS.t604 256.925
R241 VSS.n9302 VSS.t1385 248.619
R242 VSS.n1564 VSS.n132 244.691
R243 VSS.n10287 VSS.n10286 242.161
R244 VSS.n10861 VSS.t1594 219.544
R245 VSS.t1821 VSS.n10859 219.544
R246 VSS.t1077 VSS.n245 219.544
R247 VSS.t842 VSS.n10849 219.544
R248 VSS.n10697 VSS.n10696 215.996
R249 VSS.t856 VSS.t612 206.678
R250 VSS.t413 VSS.t409 206.678
R251 VSS.t411 VSS.t410 206.678
R252 VSS.t905 VSS.t1256 206.678
R253 VSS.t976 VSS.t896 206.678
R254 VSS.t333 VSS.t334 206.678
R255 VSS.t336 VSS.t335 206.678
R256 VSS.t1466 VSS.t618 206.678
R257 VSS.t944 VSS.t979 206.678
R258 VSS.t330 VSS.t329 206.678
R259 VSS.t331 VSS.t332 206.678
R260 VSS.t937 VSS.t757 206.678
R261 VSS.t1537 VSS.t772 206.678
R262 VSS.t357 VSS.t353 206.607
R263 VSS.t1360 VSS.t545 206.607
R264 VSS.t534 VSS.t891 206.607
R265 VSS.t455 VSS.t452 206.607
R266 VSS.t453 VSS.t454 206.607
R267 VSS.t571 VSS.t1315 206.607
R268 VSS.t1034 VSS.t814 206.607
R269 VSS.t285 VSS.t286 206.607
R270 VSS.t288 VSS.t287 206.607
R271 VSS.t721 VSS.t647 206.607
R272 VSS.t668 VSS.t884 206.607
R273 VSS.t352 VSS.t354 205.131
R274 VSS.t1303 VSS.t396 204.609
R275 VSS.t998 VSS.t1037 204.609
R276 VSS.t676 VSS.t1111 204.609
R277 VSS.t859 VSS.t464 204.609
R278 VSS.t392 VSS.t395 204.609
R279 VSS.t393 VSS.t394 204.609
R280 VSS.t877 VSS.t1126 204.609
R281 VSS.t808 VSS.t837 204.609
R282 VSS.t309 VSS.t308 204.609
R283 VSS.t311 VSS.t310 204.609
R284 VSS.t690 VSS.t947 204.609
R285 VSS.t1385 VSS.t1426 204.609
R286 VSS.t1294 VSS.t1025 204.541
R287 VSS.t297 VSS.t292 204.541
R288 VSS.t293 VSS.t294 204.541
R289 VSS.t684 VSS.t704 204.541
R290 VSS.t775 VSS.t644 204.541
R291 VSS.t0 VSS.t147 204.541
R292 VSS.t153 VSS.t182 204.541
R293 VSS.t501 VSS.t459 204.541
R294 VSS.t487 VSS.t1306 204.541
R295 VSS.t172 VSS.t171 204.541
R296 VSS.t162 VSS.t163 204.541
R297 VSS.t760 VSS.t792 204.541
R298 VSS.t811 VSS.t550 204.541
R299 VSS.n10850 VSS.t41 194.681
R300 VSS.n10850 VSS.t45 186.238
R301 VSS.t318 VSS.t319 175.035
R302 VSS.t323 VSS.t317 175.035
R303 VSS.t853 VSS.t641 175.035
R304 VSS.t748 VSS.t740 175.035
R305 VSS.t422 VSS.t421 175.035
R306 VSS.t424 VSS.t423 175.035
R307 VSS.t604 VSS.t1287 175.035
R308 VSS.t612 VSS.n1564 172.355
R309 VSS.t1256 VSS.n9012 172.355
R310 VSS.n9011 VSS.t976 172.355
R311 VSS.t618 VSS.n1533 172.355
R312 VSS.t979 VSS.n9112 172.355
R313 VSS.n9116 VSS.t937 172.355
R314 VSS.n9115 VSS.t1537 172.355
R315 VSS.t545 VSS.n9179 172.296
R316 VSS.n9178 VSS.t534 172.296
R317 VSS.t1315 VSS.n1517 172.296
R318 VSS.n1516 VSS.t1034 172.296
R319 VSS.t647 VSS.n9306 172.296
R320 VSS.n9305 VSS.t668 172.296
R321 VSS.n353 VSS.t676 170.631
R322 VSS.n10186 VSS.t859 170.631
R323 VSS.t1126 VSS.n10183 170.631
R324 VSS.t837 VSS.n354 170.631
R325 VSS.t947 VSS.n10177 170.631
R326 VSS.n10176 VSS.t1426 170.631
R327 VSS.n10286 VSS.t1025 170.572
R328 VSS.n281 VSS.t684 170.572
R329 VSS.n10246 VSS.t775 170.572
R330 VSS.t459 VSS.n10243 170.572
R331 VSS.t1306 VSS.n282 170.572
R332 VSS.t792 VSS.n10237 170.572
R333 VSS.n10236 VSS.t550 170.572
R334 VSS.t21 VSS.t596 163.815
R335 VSS.t29 VSS.t1104 163.815
R336 VSS.t12 VSS.t39 159.155
R337 VSS.t10 VSS.t145 159.155
R338 VSS.t884 VSS.n9304 158.827
R339 VSS.n9010 VSS.t413 148.365
R340 VSS.n9092 VSS.t334 148.365
R341 VSS.n9113 VSS.t330 148.365
R342 VSS.n9177 VSS.t354 148.315
R343 VSS.n9249 VSS.t452 148.315
R344 VSS.n9299 VSS.t286 148.315
R345 VSS.n351 VSS.t1303 146.881
R346 VSS.t395 VSS.n10185 146.881
R347 VSS.n392 VSS.t309 146.881
R348 VSS.n279 VSS.t297 146.832
R349 VSS.t147 VSS.n10245 146.832
R350 VSS.n320 VSS.t172 146.832
R351 VSS.t641 VSS.n423 145.966
R352 VSS.n10126 VSS.t748 145.966
R353 VSS.t1287 VSS.n10123 145.966
R354 VSS.t3 VSS.t1615 145.738
R355 VSS.t699 VSS.t195 145.738
R356 VSS.n9013 VSS.t411 144.674
R357 VSS.n9091 VSS.t336 144.674
R358 VSS.t332 VSS.n9114 144.674
R359 VSS.n9180 VSS.t357 144.625
R360 VSS.n9248 VSS.t453 144.625
R361 VSS.n9307 VSS.t288 144.625
R362 VSS.t1037 VSS.n352 143.227
R363 VSS.n10184 VSS.t393 143.227
R364 VSS.n10178 VSS.t311 143.227
R365 VSS.t294 VSS.n280 143.179
R366 VSS.n10244 VSS.t153 143.179
R367 VSS.n10238 VSS.t162 143.179
R368 VSS.t192 VSS.t33 142.941
R369 VSS.t193 VSS.t31 142.941
R370 VSS.n10860 VSS.t191 134.636
R371 VSS.n10847 VSS.n10846 132.153
R372 VSS.t186 VSS.n10860 128.067
R373 VSS.t319 VSS.n9301 125.65
R374 VSS.t421 VSS.n10125 125.65
R375 VSS.n9300 VSS.t323 122.525
R376 VSS.n10124 VSS.t424 122.525
R377 VSS.n1391 VSS.n424 122.525
R378 VSS.n9116 VSS.n9115 116.626
R379 VSS.n9306 VSS.n9305 116.585
R380 VSS.n10177 VSS.n10176 115.459
R381 VSS.n10237 VSS.n10236 115.419
R382 VSS.t379 VSS.t475 106.296
R383 VSS.t522 VSS.t156 106.296
R384 VSS.t1 VSS.t21 104.365
R385 VSS.t39 VSS.t1 104.365
R386 VSS.t37 VSS.t12 104.365
R387 VSS.t145 VSS.t7 104.365
R388 VSS.t7 VSS.t29 104.365
R389 VSS.n10662 VSS.t10 100.638
R390 VSS.t183 VSS.t14 88.1506
R391 VSS.t185 VSS.t18 88.1506
R392 VSS.n10696 VSS.t596 87.2188
R393 VSS.t1104 VSS.n244 87.2188
R394 VSS.t25 VSS.t165 86.287
R395 VSS.t137 VSS.t196 86.287
R396 VSS.t525 VSS.t27 83.4915
R397 VSS.n10600 VSS.t509 82.3733
R398 VSS.n9012 VSS.n9011 81.5642
R399 VSS.n9179 VSS.n9178 81.5364
R400 VSS.n10186 VSS.n353 80.7481
R401 VSS.n10246 VSS.n281 80.7209
R402 VSS.n10847 VSS.t349 75.9965
R403 VSS.t16 VSS.n10599 73.8006
R404 VSS.n10602 VSS.t190 73.8006
R405 VSS.t384 VSS.t379 72.4152
R406 VSS.n9465 VSS.t155 72.4152
R407 VSS.t1222 VSS.t522 72.4152
R408 VSS.t430 VSS.t1431 69.1825
R409 VSS.n10126 VSS.n423 69.0763
R410 VSS.n10859 VSS.n245 67.5525
R411 VSS.t553 VSS.t150 65.5106
R412 VSS.t380 VSS.n9303 63.4927
R413 VSS.t261 VSS.t337 63.4385
R414 VSS.t653 VSS.n1499 60.3892
R415 VSS.t284 VSS.t107 59.6927
R416 VSS.n1498 VSS.t1794 56.1219
R417 VSS.t397 VSS.t217 53.3171
R418 VSS.n9112 VSS.n1533 53.1461
R419 VSS.n1517 VSS.n1516 53.128
R420 VSS.n10183 VSS.n354 52.6143
R421 VSS.n10243 VSS.n282 52.5966
R422 VSS.n9347 VSS.t381 51.9839
R423 VSS.t154 VSS.n9422 51.9839
R424 VSS.n1394 VSS.t484 51.9839
R425 VSS.t264 VSS.t498 51.3247
R426 VSS.t157 VSS.n1383 50.6908
R427 VSS.t568 VSS.t105 47.579
R428 VSS.n10123 VSS.n424 45.0092
R429 VSS.n9346 VSS.t1244 44.8718
R430 VSS.t588 VSS.t528 44.6302
R431 VSS.t868 VSS.t609 44.6302
R432 VSS.t339 VSS.t340 44.6302
R433 VSS.t102 VSS.t103 44.6302
R434 VSS.t558 VSS.t1253 44.6302
R435 VSS.t681 VSS.t908 44.6302
R436 VSS.t98 VSS.t96 44.6302
R437 VSS.t281 VSS.t282 44.6302
R438 VSS.t834 VSS.t553 44.6302
R439 VSS.t156 VSS.t429 43.8373
R440 VSS.t255 VSS.t478 42.5581
R441 VSS.t745 VSS.t289 42.0799
R442 VSS.t475 VSS.t2036 41.639
R443 VSS.n1393 VSS.n1392 41.639
R444 VSS.t561 VSS.t160 40.8845
R445 VSS.t101 VSS.t168 40.486
R446 VSS.t256 VSS.t376 39.2906
R447 VSS.t490 VSS.t108 38.8124
R448 VSS.t433 VSS.t154 38.1476
R449 VSS.t506 VSS.n9524 37.2982
R450 VSS.t540 VSS.n1182 37.2982
R451 VSS.n9561 VSS.t576 37.2185
R452 VSS.n1183 VSS.t671 37.2185
R453 VSS.n565 VSS.t1064 37.2185
R454 VSS.t795 VSS.n11288 37.2185
R455 VSS.n11298 VSS.t834 37.2185
R456 VSS.t100 VSS.t591 36.3418
R457 VSS.t106 VSS.t495 36.3418
R458 VSS.t1157 VSS.t467 35.4652
R459 VSS.t638 VSS.t213 35.1464
R460 VSS.n1390 VSS.t378 34.7479
R461 VSS.t265 VSS.t687 34.5885
R462 VSS.t260 VSS.t1157 34.5885
R463 VSS.t263 VSS.t638 34.5088
R464 VSS.t283 VSS.t472 34.2697
R465 VSS.n9465 VSS.t1431 33.8803
R466 VSS.n4805 VSS.n4804 33.7899
R467 VSS.t495 VSS.t56 33.3134
R468 VSS.t399 VSS.n833 32.0383
R469 VSS.t148 VSS.n6 32.0383
R470 VSS.n10118 VSS.t377 31.2413
R471 VSS.n10067 VSS.t304 31.2413
R472 VSS.n11152 VSS.t166 31.2413
R473 VSS.t528 VSS.n1390 30.7631
R474 VSS.t259 VSS.t306 30.4443
R475 VSS.t376 VSS.t215 30.3646
R476 VSS.t467 VSS.t307 30.0459
R477 VSS.t168 VSS.t730 29.5677
R478 VSS.n10599 VSS.n10442 29.446
R479 VSS.t160 VSS.t100 29.1692
R480 VSS.n1499 VSS.n1498 28.5785
R481 VSS.t401 VSS.t257 28.2926
R482 VSS.t289 VSS.t258 27.9738
R483 VSS.n10602 VSS.n10601 26.8369
R484 VSS.t155 VSS.t2475 26.7681
R485 VSS.t149 VSS.t99 26.6986
R486 VSS.n11299 VSS.n11298 26.4596
R487 VSS.n9889 VSS.t305 25.9017
R488 VSS.t398 VSS.t601 25.5032
R489 VSS.n9526 VSS.n9525 25.1844
R490 VSS.t1064 VSS.t97 25.025
R491 VSS.t531 VSS.t101 25.025
R492 VSS.t312 VSS.t653 23.2767
R493 VSS.n9766 VSS.t229 23.1123
R494 VSS.n11279 VSS.t54 23.1123
R495 VSS.t733 VSS.t68 22.5544
R496 VSS.t150 VSS.n11297 22.4748
R497 VSS.t158 VSS.n208 22.2357
R498 VSS.n11297 VSS.t151 22.156
R499 VSS.t68 VSS.t568 22.0763
R500 VSS.n9302 VSS.t318 21.8797
R501 VSS.t215 VSS.n10117 21.5184
R502 VSS.t220 VSS.n10066 21.5184
R503 VSS.n10032 VSS.t65 21.5184
R504 VSS.n11292 VSS.t63 21.5184
R505 VSS.n10929 VSS.n217 21.2793
R506 VSS.t1237 VSS.t157 21.0784
R507 VSS.t509 VSS.t192 20.8733
R508 VSS.t31 VSS.t525 20.8733
R509 VSS.t585 VSS.n506 20.6417
R510 VSS.t266 VSS.t868 20.4824
R511 VSS.t97 VSS.t531 19.6057
R512 VSS.t340 VSS.t713 19.2072
R513 VSS.t601 VSS.t399 19.1275
R514 VSS.n1184 VSS.t224 18.8884
R515 VSS.n1394 VSS.n1393 18.6214
R516 VSS.n9013 VSS.n9010 18.4538
R517 VSS.n9092 VSS.n9091 18.4538
R518 VSS.n9114 VSS.n9113 18.4538
R519 VSS.n9180 VSS.n9177 18.4475
R520 VSS.n9249 VSS.n9248 18.4475
R521 VSS.n9307 VSS.n9299 18.4475
R522 VSS.t498 VSS.t220 18.3306
R523 VSS.t224 VSS.t537 18.3306
R524 VSS.n352 VSS.n351 18.2692
R525 VSS.n10185 VSS.n10184 18.2692
R526 VSS.n10178 VSS.n392 18.2692
R527 VSS.n280 VSS.n279 18.263
R528 VSS.n10245 VSS.n10244 18.263
R529 VSS.n10238 VSS.n320 18.263
R530 VSS.t165 VSS.t3 18.0778
R531 VSS.t196 VSS.t25 18.0778
R532 VSS.t195 VSS.t137 18.0778
R533 VSS.t105 VSS.t149 17.9321
R534 VSS.t99 VSS.t148 17.9321
R535 VSS.n566 VSS.t60 17.7727
R536 VSS.n9561 VSS.n9560 17.6133
R537 VSS.n11279 VSS.n148 17.6133
R538 VSS.n9525 VSS.t266 16.7366
R539 VSS.n11286 VSS.n93 16.7366
R540 VSS.n11361 VSS.t716 16.5773
R541 VSS.t262 VSS.t401 16.3382
R542 VSS.t257 VSS.t397 16.3382
R543 VSS.t33 VSS.t183 16.2142
R544 VSS.t14 VSS.t185 16.2142
R545 VSS.t18 VSS.t193 16.2142
R546 VSS.n11468 VSS.t481 16.0991
R547 VSS.n9301 VSS.n9300 15.6285
R548 VSS.n10125 VSS.n10124 15.6285
R549 VSS.t282 VSS.t716 15.4615
R550 VSS.n11287 VSS.t63 15.1427
R551 VSS.t151 VSS.t481 15.1427
R552 VSS.t730 VSS.t158 15.063
R553 VSS.n9564 VSS.t262 14.9036
R554 VSS.n4803 VSS.n1580 14.678
R555 VSS.n8954 VSS.n8953 14.6753
R556 VSS.t1253 VSS.t102 14.6646
R557 VSS.t304 VSS.t259 14.1864
R558 VSS.t306 VSS.t264 14.1864
R559 VSS.t54 VSS.t681 14.1067
R560 VSS.n10117 VSS.t650 13.6285
R561 VSS.t1615 VSS.t16 13.4187
R562 VSS.t190 VSS.t699 13.4187
R563 VSS.t217 VSS.t615 12.194
R564 VSS.t576 VSS.t229 12.194
R565 VSS.t713 VSS.n218 12.0346
R566 VSS.n9523 VSS.t398 11.7955
R567 VSS.n9524 VSS.n9523 11.4767
R568 VSS.n9890 VSS.n9889 11.4767
R569 VSS.n1184 VSS.n1183 11.4767
R570 VSS.n11289 VSS.n11286 11.4767
R571 VSS.n11288 VSS.n11287 11.4767
R572 VSS.t305 VSS.t585 11.397
R573 VSS.t908 VSS.t98 10.9188
R574 VSS.t338 VSS.n217 10.7595
R575 VSS.n8952 VSS.n1580 10.4817
R576 VSS.t65 VSS.t558 10.361
R577 VSS.t472 VSS.t284 10.361
R578 VSS.t687 VSS.t260 10.0422
R579 VSS.t96 VSS.t281 9.96249
R580 VSS.n10982 VSS.n208 9.8031
R581 VSS.t213 VSS.t650 9.48432
R582 VSS.n1353 VSS.t268 9.37419
R583 VSS.n9766 VSS.t615 9.32492
R584 VSS.n9143 VSS.n9142 9.30555
R585 VSS.n1491 VSS.n1490 9.30555
R586 VSS.n1211 VSS.n1210 9.30555
R587 VSS.n10949 VSS.n10948 9.30555
R588 VSS.n10995 VSS.n10994 9.30555
R589 VSS.n8976 VSS.n8975 9.30555
R590 VSS.n981 VSS.n980 9.30555
R591 VSS.n1039 VSS.n1038 9.30555
R592 VSS.n1088 VSS.n1087 9.30555
R593 VSS.n874 VSS.n873 9.30555
R594 VSS.n576 VSS.t104 9.29148
R595 VSS.n9304 VSS.t380 9.05234
R596 VSS.n1392 VSS.n1391 9.05234
R597 VSS.n9303 VSS.t381 8.92303
R598 VSS.n11309 VSS.n128 8.8165
R599 VSS.n10837 VSS.t3113 8.52542
R600 VSS.n10791 VSS.t3537 8.52542
R601 VSS.n10809 VSS.t841 8.52542
R602 VSS.n10828 VSS.t2769 8.52542
R603 VSS.n10773 VSS.t1461 8.52542
R604 VSS.n10855 VSS.t1893 8.52542
R605 VSS.n10742 VSS.t2290 8.52542
R606 VSS.n10746 VSS.t1076 8.52542
R607 VSS.n10813 VSS.t3203 8.52542
R608 VSS.n10815 VSS.t1907 8.52542
R609 VSS.n10749 VSS.t888 8.52542
R610 VSS.n10747 VSS.t580 8.52542
R611 VSS.n10736 VSS.t3543 8.52542
R612 VSS.n10784 VSS.t2232 8.52542
R613 VSS.n10737 VSS.t1262 8.52542
R614 VSS.n10778 VSS.t961 8.52542
R615 VSS.t484 VSS.t1222 8.40578
R616 VSS.t591 VSS.t106 8.28888
R617 VSS.n4803 VSS.n60 8.20625
R618 VSS.n9202 VSS.t626 8.06917
R619 VSS.n9184 VSS.t2725 8.06917
R620 VSS.n9058 VSS.t3303 8.06917
R621 VSS.n9057 VSS.t2274 8.06917
R622 VSS.n9054 VSS.t2895 8.06917
R623 VSS.n9054 VSS.t3577 8.06917
R624 VSS.n9051 VSS.t2074 8.06917
R625 VSS.n9051 VSS.t2805 8.06917
R626 VSS.n9050 VSS.t2386 8.06917
R627 VSS.n9050 VSS.t3129 8.06917
R628 VSS.n9122 VSS.t1224 8.06917
R629 VSS.n9122 VSS.t1937 8.06917
R630 VSS.n9123 VSS.t771 8.06917
R631 VSS.n9123 VSS.t1536 8.06917
R632 VSS.n9127 VSS.t2192 8.06917
R633 VSS.n9127 VSS.t2899 8.06917
R634 VSS.n9054 VSS.t1783 8.06917
R635 VSS.n9054 VSS.t1625 8.06917
R636 VSS.n9051 VSS.t936 8.06917
R637 VSS.n9051 VSS.t756 8.06917
R638 VSS.n9050 VSS.t1291 8.06917
R639 VSS.n9050 VSS.t1095 8.06917
R640 VSS.n9122 VSS.t3185 8.06917
R641 VSS.n9122 VSS.t3039 8.06917
R642 VSS.n9123 VSS.t2799 8.06917
R643 VSS.n9123 VSS.t2607 8.06917
R644 VSS.n9127 VSS.t1041 8.06917
R645 VSS.n9127 VSS.t865 8.06917
R646 VSS.n1543 VSS.t3509 8.06917
R647 VSS.n1542 VSS.t1510 8.06917
R648 VSS.n1549 VSS.t1773 8.06917
R649 VSS.n1541 VSS.t1014 8.06917
R650 VSS.n9171 VSS.t3101 8.06917
R651 VSS.n9137 VSS.t2015 8.06917
R652 VSS.n1526 VSS.t2633 8.06917
R653 VSS.n9133 VSS.t1604 8.06917
R654 VSS.n1512 VSS.t861 8.06917
R655 VSS.n9253 VSS.t2941 8.06917
R656 VSS.n9139 VSS.t1711 8.06917
R657 VSS.n9138 VSS.t2396 8.06917
R658 VSS.n9237 VSS.t2929 8.06917
R659 VSS.n9237 VSS.t1869 8.06917
R660 VSS.n9234 VSS.t2122 8.06917
R661 VSS.n9234 VSS.t1033 8.06917
R662 VSS.n9233 VSS.t2428 8.06917
R663 VSS.n9233 VSS.t1409 8.06917
R664 VSS.n9227 VSS.t1258 8.06917
R665 VSS.n9227 VSS.t3269 8.06917
R666 VSS.n9226 VSS.t813 8.06917
R667 VSS.n9226 VSS.t2891 8.06917
R668 VSS.n9223 VSS.t2212 8.06917
R669 VSS.n9223 VSS.t1146 8.06917
R670 VSS.n9237 VSS.t3333 8.06917
R671 VSS.n9237 VSS.t1366 8.06917
R672 VSS.n9234 VSS.t2563 8.06917
R673 VSS.n9234 VSS.t3629 8.06917
R674 VSS.n9233 VSS.t2907 8.06917
R675 VSS.n9233 VSS.t831 8.06917
R676 VSS.n9227 VSS.t1719 8.06917
R677 VSS.n9227 VSS.t2775 8.06917
R678 VSS.n9226 VSS.t1314 8.06917
R679 VSS.n9226 VSS.t2346 8.06917
R680 VSS.n9223 VSS.t2675 8.06917
R681 VSS.n9223 VSS.t570 8.06917
R682 VSS.n9242 VSS.t1617 8.06917
R683 VSS.n9212 VSS.t3619 8.06917
R684 VSS.n1518 VSS.t2384 8.06917
R685 VSS.n9208 VSS.t3125 8.06917
R686 VSS.n1504 VSS.t2040 8.06917
R687 VSS.n9311 VSS.t967 8.06917
R688 VSS.n9214 VSS.t1629 8.06917
R689 VSS.n9213 VSS.t2312 8.06917
R690 VSS.n9269 VSS.t2561 8.06917
R691 VSS.n9269 VSS.t1534 8.06917
R692 VSS.n9273 VSS.t1791 8.06917
R693 VSS.n9273 VSS.t667 8.06917
R694 VSS.n9274 VSS.t2100 8.06917
R695 VSS.n9274 VSS.t1004 8.06917
R696 VSS.n9282 VSS.t883 8.06917
R697 VSS.n9282 VSS.t2953 8.06917
R698 VSS.n9283 VSS.t3575 8.06917
R699 VSS.n9283 VSS.t2525 8.06917
R700 VSS.n9287 VSS.t1877 8.06917
R701 VSS.n9287 VSS.t779 8.06917
R702 VSS.n9269 VSS.t2797 8.06917
R703 VSS.n9269 VSS.t720 8.06917
R704 VSS.n9273 VSS.t1985 8.06917
R705 VSS.n9273 VSS.t3063 8.06917
R706 VSS.n9274 VSS.t2292 8.06917
R707 VSS.n9274 VSS.t3321 8.06917
R708 VSS.n9282 VSS.t1091 8.06917
R709 VSS.n9282 VSS.t2188 8.06917
R710 VSS.n9283 VSS.t646 8.06917
R711 VSS.n9283 VSS.t1785 8.06917
R712 VSS.n9287 VSS.t2068 8.06917
R713 VSS.n9287 VSS.t3143 8.06917
R714 VSS.n9293 VSS.t1368 8.06917
R715 VSS.n9263 VSS.t3343 8.06917
R716 VSS.n1508 VSS.t879 8.06917
R717 VSS.n9259 VSS.t1633 8.06917
R718 VSS.n1495 VSS.t2851 8.06917
R719 VSS.n9351 VSS.t2136 8.06917
R720 VSS.n9265 VSS.t1376 8.06917
R721 VSS.n9264 VSS.t2400 8.06917
R722 VSS.n9372 VSS.t3453 8.06917
R723 VSS.n9372 VSS.t2773 8.06917
R724 VSS.n9369 VSS.t2679 8.06917
R725 VSS.n9369 VSS.t1969 8.06917
R726 VSS.n9368 VSS.t3015 8.06917
R727 VSS.n9368 VSS.t2276 8.06917
R728 VSS.n9362 VSS.t1823 8.06917
R729 VSS.n9362 VSS.t1083 8.06917
R730 VSS.n9361 VSS.t1430 8.06917
R731 VSS.n9361 VSS.t632 8.06917
R732 VSS.n9358 VSS.t2781 8.06917
R733 VSS.n9358 VSS.t2058 8.06917
R734 VSS.n9372 VSS.t1177 8.06917
R735 VSS.n9372 VSS.t2246 8.06917
R736 VSS.n9369 VSS.t3457 8.06917
R737 VSS.n9369 VSS.t1480 8.06917
R738 VSS.n9368 VSS.t652 8.06917
R739 VSS.n9368 VSS.t1787 8.06917
R740 VSS.n9362 VSS.t2603 8.06917
R741 VSS.n9362 VSS.t474 8.06917
R742 VSS.n9361 VSS.t2208 8.06917
R743 VSS.n9361 VSS.t3249 8.06917
R744 VSS.n9358 VSS.t3561 8.06917
R745 VSS.n9358 VSS.t1567 8.06917
R746 VSS.n9340 VSS.t3533 8.06917
R747 VSS.n9321 VSS.t2847 8.06917
R748 VSS.n1500 VSS.t2048 8.06917
R749 VSS.n9317 VSS.t3131 8.06917
R750 VSS.n1476 VSS.t2597 8.06917
R751 VSS.n9384 VSS.t469 8.06917
R752 VSS.n1477 VSS.t2180 8.06917
R753 VSS.n9377 VSS.t3213 8.06917
R754 VSS.n9392 VSS.t2689 8.06917
R755 VSS.n9392 VSS.t587 8.06917
R756 VSS.n9396 VSS.t1883 8.06917
R757 VSS.n9396 VSS.t2951 8.06917
R758 VSS.n9397 VSS.t2206 8.06917
R759 VSS.n9397 VSS.t3245 8.06917
R760 VSS.n9405 VSS.t983 8.06917
R761 VSS.n9405 VSS.t2064 8.06917
R762 VSS.n9406 VSS.t527 8.06917
R763 VSS.n9406 VSS.t1685 8.06917
R764 VSS.n9410 VSS.t1977 8.06917
R765 VSS.n9410 VSS.t3059 8.06917
R766 VSS.n9392 VSS.t2011 8.06917
R767 VSS.n9392 VSS.t1325 8.06917
R768 VSS.n9396 VSS.t1221 8.06917
R769 VSS.n9396 VSS.t3583 8.06917
R770 VSS.n9397 VSS.t1561 8.06917
R771 VSS.n9397 VSS.t799 8.06917
R772 VSS.n9405 VSS.t3407 8.06917
R773 VSS.n9405 VSS.t2729 8.06917
R774 VSS.n9406 VSS.t3051 8.06917
R775 VSS.n9406 VSS.t2316 8.06917
R776 VSS.n9410 VSS.t1329 8.06917
R777 VSS.n9410 VSS.t521 8.06917
R778 VSS.n9416 VSS.t1909 8.06917
R779 VSS.n1397 VSS.t2981 8.06917
R780 VSS.n1487 VSS.t1488 8.06917
R781 VSS.n1486 VSS.t2511 8.06917
R782 VSS.n1220 VSS.t1089 8.06917
R783 VSS.n9531 VSS.t2178 8.06917
R784 VSS.n1399 VSS.t1415 8.06917
R785 VSS.n1398 VSS.t620 8.06917
R786 VSS.n1435 VSS.t1551 8.06917
R787 VSS.n1435 VSS.t2577 8.06917
R788 VSS.n1434 VSS.t1865 8.06917
R789 VSS.n1434 VSS.t2937 8.06917
R790 VSS.n1229 VSS.t608 8.06917
R791 VSS.n1229 VSS.t1749 8.06917
R792 VSS.n1228 VSS.t3313 8.06917
R793 VSS.n1228 VSS.t1335 8.06917
R794 VSS.n1225 VSS.t1653 8.06917
R795 VSS.n1225 VSS.t2709 8.06917
R796 VSS.n1435 VSS.t3501 8.06917
R797 VSS.n1435 VSS.t2817 8.06917
R798 VSS.n1434 VSS.t708 8.06917
R799 VSS.n1434 VSS.t3135 8.06917
R800 VSS.n1229 VSS.t2643 8.06917
R801 VSS.n1229 VSS.t1941 8.06917
R802 VSS.n1228 VSS.t2234 8.06917
R803 VSS.n1228 VSS.t1541 8.06917
R804 VSS.n1225 VSS.t3593 8.06917
R805 VSS.n1225 VSS.t2909 8.06917
R806 VSS.n11235 VSS.t3201 8.06917
R807 VSS.n11233 VSS.t801 8.06917
R808 VSS.n11229 VSS.t1455 8.06917
R809 VSS.n11224 VSS.t3437 8.06917
R810 VSS.n11202 VSS.t1897 8.06917
R811 VSS.n11200 VSS.t2963 8.06917
R812 VSS.n11257 VSS.t3189 8.06917
R813 VSS.n11196 VSS.t2148 8.06917
R814 VSS.n11181 VSS.t2763 8.06917
R815 VSS.n11179 VSS.t3447 8.06917
R816 VSS.n11175 VSS.t3307 8.06917
R817 VSS.n11173 VSS.t939 8.06917
R818 VSS.n153 VSS.t3047 8.06917
R819 VSS.n11164 VSS.t590 8.06917
R820 VSS.n177 VSS.t2288 8.06917
R821 VSS.n11156 VSS.t1250 8.06917
R822 VSS.n735 VSS.t1867 8.06917
R823 VSS.n731 VSS.t767 8.06917
R824 VSS.n729 VSS.t2104 8.06917
R825 VSS.n746 VSS.t3157 8.06917
R826 VSS.n705 VSS.t1351 8.06917
R827 VSS.n703 VSS.t2033 8.06917
R828 VSS.n699 VSS.t3595 8.06917
R829 VSS.n695 VSS.t1606 8.06917
R830 VSS.n692 VSS.t1861 8.06917
R831 VSS.n9835 VSS.t1123 8.06917
R832 VSS.n9830 VSS.t515 8.06917
R833 VSS.n9824 VSS.t1679 8.06917
R834 VSS.n9818 VSS.t2132 8.06917
R835 VSS.n9811 VSS.t1053 8.06917
R836 VSS.n9807 VSS.t2358 8.06917
R837 VSS.n9801 VSS.t3381 8.06917
R838 VSS.n9797 VSS.t3017 8.06917
R839 VSS.n788 VSS.t1943 8.06917
R840 VSS.n789 VSS.t3225 8.06917
R841 VSS.n9784 VSS.t1209 8.06917
R842 VSS.n9775 VSS.t2721 8.06917
R843 VSS.n9769 VSS.t2001 8.06917
R844 VSS.n9587 VSS.t2260 8.06917
R845 VSS.n9567 VSS.t1502 8.06917
R846 VSS.n830 VSS.t1769 8.06917
R847 VSS.n9600 VSS.t1006 8.06917
R848 VSS.n1442 VSS.t2322 8.06917
R849 VSS.n1440 VSS.t3357 8.06917
R850 VSS.n1453 VSS.t1226 8.06917
R851 VSS.n1455 VSS.t3587 8.06917
R852 VSS.n1424 VSS.t1812 8.06917
R853 VSS.n1467 VSS.t2879 8.06917
R854 VSS.n1471 VSS.t2090 8.06917
R855 VSS.n1417 VSS.t1411 8.06917
R856 VSS.n1154 VSS.t2420 8.06917
R857 VSS.n1154 VSS.t3483 8.06917
R858 VSS.n1155 VSS.t2761 8.06917
R859 VSS.n1155 VSS.t686 8.06917
R860 VSS.n9555 VSS.t1596 8.06917
R861 VSS.n9555 VSS.t2621 8.06917
R862 VSS.n9554 VSS.t1156 8.06917
R863 VSS.n9554 VSS.t2218 8.06917
R864 VSS.n9551 VSS.t2529 8.06917
R865 VSS.n9551 VSS.t3579 8.06917
R866 VSS.n1154 VSS.t1929 8.06917
R867 VSS.n1154 VSS.t1213 8.06917
R868 VSS.n1155 VSS.t2236 8.06917
R869 VSS.n1155 VSS.t1545 8.06917
R870 VSS.n9555 VSS.t1031 8.06917
R871 VSS.n9555 VSS.t3395 8.06917
R872 VSS.n9554 VSS.t575 8.06917
R873 VSS.n9554 VSS.t3043 8.06917
R874 VSS.n9551 VSS.t2009 8.06917
R875 VSS.n9551 VSS.t1321 8.06917
R876 VSS.n1215 VSS.t1571 8.06917
R877 VSS.n9544 VSS.t737 8.06917
R878 VSS.n1216 VSS.t1016 8.06917
R879 VSS.n9537 VSS.t3385 8.06917
R880 VSS.n1201 VSS.t1681 8.06917
R881 VSS.n1163 VSS.t2727 8.06917
R882 VSS.n1207 VSS.t2286 8.06917
R883 VSS.n1162 VSS.t1246 8.06917
R884 VSS.n213 VSS.t2927 8.06917
R885 VSS.n10933 VSS.t846 8.06917
R886 VSS.n1165 VSS.t1134 8.06917
R887 VSS.n1164 VSS.t3525 8.06917
R888 VSS.n10976 VSS.t1621 8.06917
R889 VSS.n10943 VSS.t3623 8.06917
R890 VSS.n209 VSS.t1144 8.06917
R891 VSS.n10939 VSS.t3177 8.06917
R892 VSS.n89 VSS.t2472 8.06917
R893 VSS.n11365 VSS.t1463 8.06917
R894 VSS.n10945 VSS.t2050 8.06917
R895 VSS.n10944 VSS.t2777 8.06917
R896 VSS.n84 VSS.t2967 8.06917
R897 VSS.n11378 VSS.t1901 8.06917
R898 VSS.n85 VSS.t2493 8.06917
R899 VSS.n11371 VSS.t3209 8.06917
R900 VSS.n66 VSS.t2324 8.06917
R901 VSS.n66 VSS.t3359 8.06917
R902 VSS.n67 VSS.t2657 8.06917
R903 VSS.n67 VSS.t555 8.06917
R904 VSS.n73 VSS.t1498 8.06917
R905 VSS.n73 VSS.t2523 8.06917
R906 VSS.n74 VSS.t1039 8.06917
R907 VSS.n74 VSS.t2128 8.06917
R908 VSS.n77 VSS.t2416 8.06917
R909 VSS.n77 VSS.t3475 8.06917
R910 VSS.t3233 VSS.n11458 8.06917
R911 VSS.n11459 VSS.t3233 8.06917
R912 VSS.t2450 VSS.n11456 8.06917
R913 VSS.n11457 VSS.t2450 8.06917
R914 VSS.t2589 VSS.n11454 8.06917
R915 VSS.n11455 VSS.t2589 8.06917
R916 VSS.t1827 VSS.n11452 8.06917
R917 VSS.n11453 VSS.t1827 8.06917
R918 VSS.n23 VSS.t993 8.06917
R919 VSS.t993 VSS.n18 8.06917
R920 VSS.t1152 VSS.n11442 8.06917
R921 VSS.n11443 VSS.t1152 8.06917
R922 VSS.t3435 VSS.n11440 8.06917
R923 VSS.n11441 VSS.t3435 8.06917
R924 VSS.t2693 VSS.n11438 8.06917
R925 VSS.n11439 VSS.t2693 8.06917
R926 VSS.t2985 VSS.n11436 8.06917
R927 VSS.n11437 VSS.t2985 8.06917
R928 VSS.t914 VSS.n11434 8.06917
R929 VSS.n11435 VSS.t914 8.06917
R930 VSS.t1539 VSS.n11427 8.06917
R931 VSS.n11428 VSS.t1539 8.06917
R932 VSS.t2519 VSS.n11425 8.06917
R933 VSS.n11426 VSS.t2519 8.06917
R934 VSS.t1763 VSS.n11423 8.06917
R935 VSS.n11424 VSS.t1763 8.06917
R936 VSS.t922 VSS.n11421 8.06917
R937 VSS.n11422 VSS.t922 8.06917
R938 VSS.t1072 VSS.n11419 8.06917
R939 VSS.n11420 VSS.t1072 8.06917
R940 VSS.n48 VSS.t3355 8.06917
R941 VSS.t3355 VSS.n43 8.06917
R942 VSS.t2765 VSS.n11409 8.06917
R943 VSS.n11410 VSS.t2765 8.06917
R944 VSS.t1979 VSS.n11407 8.06917
R945 VSS.n11408 VSS.t1979 8.06917
R946 VSS.t1399 VSS.n11405 8.06917
R947 VSS.n11406 VSS.t1399 8.06917
R948 VSS.t480 VSS.n11403 8.06917
R949 VSS.n11404 VSS.t480 8.06917
R950 VSS.t1689 VSS.n11401 8.06917
R951 VSS.n11402 VSS.t1689 8.06917
R952 VSS.n63 VSS.t3141 8.06917
R953 VSS.n63 VSS.t1085 8.06917
R954 VSS.n63 VSS.t461 8.06917
R955 VSS.n63 VSS.t2579 8.06917
R956 VSS.n11324 VSS.t2210 8.06917
R957 VSS.n118 VSS.t1973 8.06917
R958 VSS.n11462 VSS.t1459 8.06917
R959 VSS.n11 VSS.t1492 8.06917
R960 VSS.n11091 VSS.t1713 8.06917
R961 VSS.n11089 VSS.t624 8.06917
R962 VSS.n11084 VSS.t2885 8.06917
R963 VSS.n11079 VSS.t2913 8.06917
R964 VSS.n11058 VSS.t1319 8.06917
R965 VSS.n11056 VSS.t1043 8.06917
R966 VSS.n11113 VSS.t2456 8.06917
R967 VSS.n11052 VSS.t2481 8.06917
R968 VSS.n11034 VSS.t2739 8.06917
R969 VSS.n11032 VSS.t1745 8.06917
R970 VSS.n11028 VSS.t2667 8.06917
R971 VSS.n11025 VSS.t1671 8.06917
R972 VSS.n11132 VSS.t2302 8.06917
R973 VSS.n203 VSS.t1298 8.06917
R974 VSS.n11145 VSS.t1183 8.06917
R975 VSS.n186 VSS.t1234 8.06917
R976 VSS.n10880 VSS.t1484 8.06917
R977 VSS.n10885 VSS.t1512 8.06917
R978 VSS.n10889 VSS.t530 8.06917
R979 VSS.n10873 VSS.t3429 8.06917
R980 VSS.n237 VSS.t1397 8.06917
R981 VSS.n557 VSS.t3405 8.06917
R982 VSS.n553 VSS.t2821 8.06917
R983 VSS.n549 VSS.t2555 8.06917
R984 VSS.n10049 VSS.t2019 8.06917
R985 VSS.n544 VSS.t2849 8.06917
R986 VSS.n540 VSS.t2294 8.06917
R987 VSS.n538 VSS.t2056 8.06917
R988 VSS.n514 VSS.t2753 8.06917
R989 VSS.n529 VSS.t2801 8.06917
R990 VSS.n523 VSS.t1915 8.06917
R991 VSS.n518 VSS.t1683 8.06917
R992 VSS.n500 VSS.t1079 8.06917
R993 VSS.n498 VSS.t1108 8.06917
R994 VSS.n495 VSS.t3301 8.06917
R995 VSS.n10080 VSS.t3111 8.06917
R996 VSS.n489 VSS.t3397 8.06917
R997 VSS.n486 VSS.t1142 8.06917
R998 VSS.n478 VSS.t2547 8.06917
R999 VSS.n459 VSS.t2671 8.06917
R1000 VSS.n10098 VSS.t2134 8.06917
R1001 VSS.n456 VSS.t2949 8.06917
R1002 VSS.n452 VSS.t2046 8.06917
R1003 VSS.n450 VSS.t1829 8.06917
R1004 VSS.n10111 VSS.t2031 8.06917
R1005 VSS.n442 VSS.t2863 8.06917
R1006 VSS.n1301 VSS.t1971 8.06917
R1007 VSS.n1308 VSS.t1747 8.06917
R1008 VSS.n1297 VSS.t3455 8.06917
R1009 VSS.n1317 VSS.t1185 8.06917
R1010 VSS.n11335 VSS.t3159 8.06917
R1011 VSS.n11335 VSS.t2935 8.06917
R1012 VSS.n11333 VSS.t833 8.06917
R1013 VSS.n11333 VSS.t552 8.06917
R1014 VSS.n11332 VSS.t1289 8.06917
R1015 VSS.n11332 VSS.t1018 8.06917
R1016 VSS.n11328 VSS.t1751 8.06917
R1017 VSS.n11328 VSS.t1514 8.06917
R1018 VSS.n11327 VSS.t3567 8.06917
R1019 VSS.n11327 VSS.t3299 8.06917
R1020 VSS.n11342 VSS.t2370 8.06917
R1021 VSS.n102 VSS.t2402 8.06917
R1022 VSS.n11349 VSS.t2649 8.06917
R1023 VSS.n101 VSS.t1657 8.06917
R1024 VSS.n11355 VSS.t3377 8.06917
R1025 VSS.n97 VSS.t3419 8.06917
R1026 VSS.n10991 VSS.t513 8.06917
R1027 VSS.n10990 VSS.t2677 8.06917
R1028 VSS.n206 VSS.t2146 8.06917
R1029 VSS.n10986 VSS.t2182 8.06917
R1030 VSS.n10917 VSS.t2390 8.06917
R1031 VSS.n10916 VSS.t2422 8.06917
R1032 VSS.n10635 VSS.t3631 8.06917
R1033 VSS.n10635 VSS.t1370 8.06917
R1034 VSS.n10635 VSS.t1103 8.06917
R1035 VSS.n10635 VSS.t3485 8.06917
R1036 VSS.n10352 VSS.t1975 8.06917
R1037 VSS.n10640 VSS.t2398 8.06917
R1038 VSS.n10351 VSS.t785 8.06917
R1039 VSS.n10645 VSS.t2581 8.06917
R1040 VSS.n10350 VSS.t1647 8.06917
R1041 VSS.n10650 VSS.t2392 8.06917
R1042 VSS.n10346 VSS.t524 8.06917
R1043 VSS.n10516 VSS.t655 8.06917
R1044 VSS.n10508 VSS.t2843 8.06917
R1045 VSS.n10506 VSS.t2923 8.06917
R1046 VSS.n10502 VSS.t2282 8.06917
R1047 VSS.n10532 VSS.t1027 8.06917
R1048 VSS.n10491 VSS.t3169 8.06917
R1049 VSS.n10543 VSS.t3589 8.06917
R1050 VSS.n10487 VSS.t2625 8.06917
R1051 VSS.n10485 VSS.t1687 8.06917
R1052 VSS.n10590 VSS.t2835 8.06917
R1053 VSS.n10348 VSS.t1068 8.06917
R1054 VSS.n10510 VSS.t1165 8.06917
R1055 VSS.n10517 VSS.t872 8.06917
R1056 VSS.n10507 VSS.t565 8.06917
R1057 VSS.n10505 VSS.t2749 8.06917
R1058 VSS.n10500 VSS.t1891 8.06917
R1059 VSS.n10490 VSS.t698 8.06917
R1060 VSS.n10544 VSS.t1887 8.06917
R1061 VSS.n10486 VSS.t886 8.06917
R1062 VSS.n10484 VSS.t3055 8.06917
R1063 VSS.n10591 VSS.t1140 8.06917
R1064 VSS.n10496 VSS.t3119 8.06917
R1065 VSS.n10495 VSS.t781 8.06917
R1066 VSS.n10606 VSS.t508 8.06917
R1067 VSS.n10607 VSS.t2987 8.06917
R1068 VSS.n10609 VSS.t1470 8.06917
R1069 VSS.n10496 VSS.t1961 8.06917
R1070 VSS.n10495 VSS.t2751 8.06917
R1071 VSS.n10606 VSS.t2533 8.06917
R1072 VSS.n10607 VSS.t1833 8.06917
R1073 VSS.n10609 VSS.t3345 8.06917
R1074 VSS.n10412 VSS.t1468 8.06917
R1075 VSS.n10435 VSS.t3553 8.06917
R1076 VSS.n10413 VSS.t2575 8.06917
R1077 VSS.n10414 VSS.t657 8.06917
R1078 VSS.n10427 VSS.t2845 8.06917
R1079 VSS.n10415 VSS.t2925 8.06917
R1080 VSS.n10416 VSS.t2284 8.06917
R1081 VSS.n10420 VSS.t2366 8.06917
R1082 VSS.n10417 VSS.t1433 8.06917
R1083 VSS.n10477 VSS.t3243 8.06917
R1084 VSS.n10479 VSS.t3075 8.06917
R1085 VSS.n10480 VSS.t1695 8.06917
R1086 VSS.n10595 VSS.t2905 8.06917
R1087 VSS.n10594 VSS.t1614 8.06917
R1088 VSS.n10448 VSS.t1138 8.06917
R1089 VSS.n10457 VSS.t3255 8.06917
R1090 VSS.n10447 VSS.t3309 8.06917
R1091 VSS.n10446 VSS.t2731 8.06917
R1092 VSS.n10465 VSS.t1518 8.06917
R1093 VSS.n10445 VSS.t3599 8.06917
R1094 VSS.n10444 VSS.t920 8.06917
R1095 VSS.n10472 VSS.t3099 8.06917
R1096 VSS.n10443 VSS.t2112 8.06917
R1097 VSS.n10452 VSS.t1020 8.06917
R1098 VSS.n10450 VSS.t803 8.06917
R1099 VSS.n10449 VSS.t2539 8.06917
R1100 VSS.n10658 VSS.t622 8.06917
R1101 VSS.n10657 VSS.t2452 8.06917
R1102 VSS.n10585 VSS.t3257 8.06917
R1103 VSS.n10553 VSS.t3311 8.06917
R1104 VSS.n10554 VSS.t2733 8.06917
R1105 VSS.n10578 VSS.t2831 8.06917
R1106 VSS.n10555 VSS.t1853 8.06917
R1107 VSS.n10561 VSS.t1955 8.06917
R1108 VSS.n10559 VSS.t3173 8.06917
R1109 VSS.n10558 VSS.t850 8.06917
R1110 VSS.n10692 VSS.t595 8.06917
R1111 VSS.n10691 VSS.t3061 8.06917
R1112 VSS.n10689 VSS.t1530 8.06917
R1113 VSS.n1573 VSS.t1703 8.06917
R1114 VSS.n1573 VSS.t2745 8.06917
R1115 VSS.n1576 VSS.t855 8.06917
R1116 VSS.n1576 VSS.t1949 8.06917
R1117 VSS.n1577 VSS.t1215 8.06917
R1118 VSS.n1577 VSS.t2268 8.06917
R1119 VSS.n8958 VSS.t3121 8.06917
R1120 VSS.n8958 VSS.t1061 8.06917
R1121 VSS.n8959 VSS.t2713 8.06917
R1122 VSS.n8959 VSS.t611 8.06917
R1123 VSS.n8962 VSS.t957 8.06917
R1124 VSS.n8962 VSS.t2038 8.06917
R1125 VSS.n9035 VSS.t2873 8.06917
R1126 VSS.n9017 VSS.t797 8.06917
R1127 VSS.n1567 VSS.t1081 8.06917
R1128 VSS.n1566 VSS.t3463 8.06917
R1129 VSS.n8980 VSS.t2573 8.06917
R1130 VSS.n8980 VSS.t1814 8.06917
R1131 VSS.n8984 VSS.t1804 8.06917
R1132 VSS.n8984 VSS.t975 8.06917
R1133 VSS.n8985 VSS.t2116 8.06917
R1134 VSS.n8985 VSS.t1349 8.06917
R1135 VSS.n8993 VSS.t895 8.06917
R1136 VSS.n8993 VSS.t3223 8.06917
R1137 VSS.n8994 VSS.t3591 8.06917
R1138 VSS.n8994 VSS.t2841 8.06917
R1139 VSS.n8998 VSS.t1895 8.06917
R1140 VSS.n8998 VSS.t1087 8.06917
R1141 VSS.n8980 VSS.t3291 8.06917
R1142 VSS.n8980 VSS.t2601 8.06917
R1143 VSS.n8984 VSS.t2507 8.06917
R1144 VSS.n8984 VSS.t1818 8.06917
R1145 VSS.n8985 VSS.t2853 8.06917
R1146 VSS.n8985 VSS.t2138 8.06917
R1147 VSS.n8993 VSS.t1675 8.06917
R1148 VSS.n8993 VSS.t904 8.06917
R1149 VSS.n8994 VSS.t1255 8.06917
R1150 VSS.n8994 VSS.t3625 8.06917
R1151 VSS.n8998 VSS.t2615 8.06917
R1152 VSS.n8998 VSS.t1921 8.06917
R1153 VSS.n9004 VSS.t2170 8.06917
R1154 VSS.n8970 VSS.t3205 8.06917
R1155 VSS.n1565 VSS.t3471 8.06917
R1156 VSS.n8966 VSS.t2795 8.06917
R1157 VSS.n1553 VSS.t985 8.06917
R1158 VSS.n9096 VSS.t2066 8.06917
R1159 VSS.n8972 VSS.t1665 8.06917
R1160 VSS.n8971 VSS.t492 8.06917
R1161 VSS.n9080 VSS.t3069 8.06917
R1162 VSS.n9080 VSS.t978 8.06917
R1163 VSS.n9077 VSS.t2240 8.06917
R1164 VSS.n9077 VSS.t3283 8.06917
R1165 VSS.n9076 VSS.t2553 8.06917
R1166 VSS.n9076 VSS.t3617 8.06917
R1167 VSS.n9107 VSS.t1403 8.06917
R1168 VSS.n9107 VSS.t2426 8.06917
R1169 VSS.n9106 VSS.t943 8.06917
R1170 VSS.n9106 VSS.t2023 8.06917
R1171 VSS.n9103 VSS.t2328 8.06917
R1172 VSS.n9103 VSS.t3363 8.06917
R1173 VSS.n9080 VSS.t1504 8.06917
R1174 VSS.n9080 VSS.t3507 8.06917
R1175 VSS.n9077 VSS.t617 8.06917
R1176 VSS.n9077 VSS.t2717 8.06917
R1177 VSS.n9076 VSS.t973 8.06917
R1178 VSS.n9076 VSS.t3049 8.06917
R1179 VSS.n9107 VSS.t2919 8.06917
R1180 VSS.n9107 VSS.t1855 8.06917
R1181 VSS.n9106 VSS.t2468 8.06917
R1182 VSS.n9106 VSS.t1465 8.06917
R1183 VSS.n9103 VSS.t742 8.06917
R1184 VSS.n9103 VSS.t2825 8.06917
R1185 VSS.n9085 VSS.t1735 8.06917
R1186 VSS.n9045 VSS.t2791 8.06917
R1187 VSS.n1556 VSS.t2336 8.06917
R1188 VSS.n9041 VSS.t1296 8.06917
R1189 VSS.n9064 VSS.t1101 8.06917
R1190 VSS.n9047 VSS.t2194 8.06917
R1191 VSS.n9070 VSS.t2446 8.06917
R1192 VSS.n9046 VSS.t1767 8.06917
R1193 VSS.n962 VSS.t1293 8.06917
R1194 VSS.n962 VSS.t1024 8.06917
R1195 VSS.n960 VSS.t2088 8.06917
R1196 VSS.n960 VSS.t1857 8.06917
R1197 VSS.n959 VSS.t2491 8.06917
R1198 VSS.n959 VSS.t2266 8.06917
R1199 VSS.n10282 VSS.t2971 8.06917
R1200 VSS.n10282 VSS.t2719 8.06917
R1201 VSS.n10281 VSS.t1721 8.06917
R1202 VSS.n10281 VSS.t1496 8.06917
R1203 VSS.n10279 VSS.t3391 8.06917
R1204 VSS.n10279 VSS.t3179 8.06917
R1205 VSS.n953 VSS.t2154 8.06917
R1206 VSS.n971 VSS.t1913 8.06917
R1207 VSS.n954 VSS.t1389 8.06917
R1208 VSS.n965 VSS.t2184 8.06917
R1209 VSS.n950 VSS.t2565 8.06917
R1210 VSS.n950 VSS.t2701 8.06917
R1211 VSS.n947 VSS.t3335 8.06917
R1212 VSS.n947 VSS.t3465 8.06917
R1213 VSS.n946 VSS.t643 8.06917
R1214 VSS.n946 VSS.t774 8.06917
R1215 VSS.n10252 VSS.t1128 8.06917
R1216 VSS.n10252 VSS.t1264 8.06917
R1217 VSS.n10253 VSS.t3013 8.06917
R1218 VSS.n10253 VSS.t3115 8.06917
R1219 VSS.n10257 VSS.t1643 8.06917
R1220 VSS.n10257 VSS.t1753 8.06917
R1221 VSS.n950 VSS.t3033 8.06917
R1222 VSS.n950 VSS.t703 8.06917
R1223 VSS.n947 VSS.t683 8.06917
R1224 VSS.n947 VSS.t1553 8.06917
R1225 VSS.n946 VSS.t1132 8.06917
R1226 VSS.n946 VSS.t1957 8.06917
R1227 VSS.n10252 VSS.t1619 8.06917
R1228 VSS.n10252 VSS.t2380 8.06917
R1229 VSS.n10253 VSS.t3403 8.06917
R1230 VSS.n10253 VSS.t1148 8.06917
R1231 VSS.n10257 VSS.t2062 8.06917
R1232 VSS.n10257 VSS.t2893 8.06917
R1233 VSS.n10268 VSS.t1193 8.06917
R1234 VSS.n258 VSS.t916 8.06917
R1235 VSS.n10274 VSS.t3491 8.06917
R1236 VSS.n257 VSS.t1239 8.06917
R1237 VSS.n301 VSS.t3265 8.06917
R1238 VSS.n309 VSS.t3067 8.06917
R1239 VSS.n302 VSS.t2458 8.06917
R1240 VSS.n303 VSS.t2487 8.06917
R1241 VSS.n997 VSS.t1555 8.06917
R1242 VSS.n997 VSS.t1305 8.06917
R1243 VSS.n994 VSS.t2326 8.06917
R1244 VSS.n994 VSS.t2102 8.06917
R1245 VSS.n993 VSS.t2757 8.06917
R1246 VSS.n993 VSS.t2503 8.06917
R1247 VSS.n292 VSS.t3191 8.06917
R1248 VSS.n292 VSS.t2977 8.06917
R1249 VSS.n293 VSS.t1959 8.06917
R1250 VSS.n293 VSS.t1731 8.06917
R1251 VSS.n297 VSS.t486 8.06917
R1252 VSS.n297 VSS.t3401 8.06917
R1253 VSS.n997 VSS.t1993 8.06917
R1254 VSS.n997 VSS.t2013 8.06917
R1255 VSS.n994 VSS.t2803 8.06917
R1256 VSS.n994 VSS.t2839 8.06917
R1257 VSS.n993 VSS.t3197 8.06917
R1258 VSS.n993 VSS.t3227 8.06917
R1259 VSS.n292 VSS.t458 8.06917
R1260 VSS.n292 VSS.t500 8.06917
R1261 VSS.n293 VSS.t2394 8.06917
R1262 VSS.n293 VSS.t2430 8.06917
R1263 VSS.n297 VSS.t1008 8.06917
R1264 VSS.n297 VSS.t1055 8.06917
R1265 VSS.n942 VSS.t1115 8.06917
R1266 VSS.n987 VSS.t870 8.06917
R1267 VSS.n943 VSS.t3379 8.06917
R1268 VSS.n977 VSS.t3421 8.06917
R1269 VSS.n940 VSS.t2372 8.06917
R1270 VSS.n1008 VSS.t2162 8.06917
R1271 VSS.n941 VSS.t1631 8.06917
R1272 VSS.n1002 VSS.t2404 8.06917
R1273 VSS.n937 VSS.t3505 8.06917
R1274 VSS.n937 VSS.t2466 8.06917
R1275 VSS.n934 VSS.t1232 8.06917
R1276 VSS.n934 VSS.t3279 8.06917
R1277 VSS.n933 VSS.t1661 8.06917
R1278 VSS.n933 VSS.t549 8.06917
R1279 VSS.n10231 VSS.t2078 8.06917
R1280 VSS.n10231 VSS.t1051 8.06917
R1281 VSS.n10230 VSS.t810 8.06917
R1282 VSS.n10230 VSS.t2933 8.06917
R1283 VSS.n10227 VSS.t2549 8.06917
R1284 VSS.n10227 VSS.t1569 8.06917
R1285 VSS.n937 VSS.t3481 8.06917
R1286 VSS.n937 VSS.t2216 8.06917
R1287 VSS.n934 VSS.t1207 8.06917
R1288 VSS.n934 VSS.t3041 8.06917
R1289 VSS.n933 VSS.t1645 8.06917
R1290 VSS.n933 VSS.t3409 8.06917
R1291 VSS.n10231 VSS.t2060 8.06917
R1292 VSS.n10231 VSS.t759 8.06917
R1293 VSS.n10230 VSS.t791 8.06917
R1294 VSS.n10230 VSS.t2639 8.06917
R1295 VSS.n10227 VSS.t2535 8.06917
R1296 VSS.n10227 VSS.t1276 8.06917
R1297 VSS.n10218 VSS.t1472 8.06917
R1298 VSS.n10220 VSS.t1203 8.06917
R1299 VSS.n291 VSS.t593 8.06917
R1300 VSS.n315 VSS.t1494 8.06917
R1301 VSS.n10208 VSS.t3167 8.06917
R1302 VSS.n330 VSS.t3193 8.06917
R1303 VSS.n10214 VSS.t3399 8.06917
R1304 VSS.n329 VSS.t3443 8.06917
R1305 VSS.n1030 VSS.t2869 8.06917
R1306 VSS.n1030 VSS.t1849 8.06917
R1307 VSS.n1027 VSS.t463 8.06917
R1308 VSS.n1027 VSS.t2631 8.06917
R1309 VSS.n1026 VSS.t955 8.06917
R1310 VSS.n1026 VSS.t3089 8.06917
R1311 VSS.n10192 VSS.t1451 8.06917
R1312 VSS.n10192 VSS.t3487 8.06917
R1313 VSS.n10193 VSS.t3259 8.06917
R1314 VSS.n10193 VSS.t2262 8.06917
R1315 VSS.n10197 VSS.t1917 8.06917
R1316 VSS.n10197 VSS.t858 8.06917
R1317 VSS.n1030 VSS.t2160 8.06917
R1318 VSS.n1030 VSS.t1110 8.06917
R1319 VSS.n1027 VSS.t2969 8.06917
R1320 VSS.n1027 VSS.t1939 8.06917
R1321 VSS.n1026 VSS.t3329 8.06917
R1322 VSS.n1026 VSS.t2338 8.06917
R1323 VSS.n10192 VSS.t675 8.06917
R1324 VSS.n10192 VSS.t2813 8.06917
R1325 VSS.n10193 VSS.t2559 8.06917
R1326 VSS.n10193 VSS.t1573 8.06917
R1327 VSS.n10197 VSS.t1201 8.06917
R1328 VSS.n10197 VSS.t3261 8.06917
R1329 VSS.n929 VSS.t997 8.06917
R1330 VSS.n1020 VSS.t1036 8.06917
R1331 VSS.n930 VSS.t1302 8.06917
R1332 VSS.n1014 VSS.t1343 8.06917
R1333 VSS.n927 VSS.t2304 8.06917
R1334 VSS.n1045 VSS.t2332 8.06917
R1335 VSS.n928 VSS.t2945 8.06917
R1336 VSS.n1035 VSS.t1925 8.06917
R1337 VSS.n924 VSS.t2715 8.06917
R1338 VSS.n924 VSS.t2741 8.06917
R1339 VSS.n921 VSS.t3499 8.06917
R1340 VSS.n921 VSS.t3531 8.06917
R1341 VSS.n920 VSS.t807 8.06917
R1342 VSS.n920 VSS.t836 8.06917
R1343 VSS.n376 VSS.t1282 8.06917
R1344 VSS.n376 VSS.t1331 8.06917
R1345 VSS.n377 VSS.t3139 8.06917
R1346 VSS.n377 VSS.t3163 8.06917
R1347 VSS.n381 VSS.t1781 8.06917
R1348 VSS.n381 VSS.t1806 8.06917
R1349 VSS.n924 VSS.t1125 8.06917
R1350 VSS.n924 VSS.t876 8.06917
R1351 VSS.n921 VSS.t1947 8.06917
R1352 VSS.n921 VSS.t1715 8.06917
R1353 VSS.n920 VSS.t2352 8.06917
R1354 VSS.n920 VSS.t2126 8.06917
R1355 VSS.n376 VSS.t2823 8.06917
R1356 VSS.n376 VSS.t2557 8.06917
R1357 VSS.n377 VSS.t1589 8.06917
R1358 VSS.n377 VSS.t1337 8.06917
R1359 VSS.n381 VSS.t3271 8.06917
R1360 VSS.n381 VSS.t3073 8.06917
R1361 VSS.n364 VSS.t1387 8.06917
R1362 VSS.n372 VSS.t1421 8.06917
R1363 VSS.n365 VSS.t1983 8.06917
R1364 VSS.n366 VSS.t932 8.06917
R1365 VSS.n10158 VSS.t3373 8.06917
R1366 VSS.n10160 VSS.t3413 8.06917
R1367 VSS.n363 VSS.t503 8.06917
R1368 VSS.n387 VSS.t2669 8.06917
R1369 VSS.n1067 VSS.t1384 8.06917
R1370 VSS.n1067 VSS.t1425 8.06917
R1371 VSS.n1064 VSS.t2174 8.06917
R1372 VSS.n1064 VSS.t2204 8.06917
R1373 VSS.n1063 VSS.t2571 8.06917
R1374 VSS.n1063 VSS.t2609 8.06917
R1375 VSS.n10171 VSS.t3045 8.06917
R1376 VSS.n10171 VSS.t3093 8.06917
R1377 VSS.n10170 VSS.t1802 8.06917
R1378 VSS.n10170 VSS.t1831 8.06917
R1379 VSS.n10167 VSS.t3493 8.06917
R1380 VSS.n10167 VSS.t3527 8.06917
R1381 VSS.n1067 VSS.t2378 8.06917
R1382 VSS.n1067 VSS.t2168 8.06917
R1383 VSS.n1064 VSS.t3187 8.06917
R1384 VSS.n1064 VSS.t2973 8.06917
R1385 VSS.n1063 VSS.t3603 8.06917
R1386 VSS.n1063 VSS.t3337 8.06917
R1387 VSS.n10171 VSS.t946 8.06917
R1388 VSS.n10171 VSS.t689 8.06917
R1389 VSS.n10170 VSS.t2837 8.06917
R1390 VSS.n10170 VSS.t2567 8.06917
R1391 VSS.n10167 VSS.t1482 8.06917
R1392 VSS.n10167 VSS.t1211 8.06917
R1393 VSS.n916 VSS.t1278 8.06917
R1394 VSS.n1057 VSS.t1323 8.06917
R1395 VSS.n917 VSS.t1563 8.06917
R1396 VSS.n1051 VSS.t3605 8.06917
R1397 VSS.n914 VSS.t2673 8.06917
R1398 VSS.n1078 VSS.t3459 8.06917
R1399 VSS.n915 VSS.t2142 8.06917
R1400 VSS.n1072 VSS.t1903 8.06917
R1401 VSS.n911 VSS.t2645 8.06917
R1402 VSS.n911 VSS.t3423 8.06917
R1403 VSS.n908 VSS.t3411 8.06917
R1404 VSS.n908 VSS.t1154 8.06917
R1405 VSS.n907 VSS.t739 8.06917
R1406 VSS.n907 VSS.t1608 8.06917
R1407 VSS.n10132 VSS.t1230 8.06917
R1408 VSS.n10132 VSS.t2021 8.06917
R1409 VSS.n10133 VSS.t3097 8.06917
R1410 VSS.n10133 VSS.t747 8.06917
R1411 VSS.n10137 VSS.t1707 8.06917
R1412 VSS.n10137 VSS.t2485 8.06917
R1413 VSS.n911 VSS.t640 8.06917
R1414 VSS.n911 VSS.t3539 8.06917
R1415 VSS.n908 VSS.t1524 8.06917
R1416 VSS.n908 VSS.t1270 8.06917
R1417 VSS.n907 VSS.t1933 8.06917
R1418 VSS.n907 VSS.t1697 8.06917
R1419 VSS.n10132 VSS.t2354 8.06917
R1420 VSS.n10132 VSS.t2130 8.06917
R1421 VSS.n10133 VSS.t1099 8.06917
R1422 VSS.n10133 VSS.t852 8.06917
R1423 VSS.n10137 VSS.t2855 8.06917
R1424 VSS.n10137 VSS.t2593 8.06917
R1425 VSS.n10148 VSS.t1741 8.06917
R1426 VSS.n402 VSS.t2521 8.06917
R1427 VSS.n10154 VSS.t1181 8.06917
R1428 VSS.n401 VSS.t912 8.06917
R1429 VSS.n1283 VSS.t3315 8.06917
R1430 VSS.n1291 VSS.t3123 8.06917
R1431 VSS.n1284 VSS.t3611 8.06917
R1432 VSS.n1285 VSS.t3347 8.06917
R1433 VSS.n1104 VSS.t1272 8.06917
R1434 VSS.n1104 VSS.t989 8.06917
R1435 VSS.n1101 VSS.t2054 8.06917
R1436 VSS.n1101 VSS.t1835 8.06917
R1437 VSS.n1100 VSS.t2460 8.06917
R1438 VSS.n1100 VSS.t2238 8.06917
R1439 VSS.n1274 VSS.t2943 8.06917
R1440 VSS.n1274 VSS.t2703 8.06917
R1441 VSS.n1275 VSS.t1699 8.06917
R1442 VSS.n1275 VSS.t1474 8.06917
R1443 VSS.n1279 VSS.t3369 8.06917
R1444 VSS.n1279 VSS.t3161 8.06917
R1445 VSS.n1104 VSS.t1286 8.06917
R1446 VSS.n1104 VSS.t2096 8.06917
R1447 VSS.n1101 VSS.t2080 8.06917
R1448 VSS.n1101 VSS.t2903 8.06917
R1449 VSS.n1100 VSS.t2483 8.06917
R1450 VSS.n1100 VSS.t3287 8.06917
R1451 VSS.n1274 VSS.t2965 8.06917
R1452 VSS.n1274 VSS.t603 8.06917
R1453 VSS.n1275 VSS.t1717 8.06917
R1454 VSS.n1275 VSS.t2495 8.06917
R1455 VSS.n1279 VSS.t3387 8.06917
R1456 VSS.n1279 VSS.t1121 8.06917
R1457 VSS.n903 VSS.t1217 8.06917
R1458 VSS.n1094 VSS.t949 8.06917
R1459 VSS.n904 VSS.t1506 8.06917
R1460 VSS.n1084 VSS.t1248 8.06917
R1461 VSS.n901 VSS.t2931 8.06917
R1462 VSS.n1115 VSS.t2685 8.06917
R1463 VSS.n902 VSS.t1357 8.06917
R1464 VSS.n1109 VSS.t2150 8.06917
R1465 VSS.n878 VSS.t3503 8.06917
R1466 VSS.n1127 VSS.t3609 8.06917
R1467 VSS.n879 VSS.t3103 8.06917
R1468 VSS.n1121 VSS.t754 8.06917
R1469 VSS.n863 VSS.t2867 8.06917
R1470 VSS.n837 VSS.t2605 8.06917
R1471 VSS.n870 VSS.t2044 8.06917
R1472 VSS.n836 VSS.t2072 8.06917
R1473 VSS.n10923 VSS.t606 8.06917
R1474 VSS.n222 VSS.t3511 8.06917
R1475 VSS.n839 VSS.t2989 8.06917
R1476 VSS.n838 VSS.t630 8.06917
R1477 VSS.n858 VSS.t3235 8.06917
R1478 VSS.n858 VSS.t3027 8.06917
R1479 VSS.n855 VSS.t930 8.06917
R1480 VSS.n855 VSS.t670 8.06917
R1481 VSS.n854 VSS.t1407 8.06917
R1482 VSS.n854 VSS.t1119 8.06917
R1483 VSS.n848 VSS.t1837 8.06917
R1484 VSS.n848 VSS.t1612 8.06917
R1485 VSS.n847 VSS.t477 8.06917
R1486 VSS.n847 VSS.t3393 8.06917
R1487 VSS.n858 VSS.t536 8.06917
R1488 VSS.n858 VSS.t573 8.06917
R1489 VSS.n855 VSS.t1443 8.06917
R1490 VSS.n855 VSS.t1476 8.06917
R1491 VSS.n854 VSS.t1843 8.06917
R1492 VSS.n854 VSS.t1873 8.06917
R1493 VSS.n848 VSS.t2270 8.06917
R1494 VSS.n848 VSS.t2298 8.06917
R1495 VSS.n847 VSS.t1002 8.06917
R1496 VSS.n847 VSS.t1047 8.06917
R1497 VSS.n1135 VSS.t1197 8.06917
R1498 VSS.n1135 VSS.t926 8.06917
R1499 VSS.n1139 VSS.t1999 8.06917
R1500 VSS.n1139 VSS.t1779 8.06917
R1501 VSS.n1140 VSS.t2406 8.06917
R1502 VSS.n1140 VSS.t2190 8.06917
R1503 VSS.n1149 VSS.t2877 8.06917
R1504 VSS.n1149 VSS.t2617 8.06917
R1505 VSS.n1148 VSS.t1639 8.06917
R1506 VSS.n1148 VSS.t1405 8.06917
R1507 VSS.n1135 VSS.t1300 8.06917
R1508 VSS.n1135 VSS.t2108 8.06917
R1509 VSS.n1139 VSS.t2098 8.06917
R1510 VSS.n1139 VSS.t2911 8.06917
R1511 VSS.n1140 VSS.t2499 8.06917
R1512 VSS.n1140 VSS.t3293 8.06917
R1513 VSS.n1149 VSS.t2975 8.06917
R1514 VSS.n1149 VSS.t614 8.06917
R1515 VSS.n1148 VSS.t1729 8.06917
R1516 VSS.n1148 VSS.t2513 8.06917
R1517 VSS.n898 VSS.t3021 8.06917
R1518 VSS.n898 VSS.t2771 8.06917
R1519 VSS.n895 VSS.t665 8.06917
R1520 VSS.n895 VSS.t3557 8.06917
R1521 VSS.n894 VSS.t1113 8.06917
R1522 VSS.n894 VSS.t867 8.06917
R1523 VSS.n888 VSS.t1600 8.06917
R1524 VSS.n888 VSS.t1362 8.06917
R1525 VSS.n887 VSS.t3383 8.06917
R1526 VSS.n887 VSS.t3175 8.06917
R1527 VSS.n898 VSS.t3005 8.06917
R1528 VSS.n898 VSS.t649 8.06917
R1529 VSS.n895 VSS.t637 8.06917
R1530 VSS.n895 VSS.t1528 8.06917
R1531 VSS.n894 VSS.t1097 8.06917
R1532 VSS.n894 VSS.t1935 8.06917
R1533 VSS.n888 VSS.t1585 8.06917
R1534 VSS.n888 VSS.t2364 8.06917
R1535 VSS.n887 VSS.t3371 8.06917
R1536 VSS.n887 VSS.t1106 8.06917
R1537 VSS.n10353 VSS.t3445 8.06917
R1538 VSS.n10361 VSS.t2164 8.06917
R1539 VSS.n10354 VSS.t1175 8.06917
R1540 VSS.n10355 VSS.t1967 8.06917
R1541 VSS.n10666 VSS.t582 8.06917
R1542 VSS.n10338 VSS.t678 8.06917
R1543 VSS.n10337 VSS.t3535 8.06917
R1544 VSS.n10673 VSS.t3263 8.06917
R1545 VSS.n10336 VSS.t2300 8.06917
R1546 VSS.n10909 VSS.t1577 8.06917
R1547 VSS.n10909 VSS.t1333 8.06917
R1548 VSS.n10906 VSS.t2340 8.06917
R1549 VSS.n10906 VSS.t2124 8.06917
R1550 VSS.n10905 VSS.t2785 8.06917
R1551 VSS.n10905 VSS.t2531 8.06917
R1552 VSS.n10899 VSS.t3207 8.06917
R1553 VSS.n10899 VSS.t2993 8.06917
R1554 VSS.n10898 VSS.t1981 8.06917
R1555 VSS.n10898 VSS.t1757 8.06917
R1556 VSS.n10909 VSS.t2308 8.06917
R1557 VSS.n10909 VSS.t1317 8.06917
R1558 VSS.n10906 VSS.t3133 8.06917
R1559 VSS.n10906 VSS.t2106 8.06917
R1560 VSS.n10905 VSS.t3529 8.06917
R1561 VSS.n10905 VSS.t2509 8.06917
R1562 VSS.n10899 VSS.t863 8.06917
R1563 VSS.n10899 VSS.t2983 8.06917
R1564 VSS.n10898 VSS.t2735 8.06917
R1565 VSS.n10898 VSS.t1743 8.06917
R1566 VSS.n11003 VSS.t3601 8.06917
R1567 VSS.n11003 VSS.t2591 8.06917
R1568 VSS.n11007 VSS.t1339 8.06917
R1569 VSS.n11007 VSS.t3361 8.06917
R1570 VSS.n11008 VSS.t1765 8.06917
R1571 VSS.n11008 VSS.t680 8.06917
R1572 VSS.n11016 VSS.t2196 8.06917
R1573 VSS.n11016 VSS.t1167 8.06917
R1574 VSS.n11017 VSS.t907 8.06917
R1575 VSS.n11017 VSS.t3037 8.06917
R1576 VSS.n11003 VSS.t3241 8.06917
R1577 VSS.n11003 VSS.t2244 8.06917
R1578 VSS.n11007 VSS.t941 8.06917
R1579 VSS.n11007 VSS.t3071 8.06917
R1580 VSS.n11008 VSS.t1417 8.06917
R1581 VSS.n11008 VSS.t3433 8.06917
R1582 VSS.n11016 VSS.t1845 8.06917
R1583 VSS.n11016 VSS.t783 8.06917
R1584 VSS.n11017 VSS.t494 8.06917
R1585 VSS.n11017 VSS.t2663 8.06917
R1586 VSS.n11060 VSS.t692 8.06917
R1587 VSS.n11060 VSS.t732 8.06917
R1588 VSS.n11064 VSS.t1543 8.06917
R1589 VSS.n11064 VSS.t1581 8.06917
R1590 VSS.n11065 VSS.t1953 8.06917
R1591 VSS.n11065 VSS.t1989 8.06917
R1592 VSS.n11073 VSS.t2374 8.06917
R1593 VSS.n11073 VSS.t2412 8.06917
R1594 VSS.n11074 VSS.t1136 8.06917
R1595 VSS.n11074 VSS.t1171 8.06917
R1596 VSS.n11060 VSS.t2258 8.06917
R1597 VSS.n11060 VSS.t2005 8.06917
R1598 VSS.n11064 VSS.t3081 8.06917
R1599 VSS.n11064 VSS.t2827 8.06917
R1600 VSS.n11065 VSS.t3449 8.06917
R1601 VSS.n11065 VSS.t3219 8.06917
R1602 VSS.n11073 VSS.t794 8.06917
R1603 VSS.n11073 VSS.t489 8.06917
R1604 VSS.n11074 VSS.t2681 8.06917
R1605 VSS.n11074 VSS.t2418 8.06917
R1606 VSS.n1320 VSS.t1987 8.06917
R1607 VSS.t1987 VSS.n1319 8.06917
R1608 VSS.n1322 VSS.t1189 8.06917
R1609 VSS.t1189 VSS.n1321 8.06917
R1610 VSS.n1324 VSS.t1347 8.06917
R1611 VSS.t1347 VSS.n1323 8.06917
R1612 VSS.n1326 VSS.t3627 8.06917
R1613 VSS.t3627 VSS.n1325 8.06917
R1614 VSS.n1333 VSS.t2859 8.06917
R1615 VSS.t2859 VSS.n1332 8.06917
R1616 VSS.t2052 VSS.n9509 8.06917
R1617 VSS.n9510 VSS.t2052 8.06917
R1618 VSS.n9508 VSS.t2202 8.06917
R1619 VSS.t2202 VSS.n9507 8.06917
R1620 VSS.t1439 VSS.n9504 8.06917
R1621 VSS.n9505 VSS.t1439 8.06917
R1622 VSS.t744 VSS.n9501 8.06917
R1623 VSS.n9502 VSS.t744 8.06917
R1624 VSS.t1796 VSS.n9497 8.06917
R1625 VSS.n9498 VSS.t1796 8.06917
R1626 VSS.n1377 VSS.t2186 8.06917
R1627 VSS.t2186 VSS.n1376 8.06917
R1628 VSS.t1759 VSS.n9624 8.06917
R1629 VSS.n9625 VSS.t1759 8.06917
R1630 VSS.t1879 VSS.n9622 8.06917
R1631 VSS.n9623 VSS.t1879 8.06917
R1632 VSS.t1066 VSS.n9620 8.06917
R1633 VSS.n9621 VSS.t1066 8.06917
R1634 VSS.t3353 VSS.n9618 8.06917
R1635 VSS.n9619 VSS.t3353 8.06917
R1636 VSS.n815 VSS.t3519 8.06917
R1637 VSS.t3519 VSS.n810 8.06917
R1638 VSS.t2901 VSS.n9608 8.06917
R1639 VSS.n9609 VSS.t2901 8.06917
R1640 VSS.t2110 VSS.n9606 8.06917
R1641 VSS.n9607 VSS.t2110 8.06917
R1642 VSS.t1520 VSS.n9604 8.06917
R1643 VSS.n9605 VSS.t1520 8.06917
R1644 VSS.t663 VSS.n9602 8.06917
R1645 VSS.n9603 VSS.t663 8.06917
R1646 VSS.n9624 VSS.t542 8.06917
R1647 VSS.n9625 VSS.t542 8.06917
R1648 VSS.n9622 VSS.t723 8.06917
R1649 VSS.n9623 VSS.t723 8.06917
R1650 VSS.n9620 VSS.t3083 8.06917
R1651 VSS.n9621 VSS.t3083 8.06917
R1652 VSS.n9618 VSS.t2264 8.06917
R1653 VSS.n9619 VSS.t2264 8.06917
R1654 VSS.n815 VSS.t2382 8.06917
R1655 VSS.t2382 VSS.n810 8.06917
R1656 VSS.n9608 VSS.t1789 8.06917
R1657 VSS.n9609 VSS.t1789 8.06917
R1658 VSS.n9606 VSS.t963 8.06917
R1659 VSS.n9607 VSS.t963 8.06917
R1660 VSS.n9604 VSS.t3439 8.06917
R1661 VSS.n9605 VSS.t3439 8.06917
R1662 VSS.n9602 VSS.t2699 8.06917
R1663 VSS.n9603 VSS.t2699 8.06917
R1664 VSS.t1737 VSS.n9648 8.06917
R1665 VSS.n9649 VSS.t1737 8.06917
R1666 VSS.t1863 VSS.n9646 8.06917
R1667 VSS.n9647 VSS.t1863 8.06917
R1668 VSS.t1049 VSS.n9644 8.06917
R1669 VSS.n9645 VSS.t1049 8.06917
R1670 VSS.t3331 VSS.n649 8.06917
R1671 VSS.n9643 VSS.t3331 8.06917
R1672 VSS.n9886 VSS.t3495 8.06917
R1673 VSS.t3495 VSS.n9885 8.06917
R1674 VSS.n779 VSS.t2889 8.06917
R1675 VSS.t2889 VSS.n778 8.06917
R1676 VSS.n781 VSS.t2086 8.06917
R1677 VSS.t2086 VSS.n780 8.06917
R1678 VSS.n783 VSS.t1508 8.06917
R1679 VSS.t1508 VSS.n782 8.06917
R1680 VSS.n785 VSS.t635 8.06917
R1681 VSS.t635 VSS.n784 8.06917
R1682 VSS.n9648 VSS.t511 8.06917
R1683 VSS.n9649 VSS.t511 8.06917
R1684 VSS.n9646 VSS.t701 8.06917
R1685 VSS.n9647 VSS.t701 8.06917
R1686 VSS.n9644 VSS.t3057 8.06917
R1687 VSS.n9645 VSS.t3057 8.06917
R1688 VSS.t2254 VSS.n649 8.06917
R1689 VSS.n9643 VSS.t2254 8.06917
R1690 VSS.n9886 VSS.t2368 8.06917
R1691 VSS.n9885 VSS.t2368 8.06917
R1692 VSS.n779 VSS.t1775 8.06917
R1693 VSS.n778 VSS.t1775 8.06917
R1694 VSS.n781 VSS.t934 8.06917
R1695 VSS.n780 VSS.t934 8.06917
R1696 VSS.n783 VSS.t3415 8.06917
R1697 VSS.n782 VSS.t3415 8.06917
R1698 VSS.n785 VSS.t2661 8.06917
R1699 VSS.n784 VSS.t2661 8.06917
R1700 VSS.t1911 VSS.n9692 8.06917
R1701 VSS.n9693 VSS.t1911 8.06917
R1702 VSS.t1093 VSS.n9689 8.06917
R1703 VSS.n9690 VSS.t1093 8.06917
R1704 VSS.t3375 VSS.n9686 8.06917
R1705 VSS.n9687 VSS.t3375 8.06917
R1706 VSS.t3545 VSS.n9683 8.06917
R1707 VSS.n9684 VSS.t3545 8.06917
R1708 VSS.n1179 VSS.t2779 8.06917
R1709 VSS.t2779 VSS.n654 8.06917
R1710 VSS.t2144 VSS.n9852 8.06917
R1711 VSS.n9853 VSS.t2144 8.06917
R1712 VSS.t1372 VSS.n9849 8.06917
R1713 VSS.n9850 VSS.t1372 8.06917
R1714 VSS.t712 VSS.n9846 8.06917
R1715 VSS.n9847 VSS.t712 8.06917
R1716 VSS.t3077 VSS.n9843 8.06917
R1717 VSS.n9844 VSS.t3077 8.06917
R1718 VSS.n9691 VSS.t823 8.06917
R1719 VSS.t823 VSS.n9671 8.06917
R1720 VSS.n9688 VSS.t965 8.06917
R1721 VSS.t965 VSS.n9674 8.06917
R1722 VSS.n9685 VSS.t3277 8.06917
R1723 VSS.t3277 VSS.n9677 8.06917
R1724 VSS.t2489 VSS.n653 8.06917
R1725 VSS.n9680 VSS.t2489 8.06917
R1726 VSS.n1178 VSS.t2635 8.06917
R1727 VSS.t2635 VSS.n1177 8.06917
R1728 VSS.n9851 VSS.t2003 8.06917
R1729 VSS.t2003 VSS.n680 8.06917
R1730 VSS.n9848 VSS.t1241 8.06917
R1731 VSS.t1241 VSS.n683 8.06917
R1732 VSS.n9845 VSS.t539 8.06917
R1733 VSS.t539 VSS.n686 8.06917
R1734 VSS.n9842 VSS.t2939 8.06917
R1735 VSS.t2939 VSS.n689 8.06917
R1736 VSS.n661 VSS.t3467 8.06917
R1737 VSS.t3467 VSS.n578 8.06917
R1738 VSS.n663 VSS.t2711 8.06917
R1739 VSS.t2711 VSS.n662 8.06917
R1740 VSS.n665 VSS.t1927 8.06917
R1741 VSS.t1927 VSS.n664 8.06917
R1742 VSS.n667 VSS.t2042 8.06917
R1743 VSS.t2042 VSS.n666 8.06917
R1744 VSS.n673 VSS.t1268 8.06917
R1745 VSS.t1268 VSS.n668 8.06917
R1746 VSS.t560 VSS.n9870 8.06917
R1747 VSS.n9871 VSS.t560 8.06917
R1748 VSS.t2947 VSS.n9868 8.06917
R1749 VSS.n9869 VSS.t2947 8.06917
R1750 VSS.t2314 VSS.n9866 8.06917
R1751 VSS.n9867 VSS.t2314 8.06917
R1752 VSS.t1557 VSS.n9864 8.06917
R1753 VSS.n9865 VSS.t1557 8.06917
R1754 VSS.n661 VSS.t2348 8.06917
R1755 VSS.t2348 VSS.n578 8.06917
R1756 VSS.n663 VSS.t1598 8.06917
R1757 VSS.n662 VSS.t1598 8.06917
R1758 VSS.n665 VSS.t752 8.06917
R1759 VSS.n664 VSS.t752 8.06917
R1760 VSS.n667 VSS.t893 8.06917
R1761 VSS.n666 VSS.t893 8.06917
R1762 VSS.n673 VSS.t3217 8.06917
R1763 VSS.t3217 VSS.n668 8.06917
R1764 VSS.n9870 VSS.t2587 8.06917
R1765 VSS.n9871 VSS.t2587 8.06917
R1766 VSS.n9868 VSS.t1825 8.06917
R1767 VSS.n9869 VSS.t1825 8.06917
R1768 VSS.n9866 VSS.t1205 8.06917
R1769 VSS.n9867 VSS.t1205 8.06917
R1770 VSS.n9864 VSS.t3497 8.06917
R1771 VSS.n9865 VSS.t3497 8.06917
R1772 VSS.t2408 VSS.n9965 8.06917
R1773 VSS.n9966 VSS.t2408 8.06917
R1774 VSS.t1651 VSS.n9963 8.06917
R1775 VSS.n9964 VSS.t1651 8.06917
R1776 VSS.t819 VSS.n9961 8.06917
R1777 VSS.n9962 VSS.t819 8.06917
R1778 VSS.t953 VSS.n9959 8.06917
R1779 VSS.n9960 VSS.t953 8.06917
R1780 VSS.n141 VSS.t3267 8.06917
R1781 VSS.t3267 VSS.n140 8.06917
R1782 VSS.n11188 VSS.t2651 8.06917
R1783 VSS.t2651 VSS.n11187 8.06917
R1784 VSS.n11190 VSS.t1875 8.06917
R1785 VSS.t1875 VSS.n11189 8.06917
R1786 VSS.n11192 VSS.t1266 8.06917
R1787 VSS.t1266 VSS.n11191 8.06917
R1788 VSS.n11194 VSS.t3555 8.06917
R1789 VSS.t3555 VSS.n11193 8.06917
R1790 VSS.n9965 VSS.t1308 8.06917
R1791 VSS.n9966 VSS.t1308 8.06917
R1792 VSS.n9963 VSS.t3585 8.06917
R1793 VSS.n9964 VSS.t3585 8.06917
R1794 VSS.n9961 VSS.t2829 8.06917
R1795 VSS.n9962 VSS.t2829 8.06917
R1796 VSS.n9959 VSS.t2961 8.06917
R1797 VSS.n9960 VSS.t2961 8.06917
R1798 VSS.n141 VSS.t2172 8.06917
R1799 VSS.t2172 VSS.n140 8.06917
R1800 VSS.n11188 VSS.t1547 8.06917
R1801 VSS.n11187 VSS.t1547 8.06917
R1802 VSS.n11190 VSS.t715 8.06917
R1803 VSS.n11189 VSS.t715 8.06917
R1804 VSS.n11192 VSS.t3215 8.06917
R1805 VSS.n11191 VSS.t3215 8.06917
R1806 VSS.n11194 VSS.t2434 8.06917
R1807 VSS.n11193 VSS.t2434 8.06917
R1808 VSS.n1261 VSS.t2527 8.06917
R1809 VSS.t2527 VSS.n1260 8.06917
R1810 VSS.n1263 VSS.t1771 8.06917
R1811 VSS.t1771 VSS.n1262 8.06917
R1812 VSS.n1265 VSS.t1889 8.06917
R1813 VSS.t1889 VSS.n1264 8.06917
R1814 VSS.n1267 VSS.t1074 8.06917
R1815 VSS.t1074 VSS.n1266 8.06917
R1816 VSS.n9520 VSS.t3365 8.06917
R1817 VSS.t3365 VSS.n9519 8.06917
R1818 VSS.t2611 VSS.n1246 8.06917
R1819 VSS.n1247 VSS.t2611 8.06917
R1820 VSS.t2747 VSS.n1244 8.06917
R1821 VSS.n1245 VSS.t2747 8.06917
R1822 VSS.t1965 VSS.n1242 8.06917
R1823 VSS.n1243 VSS.t1965 8.06917
R1824 VSS.t1353 VSS.n804 8.06917
R1825 VSS.n1241 VSS.t1353 8.06917
R1826 VSS.n1261 VSS.t1413 8.06917
R1827 VSS.n1260 VSS.t1413 8.06917
R1828 VSS.n1263 VSS.t505 8.06917
R1829 VSS.n1262 VSS.t505 8.06917
R1830 VSS.n1265 VSS.t696 8.06917
R1831 VSS.n1264 VSS.t696 8.06917
R1832 VSS.n1267 VSS.t3053 8.06917
R1833 VSS.n1266 VSS.t3053 8.06917
R1834 VSS.n9520 VSS.t2252 8.06917
R1835 VSS.n9519 VSS.t2252 8.06917
R1836 VSS.n1246 VSS.t1486 8.06917
R1837 VSS.n1247 VSS.t1486 8.06917
R1838 VSS.n1244 VSS.t1627 8.06917
R1839 VSS.n1245 VSS.t1627 8.06917
R1840 VSS.n1242 VSS.t777 8.06917
R1841 VSS.n1243 VSS.t777 8.06917
R1842 VSS.t3253 VSS.n804 8.06917
R1843 VSS.n1241 VSS.t3253 8.06917
R1844 VSS.n635 VSS.t2362 8.06917
R1845 VSS.t2362 VSS.n634 8.06917
R1846 VSS.n637 VSS.t1602 8.06917
R1847 VSS.t1602 VSS.n636 8.06917
R1848 VSS.n639 VSS.t1727 8.06917
R1849 VSS.t1727 VSS.n638 8.06917
R1850 VSS.n641 VSS.t902 8.06917
R1851 VSS.t902 VSS.n640 8.06917
R1852 VSS.t3221 VSS.n9893 8.06917
R1853 VSS.n9894 VSS.t3221 8.06917
R1854 VSS.n9655 VSS.t2440 8.06917
R1855 VSS.t2440 VSS.n9654 8.06917
R1856 VSS.n9657 VSS.t2569 8.06917
R1857 VSS.t2569 VSS.n9656 8.06917
R1858 VSS.n9659 VSS.t1808 8.06917
R1859 VSS.t1808 VSS.n9658 8.06917
R1860 VSS.n9661 VSS.t1159 8.06917
R1861 VSS.t1159 VSS.n9660 8.06917
R1862 VSS.n635 VSS.t1219 8.06917
R1863 VSS.n634 VSS.t1219 8.06917
R1864 VSS.n637 VSS.t3515 8.06917
R1865 VSS.n636 VSS.t3515 8.06917
R1866 VSS.n639 VSS.t466 8.06917
R1867 VSS.n638 VSS.t466 8.06917
R1868 VSS.n641 VSS.t2881 8.06917
R1869 VSS.n640 VSS.t2881 8.06917
R1870 VSS.n9893 VSS.t2076 8.06917
R1871 VSS.n9894 VSS.t2076 8.06917
R1872 VSS.n9655 VSS.t1310 8.06917
R1873 VSS.n9654 VSS.t1310 8.06917
R1874 VSS.n9657 VSS.t1453 8.06917
R1875 VSS.n9656 VSS.t1453 8.06917
R1876 VSS.n9659 VSS.t578 8.06917
R1877 VSS.n9658 VSS.t578 8.06917
R1878 VSS.n9661 VSS.t3117 8.06917
R1879 VSS.n9660 VSS.t3117 8.06917
R1880 VSS.n601 VSS.t1659 8.06917
R1881 VSS.t1659 VSS.n546 8.06917
R1882 VSS.t821 VSS.n600 8.06917
R1883 VSS.n606 VSS.t821 8.06917
R1884 VSS.t959 VSS.n599 8.06917
R1885 VSS.n611 VSS.t959 8.06917
R1886 VSS.t3273 VSS.n598 8.06917
R1887 VSS.n616 VSS.t3273 8.06917
R1888 VSS.t2479 VSS.n9905 8.06917
R1889 VSS.n9906 VSS.t2479 8.06917
R1890 VSS.t2627 VSS.n9697 8.06917
R1891 VSS.n9698 VSS.t2627 8.06917
R1892 VSS.t1859 VSS.n9696 8.06917
R1893 VSS.n9703 VSS.t1859 8.06917
R1894 VSS.t1045 VSS.n9695 8.06917
R1895 VSS.n9708 VSS.t1045 8.06917
R1896 VSS.t1374 VSS.n9694 8.06917
R1897 VSS.n9713 VSS.t1374 8.06917
R1898 VSS.n605 VSS.t1500 8.06917
R1899 VSS.t1500 VSS.n604 8.06917
R1900 VSS.n610 VSS.t628 8.06917
R1901 VSS.t628 VSS.n609 8.06917
R1902 VSS.n615 VSS.t787 8.06917
R1903 VSS.t787 VSS.n614 8.06917
R1904 VSS.n620 VSS.t3137 8.06917
R1905 VSS.t3137 VSS.n619 8.06917
R1906 VSS.n9904 VSS.t2330 8.06917
R1907 VSS.t2330 VSS.n622 8.06917
R1908 VSS.n9702 VSS.t1579 8.06917
R1909 VSS.t1579 VSS.n9701 8.06917
R1910 VSS.n9707 VSS.t1705 8.06917
R1911 VSS.t1705 VSS.n9706 8.06917
R1912 VSS.n9712 VSS.t881 8.06917
R1913 VSS.t881 VSS.n9711 8.06917
R1914 VSS.n9717 VSS.t3323 8.06917
R1915 VSS.t3323 VSS.n9716 8.06917
R1916 VSS.n591 VSS.t2198 8.06917
R1917 VSS.t2198 VSS.n590 8.06917
R1918 VSS.n593 VSS.t1437 8.06917
R1919 VSS.t1437 VSS.n592 8.06917
R1920 VSS.n595 VSS.t1559 8.06917
R1921 VSS.t1559 VSS.n594 8.06917
R1922 VSS.n597 VSS.t725 8.06917
R1923 VSS.t725 VSS.n596 8.06917
R1924 VSS.t3087 VSS.n583 8.06917
R1925 VSS.n9917 VSS.t3087 8.06917
R1926 VSS.n9928 VSS.t3183 8.06917
R1927 VSS.t3183 VSS.n9927 8.06917
R1928 VSS.n9930 VSS.t2388 8.06917
R1929 VSS.t2388 VSS.n9929 8.06917
R1930 VSS.n9932 VSS.t1637 8.06917
R1931 VSS.t1637 VSS.n9931 8.06917
R1932 VSS.n9934 VSS.t1923 8.06917
R1933 VSS.t1923 VSS.n9933 8.06917
R1934 VSS.n591 VSS.t1010 8.06917
R1935 VSS.n590 VSS.t1010 8.06917
R1936 VSS.n593 VSS.t3305 8.06917
R1937 VSS.n592 VSS.t3305 8.06917
R1938 VSS.n595 VSS.t3461 8.06917
R1939 VSS.n594 VSS.t3461 8.06917
R1940 VSS.n597 VSS.t2707 8.06917
R1941 VSS.n596 VSS.t2707 8.06917
R1942 VSS.t1919 VSS.n583 8.06917
R1943 VSS.n9917 VSS.t1919 8.06917
R1944 VSS.n9928 VSS.t2029 8.06917
R1945 VSS.n9927 VSS.t2029 8.06917
R1946 VSS.n9930 VSS.t1260 8.06917
R1947 VSS.n9929 VSS.t1260 8.06917
R1948 VSS.n9932 VSS.t3549 8.06917
R1949 VSS.n9931 VSS.t3549 8.06917
R1950 VSS.n9934 VSS.t729 8.06917
R1951 VSS.n9933 VSS.t729 8.06917
R1952 VSS.t2815 VSS.n11049 8.06917
R1953 VSS.n11050 VSS.t2815 8.06917
R1954 VSS.t2007 VSS.n11047 8.06917
R1955 VSS.n11048 VSS.t2007 8.06917
R1956 VSS.t2156 VSS.n11045 8.06917
R1957 VSS.n11046 VSS.t2156 8.06917
R1958 VSS.t1380 VSS.n11043 8.06917
R1959 VSS.n11044 VSS.t1380 8.06917
R1960 VSS.n11282 VSS.t471 8.06917
R1961 VSS.t471 VSS.n11281 8.06917
R1962 VSS.n9948 VSS.t661 8.06917
R1963 VSS.t661 VSS.n9947 8.06917
R1964 VSS.n9950 VSS.t3031 8.06917
R1965 VSS.t3031 VSS.n9949 8.06917
R1966 VSS.n9952 VSS.t2220 8.06917
R1967 VSS.t2220 VSS.n9951 8.06917
R1968 VSS.n9954 VSS.t2505 8.06917
R1969 VSS.t2505 VSS.n9953 8.06917
R1970 VSS.n11049 VSS.t1667 8.06917
R1971 VSS.n11050 VSS.t1667 8.06917
R1972 VSS.n11047 VSS.t829 8.06917
R1973 VSS.n11048 VSS.t829 8.06917
R1974 VSS.n11045 VSS.t969 8.06917
R1975 VSS.n11046 VSS.t969 8.06917
R1976 VSS.n11043 VSS.t3281 8.06917
R1977 VSS.n11044 VSS.t3281 8.06917
R1978 VSS.n11282 VSS.t2501 8.06917
R1979 VSS.t2501 VSS.n11281 8.06917
R1980 VSS.n9948 VSS.t2647 8.06917
R1981 VSS.n9947 VSS.t2647 8.06917
R1982 VSS.n9950 VSS.t1871 8.06917
R1983 VSS.n9949 VSS.t1871 8.06917
R1984 VSS.n9952 VSS.t1057 8.06917
R1985 VSS.n9951 VSS.t1057 8.06917
R1986 VSS.n9954 VSS.t1393 8.06917
R1987 VSS.n9953 VSS.t1393 8.06917
R1988 VSS.t3231 VSS.n9476 8.06917
R1989 VSS.n9486 VSS.t3231 8.06917
R1990 VSS.t3349 VSS.n9484 8.06917
R1991 VSS.n9485 VSS.t3349 8.06917
R1992 VSS.t2583 VSS.n9482 8.06917
R1993 VSS.n9483 VSS.t2583 8.06917
R1994 VSS.t1816 VSS.n9480 8.06917
R1995 VSS.n9481 VSS.t1816 8.06917
R1996 VSS.n1387 VSS.t1945 8.06917
R1997 VSS.t1945 VSS.n1386 8.06917
R1998 VSS.n1409 VSS.t1327 8.06917
R1999 VSS.t1327 VSS.n1408 8.06917
R2000 VSS.n1411 VSS.t3607 8.06917
R2001 VSS.t3607 VSS.n1410 8.06917
R2002 VSS.n1413 VSS.t3023 8.06917
R2003 VSS.t3023 VSS.n1412 8.06917
R2004 VSS.n1415 VSS.t2214 8.06917
R2005 VSS.t2214 VSS.n1414 8.06917
R2006 VSS.n11220 VSS.t567 8.06917
R2007 VSS.n11220 VSS.t2665 8.06917
R2008 VSS.n11219 VSS.t918 8.06917
R2009 VSS.n11219 VSS.t3001 8.06917
R2010 VSS.n11213 VSS.t2875 8.06917
R2011 VSS.n11213 VSS.t1810 8.06917
R2012 VSS.n11212 VSS.t2442 8.06917
R2013 VSS.n11212 VSS.t1419 8.06917
R2014 VSS.n11209 VSS.t694 8.06917
R2015 VSS.n11209 VSS.t2767 8.06917
R2016 VSS.n11220 VSS.t1070 8.06917
R2017 VSS.n11220 VSS.t2158 8.06917
R2018 VSS.n11219 VSS.t1441 8.06917
R2019 VSS.n11219 VSS.t2454 8.06917
R2020 VSS.n11213 VSS.t3289 8.06917
R2021 VSS.n11213 VSS.t1284 8.06917
R2022 VSS.n11212 VSS.t2921 8.06917
R2023 VSS.n11212 VSS.t844 8.06917
R2024 VSS.n11209 VSS.t1179 8.06917
R2025 VSS.n11209 VSS.t2248 8.06917
R2026 VSS.n10956 VSS.t2537 8.06917
R2027 VSS.n10956 VSS.t3239 8.06917
R2028 VSS.n10957 VSS.t2883 8.06917
R2029 VSS.n10957 VSS.t3569 8.06917
R2030 VSS.n10965 VSS.t1701 8.06917
R2031 VSS.n10965 VSS.t2376 8.06917
R2032 VSS.n10966 VSS.t1280 8.06917
R2033 VSS.n10966 VSS.t1991 8.06917
R2034 VSS.n10970 VSS.t2641 8.06917
R2035 VSS.n10970 VSS.t3317 8.06917
R2036 VSS.n10956 VSS.t2222 8.06917
R2037 VSS.n10956 VSS.t2955 8.06917
R2038 VSS.n10957 VSS.t2541 8.06917
R2039 VSS.n10957 VSS.t3251 8.06917
R2040 VSS.n10965 VSS.t1395 8.06917
R2041 VSS.n10965 VSS.t2070 8.06917
R2042 VSS.n10966 VSS.t924 8.06917
R2043 VSS.n10966 VSS.t1691 8.06917
R2044 VSS.n10970 VSS.t2318 8.06917
R2045 VSS.n10970 VSS.t3065 8.06917
R2046 VSS.n722 VSS.t1312 8.06917
R2047 VSS.n722 VSS.t2342 8.06917
R2048 VSS.n721 VSS.t1641 8.06917
R2049 VSS.n721 VSS.t2695 8.06917
R2050 VSS.n715 VSS.t3517 8.06917
R2051 VSS.n715 VSS.t1516 8.06917
R2052 VSS.n714 VSS.t3127 8.06917
R2053 VSS.n714 VSS.t1063 8.06917
R2054 VSS.n711 VSS.t1423 8.06917
R2055 VSS.n711 VSS.t2448 8.06917
R2056 VSS.n722 VSS.t3615 8.06917
R2057 VSS.n722 VSS.t1252 8.06917
R2058 VSS.n721 VSS.t825 8.06917
R2059 VSS.n721 VSS.t1587 8.06917
R2060 VSS.n715 VSS.t2759 8.06917
R2061 VSS.n715 VSS.t3441 8.06917
R2062 VSS.n714 VSS.t2334 8.06917
R2063 VSS.n714 VSS.t3095 8.06917
R2064 VSS.n711 VSS.t557 8.06917
R2065 VSS.n711 VSS.t1364 8.06917
R2066 VSS.n1169 VSS.t2897 8.06917
R2067 VSS.n1169 VSS.t827 8.06917
R2068 VSS.n1170 VSS.t3199 8.06917
R2069 VSS.n1170 VSS.t1173 8.06917
R2070 VSS.n1190 VSS.t2017 8.06917
R2071 VSS.n1190 VSS.t3107 8.06917
R2072 VSS.n1191 VSS.t1635 8.06917
R2073 VSS.n1191 VSS.t2691 8.06917
R2074 VSS.n1195 VSS.t3003 8.06917
R2075 VSS.n1195 VSS.t928 8.06917
R2076 VSS.n1169 VSS.t1341 8.06917
R2077 VSS.n1169 VSS.t3319 8.06917
R2078 VSS.n1170 VSS.t1669 8.06917
R2079 VSS.n1170 VSS.t497 8.06917
R2080 VSS.n1190 VSS.t3541 8.06917
R2081 VSS.n1190 VSS.t2470 8.06917
R2082 VSS.n1191 VSS.t3149 8.06917
R2083 VSS.n1191 VSS.t2084 8.06917
R2084 VSS.n1195 VSS.t1449 8.06917
R2085 VSS.n1195 VSS.t3431 8.06917
R2086 VSS.n9147 VSS.t3009 8.06917
R2087 VSS.n9147 VSS.t533 8.06917
R2088 VSS.n9151 VSS.t2200 8.06917
R2089 VSS.n9151 VSS.t2915 8.06917
R2090 VSS.n9152 VSS.t2497 8.06917
R2091 VSS.n9152 VSS.t3211 8.06917
R2092 VSS.n9160 VSS.t1345 8.06917
R2093 VSS.n9160 VSS.t2027 8.06917
R2094 VSS.n9161 VSS.t890 8.06917
R2095 VSS.n9161 VSS.t1649 8.06917
R2096 VSS.n9165 VSS.t2278 8.06917
R2097 VSS.n9165 VSS.t3019 8.06917
R2098 VSS.n9147 VSS.t1447 8.06917
R2099 VSS.n9147 VSS.t2140 8.06917
R2100 VSS.n9151 VSS.t544 8.06917
R2101 VSS.n9151 VSS.t1359 8.06917
R2102 VSS.n9152 VSS.t910 8.06917
R2103 VSS.n9152 VSS.t1677 8.06917
R2104 VSS.n9160 VSS.t2865 8.06917
R2105 VSS.n9160 VSS.t3551 8.06917
R2106 VSS.n9161 VSS.t2436 8.06917
R2107 VSS.n9161 VSS.t3155 8.06917
R2108 VSS.n9165 VSS.t673 8.06917
R2109 VSS.n9165 VSS.t1457 8.06917
R2110 VSS.t2036 VSS.t312 7.5006
R2111 VSS.t2475 VSS.t433 7.5006
R2112 VSS.t429 VSS.t1237 7.5006
R2113 VSS.n572 VSS.t117 7.42489
R2114 VSS.t60 VSS.n565 7.41222
R2115 VSS.n9890 VSS.t307 7.25283
R2116 VSS.n11391 VSS.n60 7.08065
R2117 VSS.n10308 VSS.t280 6.72766
R2118 VSS.t337 VSS.t540 6.61526
R2119 VSS.n10760 VSS.t2917 6.60917
R2120 VSS.n10760 VSS.t1593 6.60917
R2121 VSS.n10760 VSS.t3341 6.60917
R2122 VSS.n10760 VSS.t1997 6.60917
R2123 VSS.n10760 VSS.t3035 6.60917
R2124 VSS.n10738 VSS.t563 6.60917
R2125 VSS.n10764 VSS.t659 6.60917
R2126 VSS.n10740 VSS.t718 6.60917
R2127 VSS.n10759 VSS.t789 6.60917
R2128 VSS.n10774 VSS.t3147 6.60917
R2129 VSS.n10771 VSS.t1820 6.60917
R2130 VSS.n10856 VSS.t3597 6.60917
R2131 VSS.n10854 VSS.t2226 6.60917
R2132 VSS.n10743 VSS.t3237 6.60917
R2133 VSS.n10388 VSS.t202 6.53862
R2134 VSS.n9347 VSS.n9346 6.4661
R2135 VSS.n9422 VSS.n1383 6.4661
R2136 VSS.t103 VSS.t339 6.21678
R2137 VSS.t1244 VSS.t384 5.81954
R2138 VSS.t107 VSS.t490 5.8183
R2139 VSS.t108 VSS.t795 5.8183
R2140 VSS.n10739 VSS.t187 5.49372
R2141 VSS.n10306 VSS.t199 5.47432
R2142 VSS.t377 VSS.t256 5.34013
R2143 VSS.n10032 VSS.n566 5.34013
R2144 VSS.n10301 VSS.n10300 5.31981
R2145 VSS.n10392 VSS.t30 5.28484
R2146 VSS.n10397 VSS.t128 5.28484
R2147 VSS.n10391 VSS.t212 5.28484
R2148 VSS.n10305 VSS.n10292 5.26136
R2149 VSS.n10761 VSS.t2918 5.2505
R2150 VSS.t2918 VSS.n241 5.2505
R2151 VSS.n10761 VSS.t1595 5.2505
R2152 VSS.t1595 VSS.n241 5.2505
R2153 VSS.n10761 VSS.t3342 5.2505
R2154 VSS.t3342 VSS.n241 5.2505
R2155 VSS.n10761 VSS.t1998 5.2505
R2156 VSS.t1998 VSS.n241 5.2505
R2157 VSS.n10761 VSS.t3036 5.2505
R2158 VSS.t3036 VSS.n241 5.2505
R2159 VSS.n10768 VSS.t564 5.2505
R2160 VSS.n10763 VSS.t660 5.2505
R2161 VSS.t790 VSS.n10739 5.2505
R2162 VSS.t719 VSS.n10755 5.2505
R2163 VSS.n10410 VSS.n10409 5.16888
R2164 VSS.n10374 VSS.n10373 5.15456
R2165 VSS.n10680 VSS.n10679 5.09675
R2166 VSS.t609 VSS.t506 4.94165
R2167 VSS.n10066 VSS.t537 4.78226
R2168 VSS.n10626 VSS.n10623 4.63106
R2169 VSS.n10617 VSS.n10614 4.63106
R2170 VSS.n10381 VSS.n10378 4.63106
R2171 VSS.n10302 VSS.n10301 4.61712
R2172 VSS.n10684 VSS.n10683 4.61712
R2173 VSS.n10806 VSS.n10802 4.61585
R2174 VSS.n10800 VSS.n10796 4.61585
R2175 VSS.n9196 VSS.n9195 4.61205
R2176 VSS.n9191 VSS.n9190 4.61205
R2177 VSS.n9332 VSS.n9331 4.61205
R2178 VSS.n9327 VSS.n9326 4.61205
R2179 VSS.n170 VSS.n169 4.61205
R2180 VSS.n165 VSS.n164 4.61205
R2181 VSS.n9578 VSS.n9577 4.61205
R2182 VSS.n9573 VSS.n9572 4.61205
R2183 VSS.n193 VSS.n192 4.61205
R2184 VSS.n198 VSS.n197 4.61205
R2185 VSS.n471 VSS.n470 4.61205
R2186 VSS.n476 VSS.n475 4.61205
R2187 VSS.n9029 VSS.n9028 4.61205
R2188 VSS.n9024 VSS.n9023 4.61205
R2189 VSS.n264 VSS.n263 4.61205
R2190 VSS.n269 VSS.n268 4.61205
R2191 VSS.n336 VSS.n335 4.61205
R2192 VSS.n341 VSS.n340 4.61205
R2193 VSS.n408 VSS.n407 4.61205
R2194 VSS.n413 VSS.n412 4.61205
R2195 VSS.n10630 VSS.n10628 4.61078
R2196 VSS.n10621 VSS.n10619 4.61078
R2197 VSS.n10385 VSS.n10383 4.61078
R2198 VSS.n10376 VSS.n10374 4.61078
R2199 VSS.n10682 VSS.n10681 4.61078
R2200 VSS.n10631 VSS.n10630 4.60825
R2201 VSS.n10622 VSS.n10621 4.60825
R2202 VSS.n10386 VSS.n10385 4.60825
R2203 VSS.n10377 VSS.n10376 4.60825
R2204 VSS.n10681 VSS.n10680 4.60825
R2205 VSS.n10309 VSS.n10306 4.60439
R2206 VSS.n10807 VSS.n10806 4.60318
R2207 VSS.n10801 VSS.n10800 4.60318
R2208 VSS.n10303 VSS.n10302 4.60191
R2209 VSS.n10685 VSS.n10684 4.60191
R2210 VSS.n10627 VSS.n10626 4.58796
R2211 VSS.n10618 VSS.n10617 4.58796
R2212 VSS.n10382 VSS.n10381 4.58796
R2213 VSS.n9194 VSS.n9193 4.5005
R2214 VSS.n9189 VSS.n9188 4.5005
R2215 VSS.n9330 VSS.n9329 4.5005
R2216 VSS.n9325 VSS.n9324 4.5005
R2217 VSS.n168 VSS.n167 4.5005
R2218 VSS.n163 VSS.n162 4.5005
R2219 VSS.n9576 VSS.n9575 4.5005
R2220 VSS.n9571 VSS.n9570 4.5005
R2221 VSS.n191 VSS.n190 4.5005
R2222 VSS.n196 VSS.n195 4.5005
R2223 VSS.n469 VSS.n468 4.5005
R2224 VSS.n474 VSS.n473 4.5005
R2225 VSS.n10798 VSS.n10795 4.5005
R2226 VSS.n10804 VSS.n10794 4.5005
R2227 VSS.n9027 VSS.n9026 4.5005
R2228 VSS.n9022 VSS.n9021 4.5005
R2229 VSS.n9019 VSS.n9018 4.5005
R2230 VSS.n9019 VSS.n1560 4.5005
R2231 VSS.n9034 VSS.n9033 4.5005
R2232 VSS.n9033 VSS.n9032 4.5005
R2233 VSS.n262 VSS.n261 4.5005
R2234 VSS.n267 VSS.n266 4.5005
R2235 VSS.n334 VSS.n333 4.5005
R2236 VSS.n339 VSS.n338 4.5005
R2237 VSS.n406 VSS.n405 4.5005
R2238 VSS.n411 VSS.n410 4.5005
R2239 VSS.n10144 VSS.n10143 4.5005
R2240 VSS.n10143 VSS.n403 4.5005
R2241 VSS.n10146 VSS.n10145 4.5005
R2242 VSS.n10147 VSS.n10146 4.5005
R2243 VSS.n10204 VSS.n10203 4.5005
R2244 VSS.n10203 VSS.n331 4.5005
R2245 VSS.n10206 VSS.n10205 4.5005
R2246 VSS.n10207 VSS.n10206 4.5005
R2247 VSS.n10264 VSS.n10263 4.5005
R2248 VSS.n10263 VSS.n259 4.5005
R2249 VSS.n10266 VSS.n10265 4.5005
R2250 VSS.n10267 VSS.n10266 4.5005
R2251 VSS.n10571 VSS.n10570 4.5005
R2252 VSS.n10570 VSS.n10569 4.5005
R2253 VSS.n10569 VSS.n10556 4.5005
R2254 VSS.n10563 VSS.n10556 4.5005
R2255 VSS.n10572 VSS.n10563 4.5005
R2256 VSS.n10572 VSS.n10557 4.5005
R2257 VSS.n10572 VSS.n10571 4.5005
R2258 VSS.n10375 VSS.n10372 4.5005
R2259 VSS.n10380 VSS.n10371 4.5005
R2260 VSS.n10384 VSS.n10370 4.5005
R2261 VSS.n10616 VSS.n10369 4.5005
R2262 VSS.n10620 VSS.n10368 4.5005
R2263 VSS.n10625 VSS.n10367 4.5005
R2264 VSS.n10629 VSS.n10366 4.5005
R2265 VSS.n10294 VSS.n10293 4.5005
R2266 VSS.n10297 VSS.n10295 4.5005
R2267 VSS.n10299 VSS.n10298 4.5005
R2268 VSS.n10913 VSS.n226 4.5005
R2269 VSS.n10913 VSS.n229 4.5005
R2270 VSS.n10913 VSS.n225 4.5005
R2271 VSS.n10913 VSS.n10912 4.5005
R2272 VSS.n229 VSS.n223 4.5005
R2273 VSS.n225 VSS.n223 4.5005
R2274 VSS.n10912 VSS.n223 4.5005
R2275 VSS.n11338 VSS.n108 4.5005
R2276 VSS.n11337 VSS.n103 4.5005
R2277 VSS.n11338 VSS.n106 4.5005
R2278 VSS.n11338 VSS.n109 4.5005
R2279 VSS.n11338 VSS.n11337 4.5005
R2280 VSS.n11337 VSS.n11336 4.5005
R2281 VSS.n11336 VSS.n109 4.5005
R2282 VSS.n11336 VSS.n106 4.5005
R2283 VSS.n11336 VSS.n108 4.5005
R2284 VSS.n483 VSS.n482 4.5005
R2285 VSS.n482 VSS.n466 4.5005
R2286 VSS.n480 VSS.n463 4.5005
R2287 VSS.n480 VSS.n479 4.5005
R2288 VSS.n11141 VSS.n11140 4.5005
R2289 VSS.n11140 VSS.n188 4.5005
R2290 VSS.n11143 VSS.n11142 4.5005
R2291 VSS.n11144 VSS.n11143 4.5005
R2292 VSS.n11432 VSS.n11431 4.5005
R2293 VSS.n11431 VSS.n11430 4.5005
R2294 VSS.n11429 VSS.n32 4.5005
R2295 VSS.n11430 VSS.n11429 4.5005
R2296 VSS.n11433 VSS.n32 4.5005
R2297 VSS.n11433 VSS.n30 4.5005
R2298 VSS.n11433 VSS.n11432 4.5005
R2299 VSS.n11400 VSS.n56 4.5005
R2300 VSS.n11400 VSS.n11399 4.5005
R2301 VSS.n11396 VSS.n57 4.5005
R2302 VSS.n57 VSS.n56 4.5005
R2303 VSS.n11399 VSS.n57 4.5005
R2304 VSS.n11398 VSS.n11396 4.5005
R2305 VSS.n11399 VSS.n11398 4.5005
R2306 VSS.n11384 VSS.n62 4.5005
R2307 VSS.n11387 VSS.n11383 4.5005
R2308 VSS.n11383 VSS.n78 4.5005
R2309 VSS.n11388 VSS.n78 4.5005
R2310 VSS.n11386 VSS.n78 4.5005
R2311 VSS.n11388 VSS.n11387 4.5005
R2312 VSS.n11387 VSS.n62 4.5005
R2313 VSS.n11387 VSS.n83 4.5005
R2314 VSS.n11387 VSS.n11386 4.5005
R2315 VSS.n9582 VSS.n9568 4.5005
R2316 VSS.n9583 VSS.n9582 4.5005
R2317 VSS.n9586 VSS.n9585 4.5005
R2318 VSS.n9585 VSS.n9584 4.5005
R2319 VSS.n160 VSS.n159 4.5005
R2320 VSS.n160 VSS.n157 4.5005
R2321 VSS.n176 VSS.n175 4.5005
R2322 VSS.n175 VSS.n174 4.5005
R2323 VSS.n9335 VSS.n9322 4.5005
R2324 VSS.n9336 VSS.n9335 4.5005
R2325 VSS.n9339 VSS.n9338 4.5005
R2326 VSS.n9338 VSS.n9337 4.5005
R2327 VSS.n9186 VSS.n9185 4.5005
R2328 VSS.n9186 VSS.n1522 4.5005
R2329 VSS.n9201 VSS.n9200 4.5005
R2330 VSS.n9200 VSS.n9199 4.5005
R2331 VSS.n11310 VSS.n11309 4.5005
R2332 VSS.n11305 VSS.n122 4.5005
R2333 VSS.n11305 VSS.n124 4.5005
R2334 VSS.n11309 VSS.n11308 4.5005
R2335 VSS.n11308 VSS.n11307 4.5005
R2336 VSS.n11308 VSS.n122 4.5005
R2337 VSS.n11308 VSS.n124 4.5005
R2338 VSS.n10732 VSS.n10731 4.5005
R2339 VSS.n10728 VSS.n10707 4.5005
R2340 VSS.n10729 VSS.n10728 4.5005
R2341 VSS.n10731 VSS.n10730 4.5005
R2342 VSS.n10730 VSS.n10704 4.5005
R2343 VSS.n10730 VSS.n10707 4.5005
R2344 VSS.n10730 VSS.n10729 4.5005
R2345 VSS.n10322 VSS.t206 4.41563
R2346 VSS.n10331 VSS.t34 4.41563
R2347 VSS.n10320 VSS.t143 4.41563
R2348 VSS.n10310 VSS.t142 4.41563
R2349 VSS.t1794 VSS.t633 4.2678
R2350 VSS.n10404 VSS.t11 4.22616
R2351 VSS.n10402 VSS.t179 4.22616
R2352 VSS.n10308 VSS.n10307 4.21432
R2353 VSS.n10305 VSS.n10304 4.21432
R2354 VSS.n9884 VSS.n9883 4.21138
R2355 VSS.n9881 VSS.n9880 4.21138
R2356 VSS.n9879 VSS.n9878 4.21138
R2357 VSS.n9518 VSS.n642 4.21138
R2358 VSS.n9896 VSS.n9895 4.21138
R2359 VSS.n9914 VSS.n9907 4.21138
R2360 VSS.n9919 VSS.n9918 4.21138
R2361 VSS.n678 VSS.n648 4.21074
R2362 VSS.n9859 VSS.n9854 4.21074
R2363 VSS.n9873 VSS.n9872 4.21074
R2364 VSS.n1255 VSS.n1254 4.21074
R2365 VSS.n9902 VSS.n628 4.21074
R2366 VSS.n627 VSS.n584 4.21074
R2367 VSS.n9926 VSS.n9925 4.21074
R2368 VSS.n11450 VSS.n19 4.21074
R2369 VSS.n11445 VSS.n22 4.21074
R2370 VSS.n11417 VSS.n44 4.21074
R2371 VSS.n11412 VSS.n47 4.21074
R2372 VSS.n9617 VSS.n650 4.21074
R2373 VSS.n9610 VSS.n822 4.21074
R2374 VSS.n9616 VSS.n811 4.21074
R2375 VSS.n9611 VSS.n814 4.21074
R2376 VSS.n9517 VSS.n1327 4.21074
R2377 VSS.n9512 VSS.n9511 4.21074
R2378 VSS.n9611 VSS.n9610 4.19858
R2379 VSS.n822 VSS.n648 4.19794
R2380 VSS.n9884 VSS.n650 4.19794
R2381 VSS.n679 VSS.n678 4.19794
R2382 VSS.n9883 VSS.n9882 4.19794
R2383 VSS.n9872 VSS.n9859 4.19794
R2384 VSS.n9880 VSS.n9879 4.19794
R2385 VSS.n9512 VSS.n1255 4.19794
R2386 VSS.n9518 VSS.n9517 4.19794
R2387 VSS.n1254 VSS.n628 4.19794
R2388 VSS.n9895 VSS.n642 4.19794
R2389 VSS.n9903 VSS.n9902 4.19794
R2390 VSS.n9896 VSS.n621 4.19794
R2391 VSS.n9926 VSS.n584 4.19794
R2392 VSS.n9918 VSS.n9914 4.19794
R2393 VSS.n9925 VSS.n22 4.19794
R2394 VSS.n9919 VSS.n19 4.19794
R2395 VSS.n9873 VSS.n47 4.19794
R2396 VSS.n9878 VSS.n44 4.19794
R2397 VSS.n9617 VSS.n9616 4.19794
R2398 VSS.n11445 VSS.n11444 4.19794
R2399 VSS.n11451 VSS.n11450 4.19794
R2400 VSS.n11412 VSS.n11411 4.19794
R2401 VSS.n11418 VSS.n11417 4.19794
R2402 VSS.n9192 VSS.t356 4.16335
R2403 VSS.n9187 VSS.t360 4.16335
R2404 VSS.n9328 VSS.t388 4.16335
R2405 VSS.n9323 VSS.t382 4.16335
R2406 VSS.n166 VSS.t374 4.16335
R2407 VSS.n161 VSS.t369 4.16335
R2408 VSS.n9574 VSS.t3635 4.16335
R2409 VSS.n9569 VSS.t444 4.16335
R2410 VSS.n9025 VSS.t414 4.16335
R2411 VSS.n9020 VSS.t416 4.16335
R2412 VSS.n189 VSS.t169 4.16278
R2413 VSS.n194 VSS.t189 4.16278
R2414 VSS.n467 VSS.t406 4.16278
R2415 VSS.n472 VSS.t400 4.16278
R2416 VSS.n260 VSS.t300 4.16278
R2417 VSS.n265 VSS.t303 4.16278
R2418 VSS.n332 VSS.t3639 4.16278
R2419 VSS.n337 VSS.t3643 4.16278
R2420 VSS.n404 VSS.t320 4.16278
R2421 VSS.n409 VSS.t322 4.16278
R2422 VSS.n9195 VSS.t359 4.16103
R2423 VSS.n9190 VSS.t362 4.16103
R2424 VSS.n9331 VSS.t386 4.16103
R2425 VSS.n9326 VSS.t389 4.16103
R2426 VSS.n169 VSS.t368 4.16103
R2427 VSS.n164 VSS.t371 4.16103
R2428 VSS.n9577 VSS.t3636 4.16103
R2429 VSS.n9572 VSS.t445 4.16103
R2430 VSS.n9028 VSS.t415 4.16103
R2431 VSS.n9023 VSS.t3645 4.16103
R2432 VSS.n192 VSS.t188 4.15984
R2433 VSS.n197 VSS.t167 4.15984
R2434 VSS.n470 VSS.t403 4.15984
R2435 VSS.n475 VSS.t407 4.15984
R2436 VSS.n263 VSS.t296 4.15984
R2437 VSS.n268 VSS.t301 4.15984
R2438 VSS.n335 VSS.t3640 4.15984
R2439 VSS.n340 VSS.t3644 4.15984
R2440 VSS.n407 VSS.t325 4.15984
R2441 VSS.n412 VSS.t327 4.15984
R2442 VSS.n10565 VSS.n128 4.1417
R2443 VSS.t258 VSS.n434 4.06499
R2444 VSS.n1346 VSS.t1478 4.03583
R2445 VSS.n1371 VSS.t2166 4.03583
R2446 VSS.n1348 VSS.t1761 4.03583
R2447 VSS.n1365 VSS.t995 4.03583
R2448 VSS.n1351 VSS.t2653 4.03583
R2449 VSS.n1359 VSS.t3325 4.03583
R2450 VSS.n1354 VSS.t2623 4.03583
R2451 VSS.n803 VSS.t600 4.03583
R2452 VSS.n802 VSS.t2687 4.03583
R2453 VSS.n801 VSS.t3427 4.03583
R2454 VSS.n798 VSS.t991 4.03583
R2455 VSS.n800 VSS.t3079 4.03583
R2456 VSS.n9636 VSS.t2629 4.03583
R2457 VSS.n9756 VSS.t517 4.03583
R2458 VSS.n9638 VSS.t2613 4.03583
R2459 VSS.n9662 VSS.t584 4.03583
R2460 VSS.n9663 VSS.t2655 4.03583
R2461 VSS.n9746 VSS.t1951 4.03583
R2462 VSS.n9665 VSS.t3563 4.03583
R2463 VSS.n9740 VSS.t1187 4.03583
R2464 VSS.n9668 VSS.t3165 4.03583
R2465 VSS.n9734 VSS.t2114 4.03583
R2466 VSS.n9670 VSS.t2887 4.03583
R2467 VSS.n9718 VSS.t874 4.03583
R2468 VSS.n9719 VSS.t3247 4.03583
R2469 VSS.n9724 VSS.t848 4.03583
R2470 VSS.n569 VSS.t3547 4.03583
R2471 VSS.n571 VSS.t2857 4.03583
R2472 VSS.n574 VSS.t3153 4.03583
R2473 VSS.n10021 VSS.t2092 4.03583
R2474 VSS.n577 VSS.t1378 4.03583
R2475 VSS.n9935 VSS.t2462 4.03583
R2476 VSS.n9936 VSS.t1435 4.03583
R2477 VSS.n10009 VSS.t2118 4.03583
R2478 VSS.n9938 VSS.t971 4.03583
R2479 VSS.n10003 VSS.t1798 4.03583
R2480 VSS.n9940 VSS.t1391 4.03583
R2481 VSS.n9997 VSS.t2410 4.03583
R2482 VSS.n9942 VSS.t3351 4.03583
R2483 VSS.n9967 VSS.t1445 4.03583
R2484 VSS.n9968 VSS.t3389 4.03583
R2485 VSS.n9987 VSS.t2723 4.03583
R2486 VSS.n9970 VSS.t2296 4.03583
R2487 VSS.n9981 VSS.t3029 4.03583
R2488 VSS.n9972 VSS.t1905 4.03583
R2489 VSS.n9975 VSS.t805 4.03583
R2490 VSS.n1346 VSS.t3327 4.03583
R2491 VSS.n1371 VSS.t1623 4.03583
R2492 VSS.n1348 VSS.t2683 4.03583
R2493 VSS.n1365 VSS.t2585 4.03583
R2494 VSS.n1351 VSS.t1382 4.03583
R2495 VSS.n1359 VSS.t2697 4.03583
R2496 VSS.n1354 VSS.t1169 4.03583
R2497 VSS.n803 VSS.t2320 4.03583
R2498 VSS.n802 VSS.t1885 4.03583
R2499 VSS.n801 VSS.t1059 4.03583
R2500 VSS.n798 VSS.t2230 4.03583
R2501 VSS.n800 VSS.t3195 4.03583
R2502 VSS.n9636 VSS.t1195 4.03583
R2503 VSS.n9756 VSS.t1490 4.03583
R2504 VSS.n9638 VSS.t981 4.03583
R2505 VSS.n9662 VSS.t2176 4.03583
R2506 VSS.n9663 VSS.t1723 4.03583
R2507 VSS.n9746 VSS.t1655 4.03583
R2508 VSS.n9665 VSS.t3473 4.03583
R2509 VSS.n9740 VSS.t1733 4.03583
R2510 VSS.n9668 VSS.t2515 4.03583
R2511 VSS.n9734 VSS.t3477 4.03583
R2512 VSS.n9670 VSS.t1274 4.03583
R2513 VSS.n9718 VSS.t2414 4.03583
R2514 VSS.n9719 VSS.t900 4.03583
R2515 VSS.n9724 VSS.t2242 4.03583
R2516 VSS.n569 VSS.t3295 4.03583
R2517 VSS.n571 VSS.t3229 4.03583
R2518 VSS.n574 VSS.t2344 4.03583
R2519 VSS.n10021 VSS.t3297 4.03583
R2520 VSS.n577 VSS.t1841 4.03583
R2521 VSS.n9935 VSS.t2991 4.03583
R2522 VSS.n9936 VSS.t2517 4.03583
R2523 VSS.n10009 VSS.t727 4.03583
R2524 VSS.n9938 VSS.t1583 4.03583
R2525 VSS.n10003 VSS.t735 4.03583
R2526 VSS.n9940 VSS.t1851 4.03583
R2527 VSS.n9997 VSS.t2120 4.03583
R2528 VSS.n9942 VSS.t2424 4.03583
R2529 VSS.n9967 VSS.t3571 4.03583
R2530 VSS.n9968 VSS.t3145 4.03583
R2531 VSS.n9987 VSS.t3091 4.03583
R2532 VSS.n9970 VSS.t1022 4.03583
R2533 VSS.n9981 VSS.t2356 4.03583
R2534 VSS.n9972 VSS.t3171 4.03583
R2535 VSS.n9975 VSS.t1029 4.03583
R2536 VSS.n1316 VSS.t2979 4.03583
R2537 VSS.n1312 VSS.t598 4.03583
R2538 VSS.n1307 VSS.t2959 4.03583
R2539 VSS.n1303 VSS.t706 4.03583
R2540 VSS.n443 VSS.t1777 4.03583
R2541 VSS.n447 VSS.t1847 4.03583
R2542 VSS.n449 VSS.t1000 4.03583
R2543 VSS.n453 VSS.t1839 4.03583
R2544 VSS.n10099 VSS.t2637 4.03583
R2545 VSS.n461 VSS.t2659 4.03583
R2546 VSS.n460 VSS.t2543 4.03583
R2547 VSS.n485 VSS.t2350 4.03583
R2548 VSS.n488 VSS.t2595 4.03583
R2549 VSS.n492 VSS.t3469 4.03583
R2550 VSS.n10079 VSS.t3425 4.03583
R2551 VSS.n10075 VSS.t3451 4.03583
R2552 VSS.n501 VSS.t1199 4.03583
R2553 VSS.n519 VSS.t1228 4.03583
R2554 VSS.n522 VSS.t2228 4.03583
R2555 VSS.n528 VSS.t2310 4.03583
R2556 VSS.n515 VSS.t1532 4.03583
R2557 VSS.n539 VSS.t2360 4.03583
R2558 VSS.n541 VSS.t2599 4.03583
R2559 VSS.n545 VSS.t2272 4.03583
R2560 VSS.n551 VSS.t3109 4.03583
R2561 VSS.n554 VSS.t765 4.03583
R2562 VSS.n556 VSS.t3105 4.03583
R2563 VSS.n559 VSS.t839 4.03583
R2564 VSS.n10894 VSS.t1899 4.03583
R2565 VSS.n10890 VSS.t898 4.03583
R2566 VSS.n10876 VSS.t1161 4.03583
R2567 VSS.n10879 VSS.t1963 4.03583
R2568 VSS.n187 VSS.t2793 4.03583
R2569 VSS.n11138 VSS.t2809 4.03583
R2570 VSS.n204 VSS.t1995 4.03583
R2571 VSS.n11021 VSS.t2861 4.03583
R2572 VSS.n11024 VSS.t2737 4.03583
R2573 VSS.n11029 VSS.t3613 4.03583
R2574 VSS.n11031 VSS.t3573 4.03583
R2575 VSS.n11035 VSS.t2819 4.03583
R2576 VSS.n11114 VSS.t3621 4.03583
R2577 VSS.n11055 VSS.t456 4.03583
R2578 VSS.n11057 VSS.t1591 4.03583
R2579 VSS.n11082 VSS.t2444 4.03583
R2580 VSS.n11080 VSS.t1663 4.03583
R2581 VSS.n11088 VSS.t2477 4.03583
R2582 VSS.n11090 VSS.t2743 4.03583
R2583 VSS.n10 VSS.t1725 4.03583
R2584 VSS.n1418 VSS.t2306 4.03583
R2585 VSS.n1420 VSS.t1610 4.03583
R2586 VSS.n1466 VSS.t2280 4.03583
R2587 VSS.n1462 VSS.t1881 4.03583
R2588 VSS.n1427 VSS.t1163 4.03583
R2589 VSS.n1429 VSS.t2807 4.03583
R2590 VSS.n1439 VSS.t3489 4.03583
R2591 VSS.n1443 VSS.t2783 4.03583
R2592 VSS.n829 VSS.t769 4.03583
R2593 VSS.n9589 VSS.t2833 4.03583
R2594 VSS.n9588 VSS.t3581 4.03583
R2595 VSS.n9770 VSS.t1150 4.03583
R2596 VSS.n9776 VSS.t3181 4.03583
R2597 VSS.n9782 VSS.t2787 4.03583
R2598 VSS.n790 VSS.t710 4.03583
R2599 VSS.n787 VSS.t2755 4.03583
R2600 VSS.n9796 VSS.t750 4.03583
R2601 VSS.n772 VSS.t2811 4.03583
R2602 VSS.n9806 VSS.t2082 4.03583
R2603 VSS.n770 VSS.t547 4.03583
R2604 VSS.n9817 VSS.t1355 4.03583
R2605 VSS.n765 VSS.t3285 4.03583
R2606 VSS.n9829 VSS.t2250 4.03583
R2607 VSS.n763 VSS.t3025 4.03583
R2608 VSS.n697 VSS.t1012 4.03583
R2609 VSS.n700 VSS.t3367 4.03583
R2610 VSS.n702 VSS.t987 4.03583
R2611 VSS.n706 VSS.t519 4.03583
R2612 VSS.n726 VSS.t2995 4.03583
R2613 VSS.n728 VSS.t3275 4.03583
R2614 VSS.n740 VSS.t2224 4.03583
R2615 VSS.n736 VSS.t1522 4.03583
R2616 VSS.n158 VSS.t2619 4.03583
R2617 VSS.n11162 VSS.t1565 4.03583
R2618 VSS.n155 VSS.t2256 4.03583
R2619 VSS.n154 VSS.t1117 4.03583
R2620 VSS.n11172 VSS.t1931 4.03583
R2621 VSS.n11176 VSS.t1526 4.03583
R2622 VSS.n11178 VSS.t2545 4.03583
R2623 VSS.n11182 VSS.t3521 4.03583
R2624 VSS.n11258 VSS.t1575 4.03583
R2625 VSS.n11199 VSS.t3559 4.03583
R2626 VSS.n11201 VSS.t2871 4.03583
R2627 VSS.n11227 VSS.t2438 4.03583
R2628 VSS.n11225 VSS.t3151 4.03583
R2629 VSS.n11232 VSS.t2025 4.03583
R2630 VSS.n11234 VSS.t951 4.03583
R2631 VSS.n10394 VSS.n10393 4.02484
R2632 VSS.n10396 VSS.n10395 4.02484
R2633 VSS.n10390 VSS.n10389 4.02484
R2634 VSS.n10388 VSS.n10387 4.02484
R2635 VSS.n10404 VSS.t133 4.02247
R2636 VSS.n10402 VSS.t200 4.02247
R2637 VSS.n10299 VSS.t32 4.00471
R2638 VSS.n10294 VSS.t13 4.00471
R2639 VSS.n10118 VSS.n434 3.9853
R2640 VSS.n9564 VSS.n833 3.9853
R2641 VSS.n10067 VSS.n506 3.9853
R2642 VSS.n10929 VSS.n218 3.9853
R2643 VSS.n11361 VSS.n93 3.9853
R2644 VSS.n11468 VSS.n6 3.9853
R2645 VSS.n9197 VSS.n9191 3.98482
R2646 VSS.n9333 VSS.n9327 3.98482
R2647 VSS.n171 VSS.n165 3.98482
R2648 VSS.n9579 VSS.n9573 3.98482
R2649 VSS.n199 VSS.n193 3.98482
R2650 VSS.n477 VSS.n471 3.98482
R2651 VSS.n9030 VSS.n9024 3.98482
R2652 VSS.n270 VSS.n264 3.98482
R2653 VSS.n342 VSS.n336 3.98482
R2654 VSS.n414 VSS.n408 3.98482
R2655 VSS.n10405 VSS.n10365 3.96014
R2656 VSS.n1454 VSS.t278 3.9481
R2657 VSS.n794 VSS.t269 3.9481
R2658 VSS.n9822 VSS.t277 3.9481
R2659 VSS.n11086 VSS.t116 3.9481
R2660 VSS.n11027 VSS.t109 3.9481
R2661 VSS.n10872 VSS.t113 3.9481
R2662 VSS.n1363 VSS.t274 3.9481
R2663 VSS.n9760 VSS.t271 3.9481
R2664 VSS.n9738 VSS.t279 3.9481
R2665 VSS.n9979 VSS.t120 3.9481
R2666 VSS.n10001 VSS.t111 3.9481
R2667 VSS.n10026 VSS.t121 3.9481
R2668 VSS.n189 VSS.t159 3.93054
R2669 VSS.n194 VSS.t174 3.93054
R2670 VSS.n467 VSS.t408 3.93054
R2671 VSS.n472 VSS.t404 3.93054
R2672 VSS.n260 VSS.t302 3.93054
R2673 VSS.n265 VSS.t298 3.93054
R2674 VSS.n332 VSS.t3641 3.93054
R2675 VSS.n337 VSS.t3637 3.93054
R2676 VSS.n404 VSS.t321 3.93054
R2677 VSS.n409 VSS.t328 3.93054
R2678 VSS.n9192 VSS.t355 3.92996
R2679 VSS.n9187 VSS.t361 3.92996
R2680 VSS.n9328 VSS.t387 3.92996
R2681 VSS.n9323 VSS.t383 3.92996
R2682 VSS.n166 VSS.t373 3.92996
R2683 VSS.n161 VSS.t370 3.92996
R2684 VSS.n9574 VSS.t3633 3.92996
R2685 VSS.n9569 VSS.t446 3.92996
R2686 VSS.n9025 VSS.t3648 3.92996
R2687 VSS.n9020 VSS.t3646 3.92996
R2688 VSS.n9194 VSS.t358 3.92774
R2689 VSS.n9189 VSS.t363 3.92774
R2690 VSS.n9330 VSS.t385 3.92774
R2691 VSS.n9325 VSS.t390 3.92774
R2692 VSS.n168 VSS.t375 3.92774
R2693 VSS.n163 VSS.t372 3.92774
R2694 VSS.n9576 VSS.t3634 3.92774
R2695 VSS.n9571 VSS.t447 3.92774
R2696 VSS.n191 VSS.t197 3.92774
R2697 VSS.n196 VSS.t198 3.92774
R2698 VSS.n469 VSS.t405 3.92774
R2699 VSS.n474 VSS.t402 3.92774
R2700 VSS.n9027 VSS.t412 3.92774
R2701 VSS.n9022 VSS.t3647 3.92774
R2702 VSS.n262 VSS.t299 3.92774
R2703 VSS.n267 VSS.t295 3.92774
R2704 VSS.n334 VSS.t3642 3.92774
R2705 VSS.n339 VSS.t3638 3.92774
R2706 VSS.n406 VSS.t326 3.92774
R2707 VSS.n411 VSS.t324 3.92774
R2708 VSS.t56 VSS.n148 3.9056
R2709 VSS.n10322 VSS.t47 3.833
R2710 VSS.n10331 VSS.t124 3.833
R2711 VSS.n10320 VSS.t138 3.833
R2712 VSS.n10310 VSS.t144 3.833
R2713 VSS.n10629 VSS.t36 3.81405
R2714 VSS.n10620 VSS.t50 3.81405
R2715 VSS.n10384 VSS.t177 3.81405
R2716 VSS.n10375 VSS.t140 3.81405
R2717 VSS.n10390 VSS.n10388 3.80578
R2718 VSS.n10396 VSS.n10394 3.80578
R2719 VSS.n10319 VSS.n10315 3.80578
R2720 VSS.n10330 VSS.n10326 3.80578
R2721 VSS.n754 VSS.t110 3.78612
R2722 VSS.n156 VSS.t119 3.78612
R2723 VSS.n11204 VSS.t115 3.78612
R2724 VSS.n527 VSS.t272 3.78612
R2725 VSS.n464 VSS.t276 3.78612
R2726 VSS.n1300 VSS.t273 3.78612
R2727 VSS.n9722 VSS.t118 3.78612
R2728 VSS.n10007 VSS.t112 3.78612
R2729 VSS.n9985 VSS.t114 3.78612
R2730 VSS.n9744 VSS.t270 3.78612
R2731 VSS.n9634 VSS.t275 3.78612
R2732 VSS.n1369 VSS.t267 3.78612
R2733 VSS.n10686 VSS.n10685 3.76738
R2734 VSS.n11301 VSS.t349 3.75339
R2735 VSS.t166 VSS.t561 3.74621
R2736 VSS.n9140 VSS.t342 3.73318
R2737 VSS.n9141 VSS.t344 3.73318
R2738 VSS.n1488 VSS.t365 3.73318
R2739 VSS.n1489 VSS.t367 3.73318
R2740 VSS.n1208 VSS.t175 3.73318
R2741 VSS.n1209 VSS.t194 3.73318
R2742 VSS.n10946 VSS.t441 3.73318
R2743 VSS.n10947 VSS.t440 3.73318
R2744 VSS.n10992 VSS.t426 3.73318
R2745 VSS.n10993 VSS.t425 3.73318
R2746 VSS.n8973 VSS.t450 3.73318
R2747 VSS.n8974 VSS.t448 3.73318
R2748 VSS.n978 VSS.t313 3.73318
R2749 VSS.n979 VSS.t316 3.73318
R2750 VSS.n1036 VSS.t346 3.73318
R2751 VSS.n1037 VSS.t348 3.73318
R2752 VSS.n1085 VSS.t3649 3.73318
R2753 VSS.n1086 VSS.t170 3.73318
R2754 VSS.n871 VSS.t418 3.73318
R2755 VSS.n872 VSS.t417 3.73318
R2756 VSS.n10601 VSS.t184 3.72778
R2757 VSS.n9140 VSS.t343 3.4916
R2758 VSS.n9141 VSS.t341 3.4916
R2759 VSS.n1488 VSS.t366 3.4916
R2760 VSS.n1489 VSS.t364 3.4916
R2761 VSS.n1208 VSS.t391 3.4916
R2762 VSS.n1209 VSS.t290 3.4916
R2763 VSS.n10946 VSS.t443 3.4916
R2764 VSS.n10947 VSS.t442 3.4916
R2765 VSS.n10992 VSS.t428 3.4916
R2766 VSS.n10993 VSS.t427 3.4916
R2767 VSS.n8973 VSS.t451 3.4916
R2768 VSS.n8974 VSS.t449 3.4916
R2769 VSS.n978 VSS.t315 3.4916
R2770 VSS.n979 VSS.t314 3.4916
R2771 VSS.n1036 VSS.t347 3.4916
R2772 VSS.n1037 VSS.t345 3.4916
R2773 VSS.n1085 VSS.t173 3.4916
R2774 VSS.n1086 VSS.t180 3.4916
R2775 VSS.n871 VSS.t420 3.4916
R2776 VSS.n872 VSS.t419 3.4916
R2777 VSS.t1801 VSS.n10840 3.40963
R2778 VSS.n10638 VSS.t1976 3.37683
R2779 VSS.n11324 VSS.t2211 3.36554
R2780 VSS.n10823 VSS.t1710 3.3605
R2781 VSS.t1710 VSS.n10821 3.3605
R2782 VSS.n10823 VSS.t3480 3.3605
R2783 VSS.t3480 VSS.n10821 3.3605
R2784 VSS.n10841 VSS.t1801 3.3605
R2785 VSS.n10843 VSS.t2790 3.3605
R2786 VSS.t2790 VSS.n10842 3.3605
R2787 VSS.n10712 VSS.t351 3.3605
R2788 VSS.n10713 VSS.t350 3.3605
R2789 VSS.t1429 VSS.n127 3.3605
R2790 VSS.n9205 VSS.t627 3.3605
R2791 VSS.n9183 VSS.t2726 3.3605
R2792 VSS.t3304 VSS.n1523 3.3605
R2793 VSS.n9061 VSS.t2275 3.3605
R2794 VSS.t3510 VSS.n1527 3.3605
R2795 VSS.n1546 VSS.t1511 3.3605
R2796 VSS.n1548 VSS.t1774 3.3605
R2797 VSS.n1552 VSS.t1015 3.3605
R2798 VSS.n9170 VSS.t3102 3.3605
R2799 VSS.n9174 VSS.t2016 3.3605
R2800 VSS.n9136 VSS.t2634 3.3605
R2801 VSS.n9132 VSS.t1605 3.3605
R2802 VSS.n9256 VSS.t862 3.3605
R2803 VSS.n9252 VSS.t2942 3.3605
R2804 VSS.t1712 VSS.n1513 3.3605
R2805 VSS.n9146 VSS.t2397 3.3605
R2806 VSS.n9241 VSS.t1618 3.3605
R2807 VSS.n9245 VSS.t3620 3.3605
R2808 VSS.n9211 VSS.t2385 3.3605
R2809 VSS.n9207 VSS.t3126 3.3605
R2810 VSS.n9314 VSS.t2041 3.3605
R2811 VSS.n9310 VSS.t968 3.3605
R2812 VSS.t1630 VSS.n1505 3.3605
R2813 VSS.n9217 VSS.t2313 3.3605
R2814 VSS.n9292 VSS.t1369 3.3605
R2815 VSS.n9296 VSS.t3344 3.3605
R2816 VSS.n9262 VSS.t880 3.3605
R2817 VSS.n9258 VSS.t1634 3.3605
R2818 VSS.n9354 VSS.t2852 3.3605
R2819 VSS.n9350 VSS.t2137 3.3605
R2820 VSS.t1377 VSS.n1496 3.3605
R2821 VSS.n9268 VSS.t2401 3.3605
R2822 VSS.t3534 VSS.n1478 3.3605
R2823 VSS.n9343 VSS.t2848 3.3605
R2824 VSS.n9320 VSS.t2049 3.3605
R2825 VSS.n9316 VSS.t3132 3.3605
R2826 VSS.n9387 VSS.t2598 3.3605
R2827 VSS.n9383 VSS.t470 3.3605
R2828 VSS.n9380 VSS.t2181 3.3605
R2829 VSS.n9376 VSS.t3214 3.3605
R2830 VSS.n9415 VSS.t1910 3.3605
R2831 VSS.n9419 VSS.t2982 3.3605
R2832 VSS.t1489 VSS.n1396 3.3605
R2833 VSS.n1494 VSS.t2512 3.3605
R2834 VSS.n9534 VSS.t1090 3.3605
R2835 VSS.n9530 VSS.t2179 3.3605
R2836 VSS.t1416 VSS.n1221 3.3605
R2837 VSS.n1402 VSS.t621 3.3605
R2838 VSS.n11236 VSS.t952 3.3605
R2839 VSS.n11242 VSS.t2026 3.3605
R2840 VSS.n11230 VSS.t3152 3.3605
R2841 VSS.n11248 VSS.t2439 3.3605
R2842 VSS.n11203 VSS.t2872 3.3605
R2843 VSS.n11254 VSS.t3560 3.3605
R2844 VSS.n11256 VSS.t1576 3.3605
R2845 VSS.t1576 VSS.n11197 3.3605
R2846 VSS.n11262 VSS.t3522 3.3605
R2847 VSS.t3522 VSS.n11180 3.3605
R2848 VSS.t2546 VSS.n11268 3.3605
R2849 VSS.t1527 VSS.n11174 3.3605
R2850 VSS.t1932 VSS.n11274 3.3605
R2851 VSS.t1118 VSS.n11171 3.3605
R2852 VSS.n11167 VSS.t2257 3.3605
R2853 VSS.n173 VSS.t1566 3.3605
R2854 VSS.n11158 VSS.t2620 3.3605
R2855 VSS.t2620 VSS.n11157 3.3605
R2856 VSS.n734 VSS.t1523 3.3605
R2857 VSS.t1523 VSS.n732 3.3605
R2858 VSS.n730 VSS.t2225 3.3605
R2859 VSS.n745 VSS.t3276 3.3605
R2860 VSS.t2996 VSS.n747 3.3605
R2861 VSS.t520 VSS.n704 3.3605
R2862 VSS.t988 VSS.n755 3.3605
R2863 VSS.t3368 VSS.n696 3.3605
R2864 VSS.t1013 VSS.n761 3.3605
R2865 VSS.n762 VSS.t1013 3.3605
R2866 VSS.n9837 VSS.t3026 3.3605
R2867 VSS.t3026 VSS.n9836 3.3605
R2868 VSS.n9833 VSS.t2251 3.3605
R2869 VSS.n9825 VSS.t3286 3.3605
R2870 VSS.n9821 VSS.t1356 3.3605
R2871 VSS.n9812 VSS.t548 3.3605
R2872 VSS.n9810 VSS.t2083 3.3605
R2873 VSS.n9802 VSS.t2812 3.3605
R2874 VSS.n9799 VSS.t751 3.3605
R2875 VSS.t751 VSS.n9798 3.3605
R2876 VSS.n9792 VSS.t2756 3.3605
R2877 VSS.t2756 VSS.n9791 3.3605
R2878 VSS.n9787 VSS.t711 3.3605
R2879 VSS.n9780 VSS.t2788 3.3605
R2880 VSS.n9774 VSS.t3182 3.3605
R2881 VSS.t1151 VSS.n9772 3.3605
R2882 VSS.n9581 VSS.t3582 3.3605
R2883 VSS.n9595 VSS.t2834 3.3605
R2884 VSS.t770 VSS.n9598 3.3605
R2885 VSS.n9599 VSS.t770 3.3605
R2886 VSS.t2784 VSS.n1445 3.3605
R2887 VSS.n1446 VSS.t2784 3.3605
R2888 VSS.n1441 VSS.t3490 3.3605
R2889 VSS.n1452 VSS.t2808 3.3605
R2890 VSS.n1458 VSS.t1164 3.3605
R2891 VSS.t1882 VSS.n1425 3.3605
R2892 VSS.n1423 VSS.t2281 3.3605
R2893 VSS.n1470 VSS.t1611 3.3605
R2894 VSS.n1472 VSS.t2307 3.3605
R2895 VSS.t2307 VSS.n1403 3.3605
R2896 VSS.t3202 VSS.n11237 3.3605
R2897 VSS.t802 VSS.n11231 3.3605
R2898 VSS.t1456 VSS.n11243 3.3605
R2899 VSS.t3438 VSS.n11228 3.3605
R2900 VSS.t1898 VSS.n11249 3.3605
R2901 VSS.t2964 VSS.n11198 3.3605
R2902 VSS.n11255 VSS.t3190 3.3605
R2903 VSS.n11261 VSS.t2149 3.3605
R2904 VSS.t2764 VSS.n11265 3.3605
R2905 VSS.t3448 VSS.n11177 3.3605
R2906 VSS.t3308 VSS.n11271 3.3605
R2907 VSS.t940 VSS.n152 3.3605
R2908 VSS.n11170 VSS.t3048 3.3605
R2909 VSS.n11163 VSS.t592 3.3605
R2910 VSS.n11161 VSS.t2289 3.3605
R2911 VSS.n11155 VSS.t1251 3.3605
R2912 VSS.n733 VSS.t1868 3.3605
R2913 VSS.n739 VSS.t768 3.3605
R2914 VSS.n742 VSS.t2105 3.3605
R2915 VSS.n747 VSS.t3158 3.3605
R2916 VSS.t1352 VSS.n751 3.3605
R2917 VSS.t2034 VSS.n701 3.3605
R2918 VSS.t3596 VSS.n758 3.3605
R2919 VSS.t1607 VSS.n698 3.3605
R2920 VSS.n9840 VSS.t1862 3.3605
R2921 VSS.n9834 VSS.t1124 3.3605
R2922 VSS.t516 VSS.n764 3.3605
R2923 VSS.t1680 VSS.n9826 3.3605
R2924 VSS.t2133 VSS.n769 3.3605
R2925 VSS.t1054 VSS.n9813 3.3605
R2926 VSS.t2359 VSS.n771 3.3605
R2927 VSS.t3382 VSS.n9803 3.3605
R2928 VSS.t3018 VSS.n773 3.3605
R2929 VSS.t1944 VSS.n9793 3.3605
R2930 VSS.n9790 VSS.t3226 3.3605
R2931 VSS.n9783 VSS.t1210 3.3605
R2932 VSS.n9779 VSS.t2722 3.3605
R2933 VSS.n9771 VSS.t2002 3.3605
R2934 VSS.t2261 VSS.n796 3.3605
R2935 VSS.t1503 VSS.n9590 3.3605
R2936 VSS.n9597 VSS.t1770 3.3605
R2937 VSS.t1007 VSS.n827 3.3605
R2938 VSS.n1444 VSS.t2323 3.3605
R2939 VSS.n1449 VSS.t3358 3.3605
R2940 VSS.n1428 VSS.t1227 3.3605
R2941 VSS.n1461 VSS.t3588 3.3605
R2942 VSS.t1813 VSS.n1463 3.3605
R2943 VSS.t2880 VSS.n1422 3.3605
R2944 VSS.n1419 VSS.t2091 3.3605
R2945 VSS.n1475 VSS.t1412 3.3605
R2946 VSS.n9547 VSS.t1572 3.3605
R2947 VSS.n9543 VSS.t738 3.3605
R2948 VSS.n9540 VSS.t1017 3.3605
R2949 VSS.n9536 VSS.t3386 3.3605
R2950 VSS.n1200 VSS.t1682 3.3605
R2951 VSS.n1204 VSS.t2728 3.3605
R2952 VSS.n1206 VSS.t2287 3.3605
R2953 VSS.n1214 VSS.t1247 3.3605
R2954 VSS.n10936 VSS.t2928 3.3605
R2955 VSS.n10932 VSS.t847 3.3605
R2956 VSS.t1135 VSS.n214 3.3605
R2957 VSS.n1168 VSS.t3526 3.3605
R2958 VSS.n10975 VSS.t1622 3.3605
R2959 VSS.n10979 VSS.t3624 3.3605
R2960 VSS.n10942 VSS.t1145 3.3605
R2961 VSS.n10938 VSS.t3178 3.3605
R2962 VSS.n11368 VSS.t2473 3.3605
R2963 VSS.n11364 VSS.t1464 3.3605
R2964 VSS.t2051 VSS.n90 3.3605
R2965 VSS.n10952 VSS.t2778 3.3605
R2966 VSS.n11381 VSS.t2968 3.3605
R2967 VSS.n11377 VSS.t1902 3.3605
R2968 VSS.n11374 VSS.t2494 3.3605
R2969 VSS.n11370 VSS.t3210 3.3605
R2970 VSS.t1974 VSS.n13 3.3605
R2971 VSS.n11461 VSS.t1460 3.3605
R2972 VSS.n11465 VSS.t1493 3.3605
R2973 VSS.t1714 VSS.n11093 3.3605
R2974 VSS.t625 VSS.n11087 3.3605
R2975 VSS.t2886 VSS.n11099 3.3605
R2976 VSS.t2914 VSS.n11083 3.3605
R2977 VSS.t1320 VSS.n11105 3.3605
R2978 VSS.t1044 VSS.n11054 3.3605
R2979 VSS.n11111 VSS.t2457 3.3605
R2980 VSS.n11117 VSS.t2482 3.3605
R2981 VSS.n11036 VSS.t2740 3.3605
R2982 VSS.n11122 VSS.t1746 3.3605
R2983 VSS.n11030 VSS.t2668 3.3605
R2984 VSS.n11128 VSS.t1672 3.3605
R2985 VSS.n205 VSS.t2303 3.3605
R2986 VSS.n11137 VSS.t1299 3.3605
R2987 VSS.n11139 VSS.t1184 3.3605
R2988 VSS.n11149 VSS.t1235 3.3605
R2989 VSS.n10882 VSS.t1485 3.3605
R2990 VSS.t1513 VSS.n10877 3.3605
R2991 VSS.n10875 VSS.t532 3.3605
R2992 VSS.n10893 VSS.t3430 3.3605
R2993 VSS.t1398 VSS.n10035 3.3605
R2994 VSS.t3406 VSS.n555 3.3605
R2995 VSS.t2822 VSS.n10042 3.3605
R2996 VSS.t2556 VSS.n552 3.3605
R2997 VSS.n10047 VSS.t2020 3.3605
R2998 VSS.n10053 VSS.t2850 3.3605
R2999 VSS.n542 VSS.t2295 3.3605
R3000 VSS.n10059 VSS.t2057 3.3605
R3001 VSS.n533 VSS.t2754 3.3605
R3002 VSS.t2802 VSS.n531 3.3605
R3003 VSS.t1916 VSS.n516 3.3605
R3004 VSS.t1684 VSS.n503 3.3605
R3005 VSS.n502 VSS.t1080 3.3605
R3006 VSS.n10074 VSS.t1109 3.3605
R3007 VSS.t3302 VSS.n10076 3.3605
R3008 VSS.t3112 VSS.n493 3.3605
R3009 VSS.t3398 VSS.n10084 3.3605
R3010 VSS.t1143 VSS.n484 3.3605
R3011 VSS.t2548 VSS.n10090 3.3605
R3012 VSS.t2672 VSS.n462 3.3605
R3013 VSS.n10096 VSS.t2135 3.3605
R3014 VSS.n10102 VSS.t2950 3.3605
R3015 VSS.n454 VSS.t2047 3.3605
R3016 VSS.n10107 VSS.t1830 3.3605
R3017 VSS.n446 VSS.t2032 3.3605
R3018 VSS.t2864 VSS.n441 3.3605
R3019 VSS.t1972 VSS.n1304 3.3605
R3020 VSS.t1748 VSS.n1298 3.3605
R3021 VSS.t3456 VSS.n1313 3.3605
R3022 VSS.t1186 VSS.n1296 3.3605
R3023 VSS.n12 VSS.t1726 3.3605
R3024 VSS.t1726 VSS.n9 3.3605
R3025 VSS.n11092 VSS.t2744 3.3605
R3026 VSS.n11098 VSS.t2478 3.3605
R3027 VSS.n11085 VSS.t1664 3.3605
R3028 VSS.n11104 VSS.t2445 3.3605
R3029 VSS.n11059 VSS.t1592 3.3605
R3030 VSS.n11110 VSS.t457 3.3605
R3031 VSS.n11112 VSS.t3622 3.3605
R3032 VSS.t3622 VSS.n11053 3.3605
R3033 VSS.t2820 VSS.n11118 3.3605
R3034 VSS.n11119 VSS.t2820 3.3605
R3035 VSS.n11033 VSS.t3574 3.3605
R3036 VSS.n11125 VSS.t3614 3.3605
R3037 VSS.n11026 VSS.t2738 3.3605
R3038 VSS.n11131 VSS.t2862 3.3605
R3039 VSS.n11134 VSS.t1996 3.3605
R3040 VSS.t2810 VSS.n201 3.3605
R3041 VSS.n11146 VSS.t2794 3.3605
R3042 VSS.t2794 VSS.n185 3.3605
R3043 VSS.t1964 VSS.n10883 3.3605
R3044 VSS.n10884 VSS.t1964 3.3605
R3045 VSS.t1162 VSS.n10886 3.3605
R3046 VSS.t899 VSS.n10874 3.3605
R3047 VSS.n10893 VSS.t1900 3.3605
R3048 VSS.t840 VSS.n10870 3.3605
R3049 VSS.t3106 VSS.n10039 3.3605
R3050 VSS.t766 VSS.n550 3.3605
R3051 VSS.t3110 VSS.n10045 3.3605
R3052 VSS.n10046 VSS.t3110 3.3605
R3053 VSS.n10050 VSS.t2273 3.3605
R3054 VSS.t2273 VSS.n543 3.3605
R3055 VSS.t2600 VSS.n10054 3.3605
R3056 VSS.t2361 VSS.n537 3.3605
R3057 VSS.t1533 VSS.n10061 3.3605
R3058 VSS.n530 VSS.t2311 3.3605
R3059 VSS.n526 VSS.t2229 3.3605
R3060 VSS.n517 VSS.t1229 3.3605
R3061 VSS.t1200 VSS.n10070 3.3605
R3062 VSS.n10071 VSS.t1200 3.3605
R3063 VSS.n497 VSS.t3452 3.3605
R3064 VSS.t3452 VSS.n496 3.3605
R3065 VSS.n494 VSS.t3426 3.3605
R3066 VSS.n10083 VSS.t3470 3.3605
R3067 VSS.n490 VSS.t2596 3.3605
R3068 VSS.n10089 VSS.t2351 3.3605
R3069 VSS.n465 VSS.t2544 3.3605
R3070 VSS.n10095 VSS.t2660 3.3605
R3071 VSS.n10097 VSS.t2638 3.3605
R3072 VSS.t2638 VSS.n457 3.3605
R3073 VSS.t1840 VSS.n10103 3.3605
R3074 VSS.n10104 VSS.t1840 3.3605
R3075 VSS.n451 VSS.t1001 3.3605
R3076 VSS.n10110 VSS.t1848 3.3605
R3077 VSS.t1778 VSS.n10112 3.3605
R3078 VSS.n1302 VSS.t707 3.3605
R3079 VSS.n1299 VSS.t2960 3.3605
R3080 VSS.n1311 VSS.t599 3.3605
R3081 VSS.n1273 VSS.t2980 3.3605
R3082 VSS.t2980 VSS.n1272 3.3605
R3083 VSS.n11341 VSS.t2371 3.3605
R3084 VSS.n11345 VSS.t2403 3.3605
R3085 VSS.n11348 VSS.t2650 3.3605
R3086 VSS.n11352 VSS.t1658 3.3605
R3087 VSS.n11354 VSS.t3378 3.3605
R3088 VSS.n11358 VSS.t3420 3.3605
R3089 VSS.t514 VSS.n96 3.3605
R3090 VSS.n10998 VSS.t2678 3.3605
R3091 VSS.n10989 VSS.t2147 3.3605
R3092 VSS.n10985 VSS.t2183 3.3605
R3093 VSS.t2391 VSS.n207 3.3605
R3094 VSS.n10920 VSS.t2423 3.3605
R3095 VSS.n10637 VSS.t1371 3.3605
R3096 VSS.t1371 VSS.n10636 3.3605
R3097 VSS.n10637 VSS.t1105 3.3605
R3098 VSS.n10636 VSS.t1105 3.3605
R3099 VSS.n10637 VSS.t3486 3.3605
R3100 VSS.n10636 VSS.t3486 3.3605
R3101 VSS.t1976 VSS.n10634 3.3605
R3102 VSS.t786 VSS.n10642 3.3605
R3103 VSS.n10648 VSS.t1648 3.3605
R3104 VSS.n10649 VSS.t2393 3.3605
R3105 VSS.t526 VSS.n10347 3.3605
R3106 VSS.n10511 VSS.t526 3.3605
R3107 VSS.n10513 VSS.t656 3.3605
R3108 VSS.t2924 VSS.n10504 3.3605
R3109 VSS.t2283 VSS.n10525 3.3605
R3110 VSS.t3170 VSS.n10489 3.3605
R3111 VSS.n10540 VSS.t3590 3.3605
R3112 VSS.t1688 VSS.n10483 3.3605
R3113 VSS.n10552 VSS.t2836 3.3605
R3114 VSS.t2836 VSS.n10482 3.3605
R3115 VSS.n10512 VSS.t1166 3.3605
R3116 VSS.n10515 VSS.t873 3.3605
R3117 VSS.n10524 VSS.t2750 3.3605
R3118 VSS.n10503 VSS.t1892 3.3605
R3119 VSS.t1892 VSS.n10498 3.3605
R3120 VSS.t700 VSS.n10538 3.3605
R3121 VSS.n10539 VSS.t700 3.3605
R3122 VSS.n10542 VSS.t1888 3.3605
R3123 VSS.n10551 VSS.t3056 3.3605
R3124 VSS.n10589 VSS.t1141 3.3605
R3125 VSS.n10438 VSS.t1469 3.3605
R3126 VSS.t2576 VSS.n10432 3.3605
R3127 VSS.n10431 VSS.t658 3.3605
R3128 VSS.t2926 VSS.n10424 3.3605
R3129 VSS.n10423 VSS.t2285 3.3605
R3130 VSS.t1434 VSS.n10291 3.3605
R3131 VSS.t1139 VSS.n10454 3.3605
R3132 VSS.n10460 VSS.t3310 3.3605
R3133 VSS.t2732 VSS.n10461 3.3605
R3134 VSS.n10468 VSS.t3600 3.3605
R3135 VSS.t921 VSS.n10469 3.3605
R3136 VSS.n10475 VSS.t2113 3.3605
R3137 VSS.t3312 VSS.n10582 3.3605
R3138 VSS.n10581 VSS.t2734 3.3605
R3139 VSS.t1854 VSS.n10575 3.3605
R3140 VSS.n9038 VSS.t2874 3.3605
R3141 VSS.n9016 VSS.t798 3.3605
R3142 VSS.t1082 VSS.n1561 3.3605
R3143 VSS.n1570 VSS.t3464 3.3605
R3144 VSS.n9003 VSS.t2171 3.3605
R3145 VSS.n9007 VSS.t3206 3.3605
R3146 VSS.n8969 VSS.t3472 3.3605
R3147 VSS.n8965 VSS.t2796 3.3605
R3148 VSS.n9099 VSS.t986 3.3605
R3149 VSS.n9095 VSS.t2067 3.3605
R3150 VSS.t1666 VSS.n1554 3.3605
R3151 VSS.n8979 VSS.t493 3.3605
R3152 VSS.n9084 VSS.t1736 3.3605
R3153 VSS.n9088 VSS.t2792 3.3605
R3154 VSS.n9044 VSS.t2337 3.3605
R3155 VSS.n9040 VSS.t1297 3.3605
R3156 VSS.n9063 VSS.t1102 3.3605
R3157 VSS.n9067 VSS.t2195 3.3605
R3158 VSS.n9069 VSS.t2447 3.3605
R3159 VSS.n9073 VSS.t1768 3.3605
R3160 VSS.n974 VSS.t2155 3.3605
R3161 VSS.n970 VSS.t1914 3.3605
R3162 VSS.n968 VSS.t1390 3.3605
R3163 VSS.n964 VSS.t2185 3.3605
R3164 VSS.n10262 VSS.t1194 3.3605
R3165 VSS.n10271 VSS.t917 3.3605
R3166 VSS.n10273 VSS.t3492 3.3605
R3167 VSS.n10277 VSS.t1240 3.3605
R3168 VSS.n312 VSS.t3266 3.3605
R3169 VSS.n308 VSS.t3068 3.3605
R3170 VSS.n306 VSS.t2459 3.3605
R3171 VSS.t2488 VSS.n272 3.3605
R3172 VSS.n990 VSS.t1116 3.3605
R3173 VSS.n986 VSS.t871 3.3605
R3174 VSS.n984 VSS.t3380 3.3605
R3175 VSS.n976 VSS.t3422 3.3605
R3176 VSS.n1011 VSS.t2373 3.3605
R3177 VSS.n1007 VSS.t2163 3.3605
R3178 VSS.n1005 VSS.t1632 3.3605
R3179 VSS.n1001 VSS.t2405 3.3605
R3180 VSS.n10223 VSS.t1473 3.3605
R3181 VSS.n10219 VSS.t1204 3.3605
R3182 VSS.n318 VSS.t594 3.3605
R3183 VSS.n314 VSS.t1495 3.3605
R3184 VSS.n10202 VSS.t3168 3.3605
R3185 VSS.n10211 VSS.t3194 3.3605
R3186 VSS.n10213 VSS.t3400 3.3605
R3187 VSS.n10217 VSS.t3444 3.3605
R3188 VSS.n1023 VSS.t999 3.3605
R3189 VSS.n1019 VSS.t1038 3.3605
R3190 VSS.n1017 VSS.t1304 3.3605
R3191 VSS.n1013 VSS.t1344 3.3605
R3192 VSS.n1048 VSS.t2305 3.3605
R3193 VSS.n1044 VSS.t2333 3.3605
R3194 VSS.n1042 VSS.t2946 3.3605
R3195 VSS.n1034 VSS.t1926 3.3605
R3196 VSS.n375 VSS.t1388 3.3605
R3197 VSS.n371 VSS.t1422 3.3605
R3198 VSS.n369 VSS.t1984 3.3605
R3199 VSS.t933 VSS.n344 3.3605
R3200 VSS.n10163 VSS.t3374 3.3605
R3201 VSS.n10159 VSS.t3414 3.3605
R3202 VSS.n390 VSS.t504 3.3605
R3203 VSS.n386 VSS.t2670 3.3605
R3204 VSS.n1060 VSS.t1279 3.3605
R3205 VSS.n1056 VSS.t1324 3.3605
R3206 VSS.n1054 VSS.t1564 3.3605
R3207 VSS.n1050 VSS.t3606 3.3605
R3208 VSS.n1081 VSS.t2674 3.3605
R3209 VSS.n1077 VSS.t3460 3.3605
R3210 VSS.n1075 VSS.t2143 3.3605
R3211 VSS.n1071 VSS.t1904 3.3605
R3212 VSS.n10142 VSS.t1742 3.3605
R3213 VSS.n10151 VSS.t2522 3.3605
R3214 VSS.n10153 VSS.t1182 3.3605
R3215 VSS.n10157 VSS.t913 3.3605
R3216 VSS.n1294 VSS.t3316 3.3605
R3217 VSS.n1290 VSS.t3124 3.3605
R3218 VSS.n1288 VSS.t3612 3.3605
R3219 VSS.t3348 VSS.n416 3.3605
R3220 VSS.n1097 VSS.t1218 3.3605
R3221 VSS.n1093 VSS.t950 3.3605
R3222 VSS.n1091 VSS.t1507 3.3605
R3223 VSS.n1083 VSS.t1249 3.3605
R3224 VSS.n1118 VSS.t2932 3.3605
R3225 VSS.n1114 VSS.t2686 3.3605
R3226 VSS.n1112 VSS.t1358 3.3605
R3227 VSS.n1108 VSS.t2151 3.3605
R3228 VSS.n1130 VSS.t3504 3.3605
R3229 VSS.n1126 VSS.t3610 3.3605
R3230 VSS.n1124 VSS.t3104 3.3605
R3231 VSS.n1120 VSS.t755 3.3605
R3232 VSS.n862 VSS.t2868 3.3605
R3233 VSS.n866 VSS.t2606 3.3605
R3234 VSS.n869 VSS.t2045 3.3605
R3235 VSS.n877 VSS.t2073 3.3605
R3236 VSS.n10922 VSS.t607 3.3605
R3237 VSS.n10926 VSS.t3512 3.3605
R3238 VSS.t2990 VSS.n221 3.3605
R3239 VSS.n842 VSS.t631 3.3605
R3240 VSS.n10364 VSS.t3446 3.3605
R3241 VSS.t1176 VSS.n10358 3.3605
R3242 VSS.n10357 VSS.t1968 3.3605
R3243 VSS.n10669 VSS.t679 3.3605
R3244 VSS.t3536 VSS.n10670 3.3605
R3245 VSS.n10676 VSS.t2301 3.3605
R3246 VSS.n9473 VSS.t1402 3.3605
R3247 VSS.n9469 VSS.t3008 3.3605
R3248 VSS.t3514 VSS.n1380 3.3605
R3249 VSS.n9433 VSS.t2037 3.3605
R3250 VSS.n9461 VSS.t434 3.3605
R3251 VSS.n9461 VSS.t437 3.3605
R3252 VSS.n9460 VSS.t438 3.3605
R3253 VSS.n9460 VSS.t431 3.3605
R3254 VSS.n9459 VSS.t435 3.3605
R3255 VSS.n9459 VSS.t432 3.3605
R3256 VSS.n1379 VSS.t439 3.3605
R3257 VSS.n1379 VSS.t436 3.3605
R3258 VSS.n9454 VSS.t1238 3.3605
R3259 VSS.n9458 VSS.t2476 3.3605
R3260 VSS.n9452 VSS.t1795 3.3605
R3261 VSS.n9448 VSS.t3086 3.3605
R3262 VSS.n9974 VSS.t1030 3.3605
R3263 VSS.n9978 VSS.t3172 3.3605
R3264 VSS.n9980 VSS.t2357 3.3605
R3265 VSS.n9984 VSS.t1023 3.3605
R3266 VSS.n9986 VSS.t3092 3.3605
R3267 VSS.n9990 VSS.t3146 3.3605
R3268 VSS.t3572 VSS.n9991 3.3605
R3269 VSS.n9992 VSS.t3572 3.3605
R3270 VSS.t2425 VSS.n9994 3.3605
R3271 VSS.n9995 VSS.t2425 3.3605
R3272 VSS.n9996 VSS.t2121 3.3605
R3273 VSS.n10000 VSS.t1852 3.3605
R3274 VSS.n10002 VSS.t736 3.3605
R3275 VSS.n10006 VSS.t1584 3.3605
R3276 VSS.n10008 VSS.t728 3.3605
R3277 VSS.n10012 VSS.t2518 3.3605
R3278 VSS.t2992 VSS.n10013 3.3605
R3279 VSS.n10014 VSS.t2992 3.3605
R3280 VSS.t1842 VSS.n10016 3.3605
R3281 VSS.n10017 VSS.t1842 3.3605
R3282 VSS.n10019 VSS.t3298 3.3605
R3283 VSS.n10024 VSS.t2345 3.3605
R3284 VSS.t3230 VSS.n10027 3.3605
R3285 VSS.n9721 VSS.t3296 3.3605
R3286 VSS.n9723 VSS.t2243 3.3605
R3287 VSS.n9727 VSS.t901 3.3605
R3288 VSS.t2415 VSS.n9728 3.3605
R3289 VSS.n9729 VSS.t2415 3.3605
R3290 VSS.t1275 VSS.n9731 3.3605
R3291 VSS.n9732 VSS.t1275 3.3605
R3292 VSS.n9733 VSS.t3478 3.3605
R3293 VSS.n9737 VSS.t2516 3.3605
R3294 VSS.n9739 VSS.t1734 3.3605
R3295 VSS.n9743 VSS.t3474 3.3605
R3296 VSS.n9745 VSS.t1656 3.3605
R3297 VSS.n9749 VSS.t1724 3.3605
R3298 VSS.t2177 VSS.n9750 3.3605
R3299 VSS.n9751 VSS.t2177 3.3605
R3300 VSS.t982 VSS.n9753 3.3605
R3301 VSS.n9754 VSS.t982 3.3605
R3302 VSS.n9755 VSS.t1491 3.3605
R3303 VSS.n9759 VSS.t1196 3.3605
R3304 VSS.t3196 VSS.n9761 3.3605
R3305 VSS.t2231 VSS.n9635 3.3605
R3306 VSS.n9633 VSS.t1060 3.3605
R3307 VSS.n9629 VSS.t1886 3.3605
R3308 VSS.n9628 VSS.t2321 3.3605
R3309 VSS.t2321 VSS.n9627 3.3605
R3310 VSS.t1170 VSS.n805 3.3605
R3311 VSS.n1355 VSS.t1170 3.3605
R3312 VSS.n1357 VSS.t2698 3.3605
R3313 VSS.n1362 VSS.t1383 3.3605
R3314 VSS.n1364 VSS.t2586 3.3605
R3315 VSS.n1368 VSS.t2684 3.3605
R3316 VSS.n1370 VSS.t1624 3.3605
R3317 VSS.n1374 VSS.t3328 3.3605
R3318 VSS.n9974 VSS.t806 3.3605
R3319 VSS.n9978 VSS.t1906 3.3605
R3320 VSS.n9980 VSS.t3030 3.3605
R3321 VSS.n9984 VSS.t2297 3.3605
R3322 VSS.n9986 VSS.t2724 3.3605
R3323 VSS.n9990 VSS.t3390 3.3605
R3324 VSS.n9991 VSS.t1446 3.3605
R3325 VSS.n9992 VSS.t1446 3.3605
R3326 VSS.n9994 VSS.t3352 3.3605
R3327 VSS.n9995 VSS.t3352 3.3605
R3328 VSS.n9996 VSS.t2411 3.3605
R3329 VSS.n10000 VSS.t1392 3.3605
R3330 VSS.n10002 VSS.t1799 3.3605
R3331 VSS.n10006 VSS.t972 3.3605
R3332 VSS.n10008 VSS.t2119 3.3605
R3333 VSS.n10012 VSS.t1436 3.3605
R3334 VSS.n10013 VSS.t2463 3.3605
R3335 VSS.n10014 VSS.t2463 3.3605
R3336 VSS.n10016 VSS.t1379 3.3605
R3337 VSS.n10017 VSS.t1379 3.3605
R3338 VSS.n10019 VSS.t2093 3.3605
R3339 VSS.n10024 VSS.t3154 3.3605
R3340 VSS.n10027 VSS.t2858 3.3605
R3341 VSS.n9721 VSS.t3548 3.3605
R3342 VSS.n9723 VSS.t849 3.3605
R3343 VSS.n9727 VSS.t3248 3.3605
R3344 VSS.n9728 VSS.t875 3.3605
R3345 VSS.n9729 VSS.t875 3.3605
R3346 VSS.n9731 VSS.t2888 3.3605
R3347 VSS.n9732 VSS.t2888 3.3605
R3348 VSS.n9733 VSS.t2115 3.3605
R3349 VSS.n9737 VSS.t3166 3.3605
R3350 VSS.n9739 VSS.t1188 3.3605
R3351 VSS.n9743 VSS.t3564 3.3605
R3352 VSS.n9745 VSS.t1952 3.3605
R3353 VSS.n9749 VSS.t2656 3.3605
R3354 VSS.n9750 VSS.t586 3.3605
R3355 VSS.n9751 VSS.t586 3.3605
R3356 VSS.n9753 VSS.t2614 3.3605
R3357 VSS.n9754 VSS.t2614 3.3605
R3358 VSS.n9755 VSS.t518 3.3605
R3359 VSS.n9759 VSS.t2630 3.3605
R3360 VSS.n9761 VSS.t3080 3.3605
R3361 VSS.n9635 VSS.t992 3.3605
R3362 VSS.n9633 VSS.t3428 3.3605
R3363 VSS.t2688 VSS.n9629 3.3605
R3364 VSS.n9628 VSS.t602 3.3605
R3365 VSS.n9627 VSS.t602 3.3605
R3366 VSS.t2624 VSS.n805 3.3605
R3367 VSS.n1355 VSS.t2624 3.3605
R3368 VSS.n1357 VSS.t3326 3.3605
R3369 VSS.n1362 VSS.t2654 3.3605
R3370 VSS.n1364 VSS.t996 3.3605
R3371 VSS.n1368 VSS.t1762 3.3605
R3372 VSS.n1370 VSS.t2167 3.3605
R3373 VSS.n1374 VSS.t1479 3.3605
R3374 VSS.n10822 VSS.t1429 3.3605
R3375 VSS.n9197 VSS.n9196 3.27473
R3376 VSS.n9333 VSS.n9332 3.27473
R3377 VSS.n171 VSS.n170 3.27473
R3378 VSS.n9579 VSS.n9578 3.27473
R3379 VSS.n199 VSS.n198 3.27473
R3380 VSS.n477 VSS.n476 3.27473
R3381 VSS.n9030 VSS.n9029 3.27473
R3382 VSS.n270 VSS.n269 3.27473
R3383 VSS.n342 VSS.n341 3.27473
R3384 VSS.n414 VSS.n413 3.27473
R3385 VSS.t633 VSS.t430 3.2333
R3386 VSS.n1391 VSS.t588 3.19467
R3387 VSS.n10325 VSS.n10323 3.15563
R3388 VSS.n10329 VSS.n10327 3.15563
R3389 VSS.n10318 VSS.n10316 3.15563
R3390 VSS.n10314 VSS.n10312 3.15563
R3391 VSS.n10757 VSS.n10756 3.1505
R3392 VSS.n10767 VSS.n10766 3.1505
R3393 VSS.n11289 VSS.t283 3.02895
R3394 VSS.n10309 VSS.n10308 3.02463
R3395 VSS.n10408 VSS.n10406 2.96616
R3396 VSS.n10401 VSS.n10399 2.96616
R3397 VSS.n10378 VSS.n10377 2.885
R3398 VSS.n10623 VSS.n10622 2.885
R3399 VSS.n10614 VSS.n10613 2.795
R3400 VSS.n10408 VSS.n10407 2.76247
R3401 VSS.n10401 VSS.n10400 2.76247
R3402 VSS.n10297 VSS.n10296 2.74471
R3403 VSS.n10403 VSS.n10401 2.71914
R3404 VSS.n10326 VSS.n10322 2.71872
R3405 VSS.n9526 VSS.t263 2.71016
R3406 VSS.n10818 VSS.t3204 2.6955
R3407 VSS.n10814 VSS.t1908 2.6955
R3408 VSS.n10748 VSS.t889 2.6955
R3409 VSS.n10752 VSS.t581 2.6955
R3410 VSS.n10787 VSS.t3544 2.6955
R3411 VSS.n10783 VSS.t2233 2.6955
R3412 VSS.n10781 VSS.t1263 2.6955
R3413 VSS.n10777 VSS.t962 2.6955
R3414 VSS.n9193 VSS.n9192 2.68042
R3415 VSS.n9188 VSS.n9187 2.68042
R3416 VSS.n9329 VSS.n9328 2.68042
R3417 VSS.n9324 VSS.n9323 2.68042
R3418 VSS.n167 VSS.n166 2.68042
R3419 VSS.n162 VSS.n161 2.68042
R3420 VSS.n9575 VSS.n9574 2.68042
R3421 VSS.n9570 VSS.n9569 2.68042
R3422 VSS.n9026 VSS.n9025 2.68042
R3423 VSS.n9021 VSS.n9020 2.68042
R3424 VSS.n190 VSS.n189 2.68012
R3425 VSS.n195 VSS.n194 2.68012
R3426 VSS.n468 VSS.n467 2.68012
R3427 VSS.n473 VSS.n472 2.68012
R3428 VSS.n261 VSS.n260 2.68012
R3429 VSS.n266 VSS.n265 2.68012
R3430 VSS.n333 VSS.n332 2.68012
R3431 VSS.n338 VSS.n337 2.68012
R3432 VSS.n405 VSS.n404 2.68012
R3433 VSS.n410 VSS.n409 2.68012
R3434 VSS.n4804 VSS.n4803 2.66637
R3435 VSS.n10866 VSS.n10864 2.65976
R3436 VSS.n9560 VSS.t265 2.63047
R3437 VSS.n10769 VSS.t3148 2.6255
R3438 VSS.n10772 VSS.t1822 2.6255
R3439 VSS.n10770 VSS.t3598 2.6255
R3440 VSS.n10741 VSS.t2227 2.6255
R3441 VSS.n10745 VSS.t3238 2.6255
R3442 VSS.n10663 VSS.n10662 2.60959
R3443 VSS.n9612 VSS.n813 2.58721
R3444 VSS.n9877 VSS.n669 2.58721
R3445 VSS.n656 VSS.n655 2.58721
R3446 VSS.n821 VSS.n820 2.58721
R3447 VSS.n677 VSS.n676 2.58721
R3448 VSS.n11416 VSS.n45 2.58721
R3449 VSS.n11449 VSS.n20 2.58721
R3450 VSS.n9920 VSS.n585 2.58721
R3451 VSS.n9913 VSS.n9908 2.58721
R3452 VSS.n9513 VSS.n1329 2.58721
R3453 VSS.n1253 VSS.n1252 2.58721
R3454 VSS.n9901 VSS.n9900 2.58721
R3455 VSS.n652 VSS.n651 2.58366
R3456 VSS.n817 VSS.n816 2.58366
R3457 VSS.n9858 VSS.n9857 2.58366
R3458 VSS.n9874 VSS.n670 2.58366
R3459 VSS.n11413 VSS.n46 2.58366
R3460 VSS.n11446 VSS.n21 2.58366
R3461 VSS.n9897 VSS.n629 2.58366
R3462 VSS.n1249 VSS.n1248 2.58366
R3463 VSS.n9516 VSS.n1328 2.58366
R3464 VSS.n9910 VSS.n9909 2.58366
R3465 VSS.n9924 VSS.n9923 2.58366
R3466 VSS.n9615 VSS.n812 2.58366
R3467 VSS.n10325 VSS.n10324 2.573
R3468 VSS.n10329 VSS.n10328 2.573
R3469 VSS.n10318 VSS.n10317 2.573
R3470 VSS.n10314 VSS.n10313 2.573
R3471 VSS.n10625 VSS.n10624 2.55405
R3472 VSS.n10616 VSS.n10615 2.55405
R3473 VSS.n10380 VSS.n10379 2.55405
R3474 VSS.t378 VSS.t745 2.55077
R3475 VSS.n10733 VSS.t1755 2.5394
R3476 VSS.t1243 VSS.n9434 2.53859
R3477 VSS.n9447 VSS.t2094 2.53837
R3478 VSS.n11304 VSS.t3417 2.53699
R3479 VSS.t3565 VSS.n10838 2.52844
R3480 VSS.n10839 VSS.t3565 2.52844
R3481 VSS.t816 VSS.n10835 2.52844
R3482 VSS.n10836 VSS.t816 2.52844
R3483 VSS.t2464 VSS.n10832 2.52844
R3484 VSS.n10833 VSS.t2464 2.52844
R3485 VSS.t1191 VSS.n10829 2.52844
R3486 VSS.n10830 VSS.t1191 2.52844
R3487 VSS.t3011 VSS.n10826 2.52844
R3488 VSS.n10827 VSS.t3011 2.52844
R3489 VSS.n10727 VSS.t1755 2.52844
R3490 VSS.t3523 VSS.n10725 2.52844
R3491 VSS.n10726 VSS.t3523 2.52844
R3492 VSS.t762 VSS.n10723 2.52844
R3493 VSS.n10724 VSS.t762 2.52844
R3494 VSS.t2432 VSS.n10721 2.52844
R3495 VSS.n10722 VSS.t2432 2.52844
R3496 VSS.t1130 VSS.n10718 2.52844
R3497 VSS.n10719 VSS.t1130 2.52844
R3498 VSS.n10717 VSS.t2957 2.52844
R3499 VSS.t2957 VSS.n10716 2.52844
R3500 VSS.t1673 VSS.n10714 2.52844
R3501 VSS.n10715 VSS.t1673 2.52844
R3502 VSS.t3417 VSS.n125 2.52844
R3503 VSS.n1338 VSS.t1693 2.52844
R3504 VSS.t1693 VSS.n1337 2.52844
R3505 VSS.n1341 VSS.t2551 2.52844
R3506 VSS.t2551 VSS.n1340 2.52844
R3507 VSS.n9499 VSS.t1739 2.52844
R3508 VSS.t1739 VSS.n1343 2.52844
R3509 VSS.n9496 VSS.t483 2.52844
R3510 VSS.t483 VSS.n9495 2.52844
R3511 VSS.t2999 VSS.n9491 2.52844
R3512 VSS.n9492 VSS.t2999 2.52844
R3513 VSS.t1549 VSS.n9488 2.52844
R3514 VSS.n9489 VSS.t1549 2.52844
R3515 VSS.n9445 VSS.t2094 2.52844
R3516 VSS.t2997 VSS.n9443 2.52844
R3517 VSS.n9444 VSS.t2997 2.52844
R3518 VSS.t2152 VSS.n9441 2.52844
R3519 VSS.n9442 VSS.t2152 2.52844
R3520 VSS.t3339 VSS.n9438 2.52844
R3521 VSS.n9439 VSS.t3339 2.52844
R3522 VSS.t2705 VSS.n9436 2.52844
R3523 VSS.n9437 VSS.t2705 2.52844
R3524 VSS.n9435 VSS.t1243 2.52844
R3525 VSS.n10410 VSS.n10403 2.46014
R3526 VSS.n10796 VSS.n247 2.45973
R3527 VSS.n10808 VSS.n10807 2.45073
R3528 VSS.n10333 VSS.n10321 2.38034
R3529 VSS.n10392 VSS.n10365 2.37491
R3530 VSS.n10398 VSS.n10397 2.32143
R3531 VSS.n11152 VSS.n181 2.31168
R3532 VSS.n10611 VSS.n10610 2.30076
R3533 VSS.n10018 VSS.n576 2.28095
R3534 VSS.n573 VSS.n572 2.28095
R3535 VSS.n1356 VSS.n1353 2.28095
R3536 VSS.n10020 VSS.n576 2.27641
R3537 VSS.n10025 VSS.n572 2.27641
R3538 VSS.n1358 VSS.n1353 2.27641
R3539 VSS.n228 VSS.n227 2.26832
R3540 VSS.n10679 VSS.n10303 2.26738
R3541 VSS.n5468 VSS.n2743 2.2505
R3542 VSS.n5467 VSS.n5466 2.2505
R3543 VSS.n5465 VSS.n2744 2.2505
R3544 VSS.n5464 VSS.n5463 2.2505
R3545 VSS.n5462 VSS.n2745 2.2505
R3546 VSS.n5461 VSS.n5460 2.2505
R3547 VSS.n5459 VSS.n2746 2.2505
R3548 VSS.n5458 VSS.n5457 2.2505
R3549 VSS.n5456 VSS.n2747 2.2505
R3550 VSS.n5455 VSS.n5454 2.2505
R3551 VSS.n5453 VSS.n2748 2.2505
R3552 VSS.n5452 VSS.n5451 2.2505
R3553 VSS.n5450 VSS.n2749 2.2505
R3554 VSS.n5449 VSS.n5448 2.2505
R3555 VSS.n5447 VSS.n2750 2.2505
R3556 VSS.n5446 VSS.n5445 2.2505
R3557 VSS.n5444 VSS.n2751 2.2505
R3558 VSS.n5443 VSS.n5442 2.2505
R3559 VSS.n5441 VSS.n2752 2.2505
R3560 VSS.n5440 VSS.n5439 2.2505
R3561 VSS.n5438 VSS.n2753 2.2505
R3562 VSS.n5437 VSS.n5436 2.2505
R3563 VSS.n5435 VSS.n2754 2.2505
R3564 VSS.n5434 VSS.n5433 2.2505
R3565 VSS.n5432 VSS.n2755 2.2505
R3566 VSS.n5431 VSS.n5430 2.2505
R3567 VSS.n5429 VSS.n2756 2.2505
R3568 VSS.n5428 VSS.n5427 2.2505
R3569 VSS.n5426 VSS.n2757 2.2505
R3570 VSS.n5425 VSS.n5424 2.2505
R3571 VSS.n5423 VSS.n2758 2.2505
R3572 VSS.n5422 VSS.n5421 2.2505
R3573 VSS.n5420 VSS.n2759 2.2505
R3574 VSS.n5419 VSS.n5418 2.2505
R3575 VSS.n5417 VSS.n2760 2.2505
R3576 VSS.n5416 VSS.n5415 2.2505
R3577 VSS.n5414 VSS.n2761 2.2505
R3578 VSS.n5413 VSS.n5412 2.2505
R3579 VSS.n5411 VSS.n2762 2.2505
R3580 VSS.n5410 VSS.n5409 2.2505
R3581 VSS.n5408 VSS.n2763 2.2505
R3582 VSS.n5407 VSS.n5406 2.2505
R3583 VSS.n5405 VSS.n2764 2.2505
R3584 VSS.n5404 VSS.n5403 2.2505
R3585 VSS.n5402 VSS.n2765 2.2505
R3586 VSS.n5401 VSS.n5400 2.2505
R3587 VSS.n5399 VSS.n2766 2.2505
R3588 VSS.n5398 VSS.n5397 2.2505
R3589 VSS.n5396 VSS.n2767 2.2505
R3590 VSS.n5395 VSS.n5394 2.2505
R3591 VSS.n5393 VSS.n2768 2.2505
R3592 VSS.n5392 VSS.n5391 2.2505
R3593 VSS.n5390 VSS.n2769 2.2505
R3594 VSS.n5389 VSS.n5388 2.2505
R3595 VSS.n5387 VSS.n2770 2.2505
R3596 VSS.n5386 VSS.n5385 2.2505
R3597 VSS.n5384 VSS.n2771 2.2505
R3598 VSS.n5383 VSS.n5382 2.2505
R3599 VSS.n5381 VSS.n2772 2.2505
R3600 VSS.n5380 VSS.n5379 2.2505
R3601 VSS.n5378 VSS.n2773 2.2505
R3602 VSS.n5377 VSS.n5376 2.2505
R3603 VSS.n5375 VSS.n2774 2.2505
R3604 VSS.n5374 VSS.n5373 2.2505
R3605 VSS.n5372 VSS.n2775 2.2505
R3606 VSS.n5371 VSS.n5370 2.2505
R3607 VSS.n5369 VSS.n2776 2.2505
R3608 VSS.n5368 VSS.n5367 2.2505
R3609 VSS.n5366 VSS.n2777 2.2505
R3610 VSS.n5365 VSS.n5364 2.2505
R3611 VSS.n5363 VSS.n2778 2.2505
R3612 VSS.n5362 VSS.n5361 2.2505
R3613 VSS.n5360 VSS.n2779 2.2505
R3614 VSS.n5359 VSS.n5358 2.2505
R3615 VSS.n5357 VSS.n2780 2.2505
R3616 VSS.n5356 VSS.n5355 2.2505
R3617 VSS.n5354 VSS.n2781 2.2505
R3618 VSS.n5353 VSS.n5352 2.2505
R3619 VSS.n5351 VSS.n2782 2.2505
R3620 VSS.n5350 VSS.n5349 2.2505
R3621 VSS.n5348 VSS.n2783 2.2505
R3622 VSS.n5347 VSS.n5346 2.2505
R3623 VSS.n5345 VSS.n2784 2.2505
R3624 VSS.n5344 VSS.n5343 2.2505
R3625 VSS.n5342 VSS.n2785 2.2505
R3626 VSS.n5341 VSS.n5340 2.2505
R3627 VSS.n5339 VSS.n2786 2.2505
R3628 VSS.n5338 VSS.n5337 2.2505
R3629 VSS.n5336 VSS.n2787 2.2505
R3630 VSS.n5335 VSS.n5334 2.2505
R3631 VSS.n5333 VSS.n2788 2.2505
R3632 VSS.n5332 VSS.n5331 2.2505
R3633 VSS.n5330 VSS.n2789 2.2505
R3634 VSS.n5329 VSS.n5328 2.2505
R3635 VSS.n5327 VSS.n2790 2.2505
R3636 VSS.n5326 VSS.n5325 2.2505
R3637 VSS.n5324 VSS.n2791 2.2505
R3638 VSS.n5323 VSS.n5322 2.2505
R3639 VSS.n5321 VSS.n2792 2.2505
R3640 VSS.n5320 VSS.n5319 2.2505
R3641 VSS.n5318 VSS.n2793 2.2505
R3642 VSS.n5317 VSS.n5316 2.2505
R3643 VSS.n5315 VSS.n2794 2.2505
R3644 VSS.n5314 VSS.n5313 2.2505
R3645 VSS.n5312 VSS.n2795 2.2505
R3646 VSS.n5311 VSS.n5310 2.2505
R3647 VSS.n5309 VSS.n2796 2.2505
R3648 VSS.n5308 VSS.n5307 2.2505
R3649 VSS.n5306 VSS.n2797 2.2505
R3650 VSS.n5305 VSS.n5304 2.2505
R3651 VSS.n5303 VSS.n2798 2.2505
R3652 VSS.n5302 VSS.n5301 2.2505
R3653 VSS.n5300 VSS.n2799 2.2505
R3654 VSS.n5299 VSS.n5298 2.2505
R3655 VSS.n5297 VSS.n2800 2.2505
R3656 VSS.n5296 VSS.n5295 2.2505
R3657 VSS.n5294 VSS.n2801 2.2505
R3658 VSS.n5293 VSS.n5292 2.2505
R3659 VSS.n5291 VSS.n2802 2.2505
R3660 VSS.n5290 VSS.n5289 2.2505
R3661 VSS.n5288 VSS.n2803 2.2505
R3662 VSS.n5287 VSS.n5286 2.2505
R3663 VSS.n5285 VSS.n2804 2.2505
R3664 VSS.n5284 VSS.n5283 2.2505
R3665 VSS.n5282 VSS.n2805 2.2505
R3666 VSS.n5281 VSS.n5280 2.2505
R3667 VSS.n5279 VSS.n2806 2.2505
R3668 VSS.n5278 VSS.n5277 2.2505
R3669 VSS.n5276 VSS.n2807 2.2505
R3670 VSS.n5275 VSS.n5274 2.2505
R3671 VSS.n5273 VSS.n2808 2.2505
R3672 VSS.n5272 VSS.n5271 2.2505
R3673 VSS.n5270 VSS.n2809 2.2505
R3674 VSS.n5269 VSS.n5268 2.2505
R3675 VSS.n5267 VSS.n2810 2.2505
R3676 VSS.n5266 VSS.n5265 2.2505
R3677 VSS.n5264 VSS.n2811 2.2505
R3678 VSS.n5263 VSS.n5262 2.2505
R3679 VSS.n5261 VSS.n2812 2.2505
R3680 VSS.n5260 VSS.n5259 2.2505
R3681 VSS.n5258 VSS.n2813 2.2505
R3682 VSS.n5257 VSS.n5256 2.2505
R3683 VSS.n5255 VSS.n2814 2.2505
R3684 VSS.n5254 VSS.n5253 2.2505
R3685 VSS.n5252 VSS.n2815 2.2505
R3686 VSS.n5251 VSS.n5250 2.2505
R3687 VSS.n5249 VSS.n2816 2.2505
R3688 VSS.n5248 VSS.n5247 2.2505
R3689 VSS.n5246 VSS.n2817 2.2505
R3690 VSS.n5245 VSS.n5244 2.2505
R3691 VSS.n5243 VSS.n2818 2.2505
R3692 VSS.n5242 VSS.n5241 2.2505
R3693 VSS.n5240 VSS.n2819 2.2505
R3694 VSS.n5239 VSS.n5238 2.2505
R3695 VSS.n5237 VSS.n2820 2.2505
R3696 VSS.n5236 VSS.n5235 2.2505
R3697 VSS.n5234 VSS.n2821 2.2505
R3698 VSS.n5233 VSS.n5232 2.2505
R3699 VSS.n5231 VSS.n2822 2.2505
R3700 VSS.n5230 VSS.n5229 2.2505
R3701 VSS.n5228 VSS.n2823 2.2505
R3702 VSS.n5227 VSS.n5226 2.2505
R3703 VSS.n5225 VSS.n2824 2.2505
R3704 VSS.n5224 VSS.n5223 2.2505
R3705 VSS.n5222 VSS.n2825 2.2505
R3706 VSS.n5221 VSS.n5220 2.2505
R3707 VSS.n5219 VSS.n2826 2.2505
R3708 VSS.n5218 VSS.n5217 2.2505
R3709 VSS.n5216 VSS.n2827 2.2505
R3710 VSS.n5215 VSS.n5214 2.2505
R3711 VSS.n5213 VSS.n2828 2.2505
R3712 VSS.n5212 VSS.n5211 2.2505
R3713 VSS.n5210 VSS.n2829 2.2505
R3714 VSS.n5209 VSS.n5208 2.2505
R3715 VSS.n5207 VSS.n2830 2.2505
R3716 VSS.n5206 VSS.n5205 2.2505
R3717 VSS.n5204 VSS.n2831 2.2505
R3718 VSS.n5203 VSS.n5202 2.2505
R3719 VSS.n5201 VSS.n2832 2.2505
R3720 VSS.n5200 VSS.n5199 2.2505
R3721 VSS.n5198 VSS.n2833 2.2505
R3722 VSS.n5197 VSS.n5196 2.2505
R3723 VSS.n5195 VSS.n2834 2.2505
R3724 VSS.n5194 VSS.n5193 2.2505
R3725 VSS.n5192 VSS.n2835 2.2505
R3726 VSS.n5191 VSS.n5190 2.2505
R3727 VSS.n5189 VSS.n2836 2.2505
R3728 VSS.n5188 VSS.n5187 2.2505
R3729 VSS.n5186 VSS.n2837 2.2505
R3730 VSS.n5185 VSS.n5184 2.2505
R3731 VSS.n5183 VSS.n2838 2.2505
R3732 VSS.n5182 VSS.n5181 2.2505
R3733 VSS.n5180 VSS.n2839 2.2505
R3734 VSS.n5179 VSS.n5178 2.2505
R3735 VSS.n5177 VSS.n2840 2.2505
R3736 VSS.n5176 VSS.n5175 2.2505
R3737 VSS.n5174 VSS.n2841 2.2505
R3738 VSS.n5173 VSS.n5172 2.2505
R3739 VSS.n5171 VSS.n2842 2.2505
R3740 VSS.n5170 VSS.n5169 2.2505
R3741 VSS.n5168 VSS.n2843 2.2505
R3742 VSS.n5167 VSS.n5166 2.2505
R3743 VSS.n5165 VSS.n2844 2.2505
R3744 VSS.n5164 VSS.n5163 2.2505
R3745 VSS.n5162 VSS.n2845 2.2505
R3746 VSS.n5161 VSS.n5160 2.2505
R3747 VSS.n5159 VSS.n2846 2.2505
R3748 VSS.n5158 VSS.n5157 2.2505
R3749 VSS.n5156 VSS.n2847 2.2505
R3750 VSS.n5155 VSS.n5154 2.2505
R3751 VSS.n5153 VSS.n2848 2.2505
R3752 VSS.n5152 VSS.n5151 2.2505
R3753 VSS.n5150 VSS.n2849 2.2505
R3754 VSS.n5149 VSS.n5148 2.2505
R3755 VSS.n5147 VSS.n2850 2.2505
R3756 VSS.n5146 VSS.n5145 2.2505
R3757 VSS.n5144 VSS.n2851 2.2505
R3758 VSS.n5143 VSS.n5142 2.2505
R3759 VSS.n5141 VSS.n2852 2.2505
R3760 VSS.n5140 VSS.n5139 2.2505
R3761 VSS.n5138 VSS.n2853 2.2505
R3762 VSS.n5137 VSS.n5136 2.2505
R3763 VSS.n5135 VSS.n2854 2.2505
R3764 VSS.n5134 VSS.n5133 2.2505
R3765 VSS.n5132 VSS.n2855 2.2505
R3766 VSS.n5131 VSS.n5130 2.2505
R3767 VSS.n5129 VSS.n2856 2.2505
R3768 VSS.n5128 VSS.n5127 2.2505
R3769 VSS.n5126 VSS.n2857 2.2505
R3770 VSS.n5125 VSS.n5124 2.2505
R3771 VSS.n5123 VSS.n2858 2.2505
R3772 VSS.n5122 VSS.n5121 2.2505
R3773 VSS.n5120 VSS.n2859 2.2505
R3774 VSS.n5119 VSS.n5118 2.2505
R3775 VSS.n5117 VSS.n2860 2.2505
R3776 VSS.n5116 VSS.n5115 2.2505
R3777 VSS.n5114 VSS.n2861 2.2505
R3778 VSS.n5113 VSS.n5112 2.2505
R3779 VSS.n5111 VSS.n2862 2.2505
R3780 VSS.n5110 VSS.n5109 2.2505
R3781 VSS.n5108 VSS.n2863 2.2505
R3782 VSS.n5107 VSS.n5106 2.2505
R3783 VSS.n5105 VSS.n2864 2.2505
R3784 VSS.n5104 VSS.n5103 2.2505
R3785 VSS.n5102 VSS.n2865 2.2505
R3786 VSS.n5101 VSS.n5100 2.2505
R3787 VSS.n5099 VSS.n2866 2.2505
R3788 VSS.n5098 VSS.n5097 2.2505
R3789 VSS.n5096 VSS.n2867 2.2505
R3790 VSS.n5095 VSS.n5094 2.2505
R3791 VSS.n5093 VSS.n2868 2.2505
R3792 VSS.n5092 VSS.n5091 2.2505
R3793 VSS.n5090 VSS.n2869 2.2505
R3794 VSS.n5089 VSS.n5088 2.2505
R3795 VSS.n5087 VSS.n2870 2.2505
R3796 VSS.n5086 VSS.n5085 2.2505
R3797 VSS.n5084 VSS.n2871 2.2505
R3798 VSS.n5083 VSS.n5082 2.2505
R3799 VSS.n5081 VSS.n2872 2.2505
R3800 VSS.n5080 VSS.n5079 2.2505
R3801 VSS.n5078 VSS.n2873 2.2505
R3802 VSS.n5077 VSS.n5076 2.2505
R3803 VSS.n5075 VSS.n2874 2.2505
R3804 VSS.n5074 VSS.n5073 2.2505
R3805 VSS.n5072 VSS.n2875 2.2505
R3806 VSS.n5071 VSS.n5070 2.2505
R3807 VSS.n5069 VSS.n2876 2.2505
R3808 VSS.n5068 VSS.n5067 2.2505
R3809 VSS.n5066 VSS.n2877 2.2505
R3810 VSS.n5065 VSS.n5064 2.2505
R3811 VSS.n5063 VSS.n2878 2.2505
R3812 VSS.n5062 VSS.n5061 2.2505
R3813 VSS.n5060 VSS.n2879 2.2505
R3814 VSS.n5059 VSS.n5058 2.2505
R3815 VSS.n5057 VSS.n2880 2.2505
R3816 VSS.n5056 VSS.n5055 2.2505
R3817 VSS.n5054 VSS.n2881 2.2505
R3818 VSS.n5053 VSS.n5052 2.2505
R3819 VSS.n5051 VSS.n2882 2.2505
R3820 VSS.n5050 VSS.n5049 2.2505
R3821 VSS.n5048 VSS.n2883 2.2505
R3822 VSS.n5047 VSS.n5046 2.2505
R3823 VSS.n5045 VSS.n2884 2.2505
R3824 VSS.n5044 VSS.n5043 2.2505
R3825 VSS.n5042 VSS.n2885 2.2505
R3826 VSS.n5041 VSS.n5040 2.2505
R3827 VSS.n5039 VSS.n2886 2.2505
R3828 VSS.n5038 VSS.n5037 2.2505
R3829 VSS.n5036 VSS.n2887 2.2505
R3830 VSS.n5035 VSS.n5034 2.2505
R3831 VSS.n5033 VSS.n2888 2.2505
R3832 VSS.n5032 VSS.n5031 2.2505
R3833 VSS.n5030 VSS.n2889 2.2505
R3834 VSS.n5029 VSS.n5028 2.2505
R3835 VSS.n5027 VSS.n2890 2.2505
R3836 VSS.n5026 VSS.n5025 2.2505
R3837 VSS.n5024 VSS.n2891 2.2505
R3838 VSS.n5023 VSS.n5022 2.2505
R3839 VSS.n5021 VSS.n2892 2.2505
R3840 VSS.n5020 VSS.n5019 2.2505
R3841 VSS.n5018 VSS.n2893 2.2505
R3842 VSS.n5017 VSS.n5016 2.2505
R3843 VSS.n5015 VSS.n2894 2.2505
R3844 VSS.n5014 VSS.n5013 2.2505
R3845 VSS.n5012 VSS.n2895 2.2505
R3846 VSS.n5011 VSS.n5010 2.2505
R3847 VSS.n5009 VSS.n2896 2.2505
R3848 VSS.n5008 VSS.n5007 2.2505
R3849 VSS.n5006 VSS.n2897 2.2505
R3850 VSS.n5005 VSS.n5004 2.2505
R3851 VSS.n5003 VSS.n2898 2.2505
R3852 VSS.n5002 VSS.n5001 2.2505
R3853 VSS.n5000 VSS.n2899 2.2505
R3854 VSS.n4999 VSS.n4998 2.2505
R3855 VSS.n4997 VSS.n2900 2.2505
R3856 VSS.n4996 VSS.n4995 2.2505
R3857 VSS.n4994 VSS.n2901 2.2505
R3858 VSS.n4993 VSS.n4992 2.2505
R3859 VSS.n4991 VSS.n2902 2.2505
R3860 VSS.n4990 VSS.n4989 2.2505
R3861 VSS.n4988 VSS.n2903 2.2505
R3862 VSS.n4987 VSS.n4986 2.2505
R3863 VSS.n4985 VSS.n2904 2.2505
R3864 VSS.n4984 VSS.n4983 2.2505
R3865 VSS.n4982 VSS.n2905 2.2505
R3866 VSS.n4981 VSS.n4980 2.2505
R3867 VSS.n4979 VSS.n2906 2.2505
R3868 VSS.n4978 VSS.n4977 2.2505
R3869 VSS.n4976 VSS.n2907 2.2505
R3870 VSS.n4975 VSS.n4974 2.2505
R3871 VSS.n4973 VSS.n2908 2.2505
R3872 VSS.n4972 VSS.n4971 2.2505
R3873 VSS.n4970 VSS.n2909 2.2505
R3874 VSS.n4969 VSS.n4968 2.2505
R3875 VSS.n4967 VSS.n2910 2.2505
R3876 VSS.n4966 VSS.n4965 2.2505
R3877 VSS.n4964 VSS.n2911 2.2505
R3878 VSS.n4963 VSS.n4962 2.2505
R3879 VSS.n4961 VSS.n2912 2.2505
R3880 VSS.n4960 VSS.n4959 2.2505
R3881 VSS.n4958 VSS.n2913 2.2505
R3882 VSS.n4957 VSS.n4956 2.2505
R3883 VSS.n4955 VSS.n2914 2.2505
R3884 VSS.n4954 VSS.n4953 2.2505
R3885 VSS.n4952 VSS.n2915 2.2505
R3886 VSS.n4951 VSS.n4950 2.2505
R3887 VSS.n4949 VSS.n2916 2.2505
R3888 VSS.n4948 VSS.n4947 2.2505
R3889 VSS.n4946 VSS.n2917 2.2505
R3890 VSS.n4945 VSS.n4944 2.2505
R3891 VSS.n4943 VSS.n2918 2.2505
R3892 VSS.n4942 VSS.n4941 2.2505
R3893 VSS.n4940 VSS.n2919 2.2505
R3894 VSS.n4939 VSS.n4938 2.2505
R3895 VSS.n4937 VSS.n2920 2.2505
R3896 VSS.n4936 VSS.n4935 2.2505
R3897 VSS.n4934 VSS.n2921 2.2505
R3898 VSS.n4933 VSS.n4932 2.2505
R3899 VSS.n4931 VSS.n2922 2.2505
R3900 VSS.n4930 VSS.n4929 2.2505
R3901 VSS.n4928 VSS.n2923 2.2505
R3902 VSS.n4927 VSS.n4926 2.2505
R3903 VSS.n4925 VSS.n2924 2.2505
R3904 VSS.n4924 VSS.n4923 2.2505
R3905 VSS.n4922 VSS.n2925 2.2505
R3906 VSS.n4921 VSS.n4920 2.2505
R3907 VSS.n4919 VSS.n2926 2.2505
R3908 VSS.n4918 VSS.n4917 2.2505
R3909 VSS.n4916 VSS.n2927 2.2505
R3910 VSS.n4915 VSS.n4914 2.2505
R3911 VSS.n4913 VSS.n2928 2.2505
R3912 VSS.n4912 VSS.n4911 2.2505
R3913 VSS.n4910 VSS.n2929 2.2505
R3914 VSS.n4909 VSS.n4908 2.2505
R3915 VSS.n4907 VSS.n2930 2.2505
R3916 VSS.n4906 VSS.n4905 2.2505
R3917 VSS.n4904 VSS.n2931 2.2505
R3918 VSS.n4903 VSS.n4902 2.2505
R3919 VSS.n4901 VSS.n2932 2.2505
R3920 VSS.n4900 VSS.n4899 2.2505
R3921 VSS.n4898 VSS.n2933 2.2505
R3922 VSS.n4897 VSS.n4896 2.2505
R3923 VSS.n4895 VSS.n2934 2.2505
R3924 VSS.n4894 VSS.n4893 2.2505
R3925 VSS.n4892 VSS.n2935 2.2505
R3926 VSS.n4891 VSS.n4890 2.2505
R3927 VSS.n4889 VSS.n2936 2.2505
R3928 VSS.n4888 VSS.n4887 2.2505
R3929 VSS.n4886 VSS.n2937 2.2505
R3930 VSS.n4885 VSS.n4884 2.2505
R3931 VSS.n4883 VSS.n2938 2.2505
R3932 VSS.n4882 VSS.n4881 2.2505
R3933 VSS.n4880 VSS.n2939 2.2505
R3934 VSS.n4879 VSS.n4878 2.2505
R3935 VSS.n4877 VSS.n2940 2.2505
R3936 VSS.n4876 VSS.n4875 2.2505
R3937 VSS.n4874 VSS.n2941 2.2505
R3938 VSS.n4873 VSS.n4872 2.2505
R3939 VSS.n4871 VSS.n2942 2.2505
R3940 VSS.n4870 VSS.n4869 2.2505
R3941 VSS.n4868 VSS.n2943 2.2505
R3942 VSS.n4867 VSS.n4866 2.2505
R3943 VSS.n4865 VSS.n2944 2.2505
R3944 VSS.n4864 VSS.n4863 2.2505
R3945 VSS.n4862 VSS.n2945 2.2505
R3946 VSS.n4861 VSS.n4860 2.2505
R3947 VSS.n4859 VSS.n2946 2.2505
R3948 VSS.n4858 VSS.n4857 2.2505
R3949 VSS.n4856 VSS.n2947 2.2505
R3950 VSS.n4855 VSS.n4854 2.2505
R3951 VSS.n4853 VSS.n2948 2.2505
R3952 VSS.n4852 VSS.n4851 2.2505
R3953 VSS.n4850 VSS.n2949 2.2505
R3954 VSS.n4849 VSS.n4848 2.2505
R3955 VSS.n4847 VSS.n2950 2.2505
R3956 VSS.n4846 VSS.n4845 2.2505
R3957 VSS.n4844 VSS.n2951 2.2505
R3958 VSS.n4843 VSS.n4842 2.2505
R3959 VSS.n4841 VSS.n2952 2.2505
R3960 VSS.n4840 VSS.n4839 2.2505
R3961 VSS.n4838 VSS.n2953 2.2505
R3962 VSS.n4837 VSS.n4836 2.2505
R3963 VSS.n4835 VSS.n2954 2.2505
R3964 VSS.n4834 VSS.n4833 2.2505
R3965 VSS.n4832 VSS.n2955 2.2505
R3966 VSS.n4831 VSS.n4830 2.2505
R3967 VSS.n4829 VSS.n2956 2.2505
R3968 VSS.n4828 VSS.n4827 2.2505
R3969 VSS.n4826 VSS.n2957 2.2505
R3970 VSS.n4825 VSS.n4824 2.2505
R3971 VSS.n4823 VSS.n2958 2.2505
R3972 VSS.n4822 VSS.n4821 2.2505
R3973 VSS.n4820 VSS.n2959 2.2505
R3974 VSS.n4819 VSS.n4818 2.2505
R3975 VSS.n4817 VSS.n2960 2.2505
R3976 VSS.n4816 VSS.n4815 2.2505
R3977 VSS.n4814 VSS.n2961 2.2505
R3978 VSS.n4813 VSS.n4812 2.2505
R3979 VSS.n4811 VSS.n2962 2.2505
R3980 VSS.n4810 VSS.n4809 2.2505
R3981 VSS.n4808 VSS.n2963 2.2505
R3982 VSS.n4807 VSS.n4806 2.2505
R3983 VSS.n4802 VSS.n2964 2.2505
R3984 VSS.n4801 VSS.n4800 2.2505
R3985 VSS.n4799 VSS.n2965 2.2505
R3986 VSS.n4798 VSS.n4797 2.2505
R3987 VSS.n4796 VSS.n2966 2.2505
R3988 VSS.n4795 VSS.n4794 2.2505
R3989 VSS.n4793 VSS.n2967 2.2505
R3990 VSS.n4792 VSS.n4791 2.2505
R3991 VSS.n4790 VSS.n2968 2.2505
R3992 VSS.n4789 VSS.n4788 2.2505
R3993 VSS.n4787 VSS.n2969 2.2505
R3994 VSS.n4786 VSS.n4785 2.2505
R3995 VSS.n4784 VSS.n2970 2.2505
R3996 VSS.n4783 VSS.n4782 2.2505
R3997 VSS.n4781 VSS.n2971 2.2505
R3998 VSS.n4780 VSS.n4779 2.2505
R3999 VSS.n4778 VSS.n2972 2.2505
R4000 VSS.n4777 VSS.n4776 2.2505
R4001 VSS.n4775 VSS.n2973 2.2505
R4002 VSS.n4774 VSS.n4773 2.2505
R4003 VSS.n4772 VSS.n2974 2.2505
R4004 VSS.n4771 VSS.n4770 2.2505
R4005 VSS.n4769 VSS.n2975 2.2505
R4006 VSS.n4768 VSS.n4767 2.2505
R4007 VSS.n4766 VSS.n2976 2.2505
R4008 VSS.n4765 VSS.n4764 2.2505
R4009 VSS.n4763 VSS.n2977 2.2505
R4010 VSS.n4762 VSS.n4761 2.2505
R4011 VSS.n4760 VSS.n2978 2.2505
R4012 VSS.n4759 VSS.n4758 2.2505
R4013 VSS.n4757 VSS.n2979 2.2505
R4014 VSS.n4756 VSS.n4755 2.2505
R4015 VSS.n4754 VSS.n2980 2.2505
R4016 VSS.n4753 VSS.n4752 2.2505
R4017 VSS.n4751 VSS.n2981 2.2505
R4018 VSS.n4750 VSS.n4749 2.2505
R4019 VSS.n4748 VSS.n2982 2.2505
R4020 VSS.n4747 VSS.n4746 2.2505
R4021 VSS.n4745 VSS.n2983 2.2505
R4022 VSS.n4744 VSS.n4743 2.2505
R4023 VSS.n4742 VSS.n2984 2.2505
R4024 VSS.n4741 VSS.n4740 2.2505
R4025 VSS.n4739 VSS.n2985 2.2505
R4026 VSS.n4738 VSS.n4737 2.2505
R4027 VSS.n4736 VSS.n2986 2.2505
R4028 VSS.n4735 VSS.n4734 2.2505
R4029 VSS.n4733 VSS.n2987 2.2505
R4030 VSS.n4732 VSS.n4731 2.2505
R4031 VSS.n4730 VSS.n2988 2.2505
R4032 VSS.n4729 VSS.n4728 2.2505
R4033 VSS.n4727 VSS.n2989 2.2505
R4034 VSS.n4726 VSS.n4725 2.2505
R4035 VSS.n4724 VSS.n2990 2.2505
R4036 VSS.n4723 VSS.n4722 2.2505
R4037 VSS.n4721 VSS.n2991 2.2505
R4038 VSS.n4720 VSS.n4719 2.2505
R4039 VSS.n4718 VSS.n2992 2.2505
R4040 VSS.n4717 VSS.n4716 2.2505
R4041 VSS.n4715 VSS.n2993 2.2505
R4042 VSS.n4714 VSS.n4713 2.2505
R4043 VSS.n4712 VSS.n2994 2.2505
R4044 VSS.n4711 VSS.n4710 2.2505
R4045 VSS.n4709 VSS.n2995 2.2505
R4046 VSS.n4708 VSS.n4707 2.2505
R4047 VSS.n4706 VSS.n2996 2.2505
R4048 VSS.n4705 VSS.n4704 2.2505
R4049 VSS.n4703 VSS.n2997 2.2505
R4050 VSS.n4702 VSS.n4701 2.2505
R4051 VSS.n4700 VSS.n2998 2.2505
R4052 VSS.n4699 VSS.n4698 2.2505
R4053 VSS.n4697 VSS.n2999 2.2505
R4054 VSS.n4696 VSS.n4695 2.2505
R4055 VSS.n4694 VSS.n3000 2.2505
R4056 VSS.n4693 VSS.n4692 2.2505
R4057 VSS.n4691 VSS.n3001 2.2505
R4058 VSS.n4690 VSS.n4689 2.2505
R4059 VSS.n4688 VSS.n3002 2.2505
R4060 VSS.n4687 VSS.n4686 2.2505
R4061 VSS.n4685 VSS.n3003 2.2505
R4062 VSS.n4684 VSS.n4683 2.2505
R4063 VSS.n4682 VSS.n3004 2.2505
R4064 VSS.n4681 VSS.n4680 2.2505
R4065 VSS.n4679 VSS.n3005 2.2505
R4066 VSS.n4678 VSS.n4677 2.2505
R4067 VSS.n4676 VSS.n3006 2.2505
R4068 VSS.n4675 VSS.n4674 2.2505
R4069 VSS.n4673 VSS.n3007 2.2505
R4070 VSS.n4672 VSS.n4671 2.2505
R4071 VSS.n4670 VSS.n3008 2.2505
R4072 VSS.n4669 VSS.n4668 2.2505
R4073 VSS.n4667 VSS.n3009 2.2505
R4074 VSS.n4666 VSS.n4665 2.2505
R4075 VSS.n4664 VSS.n3010 2.2505
R4076 VSS.n4663 VSS.n4662 2.2505
R4077 VSS.n4661 VSS.n3011 2.2505
R4078 VSS.n4660 VSS.n4659 2.2505
R4079 VSS.n4658 VSS.n3012 2.2505
R4080 VSS.n4657 VSS.n4656 2.2505
R4081 VSS.n4655 VSS.n3013 2.2505
R4082 VSS.n4654 VSS.n4653 2.2505
R4083 VSS.n4652 VSS.n3014 2.2505
R4084 VSS.n4651 VSS.n4650 2.2505
R4085 VSS.n4649 VSS.n3015 2.2505
R4086 VSS.n4648 VSS.n4647 2.2505
R4087 VSS.n4646 VSS.n3016 2.2505
R4088 VSS.n4645 VSS.n4644 2.2505
R4089 VSS.n4643 VSS.n3017 2.2505
R4090 VSS.n4642 VSS.n4641 2.2505
R4091 VSS.n4640 VSS.n3018 2.2505
R4092 VSS.n4639 VSS.n4638 2.2505
R4093 VSS.n4637 VSS.n3019 2.2505
R4094 VSS.n4636 VSS.n4635 2.2505
R4095 VSS.n4634 VSS.n3020 2.2505
R4096 VSS.n4633 VSS.n4632 2.2505
R4097 VSS.n4631 VSS.n3021 2.2505
R4098 VSS.n4630 VSS.n4629 2.2505
R4099 VSS.n4628 VSS.n3022 2.2505
R4100 VSS.n4627 VSS.n4626 2.2505
R4101 VSS.n4625 VSS.n3023 2.2505
R4102 VSS.n4624 VSS.n4623 2.2505
R4103 VSS.n4622 VSS.n3024 2.2505
R4104 VSS.n4621 VSS.n4620 2.2505
R4105 VSS.n4619 VSS.n3025 2.2505
R4106 VSS.n4618 VSS.n4617 2.2505
R4107 VSS.n4616 VSS.n3026 2.2505
R4108 VSS.n4615 VSS.n4614 2.2505
R4109 VSS.n4613 VSS.n3027 2.2505
R4110 VSS.n4612 VSS.n4611 2.2505
R4111 VSS.n4610 VSS.n3028 2.2505
R4112 VSS.n4609 VSS.n4608 2.2505
R4113 VSS.n4607 VSS.n3029 2.2505
R4114 VSS.n4606 VSS.n4605 2.2505
R4115 VSS.n4604 VSS.n3030 2.2505
R4116 VSS.n4603 VSS.n4602 2.2505
R4117 VSS.n4601 VSS.n3031 2.2505
R4118 VSS.n4600 VSS.n4599 2.2505
R4119 VSS.n4598 VSS.n3032 2.2505
R4120 VSS.n4597 VSS.n4596 2.2505
R4121 VSS.n4595 VSS.n3033 2.2505
R4122 VSS.n4594 VSS.n4593 2.2505
R4123 VSS.n4592 VSS.n3034 2.2505
R4124 VSS.n4591 VSS.n4590 2.2505
R4125 VSS.n4589 VSS.n3035 2.2505
R4126 VSS.n4588 VSS.n4587 2.2505
R4127 VSS.n4586 VSS.n3036 2.2505
R4128 VSS.n4585 VSS.n4584 2.2505
R4129 VSS.n4583 VSS.n3037 2.2505
R4130 VSS.n4582 VSS.n4581 2.2505
R4131 VSS.n4580 VSS.n3038 2.2505
R4132 VSS.n4579 VSS.n4578 2.2505
R4133 VSS.n4577 VSS.n3039 2.2505
R4134 VSS.n4576 VSS.n4575 2.2505
R4135 VSS.n4574 VSS.n3040 2.2505
R4136 VSS.n4573 VSS.n4572 2.2505
R4137 VSS.n4571 VSS.n3041 2.2505
R4138 VSS.n4570 VSS.n4569 2.2505
R4139 VSS.n4568 VSS.n3042 2.2505
R4140 VSS.n4567 VSS.n4566 2.2505
R4141 VSS.n4565 VSS.n3043 2.2505
R4142 VSS.n4564 VSS.n4563 2.2505
R4143 VSS.n4562 VSS.n3044 2.2505
R4144 VSS.n4561 VSS.n4560 2.2505
R4145 VSS.n4559 VSS.n3045 2.2505
R4146 VSS.n4558 VSS.n4557 2.2505
R4147 VSS.n4556 VSS.n3046 2.2505
R4148 VSS.n4555 VSS.n4554 2.2505
R4149 VSS.n4553 VSS.n3047 2.2505
R4150 VSS.n4552 VSS.n4551 2.2505
R4151 VSS.n4550 VSS.n3048 2.2505
R4152 VSS.n4549 VSS.n4548 2.2505
R4153 VSS.n4547 VSS.n3049 2.2505
R4154 VSS.n4546 VSS.n4545 2.2505
R4155 VSS.n4544 VSS.n3050 2.2505
R4156 VSS.n4543 VSS.n4542 2.2505
R4157 VSS.n4541 VSS.n3051 2.2505
R4158 VSS.n4540 VSS.n4539 2.2505
R4159 VSS.n4538 VSS.n3052 2.2505
R4160 VSS.n4537 VSS.n4536 2.2505
R4161 VSS.n4535 VSS.n3053 2.2505
R4162 VSS.n4534 VSS.n4533 2.2505
R4163 VSS.n4532 VSS.n3054 2.2505
R4164 VSS.n4531 VSS.n4530 2.2505
R4165 VSS.n4529 VSS.n3055 2.2505
R4166 VSS.n4528 VSS.n4527 2.2505
R4167 VSS.n4526 VSS.n3056 2.2505
R4168 VSS.n4525 VSS.n4524 2.2505
R4169 VSS.n4523 VSS.n3057 2.2505
R4170 VSS.n4522 VSS.n4521 2.2505
R4171 VSS.n4520 VSS.n3058 2.2505
R4172 VSS.n4519 VSS.n4518 2.2505
R4173 VSS.n4517 VSS.n3059 2.2505
R4174 VSS.n4516 VSS.n4515 2.2505
R4175 VSS.n4514 VSS.n3060 2.2505
R4176 VSS.n4513 VSS.n4512 2.2505
R4177 VSS.n4511 VSS.n3061 2.2505
R4178 VSS.n4510 VSS.n4509 2.2505
R4179 VSS.n4508 VSS.n3062 2.2505
R4180 VSS.n4507 VSS.n4506 2.2505
R4181 VSS.n4505 VSS.n3063 2.2505
R4182 VSS.n4504 VSS.n4503 2.2505
R4183 VSS.n4502 VSS.n3064 2.2505
R4184 VSS.n4501 VSS.n4500 2.2505
R4185 VSS.n4499 VSS.n3065 2.2505
R4186 VSS.n4498 VSS.n4497 2.2505
R4187 VSS.n4496 VSS.n3066 2.2505
R4188 VSS.n4495 VSS.n4494 2.2505
R4189 VSS.n4493 VSS.n3067 2.2505
R4190 VSS.n4492 VSS.n4491 2.2505
R4191 VSS.n4490 VSS.n3068 2.2505
R4192 VSS.n4489 VSS.n4488 2.2505
R4193 VSS.n4487 VSS.n3069 2.2505
R4194 VSS.n4486 VSS.n4485 2.2505
R4195 VSS.n4484 VSS.n3070 2.2505
R4196 VSS.n4483 VSS.n4482 2.2505
R4197 VSS.n4481 VSS.n3071 2.2505
R4198 VSS.n4480 VSS.n4479 2.2505
R4199 VSS.n4478 VSS.n3072 2.2505
R4200 VSS.n4477 VSS.n4476 2.2505
R4201 VSS.n4475 VSS.n3073 2.2505
R4202 VSS.n4474 VSS.n4473 2.2505
R4203 VSS.n4472 VSS.n3074 2.2505
R4204 VSS.n4471 VSS.n4470 2.2505
R4205 VSS.n4469 VSS.n3075 2.2505
R4206 VSS.n4468 VSS.n4467 2.2505
R4207 VSS.n4466 VSS.n3076 2.2505
R4208 VSS.n4465 VSS.n4464 2.2505
R4209 VSS.n4463 VSS.n3077 2.2505
R4210 VSS.n4462 VSS.n4461 2.2505
R4211 VSS.n4460 VSS.n3078 2.2505
R4212 VSS.n4459 VSS.n4458 2.2505
R4213 VSS.n4457 VSS.n3079 2.2505
R4214 VSS.n4456 VSS.n4455 2.2505
R4215 VSS.n4454 VSS.n3080 2.2505
R4216 VSS.n4453 VSS.n4452 2.2505
R4217 VSS.n4451 VSS.n3081 2.2505
R4218 VSS.n4450 VSS.n4449 2.2505
R4219 VSS.n4448 VSS.n3082 2.2505
R4220 VSS.n4447 VSS.n4446 2.2505
R4221 VSS.n4445 VSS.n3083 2.2505
R4222 VSS.n4444 VSS.n4443 2.2505
R4223 VSS.n4442 VSS.n3084 2.2505
R4224 VSS.n4441 VSS.n4440 2.2505
R4225 VSS.n4439 VSS.n3085 2.2505
R4226 VSS.n4438 VSS.n4437 2.2505
R4227 VSS.n4436 VSS.n3086 2.2505
R4228 VSS.n4435 VSS.n4434 2.2505
R4229 VSS.n4433 VSS.n3087 2.2505
R4230 VSS.n4432 VSS.n4431 2.2505
R4231 VSS.n4430 VSS.n3088 2.2505
R4232 VSS.n4429 VSS.n4428 2.2505
R4233 VSS.n4427 VSS.n3089 2.2505
R4234 VSS.n4426 VSS.n4425 2.2505
R4235 VSS.n4424 VSS.n3090 2.2505
R4236 VSS.n4423 VSS.n4422 2.2505
R4237 VSS.n4421 VSS.n3091 2.2505
R4238 VSS.n4420 VSS.n4419 2.2505
R4239 VSS.n4418 VSS.n3092 2.2505
R4240 VSS.n4417 VSS.n4416 2.2505
R4241 VSS.n4415 VSS.n3093 2.2505
R4242 VSS.n4414 VSS.n4413 2.2505
R4243 VSS.n4412 VSS.n3094 2.2505
R4244 VSS.n4411 VSS.n4410 2.2505
R4245 VSS.n4409 VSS.n3095 2.2505
R4246 VSS.n4408 VSS.n4407 2.2505
R4247 VSS.n4406 VSS.n3096 2.2505
R4248 VSS.n4405 VSS.n4404 2.2505
R4249 VSS.n4403 VSS.n3097 2.2505
R4250 VSS.n4402 VSS.n4401 2.2505
R4251 VSS.n4400 VSS.n3098 2.2505
R4252 VSS.n4399 VSS.n4398 2.2505
R4253 VSS.n4397 VSS.n3099 2.2505
R4254 VSS.n4396 VSS.n4395 2.2505
R4255 VSS.n4394 VSS.n3100 2.2505
R4256 VSS.n4393 VSS.n4392 2.2505
R4257 VSS.n4391 VSS.n3101 2.2505
R4258 VSS.n4390 VSS.n4389 2.2505
R4259 VSS.n4388 VSS.n3102 2.2505
R4260 VSS.n4387 VSS.n4386 2.2505
R4261 VSS.n4385 VSS.n3103 2.2505
R4262 VSS.n4384 VSS.n4383 2.2505
R4263 VSS.n4382 VSS.n3104 2.2505
R4264 VSS.n4381 VSS.n4380 2.2505
R4265 VSS.n4379 VSS.n3105 2.2505
R4266 VSS.n4378 VSS.n4377 2.2505
R4267 VSS.n4376 VSS.n3106 2.2505
R4268 VSS.n4375 VSS.n4374 2.2505
R4269 VSS.n4373 VSS.n3107 2.2505
R4270 VSS.n4372 VSS.n4371 2.2505
R4271 VSS.n4370 VSS.n3108 2.2505
R4272 VSS.n4369 VSS.n4368 2.2505
R4273 VSS.n4367 VSS.n3109 2.2505
R4274 VSS.n4366 VSS.n4365 2.2505
R4275 VSS.n4364 VSS.n3110 2.2505
R4276 VSS.n4363 VSS.n4362 2.2505
R4277 VSS.n4361 VSS.n3111 2.2505
R4278 VSS.n4360 VSS.n4359 2.2505
R4279 VSS.n4358 VSS.n3112 2.2505
R4280 VSS.n4357 VSS.n4356 2.2505
R4281 VSS.n4355 VSS.n3113 2.2505
R4282 VSS.n4354 VSS.n4353 2.2505
R4283 VSS.n4352 VSS.n3114 2.2505
R4284 VSS.n4351 VSS.n4350 2.2505
R4285 VSS.n4349 VSS.n3115 2.2505
R4286 VSS.n4348 VSS.n4347 2.2505
R4287 VSS.n4346 VSS.n3116 2.2505
R4288 VSS.n4345 VSS.n4344 2.2505
R4289 VSS.n4343 VSS.n3117 2.2505
R4290 VSS.n4342 VSS.n4341 2.2505
R4291 VSS.n4340 VSS.n3118 2.2505
R4292 VSS.n4339 VSS.n4338 2.2505
R4293 VSS.n4337 VSS.n3119 2.2505
R4294 VSS.n4336 VSS.n4335 2.2505
R4295 VSS.n4334 VSS.n3120 2.2505
R4296 VSS.n4333 VSS.n4332 2.2505
R4297 VSS.n4331 VSS.n3121 2.2505
R4298 VSS.n4330 VSS.n4329 2.2505
R4299 VSS.n4328 VSS.n3122 2.2505
R4300 VSS.n4327 VSS.n4326 2.2505
R4301 VSS.n4325 VSS.n3123 2.2505
R4302 VSS.n4324 VSS.n4323 2.2505
R4303 VSS.n4322 VSS.n3124 2.2505
R4304 VSS.n4321 VSS.n4320 2.2505
R4305 VSS.n4319 VSS.n3125 2.2505
R4306 VSS.n4318 VSS.n4317 2.2505
R4307 VSS.n4316 VSS.n3126 2.2505
R4308 VSS.n4315 VSS.n4314 2.2505
R4309 VSS.n4313 VSS.n3127 2.2505
R4310 VSS.n4312 VSS.n4311 2.2505
R4311 VSS.n4310 VSS.n3128 2.2505
R4312 VSS.n4309 VSS.n4308 2.2505
R4313 VSS.n4307 VSS.n3129 2.2505
R4314 VSS.n4306 VSS.n4305 2.2505
R4315 VSS.n4304 VSS.n3130 2.2505
R4316 VSS.n4303 VSS.n4302 2.2505
R4317 VSS.n4301 VSS.n3131 2.2505
R4318 VSS.n4300 VSS.n4299 2.2505
R4319 VSS.n4298 VSS.n3132 2.2505
R4320 VSS.n4297 VSS.n4296 2.2505
R4321 VSS.n4295 VSS.n3133 2.2505
R4322 VSS.n4294 VSS.n4293 2.2505
R4323 VSS.n4292 VSS.n3134 2.2505
R4324 VSS.n4291 VSS.n4290 2.2505
R4325 VSS.n4289 VSS.n3135 2.2505
R4326 VSS.n4288 VSS.n4287 2.2505
R4327 VSS.n4286 VSS.n3136 2.2505
R4328 VSS.n4285 VSS.n4284 2.2505
R4329 VSS.n4283 VSS.n3137 2.2505
R4330 VSS.n4282 VSS.n4281 2.2505
R4331 VSS.n4280 VSS.n3138 2.2505
R4332 VSS.n4279 VSS.n4278 2.2505
R4333 VSS.n4277 VSS.n3139 2.2505
R4334 VSS.n4276 VSS.n4275 2.2505
R4335 VSS.n4274 VSS.n3140 2.2505
R4336 VSS.n4273 VSS.n4272 2.2505
R4337 VSS.n4271 VSS.n3141 2.2505
R4338 VSS.n4270 VSS.n4269 2.2505
R4339 VSS.n4268 VSS.n3142 2.2505
R4340 VSS.n4267 VSS.n4266 2.2505
R4341 VSS.n4265 VSS.n3143 2.2505
R4342 VSS.n4264 VSS.n4263 2.2505
R4343 VSS.n4262 VSS.n3144 2.2505
R4344 VSS.n4261 VSS.n4260 2.2505
R4345 VSS.n4259 VSS.n3145 2.2505
R4346 VSS.n4258 VSS.n4257 2.2505
R4347 VSS.n4256 VSS.n3146 2.2505
R4348 VSS.n4255 VSS.n4254 2.2505
R4349 VSS.n4253 VSS.n3147 2.2505
R4350 VSS.n4252 VSS.n4251 2.2505
R4351 VSS.n4250 VSS.n3148 2.2505
R4352 VSS.n4249 VSS.n4248 2.2505
R4353 VSS.n4247 VSS.n3149 2.2505
R4354 VSS.n4246 VSS.n4245 2.2505
R4355 VSS.n4244 VSS.n3150 2.2505
R4356 VSS.n4243 VSS.n4242 2.2505
R4357 VSS.n4241 VSS.n3151 2.2505
R4358 VSS.n4240 VSS.n4239 2.2505
R4359 VSS.n4238 VSS.n3152 2.2505
R4360 VSS.n4237 VSS.n4236 2.2505
R4361 VSS.n4235 VSS.n3153 2.2505
R4362 VSS.n4234 VSS.n4233 2.2505
R4363 VSS.n4232 VSS.n3154 2.2505
R4364 VSS.n4231 VSS.n4230 2.2505
R4365 VSS.n4229 VSS.n3155 2.2505
R4366 VSS.n4228 VSS.n4227 2.2505
R4367 VSS.n4226 VSS.n3156 2.2505
R4368 VSS.n4225 VSS.n4224 2.2505
R4369 VSS.n4223 VSS.n3157 2.2505
R4370 VSS.n4222 VSS.n4221 2.2505
R4371 VSS.n4220 VSS.n3158 2.2505
R4372 VSS.n4219 VSS.n4218 2.2505
R4373 VSS.n4217 VSS.n3159 2.2505
R4374 VSS.n4216 VSS.n4215 2.2505
R4375 VSS.n4214 VSS.n3160 2.2505
R4376 VSS.n4213 VSS.n4212 2.2505
R4377 VSS.n4211 VSS.n3161 2.2505
R4378 VSS.n4210 VSS.n4209 2.2505
R4379 VSS.n4208 VSS.n3162 2.2505
R4380 VSS.n4207 VSS.n4206 2.2505
R4381 VSS.n4205 VSS.n3163 2.2505
R4382 VSS.n4204 VSS.n4203 2.2505
R4383 VSS.n4202 VSS.n3164 2.2505
R4384 VSS.n4201 VSS.n4200 2.2505
R4385 VSS.n4199 VSS.n3165 2.2505
R4386 VSS.n4198 VSS.n4197 2.2505
R4387 VSS.n4196 VSS.n3166 2.2505
R4388 VSS.n4195 VSS.n4194 2.2505
R4389 VSS.n4193 VSS.n3167 2.2505
R4390 VSS.n4192 VSS.n4191 2.2505
R4391 VSS.n4190 VSS.n3168 2.2505
R4392 VSS.n4189 VSS.n4188 2.2505
R4393 VSS.n4187 VSS.n3169 2.2505
R4394 VSS.n4186 VSS.n4185 2.2505
R4395 VSS.n4184 VSS.n3170 2.2505
R4396 VSS.n4183 VSS.n4182 2.2505
R4397 VSS.n4181 VSS.n3171 2.2505
R4398 VSS.n4180 VSS.n4179 2.2505
R4399 VSS.n4178 VSS.n3172 2.2505
R4400 VSS.n4177 VSS.n4176 2.2505
R4401 VSS.n4175 VSS.n3173 2.2505
R4402 VSS.n4174 VSS.n4173 2.2505
R4403 VSS.n4172 VSS.n3174 2.2505
R4404 VSS.n4171 VSS.n4170 2.2505
R4405 VSS.n4169 VSS.n3175 2.2505
R4406 VSS.n4168 VSS.n4167 2.2505
R4407 VSS.n4166 VSS.n3176 2.2505
R4408 VSS.n4165 VSS.n4164 2.2505
R4409 VSS.n4163 VSS.n3177 2.2505
R4410 VSS.n4162 VSS.n4161 2.2505
R4411 VSS.n4160 VSS.n3178 2.2505
R4412 VSS.n4159 VSS.n4158 2.2505
R4413 VSS.n4157 VSS.n3179 2.2505
R4414 VSS.n4156 VSS.n4155 2.2505
R4415 VSS.n4154 VSS.n3180 2.2505
R4416 VSS.n4153 VSS.n4152 2.2505
R4417 VSS.n4151 VSS.n3181 2.2505
R4418 VSS.n4150 VSS.n4149 2.2505
R4419 VSS.n4148 VSS.n3182 2.2505
R4420 VSS.n4147 VSS.n4146 2.2505
R4421 VSS.n4145 VSS.n3183 2.2505
R4422 VSS.n4144 VSS.n4143 2.2505
R4423 VSS.n4142 VSS.n3184 2.2505
R4424 VSS.n6907 VSS.n6906 2.2505
R4425 VSS.n6905 VSS.n2264 2.2505
R4426 VSS.n6904 VSS.n6903 2.2505
R4427 VSS.n6902 VSS.n2265 2.2505
R4428 VSS.n6901 VSS.n6900 2.2505
R4429 VSS.n6899 VSS.n2266 2.2505
R4430 VSS.n6898 VSS.n6897 2.2505
R4431 VSS.n6896 VSS.n2267 2.2505
R4432 VSS.n6895 VSS.n6894 2.2505
R4433 VSS.n6893 VSS.n2268 2.2505
R4434 VSS.n6892 VSS.n6891 2.2505
R4435 VSS.n6890 VSS.n2269 2.2505
R4436 VSS.n6889 VSS.n6888 2.2505
R4437 VSS.n6887 VSS.n2270 2.2505
R4438 VSS.n6886 VSS.n6885 2.2505
R4439 VSS.n6884 VSS.n2271 2.2505
R4440 VSS.n6883 VSS.n6882 2.2505
R4441 VSS.n6881 VSS.n2272 2.2505
R4442 VSS.n6880 VSS.n6879 2.2505
R4443 VSS.n6878 VSS.n2273 2.2505
R4444 VSS.n6877 VSS.n6876 2.2505
R4445 VSS.n6875 VSS.n2274 2.2505
R4446 VSS.n6874 VSS.n6873 2.2505
R4447 VSS.n6872 VSS.n2275 2.2505
R4448 VSS.n6871 VSS.n6870 2.2505
R4449 VSS.n6869 VSS.n2276 2.2505
R4450 VSS.n6868 VSS.n6867 2.2505
R4451 VSS.n6866 VSS.n2277 2.2505
R4452 VSS.n6865 VSS.n6864 2.2505
R4453 VSS.n6863 VSS.n2278 2.2505
R4454 VSS.n6862 VSS.n6861 2.2505
R4455 VSS.n6860 VSS.n2279 2.2505
R4456 VSS.n6859 VSS.n6858 2.2505
R4457 VSS.n6857 VSS.n2280 2.2505
R4458 VSS.n6856 VSS.n6855 2.2505
R4459 VSS.n6854 VSS.n2281 2.2505
R4460 VSS.n6853 VSS.n6852 2.2505
R4461 VSS.n6851 VSS.n2282 2.2505
R4462 VSS.n6850 VSS.n6849 2.2505
R4463 VSS.n6848 VSS.n2283 2.2505
R4464 VSS.n6847 VSS.n6846 2.2505
R4465 VSS.n6845 VSS.n2284 2.2505
R4466 VSS.n6844 VSS.n6843 2.2505
R4467 VSS.n6842 VSS.n2285 2.2505
R4468 VSS.n6841 VSS.n6840 2.2505
R4469 VSS.n6839 VSS.n2286 2.2505
R4470 VSS.n6838 VSS.n6837 2.2505
R4471 VSS.n6836 VSS.n2287 2.2505
R4472 VSS.n6835 VSS.n6834 2.2505
R4473 VSS.n6833 VSS.n2288 2.2505
R4474 VSS.n6832 VSS.n6831 2.2505
R4475 VSS.n6830 VSS.n2289 2.2505
R4476 VSS.n6829 VSS.n6828 2.2505
R4477 VSS.n6827 VSS.n2290 2.2505
R4478 VSS.n6826 VSS.n6825 2.2505
R4479 VSS.n6824 VSS.n2291 2.2505
R4480 VSS.n6823 VSS.n6822 2.2505
R4481 VSS.n6821 VSS.n2292 2.2505
R4482 VSS.n6820 VSS.n6819 2.2505
R4483 VSS.n6818 VSS.n2293 2.2505
R4484 VSS.n6817 VSS.n6816 2.2505
R4485 VSS.n6815 VSS.n2294 2.2505
R4486 VSS.n6814 VSS.n6813 2.2505
R4487 VSS.n6812 VSS.n2295 2.2505
R4488 VSS.n6811 VSS.n6810 2.2505
R4489 VSS.n6809 VSS.n2296 2.2505
R4490 VSS.n6808 VSS.n6807 2.2505
R4491 VSS.n6806 VSS.n2297 2.2505
R4492 VSS.n6805 VSS.n6804 2.2505
R4493 VSS.n6803 VSS.n2298 2.2505
R4494 VSS.n6802 VSS.n6801 2.2505
R4495 VSS.n6800 VSS.n2299 2.2505
R4496 VSS.n6799 VSS.n6798 2.2505
R4497 VSS.n6797 VSS.n2300 2.2505
R4498 VSS.n6796 VSS.n6795 2.2505
R4499 VSS.n6794 VSS.n2301 2.2505
R4500 VSS.n6793 VSS.n6792 2.2505
R4501 VSS.n6791 VSS.n2302 2.2505
R4502 VSS.n6790 VSS.n6789 2.2505
R4503 VSS.n6788 VSS.n2303 2.2505
R4504 VSS.n6787 VSS.n6786 2.2505
R4505 VSS.n6785 VSS.n2304 2.2505
R4506 VSS.n6784 VSS.n6783 2.2505
R4507 VSS.n6782 VSS.n2305 2.2505
R4508 VSS.n6781 VSS.n6780 2.2505
R4509 VSS.n6779 VSS.n2306 2.2505
R4510 VSS.n6778 VSS.n6777 2.2505
R4511 VSS.n6776 VSS.n2307 2.2505
R4512 VSS.n6775 VSS.n6774 2.2505
R4513 VSS.n6773 VSS.n2308 2.2505
R4514 VSS.n6772 VSS.n6771 2.2505
R4515 VSS.n6770 VSS.n2309 2.2505
R4516 VSS.n6769 VSS.n6768 2.2505
R4517 VSS.n6767 VSS.n2310 2.2505
R4518 VSS.n6766 VSS.n6765 2.2505
R4519 VSS.n6764 VSS.n2311 2.2505
R4520 VSS.n6763 VSS.n6762 2.2505
R4521 VSS.n6761 VSS.n2312 2.2505
R4522 VSS.n6760 VSS.n6759 2.2505
R4523 VSS.n6758 VSS.n2313 2.2505
R4524 VSS.n6757 VSS.n6756 2.2505
R4525 VSS.n6755 VSS.n2314 2.2505
R4526 VSS.n6754 VSS.n6753 2.2505
R4527 VSS.n6752 VSS.n2315 2.2505
R4528 VSS.n6751 VSS.n6750 2.2505
R4529 VSS.n6749 VSS.n2316 2.2505
R4530 VSS.n6748 VSS.n6747 2.2505
R4531 VSS.n6746 VSS.n2317 2.2505
R4532 VSS.n6745 VSS.n6744 2.2505
R4533 VSS.n6743 VSS.n2318 2.2505
R4534 VSS.n6742 VSS.n6741 2.2505
R4535 VSS.n6740 VSS.n2319 2.2505
R4536 VSS.n6739 VSS.n6738 2.2505
R4537 VSS.n6737 VSS.n2320 2.2505
R4538 VSS.n6736 VSS.n6735 2.2505
R4539 VSS.n6734 VSS.n2321 2.2505
R4540 VSS.n6733 VSS.n6732 2.2505
R4541 VSS.n6731 VSS.n2322 2.2505
R4542 VSS.n6730 VSS.n6729 2.2505
R4543 VSS.n6728 VSS.n2323 2.2505
R4544 VSS.n6727 VSS.n6726 2.2505
R4545 VSS.n6725 VSS.n2324 2.2505
R4546 VSS.n6724 VSS.n6723 2.2505
R4547 VSS.n6722 VSS.n2325 2.2505
R4548 VSS.n6721 VSS.n6720 2.2505
R4549 VSS.n6719 VSS.n2326 2.2505
R4550 VSS.n6718 VSS.n6717 2.2505
R4551 VSS.n6716 VSS.n2327 2.2505
R4552 VSS.n6715 VSS.n6714 2.2505
R4553 VSS.n6713 VSS.n2328 2.2505
R4554 VSS.n6712 VSS.n6711 2.2505
R4555 VSS.n6710 VSS.n2329 2.2505
R4556 VSS.n6709 VSS.n6708 2.2505
R4557 VSS.n6707 VSS.n2330 2.2505
R4558 VSS.n6706 VSS.n6705 2.2505
R4559 VSS.n6704 VSS.n2331 2.2505
R4560 VSS.n6703 VSS.n6702 2.2505
R4561 VSS.n6701 VSS.n2332 2.2505
R4562 VSS.n6700 VSS.n6699 2.2505
R4563 VSS.n6698 VSS.n2333 2.2505
R4564 VSS.n6697 VSS.n6696 2.2505
R4565 VSS.n6695 VSS.n2334 2.2505
R4566 VSS.n6694 VSS.n6693 2.2505
R4567 VSS.n6692 VSS.n2335 2.2505
R4568 VSS.n6691 VSS.n6690 2.2505
R4569 VSS.n6689 VSS.n2336 2.2505
R4570 VSS.n6688 VSS.n6687 2.2505
R4571 VSS.n6686 VSS.n2337 2.2505
R4572 VSS.n6685 VSS.n6684 2.2505
R4573 VSS.n6683 VSS.n2338 2.2505
R4574 VSS.n6682 VSS.n6681 2.2505
R4575 VSS.n6680 VSS.n2339 2.2505
R4576 VSS.n6679 VSS.n6678 2.2505
R4577 VSS.n6677 VSS.n2340 2.2505
R4578 VSS.n6676 VSS.n6675 2.2505
R4579 VSS.n6674 VSS.n2341 2.2505
R4580 VSS.n6673 VSS.n6672 2.2505
R4581 VSS.n6671 VSS.n2342 2.2505
R4582 VSS.n6670 VSS.n6669 2.2505
R4583 VSS.n6668 VSS.n2343 2.2505
R4584 VSS.n6667 VSS.n6666 2.2505
R4585 VSS.n6665 VSS.n2344 2.2505
R4586 VSS.n6664 VSS.n6663 2.2505
R4587 VSS.n6662 VSS.n2345 2.2505
R4588 VSS.n6661 VSS.n6660 2.2505
R4589 VSS.n6659 VSS.n2346 2.2505
R4590 VSS.n6658 VSS.n6657 2.2505
R4591 VSS.n6656 VSS.n2347 2.2505
R4592 VSS.n6655 VSS.n6654 2.2505
R4593 VSS.n6653 VSS.n2348 2.2505
R4594 VSS.n6652 VSS.n6651 2.2505
R4595 VSS.n6650 VSS.n2349 2.2505
R4596 VSS.n6649 VSS.n6648 2.2505
R4597 VSS.n6647 VSS.n2350 2.2505
R4598 VSS.n6646 VSS.n6645 2.2505
R4599 VSS.n6644 VSS.n2351 2.2505
R4600 VSS.n6643 VSS.n6642 2.2505
R4601 VSS.n6641 VSS.n2352 2.2505
R4602 VSS.n6640 VSS.n6639 2.2505
R4603 VSS.n6638 VSS.n2353 2.2505
R4604 VSS.n6637 VSS.n6636 2.2505
R4605 VSS.n6635 VSS.n2354 2.2505
R4606 VSS.n6634 VSS.n6633 2.2505
R4607 VSS.n6632 VSS.n2355 2.2505
R4608 VSS.n6631 VSS.n6630 2.2505
R4609 VSS.n6629 VSS.n2356 2.2505
R4610 VSS.n6628 VSS.n6627 2.2505
R4611 VSS.n6626 VSS.n2357 2.2505
R4612 VSS.n6625 VSS.n6624 2.2505
R4613 VSS.n6623 VSS.n2358 2.2505
R4614 VSS.n6622 VSS.n6621 2.2505
R4615 VSS.n6620 VSS.n2359 2.2505
R4616 VSS.n6619 VSS.n6618 2.2505
R4617 VSS.n6617 VSS.n2360 2.2505
R4618 VSS.n6616 VSS.n6615 2.2505
R4619 VSS.n6614 VSS.n2361 2.2505
R4620 VSS.n6613 VSS.n6612 2.2505
R4621 VSS.n6611 VSS.n2362 2.2505
R4622 VSS.n6610 VSS.n6609 2.2505
R4623 VSS.n6608 VSS.n2363 2.2505
R4624 VSS.n6607 VSS.n6606 2.2505
R4625 VSS.n6605 VSS.n2364 2.2505
R4626 VSS.n6604 VSS.n6603 2.2505
R4627 VSS.n6602 VSS.n2365 2.2505
R4628 VSS.n6601 VSS.n6600 2.2505
R4629 VSS.n6599 VSS.n2366 2.2505
R4630 VSS.n6598 VSS.n6597 2.2505
R4631 VSS.n6596 VSS.n2367 2.2505
R4632 VSS.n6595 VSS.n6594 2.2505
R4633 VSS.n6593 VSS.n2368 2.2505
R4634 VSS.n6592 VSS.n6591 2.2505
R4635 VSS.n6590 VSS.n2369 2.2505
R4636 VSS.n6589 VSS.n6588 2.2505
R4637 VSS.n6587 VSS.n2370 2.2505
R4638 VSS.n6586 VSS.n6585 2.2505
R4639 VSS.n6584 VSS.n2371 2.2505
R4640 VSS.n6583 VSS.n6582 2.2505
R4641 VSS.n6581 VSS.n2372 2.2505
R4642 VSS.n6580 VSS.n6579 2.2505
R4643 VSS.n6578 VSS.n2373 2.2505
R4644 VSS.n6577 VSS.n6576 2.2505
R4645 VSS.n6575 VSS.n2374 2.2505
R4646 VSS.n6574 VSS.n6573 2.2505
R4647 VSS.n6572 VSS.n2375 2.2505
R4648 VSS.n6571 VSS.n6570 2.2505
R4649 VSS.n6569 VSS.n2376 2.2505
R4650 VSS.n6568 VSS.n6567 2.2505
R4651 VSS.n6566 VSS.n2377 2.2505
R4652 VSS.n6565 VSS.n6564 2.2505
R4653 VSS.n6563 VSS.n2378 2.2505
R4654 VSS.n6562 VSS.n6561 2.2505
R4655 VSS.n6560 VSS.n2379 2.2505
R4656 VSS.n6559 VSS.n6558 2.2505
R4657 VSS.n6557 VSS.n2380 2.2505
R4658 VSS.n6556 VSS.n6555 2.2505
R4659 VSS.n6554 VSS.n2381 2.2505
R4660 VSS.n6553 VSS.n6552 2.2505
R4661 VSS.n6551 VSS.n2382 2.2505
R4662 VSS.n6550 VSS.n6549 2.2505
R4663 VSS.n6548 VSS.n2383 2.2505
R4664 VSS.n6547 VSS.n6546 2.2505
R4665 VSS.n6545 VSS.n2384 2.2505
R4666 VSS.n6544 VSS.n6543 2.2505
R4667 VSS.n6542 VSS.n2385 2.2505
R4668 VSS.n6541 VSS.n6540 2.2505
R4669 VSS.n6539 VSS.n2386 2.2505
R4670 VSS.n6538 VSS.n6537 2.2505
R4671 VSS.n6536 VSS.n2387 2.2505
R4672 VSS.n6535 VSS.n6534 2.2505
R4673 VSS.n6533 VSS.n2388 2.2505
R4674 VSS.n6532 VSS.n6531 2.2505
R4675 VSS.n6530 VSS.n2389 2.2505
R4676 VSS.n6529 VSS.n6528 2.2505
R4677 VSS.n6527 VSS.n2390 2.2505
R4678 VSS.n6526 VSS.n6525 2.2505
R4679 VSS.n6524 VSS.n2391 2.2505
R4680 VSS.n6523 VSS.n6522 2.2505
R4681 VSS.n6521 VSS.n2392 2.2505
R4682 VSS.n6520 VSS.n6519 2.2505
R4683 VSS.n6518 VSS.n2393 2.2505
R4684 VSS.n6517 VSS.n6516 2.2505
R4685 VSS.n6515 VSS.n2394 2.2505
R4686 VSS.n6514 VSS.n6513 2.2505
R4687 VSS.n6512 VSS.n2395 2.2505
R4688 VSS.n6511 VSS.n6510 2.2505
R4689 VSS.n6509 VSS.n2396 2.2505
R4690 VSS.n6508 VSS.n6507 2.2505
R4691 VSS.n6506 VSS.n2397 2.2505
R4692 VSS.n6505 VSS.n6504 2.2505
R4693 VSS.n6503 VSS.n2398 2.2505
R4694 VSS.n6502 VSS.n6501 2.2505
R4695 VSS.n6500 VSS.n2399 2.2505
R4696 VSS.n6499 VSS.n6498 2.2505
R4697 VSS.n6497 VSS.n2400 2.2505
R4698 VSS.n6496 VSS.n6495 2.2505
R4699 VSS.n6494 VSS.n2401 2.2505
R4700 VSS.n6493 VSS.n6492 2.2505
R4701 VSS.n6491 VSS.n2402 2.2505
R4702 VSS.n6490 VSS.n6489 2.2505
R4703 VSS.n6488 VSS.n2403 2.2505
R4704 VSS.n6487 VSS.n6486 2.2505
R4705 VSS.n6485 VSS.n2404 2.2505
R4706 VSS.n6484 VSS.n6483 2.2505
R4707 VSS.n6482 VSS.n2405 2.2505
R4708 VSS.n6481 VSS.n6480 2.2505
R4709 VSS.n6479 VSS.n2406 2.2505
R4710 VSS.n6478 VSS.n6477 2.2505
R4711 VSS.n6476 VSS.n2407 2.2505
R4712 VSS.n6475 VSS.n6474 2.2505
R4713 VSS.n6473 VSS.n2408 2.2505
R4714 VSS.n6472 VSS.n6471 2.2505
R4715 VSS.n6470 VSS.n2409 2.2505
R4716 VSS.n6469 VSS.n6468 2.2505
R4717 VSS.n6467 VSS.n2410 2.2505
R4718 VSS.n6466 VSS.n6465 2.2505
R4719 VSS.n6464 VSS.n2411 2.2505
R4720 VSS.n6463 VSS.n6462 2.2505
R4721 VSS.n6461 VSS.n2412 2.2505
R4722 VSS.n6460 VSS.n6459 2.2505
R4723 VSS.n6458 VSS.n2413 2.2505
R4724 VSS.n6457 VSS.n6456 2.2505
R4725 VSS.n6455 VSS.n2414 2.2505
R4726 VSS.n6454 VSS.n6453 2.2505
R4727 VSS.n6452 VSS.n2415 2.2505
R4728 VSS.n6451 VSS.n6450 2.2505
R4729 VSS.n6449 VSS.n2416 2.2505
R4730 VSS.n6448 VSS.n6447 2.2505
R4731 VSS.n6446 VSS.n2417 2.2505
R4732 VSS.n6445 VSS.n6444 2.2505
R4733 VSS.n6443 VSS.n2418 2.2505
R4734 VSS.n6442 VSS.n6441 2.2505
R4735 VSS.n6440 VSS.n2419 2.2505
R4736 VSS.n6439 VSS.n6438 2.2505
R4737 VSS.n6437 VSS.n2420 2.2505
R4738 VSS.n6436 VSS.n6435 2.2505
R4739 VSS.n6434 VSS.n2421 2.2505
R4740 VSS.n6433 VSS.n6432 2.2505
R4741 VSS.n6431 VSS.n2422 2.2505
R4742 VSS.n6430 VSS.n6429 2.2505
R4743 VSS.n6428 VSS.n2423 2.2505
R4744 VSS.n6427 VSS.n6426 2.2505
R4745 VSS.n6425 VSS.n2424 2.2505
R4746 VSS.n6424 VSS.n6423 2.2505
R4747 VSS.n6422 VSS.n2425 2.2505
R4748 VSS.n6421 VSS.n6420 2.2505
R4749 VSS.n6419 VSS.n2426 2.2505
R4750 VSS.n6418 VSS.n6417 2.2505
R4751 VSS.n6416 VSS.n2427 2.2505
R4752 VSS.n6415 VSS.n6414 2.2505
R4753 VSS.n6413 VSS.n2428 2.2505
R4754 VSS.n6412 VSS.n6411 2.2505
R4755 VSS.n6410 VSS.n2429 2.2505
R4756 VSS.n6409 VSS.n6408 2.2505
R4757 VSS.n6407 VSS.n2430 2.2505
R4758 VSS.n6406 VSS.n6405 2.2505
R4759 VSS.n6404 VSS.n2431 2.2505
R4760 VSS.n6403 VSS.n6402 2.2505
R4761 VSS.n6401 VSS.n2432 2.2505
R4762 VSS.n6400 VSS.n6399 2.2505
R4763 VSS.n6398 VSS.n2433 2.2505
R4764 VSS.n6397 VSS.n6396 2.2505
R4765 VSS.n6395 VSS.n2434 2.2505
R4766 VSS.n6394 VSS.n6393 2.2505
R4767 VSS.n6392 VSS.n2435 2.2505
R4768 VSS.n6391 VSS.n6390 2.2505
R4769 VSS.n6389 VSS.n2436 2.2505
R4770 VSS.n6388 VSS.n6387 2.2505
R4771 VSS.n6386 VSS.n2437 2.2505
R4772 VSS.n6385 VSS.n6384 2.2505
R4773 VSS.n6383 VSS.n2438 2.2505
R4774 VSS.n6382 VSS.n6381 2.2505
R4775 VSS.n6380 VSS.n2439 2.2505
R4776 VSS.n6379 VSS.n6378 2.2505
R4777 VSS.n6377 VSS.n2440 2.2505
R4778 VSS.n6376 VSS.n6375 2.2505
R4779 VSS.n6374 VSS.n2441 2.2505
R4780 VSS.n6373 VSS.n6372 2.2505
R4781 VSS.n6371 VSS.n2442 2.2505
R4782 VSS.n6370 VSS.n6369 2.2505
R4783 VSS.n6368 VSS.n2443 2.2505
R4784 VSS.n6367 VSS.n6366 2.2505
R4785 VSS.n6365 VSS.n2444 2.2505
R4786 VSS.n6364 VSS.n6363 2.2505
R4787 VSS.n6362 VSS.n2445 2.2505
R4788 VSS.n6361 VSS.n6360 2.2505
R4789 VSS.n6359 VSS.n2446 2.2505
R4790 VSS.n6358 VSS.n6357 2.2505
R4791 VSS.n6356 VSS.n2447 2.2505
R4792 VSS.n6355 VSS.n6354 2.2505
R4793 VSS.n6353 VSS.n2448 2.2505
R4794 VSS.n6352 VSS.n6351 2.2505
R4795 VSS.n6350 VSS.n2449 2.2505
R4796 VSS.n6349 VSS.n6348 2.2505
R4797 VSS.n6347 VSS.n2450 2.2505
R4798 VSS.n6346 VSS.n6345 2.2505
R4799 VSS.n6344 VSS.n2451 2.2505
R4800 VSS.n6343 VSS.n6342 2.2505
R4801 VSS.n6341 VSS.n2452 2.2505
R4802 VSS.n6340 VSS.n6339 2.2505
R4803 VSS.n6338 VSS.n2453 2.2505
R4804 VSS.n6337 VSS.n6336 2.2505
R4805 VSS.n6335 VSS.n2454 2.2505
R4806 VSS.n6334 VSS.n6333 2.2505
R4807 VSS.n6332 VSS.n2455 2.2505
R4808 VSS.n6331 VSS.n6330 2.2505
R4809 VSS.n6329 VSS.n2456 2.2505
R4810 VSS.n6328 VSS.n6327 2.2505
R4811 VSS.n6326 VSS.n2457 2.2505
R4812 VSS.n6325 VSS.n6324 2.2505
R4813 VSS.n6323 VSS.n2458 2.2505
R4814 VSS.n6322 VSS.n6321 2.2505
R4815 VSS.n6320 VSS.n2459 2.2505
R4816 VSS.n6319 VSS.n6318 2.2505
R4817 VSS.n6317 VSS.n2460 2.2505
R4818 VSS.n6316 VSS.n6315 2.2505
R4819 VSS.n6314 VSS.n2461 2.2505
R4820 VSS.n6313 VSS.n6312 2.2505
R4821 VSS.n6311 VSS.n2462 2.2505
R4822 VSS.n6310 VSS.n6309 2.2505
R4823 VSS.n6308 VSS.n2463 2.2505
R4824 VSS.n6307 VSS.n6306 2.2505
R4825 VSS.n6305 VSS.n2464 2.2505
R4826 VSS.n6304 VSS.n6303 2.2505
R4827 VSS.n6302 VSS.n2465 2.2505
R4828 VSS.n6301 VSS.n6300 2.2505
R4829 VSS.n6299 VSS.n2466 2.2505
R4830 VSS.n6298 VSS.n6297 2.2505
R4831 VSS.n6296 VSS.n2467 2.2505
R4832 VSS.n6295 VSS.n6294 2.2505
R4833 VSS.n6293 VSS.n2468 2.2505
R4834 VSS.n6292 VSS.n6291 2.2505
R4835 VSS.n6290 VSS.n2469 2.2505
R4836 VSS.n6289 VSS.n6288 2.2505
R4837 VSS.n6287 VSS.n2470 2.2505
R4838 VSS.n6286 VSS.n6285 2.2505
R4839 VSS.n6284 VSS.n2471 2.2505
R4840 VSS.n6283 VSS.n6282 2.2505
R4841 VSS.n6281 VSS.n2472 2.2505
R4842 VSS.n6280 VSS.n6279 2.2505
R4843 VSS.n6278 VSS.n2473 2.2505
R4844 VSS.n6277 VSS.n6276 2.2505
R4845 VSS.n6275 VSS.n2474 2.2505
R4846 VSS.n6274 VSS.n6273 2.2505
R4847 VSS.n6272 VSS.n2475 2.2505
R4848 VSS.n6271 VSS.n6270 2.2505
R4849 VSS.n6269 VSS.n2476 2.2505
R4850 VSS.n6268 VSS.n6267 2.2505
R4851 VSS.n6266 VSS.n2477 2.2505
R4852 VSS.n6265 VSS.n6264 2.2505
R4853 VSS.n6263 VSS.n2478 2.2505
R4854 VSS.n6262 VSS.n6261 2.2505
R4855 VSS.n6260 VSS.n2479 2.2505
R4856 VSS.n6259 VSS.n6258 2.2505
R4857 VSS.n6257 VSS.n2480 2.2505
R4858 VSS.n6256 VSS.n6255 2.2505
R4859 VSS.n6254 VSS.n2481 2.2505
R4860 VSS.n6253 VSS.n6252 2.2505
R4861 VSS.n6251 VSS.n2482 2.2505
R4862 VSS.n6250 VSS.n6249 2.2505
R4863 VSS.n6248 VSS.n2483 2.2505
R4864 VSS.n6247 VSS.n6246 2.2505
R4865 VSS.n6245 VSS.n2484 2.2505
R4866 VSS.n6244 VSS.n6243 2.2505
R4867 VSS.n6242 VSS.n2485 2.2505
R4868 VSS.n6241 VSS.n6240 2.2505
R4869 VSS.n6239 VSS.n2486 2.2505
R4870 VSS.n6238 VSS.n6237 2.2505
R4871 VSS.n6236 VSS.n2487 2.2505
R4872 VSS.n6235 VSS.n6234 2.2505
R4873 VSS.n6233 VSS.n2488 2.2505
R4874 VSS.n6232 VSS.n6231 2.2505
R4875 VSS.n6230 VSS.n2489 2.2505
R4876 VSS.n6229 VSS.n6228 2.2505
R4877 VSS.n6227 VSS.n2490 2.2505
R4878 VSS.n6226 VSS.n6225 2.2505
R4879 VSS.n6224 VSS.n2491 2.2505
R4880 VSS.n6223 VSS.n6222 2.2505
R4881 VSS.n6221 VSS.n2492 2.2505
R4882 VSS.n6220 VSS.n6219 2.2505
R4883 VSS.n6218 VSS.n2493 2.2505
R4884 VSS.n6217 VSS.n6216 2.2505
R4885 VSS.n6215 VSS.n2494 2.2505
R4886 VSS.n6214 VSS.n6213 2.2505
R4887 VSS.n6212 VSS.n2495 2.2505
R4888 VSS.n6211 VSS.n6210 2.2505
R4889 VSS.n6209 VSS.n2496 2.2505
R4890 VSS.n6208 VSS.n6207 2.2505
R4891 VSS.n6206 VSS.n2497 2.2505
R4892 VSS.n6205 VSS.n6204 2.2505
R4893 VSS.n6203 VSS.n2498 2.2505
R4894 VSS.n6202 VSS.n6201 2.2505
R4895 VSS.n6200 VSS.n2499 2.2505
R4896 VSS.n6199 VSS.n6198 2.2505
R4897 VSS.n6197 VSS.n2500 2.2505
R4898 VSS.n6196 VSS.n6195 2.2505
R4899 VSS.n6194 VSS.n2501 2.2505
R4900 VSS.n6193 VSS.n6192 2.2505
R4901 VSS.n6191 VSS.n2502 2.2505
R4902 VSS.n6190 VSS.n6189 2.2505
R4903 VSS.n6188 VSS.n2503 2.2505
R4904 VSS.n6187 VSS.n6186 2.2505
R4905 VSS.n6185 VSS.n2504 2.2505
R4906 VSS.n6184 VSS.n6183 2.2505
R4907 VSS.n6182 VSS.n2505 2.2505
R4908 VSS.n6181 VSS.n6180 2.2505
R4909 VSS.n6179 VSS.n2506 2.2505
R4910 VSS.n6178 VSS.n6177 2.2505
R4911 VSS.n6176 VSS.n2507 2.2505
R4912 VSS.n6175 VSS.n6174 2.2505
R4913 VSS.n6173 VSS.n2508 2.2505
R4914 VSS.n6172 VSS.n6171 2.2505
R4915 VSS.n6170 VSS.n2509 2.2505
R4916 VSS.n6169 VSS.n6168 2.2505
R4917 VSS.n6167 VSS.n2510 2.2505
R4918 VSS.n6166 VSS.n6165 2.2505
R4919 VSS.n6164 VSS.n2511 2.2505
R4920 VSS.n6163 VSS.n6162 2.2505
R4921 VSS.n6161 VSS.n2512 2.2505
R4922 VSS.n6160 VSS.n6159 2.2505
R4923 VSS.n6158 VSS.n2513 2.2505
R4924 VSS.n6157 VSS.n6156 2.2505
R4925 VSS.n6155 VSS.n2514 2.2505
R4926 VSS.n6154 VSS.n6153 2.2505
R4927 VSS.n6152 VSS.n2515 2.2505
R4928 VSS.n6151 VSS.n6150 2.2505
R4929 VSS.n6149 VSS.n2516 2.2505
R4930 VSS.n6148 VSS.n6147 2.2505
R4931 VSS.n6146 VSS.n2517 2.2505
R4932 VSS.n6145 VSS.n6144 2.2505
R4933 VSS.n6143 VSS.n2518 2.2505
R4934 VSS.n6142 VSS.n6141 2.2505
R4935 VSS.n6140 VSS.n2519 2.2505
R4936 VSS.n6139 VSS.n6138 2.2505
R4937 VSS.n6137 VSS.n2520 2.2505
R4938 VSS.n6136 VSS.n6135 2.2505
R4939 VSS.n6134 VSS.n2521 2.2505
R4940 VSS.n6133 VSS.n6132 2.2505
R4941 VSS.n6131 VSS.n2522 2.2505
R4942 VSS.n6130 VSS.n6129 2.2505
R4943 VSS.n6128 VSS.n2523 2.2505
R4944 VSS.n6127 VSS.n6126 2.2505
R4945 VSS.n6125 VSS.n2524 2.2505
R4946 VSS.n6124 VSS.n6123 2.2505
R4947 VSS.n6122 VSS.n2525 2.2505
R4948 VSS.n6121 VSS.n6120 2.2505
R4949 VSS.n6119 VSS.n2526 2.2505
R4950 VSS.n6118 VSS.n6117 2.2505
R4951 VSS.n6116 VSS.n2527 2.2505
R4952 VSS.n6115 VSS.n6114 2.2505
R4953 VSS.n6113 VSS.n2528 2.2505
R4954 VSS.n6112 VSS.n6111 2.2505
R4955 VSS.n6110 VSS.n2529 2.2505
R4956 VSS.n6109 VSS.n6108 2.2505
R4957 VSS.n6107 VSS.n2530 2.2505
R4958 VSS.n6106 VSS.n6105 2.2505
R4959 VSS.n6104 VSS.n2531 2.2505
R4960 VSS.n6103 VSS.n6102 2.2505
R4961 VSS.n6101 VSS.n2532 2.2505
R4962 VSS.n6100 VSS.n6099 2.2505
R4963 VSS.n6098 VSS.n2533 2.2505
R4964 VSS.n6097 VSS.n6096 2.2505
R4965 VSS.n6095 VSS.n2534 2.2505
R4966 VSS.n6094 VSS.n6093 2.2505
R4967 VSS.n6092 VSS.n2535 2.2505
R4968 VSS.n6091 VSS.n6090 2.2505
R4969 VSS.n6089 VSS.n2536 2.2505
R4970 VSS.n6088 VSS.n6087 2.2505
R4971 VSS.n6086 VSS.n2537 2.2505
R4972 VSS.n6085 VSS.n6084 2.2505
R4973 VSS.n6083 VSS.n2538 2.2505
R4974 VSS.n6082 VSS.n6081 2.2505
R4975 VSS.n6080 VSS.n2539 2.2505
R4976 VSS.n6079 VSS.n6078 2.2505
R4977 VSS.n6077 VSS.n2540 2.2505
R4978 VSS.n6076 VSS.n6075 2.2505
R4979 VSS.n6074 VSS.n2541 2.2505
R4980 VSS.n6073 VSS.n6072 2.2505
R4981 VSS.n6071 VSS.n2542 2.2505
R4982 VSS.n6070 VSS.n6069 2.2505
R4983 VSS.n6068 VSS.n2543 2.2505
R4984 VSS.n6067 VSS.n6066 2.2505
R4985 VSS.n6065 VSS.n2544 2.2505
R4986 VSS.n6064 VSS.n6063 2.2505
R4987 VSS.n6062 VSS.n2545 2.2505
R4988 VSS.n6061 VSS.n6060 2.2505
R4989 VSS.n6059 VSS.n2546 2.2505
R4990 VSS.n6058 VSS.n6057 2.2505
R4991 VSS.n6056 VSS.n2547 2.2505
R4992 VSS.n6055 VSS.n6054 2.2505
R4993 VSS.n6053 VSS.n2548 2.2505
R4994 VSS.n6052 VSS.n6051 2.2505
R4995 VSS.n6050 VSS.n2549 2.2505
R4996 VSS.n6049 VSS.n6048 2.2505
R4997 VSS.n6047 VSS.n2550 2.2505
R4998 VSS.n6046 VSS.n6045 2.2505
R4999 VSS.n6044 VSS.n2551 2.2505
R5000 VSS.n6043 VSS.n6042 2.2505
R5001 VSS.n6041 VSS.n2552 2.2505
R5002 VSS.n6040 VSS.n6039 2.2505
R5003 VSS.n6038 VSS.n2553 2.2505
R5004 VSS.n6037 VSS.n6036 2.2505
R5005 VSS.n6035 VSS.n2554 2.2505
R5006 VSS.n6034 VSS.n6033 2.2505
R5007 VSS.n6032 VSS.n2555 2.2505
R5008 VSS.n6031 VSS.n6030 2.2505
R5009 VSS.n6029 VSS.n2556 2.2505
R5010 VSS.n6028 VSS.n6027 2.2505
R5011 VSS.n6026 VSS.n2557 2.2505
R5012 VSS.n6025 VSS.n6024 2.2505
R5013 VSS.n6023 VSS.n2558 2.2505
R5014 VSS.n6022 VSS.n6021 2.2505
R5015 VSS.n6020 VSS.n2559 2.2505
R5016 VSS.n6019 VSS.n6018 2.2505
R5017 VSS.n6017 VSS.n2560 2.2505
R5018 VSS.n6016 VSS.n6015 2.2505
R5019 VSS.n6014 VSS.n2561 2.2505
R5020 VSS.n6013 VSS.n6012 2.2505
R5021 VSS.n6011 VSS.n2562 2.2505
R5022 VSS.n6010 VSS.n6009 2.2505
R5023 VSS.n6008 VSS.n2563 2.2505
R5024 VSS.n6007 VSS.n6006 2.2505
R5025 VSS.n6005 VSS.n2564 2.2505
R5026 VSS.n6004 VSS.n6003 2.2505
R5027 VSS.n6002 VSS.n2565 2.2505
R5028 VSS.n6001 VSS.n6000 2.2505
R5029 VSS.n5999 VSS.n2566 2.2505
R5030 VSS.n5998 VSS.n5997 2.2505
R5031 VSS.n5996 VSS.n2567 2.2505
R5032 VSS.n5995 VSS.n5994 2.2505
R5033 VSS.n5993 VSS.n2568 2.2505
R5034 VSS.n5992 VSS.n5991 2.2505
R5035 VSS.n5990 VSS.n2569 2.2505
R5036 VSS.n5989 VSS.n5988 2.2505
R5037 VSS.n5987 VSS.n2570 2.2505
R5038 VSS.n5986 VSS.n5985 2.2505
R5039 VSS.n5984 VSS.n2571 2.2505
R5040 VSS.n5983 VSS.n5982 2.2505
R5041 VSS.n5981 VSS.n2572 2.2505
R5042 VSS.n5980 VSS.n5979 2.2505
R5043 VSS.n5978 VSS.n2573 2.2505
R5044 VSS.n5977 VSS.n5976 2.2505
R5045 VSS.n5975 VSS.n2574 2.2505
R5046 VSS.n5974 VSS.n5973 2.2505
R5047 VSS.n5972 VSS.n2575 2.2505
R5048 VSS.n5971 VSS.n5970 2.2505
R5049 VSS.n5969 VSS.n2576 2.2505
R5050 VSS.n5968 VSS.n5967 2.2505
R5051 VSS.n5966 VSS.n2577 2.2505
R5052 VSS.n5965 VSS.n5964 2.2505
R5053 VSS.n5963 VSS.n2578 2.2505
R5054 VSS.n5962 VSS.n5961 2.2505
R5055 VSS.n5960 VSS.n2579 2.2505
R5056 VSS.n5959 VSS.n5958 2.2505
R5057 VSS.n5957 VSS.n2580 2.2505
R5058 VSS.n5956 VSS.n5955 2.2505
R5059 VSS.n5954 VSS.n2581 2.2505
R5060 VSS.n5953 VSS.n5952 2.2505
R5061 VSS.n5951 VSS.n2582 2.2505
R5062 VSS.n5950 VSS.n5949 2.2505
R5063 VSS.n5948 VSS.n2583 2.2505
R5064 VSS.n5947 VSS.n5946 2.2505
R5065 VSS.n5945 VSS.n2584 2.2505
R5066 VSS.n5944 VSS.n5943 2.2505
R5067 VSS.n5942 VSS.n2585 2.2505
R5068 VSS.n5941 VSS.n5940 2.2505
R5069 VSS.n5939 VSS.n2586 2.2505
R5070 VSS.n5938 VSS.n5937 2.2505
R5071 VSS.n5936 VSS.n2587 2.2505
R5072 VSS.n5935 VSS.n5934 2.2505
R5073 VSS.n5933 VSS.n2588 2.2505
R5074 VSS.n5932 VSS.n5931 2.2505
R5075 VSS.n5930 VSS.n2589 2.2505
R5076 VSS.n5929 VSS.n5928 2.2505
R5077 VSS.n5927 VSS.n2590 2.2505
R5078 VSS.n5926 VSS.n5925 2.2505
R5079 VSS.n5924 VSS.n2591 2.2505
R5080 VSS.n5923 VSS.n5922 2.2505
R5081 VSS.n5921 VSS.n2592 2.2505
R5082 VSS.n5920 VSS.n5919 2.2505
R5083 VSS.n5918 VSS.n2593 2.2505
R5084 VSS.n5917 VSS.n5916 2.2505
R5085 VSS.n5915 VSS.n2594 2.2505
R5086 VSS.n5914 VSS.n5913 2.2505
R5087 VSS.n5912 VSS.n2595 2.2505
R5088 VSS.n5911 VSS.n5910 2.2505
R5089 VSS.n5909 VSS.n2596 2.2505
R5090 VSS.n5908 VSS.n5907 2.2505
R5091 VSS.n5906 VSS.n2597 2.2505
R5092 VSS.n5905 VSS.n5904 2.2505
R5093 VSS.n5903 VSS.n2598 2.2505
R5094 VSS.n5902 VSS.n5901 2.2505
R5095 VSS.n5900 VSS.n2599 2.2505
R5096 VSS.n5899 VSS.n5898 2.2505
R5097 VSS.n5897 VSS.n2600 2.2505
R5098 VSS.n5896 VSS.n5895 2.2505
R5099 VSS.n5894 VSS.n2601 2.2505
R5100 VSS.n5893 VSS.n5892 2.2505
R5101 VSS.n5891 VSS.n2602 2.2505
R5102 VSS.n5890 VSS.n5889 2.2505
R5103 VSS.n5888 VSS.n2603 2.2505
R5104 VSS.n5887 VSS.n5886 2.2505
R5105 VSS.n5885 VSS.n2604 2.2505
R5106 VSS.n5884 VSS.n5883 2.2505
R5107 VSS.n5882 VSS.n2605 2.2505
R5108 VSS.n5881 VSS.n5880 2.2505
R5109 VSS.n5879 VSS.n2606 2.2505
R5110 VSS.n5878 VSS.n5877 2.2505
R5111 VSS.n5876 VSS.n2607 2.2505
R5112 VSS.n5875 VSS.n5874 2.2505
R5113 VSS.n5873 VSS.n2608 2.2505
R5114 VSS.n5872 VSS.n5871 2.2505
R5115 VSS.n5870 VSS.n2609 2.2505
R5116 VSS.n5869 VSS.n5868 2.2505
R5117 VSS.n5867 VSS.n2610 2.2505
R5118 VSS.n5866 VSS.n5865 2.2505
R5119 VSS.n5864 VSS.n2611 2.2505
R5120 VSS.n5863 VSS.n5862 2.2505
R5121 VSS.n5861 VSS.n2612 2.2505
R5122 VSS.n5860 VSS.n5859 2.2505
R5123 VSS.n5858 VSS.n2613 2.2505
R5124 VSS.n5857 VSS.n5856 2.2505
R5125 VSS.n5855 VSS.n2614 2.2505
R5126 VSS.n5854 VSS.n5853 2.2505
R5127 VSS.n5852 VSS.n2615 2.2505
R5128 VSS.n5851 VSS.n5850 2.2505
R5129 VSS.n5849 VSS.n2616 2.2505
R5130 VSS.n5848 VSS.n5847 2.2505
R5131 VSS.n5846 VSS.n2617 2.2505
R5132 VSS.n5845 VSS.n5844 2.2505
R5133 VSS.n5843 VSS.n2618 2.2505
R5134 VSS.n5842 VSS.n5841 2.2505
R5135 VSS.n5840 VSS.n2619 2.2505
R5136 VSS.n5839 VSS.n5838 2.2505
R5137 VSS.n5837 VSS.n2620 2.2505
R5138 VSS.n5836 VSS.n5835 2.2505
R5139 VSS.n5834 VSS.n2621 2.2505
R5140 VSS.n5833 VSS.n5832 2.2505
R5141 VSS.n5831 VSS.n2622 2.2505
R5142 VSS.n5830 VSS.n5829 2.2505
R5143 VSS.n5828 VSS.n2623 2.2505
R5144 VSS.n5827 VSS.n5826 2.2505
R5145 VSS.n5825 VSS.n2624 2.2505
R5146 VSS.n5824 VSS.n5823 2.2505
R5147 VSS.n5822 VSS.n2625 2.2505
R5148 VSS.n5821 VSS.n5820 2.2505
R5149 VSS.n5819 VSS.n2626 2.2505
R5150 VSS.n5818 VSS.n5817 2.2505
R5151 VSS.n5816 VSS.n2627 2.2505
R5152 VSS.n5815 VSS.n5814 2.2505
R5153 VSS.n5813 VSS.n2628 2.2505
R5154 VSS.n5812 VSS.n5811 2.2505
R5155 VSS.n5810 VSS.n2629 2.2505
R5156 VSS.n5809 VSS.n5808 2.2505
R5157 VSS.n5807 VSS.n2630 2.2505
R5158 VSS.n5806 VSS.n5805 2.2505
R5159 VSS.n5804 VSS.n2631 2.2505
R5160 VSS.n5803 VSS.n5802 2.2505
R5161 VSS.n5801 VSS.n2632 2.2505
R5162 VSS.n5800 VSS.n5799 2.2505
R5163 VSS.n5798 VSS.n2633 2.2505
R5164 VSS.n5797 VSS.n5796 2.2505
R5165 VSS.n5795 VSS.n2634 2.2505
R5166 VSS.n5794 VSS.n5793 2.2505
R5167 VSS.n5792 VSS.n2635 2.2505
R5168 VSS.n5791 VSS.n5790 2.2505
R5169 VSS.n5789 VSS.n2636 2.2505
R5170 VSS.n5788 VSS.n5787 2.2505
R5171 VSS.n5786 VSS.n2637 2.2505
R5172 VSS.n5785 VSS.n5784 2.2505
R5173 VSS.n5783 VSS.n2638 2.2505
R5174 VSS.n5782 VSS.n5781 2.2505
R5175 VSS.n5780 VSS.n2639 2.2505
R5176 VSS.n5779 VSS.n5778 2.2505
R5177 VSS.n5777 VSS.n2640 2.2505
R5178 VSS.n5776 VSS.n5775 2.2505
R5179 VSS.n5774 VSS.n2641 2.2505
R5180 VSS.n5773 VSS.n5772 2.2505
R5181 VSS.n5771 VSS.n2642 2.2505
R5182 VSS.n5770 VSS.n5769 2.2505
R5183 VSS.n5768 VSS.n2643 2.2505
R5184 VSS.n5767 VSS.n5766 2.2505
R5185 VSS.n5765 VSS.n2644 2.2505
R5186 VSS.n5764 VSS.n5763 2.2505
R5187 VSS.n5762 VSS.n2645 2.2505
R5188 VSS.n5761 VSS.n5760 2.2505
R5189 VSS.n5759 VSS.n2646 2.2505
R5190 VSS.n5758 VSS.n5757 2.2505
R5191 VSS.n5756 VSS.n2647 2.2505
R5192 VSS.n5755 VSS.n5754 2.2505
R5193 VSS.n5753 VSS.n2648 2.2505
R5194 VSS.n5752 VSS.n5751 2.2505
R5195 VSS.n5750 VSS.n2649 2.2505
R5196 VSS.n5749 VSS.n5748 2.2505
R5197 VSS.n5747 VSS.n2650 2.2505
R5198 VSS.n5746 VSS.n5745 2.2505
R5199 VSS.n5744 VSS.n2651 2.2505
R5200 VSS.n5743 VSS.n5742 2.2505
R5201 VSS.n5741 VSS.n2652 2.2505
R5202 VSS.n5740 VSS.n5739 2.2505
R5203 VSS.n5738 VSS.n2653 2.2505
R5204 VSS.n5737 VSS.n5736 2.2505
R5205 VSS.n5735 VSS.n2654 2.2505
R5206 VSS.n5734 VSS.n5733 2.2505
R5207 VSS.n5732 VSS.n2655 2.2505
R5208 VSS.n5731 VSS.n5730 2.2505
R5209 VSS.n5729 VSS.n2656 2.2505
R5210 VSS.n5728 VSS.n5727 2.2505
R5211 VSS.n5726 VSS.n2657 2.2505
R5212 VSS.n5725 VSS.n5724 2.2505
R5213 VSS.n5723 VSS.n2658 2.2505
R5214 VSS.n5722 VSS.n5721 2.2505
R5215 VSS.n5720 VSS.n2659 2.2505
R5216 VSS.n5719 VSS.n5718 2.2505
R5217 VSS.n5717 VSS.n2660 2.2505
R5218 VSS.n5716 VSS.n5715 2.2505
R5219 VSS.n5714 VSS.n2661 2.2505
R5220 VSS.n5713 VSS.n5712 2.2505
R5221 VSS.n5711 VSS.n2662 2.2505
R5222 VSS.n5710 VSS.n5709 2.2505
R5223 VSS.n5708 VSS.n2663 2.2505
R5224 VSS.n5707 VSS.n5706 2.2505
R5225 VSS.n5705 VSS.n2664 2.2505
R5226 VSS.n5704 VSS.n5703 2.2505
R5227 VSS.n5702 VSS.n2665 2.2505
R5228 VSS.n5701 VSS.n5700 2.2505
R5229 VSS.n5699 VSS.n2666 2.2505
R5230 VSS.n5698 VSS.n5697 2.2505
R5231 VSS.n5696 VSS.n2667 2.2505
R5232 VSS.n5695 VSS.n5694 2.2505
R5233 VSS.n5693 VSS.n2668 2.2505
R5234 VSS.n5692 VSS.n5691 2.2505
R5235 VSS.n5690 VSS.n2669 2.2505
R5236 VSS.n5689 VSS.n5688 2.2505
R5237 VSS.n5687 VSS.n2670 2.2505
R5238 VSS.n5686 VSS.n5685 2.2505
R5239 VSS.n5684 VSS.n2671 2.2505
R5240 VSS.n5683 VSS.n5682 2.2505
R5241 VSS.n5681 VSS.n2672 2.2505
R5242 VSS.n5680 VSS.n5679 2.2505
R5243 VSS.n5678 VSS.n2673 2.2505
R5244 VSS.n5677 VSS.n5676 2.2505
R5245 VSS.n5675 VSS.n2674 2.2505
R5246 VSS.n5674 VSS.n5673 2.2505
R5247 VSS.n5672 VSS.n2675 2.2505
R5248 VSS.n5671 VSS.n5670 2.2505
R5249 VSS.n5669 VSS.n2676 2.2505
R5250 VSS.n5668 VSS.n5667 2.2505
R5251 VSS.n5666 VSS.n2677 2.2505
R5252 VSS.n5665 VSS.n5664 2.2505
R5253 VSS.n5663 VSS.n2678 2.2505
R5254 VSS.n5662 VSS.n5661 2.2505
R5255 VSS.n5660 VSS.n2679 2.2505
R5256 VSS.n5659 VSS.n5658 2.2505
R5257 VSS.n5657 VSS.n2680 2.2505
R5258 VSS.n5656 VSS.n5655 2.2505
R5259 VSS.n5654 VSS.n2681 2.2505
R5260 VSS.n5653 VSS.n5652 2.2505
R5261 VSS.n5651 VSS.n2682 2.2505
R5262 VSS.n5650 VSS.n5649 2.2505
R5263 VSS.n5648 VSS.n2683 2.2505
R5264 VSS.n5647 VSS.n5646 2.2505
R5265 VSS.n5645 VSS.n2684 2.2505
R5266 VSS.n5644 VSS.n5643 2.2505
R5267 VSS.n5642 VSS.n2685 2.2505
R5268 VSS.n5641 VSS.n5640 2.2505
R5269 VSS.n5639 VSS.n2686 2.2505
R5270 VSS.n5638 VSS.n5637 2.2505
R5271 VSS.n5636 VSS.n2687 2.2505
R5272 VSS.n5635 VSS.n5634 2.2505
R5273 VSS.n5633 VSS.n2688 2.2505
R5274 VSS.n5632 VSS.n5631 2.2505
R5275 VSS.n5630 VSS.n2689 2.2505
R5276 VSS.n5629 VSS.n5628 2.2505
R5277 VSS.n5627 VSS.n2690 2.2505
R5278 VSS.n5626 VSS.n5625 2.2505
R5279 VSS.n5624 VSS.n2691 2.2505
R5280 VSS.n5623 VSS.n5622 2.2505
R5281 VSS.n5621 VSS.n2692 2.2505
R5282 VSS.n5620 VSS.n5619 2.2505
R5283 VSS.n5618 VSS.n2693 2.2505
R5284 VSS.n5617 VSS.n5616 2.2505
R5285 VSS.n5615 VSS.n2694 2.2505
R5286 VSS.n5614 VSS.n5613 2.2505
R5287 VSS.n5612 VSS.n2695 2.2505
R5288 VSS.n5611 VSS.n5610 2.2505
R5289 VSS.n5609 VSS.n2696 2.2505
R5290 VSS.n5608 VSS.n5607 2.2505
R5291 VSS.n5606 VSS.n2697 2.2505
R5292 VSS.n5605 VSS.n5604 2.2505
R5293 VSS.n5603 VSS.n2698 2.2505
R5294 VSS.n5602 VSS.n5601 2.2505
R5295 VSS.n5600 VSS.n2699 2.2505
R5296 VSS.n5599 VSS.n5598 2.2505
R5297 VSS.n5597 VSS.n2700 2.2505
R5298 VSS.n5596 VSS.n5595 2.2505
R5299 VSS.n5594 VSS.n2701 2.2505
R5300 VSS.n5593 VSS.n5592 2.2505
R5301 VSS.n5591 VSS.n2702 2.2505
R5302 VSS.n5590 VSS.n5589 2.2505
R5303 VSS.n5588 VSS.n2703 2.2505
R5304 VSS.n5587 VSS.n5586 2.2505
R5305 VSS.n5585 VSS.n2704 2.2505
R5306 VSS.n5584 VSS.n5583 2.2505
R5307 VSS.n5582 VSS.n2705 2.2505
R5308 VSS.n5581 VSS.n5580 2.2505
R5309 VSS.n5579 VSS.n2706 2.2505
R5310 VSS.n5578 VSS.n5577 2.2505
R5311 VSS.n5576 VSS.n2707 2.2505
R5312 VSS.n5575 VSS.n5574 2.2505
R5313 VSS.n5573 VSS.n2708 2.2505
R5314 VSS.n5572 VSS.n5571 2.2505
R5315 VSS.n5570 VSS.n2709 2.2505
R5316 VSS.n5569 VSS.n5568 2.2505
R5317 VSS.n5567 VSS.n2710 2.2505
R5318 VSS.n5566 VSS.n5565 2.2505
R5319 VSS.n5564 VSS.n2711 2.2505
R5320 VSS.n5563 VSS.n5562 2.2505
R5321 VSS.n5561 VSS.n2712 2.2505
R5322 VSS.n5560 VSS.n5559 2.2505
R5323 VSS.n5558 VSS.n2713 2.2505
R5324 VSS.n5557 VSS.n5556 2.2505
R5325 VSS.n5555 VSS.n2714 2.2505
R5326 VSS.n5554 VSS.n5553 2.2505
R5327 VSS.n5552 VSS.n2715 2.2505
R5328 VSS.n5551 VSS.n5550 2.2505
R5329 VSS.n5549 VSS.n2716 2.2505
R5330 VSS.n5548 VSS.n5547 2.2505
R5331 VSS.n5546 VSS.n2717 2.2505
R5332 VSS.n5545 VSS.n5544 2.2505
R5333 VSS.n5543 VSS.n2718 2.2505
R5334 VSS.n5542 VSS.n5541 2.2505
R5335 VSS.n5540 VSS.n2719 2.2505
R5336 VSS.n5539 VSS.n5538 2.2505
R5337 VSS.n5537 VSS.n2720 2.2505
R5338 VSS.n5536 VSS.n5535 2.2505
R5339 VSS.n5534 VSS.n2721 2.2505
R5340 VSS.n5533 VSS.n5532 2.2505
R5341 VSS.n5531 VSS.n2722 2.2505
R5342 VSS.n5530 VSS.n5529 2.2505
R5343 VSS.n5528 VSS.n2723 2.2505
R5344 VSS.n5527 VSS.n5526 2.2505
R5345 VSS.n5525 VSS.n2724 2.2505
R5346 VSS.n5524 VSS.n5523 2.2505
R5347 VSS.n5522 VSS.n2725 2.2505
R5348 VSS.n5521 VSS.n5520 2.2505
R5349 VSS.n5519 VSS.n2726 2.2505
R5350 VSS.n5518 VSS.n5517 2.2505
R5351 VSS.n5516 VSS.n2727 2.2505
R5352 VSS.n5515 VSS.n5514 2.2505
R5353 VSS.n5513 VSS.n2728 2.2505
R5354 VSS.n5512 VSS.n5511 2.2505
R5355 VSS.n5510 VSS.n2729 2.2505
R5356 VSS.n5509 VSS.n5508 2.2505
R5357 VSS.n5507 VSS.n2730 2.2505
R5358 VSS.n5506 VSS.n5505 2.2505
R5359 VSS.n5504 VSS.n2731 2.2505
R5360 VSS.n5503 VSS.n5502 2.2505
R5361 VSS.n5501 VSS.n2732 2.2505
R5362 VSS.n5500 VSS.n5499 2.2505
R5363 VSS.n5498 VSS.n2733 2.2505
R5364 VSS.n5497 VSS.n5496 2.2505
R5365 VSS.n5495 VSS.n2734 2.2505
R5366 VSS.n5494 VSS.n5493 2.2505
R5367 VSS.n5492 VSS.n2735 2.2505
R5368 VSS.n5491 VSS.n5490 2.2505
R5369 VSS.n5489 VSS.n2736 2.2505
R5370 VSS.n5488 VSS.n5487 2.2505
R5371 VSS.n5486 VSS.n2737 2.2505
R5372 VSS.n5485 VSS.n5484 2.2505
R5373 VSS.n5483 VSS.n2738 2.2505
R5374 VSS.n5482 VSS.n5481 2.2505
R5375 VSS.n5480 VSS.n2739 2.2505
R5376 VSS.n5479 VSS.n5478 2.2505
R5377 VSS.n5477 VSS.n2740 2.2505
R5378 VSS.n5476 VSS.n5475 2.2505
R5379 VSS.n5474 VSS.n2741 2.2505
R5380 VSS.n5473 VSS.n5472 2.2505
R5381 VSS.n5471 VSS.n2742 2.2505
R5382 VSS.n5470 VSS.n5469 2.2505
R5383 VSS.n6908 VSS.n2263 2.2505
R5384 VSS.n6910 VSS.n6909 2.2505
R5385 VSS.n6911 VSS.n2262 2.2505
R5386 VSS.n6913 VSS.n6912 2.2505
R5387 VSS.n6914 VSS.n2261 2.2505
R5388 VSS.n6916 VSS.n6915 2.2505
R5389 VSS.n6917 VSS.n2260 2.2505
R5390 VSS.n6919 VSS.n6918 2.2505
R5391 VSS.n6920 VSS.n2259 2.2505
R5392 VSS.n6922 VSS.n6921 2.2505
R5393 VSS.n6923 VSS.n2258 2.2505
R5394 VSS.n6925 VSS.n6924 2.2505
R5395 VSS.n6926 VSS.n2257 2.2505
R5396 VSS.n6928 VSS.n6927 2.2505
R5397 VSS.n6929 VSS.n2256 2.2505
R5398 VSS.n6931 VSS.n6930 2.2505
R5399 VSS.n6932 VSS.n2255 2.2505
R5400 VSS.n6934 VSS.n6933 2.2505
R5401 VSS.n6935 VSS.n2254 2.2505
R5402 VSS.n6937 VSS.n6936 2.2505
R5403 VSS.n6938 VSS.n2253 2.2505
R5404 VSS.n6940 VSS.n6939 2.2505
R5405 VSS.n6941 VSS.n2252 2.2505
R5406 VSS.n6943 VSS.n6942 2.2505
R5407 VSS.n6944 VSS.n2251 2.2505
R5408 VSS.n6946 VSS.n6945 2.2505
R5409 VSS.n6947 VSS.n2250 2.2505
R5410 VSS.n6949 VSS.n6948 2.2505
R5411 VSS.n6950 VSS.n2249 2.2505
R5412 VSS.n6952 VSS.n6951 2.2505
R5413 VSS.n6953 VSS.n2248 2.2505
R5414 VSS.n6955 VSS.n6954 2.2505
R5415 VSS.n6956 VSS.n2247 2.2505
R5416 VSS.n6958 VSS.n6957 2.2505
R5417 VSS.n6959 VSS.n2246 2.2505
R5418 VSS.n6961 VSS.n6960 2.2505
R5419 VSS.n6962 VSS.n2245 2.2505
R5420 VSS.n6964 VSS.n6963 2.2505
R5421 VSS.n6965 VSS.n2244 2.2505
R5422 VSS.n6967 VSS.n6966 2.2505
R5423 VSS.n6968 VSS.n2243 2.2505
R5424 VSS.n6970 VSS.n6969 2.2505
R5425 VSS.n6971 VSS.n2242 2.2505
R5426 VSS.n6973 VSS.n6972 2.2505
R5427 VSS.n6974 VSS.n2241 2.2505
R5428 VSS.n6976 VSS.n6975 2.2505
R5429 VSS.n6977 VSS.n2240 2.2505
R5430 VSS.n6979 VSS.n6978 2.2505
R5431 VSS.n6980 VSS.n2239 2.2505
R5432 VSS.n6982 VSS.n6981 2.2505
R5433 VSS.n6983 VSS.n2238 2.2505
R5434 VSS.n6985 VSS.n6984 2.2505
R5435 VSS.n6986 VSS.n2237 2.2505
R5436 VSS.n6988 VSS.n6987 2.2505
R5437 VSS.n6989 VSS.n2236 2.2505
R5438 VSS.n6991 VSS.n6990 2.2505
R5439 VSS.n6992 VSS.n2235 2.2505
R5440 VSS.n6994 VSS.n6993 2.2505
R5441 VSS.n6995 VSS.n2234 2.2505
R5442 VSS.n6997 VSS.n6996 2.2505
R5443 VSS.n6998 VSS.n2233 2.2505
R5444 VSS.n7000 VSS.n6999 2.2505
R5445 VSS.n7001 VSS.n2232 2.2505
R5446 VSS.n7003 VSS.n7002 2.2505
R5447 VSS.n7004 VSS.n2231 2.2505
R5448 VSS.n7006 VSS.n7005 2.2505
R5449 VSS.n7007 VSS.n2230 2.2505
R5450 VSS.n7009 VSS.n7008 2.2505
R5451 VSS.n7010 VSS.n2229 2.2505
R5452 VSS.n7012 VSS.n7011 2.2505
R5453 VSS.n7013 VSS.n2228 2.2505
R5454 VSS.n7015 VSS.n7014 2.2505
R5455 VSS.n7016 VSS.n2227 2.2505
R5456 VSS.n7018 VSS.n7017 2.2505
R5457 VSS.n7019 VSS.n2226 2.2505
R5458 VSS.n7021 VSS.n7020 2.2505
R5459 VSS.n7022 VSS.n2225 2.2505
R5460 VSS.n7024 VSS.n7023 2.2505
R5461 VSS.n7025 VSS.n2224 2.2505
R5462 VSS.n7027 VSS.n7026 2.2505
R5463 VSS.n7028 VSS.n2223 2.2505
R5464 VSS.n7030 VSS.n7029 2.2505
R5465 VSS.n7031 VSS.n2222 2.2505
R5466 VSS.n7033 VSS.n7032 2.2505
R5467 VSS.n7034 VSS.n2221 2.2505
R5468 VSS.n7036 VSS.n7035 2.2505
R5469 VSS.n7037 VSS.n2220 2.2505
R5470 VSS.n7039 VSS.n7038 2.2505
R5471 VSS.n7040 VSS.n2219 2.2505
R5472 VSS.n7042 VSS.n7041 2.2505
R5473 VSS.n7043 VSS.n2218 2.2505
R5474 VSS.n7045 VSS.n7044 2.2505
R5475 VSS.n7046 VSS.n2217 2.2505
R5476 VSS.n7048 VSS.n7047 2.2505
R5477 VSS.n7049 VSS.n2216 2.2505
R5478 VSS.n7051 VSS.n7050 2.2505
R5479 VSS.n7052 VSS.n2215 2.2505
R5480 VSS.n7054 VSS.n7053 2.2505
R5481 VSS.n7055 VSS.n2214 2.2505
R5482 VSS.n7057 VSS.n7056 2.2505
R5483 VSS.n7058 VSS.n2213 2.2505
R5484 VSS.n7060 VSS.n7059 2.2505
R5485 VSS.n7061 VSS.n2212 2.2505
R5486 VSS.n7063 VSS.n7062 2.2505
R5487 VSS.n7064 VSS.n2211 2.2505
R5488 VSS.n7066 VSS.n7065 2.2505
R5489 VSS.n7067 VSS.n2210 2.2505
R5490 VSS.n7069 VSS.n7068 2.2505
R5491 VSS.n7070 VSS.n2209 2.2505
R5492 VSS.n7072 VSS.n7071 2.2505
R5493 VSS.n7073 VSS.n2208 2.2505
R5494 VSS.n7075 VSS.n7074 2.2505
R5495 VSS.n7076 VSS.n2207 2.2505
R5496 VSS.n7078 VSS.n7077 2.2505
R5497 VSS.n7079 VSS.n2206 2.2505
R5498 VSS.n7081 VSS.n7080 2.2505
R5499 VSS.n7082 VSS.n2205 2.2505
R5500 VSS.n7084 VSS.n7083 2.2505
R5501 VSS.n7085 VSS.n2204 2.2505
R5502 VSS.n7087 VSS.n7086 2.2505
R5503 VSS.n7088 VSS.n2203 2.2505
R5504 VSS.n7090 VSS.n7089 2.2505
R5505 VSS.n7091 VSS.n2202 2.2505
R5506 VSS.n7093 VSS.n7092 2.2505
R5507 VSS.n7094 VSS.n2201 2.2505
R5508 VSS.n7096 VSS.n7095 2.2505
R5509 VSS.n7097 VSS.n2200 2.2505
R5510 VSS.n7099 VSS.n7098 2.2505
R5511 VSS.n7100 VSS.n2199 2.2505
R5512 VSS.n7102 VSS.n7101 2.2505
R5513 VSS.n7103 VSS.n2198 2.2505
R5514 VSS.n7105 VSS.n7104 2.2505
R5515 VSS.n7106 VSS.n2197 2.2505
R5516 VSS.n7108 VSS.n7107 2.2505
R5517 VSS.n7109 VSS.n2196 2.2505
R5518 VSS.n7111 VSS.n7110 2.2505
R5519 VSS.n7112 VSS.n2195 2.2505
R5520 VSS.n7114 VSS.n7113 2.2505
R5521 VSS.n7115 VSS.n2194 2.2505
R5522 VSS.n7117 VSS.n7116 2.2505
R5523 VSS.n7118 VSS.n2193 2.2505
R5524 VSS.n7120 VSS.n7119 2.2505
R5525 VSS.n7121 VSS.n2192 2.2505
R5526 VSS.n7123 VSS.n7122 2.2505
R5527 VSS.n7124 VSS.n2191 2.2505
R5528 VSS.n7126 VSS.n7125 2.2505
R5529 VSS.n7127 VSS.n2190 2.2505
R5530 VSS.n7129 VSS.n7128 2.2505
R5531 VSS.n7130 VSS.n2189 2.2505
R5532 VSS.n7132 VSS.n7131 2.2505
R5533 VSS.n7133 VSS.n2188 2.2505
R5534 VSS.n7135 VSS.n7134 2.2505
R5535 VSS.n7136 VSS.n2187 2.2505
R5536 VSS.n7138 VSS.n7137 2.2505
R5537 VSS.n7139 VSS.n2186 2.2505
R5538 VSS.n7141 VSS.n7140 2.2505
R5539 VSS.n7142 VSS.n2185 2.2505
R5540 VSS.n7144 VSS.n7143 2.2505
R5541 VSS.n7145 VSS.n2184 2.2505
R5542 VSS.n7147 VSS.n7146 2.2505
R5543 VSS.n7148 VSS.n2183 2.2505
R5544 VSS.n7150 VSS.n7149 2.2505
R5545 VSS.n7151 VSS.n2182 2.2505
R5546 VSS.n7153 VSS.n7152 2.2505
R5547 VSS.n7154 VSS.n2181 2.2505
R5548 VSS.n7156 VSS.n7155 2.2505
R5549 VSS.n7157 VSS.n2180 2.2505
R5550 VSS.n7159 VSS.n7158 2.2505
R5551 VSS.n7160 VSS.n2179 2.2505
R5552 VSS.n7162 VSS.n7161 2.2505
R5553 VSS.n7163 VSS.n2178 2.2505
R5554 VSS.n7165 VSS.n7164 2.2505
R5555 VSS.n7166 VSS.n2177 2.2505
R5556 VSS.n7168 VSS.n7167 2.2505
R5557 VSS.n7169 VSS.n2176 2.2505
R5558 VSS.n7171 VSS.n7170 2.2505
R5559 VSS.n7172 VSS.n2175 2.2505
R5560 VSS.n7174 VSS.n7173 2.2505
R5561 VSS.n7175 VSS.n2174 2.2505
R5562 VSS.n7177 VSS.n7176 2.2505
R5563 VSS.n7178 VSS.n2173 2.2505
R5564 VSS.n7180 VSS.n7179 2.2505
R5565 VSS.n7181 VSS.n2172 2.2505
R5566 VSS.n7183 VSS.n7182 2.2505
R5567 VSS.n7184 VSS.n2171 2.2505
R5568 VSS.n7186 VSS.n7185 2.2505
R5569 VSS.n7187 VSS.n2170 2.2505
R5570 VSS.n7189 VSS.n7188 2.2505
R5571 VSS.n7190 VSS.n2169 2.2505
R5572 VSS.n7192 VSS.n7191 2.2505
R5573 VSS.n7193 VSS.n2168 2.2505
R5574 VSS.n7195 VSS.n7194 2.2505
R5575 VSS.n7196 VSS.n2167 2.2505
R5576 VSS.n7198 VSS.n7197 2.2505
R5577 VSS.n7199 VSS.n2166 2.2505
R5578 VSS.n7201 VSS.n7200 2.2505
R5579 VSS.n7202 VSS.n2165 2.2505
R5580 VSS.n7204 VSS.n7203 2.2505
R5581 VSS.n7205 VSS.n2164 2.2505
R5582 VSS.n7207 VSS.n7206 2.2505
R5583 VSS.n7208 VSS.n2163 2.2505
R5584 VSS.n7210 VSS.n7209 2.2505
R5585 VSS.n7211 VSS.n2162 2.2505
R5586 VSS.n7213 VSS.n7212 2.2505
R5587 VSS.n7214 VSS.n2161 2.2505
R5588 VSS.n7216 VSS.n7215 2.2505
R5589 VSS.n7217 VSS.n2160 2.2505
R5590 VSS.n7219 VSS.n7218 2.2505
R5591 VSS.n7220 VSS.n2159 2.2505
R5592 VSS.n7222 VSS.n7221 2.2505
R5593 VSS.n7223 VSS.n2158 2.2505
R5594 VSS.n7225 VSS.n7224 2.2505
R5595 VSS.n7226 VSS.n2157 2.2505
R5596 VSS.n7228 VSS.n7227 2.2505
R5597 VSS.n7229 VSS.n2156 2.2505
R5598 VSS.n7231 VSS.n7230 2.2505
R5599 VSS.n7232 VSS.n2155 2.2505
R5600 VSS.n7234 VSS.n7233 2.2505
R5601 VSS.n7235 VSS.n2154 2.2505
R5602 VSS.n7237 VSS.n7236 2.2505
R5603 VSS.n7238 VSS.n2153 2.2505
R5604 VSS.n7240 VSS.n7239 2.2505
R5605 VSS.n7241 VSS.n2152 2.2505
R5606 VSS.n7243 VSS.n7242 2.2505
R5607 VSS.n7244 VSS.n2151 2.2505
R5608 VSS.n7246 VSS.n7245 2.2505
R5609 VSS.n7247 VSS.n2150 2.2505
R5610 VSS.n7249 VSS.n7248 2.2505
R5611 VSS.n7250 VSS.n2149 2.2505
R5612 VSS.n7252 VSS.n7251 2.2505
R5613 VSS.n7253 VSS.n2148 2.2505
R5614 VSS.n7255 VSS.n7254 2.2505
R5615 VSS.n7256 VSS.n2147 2.2505
R5616 VSS.n7258 VSS.n7257 2.2505
R5617 VSS.n7259 VSS.n2146 2.2505
R5618 VSS.n7261 VSS.n7260 2.2505
R5619 VSS.n7262 VSS.n2145 2.2505
R5620 VSS.n7264 VSS.n7263 2.2505
R5621 VSS.n7265 VSS.n2144 2.2505
R5622 VSS.n7267 VSS.n7266 2.2505
R5623 VSS.n7268 VSS.n2143 2.2505
R5624 VSS.n7270 VSS.n7269 2.2505
R5625 VSS.n7271 VSS.n2142 2.2505
R5626 VSS.n7273 VSS.n7272 2.2505
R5627 VSS.n7274 VSS.n2141 2.2505
R5628 VSS.n7276 VSS.n7275 2.2505
R5629 VSS.n7277 VSS.n2140 2.2505
R5630 VSS.n7279 VSS.n7278 2.2505
R5631 VSS.n7280 VSS.n2139 2.2505
R5632 VSS.n7282 VSS.n7281 2.2505
R5633 VSS.n7283 VSS.n2138 2.2505
R5634 VSS.n7285 VSS.n7284 2.2505
R5635 VSS.n7286 VSS.n2137 2.2505
R5636 VSS.n7288 VSS.n7287 2.2505
R5637 VSS.n7289 VSS.n2136 2.2505
R5638 VSS.n7291 VSS.n7290 2.2505
R5639 VSS.n7292 VSS.n2135 2.2505
R5640 VSS.n7294 VSS.n7293 2.2505
R5641 VSS.n7295 VSS.n2134 2.2505
R5642 VSS.n7297 VSS.n7296 2.2505
R5643 VSS.n7298 VSS.n2133 2.2505
R5644 VSS.n7300 VSS.n7299 2.2505
R5645 VSS.n7301 VSS.n2132 2.2505
R5646 VSS.n7303 VSS.n7302 2.2505
R5647 VSS.n7304 VSS.n2131 2.2505
R5648 VSS.n7306 VSS.n7305 2.2505
R5649 VSS.n7307 VSS.n2130 2.2505
R5650 VSS.n7309 VSS.n7308 2.2505
R5651 VSS.n7310 VSS.n2129 2.2505
R5652 VSS.n7312 VSS.n7311 2.2505
R5653 VSS.n7313 VSS.n2128 2.2505
R5654 VSS.n7315 VSS.n7314 2.2505
R5655 VSS.n7316 VSS.n2127 2.2505
R5656 VSS.n7318 VSS.n7317 2.2505
R5657 VSS.n7319 VSS.n2126 2.2505
R5658 VSS.n7321 VSS.n7320 2.2505
R5659 VSS.n7322 VSS.n2125 2.2505
R5660 VSS.n7324 VSS.n7323 2.2505
R5661 VSS.n7325 VSS.n2124 2.2505
R5662 VSS.n7327 VSS.n7326 2.2505
R5663 VSS.n7328 VSS.n2123 2.2505
R5664 VSS.n7330 VSS.n7329 2.2505
R5665 VSS.n7331 VSS.n2122 2.2505
R5666 VSS.n7333 VSS.n7332 2.2505
R5667 VSS.n7334 VSS.n2121 2.2505
R5668 VSS.n7336 VSS.n7335 2.2505
R5669 VSS.n7337 VSS.n2120 2.2505
R5670 VSS.n7339 VSS.n7338 2.2505
R5671 VSS.n7340 VSS.n2119 2.2505
R5672 VSS.n7342 VSS.n7341 2.2505
R5673 VSS.n7343 VSS.n2118 2.2505
R5674 VSS.n7345 VSS.n7344 2.2505
R5675 VSS.n7346 VSS.n2117 2.2505
R5676 VSS.n7348 VSS.n7347 2.2505
R5677 VSS.n7349 VSS.n2116 2.2505
R5678 VSS.n7351 VSS.n7350 2.2505
R5679 VSS.n7352 VSS.n2115 2.2505
R5680 VSS.n7354 VSS.n7353 2.2505
R5681 VSS.n7355 VSS.n2114 2.2505
R5682 VSS.n7357 VSS.n7356 2.2505
R5683 VSS.n7358 VSS.n2113 2.2505
R5684 VSS.n7360 VSS.n7359 2.2505
R5685 VSS.n7361 VSS.n2112 2.2505
R5686 VSS.n7363 VSS.n7362 2.2505
R5687 VSS.n7364 VSS.n2111 2.2505
R5688 VSS.n7366 VSS.n7365 2.2505
R5689 VSS.n7367 VSS.n2110 2.2505
R5690 VSS.n7369 VSS.n7368 2.2505
R5691 VSS.n7370 VSS.n2109 2.2505
R5692 VSS.n7372 VSS.n7371 2.2505
R5693 VSS.n7373 VSS.n2108 2.2505
R5694 VSS.n7375 VSS.n7374 2.2505
R5695 VSS.n7376 VSS.n2107 2.2505
R5696 VSS.n7378 VSS.n7377 2.2505
R5697 VSS.n7379 VSS.n2106 2.2505
R5698 VSS.n7381 VSS.n7380 2.2505
R5699 VSS.n7382 VSS.n2105 2.2505
R5700 VSS.n7384 VSS.n7383 2.2505
R5701 VSS.n7385 VSS.n2104 2.2505
R5702 VSS.n7387 VSS.n7386 2.2505
R5703 VSS.n7388 VSS.n2103 2.2505
R5704 VSS.n7390 VSS.n7389 2.2505
R5705 VSS.n7391 VSS.n2102 2.2505
R5706 VSS.n7393 VSS.n7392 2.2505
R5707 VSS.n7394 VSS.n2101 2.2505
R5708 VSS.n7396 VSS.n7395 2.2505
R5709 VSS.n7397 VSS.n2100 2.2505
R5710 VSS.n7399 VSS.n7398 2.2505
R5711 VSS.n7400 VSS.n2099 2.2505
R5712 VSS.n7402 VSS.n7401 2.2505
R5713 VSS.n7403 VSS.n2098 2.2505
R5714 VSS.n7405 VSS.n7404 2.2505
R5715 VSS.n7406 VSS.n2097 2.2505
R5716 VSS.n7408 VSS.n7407 2.2505
R5717 VSS.n7409 VSS.n2096 2.2505
R5718 VSS.n7411 VSS.n7410 2.2505
R5719 VSS.n7412 VSS.n2095 2.2505
R5720 VSS.n7414 VSS.n7413 2.2505
R5721 VSS.n7415 VSS.n2094 2.2505
R5722 VSS.n7417 VSS.n7416 2.2505
R5723 VSS.n7418 VSS.n2093 2.2505
R5724 VSS.n7420 VSS.n7419 2.2505
R5725 VSS.n7421 VSS.n2092 2.2505
R5726 VSS.n7423 VSS.n7422 2.2505
R5727 VSS.n7424 VSS.n2091 2.2505
R5728 VSS.n7426 VSS.n7425 2.2505
R5729 VSS.n7427 VSS.n2090 2.2505
R5730 VSS.n7429 VSS.n7428 2.2505
R5731 VSS.n7430 VSS.n2089 2.2505
R5732 VSS.n7432 VSS.n7431 2.2505
R5733 VSS.n7433 VSS.n2088 2.2505
R5734 VSS.n7435 VSS.n7434 2.2505
R5735 VSS.n7436 VSS.n2087 2.2505
R5736 VSS.n7438 VSS.n7437 2.2505
R5737 VSS.n7439 VSS.n2086 2.2505
R5738 VSS.n7441 VSS.n7440 2.2505
R5739 VSS.n7442 VSS.n2085 2.2505
R5740 VSS.n7444 VSS.n7443 2.2505
R5741 VSS.n7445 VSS.n2084 2.2505
R5742 VSS.n7447 VSS.n7446 2.2505
R5743 VSS.n7448 VSS.n2083 2.2505
R5744 VSS.n7450 VSS.n7449 2.2505
R5745 VSS.n7451 VSS.n2082 2.2505
R5746 VSS.n7453 VSS.n7452 2.2505
R5747 VSS.n7454 VSS.n2081 2.2505
R5748 VSS.n7456 VSS.n7455 2.2505
R5749 VSS.n7457 VSS.n2080 2.2505
R5750 VSS.n7459 VSS.n7458 2.2505
R5751 VSS.n7460 VSS.n2079 2.2505
R5752 VSS.n7462 VSS.n7461 2.2505
R5753 VSS.n7463 VSS.n2078 2.2505
R5754 VSS.n7465 VSS.n7464 2.2505
R5755 VSS.n7466 VSS.n2077 2.2505
R5756 VSS.n7468 VSS.n7467 2.2505
R5757 VSS.n7469 VSS.n2076 2.2505
R5758 VSS.n7471 VSS.n7470 2.2505
R5759 VSS.n7472 VSS.n2075 2.2505
R5760 VSS.n7474 VSS.n7473 2.2505
R5761 VSS.n7475 VSS.n2074 2.2505
R5762 VSS.n7477 VSS.n7476 2.2505
R5763 VSS.n7478 VSS.n2073 2.2505
R5764 VSS.n7480 VSS.n7479 2.2505
R5765 VSS.n7481 VSS.n2072 2.2505
R5766 VSS.n7483 VSS.n7482 2.2505
R5767 VSS.n7484 VSS.n2071 2.2505
R5768 VSS.n7486 VSS.n7485 2.2505
R5769 VSS.n7487 VSS.n2070 2.2505
R5770 VSS.n7489 VSS.n7488 2.2505
R5771 VSS.n7490 VSS.n2069 2.2505
R5772 VSS.n7492 VSS.n7491 2.2505
R5773 VSS.n7493 VSS.n2068 2.2505
R5774 VSS.n7495 VSS.n7494 2.2505
R5775 VSS.n7496 VSS.n2067 2.2505
R5776 VSS.n7498 VSS.n7497 2.2505
R5777 VSS.n7499 VSS.n2066 2.2505
R5778 VSS.n7501 VSS.n7500 2.2505
R5779 VSS.n7502 VSS.n2065 2.2505
R5780 VSS.n7504 VSS.n7503 2.2505
R5781 VSS.n7505 VSS.n2064 2.2505
R5782 VSS.n7507 VSS.n7506 2.2505
R5783 VSS.n7508 VSS.n2063 2.2505
R5784 VSS.n7510 VSS.n7509 2.2505
R5785 VSS.n7511 VSS.n2062 2.2505
R5786 VSS.n7513 VSS.n7512 2.2505
R5787 VSS.n7514 VSS.n2061 2.2505
R5788 VSS.n7516 VSS.n7515 2.2505
R5789 VSS.n7517 VSS.n2060 2.2505
R5790 VSS.n7519 VSS.n7518 2.2505
R5791 VSS.n7520 VSS.n2059 2.2505
R5792 VSS.n7522 VSS.n7521 2.2505
R5793 VSS.n7523 VSS.n2058 2.2505
R5794 VSS.n7525 VSS.n7524 2.2505
R5795 VSS.n7526 VSS.n2057 2.2505
R5796 VSS.n7528 VSS.n7527 2.2505
R5797 VSS.n7529 VSS.n2056 2.2505
R5798 VSS.n7531 VSS.n7530 2.2505
R5799 VSS.n7532 VSS.n2055 2.2505
R5800 VSS.n7534 VSS.n7533 2.2505
R5801 VSS.n7535 VSS.n2054 2.2505
R5802 VSS.n7537 VSS.n7536 2.2505
R5803 VSS.n7538 VSS.n2053 2.2505
R5804 VSS.n7540 VSS.n7539 2.2505
R5805 VSS.n7541 VSS.n2052 2.2505
R5806 VSS.n7543 VSS.n7542 2.2505
R5807 VSS.n7544 VSS.n2051 2.2505
R5808 VSS.n7546 VSS.n7545 2.2505
R5809 VSS.n7547 VSS.n2050 2.2505
R5810 VSS.n7549 VSS.n7548 2.2505
R5811 VSS.n7550 VSS.n2049 2.2505
R5812 VSS.n7552 VSS.n7551 2.2505
R5813 VSS.n7553 VSS.n2048 2.2505
R5814 VSS.n7555 VSS.n7554 2.2505
R5815 VSS.n7556 VSS.n2047 2.2505
R5816 VSS.n7558 VSS.n7557 2.2505
R5817 VSS.n7559 VSS.n2046 2.2505
R5818 VSS.n7561 VSS.n7560 2.2505
R5819 VSS.n7562 VSS.n2045 2.2505
R5820 VSS.n7564 VSS.n7563 2.2505
R5821 VSS.n7565 VSS.n2044 2.2505
R5822 VSS.n7567 VSS.n7566 2.2505
R5823 VSS.n7568 VSS.n2043 2.2505
R5824 VSS.n7570 VSS.n7569 2.2505
R5825 VSS.n7571 VSS.n2042 2.2505
R5826 VSS.n7573 VSS.n7572 2.2505
R5827 VSS.n7574 VSS.n2041 2.2505
R5828 VSS.n7576 VSS.n7575 2.2505
R5829 VSS.n7577 VSS.n2040 2.2505
R5830 VSS.n7579 VSS.n7578 2.2505
R5831 VSS.n7580 VSS.n2039 2.2505
R5832 VSS.n7582 VSS.n7581 2.2505
R5833 VSS.n7583 VSS.n2038 2.2505
R5834 VSS.n7585 VSS.n7584 2.2505
R5835 VSS.n7586 VSS.n2037 2.2505
R5836 VSS.n7588 VSS.n7587 2.2505
R5837 VSS.n7589 VSS.n2036 2.2505
R5838 VSS.n7591 VSS.n7590 2.2505
R5839 VSS.n7592 VSS.n2035 2.2505
R5840 VSS.n7594 VSS.n7593 2.2505
R5841 VSS.n7595 VSS.n2034 2.2505
R5842 VSS.n7597 VSS.n7596 2.2505
R5843 VSS.n7598 VSS.n2033 2.2505
R5844 VSS.n7600 VSS.n7599 2.2505
R5845 VSS.n7601 VSS.n2032 2.2505
R5846 VSS.n7603 VSS.n7602 2.2505
R5847 VSS.n7604 VSS.n2031 2.2505
R5848 VSS.n7606 VSS.n7605 2.2505
R5849 VSS.n7607 VSS.n2030 2.2505
R5850 VSS.n7609 VSS.n7608 2.2505
R5851 VSS.n7610 VSS.n2029 2.2505
R5852 VSS.n7612 VSS.n7611 2.2505
R5853 VSS.n7613 VSS.n2028 2.2505
R5854 VSS.n7615 VSS.n7614 2.2505
R5855 VSS.n7616 VSS.n2027 2.2505
R5856 VSS.n7618 VSS.n7617 2.2505
R5857 VSS.n7619 VSS.n2026 2.2505
R5858 VSS.n7621 VSS.n7620 2.2505
R5859 VSS.n7622 VSS.n2025 2.2505
R5860 VSS.n7624 VSS.n7623 2.2505
R5861 VSS.n7625 VSS.n2024 2.2505
R5862 VSS.n7627 VSS.n7626 2.2505
R5863 VSS.n7628 VSS.n2023 2.2505
R5864 VSS.n7630 VSS.n7629 2.2505
R5865 VSS.n7631 VSS.n2022 2.2505
R5866 VSS.n7633 VSS.n7632 2.2505
R5867 VSS.n7634 VSS.n2021 2.2505
R5868 VSS.n7636 VSS.n7635 2.2505
R5869 VSS.n7637 VSS.n2020 2.2505
R5870 VSS.n7639 VSS.n7638 2.2505
R5871 VSS.n7640 VSS.n2019 2.2505
R5872 VSS.n7642 VSS.n7641 2.2505
R5873 VSS.n7643 VSS.n2018 2.2505
R5874 VSS.n7645 VSS.n7644 2.2505
R5875 VSS.n7646 VSS.n2017 2.2505
R5876 VSS.n7648 VSS.n7647 2.2505
R5877 VSS.n7649 VSS.n2016 2.2505
R5878 VSS.n7651 VSS.n7650 2.2505
R5879 VSS.n7652 VSS.n2015 2.2505
R5880 VSS.n7654 VSS.n7653 2.2505
R5881 VSS.n7655 VSS.n2014 2.2505
R5882 VSS.n7657 VSS.n7656 2.2505
R5883 VSS.n7658 VSS.n2013 2.2505
R5884 VSS.n7660 VSS.n7659 2.2505
R5885 VSS.n7661 VSS.n2012 2.2505
R5886 VSS.n7663 VSS.n7662 2.2505
R5887 VSS.n7664 VSS.n2011 2.2505
R5888 VSS.n7666 VSS.n7665 2.2505
R5889 VSS.n7667 VSS.n2010 2.2505
R5890 VSS.n7669 VSS.n7668 2.2505
R5891 VSS.n7670 VSS.n2009 2.2505
R5892 VSS.n7672 VSS.n7671 2.2505
R5893 VSS.n7673 VSS.n2008 2.2505
R5894 VSS.n7675 VSS.n7674 2.2505
R5895 VSS.n7676 VSS.n2007 2.2505
R5896 VSS.n7678 VSS.n7677 2.2505
R5897 VSS.n7679 VSS.n2006 2.2505
R5898 VSS.n7681 VSS.n7680 2.2505
R5899 VSS.n7682 VSS.n2005 2.2505
R5900 VSS.n7684 VSS.n7683 2.2505
R5901 VSS.n7685 VSS.n2004 2.2505
R5902 VSS.n7687 VSS.n7686 2.2505
R5903 VSS.n7688 VSS.n2003 2.2505
R5904 VSS.n7690 VSS.n7689 2.2505
R5905 VSS.n7691 VSS.n2002 2.2505
R5906 VSS.n7693 VSS.n7692 2.2505
R5907 VSS.n7694 VSS.n2001 2.2505
R5908 VSS.n7696 VSS.n7695 2.2505
R5909 VSS.n7697 VSS.n2000 2.2505
R5910 VSS.n7699 VSS.n7698 2.2505
R5911 VSS.n7700 VSS.n1999 2.2505
R5912 VSS.n7702 VSS.n7701 2.2505
R5913 VSS.n7703 VSS.n1998 2.2505
R5914 VSS.n7705 VSS.n7704 2.2505
R5915 VSS.n7706 VSS.n1997 2.2505
R5916 VSS.n7708 VSS.n7707 2.2505
R5917 VSS.n7709 VSS.n1996 2.2505
R5918 VSS.n7711 VSS.n7710 2.2505
R5919 VSS.n7712 VSS.n1995 2.2505
R5920 VSS.n7714 VSS.n7713 2.2505
R5921 VSS.n7715 VSS.n1994 2.2505
R5922 VSS.n7717 VSS.n7716 2.2505
R5923 VSS.n7718 VSS.n1993 2.2505
R5924 VSS.n7720 VSS.n7719 2.2505
R5925 VSS.n7721 VSS.n1992 2.2505
R5926 VSS.n7723 VSS.n7722 2.2505
R5927 VSS.n7724 VSS.n1991 2.2505
R5928 VSS.n7726 VSS.n7725 2.2505
R5929 VSS.n7727 VSS.n1990 2.2505
R5930 VSS.n7729 VSS.n7728 2.2505
R5931 VSS.n7730 VSS.n1989 2.2505
R5932 VSS.n7732 VSS.n7731 2.2505
R5933 VSS.n7733 VSS.n1988 2.2505
R5934 VSS.n7735 VSS.n7734 2.2505
R5935 VSS.n7736 VSS.n1987 2.2505
R5936 VSS.n7738 VSS.n7737 2.2505
R5937 VSS.n7739 VSS.n1986 2.2505
R5938 VSS.n7741 VSS.n7740 2.2505
R5939 VSS.n7742 VSS.n1985 2.2505
R5940 VSS.n7744 VSS.n7743 2.2505
R5941 VSS.n7745 VSS.n1984 2.2505
R5942 VSS.n7747 VSS.n7746 2.2505
R5943 VSS.n7748 VSS.n1983 2.2505
R5944 VSS.n7750 VSS.n7749 2.2505
R5945 VSS.n7751 VSS.n1982 2.2505
R5946 VSS.n7753 VSS.n7752 2.2505
R5947 VSS.n7754 VSS.n1981 2.2505
R5948 VSS.n7756 VSS.n7755 2.2505
R5949 VSS.n7757 VSS.n1980 2.2505
R5950 VSS.n7759 VSS.n7758 2.2505
R5951 VSS.n7760 VSS.n1979 2.2505
R5952 VSS.n7762 VSS.n7761 2.2505
R5953 VSS.n7763 VSS.n1978 2.2505
R5954 VSS.n7765 VSS.n7764 2.2505
R5955 VSS.n7766 VSS.n1977 2.2505
R5956 VSS.n7768 VSS.n7767 2.2505
R5957 VSS.n7769 VSS.n1976 2.2505
R5958 VSS.n7771 VSS.n7770 2.2505
R5959 VSS.n7772 VSS.n1975 2.2505
R5960 VSS.n7774 VSS.n7773 2.2505
R5961 VSS.n7775 VSS.n1974 2.2505
R5962 VSS.n7777 VSS.n7776 2.2505
R5963 VSS.n7778 VSS.n1973 2.2505
R5964 VSS.n7780 VSS.n7779 2.2505
R5965 VSS.n7781 VSS.n1972 2.2505
R5966 VSS.n7783 VSS.n7782 2.2505
R5967 VSS.n7784 VSS.n1971 2.2505
R5968 VSS.n7786 VSS.n7785 2.2505
R5969 VSS.n7787 VSS.n1970 2.2505
R5970 VSS.n7789 VSS.n7788 2.2505
R5971 VSS.n7790 VSS.n1969 2.2505
R5972 VSS.n7792 VSS.n7791 2.2505
R5973 VSS.n7793 VSS.n1968 2.2505
R5974 VSS.n7795 VSS.n7794 2.2505
R5975 VSS.n7796 VSS.n1967 2.2505
R5976 VSS.n7798 VSS.n7797 2.2505
R5977 VSS.n7799 VSS.n1966 2.2505
R5978 VSS.n7801 VSS.n7800 2.2505
R5979 VSS.n7802 VSS.n1965 2.2505
R5980 VSS.n7804 VSS.n7803 2.2505
R5981 VSS.n7805 VSS.n1964 2.2505
R5982 VSS.n7807 VSS.n7806 2.2505
R5983 VSS.n7808 VSS.n1963 2.2505
R5984 VSS.n7810 VSS.n7809 2.2505
R5985 VSS.n7811 VSS.n1962 2.2505
R5986 VSS.n7813 VSS.n7812 2.2505
R5987 VSS.n7814 VSS.n1961 2.2505
R5988 VSS.n7816 VSS.n7815 2.2505
R5989 VSS.n7817 VSS.n1960 2.2505
R5990 VSS.n7819 VSS.n7818 2.2505
R5991 VSS.n7820 VSS.n1959 2.2505
R5992 VSS.n7822 VSS.n7821 2.2505
R5993 VSS.n7823 VSS.n1958 2.2505
R5994 VSS.n7825 VSS.n7824 2.2505
R5995 VSS.n7826 VSS.n1957 2.2505
R5996 VSS.n7828 VSS.n7827 2.2505
R5997 VSS.n7829 VSS.n1956 2.2505
R5998 VSS.n7831 VSS.n7830 2.2505
R5999 VSS.n7832 VSS.n1955 2.2505
R6000 VSS.n7834 VSS.n7833 2.2505
R6001 VSS.n7835 VSS.n1954 2.2505
R6002 VSS.n7837 VSS.n7836 2.2505
R6003 VSS.n7838 VSS.n1953 2.2505
R6004 VSS.n7840 VSS.n7839 2.2505
R6005 VSS.n7841 VSS.n1952 2.2505
R6006 VSS.n7843 VSS.n7842 2.2505
R6007 VSS.n7844 VSS.n1951 2.2505
R6008 VSS.n7846 VSS.n7845 2.2505
R6009 VSS.n7847 VSS.n1950 2.2505
R6010 VSS.n7849 VSS.n7848 2.2505
R6011 VSS.n7850 VSS.n1949 2.2505
R6012 VSS.n7852 VSS.n7851 2.2505
R6013 VSS.n7853 VSS.n1948 2.2505
R6014 VSS.n7855 VSS.n7854 2.2505
R6015 VSS.n7856 VSS.n1947 2.2505
R6016 VSS.n7858 VSS.n7857 2.2505
R6017 VSS.n7859 VSS.n1946 2.2505
R6018 VSS.n7861 VSS.n7860 2.2505
R6019 VSS.n7862 VSS.n1945 2.2505
R6020 VSS.n7864 VSS.n7863 2.2505
R6021 VSS.n7865 VSS.n1944 2.2505
R6022 VSS.n7867 VSS.n7866 2.2505
R6023 VSS.n7868 VSS.n1943 2.2505
R6024 VSS.n7870 VSS.n7869 2.2505
R6025 VSS.n7871 VSS.n1942 2.2505
R6026 VSS.n7873 VSS.n7872 2.2505
R6027 VSS.n7874 VSS.n1941 2.2505
R6028 VSS.n7876 VSS.n7875 2.2505
R6029 VSS.n7877 VSS.n1940 2.2505
R6030 VSS.n7879 VSS.n7878 2.2505
R6031 VSS.n7880 VSS.n1939 2.2505
R6032 VSS.n7882 VSS.n7881 2.2505
R6033 VSS.n7883 VSS.n1938 2.2505
R6034 VSS.n7885 VSS.n7884 2.2505
R6035 VSS.n7886 VSS.n1937 2.2505
R6036 VSS.n7888 VSS.n7887 2.2505
R6037 VSS.n7889 VSS.n1936 2.2505
R6038 VSS.n7891 VSS.n7890 2.2505
R6039 VSS.n7892 VSS.n1935 2.2505
R6040 VSS.n7894 VSS.n7893 2.2505
R6041 VSS.n7895 VSS.n1934 2.2505
R6042 VSS.n7897 VSS.n7896 2.2505
R6043 VSS.n7898 VSS.n1933 2.2505
R6044 VSS.n7900 VSS.n7899 2.2505
R6045 VSS.n7901 VSS.n1932 2.2505
R6046 VSS.n7903 VSS.n7902 2.2505
R6047 VSS.n7904 VSS.n1931 2.2505
R6048 VSS.n7906 VSS.n7905 2.2505
R6049 VSS.n7907 VSS.n1930 2.2505
R6050 VSS.n7909 VSS.n7908 2.2505
R6051 VSS.n7910 VSS.n1929 2.2505
R6052 VSS.n7912 VSS.n7911 2.2505
R6053 VSS.n7913 VSS.n1928 2.2505
R6054 VSS.n7915 VSS.n7914 2.2505
R6055 VSS.n7916 VSS.n1927 2.2505
R6056 VSS.n7918 VSS.n7917 2.2505
R6057 VSS.n7919 VSS.n1926 2.2505
R6058 VSS.n7921 VSS.n7920 2.2505
R6059 VSS.n7922 VSS.n1925 2.2505
R6060 VSS.n7924 VSS.n7923 2.2505
R6061 VSS.n7925 VSS.n1924 2.2505
R6062 VSS.n7927 VSS.n7926 2.2505
R6063 VSS.n7928 VSS.n1923 2.2505
R6064 VSS.n7930 VSS.n7929 2.2505
R6065 VSS.n7931 VSS.n1922 2.2505
R6066 VSS.n7933 VSS.n7932 2.2505
R6067 VSS.n7934 VSS.n1921 2.2505
R6068 VSS.n7936 VSS.n7935 2.2505
R6069 VSS.n7937 VSS.n1920 2.2505
R6070 VSS.n7939 VSS.n7938 2.2505
R6071 VSS.n7940 VSS.n1919 2.2505
R6072 VSS.n7942 VSS.n7941 2.2505
R6073 VSS.n7943 VSS.n1918 2.2505
R6074 VSS.n7945 VSS.n7944 2.2505
R6075 VSS.n7946 VSS.n1917 2.2505
R6076 VSS.n7948 VSS.n7947 2.2505
R6077 VSS.n7949 VSS.n1916 2.2505
R6078 VSS.n7951 VSS.n7950 2.2505
R6079 VSS.n7952 VSS.n1915 2.2505
R6080 VSS.n7954 VSS.n7953 2.2505
R6081 VSS.n7955 VSS.n1914 2.2505
R6082 VSS.n7957 VSS.n7956 2.2505
R6083 VSS.n7958 VSS.n1913 2.2505
R6084 VSS.n7960 VSS.n7959 2.2505
R6085 VSS.n7961 VSS.n1912 2.2505
R6086 VSS.n7963 VSS.n7962 2.2505
R6087 VSS.n7964 VSS.n1911 2.2505
R6088 VSS.n7966 VSS.n7965 2.2505
R6089 VSS.n7967 VSS.n1910 2.2505
R6090 VSS.n7969 VSS.n7968 2.2505
R6091 VSS.n7970 VSS.n1909 2.2505
R6092 VSS.n7972 VSS.n7971 2.2505
R6093 VSS.n7973 VSS.n1908 2.2505
R6094 VSS.n7975 VSS.n7974 2.2505
R6095 VSS.n7976 VSS.n1907 2.2505
R6096 VSS.n7978 VSS.n7977 2.2505
R6097 VSS.n7979 VSS.n1906 2.2505
R6098 VSS.n7981 VSS.n7980 2.2505
R6099 VSS.n7982 VSS.n1905 2.2505
R6100 VSS.n7984 VSS.n7983 2.2505
R6101 VSS.n7985 VSS.n1904 2.2505
R6102 VSS.n7987 VSS.n7986 2.2505
R6103 VSS.n7988 VSS.n1903 2.2505
R6104 VSS.n7990 VSS.n7989 2.2505
R6105 VSS.n7991 VSS.n1902 2.2505
R6106 VSS.n7993 VSS.n7992 2.2505
R6107 VSS.n7994 VSS.n1901 2.2505
R6108 VSS.n7996 VSS.n7995 2.2505
R6109 VSS.n7997 VSS.n1900 2.2505
R6110 VSS.n7999 VSS.n7998 2.2505
R6111 VSS.n8000 VSS.n1899 2.2505
R6112 VSS.n8002 VSS.n8001 2.2505
R6113 VSS.n8003 VSS.n1898 2.2505
R6114 VSS.n8005 VSS.n8004 2.2505
R6115 VSS.n8006 VSS.n1897 2.2505
R6116 VSS.n8008 VSS.n8007 2.2505
R6117 VSS.n8009 VSS.n1896 2.2505
R6118 VSS.n8011 VSS.n8010 2.2505
R6119 VSS.n8012 VSS.n1895 2.2505
R6120 VSS.n8014 VSS.n8013 2.2505
R6121 VSS.n8015 VSS.n1894 2.2505
R6122 VSS.n8017 VSS.n8016 2.2505
R6123 VSS.n8018 VSS.n1893 2.2505
R6124 VSS.n8020 VSS.n8019 2.2505
R6125 VSS.n8021 VSS.n1892 2.2505
R6126 VSS.n8023 VSS.n8022 2.2505
R6127 VSS.n8024 VSS.n1891 2.2505
R6128 VSS.n8026 VSS.n8025 2.2505
R6129 VSS.n8027 VSS.n1890 2.2505
R6130 VSS.n8029 VSS.n8028 2.2505
R6131 VSS.n8030 VSS.n1889 2.2505
R6132 VSS.n8032 VSS.n8031 2.2505
R6133 VSS.n8033 VSS.n1888 2.2505
R6134 VSS.n8035 VSS.n8034 2.2505
R6135 VSS.n8036 VSS.n1887 2.2505
R6136 VSS.n8038 VSS.n8037 2.2505
R6137 VSS.n8039 VSS.n1886 2.2505
R6138 VSS.n8041 VSS.n8040 2.2505
R6139 VSS.n8042 VSS.n1885 2.2505
R6140 VSS.n8044 VSS.n8043 2.2505
R6141 VSS.n8045 VSS.n1884 2.2505
R6142 VSS.n8047 VSS.n8046 2.2505
R6143 VSS.n8048 VSS.n1883 2.2505
R6144 VSS.n8050 VSS.n8049 2.2505
R6145 VSS.n8051 VSS.n1882 2.2505
R6146 VSS.n8053 VSS.n8052 2.2505
R6147 VSS.n8054 VSS.n1881 2.2505
R6148 VSS.n8056 VSS.n8055 2.2505
R6149 VSS.n8057 VSS.n1880 2.2505
R6150 VSS.n8059 VSS.n8058 2.2505
R6151 VSS.n8060 VSS.n1879 2.2505
R6152 VSS.n8062 VSS.n8061 2.2505
R6153 VSS.n8063 VSS.n1878 2.2505
R6154 VSS.n8065 VSS.n8064 2.2505
R6155 VSS.n8066 VSS.n1877 2.2505
R6156 VSS.n8068 VSS.n8067 2.2505
R6157 VSS.n8069 VSS.n1876 2.2505
R6158 VSS.n8071 VSS.n8070 2.2505
R6159 VSS.n8072 VSS.n1875 2.2505
R6160 VSS.n8074 VSS.n8073 2.2505
R6161 VSS.n8075 VSS.n1874 2.2505
R6162 VSS.n8077 VSS.n8076 2.2505
R6163 VSS.n8078 VSS.n1873 2.2505
R6164 VSS.n8080 VSS.n8079 2.2505
R6165 VSS.n8081 VSS.n1872 2.2505
R6166 VSS.n8083 VSS.n8082 2.2505
R6167 VSS.n8084 VSS.n1871 2.2505
R6168 VSS.n8086 VSS.n8085 2.2505
R6169 VSS.n8087 VSS.n1870 2.2505
R6170 VSS.n8089 VSS.n8088 2.2505
R6171 VSS.n8090 VSS.n1869 2.2505
R6172 VSS.n8092 VSS.n8091 2.2505
R6173 VSS.n8093 VSS.n1868 2.2505
R6174 VSS.n8095 VSS.n8094 2.2505
R6175 VSS.n8096 VSS.n1867 2.2505
R6176 VSS.n8098 VSS.n8097 2.2505
R6177 VSS.n8099 VSS.n1866 2.2505
R6178 VSS.n8101 VSS.n8100 2.2505
R6179 VSS.n8102 VSS.n1865 2.2505
R6180 VSS.n8104 VSS.n8103 2.2505
R6181 VSS.n8105 VSS.n1864 2.2505
R6182 VSS.n8107 VSS.n8106 2.2505
R6183 VSS.n8108 VSS.n1863 2.2505
R6184 VSS.n8110 VSS.n8109 2.2505
R6185 VSS.n8111 VSS.n1862 2.2505
R6186 VSS.n8113 VSS.n8112 2.2505
R6187 VSS.n8114 VSS.n1861 2.2505
R6188 VSS.n8116 VSS.n8115 2.2505
R6189 VSS.n8117 VSS.n1860 2.2505
R6190 VSS.n8119 VSS.n8118 2.2505
R6191 VSS.n8120 VSS.n1859 2.2505
R6192 VSS.n8122 VSS.n8121 2.2505
R6193 VSS.n8123 VSS.n1858 2.2505
R6194 VSS.n8125 VSS.n8124 2.2505
R6195 VSS.n8126 VSS.n1857 2.2505
R6196 VSS.n8128 VSS.n8127 2.2505
R6197 VSS.n8129 VSS.n1856 2.2505
R6198 VSS.n8131 VSS.n8130 2.2505
R6199 VSS.n8132 VSS.n1855 2.2505
R6200 VSS.n8134 VSS.n8133 2.2505
R6201 VSS.n8135 VSS.n1854 2.2505
R6202 VSS.n8137 VSS.n8136 2.2505
R6203 VSS.n8138 VSS.n1853 2.2505
R6204 VSS.n8140 VSS.n8139 2.2505
R6205 VSS.n8141 VSS.n1852 2.2505
R6206 VSS.n8143 VSS.n8142 2.2505
R6207 VSS.n8144 VSS.n1851 2.2505
R6208 VSS.n8146 VSS.n8145 2.2505
R6209 VSS.n8147 VSS.n1850 2.2505
R6210 VSS.n8149 VSS.n8148 2.2505
R6211 VSS.n8150 VSS.n1849 2.2505
R6212 VSS.n8152 VSS.n8151 2.2505
R6213 VSS.n8153 VSS.n1848 2.2505
R6214 VSS.n8155 VSS.n8154 2.2505
R6215 VSS.n8156 VSS.n1847 2.2505
R6216 VSS.n8158 VSS.n8157 2.2505
R6217 VSS.n8159 VSS.n1846 2.2505
R6218 VSS.n8161 VSS.n8160 2.2505
R6219 VSS.n8162 VSS.n1845 2.2505
R6220 VSS.n8164 VSS.n8163 2.2505
R6221 VSS.n8165 VSS.n1844 2.2505
R6222 VSS.n8167 VSS.n8166 2.2505
R6223 VSS.n8168 VSS.n1843 2.2505
R6224 VSS.n8170 VSS.n8169 2.2505
R6225 VSS.n8171 VSS.n1842 2.2505
R6226 VSS.n8173 VSS.n8172 2.2505
R6227 VSS.n8174 VSS.n1841 2.2505
R6228 VSS.n8176 VSS.n8175 2.2505
R6229 VSS.n8177 VSS.n1840 2.2505
R6230 VSS.n8179 VSS.n8178 2.2505
R6231 VSS.n8180 VSS.n1839 2.2505
R6232 VSS.n8182 VSS.n8181 2.2505
R6233 VSS.n8183 VSS.n1838 2.2505
R6234 VSS.n8185 VSS.n8184 2.2505
R6235 VSS.n8186 VSS.n1837 2.2505
R6236 VSS.n8188 VSS.n8187 2.2505
R6237 VSS.n8189 VSS.n1836 2.2505
R6238 VSS.n8191 VSS.n8190 2.2505
R6239 VSS.n8192 VSS.n1835 2.2505
R6240 VSS.n8194 VSS.n8193 2.2505
R6241 VSS.n8195 VSS.n1834 2.2505
R6242 VSS.n8197 VSS.n8196 2.2505
R6243 VSS.n8198 VSS.n1833 2.2505
R6244 VSS.n8200 VSS.n8199 2.2505
R6245 VSS.n8201 VSS.n1832 2.2505
R6246 VSS.n8203 VSS.n8202 2.2505
R6247 VSS.n8204 VSS.n1831 2.2505
R6248 VSS.n8206 VSS.n8205 2.2505
R6249 VSS.n8207 VSS.n1830 2.2505
R6250 VSS.n8209 VSS.n8208 2.2505
R6251 VSS.n8210 VSS.n1829 2.2505
R6252 VSS.n8212 VSS.n8211 2.2505
R6253 VSS.n8213 VSS.n1828 2.2505
R6254 VSS.n8215 VSS.n8214 2.2505
R6255 VSS.n8216 VSS.n1827 2.2505
R6256 VSS.n8218 VSS.n8217 2.2505
R6257 VSS.n8219 VSS.n1826 2.2505
R6258 VSS.n8221 VSS.n8220 2.2505
R6259 VSS.n8222 VSS.n1825 2.2505
R6260 VSS.n8224 VSS.n8223 2.2505
R6261 VSS.n8225 VSS.n1824 2.2505
R6262 VSS.n8227 VSS.n8226 2.2505
R6263 VSS.n8228 VSS.n1823 2.2505
R6264 VSS.n8230 VSS.n8229 2.2505
R6265 VSS.n8231 VSS.n1822 2.2505
R6266 VSS.n4141 VSS.n4140 2.2505
R6267 VSS.n4139 VSS.n3185 2.2505
R6268 VSS.n4138 VSS.n4137 2.2505
R6269 VSS.n4136 VSS.n3186 2.2505
R6270 VSS.n4135 VSS.n4134 2.2505
R6271 VSS.n4133 VSS.n3187 2.2505
R6272 VSS.n4132 VSS.n4131 2.2505
R6273 VSS.n4130 VSS.n3188 2.2505
R6274 VSS.n4129 VSS.n4128 2.2505
R6275 VSS.n4127 VSS.n3189 2.2505
R6276 VSS.n4126 VSS.n4125 2.2505
R6277 VSS.n4124 VSS.n3190 2.2505
R6278 VSS.n4123 VSS.n4122 2.2505
R6279 VSS.n4121 VSS.n3191 2.2505
R6280 VSS.n4120 VSS.n4119 2.2505
R6281 VSS.n4118 VSS.n3192 2.2505
R6282 VSS.n4117 VSS.n4116 2.2505
R6283 VSS.n4115 VSS.n3193 2.2505
R6284 VSS.n4114 VSS.n4113 2.2505
R6285 VSS.n4112 VSS.n3194 2.2505
R6286 VSS.n4111 VSS.n4110 2.2505
R6287 VSS.n4109 VSS.n3195 2.2505
R6288 VSS.n4108 VSS.n4107 2.2505
R6289 VSS.n4106 VSS.n3196 2.2505
R6290 VSS.n4105 VSS.n4104 2.2505
R6291 VSS.n4103 VSS.n3197 2.2505
R6292 VSS.n4102 VSS.n4101 2.2505
R6293 VSS.n4100 VSS.n3198 2.2505
R6294 VSS.n4099 VSS.n4098 2.2505
R6295 VSS.n4097 VSS.n3199 2.2505
R6296 VSS.n4096 VSS.n4095 2.2505
R6297 VSS.n4094 VSS.n3200 2.2505
R6298 VSS.n4093 VSS.n4092 2.2505
R6299 VSS.n4091 VSS.n3201 2.2505
R6300 VSS.n4090 VSS.n4089 2.2505
R6301 VSS.n4088 VSS.n3202 2.2505
R6302 VSS.n4087 VSS.n4086 2.2505
R6303 VSS.n4085 VSS.n3203 2.2505
R6304 VSS.n4084 VSS.n4083 2.2505
R6305 VSS.n4082 VSS.n3204 2.2505
R6306 VSS.n4081 VSS.n4080 2.2505
R6307 VSS.n4079 VSS.n3205 2.2505
R6308 VSS.n4078 VSS.n4077 2.2505
R6309 VSS.n4076 VSS.n3206 2.2505
R6310 VSS.n4075 VSS.n4074 2.2505
R6311 VSS.n4073 VSS.n3207 2.2505
R6312 VSS.n4072 VSS.n4071 2.2505
R6313 VSS.n4070 VSS.n3208 2.2505
R6314 VSS.n4069 VSS.n4068 2.2505
R6315 VSS.n4067 VSS.n3209 2.2505
R6316 VSS.n4066 VSS.n4065 2.2505
R6317 VSS.n4064 VSS.n3210 2.2505
R6318 VSS.n4063 VSS.n4062 2.2505
R6319 VSS.n4061 VSS.n3211 2.2505
R6320 VSS.n4060 VSS.n4059 2.2505
R6321 VSS.n4058 VSS.n3212 2.2505
R6322 VSS.n4057 VSS.n4056 2.2505
R6323 VSS.n4055 VSS.n3213 2.2505
R6324 VSS.n4054 VSS.n4053 2.2505
R6325 VSS.n4052 VSS.n3214 2.2505
R6326 VSS.n4051 VSS.n4050 2.2505
R6327 VSS.n4049 VSS.n3215 2.2505
R6328 VSS.n4048 VSS.n4047 2.2505
R6329 VSS.n4046 VSS.n3216 2.2505
R6330 VSS.n4045 VSS.n4044 2.2505
R6331 VSS.n4043 VSS.n3217 2.2505
R6332 VSS.n4042 VSS.n4041 2.2505
R6333 VSS.n4040 VSS.n3218 2.2505
R6334 VSS.n4039 VSS.n4038 2.2505
R6335 VSS.n4037 VSS.n3219 2.2505
R6336 VSS.n4036 VSS.n4035 2.2505
R6337 VSS.n4034 VSS.n3220 2.2505
R6338 VSS.n4033 VSS.n4032 2.2505
R6339 VSS.n4031 VSS.n3221 2.2505
R6340 VSS.n4030 VSS.n4029 2.2505
R6341 VSS.n4028 VSS.n3222 2.2505
R6342 VSS.n4027 VSS.n4026 2.2505
R6343 VSS.n4025 VSS.n3223 2.2505
R6344 VSS.n4024 VSS.n4023 2.2505
R6345 VSS.n4022 VSS.n3224 2.2505
R6346 VSS.n4021 VSS.n4020 2.2505
R6347 VSS.n4019 VSS.n3225 2.2505
R6348 VSS.n4018 VSS.n4017 2.2505
R6349 VSS.n4016 VSS.n3226 2.2505
R6350 VSS.n4015 VSS.n4014 2.2505
R6351 VSS.n4013 VSS.n3227 2.2505
R6352 VSS.n4012 VSS.n4011 2.2505
R6353 VSS.n4010 VSS.n3228 2.2505
R6354 VSS.n4009 VSS.n4008 2.2505
R6355 VSS.n4007 VSS.n3229 2.2505
R6356 VSS.n4006 VSS.n4005 2.2505
R6357 VSS.n4004 VSS.n3230 2.2505
R6358 VSS.n4003 VSS.n4002 2.2505
R6359 VSS.n4001 VSS.n3231 2.2505
R6360 VSS.n4000 VSS.n3999 2.2505
R6361 VSS.n3998 VSS.n3232 2.2505
R6362 VSS.n3997 VSS.n3996 2.2505
R6363 VSS.n3995 VSS.n3233 2.2505
R6364 VSS.n3994 VSS.n3993 2.2505
R6365 VSS.n3992 VSS.n3234 2.2505
R6366 VSS.n3991 VSS.n3990 2.2505
R6367 VSS.n3989 VSS.n3235 2.2505
R6368 VSS.n3988 VSS.n3987 2.2505
R6369 VSS.n3986 VSS.n3236 2.2505
R6370 VSS.n3985 VSS.n3984 2.2505
R6371 VSS.n3983 VSS.n3237 2.2505
R6372 VSS.n3982 VSS.n3981 2.2505
R6373 VSS.n3980 VSS.n3238 2.2505
R6374 VSS.n3979 VSS.n3978 2.2505
R6375 VSS.n3977 VSS.n3239 2.2505
R6376 VSS.n3976 VSS.n3975 2.2505
R6377 VSS.n3974 VSS.n3240 2.2505
R6378 VSS.n3973 VSS.n3972 2.2505
R6379 VSS.n3971 VSS.n3241 2.2505
R6380 VSS.n3970 VSS.n3969 2.2505
R6381 VSS.n3968 VSS.n3242 2.2505
R6382 VSS.n3967 VSS.n3966 2.2505
R6383 VSS.n3965 VSS.n3243 2.2505
R6384 VSS.n3964 VSS.n3963 2.2505
R6385 VSS.n3962 VSS.n3244 2.2505
R6386 VSS.n3961 VSS.n3960 2.2505
R6387 VSS.n3959 VSS.n3245 2.2505
R6388 VSS.n3958 VSS.n3957 2.2505
R6389 VSS.n3956 VSS.n3246 2.2505
R6390 VSS.n3955 VSS.n3954 2.2505
R6391 VSS.n3953 VSS.n3247 2.2505
R6392 VSS.n3952 VSS.n3951 2.2505
R6393 VSS.n3950 VSS.n3248 2.2505
R6394 VSS.n3949 VSS.n3948 2.2505
R6395 VSS.n3947 VSS.n3249 2.2505
R6396 VSS.n3946 VSS.n3945 2.2505
R6397 VSS.n3944 VSS.n3250 2.2505
R6398 VSS.n3943 VSS.n3942 2.2505
R6399 VSS.n3941 VSS.n3251 2.2505
R6400 VSS.n3940 VSS.n3939 2.2505
R6401 VSS.n3938 VSS.n3252 2.2505
R6402 VSS.n3937 VSS.n3936 2.2505
R6403 VSS.n3935 VSS.n3253 2.2505
R6404 VSS.n3934 VSS.n3933 2.2505
R6405 VSS.n3932 VSS.n3254 2.2505
R6406 VSS.n3931 VSS.n3930 2.2505
R6407 VSS.n3929 VSS.n3255 2.2505
R6408 VSS.n3928 VSS.n3927 2.2505
R6409 VSS.n3926 VSS.n3256 2.2505
R6410 VSS.n3925 VSS.n3924 2.2505
R6411 VSS.n3923 VSS.n3257 2.2505
R6412 VSS.n3922 VSS.n3921 2.2505
R6413 VSS.n3920 VSS.n3258 2.2505
R6414 VSS.n3919 VSS.n3918 2.2505
R6415 VSS.n3917 VSS.n3259 2.2505
R6416 VSS.n3916 VSS.n3915 2.2505
R6417 VSS.n3914 VSS.n3260 2.2505
R6418 VSS.n3913 VSS.n3912 2.2505
R6419 VSS.n3911 VSS.n3261 2.2505
R6420 VSS.n3910 VSS.n3909 2.2505
R6421 VSS.n3908 VSS.n3262 2.2505
R6422 VSS.n3907 VSS.n3906 2.2505
R6423 VSS.n3905 VSS.n3263 2.2505
R6424 VSS.n3904 VSS.n3903 2.2505
R6425 VSS.n3902 VSS.n3264 2.2505
R6426 VSS.n3901 VSS.n3900 2.2505
R6427 VSS.n3899 VSS.n3265 2.2505
R6428 VSS.n3898 VSS.n3897 2.2505
R6429 VSS.n3896 VSS.n3266 2.2505
R6430 VSS.n3895 VSS.n3894 2.2505
R6431 VSS.n3893 VSS.n3267 2.2505
R6432 VSS.n3892 VSS.n3891 2.2505
R6433 VSS.n3890 VSS.n3268 2.2505
R6434 VSS.n3889 VSS.n3888 2.2505
R6435 VSS.n3887 VSS.n3269 2.2505
R6436 VSS.n3886 VSS.n3885 2.2505
R6437 VSS.n3884 VSS.n3270 2.2505
R6438 VSS.n3883 VSS.n3882 2.2505
R6439 VSS.n3881 VSS.n3271 2.2505
R6440 VSS.n3880 VSS.n3879 2.2505
R6441 VSS.n3878 VSS.n3272 2.2505
R6442 VSS.n3877 VSS.n3876 2.2505
R6443 VSS.n3875 VSS.n3273 2.2505
R6444 VSS.n3874 VSS.n3873 2.2505
R6445 VSS.n3872 VSS.n3274 2.2505
R6446 VSS.n3871 VSS.n3870 2.2505
R6447 VSS.n3869 VSS.n3275 2.2505
R6448 VSS.n3868 VSS.n3867 2.2505
R6449 VSS.n3866 VSS.n3276 2.2505
R6450 VSS.n3865 VSS.n3864 2.2505
R6451 VSS.n3863 VSS.n3277 2.2505
R6452 VSS.n3862 VSS.n3861 2.2505
R6453 VSS.n3860 VSS.n3278 2.2505
R6454 VSS.n3859 VSS.n3858 2.2505
R6455 VSS.n3857 VSS.n3279 2.2505
R6456 VSS.n3856 VSS.n3855 2.2505
R6457 VSS.n3854 VSS.n3280 2.2505
R6458 VSS.n3853 VSS.n3852 2.2505
R6459 VSS.n3851 VSS.n3281 2.2505
R6460 VSS.n3850 VSS.n3849 2.2505
R6461 VSS.n3848 VSS.n3282 2.2505
R6462 VSS.n3847 VSS.n3846 2.2505
R6463 VSS.n3845 VSS.n3283 2.2505
R6464 VSS.n3844 VSS.n3843 2.2505
R6465 VSS.n3842 VSS.n3284 2.2505
R6466 VSS.n3841 VSS.n3840 2.2505
R6467 VSS.n3839 VSS.n3285 2.2505
R6468 VSS.n3838 VSS.n3837 2.2505
R6469 VSS.n3836 VSS.n3286 2.2505
R6470 VSS.n3835 VSS.n3834 2.2505
R6471 VSS.n3833 VSS.n3287 2.2505
R6472 VSS.n3832 VSS.n3831 2.2505
R6473 VSS.n3830 VSS.n3288 2.2505
R6474 VSS.n3829 VSS.n3828 2.2505
R6475 VSS.n3827 VSS.n3289 2.2505
R6476 VSS.n3826 VSS.n3825 2.2505
R6477 VSS.n3824 VSS.n3290 2.2505
R6478 VSS.n3823 VSS.n3822 2.2505
R6479 VSS.n3821 VSS.n3291 2.2505
R6480 VSS.n3820 VSS.n3819 2.2505
R6481 VSS.n3818 VSS.n3292 2.2505
R6482 VSS.n3817 VSS.n3816 2.2505
R6483 VSS.n3815 VSS.n3293 2.2505
R6484 VSS.n3814 VSS.n3813 2.2505
R6485 VSS.n3812 VSS.n3294 2.2505
R6486 VSS.n3811 VSS.n3810 2.2505
R6487 VSS.n3809 VSS.n3295 2.2505
R6488 VSS.n3808 VSS.n3807 2.2505
R6489 VSS.n3806 VSS.n3296 2.2505
R6490 VSS.n3805 VSS.n3804 2.2505
R6491 VSS.n3803 VSS.n3297 2.2505
R6492 VSS.n3802 VSS.n3801 2.2505
R6493 VSS.n3800 VSS.n3298 2.2505
R6494 VSS.n3799 VSS.n3798 2.2505
R6495 VSS.n3797 VSS.n3299 2.2505
R6496 VSS.n3796 VSS.n3795 2.2505
R6497 VSS.n3794 VSS.n3300 2.2505
R6498 VSS.n3793 VSS.n3792 2.2505
R6499 VSS.n3791 VSS.n3301 2.2505
R6500 VSS.n3790 VSS.n3789 2.2505
R6501 VSS.n3788 VSS.n3302 2.2505
R6502 VSS.n3787 VSS.n3786 2.2505
R6503 VSS.n3785 VSS.n3303 2.2505
R6504 VSS.n3784 VSS.n3783 2.2505
R6505 VSS.n3782 VSS.n3304 2.2505
R6506 VSS.n3781 VSS.n3780 2.2505
R6507 VSS.n3779 VSS.n3305 2.2505
R6508 VSS.n3778 VSS.n3777 2.2505
R6509 VSS.n3776 VSS.n3306 2.2505
R6510 VSS.n3775 VSS.n3774 2.2505
R6511 VSS.n3773 VSS.n3307 2.2505
R6512 VSS.n3772 VSS.n3771 2.2505
R6513 VSS.n3770 VSS.n3308 2.2505
R6514 VSS.n3769 VSS.n3768 2.2505
R6515 VSS.n3767 VSS.n3309 2.2505
R6516 VSS.n3766 VSS.n3765 2.2505
R6517 VSS.n3764 VSS.n3310 2.2505
R6518 VSS.n3763 VSS.n3762 2.2505
R6519 VSS.n3761 VSS.n3311 2.2505
R6520 VSS.n3760 VSS.n3759 2.2505
R6521 VSS.n3758 VSS.n3312 2.2505
R6522 VSS.n3757 VSS.n3756 2.2505
R6523 VSS.n3755 VSS.n3313 2.2505
R6524 VSS.n3754 VSS.n3753 2.2505
R6525 VSS.n3752 VSS.n3314 2.2505
R6526 VSS.n3751 VSS.n3750 2.2505
R6527 VSS.n3749 VSS.n3315 2.2505
R6528 VSS.n3748 VSS.n3747 2.2505
R6529 VSS.n3746 VSS.n3316 2.2505
R6530 VSS.n3745 VSS.n3744 2.2505
R6531 VSS.n3743 VSS.n3317 2.2505
R6532 VSS.n3742 VSS.n3741 2.2505
R6533 VSS.n3740 VSS.n3318 2.2505
R6534 VSS.n3739 VSS.n3738 2.2505
R6535 VSS.n3737 VSS.n3319 2.2505
R6536 VSS.n3736 VSS.n3735 2.2505
R6537 VSS.n3734 VSS.n3320 2.2505
R6538 VSS.n3733 VSS.n3732 2.2505
R6539 VSS.n3731 VSS.n3321 2.2505
R6540 VSS.n3730 VSS.n3729 2.2505
R6541 VSS.n3728 VSS.n3322 2.2505
R6542 VSS.n3727 VSS.n3726 2.2505
R6543 VSS.n3725 VSS.n3323 2.2505
R6544 VSS.n3724 VSS.n3723 2.2505
R6545 VSS.n3722 VSS.n3324 2.2505
R6546 VSS.n3721 VSS.n3720 2.2505
R6547 VSS.n3719 VSS.n3325 2.2505
R6548 VSS.n3718 VSS.n3717 2.2505
R6549 VSS.n3716 VSS.n3326 2.2505
R6550 VSS.n3715 VSS.n3714 2.2505
R6551 VSS.n3713 VSS.n3327 2.2505
R6552 VSS.n3712 VSS.n3711 2.2505
R6553 VSS.n3710 VSS.n3328 2.2505
R6554 VSS.n3709 VSS.n3708 2.2505
R6555 VSS.n3707 VSS.n3329 2.2505
R6556 VSS.n3706 VSS.n3705 2.2505
R6557 VSS.n3704 VSS.n3330 2.2505
R6558 VSS.n3703 VSS.n3702 2.2505
R6559 VSS.n3701 VSS.n3331 2.2505
R6560 VSS.n3700 VSS.n3699 2.2505
R6561 VSS.n3698 VSS.n3332 2.2505
R6562 VSS.n3697 VSS.n3696 2.2505
R6563 VSS.n3695 VSS.n3333 2.2505
R6564 VSS.n3694 VSS.n3693 2.2505
R6565 VSS.n3692 VSS.n3334 2.2505
R6566 VSS.n3691 VSS.n3690 2.2505
R6567 VSS.n3689 VSS.n3335 2.2505
R6568 VSS.n3688 VSS.n3687 2.2505
R6569 VSS.n3686 VSS.n3336 2.2505
R6570 VSS.n3685 VSS.n3684 2.2505
R6571 VSS.n3683 VSS.n3337 2.2505
R6572 VSS.n3682 VSS.n3681 2.2505
R6573 VSS.n3680 VSS.n3338 2.2505
R6574 VSS.n3679 VSS.n3678 2.2505
R6575 VSS.n3677 VSS.n3339 2.2505
R6576 VSS.n3676 VSS.n3675 2.2505
R6577 VSS.n3674 VSS.n3340 2.2505
R6578 VSS.n3673 VSS.n3672 2.2505
R6579 VSS.n3671 VSS.n3341 2.2505
R6580 VSS.n3670 VSS.n3669 2.2505
R6581 VSS.n3668 VSS.n3342 2.2505
R6582 VSS.n3667 VSS.n3666 2.2505
R6583 VSS.n3665 VSS.n3343 2.2505
R6584 VSS.n3664 VSS.n3663 2.2505
R6585 VSS.n3662 VSS.n3344 2.2505
R6586 VSS.n3661 VSS.n3660 2.2505
R6587 VSS.n3659 VSS.n3345 2.2505
R6588 VSS.n3658 VSS.n3657 2.2505
R6589 VSS.n3656 VSS.n3346 2.2505
R6590 VSS.n3655 VSS.n3654 2.2505
R6591 VSS.n3653 VSS.n3347 2.2505
R6592 VSS.n3652 VSS.n3651 2.2505
R6593 VSS.n3650 VSS.n3348 2.2505
R6594 VSS.n3649 VSS.n3648 2.2505
R6595 VSS.n3647 VSS.n3349 2.2505
R6596 VSS.n3646 VSS.n3645 2.2505
R6597 VSS.n3644 VSS.n3350 2.2505
R6598 VSS.n3643 VSS.n3642 2.2505
R6599 VSS.n3641 VSS.n3351 2.2505
R6600 VSS.n3640 VSS.n3639 2.2505
R6601 VSS.n3638 VSS.n3352 2.2505
R6602 VSS.n3637 VSS.n3636 2.2505
R6603 VSS.n3635 VSS.n3353 2.2505
R6604 VSS.n3634 VSS.n3633 2.2505
R6605 VSS.n3632 VSS.n3354 2.2505
R6606 VSS.n3631 VSS.n3630 2.2505
R6607 VSS.n3629 VSS.n3355 2.2505
R6608 VSS.n3628 VSS.n3627 2.2505
R6609 VSS.n3626 VSS.n3356 2.2505
R6610 VSS.n3625 VSS.n3624 2.2505
R6611 VSS.n3623 VSS.n3357 2.2505
R6612 VSS.n3622 VSS.n3621 2.2505
R6613 VSS.n3620 VSS.n3358 2.2505
R6614 VSS.n3619 VSS.n3618 2.2505
R6615 VSS.n3617 VSS.n3359 2.2505
R6616 VSS.n3616 VSS.n3615 2.2505
R6617 VSS.n3614 VSS.n3360 2.2505
R6618 VSS.n3613 VSS.n3612 2.2505
R6619 VSS.n3611 VSS.n3361 2.2505
R6620 VSS.n3610 VSS.n3609 2.2505
R6621 VSS.n3608 VSS.n3362 2.2505
R6622 VSS.n3607 VSS.n3606 2.2505
R6623 VSS.n3605 VSS.n3363 2.2505
R6624 VSS.n3604 VSS.n3603 2.2505
R6625 VSS.n3602 VSS.n3364 2.2505
R6626 VSS.n3601 VSS.n3600 2.2505
R6627 VSS.n3599 VSS.n3365 2.2505
R6628 VSS.n3598 VSS.n3597 2.2505
R6629 VSS.n3596 VSS.n3366 2.2505
R6630 VSS.n3595 VSS.n3594 2.2505
R6631 VSS.n3593 VSS.n3367 2.2505
R6632 VSS.n3592 VSS.n3591 2.2505
R6633 VSS.n3590 VSS.n3368 2.2505
R6634 VSS.n3589 VSS.n3588 2.2505
R6635 VSS.n3587 VSS.n3369 2.2505
R6636 VSS.n3586 VSS.n3585 2.2505
R6637 VSS.n3584 VSS.n3370 2.2505
R6638 VSS.n3583 VSS.n3582 2.2505
R6639 VSS.n3581 VSS.n3371 2.2505
R6640 VSS.n3580 VSS.n3579 2.2505
R6641 VSS.n3578 VSS.n3372 2.2505
R6642 VSS.n3577 VSS.n3576 2.2505
R6643 VSS.n3575 VSS.n3373 2.2505
R6644 VSS.n3574 VSS.n3573 2.2505
R6645 VSS.n3572 VSS.n3374 2.2505
R6646 VSS.n3571 VSS.n3570 2.2505
R6647 VSS.n3569 VSS.n3375 2.2505
R6648 VSS.n3568 VSS.n3567 2.2505
R6649 VSS.n3566 VSS.n3376 2.2505
R6650 VSS.n3565 VSS.n3564 2.2505
R6651 VSS.n3563 VSS.n3377 2.2505
R6652 VSS.n3562 VSS.n3561 2.2505
R6653 VSS.n3560 VSS.n3378 2.2505
R6654 VSS.n3559 VSS.n3558 2.2505
R6655 VSS.n3557 VSS.n3379 2.2505
R6656 VSS.n3556 VSS.n3555 2.2505
R6657 VSS.n3554 VSS.n3380 2.2505
R6658 VSS.n3553 VSS.n3552 2.2505
R6659 VSS.n3551 VSS.n3381 2.2505
R6660 VSS.n3550 VSS.n3549 2.2505
R6661 VSS.n3548 VSS.n3382 2.2505
R6662 VSS.n3547 VSS.n3546 2.2505
R6663 VSS.n3545 VSS.n3383 2.2505
R6664 VSS.n3544 VSS.n3543 2.2505
R6665 VSS.n3542 VSS.n3384 2.2505
R6666 VSS.n3541 VSS.n3540 2.2505
R6667 VSS.n3539 VSS.n3385 2.2505
R6668 VSS.n3538 VSS.n3537 2.2505
R6669 VSS.n3536 VSS.n3386 2.2505
R6670 VSS.n3535 VSS.n3534 2.2505
R6671 VSS.n3533 VSS.n3387 2.2505
R6672 VSS.n3532 VSS.n3531 2.2505
R6673 VSS.n3530 VSS.n3388 2.2505
R6674 VSS.n3529 VSS.n3528 2.2505
R6675 VSS.n3527 VSS.n3389 2.2505
R6676 VSS.n3526 VSS.n3525 2.2505
R6677 VSS.n3524 VSS.n3390 2.2505
R6678 VSS.n3523 VSS.n3522 2.2505
R6679 VSS.n3521 VSS.n3391 2.2505
R6680 VSS.n3520 VSS.n3519 2.2505
R6681 VSS.n3518 VSS.n3392 2.2505
R6682 VSS.n3517 VSS.n3516 2.2505
R6683 VSS.n3515 VSS.n3393 2.2505
R6684 VSS.n3514 VSS.n3513 2.2505
R6685 VSS.n3512 VSS.n3394 2.2505
R6686 VSS.n3511 VSS.n3510 2.2505
R6687 VSS.n3509 VSS.n3395 2.2505
R6688 VSS.n3508 VSS.n3507 2.2505
R6689 VSS.n3506 VSS.n3396 2.2505
R6690 VSS.n3505 VSS.n3504 2.2505
R6691 VSS.n3503 VSS.n3397 2.2505
R6692 VSS.n3502 VSS.n3501 2.2505
R6693 VSS.n3500 VSS.n3398 2.2505
R6694 VSS.n3499 VSS.n3498 2.2505
R6695 VSS.n3497 VSS.n3399 2.2505
R6696 VSS.n3496 VSS.n3495 2.2505
R6697 VSS.n3494 VSS.n3400 2.2505
R6698 VSS.n3493 VSS.n3492 2.2505
R6699 VSS.n3491 VSS.n3401 2.2505
R6700 VSS.n3490 VSS.n3489 2.2505
R6701 VSS.n3488 VSS.n3402 2.2505
R6702 VSS.n3487 VSS.n3486 2.2505
R6703 VSS.n3485 VSS.n3403 2.2505
R6704 VSS.n3484 VSS.n3483 2.2505
R6705 VSS.n3482 VSS.n3404 2.2505
R6706 VSS.n3481 VSS.n3480 2.2505
R6707 VSS.n3479 VSS.n3405 2.2505
R6708 VSS.n3478 VSS.n3477 2.2505
R6709 VSS.n3476 VSS.n3406 2.2505
R6710 VSS.n3475 VSS.n3474 2.2505
R6711 VSS.n3473 VSS.n3407 2.2505
R6712 VSS.n3472 VSS.n3471 2.2505
R6713 VSS.n3470 VSS.n3408 2.2505
R6714 VSS.n3469 VSS.n3468 2.2505
R6715 VSS.n3467 VSS.n3409 2.2505
R6716 VSS.n3466 VSS.n3465 2.2505
R6717 VSS.n3464 VSS.n3410 2.2505
R6718 VSS.n3463 VSS.n3462 2.2505
R6719 VSS.n3461 VSS.n3411 2.2505
R6720 VSS.n3460 VSS.n3459 2.2505
R6721 VSS.n3458 VSS.n3412 2.2505
R6722 VSS.n3457 VSS.n3456 2.2505
R6723 VSS.n3455 VSS.n3413 2.2505
R6724 VSS.n3454 VSS.n3453 2.2505
R6725 VSS.n3452 VSS.n3414 2.2505
R6726 VSS.n3451 VSS.n3450 2.2505
R6727 VSS.n3449 VSS.n3415 2.2505
R6728 VSS.n3448 VSS.n3447 2.2505
R6729 VSS.n3446 VSS.n3416 2.2505
R6730 VSS.n3445 VSS.n3444 2.2505
R6731 VSS.n3443 VSS.n3417 2.2505
R6732 VSS.n3442 VSS.n3441 2.2505
R6733 VSS.n3440 VSS.n3418 2.2505
R6734 VSS.n3439 VSS.n3438 2.2505
R6735 VSS.n3437 VSS.n3419 2.2505
R6736 VSS.n3436 VSS.n3435 2.2505
R6737 VSS.n3434 VSS.n3420 2.2505
R6738 VSS.n3433 VSS.n3432 2.2505
R6739 VSS.n3431 VSS.n3421 2.2505
R6740 VSS.n3430 VSS.n3429 2.2505
R6741 VSS.n3428 VSS.n3422 2.2505
R6742 VSS.n3427 VSS.n3426 2.2505
R6743 VSS.n3425 VSS.n3423 2.2505
R6744 VSS.n3424 VSS.n1581 2.2505
R6745 VSS.n8951 VSS.n1582 2.2505
R6746 VSS.n8950 VSS.n8949 2.2505
R6747 VSS.n8948 VSS.n1583 2.2505
R6748 VSS.n8947 VSS.n8946 2.2505
R6749 VSS.n8945 VSS.n1584 2.2505
R6750 VSS.n8944 VSS.n8943 2.2505
R6751 VSS.n8942 VSS.n1585 2.2505
R6752 VSS.n8941 VSS.n8940 2.2505
R6753 VSS.n8939 VSS.n1586 2.2505
R6754 VSS.n8938 VSS.n8937 2.2505
R6755 VSS.n8936 VSS.n1587 2.2505
R6756 VSS.n8935 VSS.n8934 2.2505
R6757 VSS.n8933 VSS.n1588 2.2505
R6758 VSS.n8932 VSS.n8931 2.2505
R6759 VSS.n8930 VSS.n1589 2.2505
R6760 VSS.n8929 VSS.n8928 2.2505
R6761 VSS.n8927 VSS.n1590 2.2505
R6762 VSS.n8926 VSS.n8925 2.2505
R6763 VSS.n8924 VSS.n1591 2.2505
R6764 VSS.n8923 VSS.n8922 2.2505
R6765 VSS.n8921 VSS.n1592 2.2505
R6766 VSS.n8920 VSS.n8919 2.2505
R6767 VSS.n8918 VSS.n1593 2.2505
R6768 VSS.n8917 VSS.n8916 2.2505
R6769 VSS.n8915 VSS.n1594 2.2505
R6770 VSS.n8914 VSS.n8913 2.2505
R6771 VSS.n8912 VSS.n1595 2.2505
R6772 VSS.n8911 VSS.n8910 2.2505
R6773 VSS.n8909 VSS.n1596 2.2505
R6774 VSS.n8908 VSS.n8907 2.2505
R6775 VSS.n8906 VSS.n1597 2.2505
R6776 VSS.n8905 VSS.n8904 2.2505
R6777 VSS.n8903 VSS.n1598 2.2505
R6778 VSS.n8902 VSS.n8901 2.2505
R6779 VSS.n8900 VSS.n1599 2.2505
R6780 VSS.n8899 VSS.n8898 2.2505
R6781 VSS.n8897 VSS.n1600 2.2505
R6782 VSS.n8896 VSS.n8895 2.2505
R6783 VSS.n8894 VSS.n1601 2.2505
R6784 VSS.n8893 VSS.n8892 2.2505
R6785 VSS.n8891 VSS.n1602 2.2505
R6786 VSS.n8890 VSS.n8889 2.2505
R6787 VSS.n8888 VSS.n1603 2.2505
R6788 VSS.n8887 VSS.n8886 2.2505
R6789 VSS.n8885 VSS.n1604 2.2505
R6790 VSS.n8884 VSS.n8883 2.2505
R6791 VSS.n8882 VSS.n1605 2.2505
R6792 VSS.n8881 VSS.n8880 2.2505
R6793 VSS.n8879 VSS.n1606 2.2505
R6794 VSS.n8878 VSS.n8877 2.2505
R6795 VSS.n8876 VSS.n1607 2.2505
R6796 VSS.n8875 VSS.n8874 2.2505
R6797 VSS.n8873 VSS.n1608 2.2505
R6798 VSS.n8872 VSS.n8871 2.2505
R6799 VSS.n8870 VSS.n1609 2.2505
R6800 VSS.n8869 VSS.n8868 2.2505
R6801 VSS.n8867 VSS.n1610 2.2505
R6802 VSS.n8866 VSS.n8865 2.2505
R6803 VSS.n8864 VSS.n1611 2.2505
R6804 VSS.n8863 VSS.n8862 2.2505
R6805 VSS.n8861 VSS.n1612 2.2505
R6806 VSS.n8860 VSS.n8859 2.2505
R6807 VSS.n8858 VSS.n1613 2.2505
R6808 VSS.n8857 VSS.n8856 2.2505
R6809 VSS.n8855 VSS.n1614 2.2505
R6810 VSS.n8854 VSS.n8853 2.2505
R6811 VSS.n8852 VSS.n1615 2.2505
R6812 VSS.n8851 VSS.n8850 2.2505
R6813 VSS.n8849 VSS.n1616 2.2505
R6814 VSS.n8848 VSS.n8847 2.2505
R6815 VSS.n8846 VSS.n1617 2.2505
R6816 VSS.n8845 VSS.n8844 2.2505
R6817 VSS.n8843 VSS.n1618 2.2505
R6818 VSS.n8842 VSS.n8841 2.2505
R6819 VSS.n8840 VSS.n1619 2.2505
R6820 VSS.n8839 VSS.n8838 2.2505
R6821 VSS.n8837 VSS.n1620 2.2505
R6822 VSS.n8836 VSS.n8835 2.2505
R6823 VSS.n8834 VSS.n1621 2.2505
R6824 VSS.n8833 VSS.n8832 2.2505
R6825 VSS.n8831 VSS.n1622 2.2505
R6826 VSS.n8830 VSS.n8829 2.2505
R6827 VSS.n8828 VSS.n1623 2.2505
R6828 VSS.n8827 VSS.n8826 2.2505
R6829 VSS.n8825 VSS.n1624 2.2505
R6830 VSS.n8824 VSS.n8823 2.2505
R6831 VSS.n8822 VSS.n1625 2.2505
R6832 VSS.n8821 VSS.n8820 2.2505
R6833 VSS.n8819 VSS.n1626 2.2505
R6834 VSS.n8818 VSS.n8817 2.2505
R6835 VSS.n8816 VSS.n1627 2.2505
R6836 VSS.n8815 VSS.n8814 2.2505
R6837 VSS.n8813 VSS.n1628 2.2505
R6838 VSS.n8812 VSS.n8811 2.2505
R6839 VSS.n8810 VSS.n1629 2.2505
R6840 VSS.n8809 VSS.n8808 2.2505
R6841 VSS.n8807 VSS.n1630 2.2505
R6842 VSS.n8806 VSS.n8805 2.2505
R6843 VSS.n8804 VSS.n1631 2.2505
R6844 VSS.n8803 VSS.n8802 2.2505
R6845 VSS.n8801 VSS.n1632 2.2505
R6846 VSS.n8800 VSS.n8799 2.2505
R6847 VSS.n8798 VSS.n1633 2.2505
R6848 VSS.n8797 VSS.n8796 2.2505
R6849 VSS.n8795 VSS.n1634 2.2505
R6850 VSS.n8794 VSS.n8793 2.2505
R6851 VSS.n8792 VSS.n1635 2.2505
R6852 VSS.n8791 VSS.n8790 2.2505
R6853 VSS.n8789 VSS.n1636 2.2505
R6854 VSS.n8788 VSS.n8787 2.2505
R6855 VSS.n8786 VSS.n1637 2.2505
R6856 VSS.n8785 VSS.n8784 2.2505
R6857 VSS.n8783 VSS.n1638 2.2505
R6858 VSS.n8782 VSS.n8781 2.2505
R6859 VSS.n8780 VSS.n1639 2.2505
R6860 VSS.n8779 VSS.n8778 2.2505
R6861 VSS.n8777 VSS.n1640 2.2505
R6862 VSS.n8776 VSS.n8775 2.2505
R6863 VSS.n8774 VSS.n1641 2.2505
R6864 VSS.n8773 VSS.n8772 2.2505
R6865 VSS.n8771 VSS.n1642 2.2505
R6866 VSS.n8770 VSS.n8769 2.2505
R6867 VSS.n8768 VSS.n1643 2.2505
R6868 VSS.n8767 VSS.n8766 2.2505
R6869 VSS.n8765 VSS.n1644 2.2505
R6870 VSS.n8764 VSS.n8763 2.2505
R6871 VSS.n8762 VSS.n1645 2.2505
R6872 VSS.n8761 VSS.n8760 2.2505
R6873 VSS.n8759 VSS.n1646 2.2505
R6874 VSS.n8758 VSS.n8757 2.2505
R6875 VSS.n8756 VSS.n1647 2.2505
R6876 VSS.n8755 VSS.n8754 2.2505
R6877 VSS.n8753 VSS.n1648 2.2505
R6878 VSS.n8752 VSS.n8751 2.2505
R6879 VSS.n8750 VSS.n1649 2.2505
R6880 VSS.n8749 VSS.n8748 2.2505
R6881 VSS.n8747 VSS.n1650 2.2505
R6882 VSS.n8746 VSS.n8745 2.2505
R6883 VSS.n8744 VSS.n1651 2.2505
R6884 VSS.n8743 VSS.n8742 2.2505
R6885 VSS.n8741 VSS.n1652 2.2505
R6886 VSS.n8740 VSS.n8739 2.2505
R6887 VSS.n8738 VSS.n1653 2.2505
R6888 VSS.n8737 VSS.n8736 2.2505
R6889 VSS.n8735 VSS.n1654 2.2505
R6890 VSS.n8734 VSS.n8733 2.2505
R6891 VSS.n8732 VSS.n1655 2.2505
R6892 VSS.n8731 VSS.n8730 2.2505
R6893 VSS.n8729 VSS.n1656 2.2505
R6894 VSS.n8728 VSS.n8727 2.2505
R6895 VSS.n8726 VSS.n1657 2.2505
R6896 VSS.n8725 VSS.n8724 2.2505
R6897 VSS.n8723 VSS.n1658 2.2505
R6898 VSS.n8722 VSS.n8721 2.2505
R6899 VSS.n8720 VSS.n1659 2.2505
R6900 VSS.n8719 VSS.n8718 2.2505
R6901 VSS.n8717 VSS.n1660 2.2505
R6902 VSS.n8716 VSS.n8715 2.2505
R6903 VSS.n8714 VSS.n1661 2.2505
R6904 VSS.n8713 VSS.n8712 2.2505
R6905 VSS.n8711 VSS.n1662 2.2505
R6906 VSS.n8710 VSS.n8709 2.2505
R6907 VSS.n8708 VSS.n1663 2.2505
R6908 VSS.n8707 VSS.n8706 2.2505
R6909 VSS.n8705 VSS.n1664 2.2505
R6910 VSS.n8704 VSS.n8703 2.2505
R6911 VSS.n8702 VSS.n1665 2.2505
R6912 VSS.n8701 VSS.n8700 2.2505
R6913 VSS.n8699 VSS.n1666 2.2505
R6914 VSS.n8698 VSS.n8697 2.2505
R6915 VSS.n8696 VSS.n1667 2.2505
R6916 VSS.n8695 VSS.n8694 2.2505
R6917 VSS.n8693 VSS.n1668 2.2505
R6918 VSS.n8692 VSS.n8691 2.2505
R6919 VSS.n8690 VSS.n1669 2.2505
R6920 VSS.n8689 VSS.n8688 2.2505
R6921 VSS.n8687 VSS.n1670 2.2505
R6922 VSS.n8686 VSS.n8685 2.2505
R6923 VSS.n8684 VSS.n1671 2.2505
R6924 VSS.n8683 VSS.n8682 2.2505
R6925 VSS.n8681 VSS.n1672 2.2505
R6926 VSS.n8680 VSS.n8679 2.2505
R6927 VSS.n8678 VSS.n1673 2.2505
R6928 VSS.n8677 VSS.n8676 2.2505
R6929 VSS.n8675 VSS.n1674 2.2505
R6930 VSS.n8674 VSS.n8673 2.2505
R6931 VSS.n8672 VSS.n1675 2.2505
R6932 VSS.n8671 VSS.n8670 2.2505
R6933 VSS.n8669 VSS.n1676 2.2505
R6934 VSS.n8668 VSS.n8667 2.2505
R6935 VSS.n8666 VSS.n1677 2.2505
R6936 VSS.n8665 VSS.n8664 2.2505
R6937 VSS.n8663 VSS.n1678 2.2505
R6938 VSS.n8662 VSS.n8661 2.2505
R6939 VSS.n8660 VSS.n1679 2.2505
R6940 VSS.n8659 VSS.n8658 2.2505
R6941 VSS.n8657 VSS.n1680 2.2505
R6942 VSS.n8656 VSS.n8655 2.2505
R6943 VSS.n8654 VSS.n1681 2.2505
R6944 VSS.n8653 VSS.n8652 2.2505
R6945 VSS.n8651 VSS.n1682 2.2505
R6946 VSS.n8650 VSS.n8649 2.2505
R6947 VSS.n8648 VSS.n1683 2.2505
R6948 VSS.n8647 VSS.n8646 2.2505
R6949 VSS.n8645 VSS.n1684 2.2505
R6950 VSS.n8644 VSS.n8643 2.2505
R6951 VSS.n8642 VSS.n1685 2.2505
R6952 VSS.n8641 VSS.n8640 2.2505
R6953 VSS.n8639 VSS.n1686 2.2505
R6954 VSS.n8638 VSS.n8637 2.2505
R6955 VSS.n8636 VSS.n1687 2.2505
R6956 VSS.n8635 VSS.n8634 2.2505
R6957 VSS.n8633 VSS.n1688 2.2505
R6958 VSS.n8632 VSS.n8631 2.2505
R6959 VSS.n8630 VSS.n1689 2.2505
R6960 VSS.n8629 VSS.n8628 2.2505
R6961 VSS.n8627 VSS.n1690 2.2505
R6962 VSS.n8626 VSS.n8625 2.2505
R6963 VSS.n8624 VSS.n1691 2.2505
R6964 VSS.n8623 VSS.n8622 2.2505
R6965 VSS.n8621 VSS.n1692 2.2505
R6966 VSS.n8620 VSS.n8619 2.2505
R6967 VSS.n8618 VSS.n1693 2.2505
R6968 VSS.n8617 VSS.n8616 2.2505
R6969 VSS.n8615 VSS.n1694 2.2505
R6970 VSS.n8614 VSS.n8613 2.2505
R6971 VSS.n8612 VSS.n1695 2.2505
R6972 VSS.n8611 VSS.n8610 2.2505
R6973 VSS.n8609 VSS.n1696 2.2505
R6974 VSS.n8608 VSS.n8607 2.2505
R6975 VSS.n8606 VSS.n1697 2.2505
R6976 VSS.n8605 VSS.n8604 2.2505
R6977 VSS.n8603 VSS.n1698 2.2505
R6978 VSS.n8602 VSS.n8601 2.2505
R6979 VSS.n8600 VSS.n1699 2.2505
R6980 VSS.n8599 VSS.n8598 2.2505
R6981 VSS.n8597 VSS.n1700 2.2505
R6982 VSS.n8596 VSS.n8595 2.2505
R6983 VSS.n8594 VSS.n1701 2.2505
R6984 VSS.n8593 VSS.n8592 2.2505
R6985 VSS.n8591 VSS.n1702 2.2505
R6986 VSS.n8590 VSS.n8589 2.2505
R6987 VSS.n8588 VSS.n1703 2.2505
R6988 VSS.n8587 VSS.n8586 2.2505
R6989 VSS.n8585 VSS.n1704 2.2505
R6990 VSS.n8584 VSS.n8583 2.2505
R6991 VSS.n8582 VSS.n1705 2.2505
R6992 VSS.n8581 VSS.n8580 2.2505
R6993 VSS.n8579 VSS.n1706 2.2505
R6994 VSS.n8578 VSS.n8577 2.2505
R6995 VSS.n8576 VSS.n1707 2.2505
R6996 VSS.n8575 VSS.n8574 2.2505
R6997 VSS.n8573 VSS.n1708 2.2505
R6998 VSS.n8572 VSS.n8571 2.2505
R6999 VSS.n8570 VSS.n1709 2.2505
R7000 VSS.n8569 VSS.n8568 2.2505
R7001 VSS.n8567 VSS.n1710 2.2505
R7002 VSS.n8566 VSS.n8565 2.2505
R7003 VSS.n8564 VSS.n1711 2.2505
R7004 VSS.n8563 VSS.n8562 2.2505
R7005 VSS.n8561 VSS.n1712 2.2505
R7006 VSS.n8560 VSS.n8559 2.2505
R7007 VSS.n8558 VSS.n1713 2.2505
R7008 VSS.n8557 VSS.n8556 2.2505
R7009 VSS.n8555 VSS.n1714 2.2505
R7010 VSS.n8554 VSS.n8553 2.2505
R7011 VSS.n8552 VSS.n1715 2.2505
R7012 VSS.n8551 VSS.n8550 2.2505
R7013 VSS.n8549 VSS.n1716 2.2505
R7014 VSS.n8548 VSS.n8547 2.2505
R7015 VSS.n8546 VSS.n1717 2.2505
R7016 VSS.n8545 VSS.n8544 2.2505
R7017 VSS.n8543 VSS.n1718 2.2505
R7018 VSS.n8542 VSS.n8541 2.2505
R7019 VSS.n8540 VSS.n1719 2.2505
R7020 VSS.n8539 VSS.n8538 2.2505
R7021 VSS.n8537 VSS.n1720 2.2505
R7022 VSS.n8536 VSS.n8535 2.2505
R7023 VSS.n8534 VSS.n1721 2.2505
R7024 VSS.n8533 VSS.n8532 2.2505
R7025 VSS.n8531 VSS.n1722 2.2505
R7026 VSS.n8530 VSS.n8529 2.2505
R7027 VSS.n8528 VSS.n1723 2.2505
R7028 VSS.n8527 VSS.n8526 2.2505
R7029 VSS.n8525 VSS.n1724 2.2505
R7030 VSS.n8524 VSS.n8523 2.2505
R7031 VSS.n8522 VSS.n1725 2.2505
R7032 VSS.n8521 VSS.n8520 2.2505
R7033 VSS.n8519 VSS.n1726 2.2505
R7034 VSS.n8518 VSS.n8517 2.2505
R7035 VSS.n8516 VSS.n1727 2.2505
R7036 VSS.n8515 VSS.n8514 2.2505
R7037 VSS.n8513 VSS.n1728 2.2505
R7038 VSS.n8512 VSS.n8511 2.2505
R7039 VSS.n8510 VSS.n1729 2.2505
R7040 VSS.n8509 VSS.n8508 2.2505
R7041 VSS.n8507 VSS.n1730 2.2505
R7042 VSS.n8506 VSS.n8505 2.2505
R7043 VSS.n8504 VSS.n1731 2.2505
R7044 VSS.n8503 VSS.n8502 2.2505
R7045 VSS.n8501 VSS.n1732 2.2505
R7046 VSS.n8500 VSS.n8499 2.2505
R7047 VSS.n8498 VSS.n1733 2.2505
R7048 VSS.n8497 VSS.n8496 2.2505
R7049 VSS.n8495 VSS.n1734 2.2505
R7050 VSS.n8494 VSS.n8493 2.2505
R7051 VSS.n8492 VSS.n1735 2.2505
R7052 VSS.n8491 VSS.n8490 2.2505
R7053 VSS.n8489 VSS.n1736 2.2505
R7054 VSS.n8488 VSS.n8487 2.2505
R7055 VSS.n8486 VSS.n1737 2.2505
R7056 VSS.n8485 VSS.n8484 2.2505
R7057 VSS.n8483 VSS.n1738 2.2505
R7058 VSS.n8482 VSS.n8481 2.2505
R7059 VSS.n8480 VSS.n1739 2.2505
R7060 VSS.n8479 VSS.n8478 2.2505
R7061 VSS.n8477 VSS.n1740 2.2505
R7062 VSS.n8476 VSS.n8475 2.2505
R7063 VSS.n8474 VSS.n1741 2.2505
R7064 VSS.n8473 VSS.n8472 2.2505
R7065 VSS.n8471 VSS.n1742 2.2505
R7066 VSS.n8470 VSS.n8469 2.2505
R7067 VSS.n8468 VSS.n1743 2.2505
R7068 VSS.n8467 VSS.n8466 2.2505
R7069 VSS.n8465 VSS.n1744 2.2505
R7070 VSS.n8464 VSS.n8463 2.2505
R7071 VSS.n8462 VSS.n1745 2.2505
R7072 VSS.n8461 VSS.n8460 2.2505
R7073 VSS.n8459 VSS.n1746 2.2505
R7074 VSS.n8458 VSS.n8457 2.2505
R7075 VSS.n8456 VSS.n1747 2.2505
R7076 VSS.n8455 VSS.n8454 2.2505
R7077 VSS.n8453 VSS.n1748 2.2505
R7078 VSS.n8452 VSS.n8451 2.2505
R7079 VSS.n8450 VSS.n1749 2.2505
R7080 VSS.n8449 VSS.n8448 2.2505
R7081 VSS.n8447 VSS.n1750 2.2505
R7082 VSS.n8446 VSS.n8445 2.2505
R7083 VSS.n8444 VSS.n1751 2.2505
R7084 VSS.n8443 VSS.n8442 2.2505
R7085 VSS.n8441 VSS.n1752 2.2505
R7086 VSS.n8440 VSS.n8439 2.2505
R7087 VSS.n8438 VSS.n1753 2.2505
R7088 VSS.n8437 VSS.n8436 2.2505
R7089 VSS.n8435 VSS.n1754 2.2505
R7090 VSS.n8434 VSS.n8433 2.2505
R7091 VSS.n8432 VSS.n1755 2.2505
R7092 VSS.n8431 VSS.n8430 2.2505
R7093 VSS.n8429 VSS.n1756 2.2505
R7094 VSS.n8428 VSS.n8427 2.2505
R7095 VSS.n8426 VSS.n1757 2.2505
R7096 VSS.n8425 VSS.n8424 2.2505
R7097 VSS.n8423 VSS.n1758 2.2505
R7098 VSS.n8422 VSS.n8421 2.2505
R7099 VSS.n8420 VSS.n1759 2.2505
R7100 VSS.n8419 VSS.n8418 2.2505
R7101 VSS.n8417 VSS.n1760 2.2505
R7102 VSS.n8416 VSS.n8415 2.2505
R7103 VSS.n8414 VSS.n1761 2.2505
R7104 VSS.n8413 VSS.n8412 2.2505
R7105 VSS.n8411 VSS.n1762 2.2505
R7106 VSS.n8410 VSS.n8409 2.2505
R7107 VSS.n8408 VSS.n1763 2.2505
R7108 VSS.n8407 VSS.n8406 2.2505
R7109 VSS.n8405 VSS.n1764 2.2505
R7110 VSS.n8404 VSS.n8403 2.2505
R7111 VSS.n8402 VSS.n1765 2.2505
R7112 VSS.n8401 VSS.n8400 2.2505
R7113 VSS.n8399 VSS.n1766 2.2505
R7114 VSS.n8398 VSS.n8397 2.2505
R7115 VSS.n8396 VSS.n1767 2.2505
R7116 VSS.n8395 VSS.n8394 2.2505
R7117 VSS.n8393 VSS.n1768 2.2505
R7118 VSS.n8392 VSS.n8391 2.2505
R7119 VSS.n8390 VSS.n1769 2.2505
R7120 VSS.n8389 VSS.n8388 2.2505
R7121 VSS.n8387 VSS.n1770 2.2505
R7122 VSS.n8386 VSS.n8385 2.2505
R7123 VSS.n8384 VSS.n1771 2.2505
R7124 VSS.n8383 VSS.n8382 2.2505
R7125 VSS.n8381 VSS.n1772 2.2505
R7126 VSS.n8380 VSS.n8379 2.2505
R7127 VSS.n8378 VSS.n1773 2.2505
R7128 VSS.n8377 VSS.n8376 2.2505
R7129 VSS.n8375 VSS.n1774 2.2505
R7130 VSS.n8374 VSS.n8373 2.2505
R7131 VSS.n8372 VSS.n1775 2.2505
R7132 VSS.n8371 VSS.n8370 2.2505
R7133 VSS.n8369 VSS.n1776 2.2505
R7134 VSS.n8368 VSS.n8367 2.2505
R7135 VSS.n8366 VSS.n1777 2.2505
R7136 VSS.n8365 VSS.n8364 2.2505
R7137 VSS.n8363 VSS.n1778 2.2505
R7138 VSS.n8362 VSS.n8361 2.2505
R7139 VSS.n8360 VSS.n1779 2.2505
R7140 VSS.n8359 VSS.n8358 2.2505
R7141 VSS.n8357 VSS.n1780 2.2505
R7142 VSS.n8356 VSS.n8355 2.2505
R7143 VSS.n8354 VSS.n1781 2.2505
R7144 VSS.n8353 VSS.n8352 2.2505
R7145 VSS.n8351 VSS.n1782 2.2505
R7146 VSS.n8350 VSS.n8349 2.2505
R7147 VSS.n8348 VSS.n1783 2.2505
R7148 VSS.n8347 VSS.n8346 2.2505
R7149 VSS.n8345 VSS.n1784 2.2505
R7150 VSS.n8344 VSS.n8343 2.2505
R7151 VSS.n8342 VSS.n1785 2.2505
R7152 VSS.n8341 VSS.n8340 2.2505
R7153 VSS.n8339 VSS.n1786 2.2505
R7154 VSS.n8338 VSS.n8337 2.2505
R7155 VSS.n8336 VSS.n1787 2.2505
R7156 VSS.n8335 VSS.n8334 2.2505
R7157 VSS.n8333 VSS.n1788 2.2505
R7158 VSS.n8332 VSS.n8331 2.2505
R7159 VSS.n8330 VSS.n1789 2.2505
R7160 VSS.n8329 VSS.n8328 2.2505
R7161 VSS.n8327 VSS.n1790 2.2505
R7162 VSS.n8326 VSS.n8325 2.2505
R7163 VSS.n8324 VSS.n1791 2.2505
R7164 VSS.n8323 VSS.n8322 2.2505
R7165 VSS.n8321 VSS.n1792 2.2505
R7166 VSS.n8320 VSS.n8319 2.2505
R7167 VSS.n8318 VSS.n1793 2.2505
R7168 VSS.n8317 VSS.n8316 2.2505
R7169 VSS.n8315 VSS.n1794 2.2505
R7170 VSS.n8314 VSS.n8313 2.2505
R7171 VSS.n8312 VSS.n1795 2.2505
R7172 VSS.n8311 VSS.n8310 2.2505
R7173 VSS.n8309 VSS.n1796 2.2505
R7174 VSS.n8308 VSS.n8307 2.2505
R7175 VSS.n8306 VSS.n1797 2.2505
R7176 VSS.n8305 VSS.n8304 2.2505
R7177 VSS.n8303 VSS.n1798 2.2505
R7178 VSS.n8302 VSS.n8301 2.2505
R7179 VSS.n8300 VSS.n1799 2.2505
R7180 VSS.n8299 VSS.n8298 2.2505
R7181 VSS.n8297 VSS.n1800 2.2505
R7182 VSS.n8296 VSS.n8295 2.2505
R7183 VSS.n8294 VSS.n1801 2.2505
R7184 VSS.n8293 VSS.n8292 2.2505
R7185 VSS.n8291 VSS.n1802 2.2505
R7186 VSS.n8290 VSS.n8289 2.2505
R7187 VSS.n8288 VSS.n1803 2.2505
R7188 VSS.n8287 VSS.n8286 2.2505
R7189 VSS.n8285 VSS.n1804 2.2505
R7190 VSS.n8284 VSS.n8283 2.2505
R7191 VSS.n8282 VSS.n1805 2.2505
R7192 VSS.n8281 VSS.n8280 2.2505
R7193 VSS.n8279 VSS.n1806 2.2505
R7194 VSS.n8278 VSS.n8277 2.2505
R7195 VSS.n8276 VSS.n1807 2.2505
R7196 VSS.n8275 VSS.n8274 2.2505
R7197 VSS.n8273 VSS.n1808 2.2505
R7198 VSS.n8272 VSS.n8271 2.2505
R7199 VSS.n8270 VSS.n1809 2.2505
R7200 VSS.n8269 VSS.n8268 2.2505
R7201 VSS.n8267 VSS.n1810 2.2505
R7202 VSS.n8266 VSS.n8265 2.2505
R7203 VSS.n8264 VSS.n1811 2.2505
R7204 VSS.n8263 VSS.n8262 2.2505
R7205 VSS.n8261 VSS.n1812 2.2505
R7206 VSS.n8260 VSS.n8259 2.2505
R7207 VSS.n8258 VSS.n1813 2.2505
R7208 VSS.n8257 VSS.n8256 2.2505
R7209 VSS.n8255 VSS.n1814 2.2505
R7210 VSS.n8254 VSS.n8253 2.2505
R7211 VSS.n8252 VSS.n1815 2.2505
R7212 VSS.n8251 VSS.n8250 2.2505
R7213 VSS.n8249 VSS.n1816 2.2505
R7214 VSS.n8248 VSS.n8247 2.2505
R7215 VSS.n8246 VSS.n1817 2.2505
R7216 VSS.n8245 VSS.n8244 2.2505
R7217 VSS.n8243 VSS.n1818 2.2505
R7218 VSS.n8242 VSS.n8241 2.2505
R7219 VSS.n8240 VSS.n1819 2.2505
R7220 VSS.n8239 VSS.n8238 2.2505
R7221 VSS.n8237 VSS.n1820 2.2505
R7222 VSS.n8236 VSS.n8235 2.2505
R7223 VSS.n8234 VSS.n1821 2.2505
R7224 VSS.n8233 VSS.n8232 2.2505
R7225 VSS.n36 VSS.n35 2.25016
R7226 VSS.n58 VSS.n54 2.25016
R7227 VSS.n11395 VSS.n11394 2.25016
R7228 VSS.n11312 VSS.n123 2.2497
R7229 VSS.n10705 VSS.n10703 2.24949
R7230 VSS.n111 VSS.n105 2.24922
R7231 VSS.n10567 VSS.n10566 2.24813
R7232 VSS.n10570 VSS.n10568 2.24218
R7233 VSS.n10572 VSS.n10562 2.24218
R7234 VSS.n10564 VSS.n10556 2.24218
R7235 VSS.n227 VSS.n223 2.24218
R7236 VSS.n10910 VSS.n230 2.24218
R7237 VSS.n10911 VSS.n10910 2.24218
R7238 VSS.n107 VSS.n103 2.24218
R7239 VSS.n110 VSS.n103 2.24218
R7240 VSS.n11431 VSS.n37 2.24218
R7241 VSS.n11429 VSS.n33 2.24218
R7242 VSS.n11433 VSS.n29 2.24218
R7243 VSS.n11400 VSS.n55 2.24218
R7244 VSS.n11398 VSS.n11397 2.24218
R7245 VSS.n11385 VSS.n11384 2.24218
R7246 VSS.n11384 VSS.n79 2.24218
R7247 VSS.n82 VSS.n78 2.24218
R7248 VSS.n11311 VSS.n11310 2.24218
R7249 VSS.n11310 VSS.n126 2.24218
R7250 VSS.n11306 VSS.n11305 2.24218
R7251 VSS.n10732 VSS.n10700 2.24218
R7252 VSS.n10732 VSS.n10699 2.24218
R7253 VSS.n10728 VSS.n10702 2.24218
R7254 VSS.n10334 VSS.n10309 2.23722
R7255 VSS.n10804 VSS.n10803 2.15932
R7256 VSS.n10798 VSS.n10797 2.15932
R7257 VSS.n10806 VSS.n10805 2.15458
R7258 VSS.n10800 VSS.n10799 2.15458
R7259 VSS.n10411 VSS.n10398 2.13932
R7260 VSS.n10767 VSS.t660 2.1005
R7261 VSS.t564 VSS.n10767 2.1005
R7262 VSS.n10756 VSS.t790 2.1005
R7263 VSS.n10756 VSS.t719 2.1005
R7264 VSS.n10474 VSS.n10473 2.1005
R7265 VSS.n10471 VSS.n10470 2.1005
R7266 VSS.n10467 VSS.n10466 2.1005
R7267 VSS.n10463 VSS.n10462 2.1005
R7268 VSS.n10459 VSS.n10458 2.1005
R7269 VSS.n10456 VSS.n10455 2.1005
R7270 VSS.n9072 VSS.n9071 2.1005
R7271 VSS.n9066 VSS.n9065 2.1005
R7272 VSS.n9043 VSS.n9042 2.1005
R7273 VSS.n9087 VSS.n9086 2.1005
R7274 VSS.n8978 VSS.n8977 2.1005
R7275 VSS.n9098 VSS.n9097 2.1005
R7276 VSS.n8968 VSS.n8967 2.1005
R7277 VSS.n9006 VSS.n9005 2.1005
R7278 VSS.n1569 VSS.n1568 2.1005
R7279 VSS.n9037 VSS.n9036 2.1005
R7280 VSS.n841 VSS.n840 2.1005
R7281 VSS.n10925 VSS.n10924 2.1005
R7282 VSS.n876 VSS.n875 2.1005
R7283 VSS.n865 VSS.n864 2.1005
R7284 VSS.n1123 VSS.n1122 2.1005
R7285 VSS.n1129 VSS.n1128 2.1005
R7286 VSS.n1111 VSS.n1110 2.1005
R7287 VSS.n1117 VSS.n1116 2.1005
R7288 VSS.n1090 VSS.n1089 2.1005
R7289 VSS.n1096 VSS.n1095 2.1005
R7290 VSS.n1287 VSS.n1286 2.1005
R7291 VSS.n1293 VSS.n1292 2.1005
R7292 VSS.n10156 VSS.n10155 2.1005
R7293 VSS.n10150 VSS.n10149 2.1005
R7294 VSS.n1074 VSS.n1073 2.1005
R7295 VSS.n1080 VSS.n1079 2.1005
R7296 VSS.n1053 VSS.n1052 2.1005
R7297 VSS.n1059 VSS.n1058 2.1005
R7298 VSS.n389 VSS.n388 2.1005
R7299 VSS.n10162 VSS.n10161 2.1005
R7300 VSS.n368 VSS.n367 2.1005
R7301 VSS.n374 VSS.n373 2.1005
R7302 VSS.n1041 VSS.n1040 2.1005
R7303 VSS.n1047 VSS.n1046 2.1005
R7304 VSS.n1016 VSS.n1015 2.1005
R7305 VSS.n1022 VSS.n1021 2.1005
R7306 VSS.n10216 VSS.n10215 2.1005
R7307 VSS.n10210 VSS.n10209 2.1005
R7308 VSS.n317 VSS.n316 2.1005
R7309 VSS.n10222 VSS.n10221 2.1005
R7310 VSS.n1004 VSS.n1003 2.1005
R7311 VSS.n1010 VSS.n1009 2.1005
R7312 VSS.n983 VSS.n982 2.1005
R7313 VSS.n989 VSS.n988 2.1005
R7314 VSS.n305 VSS.n304 2.1005
R7315 VSS.n311 VSS.n310 2.1005
R7316 VSS.n10276 VSS.n10275 2.1005
R7317 VSS.n10270 VSS.n10269 2.1005
R7318 VSS.n967 VSS.n966 2.1005
R7319 VSS.n973 VSS.n972 2.1005
R7320 VSS.n10577 VSS.n10576 2.1005
R7321 VSS.n10580 VSS.n10579 2.1005
R7322 VSS.n10584 VSS.n10583 2.1005
R7323 VSS.n10675 VSS.n10674 2.1005
R7324 VSS.n10672 VSS.n10671 2.1005
R7325 VSS.n10668 VSS.n10667 2.1005
R7326 VSS.n10356 VSS.n10339 2.1005
R7327 VSS.n10360 VSS.n10359 2.1005
R7328 VSS.n10363 VSS.n10362 2.1005
R7329 VSS.n10419 VSS.n10418 2.1005
R7330 VSS.n10422 VSS.n10421 2.1005
R7331 VSS.n10426 VSS.n10425 2.1005
R7332 VSS.n10430 VSS.n10429 2.1005
R7333 VSS.n10434 VSS.n10433 2.1005
R7334 VSS.n10437 VSS.n10436 2.1005
R7335 VSS.n10588 VSS.n10587 2.1005
R7336 VSS.n10550 VSS.n10549 2.1005
R7337 VSS.n10541 VSS.n10488 2.1005
R7338 VSS.n10523 VSS.n10522 2.1005
R7339 VSS.n10514 VSS.n10509 2.1005
R7340 VSS.n10654 VSS.n10653 2.1005
R7341 VSS.n10548 VSS.n10547 2.1005
R7342 VSS.n10546 VSS.n10545 2.1005
R7343 VSS.n10501 VSS.n10492 2.1005
R7344 VSS.n10527 VSS.n10526 2.1005
R7345 VSS.n10521 VSS.n10520 2.1005
R7346 VSS.n10519 VSS.n10518 2.1005
R7347 VSS.n10652 VSS.n10651 2.1005
R7348 VSS.n10647 VSS.n10646 2.1005
R7349 VSS.n10644 VSS.n10643 2.1005
R7350 VSS.n10919 VSS.n10918 2.1005
R7351 VSS.n10988 VSS.n10987 2.1005
R7352 VSS.n10997 VSS.n10996 2.1005
R7353 VSS.n11357 VSS.n11356 2.1005
R7354 VSS.n11351 VSS.n11350 2.1005
R7355 VSS.n11344 VSS.n11343 2.1005
R7356 VSS.n9451 VSS.n9450 2.1005
R7357 VSS.n9457 VSS.n9456 2.1005
R7358 VSS.n9432 VSS.n9431 2.1005
R7359 VSS.n9472 VSS.n9471 2.1005
R7360 VSS.n819 VSS.n818 2.1005
R7361 VSS.n675 VSS.n674 2.1005
R7362 VSS.n9856 VSS.n9855 2.1005
R7363 VSS.n9876 VSS.n9875 2.1005
R7364 VSS.n11415 VSS.n11414 2.1005
R7365 VSS.n11448 VSS.n11447 2.1005
R7366 VSS.n9515 VSS.n9514 2.1005
R7367 VSS.n1251 VSS.n1250 2.1005
R7368 VSS.n9899 VSS.n9898 2.1005
R7369 VSS.n9912 VSS.n9911 2.1005
R7370 VSS.n9922 VSS.n9921 2.1005
R7371 VSS.n1372 VSS.n1347 2.1005
R7372 VSS.n1366 VSS.n1350 2.1005
R7373 VSS.n1360 VSS.n1352 2.1005
R7374 VSS.n9631 VSS.n9630 2.1005
R7375 VSS.n9763 VSS.n799 2.1005
R7376 VSS.n9757 VSS.n9637 2.1005
R7377 VSS.n9747 VSS.n9664 2.1005
R7378 VSS.n9741 VSS.n9667 2.1005
R7379 VSS.n9735 VSS.n9669 2.1005
R7380 VSS.n9725 VSS.n9720 2.1005
R7381 VSS.n10029 VSS.n570 2.1005
R7382 VSS.n10022 VSS.n575 2.1005
R7383 VSS.n10010 VSS.n9937 2.1005
R7384 VSS.n10004 VSS.n9939 2.1005
R7385 VSS.n9998 VSS.n9941 2.1005
R7386 VSS.n9988 VSS.n9969 2.1005
R7387 VSS.n9982 VSS.n9971 2.1005
R7388 VSS.n9976 VSS.n9973 2.1005
R7389 VSS.n1373 VSS.n1372 2.1005
R7390 VSS.n1367 VSS.n1366 2.1005
R7391 VSS.n1361 VSS.n1360 2.1005
R7392 VSS.n9632 VSS.n9631 2.1005
R7393 VSS.n9763 VSS.n9762 2.1005
R7394 VSS.n9758 VSS.n9757 2.1005
R7395 VSS.n9748 VSS.n9747 2.1005
R7396 VSS.n9742 VSS.n9741 2.1005
R7397 VSS.n9736 VSS.n9735 2.1005
R7398 VSS.n9726 VSS.n9725 2.1005
R7399 VSS.n10029 VSS.n10028 2.1005
R7400 VSS.n10023 VSS.n10022 2.1005
R7401 VSS.n10011 VSS.n10010 2.1005
R7402 VSS.n10005 VSS.n10004 2.1005
R7403 VSS.n9999 VSS.n9998 2.1005
R7404 VSS.n9989 VSS.n9988 2.1005
R7405 VSS.n9983 VSS.n9982 2.1005
R7406 VSS.n9977 VSS.n9976 2.1005
R7407 VSS.n9614 VSS.n9613 2.1005
R7408 VSS.n1310 VSS.n1309 2.1005
R7409 VSS.n10114 VSS.n10113 2.1005
R7410 VSS.n10109 VSS.n10108 2.1005
R7411 VSS.n10094 VSS.n10093 2.1005
R7412 VSS.n10088 VSS.n10087 2.1005
R7413 VSS.n10082 VSS.n10081 2.1005
R7414 VSS.n525 VSS.n524 2.1005
R7415 VSS.n10063 VSS.n10062 2.1005
R7416 VSS.n10056 VSS.n10055 2.1005
R7417 VSS.n10041 VSS.n10040 2.1005
R7418 VSS.n10871 VSS.n235 2.1005
R7419 VSS.n10888 VSS.n10887 2.1005
R7420 VSS.n11133 VSS.n202 2.1005
R7421 VSS.n11130 VSS.n11129 2.1005
R7422 VSS.n11124 VSS.n11123 2.1005
R7423 VSS.n11109 VSS.n11108 2.1005
R7424 VSS.n11103 VSS.n11102 2.1005
R7425 VSS.n11097 VSS.n11096 2.1005
R7426 VSS.n1315 VSS.n1314 2.1005
R7427 VSS.n1306 VSS.n1305 2.1005
R7428 VSS.n445 VSS.n444 2.1005
R7429 VSS.n10106 VSS.n10105 2.1005
R7430 VSS.n10101 VSS.n10100 2.1005
R7431 VSS.n10092 VSS.n10091 2.1005
R7432 VSS.n10086 VSS.n10085 2.1005
R7433 VSS.n10078 VSS.n10077 2.1005
R7434 VSS.n10073 VSS.n10072 2.1005
R7435 VSS.n521 VSS.n520 2.1005
R7436 VSS.n532 VSS.n513 2.1005
R7437 VSS.n10058 VSS.n10057 2.1005
R7438 VSS.n10052 VSS.n10051 2.1005
R7439 VSS.n10044 VSS.n10043 2.1005
R7440 VSS.n10037 VSS.n10036 2.1005
R7441 VSS.n10892 VSS.n10891 2.1005
R7442 VSS.n10881 VSS.n10878 2.1005
R7443 VSS.n11148 VSS.n11147 2.1005
R7444 VSS.n11136 VSS.n11135 2.1005
R7445 VSS.n11127 VSS.n11126 2.1005
R7446 VSS.n11121 VSS.n11120 2.1005
R7447 VSS.n11116 VSS.n11115 2.1005
R7448 VSS.n11107 VSS.n11106 2.1005
R7449 VSS.n11101 VSS.n11100 2.1005
R7450 VSS.n11095 VSS.n11094 2.1005
R7451 VSS.n11464 VSS.n11463 2.1005
R7452 VSS.n11323 VSS.n11322 2.1005
R7453 VSS.n11373 VSS.n11372 2.1005
R7454 VSS.n11380 VSS.n11379 2.1005
R7455 VSS.n10951 VSS.n10950 2.1005
R7456 VSS.n11367 VSS.n11366 2.1005
R7457 VSS.n10941 VSS.n10940 2.1005
R7458 VSS.n10978 VSS.n10977 2.1005
R7459 VSS.n1167 VSS.n1166 2.1005
R7460 VSS.n10935 VSS.n10934 2.1005
R7461 VSS.n1213 VSS.n1212 2.1005
R7462 VSS.n1203 VSS.n1202 2.1005
R7463 VSS.n9539 VSS.n9538 2.1005
R7464 VSS.n9546 VSS.n9545 2.1005
R7465 VSS.n1474 VSS.n1473 2.1005
R7466 VSS.n1465 VSS.n1464 2.1005
R7467 VSS.n1460 VSS.n1459 2.1005
R7468 VSS.n1448 VSS.n1447 2.1005
R7469 VSS.n9596 VSS.n828 2.1005
R7470 VSS.n9592 VSS.n9591 2.1005
R7471 VSS.n9778 VSS.n9777 2.1005
R7472 VSS.n9789 VSS.n9788 2.1005
R7473 VSS.n9795 VSS.n9794 2.1005
R7474 VSS.n9805 VSS.n9804 2.1005
R7475 VSS.n9815 VSS.n9814 2.1005
R7476 VSS.n9828 VSS.n9827 2.1005
R7477 VSS.n9839 VSS.n9838 2.1005
R7478 VSS.n760 VSS.n759 2.1005
R7479 VSS.n753 VSS.n752 2.1005
R7480 VSS.n741 VSS.n727 2.1005
R7481 VSS.n738 VSS.n737 2.1005
R7482 VSS.n11160 VSS.n11159 2.1005
R7483 VSS.n11169 VSS.n11168 2.1005
R7484 VSS.n11273 VSS.n11272 2.1005
R7485 VSS.n11267 VSS.n11266 2.1005
R7486 VSS.n11260 VSS.n11259 2.1005
R7487 VSS.n11251 VSS.n11250 2.1005
R7488 VSS.n11245 VSS.n11244 2.1005
R7489 VSS.n11239 VSS.n11238 2.1005
R7490 VSS.n1469 VSS.n1468 2.1005
R7491 VSS.n1457 VSS.n1456 2.1005
R7492 VSS.n1451 VSS.n1450 2.1005
R7493 VSS.n9594 VSS.n9593 2.1005
R7494 VSS.n9773 VSS.n795 2.1005
R7495 VSS.n9786 VSS.n9785 2.1005
R7496 VSS.n9809 VSS.n9808 2.1005
R7497 VSS.n9820 VSS.n9819 2.1005
R7498 VSS.n9832 VSS.n9831 2.1005
R7499 VSS.n757 VSS.n756 2.1005
R7500 VSS.n749 VSS.n748 2.1005
R7501 VSS.n744 VSS.n743 2.1005
R7502 VSS.n11166 VSS.n11165 2.1005
R7503 VSS.n11276 VSS.n11275 2.1005
R7504 VSS.n11270 VSS.n11269 2.1005
R7505 VSS.n11253 VSS.n11252 2.1005
R7506 VSS.n11247 VSS.n11246 2.1005
R7507 VSS.n11241 VSS.n11240 2.1005
R7508 VSS.n1401 VSS.n1400 2.1005
R7509 VSS.n9533 VSS.n9532 2.1005
R7510 VSS.n1493 VSS.n1492 2.1005
R7511 VSS.n9418 VSS.n9417 2.1005
R7512 VSS.n9379 VSS.n9378 2.1005
R7513 VSS.n9386 VSS.n9385 2.1005
R7514 VSS.n9319 VSS.n9318 2.1005
R7515 VSS.n9342 VSS.n9341 2.1005
R7516 VSS.n9267 VSS.n9266 2.1005
R7517 VSS.n9353 VSS.n9352 2.1005
R7518 VSS.n9261 VSS.n9260 2.1005
R7519 VSS.n9295 VSS.n9294 2.1005
R7520 VSS.n9216 VSS.n9215 2.1005
R7521 VSS.n9313 VSS.n9312 2.1005
R7522 VSS.n9210 VSS.n9209 2.1005
R7523 VSS.n9244 VSS.n9243 2.1005
R7524 VSS.n9145 VSS.n9144 2.1005
R7525 VSS.n9255 VSS.n9254 2.1005
R7526 VSS.n9135 VSS.n9134 2.1005
R7527 VSS.n9173 VSS.n9172 2.1005
R7528 VSS.n1551 VSS.n1550 2.1005
R7529 VSS.n1545 VSS.n1544 2.1005
R7530 VSS.n9060 VSS.n9059 2.1005
R7531 VSS.n9204 VSS.n9203 2.1005
R7532 VSS.n11392 VSS.n59 2.08328
R7533 VSS.n11390 VSS.n61 2.08259
R7534 VSS.t671 VSS.t255 2.07259
R7535 VSS.t478 VSS.t261 2.07259
R7536 VSS.n10499 VSS.n128 1.97855
R7537 VSS.n8953 VSS.n8952 1.87288
R7538 VSS.n8953 VSS.n253 1.8724
R7539 VSS.n11318 VSS.n11317 1.8392
R7540 VSS.n10633 VSS.n10632 1.7274
R7541 VSS.n9198 VSS.n9197 1.69669
R7542 VSS.n9334 VSS.n9333 1.69669
R7543 VSS.n172 VSS.n171 1.69669
R7544 VSS.n9580 VSS.n9579 1.69669
R7545 VSS.n200 VSS.n199 1.69669
R7546 VSS.n481 VSS.n477 1.69669
R7547 VSS.n9031 VSS.n9030 1.69669
R7548 VSS.n271 VSS.n270 1.69669
R7549 VSS.n343 VSS.n342 1.69669
R7550 VSS.n415 VSS.n414 1.69669
R7551 VSS.n10735 VSS.t3566 1.6805
R7552 VSS.n10790 VSS.t818 1.6805
R7553 VSS.n10792 VSS.t2465 1.6805
R7554 VSS.n10811 VSS.t1192 1.6805
R7555 VSS.n10820 VSS.t3012 1.6805
R7556 VSS.n10701 VSS.t1756 1.6805
R7557 VSS.n10708 VSS.t3524 1.6805
R7558 VSS.n10709 VSS.t764 1.6805
R7559 VSS.n10710 VSS.t2433 1.6805
R7560 VSS.n10711 VSS.t1131 1.6805
R7561 VSS.n10712 VSS.t2958 1.6805
R7562 VSS.n10713 VSS.t1674 1.6805
R7563 VSS.n127 VSS.t3418 1.6805
R7564 VSS.n14 VSS.t3234 1.6805
R7565 VSS.n15 VSS.t2451 1.6805
R7566 VSS.n16 VSS.t2590 1.6805
R7567 VSS.n17 VSS.t1828 1.6805
R7568 VSS.n11294 VSS.t994 1.6805
R7569 VSS.n24 VSS.t1153 1.6805
R7570 VSS.n25 VSS.t3436 1.6805
R7571 VSS.n26 VSS.t2694 1.6805
R7572 VSS.n27 VSS.t2986 1.6805
R7573 VSS.n28 VSS.t915 1.6805
R7574 VSS.n38 VSS.t1540 1.6805
R7575 VSS.n39 VSS.t2520 1.6805
R7576 VSS.n40 VSS.t1764 1.6805
R7577 VSS.n41 VSS.t923 1.6805
R7578 VSS.n42 VSS.t1073 1.6805
R7579 VSS.n133 VSS.t3356 1.6805
R7580 VSS.n49 VSS.t2766 1.6805
R7581 VSS.n50 VSS.t1980 1.6805
R7582 VSS.n51 VSS.t1400 1.6805
R7583 VSS.n52 VSS.t482 1.6805
R7584 VSS.n53 VSS.t1690 1.6805
R7585 VSS.n10641 VSS.t2399 1.6805
R7586 VSS.n10639 VSS.t3632 1.6805
R7587 VSS.n10497 VSS.t3120 1.6805
R7588 VSS.n10494 VSS.t782 1.6805
R7589 VSS.n10605 VSS.t510 1.6805
R7590 VSS.n10608 VSS.t2988 1.6805
R7591 VSS.n10440 VSS.t1471 1.6805
R7592 VSS.n10497 VSS.t1962 1.6805
R7593 VSS.n10494 VSS.t2752 1.6805
R7594 VSS.n10605 VSS.t2534 1.6805
R7595 VSS.n10608 VSS.t1834 1.6805
R7596 VSS.n10440 VSS.t3346 1.6805
R7597 VSS.n10476 VSS.t3244 1.6805
R7598 VSS.n10478 VSS.t3076 1.6805
R7599 VSS.n10481 VSS.t1696 1.6805
R7600 VSS.n10596 VSS.t2906 1.6805
R7601 VSS.n10593 VSS.t1616 1.6805
R7602 VSS.n10453 VSS.t1021 1.6805
R7603 VSS.n10451 VSS.t804 1.6805
R7604 VSS.n10345 VSS.t2540 1.6805
R7605 VSS.n10659 VSS.t623 1.6805
R7606 VSS.n10656 VSS.t2453 1.6805
R7607 VSS.n10573 VSS.t1956 1.6805
R7608 VSS.n10560 VSS.t3174 1.6805
R7609 VSS.n10290 VSS.t851 1.6805
R7610 VSS.n10693 VSS.t597 1.6805
R7611 VSS.n10690 VSS.t3062 1.6805
R7612 VSS.n10688 VSS.t1531 1.6805
R7613 VSS.n1271 VSS.t1988 1.6805
R7614 VSS.n1270 VSS.t1190 1.6805
R7615 VSS.n1269 VSS.t1348 1.6805
R7616 VSS.n1268 VSS.t3628 1.6805
R7617 VSS.n1331 VSS.t2860 1.6805
R7618 VSS.n1334 VSS.t2053 1.6805
R7619 VSS.n1335 VSS.t2203 1.6805
R7620 VSS.n1339 VSS.t1440 1.6805
R7621 VSS.n1342 VSS.t746 1.6805
R7622 VSS.n9494 VSS.t1797 1.6805
R7623 VSS.n9490 VSS.t2187 1.6805
R7624 VSS.n9487 VSS.t3232 1.6805
R7625 VSS.n9506 VSS.t1694 1.6805
R7626 VSS.n9503 VSS.t2552 1.6805
R7627 VSS.n9500 VSS.t1740 1.6805
R7628 VSS.n1345 VSS.t485 1.6805
R7629 VSS.n1375 VSS.t3000 1.6805
R7630 VSS.n9474 VSS.t1550 1.6805
R7631 VSS.n9446 VSS.t2095 1.6805
R7632 VSS.n9424 VSS.t2998 1.6805
R7633 VSS.n9425 VSS.t2153 1.6805
R7634 VSS.n9426 VSS.t3340 1.6805
R7635 VSS.n9427 VSS.t2706 1.6805
R7636 VSS.n9428 VSS.t1245 1.6805
R7637 VSS.n806 VSS.t1760 1.6805
R7638 VSS.n807 VSS.t1880 1.6805
R7639 VSS.n808 VSS.t1067 1.6805
R7640 VSS.n809 VSS.t3354 1.6805
R7641 VSS.n1233 VSS.t3520 1.6805
R7642 VSS.n823 VSS.t2902 1.6805
R7643 VSS.n824 VSS.t2111 1.6805
R7644 VSS.n825 VSS.t1521 1.6805
R7645 VSS.n826 VSS.t664 1.6805
R7646 VSS.n806 VSS.t543 1.6805
R7647 VSS.n807 VSS.t724 1.6805
R7648 VSS.n808 VSS.t3084 1.6805
R7649 VSS.n809 VSS.t2265 1.6805
R7650 VSS.n1233 VSS.t2383 1.6805
R7651 VSS.n823 VSS.t1790 1.6805
R7652 VSS.n824 VSS.t964 1.6805
R7653 VSS.n825 VSS.t3440 1.6805
R7654 VSS.n826 VSS.t2700 1.6805
R7655 VSS.n9639 VSS.t1738 1.6805
R7656 VSS.n9640 VSS.t1864 1.6805
R7657 VSS.n9641 VSS.t1050 1.6805
R7658 VSS.n9642 VSS.t3332 1.6805
R7659 VSS.n647 VSS.t3496 1.6805
R7660 VSS.n777 VSS.t2890 1.6805
R7661 VSS.n776 VSS.t2087 1.6805
R7662 VSS.n775 VSS.t1509 1.6805
R7663 VSS.n774 VSS.t636 1.6805
R7664 VSS.n9639 VSS.t512 1.6805
R7665 VSS.n9640 VSS.t702 1.6805
R7666 VSS.n9641 VSS.t3058 1.6805
R7667 VSS.n9642 VSS.t2255 1.6805
R7668 VSS.n647 VSS.t2369 1.6805
R7669 VSS.n777 VSS.t1776 1.6805
R7670 VSS.n776 VSS.t935 1.6805
R7671 VSS.n775 VSS.t3416 1.6805
R7672 VSS.n774 VSS.t2662 1.6805
R7673 VSS.n9672 VSS.t1912 1.6805
R7674 VSS.n9675 VSS.t1094 1.6805
R7675 VSS.n9678 VSS.t3376 1.6805
R7676 VSS.n9681 VSS.t3546 1.6805
R7677 VSS.n1175 VSS.t2780 1.6805
R7678 VSS.n681 VSS.t2145 1.6805
R7679 VSS.n684 VSS.t1373 1.6805
R7680 VSS.n687 VSS.t714 1.6805
R7681 VSS.n690 VSS.t3078 1.6805
R7682 VSS.n9673 VSS.t824 1.6805
R7683 VSS.n9676 VSS.t966 1.6805
R7684 VSS.n9679 VSS.t3278 1.6805
R7685 VSS.n9682 VSS.t2490 1.6805
R7686 VSS.n1174 VSS.t2636 1.6805
R7687 VSS.n682 VSS.t2004 1.6805
R7688 VSS.n685 VSS.t1242 1.6805
R7689 VSS.n688 VSS.t541 1.6805
R7690 VSS.n691 VSS.t2940 1.6805
R7691 VSS.n660 VSS.t3468 1.6805
R7692 VSS.n659 VSS.t2712 1.6805
R7693 VSS.n658 VSS.t1928 1.6805
R7694 VSS.n657 VSS.t2043 1.6805
R7695 VSS.n672 VSS.t1269 1.6805
R7696 VSS.n9860 VSS.t562 1.6805
R7697 VSS.n9861 VSS.t2948 1.6805
R7698 VSS.n9862 VSS.t2315 1.6805
R7699 VSS.n9863 VSS.t1558 1.6805
R7700 VSS.n660 VSS.t2349 1.6805
R7701 VSS.n659 VSS.t1599 1.6805
R7702 VSS.n658 VSS.t753 1.6805
R7703 VSS.n657 VSS.t894 1.6805
R7704 VSS.n672 VSS.t3218 1.6805
R7705 VSS.n9860 VSS.t2588 1.6805
R7706 VSS.n9861 VSS.t1826 1.6805
R7707 VSS.n9862 VSS.t1206 1.6805
R7708 VSS.n9863 VSS.t3498 1.6805
R7709 VSS.n9955 VSS.t2409 1.6805
R7710 VSS.n9956 VSS.t1652 1.6805
R7711 VSS.n9957 VSS.t820 1.6805
R7712 VSS.n9958 VSS.t954 1.6805
R7713 VSS.n142 VSS.t3268 1.6805
R7714 VSS.n11186 VSS.t2652 1.6805
R7715 VSS.n11185 VSS.t1876 1.6805
R7716 VSS.n11184 VSS.t1267 1.6805
R7717 VSS.n11183 VSS.t3556 1.6805
R7718 VSS.n9955 VSS.t1309 1.6805
R7719 VSS.n9956 VSS.t3586 1.6805
R7720 VSS.n9957 VSS.t2830 1.6805
R7721 VSS.n9958 VSS.t2962 1.6805
R7722 VSS.n142 VSS.t2173 1.6805
R7723 VSS.n11186 VSS.t1548 1.6805
R7724 VSS.n11185 VSS.t717 1.6805
R7725 VSS.n11184 VSS.t3216 1.6805
R7726 VSS.n11183 VSS.t2435 1.6805
R7727 VSS.n1259 VSS.t2528 1.6805
R7728 VSS.n1258 VSS.t1772 1.6805
R7729 VSS.n1257 VSS.t1890 1.6805
R7730 VSS.n1256 VSS.t1075 1.6805
R7731 VSS.n1236 VSS.t3366 1.6805
R7732 VSS.n1237 VSS.t2612 1.6805
R7733 VSS.n1238 VSS.t2748 1.6805
R7734 VSS.n1239 VSS.t1966 1.6805
R7735 VSS.n1240 VSS.t1354 1.6805
R7736 VSS.n1259 VSS.t1414 1.6805
R7737 VSS.n1258 VSS.t507 1.6805
R7738 VSS.n1257 VSS.t697 1.6805
R7739 VSS.n1256 VSS.t3054 1.6805
R7740 VSS.n1236 VSS.t2253 1.6805
R7741 VSS.n1237 VSS.t1487 1.6805
R7742 VSS.n1238 VSS.t1628 1.6805
R7743 VSS.n1239 VSS.t778 1.6805
R7744 VSS.n1240 VSS.t3254 1.6805
R7745 VSS.n633 VSS.t2363 1.6805
R7746 VSS.n632 VSS.t1603 1.6805
R7747 VSS.n631 VSS.t1728 1.6805
R7748 VSS.n630 VSS.t903 1.6805
R7749 VSS.n643 VSS.t3222 1.6805
R7750 VSS.n9653 VSS.t2441 1.6805
R7751 VSS.n9652 VSS.t2570 1.6805
R7752 VSS.n9651 VSS.t1809 1.6805
R7753 VSS.n9650 VSS.t1160 1.6805
R7754 VSS.n633 VSS.t1220 1.6805
R7755 VSS.n632 VSS.t3516 1.6805
R7756 VSS.n631 VSS.t468 1.6805
R7757 VSS.n630 VSS.t2882 1.6805
R7758 VSS.n643 VSS.t2077 1.6805
R7759 VSS.n9653 VSS.t1311 1.6805
R7760 VSS.n9652 VSS.t1454 1.6805
R7761 VSS.n9651 VSS.t579 1.6805
R7762 VSS.n9650 VSS.t3118 1.6805
R7763 VSS.n603 VSS.t1660 1.6805
R7764 VSS.n608 VSS.t822 1.6805
R7765 VSS.n613 VSS.t960 1.6805
R7766 VSS.n618 VSS.t3274 1.6805
R7767 VSS.n624 VSS.t2480 1.6805
R7768 VSS.n9700 VSS.t2628 1.6805
R7769 VSS.n9705 VSS.t1860 1.6805
R7770 VSS.n9710 VSS.t1046 1.6805
R7771 VSS.n9715 VSS.t1375 1.6805
R7772 VSS.n602 VSS.t1501 1.6805
R7773 VSS.n607 VSS.t629 1.6805
R7774 VSS.n612 VSS.t788 1.6805
R7775 VSS.n617 VSS.t3138 1.6805
R7776 VSS.n625 VSS.t2331 1.6805
R7777 VSS.n9699 VSS.t1580 1.6805
R7778 VSS.n9704 VSS.t1706 1.6805
R7779 VSS.n9709 VSS.t882 1.6805
R7780 VSS.n9714 VSS.t3324 1.6805
R7781 VSS.n589 VSS.t2199 1.6805
R7782 VSS.n588 VSS.t1438 1.6805
R7783 VSS.n587 VSS.t1560 1.6805
R7784 VSS.n586 VSS.t726 1.6805
R7785 VSS.n9915 VSS.t3088 1.6805
R7786 VSS.n582 VSS.t3184 1.6805
R7787 VSS.n581 VSS.t2389 1.6805
R7788 VSS.n580 VSS.t1638 1.6805
R7789 VSS.n579 VSS.t1924 1.6805
R7790 VSS.n589 VSS.t1011 1.6805
R7791 VSS.n588 VSS.t3306 1.6805
R7792 VSS.n587 VSS.t3462 1.6805
R7793 VSS.n586 VSS.t2708 1.6805
R7794 VSS.n9915 VSS.t1920 1.6805
R7795 VSS.n582 VSS.t2030 1.6805
R7796 VSS.n581 VSS.t1261 1.6805
R7797 VSS.n580 VSS.t3550 1.6805
R7798 VSS.n579 VSS.t731 1.6805
R7799 VSS.n11039 VSS.t2816 1.6805
R7800 VSS.n11040 VSS.t2008 1.6805
R7801 VSS.n11041 VSS.t2157 1.6805
R7802 VSS.n11042 VSS.t1381 1.6805
R7803 VSS.n11283 VSS.t473 1.6805
R7804 VSS.n9946 VSS.t662 1.6805
R7805 VSS.n9945 VSS.t3032 1.6805
R7806 VSS.n9944 VSS.t2221 1.6805
R7807 VSS.n9943 VSS.t2506 1.6805
R7808 VSS.n11039 VSS.t1668 1.6805
R7809 VSS.n11040 VSS.t830 1.6805
R7810 VSS.n11041 VSS.t970 1.6805
R7811 VSS.n11042 VSS.t3282 1.6805
R7812 VSS.n11283 VSS.t2502 1.6805
R7813 VSS.n9946 VSS.t2648 1.6805
R7814 VSS.n9945 VSS.t1872 1.6805
R7815 VSS.n9944 VSS.t1058 1.6805
R7816 VSS.n9943 VSS.t1394 1.6805
R7817 VSS.n9477 VSS.t3350 1.6805
R7818 VSS.n9478 VSS.t2584 1.6805
R7819 VSS.n9479 VSS.t1817 1.6805
R7820 VSS.n1385 VSS.t1946 1.6805
R7821 VSS.n1407 VSS.t1328 1.6805
R7822 VSS.n1406 VSS.t3608 1.6805
R7823 VSS.n1405 VSS.t3024 1.6805
R7824 VSS.n1404 VSS.t2215 1.6805
R7825 VSS.n10687 VSS.n10686 1.67828
R7826 VSS.n10678 VSS.n10677 1.67828
R7827 VSS.n10311 VSS.n10292 1.67718
R7828 VSS.n10982 VSS.n181 1.67411
R7829 VSS.n11318 VSS.n11316 1.65519
R7830 VSS.n10632 VSS.n10631 1.60175
R7831 VSS.n10751 VSS.n10750 1.5755
R7832 VSS.n10817 VSS.n10816 1.5755
R7833 VSS.n10780 VSS.n10779 1.5755
R7834 VSS.n10786 VSS.n10785 1.5755
R7835 VSS.n10038 VSS.n238 1.53593
R7836 VSS.n560 VSS.n239 1.53593
R7837 VSS.n11320 VSS.n116 1.53593
R7838 VSS.n10537 VSS.n10536 1.53593
R7839 VSS.n10529 VSS.n10528 1.53593
R7840 VSS.n10613 VSS.n10612 1.5005
R7841 VSS.n10411 VSS.n10410 1.5005
R7842 VSS.n10679 VSS.n10678 1.5005
R7843 VSS.n10334 VSS.n10333 1.5005
R7844 VSS.n10536 VSS.n10535 1.5005
R7845 VSS.n10533 VSS.n10493 1.5005
R7846 VSS.n10530 VSS.n10529 1.5005
R7847 VSS.n558 VSS.n239 1.5005
R7848 VSS.n10869 VSS.n10868 1.5005
R7849 VSS.n238 VSS.n236 1.5005
R7850 VSS.n120 VSS.n117 1.5005
R7851 VSS.n11321 VSS.n11320 1.5005
R7852 VSS.n817 VSS.n650 1.47409
R7853 VSS.n822 VSS.n821 1.47409
R7854 VSS.n9883 VSS.n652 1.47409
R7855 VSS.n678 VSS.n677 1.47409
R7856 VSS.n9880 VSS.n656 1.47409
R7857 VSS.n9859 VSS.n9858 1.47409
R7858 VSS.n9878 VSS.n9877 1.47409
R7859 VSS.n9874 VSS.n9873 1.47409
R7860 VSS.n11413 VSS.n11412 1.47409
R7861 VSS.n11417 VSS.n11416 1.47409
R7862 VSS.n11446 VSS.n11445 1.47409
R7863 VSS.n11450 VSS.n11449 1.47409
R7864 VSS.n9517 VSS.n9516 1.47409
R7865 VSS.n9513 VSS.n9512 1.47409
R7866 VSS.n1249 VSS.n642 1.47409
R7867 VSS.n1254 VSS.n1253 1.47409
R7868 VSS.n9897 VSS.n9896 1.47409
R7869 VSS.n9902 VSS.n9901 1.47409
R7870 VSS.n9914 VSS.n9913 1.47409
R7871 VSS.n9910 VSS.n584 1.47409
R7872 VSS.n9920 VSS.n9919 1.47409
R7873 VSS.n9925 VSS.n9924 1.47409
R7874 VSS.n9612 VSS.n9611 1.47409
R7875 VSS.n9616 VSS.n9615 1.47409
R7876 VSS.n10405 VSS.n10404 1.46537
R7877 VSS.n10409 VSS.n10408 1.46537
R7878 VSS.n10403 VSS.n10402 1.46537
R7879 VSS.n10326 VSS.n10325 1.46537
R7880 VSS.n10330 VSS.n10329 1.46537
R7881 VSS.n10332 VSS.n10331 1.46537
R7882 VSS.n10321 VSS.n10320 1.46537
R7883 VSS.n10319 VSS.n10318 1.46537
R7884 VSS.n10315 VSS.n10314 1.46537
R7885 VSS.n10311 VSS.n10310 1.46537
R7886 VSS.n11316 VSS.n11314 1.37022
R7887 VSS.n10789 VSS.t3114 1.348
R7888 VSS.n10834 VSS.t3538 1.348
R7889 VSS.n10810 VSS.t843 1.348
R7890 VSS.n10812 VSS.t2770 1.348
R7891 VSS.n10775 VSS.t1462 1.348
R7892 VSS.n246 VSS.t1894 1.348
R7893 VSS.n10744 VSS.t2291 1.348
R7894 VSS.n10753 VSS.t1078 1.348
R7895 VSS.n9449 VSS.t3085 1.26547
R7896 VSS.n9423 VSS.t1793 1.26547
R7897 VSS.n9453 VSS.t2474 1.26547
R7898 VSS.n9455 VSS.t1236 1.26547
R7899 VSS.n9429 VSS.t2035 1.26547
R7900 VSS.n9430 VSS.t3513 1.26547
R7901 VSS.n9470 VSS.t3007 1.26547
R7902 VSS.n1378 VSS.t1401 1.26547
R7903 VSS.n129 VSS.t1428 1.26547
R7904 VSS.n10698 VSS.t2789 1.26547
R7905 VSS.n10734 VSS.t1800 1.26547
R7906 VSS.n10824 VSS.t3479 1.26547
R7907 VSS.n10824 VSS.t1709 1.26547
R7908 VSS.n10867 VSS.n10866 1.26528
R7909 VSS.n10802 VSS.n10801 1.265
R7910 VSS.n9204 VSS.t2726 1.2605
R7911 VSS.t627 VSS.n9204 1.2605
R7912 VSS.t2275 VSS.n9060 1.2605
R7913 VSS.n9060 VSS.t3304 1.2605
R7914 VSS.t1511 VSS.n1545 1.2605
R7915 VSS.n1545 VSS.t3510 1.2605
R7916 VSS.t1015 VSS.n1551 1.2605
R7917 VSS.n1551 VSS.t1774 1.2605
R7918 VSS.t2016 VSS.n9173 1.2605
R7919 VSS.n9173 VSS.t3102 1.2605
R7920 VSS.n9135 VSS.t1605 1.2605
R7921 VSS.t2634 VSS.n9135 1.2605
R7922 VSS.n9255 VSS.t2942 1.2605
R7923 VSS.t862 VSS.n9255 1.2605
R7924 VSS.t2397 VSS.n9145 1.2605
R7925 VSS.n9145 VSS.t1712 1.2605
R7926 VSS.t3620 VSS.n9244 1.2605
R7927 VSS.n9244 VSS.t1618 1.2605
R7928 VSS.n9210 VSS.t3126 1.2605
R7929 VSS.t2385 VSS.n9210 1.2605
R7930 VSS.n9313 VSS.t968 1.2605
R7931 VSS.t2041 VSS.n9313 1.2605
R7932 VSS.t2313 VSS.n9216 1.2605
R7933 VSS.n9216 VSS.t1630 1.2605
R7934 VSS.t3344 VSS.n9295 1.2605
R7935 VSS.n9295 VSS.t1369 1.2605
R7936 VSS.n9261 VSS.t1634 1.2605
R7937 VSS.t880 VSS.n9261 1.2605
R7938 VSS.n9353 VSS.t2137 1.2605
R7939 VSS.t2852 VSS.n9353 1.2605
R7940 VSS.t2401 VSS.n9267 1.2605
R7941 VSS.n9267 VSS.t1377 1.2605
R7942 VSS.t2848 VSS.n9342 1.2605
R7943 VSS.n9342 VSS.t3534 1.2605
R7944 VSS.n9319 VSS.t3132 1.2605
R7945 VSS.t2049 VSS.n9319 1.2605
R7946 VSS.n9386 VSS.t470 1.2605
R7947 VSS.t2598 VSS.n9386 1.2605
R7948 VSS.n9379 VSS.t3214 1.2605
R7949 VSS.t2181 VSS.n9379 1.2605
R7950 VSS.t2982 VSS.n9418 1.2605
R7951 VSS.n9418 VSS.t1910 1.2605
R7952 VSS.t2512 VSS.n1493 1.2605
R7953 VSS.n1493 VSS.t1489 1.2605
R7954 VSS.n9533 VSS.t2179 1.2605
R7955 VSS.t1090 VSS.n9533 1.2605
R7956 VSS.t621 VSS.n1401 1.2605
R7957 VSS.n1401 VSS.t1416 1.2605
R7958 VSS.t2026 VSS.n11241 1.2605
R7959 VSS.n11241 VSS.t952 1.2605
R7960 VSS.t2439 VSS.n11247 1.2605
R7961 VSS.n11247 VSS.t3152 1.2605
R7962 VSS.t3560 VSS.n11253 1.2605
R7963 VSS.n11253 VSS.t2872 1.2605
R7964 VSS.n11269 VSS.t1527 1.2605
R7965 VSS.n11269 VSS.t2546 1.2605
R7966 VSS.n11275 VSS.t1118 1.2605
R7967 VSS.n11275 VSS.t1932 1.2605
R7968 VSS.n11166 VSS.t1566 1.2605
R7969 VSS.t2257 VSS.n11166 1.2605
R7970 VSS.t3276 VSS.n744 1.2605
R7971 VSS.n744 VSS.t2225 1.2605
R7972 VSS.n748 VSS.t520 1.2605
R7973 VSS.n748 VSS.t2996 1.2605
R7974 VSS.n756 VSS.t3368 1.2605
R7975 VSS.n756 VSS.t988 1.2605
R7976 VSS.n9832 VSS.t3286 1.2605
R7977 VSS.t2251 VSS.n9832 1.2605
R7978 VSS.n9820 VSS.t548 1.2605
R7979 VSS.t1356 VSS.n9820 1.2605
R7980 VSS.n9809 VSS.t2812 1.2605
R7981 VSS.t2083 VSS.n9809 1.2605
R7982 VSS.n9786 VSS.t2788 1.2605
R7983 VSS.t711 VSS.n9786 1.2605
R7984 VSS.n9773 VSS.t1151 1.2605
R7985 VSS.t3182 VSS.n9773 1.2605
R7986 VSS.t2834 VSS.n9594 1.2605
R7987 VSS.n9594 VSS.t3582 1.2605
R7988 VSS.t2808 VSS.n1451 1.2605
R7989 VSS.n1451 VSS.t3490 1.2605
R7990 VSS.n1457 VSS.t1882 1.2605
R7991 VSS.t1164 VSS.n1457 1.2605
R7992 VSS.t1611 VSS.n1469 1.2605
R7993 VSS.n1469 VSS.t2281 1.2605
R7994 VSS.n11238 VSS.t802 1.2605
R7995 VSS.n11238 VSS.t3202 1.2605
R7996 VSS.n11244 VSS.t3438 1.2605
R7997 VSS.n11244 VSS.t1456 1.2605
R7998 VSS.n11250 VSS.t2964 1.2605
R7999 VSS.n11250 VSS.t1898 1.2605
R8000 VSS.t2149 VSS.n11260 1.2605
R8001 VSS.n11260 VSS.t3190 1.2605
R8002 VSS.n11266 VSS.t3448 1.2605
R8003 VSS.n11266 VSS.t2764 1.2605
R8004 VSS.n11272 VSS.t940 1.2605
R8005 VSS.n11272 VSS.t3308 1.2605
R8006 VSS.n11169 VSS.t592 1.2605
R8007 VSS.t3048 VSS.n11169 1.2605
R8008 VSS.n11160 VSS.t1251 1.2605
R8009 VSS.t2289 VSS.n11160 1.2605
R8010 VSS.t768 VSS.n738 1.2605
R8011 VSS.n738 VSS.t1868 1.2605
R8012 VSS.n741 VSS.t3158 1.2605
R8013 VSS.t2105 VSS.n741 1.2605
R8014 VSS.n752 VSS.t2034 1.2605
R8015 VSS.n752 VSS.t1352 1.2605
R8016 VSS.n759 VSS.t1607 1.2605
R8017 VSS.n759 VSS.t3596 1.2605
R8018 VSS.n9839 VSS.t1124 1.2605
R8019 VSS.t1862 VSS.n9839 1.2605
R8020 VSS.n9827 VSS.t1680 1.2605
R8021 VSS.n9827 VSS.t516 1.2605
R8022 VSS.n9814 VSS.t1054 1.2605
R8023 VSS.n9814 VSS.t2133 1.2605
R8024 VSS.n9804 VSS.t3382 1.2605
R8025 VSS.n9804 VSS.t2359 1.2605
R8026 VSS.n9794 VSS.t1944 1.2605
R8027 VSS.n9794 VSS.t3018 1.2605
R8028 VSS.n9789 VSS.t1210 1.2605
R8029 VSS.t3226 VSS.n9789 1.2605
R8030 VSS.n9778 VSS.t2002 1.2605
R8031 VSS.t2722 VSS.n9778 1.2605
R8032 VSS.n9591 VSS.t1503 1.2605
R8033 VSS.n9591 VSS.t2261 1.2605
R8034 VSS.n9596 VSS.t1007 1.2605
R8035 VSS.t1770 VSS.n9596 1.2605
R8036 VSS.t3358 VSS.n1448 1.2605
R8037 VSS.n1448 VSS.t2323 1.2605
R8038 VSS.t3588 VSS.n1460 1.2605
R8039 VSS.n1460 VSS.t1227 1.2605
R8040 VSS.n1464 VSS.t2880 1.2605
R8041 VSS.n1464 VSS.t1813 1.2605
R8042 VSS.t1412 VSS.n1474 1.2605
R8043 VSS.n1474 VSS.t2091 1.2605
R8044 VSS.n9546 VSS.t738 1.2605
R8045 VSS.t1572 VSS.n9546 1.2605
R8046 VSS.n9539 VSS.t3386 1.2605
R8047 VSS.t1017 VSS.n9539 1.2605
R8048 VSS.t2728 VSS.n1203 1.2605
R8049 VSS.n1203 VSS.t1682 1.2605
R8050 VSS.t1247 VSS.n1213 1.2605
R8051 VSS.n1213 VSS.t2287 1.2605
R8052 VSS.n10935 VSS.t847 1.2605
R8053 VSS.t2928 VSS.n10935 1.2605
R8054 VSS.t3526 VSS.n1167 1.2605
R8055 VSS.n1167 VSS.t1135 1.2605
R8056 VSS.t3624 VSS.n10978 1.2605
R8057 VSS.n10978 VSS.t1622 1.2605
R8058 VSS.n10941 VSS.t3178 1.2605
R8059 VSS.t1145 VSS.n10941 1.2605
R8060 VSS.n11367 VSS.t1464 1.2605
R8061 VSS.t2473 VSS.n11367 1.2605
R8062 VSS.t2778 VSS.n10951 1.2605
R8063 VSS.n10951 VSS.t2051 1.2605
R8064 VSS.n11380 VSS.t1902 1.2605
R8065 VSS.t2968 VSS.n11380 1.2605
R8066 VSS.n11373 VSS.t3210 1.2605
R8067 VSS.t2494 VSS.n11373 1.2605
R8068 VSS.n11323 VSS.t1974 1.2605
R8069 VSS.t2211 VSS.n11323 1.2605
R8070 VSS.t1493 VSS.n11464 1.2605
R8071 VSS.n11464 VSS.t1460 1.2605
R8072 VSS.n11094 VSS.t625 1.2605
R8073 VSS.n11094 VSS.t1714 1.2605
R8074 VSS.n11100 VSS.t2914 1.2605
R8075 VSS.n11100 VSS.t2886 1.2605
R8076 VSS.n11106 VSS.t1044 1.2605
R8077 VSS.n11106 VSS.t1320 1.2605
R8078 VSS.t2482 VSS.n11116 1.2605
R8079 VSS.n11116 VSS.t2457 1.2605
R8080 VSS.t1746 VSS.n11121 1.2605
R8081 VSS.n11121 VSS.t2740 1.2605
R8082 VSS.t1672 VSS.n11127 1.2605
R8083 VSS.n11127 VSS.t2668 1.2605
R8084 VSS.t1299 VSS.n11136 1.2605
R8085 VSS.n11136 VSS.t2303 1.2605
R8086 VSS.t1235 VSS.n11148 1.2605
R8087 VSS.n11148 VSS.t1184 1.2605
R8088 VSS.n10881 VSS.t1513 1.2605
R8089 VSS.t1485 VSS.n10881 1.2605
R8090 VSS.t3430 VSS.n10892 1.2605
R8091 VSS.n10892 VSS.t532 1.2605
R8092 VSS.n10036 VSS.t3406 1.2605
R8093 VSS.n10036 VSS.t1398 1.2605
R8094 VSS.n10043 VSS.t2556 1.2605
R8095 VSS.n10043 VSS.t2822 1.2605
R8096 VSS.t2850 VSS.n10052 1.2605
R8097 VSS.n10052 VSS.t2020 1.2605
R8098 VSS.t2057 VSS.n10058 1.2605
R8099 VSS.n10058 VSS.t2295 1.2605
R8100 VSS.n532 VSS.t2802 1.2605
R8101 VSS.t2754 VSS.n532 1.2605
R8102 VSS.n520 VSS.t1684 1.2605
R8103 VSS.n520 VSS.t1916 1.2605
R8104 VSS.t1109 VSS.n10073 1.2605
R8105 VSS.n10073 VSS.t1080 1.2605
R8106 VSS.n10077 VSS.t3112 1.2605
R8107 VSS.n10077 VSS.t3302 1.2605
R8108 VSS.n10085 VSS.t1143 1.2605
R8109 VSS.n10085 VSS.t3398 1.2605
R8110 VSS.n10091 VSS.t2672 1.2605
R8111 VSS.n10091 VSS.t2548 1.2605
R8112 VSS.t2950 VSS.n10101 1.2605
R8113 VSS.n10101 VSS.t2135 1.2605
R8114 VSS.t1830 VSS.n10106 1.2605
R8115 VSS.n10106 VSS.t2047 1.2605
R8116 VSS.n445 VSS.t2864 1.2605
R8117 VSS.t2032 VSS.n445 1.2605
R8118 VSS.n1305 VSS.t1748 1.2605
R8119 VSS.n1305 VSS.t1972 1.2605
R8120 VSS.n1314 VSS.t1186 1.2605
R8121 VSS.n1314 VSS.t3456 1.2605
R8122 VSS.t2478 VSS.n11097 1.2605
R8123 VSS.n11097 VSS.t2744 1.2605
R8124 VSS.t2445 VSS.n11103 1.2605
R8125 VSS.n11103 VSS.t1664 1.2605
R8126 VSS.t457 VSS.n11109 1.2605
R8127 VSS.n11109 VSS.t1592 1.2605
R8128 VSS.t3614 VSS.n11124 1.2605
R8129 VSS.n11124 VSS.t3574 1.2605
R8130 VSS.t2862 VSS.n11130 1.2605
R8131 VSS.n11130 VSS.t2738 1.2605
R8132 VSS.n11133 VSS.t2810 1.2605
R8133 VSS.t1996 VSS.n11133 1.2605
R8134 VSS.n10887 VSS.t899 1.2605
R8135 VSS.n10887 VSS.t1162 1.2605
R8136 VSS.n10871 VSS.t840 1.2605
R8137 VSS.t1900 VSS.n10871 1.2605
R8138 VSS.n10040 VSS.t766 1.2605
R8139 VSS.n10040 VSS.t3106 1.2605
R8140 VSS.n10055 VSS.t2361 1.2605
R8141 VSS.n10055 VSS.t2600 1.2605
R8142 VSS.n10062 VSS.t2311 1.2605
R8143 VSS.n10062 VSS.t1533 1.2605
R8144 VSS.n525 VSS.t1229 1.2605
R8145 VSS.t2229 VSS.n525 1.2605
R8146 VSS.t3470 VSS.n10082 1.2605
R8147 VSS.n10082 VSS.t3426 1.2605
R8148 VSS.t2351 VSS.n10088 1.2605
R8149 VSS.n10088 VSS.t2596 1.2605
R8150 VSS.t2660 VSS.n10094 1.2605
R8151 VSS.n10094 VSS.t2544 1.2605
R8152 VSS.t1848 VSS.n10109 1.2605
R8153 VSS.n10109 VSS.t1001 1.2605
R8154 VSS.n10113 VSS.t707 1.2605
R8155 VSS.n10113 VSS.t1778 1.2605
R8156 VSS.t599 VSS.n1310 1.2605
R8157 VSS.n1310 VSS.t2960 1.2605
R8158 VSS.t2403 VSS.n11344 1.2605
R8159 VSS.n11344 VSS.t2371 1.2605
R8160 VSS.t1658 VSS.n11351 1.2605
R8161 VSS.n11351 VSS.t2650 1.2605
R8162 VSS.t3420 VSS.n11357 1.2605
R8163 VSS.n11357 VSS.t3378 1.2605
R8164 VSS.t2678 VSS.n10997 1.2605
R8165 VSS.n10997 VSS.t514 1.2605
R8166 VSS.n10988 VSS.t2183 1.2605
R8167 VSS.t2147 VSS.n10988 1.2605
R8168 VSS.t2423 VSS.n10919 1.2605
R8169 VSS.n10919 VSS.t2391 1.2605
R8170 VSS.n10643 VSS.t2582 1.2605
R8171 VSS.n10643 VSS.t786 1.2605
R8172 VSS.t1648 VSS.n10647 1.2605
R8173 VSS.n10647 VSS.t2582 1.2605
R8174 VSS.t1069 VSS.n10652 1.2605
R8175 VSS.n10652 VSS.t2393 1.2605
R8176 VSS.t2844 VSS.n10519 1.2605
R8177 VSS.n10519 VSS.t656 1.2605
R8178 VSS.n10520 VSS.t2924 1.2605
R8179 VSS.n10520 VSS.t2844 1.2605
R8180 VSS.n10526 VSS.t1028 1.2605
R8181 VSS.n10526 VSS.t2283 1.2605
R8182 VSS.n10501 VSS.t3170 1.2605
R8183 VSS.t1028 VSS.n10501 1.2605
R8184 VSS.t2626 VSS.n10546 1.2605
R8185 VSS.n10546 VSS.t3590 1.2605
R8186 VSS.n10547 VSS.t1688 1.2605
R8187 VSS.n10547 VSS.t2626 1.2605
R8188 VSS.n10653 VSS.t1166 1.2605
R8189 VSS.n10653 VSS.t1069 1.2605
R8190 VSS.n10514 VSS.t566 1.2605
R8191 VSS.t873 VSS.n10514 1.2605
R8192 VSS.t2750 VSS.n10523 1.2605
R8193 VSS.n10523 VSS.t566 1.2605
R8194 VSS.n10541 VSS.t887 1.2605
R8195 VSS.t1888 VSS.n10541 1.2605
R8196 VSS.t3056 VSS.n10550 1.2605
R8197 VSS.n10550 VSS.t887 1.2605
R8198 VSS.n10588 VSS.t3258 1.2605
R8199 VSS.t1141 VSS.n10588 1.2605
R8200 VSS.n10437 VSS.t3554 1.2605
R8201 VSS.t1469 VSS.n10437 1.2605
R8202 VSS.n10433 VSS.t2576 1.2605
R8203 VSS.n10433 VSS.t3554 1.2605
R8204 VSS.n10430 VSS.t2846 1.2605
R8205 VSS.t658 VSS.n10430 1.2605
R8206 VSS.n10425 VSS.t2926 1.2605
R8207 VSS.n10425 VSS.t2846 1.2605
R8208 VSS.n10422 VSS.t2367 1.2605
R8209 VSS.t2285 VSS.n10422 1.2605
R8210 VSS.n10418 VSS.t1434 1.2605
R8211 VSS.n10418 VSS.t2367 1.2605
R8212 VSS.n10455 VSS.t3256 1.2605
R8213 VSS.n10455 VSS.t1139 1.2605
R8214 VSS.t3310 VSS.n10459 1.2605
R8215 VSS.n10459 VSS.t3256 1.2605
R8216 VSS.n10462 VSS.t1519 1.2605
R8217 VSS.n10462 VSS.t2732 1.2605
R8218 VSS.t3600 VSS.n10467 1.2605
R8219 VSS.n10467 VSS.t1519 1.2605
R8220 VSS.n10470 VSS.t3100 1.2605
R8221 VSS.n10470 VSS.t921 1.2605
R8222 VSS.t2113 VSS.n10474 1.2605
R8223 VSS.n10474 VSS.t3100 1.2605
R8224 VSS.n10583 VSS.t3312 1.2605
R8225 VSS.n10583 VSS.t3258 1.2605
R8226 VSS.n10580 VSS.t2832 1.2605
R8227 VSS.t2734 VSS.n10580 1.2605
R8228 VSS.n10576 VSS.t1854 1.2605
R8229 VSS.n10576 VSS.t2832 1.2605
R8230 VSS.n9037 VSS.t798 1.2605
R8231 VSS.t2874 VSS.n9037 1.2605
R8232 VSS.t3464 VSS.n1569 1.2605
R8233 VSS.n1569 VSS.t1082 1.2605
R8234 VSS.t3206 VSS.n9006 1.2605
R8235 VSS.n9006 VSS.t2171 1.2605
R8236 VSS.n8968 VSS.t2796 1.2605
R8237 VSS.t3472 VSS.n8968 1.2605
R8238 VSS.n9098 VSS.t2067 1.2605
R8239 VSS.t986 VSS.n9098 1.2605
R8240 VSS.t493 VSS.n8978 1.2605
R8241 VSS.n8978 VSS.t1666 1.2605
R8242 VSS.t2792 VSS.n9087 1.2605
R8243 VSS.n9087 VSS.t1736 1.2605
R8244 VSS.n9043 VSS.t1297 1.2605
R8245 VSS.t2337 VSS.n9043 1.2605
R8246 VSS.t2195 VSS.n9066 1.2605
R8247 VSS.n9066 VSS.t1102 1.2605
R8248 VSS.t1768 VSS.n9072 1.2605
R8249 VSS.n9072 VSS.t2447 1.2605
R8250 VSS.n973 VSS.t1914 1.2605
R8251 VSS.t2155 VSS.n973 1.2605
R8252 VSS.n967 VSS.t2185 1.2605
R8253 VSS.t1390 VSS.n967 1.2605
R8254 VSS.t917 VSS.n10270 1.2605
R8255 VSS.n10270 VSS.t1194 1.2605
R8256 VSS.t1240 VSS.n10276 1.2605
R8257 VSS.n10276 VSS.t3492 1.2605
R8258 VSS.n311 VSS.t3068 1.2605
R8259 VSS.t3266 VSS.n311 1.2605
R8260 VSS.n305 VSS.t2488 1.2605
R8261 VSS.t2459 VSS.n305 1.2605
R8262 VSS.n989 VSS.t871 1.2605
R8263 VSS.t1116 VSS.n989 1.2605
R8264 VSS.n983 VSS.t3422 1.2605
R8265 VSS.t3380 VSS.n983 1.2605
R8266 VSS.n1010 VSS.t2163 1.2605
R8267 VSS.t2373 VSS.n1010 1.2605
R8268 VSS.n1004 VSS.t2405 1.2605
R8269 VSS.t1632 VSS.n1004 1.2605
R8270 VSS.n10222 VSS.t1204 1.2605
R8271 VSS.t1473 VSS.n10222 1.2605
R8272 VSS.n317 VSS.t1495 1.2605
R8273 VSS.t594 VSS.n317 1.2605
R8274 VSS.t3194 VSS.n10210 1.2605
R8275 VSS.n10210 VSS.t3168 1.2605
R8276 VSS.t3444 VSS.n10216 1.2605
R8277 VSS.n10216 VSS.t3400 1.2605
R8278 VSS.n1022 VSS.t1038 1.2605
R8279 VSS.t999 VSS.n1022 1.2605
R8280 VSS.n1016 VSS.t1344 1.2605
R8281 VSS.t1304 VSS.n1016 1.2605
R8282 VSS.n1047 VSS.t2333 1.2605
R8283 VSS.t2305 VSS.n1047 1.2605
R8284 VSS.n1041 VSS.t1926 1.2605
R8285 VSS.t2946 VSS.n1041 1.2605
R8286 VSS.n374 VSS.t1422 1.2605
R8287 VSS.t1388 VSS.n374 1.2605
R8288 VSS.n368 VSS.t933 1.2605
R8289 VSS.t1984 VSS.n368 1.2605
R8290 VSS.n10162 VSS.t3414 1.2605
R8291 VSS.t3374 VSS.n10162 1.2605
R8292 VSS.n389 VSS.t2670 1.2605
R8293 VSS.t504 VSS.n389 1.2605
R8294 VSS.n1059 VSS.t1324 1.2605
R8295 VSS.t1279 VSS.n1059 1.2605
R8296 VSS.n1053 VSS.t3606 1.2605
R8297 VSS.t1564 VSS.n1053 1.2605
R8298 VSS.n1080 VSS.t3460 1.2605
R8299 VSS.t2674 VSS.n1080 1.2605
R8300 VSS.n1074 VSS.t1904 1.2605
R8301 VSS.t2143 VSS.n1074 1.2605
R8302 VSS.t2522 VSS.n10150 1.2605
R8303 VSS.n10150 VSS.t1742 1.2605
R8304 VSS.t913 VSS.n10156 1.2605
R8305 VSS.n10156 VSS.t1182 1.2605
R8306 VSS.n1293 VSS.t3124 1.2605
R8307 VSS.t3316 VSS.n1293 1.2605
R8308 VSS.n1287 VSS.t3348 1.2605
R8309 VSS.t3612 VSS.n1287 1.2605
R8310 VSS.n1096 VSS.t950 1.2605
R8311 VSS.t1218 VSS.n1096 1.2605
R8312 VSS.n1090 VSS.t1249 1.2605
R8313 VSS.t1507 VSS.n1090 1.2605
R8314 VSS.n1117 VSS.t2686 1.2605
R8315 VSS.t2932 VSS.n1117 1.2605
R8316 VSS.n1111 VSS.t2151 1.2605
R8317 VSS.t1358 VSS.n1111 1.2605
R8318 VSS.n1129 VSS.t3610 1.2605
R8319 VSS.t3504 VSS.n1129 1.2605
R8320 VSS.n1123 VSS.t755 1.2605
R8321 VSS.t3104 VSS.n1123 1.2605
R8322 VSS.t2606 VSS.n865 1.2605
R8323 VSS.n865 VSS.t2868 1.2605
R8324 VSS.t2073 VSS.n876 1.2605
R8325 VSS.n876 VSS.t2045 1.2605
R8326 VSS.t3512 VSS.n10925 1.2605
R8327 VSS.n10925 VSS.t607 1.2605
R8328 VSS.t631 VSS.n841 1.2605
R8329 VSS.n841 VSS.t2990 1.2605
R8330 VSS.n10363 VSS.t2165 1.2605
R8331 VSS.t3446 VSS.n10363 1.2605
R8332 VSS.n10359 VSS.t1176 1.2605
R8333 VSS.n10359 VSS.t2165 1.2605
R8334 VSS.n10356 VSS.t583 1.2605
R8335 VSS.t1968 VSS.n10356 1.2605
R8336 VSS.t679 VSS.n10668 1.2605
R8337 VSS.n10668 VSS.t583 1.2605
R8338 VSS.n10671 VSS.t3264 1.2605
R8339 VSS.n10671 VSS.t3536 1.2605
R8340 VSS.t2301 VSS.n10675 1.2605
R8341 VSS.n10675 VSS.t3264 1.2605
R8342 VSS.n10406 VSS.t204 1.2605
R8343 VSS.n10406 VSS.t181 1.2605
R8344 VSS.n10407 VSS.t201 1.2605
R8345 VSS.n10407 VSS.t291 1.2605
R8346 VSS.n10399 VSS.t23 1.2605
R8347 VSS.n10399 VSS.t38 1.2605
R8348 VSS.n10400 VSS.t53 1.2605
R8349 VSS.n10400 VSS.t43 1.2605
R8350 VSS.n10393 VSS.t208 1.2605
R8351 VSS.n10393 VSS.t139 1.2605
R8352 VSS.n10395 VSS.t52 1.2605
R8353 VSS.n10395 VSS.t35 1.2605
R8354 VSS.n10389 VSS.t134 1.2605
R8355 VSS.n10389 VSS.t49 1.2605
R8356 VSS.n10387 VSS.t131 1.2605
R8357 VSS.n10387 VSS.t127 1.2605
R8358 VSS.n10624 VSS.t178 1.2605
R8359 VSS.n10624 VSS.t136 1.2605
R8360 VSS.n10615 VSS.t141 1.2605
R8361 VSS.n10615 VSS.t210 1.2605
R8362 VSS.n10379 VSS.t132 1.2605
R8363 VSS.n10379 VSS.t26 1.2605
R8364 VSS.n10373 VSS.t22 1.2605
R8365 VSS.n10373 VSS.t135 1.2605
R8366 VSS.n10300 VSS.t28 1.2605
R8367 VSS.n10300 VSS.t152 1.2605
R8368 VSS.n10296 VSS.t126 1.2605
R8369 VSS.n10296 VSS.t17 1.2605
R8370 VSS.n10323 VSS.t146 1.2605
R8371 VSS.n10323 VSS.t8 1.2605
R8372 VSS.n10324 VSS.t176 1.2605
R8373 VSS.n10324 VSS.t9 1.2605
R8374 VSS.n10327 VSS.t15 1.2605
R8375 VSS.n10327 VSS.t24 1.2605
R8376 VSS.n10328 VSS.t164 1.2605
R8377 VSS.n10328 VSS.t19 1.2605
R8378 VSS.n10316 VSS.t20 1.2605
R8379 VSS.n10316 VSS.t44 1.2605
R8380 VSS.n10317 VSS.t4 1.2605
R8381 VSS.n10317 VSS.t207 1.2605
R8382 VSS.n10312 VSS.t2 1.2605
R8383 VSS.n10312 VSS.t40 1.2605
R8384 VSS.n10313 VSS.t48 1.2605
R8385 VSS.n10313 VSS.t123 1.2605
R8386 VSS.n10307 VSS.t161 1.2605
R8387 VSS.n10307 VSS.t51 1.2605
R8388 VSS.n10304 VSS.t125 1.2605
R8389 VSS.n10304 VSS.t122 1.2605
R8390 VSS.n9472 VSS.t3008 1.2605
R8391 VSS.t1402 VSS.n9472 1.2605
R8392 VSS.t2037 VSS.n9432 1.2605
R8393 VSS.n9432 VSS.t3514 1.2605
R8394 VSS.t2476 VSS.n9457 1.2605
R8395 VSS.n9457 VSS.t1238 1.2605
R8396 VSS.n9451 VSS.t3086 1.2605
R8397 VSS.t1795 VSS.n9451 1.2605
R8398 VSS.n9613 VSS.t235 1.2605
R8399 VSS.n9613 VSS.t223 1.2605
R8400 VSS.n813 VSS.t226 1.2605
R8401 VSS.n813 VSS.t249 1.2605
R8402 VSS.t3172 VSS.n9977 1.2605
R8403 VSS.n9977 VSS.t1030 1.2605
R8404 VSS.t1023 VSS.n9983 1.2605
R8405 VSS.n9983 VSS.t2357 1.2605
R8406 VSS.t3146 VSS.n9989 1.2605
R8407 VSS.n9989 VSS.t3092 1.2605
R8408 VSS.t1852 VSS.n9999 1.2605
R8409 VSS.n9999 VSS.t2121 1.2605
R8410 VSS.t1584 VSS.n10005 1.2605
R8411 VSS.n10005 VSS.t736 1.2605
R8412 VSS.t2518 VSS.n10011 1.2605
R8413 VSS.n10011 VSS.t728 1.2605
R8414 VSS.t2345 VSS.n10023 1.2605
R8415 VSS.n10023 VSS.t3298 1.2605
R8416 VSS.n10028 VSS.t3296 1.2605
R8417 VSS.n10028 VSS.t3230 1.2605
R8418 VSS.t901 VSS.n9726 1.2605
R8419 VSS.n9726 VSS.t2243 1.2605
R8420 VSS.t2516 VSS.n9736 1.2605
R8421 VSS.n9736 VSS.t3478 1.2605
R8422 VSS.t3474 VSS.n9742 1.2605
R8423 VSS.n9742 VSS.t1734 1.2605
R8424 VSS.t1724 VSS.n9748 1.2605
R8425 VSS.n9748 VSS.t1656 1.2605
R8426 VSS.t1196 VSS.n9758 1.2605
R8427 VSS.n9758 VSS.t1491 1.2605
R8428 VSS.n9762 VSS.t2231 1.2605
R8429 VSS.n9762 VSS.t3196 1.2605
R8430 VSS.n9632 VSS.t1886 1.2605
R8431 VSS.t1060 VSS.n9632 1.2605
R8432 VSS.t1383 VSS.n1361 1.2605
R8433 VSS.n1361 VSS.t2698 1.2605
R8434 VSS.t2684 VSS.n1367 1.2605
R8435 VSS.n1367 VSS.t2586 1.2605
R8436 VSS.t3328 VSS.n1373 1.2605
R8437 VSS.n1373 VSS.t1624 1.2605
R8438 VSS.n9973 VSS.t1906 1.2605
R8439 VSS.t806 VSS.n9973 1.2605
R8440 VSS.n9971 VSS.t2297 1.2605
R8441 VSS.t3030 VSS.n9971 1.2605
R8442 VSS.n9969 VSS.t3390 1.2605
R8443 VSS.t2724 VSS.n9969 1.2605
R8444 VSS.n9941 VSS.t1392 1.2605
R8445 VSS.t2411 VSS.n9941 1.2605
R8446 VSS.n9939 VSS.t972 1.2605
R8447 VSS.t1799 VSS.n9939 1.2605
R8448 VSS.n9937 VSS.t1436 1.2605
R8449 VSS.t2119 VSS.n9937 1.2605
R8450 VSS.n575 VSS.t3154 1.2605
R8451 VSS.t2093 VSS.n575 1.2605
R8452 VSS.t3548 VSS.n570 1.2605
R8453 VSS.t2858 VSS.n570 1.2605
R8454 VSS.n9720 VSS.t3248 1.2605
R8455 VSS.t849 VSS.n9720 1.2605
R8456 VSS.n9669 VSS.t3166 1.2605
R8457 VSS.t2115 VSS.n9669 1.2605
R8458 VSS.n9667 VSS.t3564 1.2605
R8459 VSS.t1188 VSS.n9667 1.2605
R8460 VSS.n9664 VSS.t2656 1.2605
R8461 VSS.t1952 VSS.n9664 1.2605
R8462 VSS.n9637 VSS.t2630 1.2605
R8463 VSS.t518 VSS.n9637 1.2605
R8464 VSS.t992 VSS.n799 1.2605
R8465 VSS.t3080 VSS.n799 1.2605
R8466 VSS.n9630 VSS.t2688 1.2605
R8467 VSS.n9630 VSS.t3428 1.2605
R8468 VSS.n1352 VSS.t2654 1.2605
R8469 VSS.t3326 VSS.n1352 1.2605
R8470 VSS.n1350 VSS.t1762 1.2605
R8471 VSS.t996 VSS.n1350 1.2605
R8472 VSS.n1347 VSS.t1479 1.2605
R8473 VSS.t2167 VSS.n1347 1.2605
R8474 VSS.n670 VSS.t80 1.2605
R8475 VSS.n670 VSS.t88 1.2605
R8476 VSS.n9875 VSS.t87 1.2605
R8477 VSS.n9875 VSS.t55 1.2605
R8478 VSS.n669 VSS.t57 1.2605
R8479 VSS.n669 VSS.t71 1.2605
R8480 VSS.n9857 VSS.t75 1.2605
R8481 VSS.n9857 VSS.t61 1.2605
R8482 VSS.n9855 VSS.t81 1.2605
R8483 VSS.n9855 VSS.t72 1.2605
R8484 VSS.n655 VSS.t89 1.2605
R8485 VSS.n655 VSS.t82 1.2605
R8486 VSS.n676 VSS.t242 1.2605
R8487 VSS.n676 VSS.t252 1.2605
R8488 VSS.n674 VSS.t251 1.2605
R8489 VSS.n674 VSS.t227 1.2605
R8490 VSS.n651 VSS.t247 1.2605
R8491 VSS.n651 VSS.t225 1.2605
R8492 VSS.n820 VSS.t248 1.2605
R8493 VSS.n820 VSS.t238 1.2605
R8494 VSS.n818 VSS.t222 1.2605
R8495 VSS.n818 VSS.t244 1.2605
R8496 VSS.n816 VSS.t218 1.2605
R8497 VSS.n816 VSS.t241 1.2605
R8498 VSS.n11414 VSS.t64 1.2605
R8499 VSS.n11414 VSS.t77 1.2605
R8500 VSS.n46 VSS.t95 1.2605
R8501 VSS.n46 VSS.t69 1.2605
R8502 VSS.n45 VSS.t78 1.2605
R8503 VSS.n45 VSS.t85 1.2605
R8504 VSS.n11447 VSS.t67 1.2605
R8505 VSS.n11447 VSS.t84 1.2605
R8506 VSS.n21 VSS.t70 1.2605
R8507 VSS.n21 VSS.t86 1.2605
R8508 VSS.n20 VSS.t79 1.2605
R8509 VSS.n20 VSS.t90 1.2605
R8510 VSS.n9923 VSS.t76 1.2605
R8511 VSS.n9923 VSS.t59 1.2605
R8512 VSS.n9921 VSS.t74 1.2605
R8513 VSS.n9921 VSS.t58 1.2605
R8514 VSS.n585 VSS.t83 1.2605
R8515 VSS.n585 VSS.t73 1.2605
R8516 VSS.n9909 VSS.t94 1.2605
R8517 VSS.n9909 VSS.t93 1.2605
R8518 VSS.n9911 VSS.t92 1.2605
R8519 VSS.n9911 VSS.t91 1.2605
R8520 VSS.n9908 VSS.t66 1.2605
R8521 VSS.n9908 VSS.t62 1.2605
R8522 VSS.n9900 VSS.t221 1.2605
R8523 VSS.n9900 VSS.t237 1.2605
R8524 VSS.n9898 VSS.t234 1.2605
R8525 VSS.n9898 VSS.t243 1.2605
R8526 VSS.n629 VSS.t239 1.2605
R8527 VSS.n629 VSS.t254 1.2605
R8528 VSS.n1252 VSS.t240 1.2605
R8529 VSS.n1252 VSS.t253 1.2605
R8530 VSS.n1250 VSS.t250 1.2605
R8531 VSS.n1250 VSS.t230 1.2605
R8532 VSS.n1248 VSS.t228 1.2605
R8533 VSS.n1248 VSS.t236 1.2605
R8534 VSS.n1329 VSS.t246 1.2605
R8535 VSS.n1329 VSS.t245 1.2605
R8536 VSS.n9514 VSS.t216 1.2605
R8537 VSS.n9514 VSS.t214 1.2605
R8538 VSS.n1328 VSS.t233 1.2605
R8539 VSS.n1328 VSS.t231 1.2605
R8540 VSS.n812 VSS.t232 1.2605
R8541 VSS.n812 VSS.t219 1.2605
R8542 VSS.n10391 VSS.n10390 1.25428
R8543 VSS.n10397 VSS.n10396 1.25428
R8544 VSS.n10394 VSS.n10392 1.25428
R8545 VSS.n10409 VSS.n10405 1.25428
R8546 VSS.n10315 VSS.n10311 1.25428
R8547 VSS.n10321 VSS.n10319 1.25428
R8548 VSS.n10332 VSS.n10330 1.25428
R8549 VSS.n10306 VSS.n10305 1.25428
R8550 VSS.n11392 VSS.n11391 1.21249
R8551 VSS.n10611 VSS.n10439 1.13691
R8552 VSS.n10803 VSS.t42 1.1205
R8553 VSS.n10803 VSS.t130 1.1205
R8554 VSS.n10805 VSS.t211 1.1205
R8555 VSS.n10805 VSS.t205 1.1205
R8556 VSS.n10797 VSS.t203 1.1205
R8557 VSS.n10797 VSS.t209 1.1205
R8558 VSS.n10799 VSS.t6 1.1205
R8559 VSS.n10799 VSS.t46 1.1205
R8560 VSS.n10817 VSS.t1908 1.1205
R8561 VSS.t3204 VSS.n10817 1.1205
R8562 VSS.t581 VSS.n10751 1.1205
R8563 VSS.n10751 VSS.t889 1.1205
R8564 VSS.n10786 VSS.t2233 1.1205
R8565 VSS.t3544 VSS.n10786 1.1205
R8566 VSS.n10780 VSS.t962 1.1205
R8567 VSS.t1263 VSS.n10780 1.1205
R8568 VSS.n10442 VSS.t37 1.11868
R8569 VSS.t184 VSS.n10600 1.11868
R8570 VSS.n10663 VSS.t27 1.11868
R8571 VSS.n10383 VSS.n10382 0.9995
R8572 VSS.n10619 VSS.n10618 0.9995
R8573 VSS.n10628 VSS.n10627 0.9995
R8574 VSS.n10683 VSS.n10682 0.973625
R8575 VSS.n10612 VSS.n10611 0.970331
R8576 VSS.n9048 VSS.t3578 0.918039
R8577 VSS.n9049 VSS.t2806 0.918039
R8578 VSS.n1528 VSS.t3130 0.918039
R8579 VSS.n9119 VSS.t1938 0.918039
R8580 VSS.n9124 VSS.t1538 0.918039
R8581 VSS.n9128 VSS.t2900 0.918039
R8582 VSS.n9055 VSS.t1626 0.918039
R8583 VSS.n9052 VSS.t758 0.918039
R8584 VSS.n1529 VSS.t1096 0.918039
R8585 VSS.n9120 VSS.t3040 0.918039
R8586 VSS.n9125 VSS.t2608 0.918039
R8587 VSS.n9129 VSS.t866 0.918039
R8588 VSS.n9218 VSS.t1870 0.918039
R8589 VSS.n9219 VSS.t1035 0.918039
R8590 VSS.n9220 VSS.t1410 0.918039
R8591 VSS.n9221 VSS.t3270 0.918039
R8592 VSS.n9222 VSS.t2892 0.918039
R8593 VSS.n1509 VSS.t1147 0.918039
R8594 VSS.n9238 VSS.t1367 0.918039
R8595 VSS.n9235 VSS.t3630 0.918039
R8596 VSS.n9231 VSS.t832 0.918039
R8597 VSS.n9228 VSS.t2776 0.918039
R8598 VSS.n9224 VSS.t2347 0.918039
R8599 VSS.n1510 VSS.t572 0.918039
R8600 VSS.n1501 VSS.t1535 0.918039
R8601 VSS.n9270 VSS.t669 0.918039
R8602 VSS.n9275 VSS.t1005 0.918039
R8603 VSS.n9279 VSS.t2954 0.918039
R8604 VSS.n9284 VSS.t2526 0.918039
R8605 VSS.n9288 VSS.t780 0.918039
R8606 VSS.n1502 VSS.t722 0.918039
R8607 VSS.n9271 VSS.t3064 0.918039
R8608 VSS.n9276 VSS.t3322 0.918039
R8609 VSS.n9280 VSS.t2189 0.918039
R8610 VSS.n9285 VSS.t1786 0.918039
R8611 VSS.n9289 VSS.t3144 0.918039
R8612 VSS.n1479 VSS.t2774 0.918039
R8613 VSS.n1480 VSS.t1970 0.918039
R8614 VSS.n1481 VSS.t2277 0.918039
R8615 VSS.n1483 VSS.t1084 0.918039
R8616 VSS.n1484 VSS.t634 0.918039
R8617 VSS.n1485 VSS.t2059 0.918039
R8618 VSS.n9373 VSS.t2247 0.918039
R8619 VSS.n9370 VSS.t1481 0.918039
R8620 VSS.n9366 VSS.t1788 0.918039
R8621 VSS.n9363 VSS.t476 0.918039
R8622 VSS.n9359 VSS.t3250 0.918039
R8623 VSS.n9356 VSS.t1568 0.918039
R8624 VSS.n9389 VSS.t589 0.918039
R8625 VSS.n9393 VSS.t2952 0.918039
R8626 VSS.n9398 VSS.t3246 0.918039
R8627 VSS.n9402 VSS.t2065 0.918039
R8628 VSS.n9407 VSS.t1686 0.918039
R8629 VSS.n9411 VSS.t3060 0.918039
R8630 VSS.n9390 VSS.t1326 0.918039
R8631 VSS.n9394 VSS.t3584 0.918039
R8632 VSS.n9399 VSS.t800 0.918039
R8633 VSS.n9403 VSS.t2730 0.918039
R8634 VSS.n9408 VSS.t2317 0.918039
R8635 VSS.n9412 VSS.t523 0.918039
R8636 VSS.n1430 VSS.t2578 0.918039
R8637 VSS.n1431 VSS.t2938 0.918039
R8638 VSS.n1223 VSS.t1750 0.918039
R8639 VSS.n1224 VSS.t1336 0.918039
R8640 VSS.n1217 VSS.t2710 0.918039
R8641 VSS.n1436 VSS.t2818 0.918039
R8642 VSS.n1432 VSS.t3136 0.918039
R8643 VSS.n1230 VSS.t1942 0.918039
R8644 VSS.n1226 VSS.t1542 0.918039
R8645 VSS.n1218 VSS.t2910 0.918039
R8646 VSS.n791 VSS.t3484 0.918039
R8647 VSS.n1156 VSS.t688 0.918039
R8648 VSS.n1159 VSS.t2622 0.918039
R8649 VSS.n1160 VSS.t2219 0.918039
R8650 VSS.n1161 VSS.t3580 0.918039
R8651 VSS.n792 VSS.t1214 0.918039
R8652 VSS.n1157 VSS.t1546 0.918039
R8653 VSS.n9556 VSS.t3396 0.918039
R8654 VSS.n9552 VSS.t3044 0.918039
R8655 VSS.n9549 VSS.t1322 0.918039
R8656 VSS.n64 VSS.t3360 0.918039
R8657 VSS.n68 VSS.t556 0.918039
R8658 VSS.n71 VSS.t2524 0.918039
R8659 VSS.n75 VSS.t2129 0.918039
R8660 VSS.n80 VSS.t3476 0.918039
R8661 VSS.n1 VSS.t1086 0.918039
R8662 VSS.n2 VSS.t2580 0.918039
R8663 VSS.n104 VSS.t2936 0.918039
R8664 VSS.n112 VSS.t554 0.918039
R8665 VSS.n113 VSS.t1019 0.918039
R8666 VSS.n114 VSS.t1515 0.918039
R8667 VSS.n115 VSS.t3300 0.918039
R8668 VSS.n1571 VSS.t2746 0.918039
R8669 VSS.n1574 VSS.t1950 0.918039
R8670 VSS.n1578 VSS.t2269 0.918039
R8671 VSS.n8956 VSS.t1062 0.918039
R8672 VSS.n8960 VSS.t613 0.918039
R8673 VSS.n8963 VSS.t2039 0.918039
R8674 VSS.n1557 VSS.t1815 0.918039
R8675 VSS.n8981 VSS.t977 0.918039
R8676 VSS.n8986 VSS.t1350 0.918039
R8677 VSS.n8990 VSS.t3224 0.918039
R8678 VSS.n8995 VSS.t2842 0.918039
R8679 VSS.n8999 VSS.t1088 0.918039
R8680 VSS.n1558 VSS.t2602 0.918039
R8681 VSS.n8982 VSS.t1819 0.918039
R8682 VSS.n8987 VSS.t2139 0.918039
R8683 VSS.n8991 VSS.t906 0.918039
R8684 VSS.n8996 VSS.t3626 0.918039
R8685 VSS.n9000 VSS.t1922 0.918039
R8686 VSS.n9074 VSS.t980 0.918039
R8687 VSS.n9075 VSS.t3284 0.918039
R8688 VSS.n1534 VSS.t3618 0.918039
R8689 VSS.n1538 VSS.t2427 0.918039
R8690 VSS.n1539 VSS.t2024 0.918039
R8691 VSS.n1540 VSS.t3364 0.918039
R8692 VSS.n9081 VSS.t3508 0.918039
R8693 VSS.n9078 VSS.t2718 0.918039
R8694 VSS.n1535 VSS.t3050 0.918039
R8695 VSS.n9108 VSS.t1856 0.918039
R8696 VSS.n9104 VSS.t1467 0.918039
R8697 VSS.n9101 VSS.t2826 0.918039
R8698 VSS.n955 VSS.t1026 0.918039
R8699 VSS.n956 VSS.t1858 0.918039
R8700 VSS.n957 VSS.t2267 0.918039
R8701 VSS.n254 VSS.t2720 0.918039
R8702 VSS.n255 VSS.t1497 0.918039
R8703 VSS.n256 VSS.t3180 0.918039
R8704 VSS.n944 VSS.t2702 0.918039
R8705 VSS.n945 VSS.t3466 0.918039
R8706 VSS.n273 VSS.t776 0.918039
R8707 VSS.n10249 VSS.t1265 0.918039
R8708 VSS.n10254 VSS.t3116 0.918039
R8709 VSS.n10258 VSS.t1754 0.918039
R8710 VSS.n951 VSS.t705 0.918039
R8711 VSS.n948 VSS.t1554 0.918039
R8712 VSS.n274 VSS.t1958 0.918039
R8713 VSS.n10250 VSS.t2381 0.918039
R8714 VSS.n10255 VSS.t1149 0.918039
R8715 VSS.n10259 VSS.t2894 0.918039
R8716 VSS.n991 VSS.t1307 0.918039
R8717 VSS.n992 VSS.t2103 0.918039
R8718 VSS.n283 VSS.t2504 0.918039
R8719 VSS.n286 VSS.t2978 0.918039
R8720 VSS.n294 VSS.t1732 0.918039
R8721 VSS.n298 VSS.t3402 0.918039
R8722 VSS.n998 VSS.t2014 0.918039
R8723 VSS.n995 VSS.t2840 0.918039
R8724 VSS.n284 VSS.t3228 0.918039
R8725 VSS.n287 VSS.t502 0.918039
R8726 VSS.n295 VSS.t2431 0.918039
R8727 VSS.n299 VSS.t1056 0.918039
R8728 VSS.n931 VSS.t2467 0.918039
R8729 VSS.n932 VSS.t3280 0.918039
R8730 VSS.n323 VSS.t551 0.918039
R8731 VSS.n326 VSS.t1052 0.918039
R8732 VSS.n327 VSS.t2934 0.918039
R8733 VSS.n328 VSS.t1570 0.918039
R8734 VSS.n938 VSS.t2217 0.918039
R8735 VSS.n935 VSS.t3042 0.918039
R8736 VSS.n324 VSS.t3410 0.918039
R8737 VSS.n10232 VSS.t761 0.918039
R8738 VSS.n10228 VSS.t2640 0.918039
R8739 VSS.n10225 VSS.t1277 0.918039
R8740 VSS.n1024 VSS.t1850 0.918039
R8741 VSS.n1025 VSS.t2632 0.918039
R8742 VSS.n345 VSS.t3090 0.918039
R8743 VSS.n10189 VSS.t3488 0.918039
R8744 VSS.n10194 VSS.t2263 0.918039
R8745 VSS.n10198 VSS.t860 0.918039
R8746 VSS.n1031 VSS.t1112 0.918039
R8747 VSS.n1028 VSS.t1940 0.918039
R8748 VSS.n346 VSS.t2339 0.918039
R8749 VSS.n10190 VSS.t2814 0.918039
R8750 VSS.n10195 VSS.t1574 0.918039
R8751 VSS.n10199 VSS.t3262 0.918039
R8752 VSS.n918 VSS.t2742 0.918039
R8753 VSS.n919 VSS.t3532 0.918039
R8754 VSS.n355 VSS.t838 0.918039
R8755 VSS.n358 VSS.t1332 0.918039
R8756 VSS.n378 VSS.t3164 0.918039
R8757 VSS.n382 VSS.t1807 0.918039
R8758 VSS.n925 VSS.t878 0.918039
R8759 VSS.n922 VSS.t1716 0.918039
R8760 VSS.n356 VSS.t2127 0.918039
R8761 VSS.n359 VSS.t2558 0.918039
R8762 VSS.n379 VSS.t1338 0.918039
R8763 VSS.n383 VSS.t3074 0.918039
R8764 VSS.n1061 VSS.t1427 0.918039
R8765 VSS.n1062 VSS.t2205 0.918039
R8766 VSS.n395 VSS.t2610 0.918039
R8767 VSS.n398 VSS.t3094 0.918039
R8768 VSS.n399 VSS.t1832 0.918039
R8769 VSS.n400 VSS.t3528 0.918039
R8770 VSS.n1068 VSS.t2169 0.918039
R8771 VSS.n1065 VSS.t2974 0.918039
R8772 VSS.n396 VSS.t3338 0.918039
R8773 VSS.n10172 VSS.t691 0.918039
R8774 VSS.n10168 VSS.t2568 0.918039
R8775 VSS.n10165 VSS.t1212 0.918039
R8776 VSS.n905 VSS.t3424 0.918039
R8777 VSS.n906 VSS.t1155 0.918039
R8778 VSS.n417 VSS.t1609 0.918039
R8779 VSS.n10129 VSS.t2022 0.918039
R8780 VSS.n10134 VSS.t749 0.918039
R8781 VSS.n10138 VSS.t2486 0.918039
R8782 VSS.n912 VSS.t3540 0.918039
R8783 VSS.n909 VSS.t1271 0.918039
R8784 VSS.n418 VSS.t1698 0.918039
R8785 VSS.n10130 VSS.t2131 0.918039
R8786 VSS.n10135 VSS.t854 0.918039
R8787 VSS.n10139 VSS.t2594 0.918039
R8788 VSS.n1098 VSS.t990 0.918039
R8789 VSS.n1099 VSS.t1836 0.918039
R8790 VSS.n425 VSS.t2239 0.918039
R8791 VSS.n428 VSS.t2704 0.918039
R8792 VSS.n1276 VSS.t1475 0.918039
R8793 VSS.n1280 VSS.t3162 0.918039
R8794 VSS.n1105 VSS.t2097 0.918039
R8795 VSS.n1102 VSS.t2904 0.918039
R8796 VSS.n426 VSS.t3288 0.918039
R8797 VSS.n429 VSS.t605 0.918039
R8798 VSS.n1277 VSS.t2496 0.918039
R8799 VSS.n1281 VSS.t1122 0.918039
R8800 VSS.n843 VSS.t3028 0.918039
R8801 VSS.n844 VSS.t672 0.918039
R8802 VSS.n845 VSS.t1120 0.918039
R8803 VSS.n846 VSS.t1613 0.918039
R8804 VSS.n534 VSS.t3394 0.918039
R8805 VSS.n859 VSS.t574 0.918039
R8806 VSS.n856 VSS.t1477 0.918039
R8807 VSS.n852 VSS.t1874 0.918039
R8808 VSS.n849 VSS.t2299 0.918039
R8809 VSS.n535 VSS.t1048 0.918039
R8810 VSS.n1132 VSS.t927 0.918039
R8811 VSS.n1136 VSS.t1780 0.918039
R8812 VSS.n1141 VSS.t2191 0.918039
R8813 VSS.n1144 VSS.t2618 0.918039
R8814 VSS.n1145 VSS.t1406 0.918039
R8815 VSS.n1133 VSS.t2109 0.918039
R8816 VSS.n1137 VSS.t2912 0.918039
R8817 VSS.n1142 VSS.t3294 0.918039
R8818 VSS.n1150 VSS.t616 0.918039
R8819 VSS.n1146 VSS.t2514 0.918039
R8820 VSS.n880 VSS.t2772 0.918039
R8821 VSS.n881 VSS.t3558 0.918039
R8822 VSS.n882 VSS.t869 0.918039
R8823 VSS.n883 VSS.t1363 0.918039
R8824 VSS.n884 VSS.t3176 0.918039
R8825 VSS.n899 VSS.t651 0.918039
R8826 VSS.n896 VSS.t1529 0.918039
R8827 VSS.n892 VSS.t1936 0.918039
R8828 VSS.n889 VSS.t2365 0.918039
R8829 VSS.n885 VSS.t1107 0.918039
R8830 VSS.n224 VSS.t1334 0.918039
R8831 VSS.n231 VSS.t2125 0.918039
R8832 VSS.n232 VSS.t2532 0.918039
R8833 VSS.n233 VSS.t2994 0.918039
R8834 VSS.n234 VSS.t1758 0.918039
R8835 VSS.n10914 VSS.t1318 0.918039
R8836 VSS.n10907 VSS.t2107 0.918039
R8837 VSS.n10903 VSS.t2510 0.918039
R8838 VSS.n10900 VSS.t2984 0.918039
R8839 VSS.n10896 VSS.t1744 0.918039
R8840 VSS.n11000 VSS.t2592 0.918039
R8841 VSS.n11004 VSS.t3362 0.918039
R8842 VSS.n11009 VSS.t682 0.918039
R8843 VSS.n11013 VSS.t1168 0.918039
R8844 VSS.n11018 VSS.t3038 0.918039
R8845 VSS.n11001 VSS.t2245 0.918039
R8846 VSS.n11005 VSS.t3072 0.918039
R8847 VSS.n11010 VSS.t3434 0.918039
R8848 VSS.n11014 VSS.t784 0.918039
R8849 VSS.n11019 VSS.t2664 0.918039
R8850 VSS.n98 VSS.t734 0.918039
R8851 VSS.n11061 VSS.t1582 0.918039
R8852 VSS.n11066 VSS.t1990 0.918039
R8853 VSS.n11070 VSS.t2413 0.918039
R8854 VSS.n11075 VSS.t1172 0.918039
R8855 VSS.n99 VSS.t2006 0.918039
R8856 VSS.n11062 VSS.t2828 0.918039
R8857 VSS.n11067 VSS.t3220 0.918039
R8858 VSS.n11071 VSS.t491 0.918039
R8859 VSS.n11076 VSS.t2419 0.918039
R8860 VSS.n11205 VSS.t2666 0.918039
R8861 VSS.n11206 VSS.t3002 0.918039
R8862 VSS.n11207 VSS.t1811 0.918039
R8863 VSS.n11208 VSS.t1420 0.918039
R8864 VSS.n86 VSS.t2768 0.918039
R8865 VSS.n11221 VSS.t2159 0.918039
R8866 VSS.n11217 VSS.t2455 0.918039
R8867 VSS.n11214 VSS.t1285 0.918039
R8868 VSS.n11210 VSS.t845 0.918039
R8869 VSS.n87 VSS.t2249 0.918039
R8870 VSS.n10953 VSS.t3240 0.918039
R8871 VSS.n10958 VSS.t3570 0.918039
R8872 VSS.n10962 VSS.t2377 0.918039
R8873 VSS.n10967 VSS.t1992 0.918039
R8874 VSS.n10971 VSS.t3318 0.918039
R8875 VSS.n10954 VSS.t2956 0.918039
R8876 VSS.n10959 VSS.t3252 0.918039
R8877 VSS.n10963 VSS.t2071 0.918039
R8878 VSS.n10968 VSS.t1692 0.918039
R8879 VSS.n10972 VSS.t3066 0.918039
R8880 VSS.n707 VSS.t2343 0.918039
R8881 VSS.n708 VSS.t2696 0.918039
R8882 VSS.n709 VSS.t1517 0.918039
R8883 VSS.n710 VSS.t1065 0.918039
R8884 VSS.n210 VSS.t2449 0.918039
R8885 VSS.n723 VSS.t1254 0.918039
R8886 VSS.n719 VSS.t1588 0.918039
R8887 VSS.n716 VSS.t3442 0.918039
R8888 VSS.n712 VSS.t3096 0.918039
R8889 VSS.n211 VSS.t1365 0.918039
R8890 VSS.n766 VSS.t828 0.918039
R8891 VSS.n1171 VSS.t1174 0.918039
R8892 VSS.n1187 VSS.t3108 0.918039
R8893 VSS.n1192 VSS.t2692 0.918039
R8894 VSS.n1196 VSS.t929 0.918039
R8895 VSS.n767 VSS.t3320 0.918039
R8896 VSS.n1172 VSS.t499 0.918039
R8897 VSS.n1188 VSS.t2471 0.918039
R8898 VSS.n1193 VSS.t2085 0.918039
R8899 VSS.n1197 VSS.t3432 0.918039
R8900 VSS.n1519 VSS.t535 0.918039
R8901 VSS.n9148 VSS.t2916 0.918039
R8902 VSS.n9153 VSS.t3212 0.918039
R8903 VSS.n9157 VSS.t2028 0.918039
R8904 VSS.n9162 VSS.t1650 0.918039
R8905 VSS.n9166 VSS.t3020 0.918039
R8906 VSS.n1520 VSS.t2141 0.918039
R8907 VSS.n9149 VSS.t1361 0.918039
R8908 VSS.n9154 VSS.t1678 0.918039
R8909 VSS.n9158 VSS.t3552 0.918039
R8910 VSS.n9163 VSS.t3156 0.918039
R8911 VSS.n9167 VSS.t1458 0.918039
R8912 VSS.n9048 VSS.t2896 0.91749
R8913 VSS.n9049 VSS.t2075 0.91749
R8914 VSS.n1528 VSS.t2387 0.91749
R8915 VSS.n9119 VSS.t1225 0.91749
R8916 VSS.n9124 VSS.t773 0.91749
R8917 VSS.n9128 VSS.t2193 0.91749
R8918 VSS.n9055 VSS.t1784 0.91749
R8919 VSS.n9052 VSS.t938 0.91749
R8920 VSS.n1529 VSS.t1292 0.91749
R8921 VSS.n9120 VSS.t3186 0.91749
R8922 VSS.n9125 VSS.t2800 0.91749
R8923 VSS.n9129 VSS.t1042 0.91749
R8924 VSS.n9218 VSS.t2930 0.91749
R8925 VSS.n9219 VSS.t2123 0.91749
R8926 VSS.n9220 VSS.t2429 0.91749
R8927 VSS.n9221 VSS.t1259 0.91749
R8928 VSS.n9222 VSS.t815 0.91749
R8929 VSS.n1509 VSS.t2213 0.91749
R8930 VSS.n9238 VSS.t3334 0.91749
R8931 VSS.n9235 VSS.t2564 0.91749
R8932 VSS.n9231 VSS.t2908 0.91749
R8933 VSS.n9228 VSS.t1720 0.91749
R8934 VSS.n9224 VSS.t1316 0.91749
R8935 VSS.n1510 VSS.t2676 0.91749
R8936 VSS.n1501 VSS.t2562 0.91749
R8937 VSS.n9270 VSS.t1792 0.91749
R8938 VSS.n9275 VSS.t2101 0.91749
R8939 VSS.n9279 VSS.t885 0.91749
R8940 VSS.n9284 VSS.t3576 0.91749
R8941 VSS.n9288 VSS.t1878 0.91749
R8942 VSS.n1502 VSS.t2798 0.91749
R8943 VSS.n9271 VSS.t1986 0.91749
R8944 VSS.n9276 VSS.t2293 0.91749
R8945 VSS.n9280 VSS.t1092 0.91749
R8946 VSS.n9285 VSS.t648 0.91749
R8947 VSS.n9289 VSS.t2069 0.91749
R8948 VSS.n1479 VSS.t3454 0.91749
R8949 VSS.n1480 VSS.t2680 0.91749
R8950 VSS.n1481 VSS.t3016 0.91749
R8951 VSS.n1483 VSS.t1824 0.91749
R8952 VSS.n1484 VSS.t1432 0.91749
R8953 VSS.n1485 VSS.t2782 0.91749
R8954 VSS.n9373 VSS.t1178 0.91749
R8955 VSS.n9370 VSS.t3458 0.91749
R8956 VSS.n9366 VSS.t654 0.91749
R8957 VSS.n9363 VSS.t2604 0.91749
R8958 VSS.n9359 VSS.t2209 0.91749
R8959 VSS.n9356 VSS.t3562 0.91749
R8960 VSS.n9389 VSS.t2690 0.91749
R8961 VSS.n9393 VSS.t1884 0.91749
R8962 VSS.n9398 VSS.t2207 0.91749
R8963 VSS.n9402 VSS.t984 0.91749
R8964 VSS.n9407 VSS.t529 0.91749
R8965 VSS.n9411 VSS.t1978 0.91749
R8966 VSS.n9390 VSS.t2012 0.91749
R8967 VSS.n9394 VSS.t1223 0.91749
R8968 VSS.n9399 VSS.t1562 0.91749
R8969 VSS.n9403 VSS.t3408 0.91749
R8970 VSS.n9408 VSS.t3052 0.91749
R8971 VSS.n9412 VSS.t1330 0.91749
R8972 VSS.n1430 VSS.t1552 0.91749
R8973 VSS.n1431 VSS.t1866 0.91749
R8974 VSS.n1223 VSS.t610 0.91749
R8975 VSS.n1224 VSS.t3314 0.91749
R8976 VSS.n1217 VSS.t1654 0.91749
R8977 VSS.n1436 VSS.t3502 0.91749
R8978 VSS.n1432 VSS.t709 0.91749
R8979 VSS.n1230 VSS.t2644 0.91749
R8980 VSS.n1226 VSS.t2235 0.91749
R8981 VSS.n1218 VSS.t3594 0.91749
R8982 VSS.n791 VSS.t2421 0.91749
R8983 VSS.n1156 VSS.t2762 0.91749
R8984 VSS.n1159 VSS.t1597 0.91749
R8985 VSS.n1160 VSS.t1158 0.91749
R8986 VSS.n1161 VSS.t2530 0.91749
R8987 VSS.n792 VSS.t1930 0.91749
R8988 VSS.n1157 VSS.t2237 0.91749
R8989 VSS.n9556 VSS.t1032 0.91749
R8990 VSS.n9552 VSS.t577 0.91749
R8991 VSS.n9549 VSS.t2010 0.91749
R8992 VSS.n64 VSS.t2325 0.91749
R8993 VSS.n68 VSS.t2658 0.91749
R8994 VSS.n71 VSS.t1499 0.91749
R8995 VSS.n75 VSS.t1040 0.91749
R8996 VSS.n80 VSS.t2417 0.91749
R8997 VSS.n1 VSS.t3142 0.91749
R8998 VSS.n2 VSS.t462 0.91749
R8999 VSS.n104 VSS.t3160 0.91749
R9000 VSS.n112 VSS.t835 0.91749
R9001 VSS.n113 VSS.t1290 0.91749
R9002 VSS.n114 VSS.t1752 0.91749
R9003 VSS.n115 VSS.t3568 0.91749
R9004 VSS.n1571 VSS.t1704 0.91749
R9005 VSS.n1574 VSS.t857 0.91749
R9006 VSS.n1578 VSS.t1216 0.91749
R9007 VSS.n8956 VSS.t3122 0.91749
R9008 VSS.n8960 VSS.t2714 0.91749
R9009 VSS.n8963 VSS.t958 0.91749
R9010 VSS.n1557 VSS.t2574 0.91749
R9011 VSS.n8981 VSS.t1805 0.91749
R9012 VSS.n8986 VSS.t2117 0.91749
R9013 VSS.n8990 VSS.t897 0.91749
R9014 VSS.n8995 VSS.t3592 0.91749
R9015 VSS.n8999 VSS.t1896 0.91749
R9016 VSS.n1558 VSS.t3292 0.91749
R9017 VSS.n8982 VSS.t2508 0.91749
R9018 VSS.n8987 VSS.t2854 0.91749
R9019 VSS.n8991 VSS.t1676 0.91749
R9020 VSS.n8996 VSS.t1257 0.91749
R9021 VSS.n9000 VSS.t2616 0.91749
R9022 VSS.n9074 VSS.t3070 0.91749
R9023 VSS.n9075 VSS.t2241 0.91749
R9024 VSS.n1534 VSS.t2554 0.91749
R9025 VSS.n1538 VSS.t1404 0.91749
R9026 VSS.n1539 VSS.t945 0.91749
R9027 VSS.n1540 VSS.t2329 0.91749
R9028 VSS.n9081 VSS.t1505 0.91749
R9029 VSS.n9078 VSS.t619 0.91749
R9030 VSS.n1535 VSS.t974 0.91749
R9031 VSS.n9108 VSS.t2920 0.91749
R9032 VSS.n9104 VSS.t2469 0.91749
R9033 VSS.n9101 VSS.t743 0.91749
R9034 VSS.n955 VSS.t1295 0.91749
R9035 VSS.n956 VSS.t2089 0.91749
R9036 VSS.n957 VSS.t2492 0.91749
R9037 VSS.n254 VSS.t2972 0.91749
R9038 VSS.n255 VSS.t1722 0.91749
R9039 VSS.n256 VSS.t3392 0.91749
R9040 VSS.n944 VSS.t2566 0.91749
R9041 VSS.n945 VSS.t3336 0.91749
R9042 VSS.n273 VSS.t645 0.91749
R9043 VSS.n10249 VSS.t1129 0.91749
R9044 VSS.n10254 VSS.t3014 0.91749
R9045 VSS.n10258 VSS.t1644 0.91749
R9046 VSS.n951 VSS.t3034 0.91749
R9047 VSS.n948 VSS.t685 0.91749
R9048 VSS.n274 VSS.t1133 0.91749
R9049 VSS.n10250 VSS.t1620 0.91749
R9050 VSS.n10255 VSS.t3404 0.91749
R9051 VSS.n10259 VSS.t2063 0.91749
R9052 VSS.n991 VSS.t1556 0.91749
R9053 VSS.n992 VSS.t2327 0.91749
R9054 VSS.n283 VSS.t2758 0.91749
R9055 VSS.n286 VSS.t3192 0.91749
R9056 VSS.n294 VSS.t1960 0.91749
R9057 VSS.n298 VSS.t488 0.91749
R9058 VSS.n998 VSS.t1994 0.91749
R9059 VSS.n995 VSS.t2804 0.91749
R9060 VSS.n284 VSS.t3198 0.91749
R9061 VSS.n287 VSS.t460 0.91749
R9062 VSS.n295 VSS.t2395 0.91749
R9063 VSS.n299 VSS.t1009 0.91749
R9064 VSS.n931 VSS.t3506 0.91749
R9065 VSS.n932 VSS.t1233 0.91749
R9066 VSS.n323 VSS.t1662 0.91749
R9067 VSS.n326 VSS.t2079 0.91749
R9068 VSS.n327 VSS.t812 0.91749
R9069 VSS.n328 VSS.t2550 0.91749
R9070 VSS.n938 VSS.t3482 0.91749
R9071 VSS.n935 VSS.t1208 0.91749
R9072 VSS.n324 VSS.t1646 0.91749
R9073 VSS.n10232 VSS.t2061 0.91749
R9074 VSS.n10228 VSS.t793 0.91749
R9075 VSS.n10225 VSS.t2536 0.91749
R9076 VSS.n1024 VSS.t2870 0.91749
R9077 VSS.n1025 VSS.t465 0.91749
R9078 VSS.n345 VSS.t956 0.91749
R9079 VSS.n10189 VSS.t1452 0.91749
R9080 VSS.n10194 VSS.t3260 0.91749
R9081 VSS.n10198 VSS.t1918 0.91749
R9082 VSS.n1031 VSS.t2161 0.91749
R9083 VSS.n1028 VSS.t2970 0.91749
R9084 VSS.n346 VSS.t3330 0.91749
R9085 VSS.n10190 VSS.t677 0.91749
R9086 VSS.n10195 VSS.t2560 0.91749
R9087 VSS.n10199 VSS.t1202 0.91749
R9088 VSS.n918 VSS.t2716 0.91749
R9089 VSS.n919 VSS.t3500 0.91749
R9090 VSS.n355 VSS.t809 0.91749
R9091 VSS.n358 VSS.t1283 0.91749
R9092 VSS.n378 VSS.t3140 0.91749
R9093 VSS.n382 VSS.t1782 0.91749
R9094 VSS.n925 VSS.t1127 0.91749
R9095 VSS.n922 VSS.t1948 0.91749
R9096 VSS.n356 VSS.t2353 0.91749
R9097 VSS.n359 VSS.t2824 0.91749
R9098 VSS.n379 VSS.t1590 0.91749
R9099 VSS.n383 VSS.t3272 0.91749
R9100 VSS.n1061 VSS.t1386 0.91749
R9101 VSS.n1062 VSS.t2175 0.91749
R9102 VSS.n395 VSS.t2572 0.91749
R9103 VSS.n398 VSS.t3046 0.91749
R9104 VSS.n399 VSS.t1803 0.91749
R9105 VSS.n400 VSS.t3494 0.91749
R9106 VSS.n1068 VSS.t2379 0.91749
R9107 VSS.n1065 VSS.t3188 0.91749
R9108 VSS.n396 VSS.t3604 0.91749
R9109 VSS.n10172 VSS.t948 0.91749
R9110 VSS.n10168 VSS.t2838 0.91749
R9111 VSS.n10165 VSS.t1483 0.91749
R9112 VSS.n905 VSS.t2646 0.91749
R9113 VSS.n906 VSS.t3412 0.91749
R9114 VSS.n417 VSS.t741 0.91749
R9115 VSS.n10129 VSS.t1231 0.91749
R9116 VSS.n10134 VSS.t3098 0.91749
R9117 VSS.n10138 VSS.t1708 0.91749
R9118 VSS.n912 VSS.t642 0.91749
R9119 VSS.n909 VSS.t1525 0.91749
R9120 VSS.n418 VSS.t1934 0.91749
R9121 VSS.n10130 VSS.t2355 0.91749
R9122 VSS.n10135 VSS.t1100 0.91749
R9123 VSS.n10139 VSS.t2856 0.91749
R9124 VSS.n1098 VSS.t1273 0.91749
R9125 VSS.n1099 VSS.t2055 0.91749
R9126 VSS.n425 VSS.t2461 0.91749
R9127 VSS.n428 VSS.t2944 0.91749
R9128 VSS.n1276 VSS.t1700 0.91749
R9129 VSS.n1280 VSS.t3370 0.91749
R9130 VSS.n1105 VSS.t1288 0.91749
R9131 VSS.n1102 VSS.t2081 0.91749
R9132 VSS.n426 VSS.t2484 0.91749
R9133 VSS.n429 VSS.t2966 0.91749
R9134 VSS.n1277 VSS.t1718 0.91749
R9135 VSS.n1281 VSS.t3388 0.91749
R9136 VSS.n843 VSS.t3236 0.91749
R9137 VSS.n844 VSS.t931 0.91749
R9138 VSS.n845 VSS.t1408 0.91749
R9139 VSS.n846 VSS.t1838 0.91749
R9140 VSS.n534 VSS.t479 0.91749
R9141 VSS.n859 VSS.t538 0.91749
R9142 VSS.n856 VSS.t1444 0.91749
R9143 VSS.n852 VSS.t1844 0.91749
R9144 VSS.n849 VSS.t2271 0.91749
R9145 VSS.n535 VSS.t1003 0.91749
R9146 VSS.n1132 VSS.t1198 0.91749
R9147 VSS.n1136 VSS.t2000 0.91749
R9148 VSS.n1141 VSS.t2407 0.91749
R9149 VSS.n1144 VSS.t2878 0.91749
R9150 VSS.n1145 VSS.t1640 0.91749
R9151 VSS.n1133 VSS.t1301 0.91749
R9152 VSS.n1137 VSS.t2099 0.91749
R9153 VSS.n1142 VSS.t2500 0.91749
R9154 VSS.n1150 VSS.t2976 0.91749
R9155 VSS.n1146 VSS.t1730 0.91749
R9156 VSS.n880 VSS.t3022 0.91749
R9157 VSS.n881 VSS.t666 0.91749
R9158 VSS.n882 VSS.t1114 0.91749
R9159 VSS.n883 VSS.t1601 0.91749
R9160 VSS.n884 VSS.t3384 0.91749
R9161 VSS.n899 VSS.t3006 0.91749
R9162 VSS.n896 VSS.t639 0.91749
R9163 VSS.n892 VSS.t1098 0.91749
R9164 VSS.n889 VSS.t1586 0.91749
R9165 VSS.n885 VSS.t3372 0.91749
R9166 VSS.n224 VSS.t1578 0.91749
R9167 VSS.n231 VSS.t2341 0.91749
R9168 VSS.n232 VSS.t2786 0.91749
R9169 VSS.n233 VSS.t3208 0.91749
R9170 VSS.n234 VSS.t1982 0.91749
R9171 VSS.n10914 VSS.t2309 0.91749
R9172 VSS.n10907 VSS.t3134 0.91749
R9173 VSS.n10903 VSS.t3530 0.91749
R9174 VSS.n10900 VSS.t864 0.91749
R9175 VSS.n10896 VSS.t2736 0.91749
R9176 VSS.n11000 VSS.t3602 0.91749
R9177 VSS.n11004 VSS.t1340 0.91749
R9178 VSS.n11009 VSS.t1766 0.91749
R9179 VSS.n11013 VSS.t2197 0.91749
R9180 VSS.n11018 VSS.t909 0.91749
R9181 VSS.n11001 VSS.t3242 0.91749
R9182 VSS.n11005 VSS.t942 0.91749
R9183 VSS.n11010 VSS.t1418 0.91749
R9184 VSS.n11014 VSS.t1846 0.91749
R9185 VSS.n11019 VSS.t496 0.91749
R9186 VSS.n98 VSS.t693 0.91749
R9187 VSS.n11061 VSS.t1544 0.91749
R9188 VSS.n11066 VSS.t1954 0.91749
R9189 VSS.n11070 VSS.t2375 0.91749
R9190 VSS.n11075 VSS.t1137 0.91749
R9191 VSS.n99 VSS.t2259 0.91749
R9192 VSS.n11062 VSS.t3082 0.91749
R9193 VSS.n11067 VSS.t3450 0.91749
R9194 VSS.n11071 VSS.t796 0.91749
R9195 VSS.n11076 VSS.t2682 0.91749
R9196 VSS.n11205 VSS.t569 0.91749
R9197 VSS.n11206 VSS.t919 0.91749
R9198 VSS.n11207 VSS.t2876 0.91749
R9199 VSS.n11208 VSS.t2443 0.91749
R9200 VSS.n86 VSS.t695 0.91749
R9201 VSS.n11221 VSS.t1071 0.91749
R9202 VSS.n11217 VSS.t1442 0.91749
R9203 VSS.n11214 VSS.t3290 0.91749
R9204 VSS.n11210 VSS.t2922 0.91749
R9205 VSS.n87 VSS.t1180 0.91749
R9206 VSS.n10953 VSS.t2538 0.91749
R9207 VSS.n10958 VSS.t2884 0.91749
R9208 VSS.n10962 VSS.t1702 0.91749
R9209 VSS.n10967 VSS.t1281 0.91749
R9210 VSS.n10971 VSS.t2642 0.91749
R9211 VSS.n10954 VSS.t2223 0.91749
R9212 VSS.n10959 VSS.t2542 0.91749
R9213 VSS.n10963 VSS.t1396 0.91749
R9214 VSS.n10968 VSS.t925 0.91749
R9215 VSS.n10972 VSS.t2319 0.91749
R9216 VSS.n707 VSS.t1313 0.91749
R9217 VSS.n708 VSS.t1642 0.91749
R9218 VSS.n709 VSS.t3518 0.91749
R9219 VSS.n710 VSS.t3128 0.91749
R9220 VSS.n210 VSS.t1424 0.91749
R9221 VSS.n723 VSS.t3616 0.91749
R9222 VSS.n719 VSS.t826 0.91749
R9223 VSS.n716 VSS.t2760 0.91749
R9224 VSS.n712 VSS.t2335 0.91749
R9225 VSS.n211 VSS.t559 0.91749
R9226 VSS.n766 VSS.t2898 0.91749
R9227 VSS.n1171 VSS.t3200 0.91749
R9228 VSS.n1187 VSS.t2018 0.91749
R9229 VSS.n1192 VSS.t1636 0.91749
R9230 VSS.n1196 VSS.t3004 0.91749
R9231 VSS.n767 VSS.t1342 0.91749
R9232 VSS.n1172 VSS.t1670 0.91749
R9233 VSS.n1188 VSS.t3542 0.91749
R9234 VSS.n1193 VSS.t3150 0.91749
R9235 VSS.n1197 VSS.t1450 0.91749
R9236 VSS.n1519 VSS.t3010 0.91749
R9237 VSS.n9148 VSS.t2201 0.91749
R9238 VSS.n9153 VSS.t2498 0.91749
R9239 VSS.n9157 VSS.t1346 0.91749
R9240 VSS.n9162 VSS.t892 0.91749
R9241 VSS.n9166 VSS.t2279 0.91749
R9242 VSS.n1520 VSS.t1448 0.91749
R9243 VSS.n9149 VSS.t546 0.91749
R9244 VSS.n9154 VSS.t911 0.91749
R9245 VSS.n9158 VSS.t2866 0.91749
R9246 VSS.n9163 VSS.t2437 0.91749
R9247 VSS.n9167 VSS.t674 0.91749
R9248 VSS.n10706 VSS.n121 0.823492
R9249 VSS.n120 VSS.n119 0.794733
R9250 VSS.n1182 VSS.t338 0.717763
R9251 VSS.n10612 VSS.n10411 0.585196
R9252 VSS.n10632 VSS.n10365 0.585196
R9253 VSS.n10686 VSS.n10292 0.585196
R9254 VSS.n10678 VSS.n10334 0.585196
R9255 VSS.n9102 VSS.n9101 0.582999
R9256 VSS.n9105 VSS.n9104 0.582999
R9257 VSS.n9109 VSS.n9108 0.582999
R9258 VSS.n1536 VSS.n1535 0.582999
R9259 VSS.n9079 VSS.n9078 0.582999
R9260 VSS.n9082 VSS.n9081 0.582999
R9261 VSS.n9102 VSS.n1540 0.582999
R9262 VSS.n9105 VSS.n1539 0.582999
R9263 VSS.n9109 VSS.n1538 0.582999
R9264 VSS.n1536 VSS.n1534 0.582999
R9265 VSS.n9079 VSS.n9075 0.582999
R9266 VSS.n9082 VSS.n9074 0.582999
R9267 VSS.n9001 VSS.n9000 0.582999
R9268 VSS.n8997 VSS.n8996 0.582999
R9269 VSS.n8992 VSS.n8991 0.582999
R9270 VSS.n8988 VSS.n8987 0.582999
R9271 VSS.n8983 VSS.n8982 0.582999
R9272 VSS.n1559 VSS.n1558 0.582999
R9273 VSS.n9001 VSS.n8999 0.582999
R9274 VSS.n8997 VSS.n8995 0.582999
R9275 VSS.n8992 VSS.n8990 0.582999
R9276 VSS.n8988 VSS.n8986 0.582999
R9277 VSS.n8983 VSS.n8981 0.582999
R9278 VSS.n1559 VSS.n1557 0.582999
R9279 VSS.n8964 VSS.n8963 0.582999
R9280 VSS.n8961 VSS.n8960 0.582999
R9281 VSS.n8957 VSS.n8956 0.582999
R9282 VSS.n1579 VSS.n1578 0.582999
R9283 VSS.n1575 VSS.n1574 0.582999
R9284 VSS.n1572 VSS.n1571 0.582999
R9285 VSS.n536 VSS.n535 0.582999
R9286 VSS.n850 VSS.n849 0.582999
R9287 VSS.n853 VSS.n852 0.582999
R9288 VSS.n857 VSS.n856 0.582999
R9289 VSS.n860 VSS.n859 0.582999
R9290 VSS.n536 VSS.n534 0.582999
R9291 VSS.n850 VSS.n846 0.582999
R9292 VSS.n853 VSS.n845 0.582999
R9293 VSS.n857 VSS.n844 0.582999
R9294 VSS.n860 VSS.n843 0.582999
R9295 VSS.n1147 VSS.n1146 0.582999
R9296 VSS.n1151 VSS.n1150 0.582999
R9297 VSS.n1143 VSS.n1142 0.582999
R9298 VSS.n1138 VSS.n1137 0.582999
R9299 VSS.n1134 VSS.n1133 0.582999
R9300 VSS.n1147 VSS.n1145 0.582999
R9301 VSS.n1151 VSS.n1144 0.582999
R9302 VSS.n1143 VSS.n1141 0.582999
R9303 VSS.n1138 VSS.n1136 0.582999
R9304 VSS.n1134 VSS.n1132 0.582999
R9305 VSS.n886 VSS.n885 0.582999
R9306 VSS.n890 VSS.n889 0.582999
R9307 VSS.n893 VSS.n892 0.582999
R9308 VSS.n897 VSS.n896 0.582999
R9309 VSS.n900 VSS.n899 0.582999
R9310 VSS.n886 VSS.n884 0.582999
R9311 VSS.n890 VSS.n883 0.582999
R9312 VSS.n893 VSS.n882 0.582999
R9313 VSS.n897 VSS.n881 0.582999
R9314 VSS.n900 VSS.n880 0.582999
R9315 VSS.n1282 VSS.n1281 0.582999
R9316 VSS.n1278 VSS.n1277 0.582999
R9317 VSS.n430 VSS.n429 0.582999
R9318 VSS.n427 VSS.n426 0.582999
R9319 VSS.n1103 VSS.n1102 0.582999
R9320 VSS.n1106 VSS.n1105 0.582999
R9321 VSS.n1282 VSS.n1280 0.582999
R9322 VSS.n1278 VSS.n1276 0.582999
R9323 VSS.n430 VSS.n428 0.582999
R9324 VSS.n427 VSS.n425 0.582999
R9325 VSS.n1103 VSS.n1099 0.582999
R9326 VSS.n1106 VSS.n1098 0.582999
R9327 VSS.n10140 VSS.n10139 0.582999
R9328 VSS.n10136 VSS.n10135 0.582999
R9329 VSS.n10131 VSS.n10130 0.582999
R9330 VSS.n419 VSS.n418 0.582999
R9331 VSS.n910 VSS.n909 0.582999
R9332 VSS.n913 VSS.n912 0.582999
R9333 VSS.n10140 VSS.n10138 0.582999
R9334 VSS.n10136 VSS.n10134 0.582999
R9335 VSS.n10131 VSS.n10129 0.582999
R9336 VSS.n419 VSS.n417 0.582999
R9337 VSS.n910 VSS.n906 0.582999
R9338 VSS.n913 VSS.n905 0.582999
R9339 VSS.n10166 VSS.n10165 0.582999
R9340 VSS.n10169 VSS.n10168 0.582999
R9341 VSS.n10173 VSS.n10172 0.582999
R9342 VSS.n397 VSS.n396 0.582999
R9343 VSS.n1066 VSS.n1065 0.582999
R9344 VSS.n1069 VSS.n1068 0.582999
R9345 VSS.n10166 VSS.n400 0.582999
R9346 VSS.n10169 VSS.n399 0.582999
R9347 VSS.n10173 VSS.n398 0.582999
R9348 VSS.n397 VSS.n395 0.582999
R9349 VSS.n1066 VSS.n1062 0.582999
R9350 VSS.n1069 VSS.n1061 0.582999
R9351 VSS.n384 VSS.n383 0.582999
R9352 VSS.n380 VSS.n379 0.582999
R9353 VSS.n360 VSS.n359 0.582999
R9354 VSS.n357 VSS.n356 0.582999
R9355 VSS.n923 VSS.n922 0.582999
R9356 VSS.n926 VSS.n925 0.582999
R9357 VSS.n384 VSS.n382 0.582999
R9358 VSS.n380 VSS.n378 0.582999
R9359 VSS.n360 VSS.n358 0.582999
R9360 VSS.n357 VSS.n355 0.582999
R9361 VSS.n923 VSS.n919 0.582999
R9362 VSS.n926 VSS.n918 0.582999
R9363 VSS.n10200 VSS.n10199 0.582999
R9364 VSS.n10196 VSS.n10195 0.582999
R9365 VSS.n10191 VSS.n10190 0.582999
R9366 VSS.n347 VSS.n346 0.582999
R9367 VSS.n1029 VSS.n1028 0.582999
R9368 VSS.n1032 VSS.n1031 0.582999
R9369 VSS.n10200 VSS.n10198 0.582999
R9370 VSS.n10196 VSS.n10194 0.582999
R9371 VSS.n10191 VSS.n10189 0.582999
R9372 VSS.n347 VSS.n345 0.582999
R9373 VSS.n1029 VSS.n1025 0.582999
R9374 VSS.n1032 VSS.n1024 0.582999
R9375 VSS.n10226 VSS.n10225 0.582999
R9376 VSS.n10229 VSS.n10228 0.582999
R9377 VSS.n10233 VSS.n10232 0.582999
R9378 VSS.n325 VSS.n324 0.582999
R9379 VSS.n936 VSS.n935 0.582999
R9380 VSS.n939 VSS.n938 0.582999
R9381 VSS.n10226 VSS.n328 0.582999
R9382 VSS.n10229 VSS.n327 0.582999
R9383 VSS.n10233 VSS.n326 0.582999
R9384 VSS.n325 VSS.n323 0.582999
R9385 VSS.n936 VSS.n932 0.582999
R9386 VSS.n939 VSS.n931 0.582999
R9387 VSS.n300 VSS.n299 0.582999
R9388 VSS.n296 VSS.n295 0.582999
R9389 VSS.n288 VSS.n287 0.582999
R9390 VSS.n285 VSS.n284 0.582999
R9391 VSS.n996 VSS.n995 0.582999
R9392 VSS.n999 VSS.n998 0.582999
R9393 VSS.n300 VSS.n298 0.582999
R9394 VSS.n296 VSS.n294 0.582999
R9395 VSS.n288 VSS.n286 0.582999
R9396 VSS.n285 VSS.n283 0.582999
R9397 VSS.n996 VSS.n992 0.582999
R9398 VSS.n999 VSS.n991 0.582999
R9399 VSS.n10260 VSS.n10259 0.582999
R9400 VSS.n10256 VSS.n10255 0.582999
R9401 VSS.n10251 VSS.n10250 0.582999
R9402 VSS.n275 VSS.n274 0.582999
R9403 VSS.n949 VSS.n948 0.582999
R9404 VSS.n952 VSS.n951 0.582999
R9405 VSS.n10260 VSS.n10258 0.582999
R9406 VSS.n10256 VSS.n10254 0.582999
R9407 VSS.n10251 VSS.n10249 0.582999
R9408 VSS.n275 VSS.n273 0.582999
R9409 VSS.n949 VSS.n945 0.582999
R9410 VSS.n952 VSS.n944 0.582999
R9411 VSS.n10278 VSS.n256 0.582999
R9412 VSS.n10280 VSS.n255 0.582999
R9413 VSS.n10283 VSS.n254 0.582999
R9414 VSS.n958 VSS.n957 0.582999
R9415 VSS.n961 VSS.n956 0.582999
R9416 VSS.n963 VSS.n955 0.582999
R9417 VSS.n10897 VSS.n10896 0.582999
R9418 VSS.n10901 VSS.n10900 0.582999
R9419 VSS.n10904 VSS.n10903 0.582999
R9420 VSS.n10908 VSS.n10907 0.582999
R9421 VSS.n10915 VSS.n10914 0.582999
R9422 VSS.n10897 VSS.n234 0.582999
R9423 VSS.n10901 VSS.n233 0.582999
R9424 VSS.n10904 VSS.n232 0.582999
R9425 VSS.n10908 VSS.n231 0.582999
R9426 VSS.n10915 VSS.n224 0.582999
R9427 VSS.n11020 VSS.n11019 0.582999
R9428 VSS.n11015 VSS.n11014 0.582999
R9429 VSS.n11011 VSS.n11010 0.582999
R9430 VSS.n11006 VSS.n11005 0.582999
R9431 VSS.n11002 VSS.n11001 0.582999
R9432 VSS.n11020 VSS.n11018 0.582999
R9433 VSS.n11015 VSS.n11013 0.582999
R9434 VSS.n11011 VSS.n11009 0.582999
R9435 VSS.n11006 VSS.n11004 0.582999
R9436 VSS.n11002 VSS.n11000 0.582999
R9437 VSS.n11077 VSS.n11076 0.582999
R9438 VSS.n11072 VSS.n11071 0.582999
R9439 VSS.n11068 VSS.n11067 0.582999
R9440 VSS.n11063 VSS.n11062 0.582999
R9441 VSS.n100 VSS.n99 0.582999
R9442 VSS.n11077 VSS.n11075 0.582999
R9443 VSS.n11072 VSS.n11070 0.582999
R9444 VSS.n11068 VSS.n11066 0.582999
R9445 VSS.n11063 VSS.n11061 0.582999
R9446 VSS.n100 VSS.n98 0.582999
R9447 VSS.n11326 VSS.n115 0.582999
R9448 VSS.n11329 VSS.n114 0.582999
R9449 VSS.n11331 VSS.n113 0.582999
R9450 VSS.n11334 VSS.n112 0.582999
R9451 VSS.n11339 VSS.n104 0.582999
R9452 VSS.n3 VSS.n2 0.582999
R9453 VSS.n3 VSS.n1 0.582999
R9454 VSS.n81 VSS.n80 0.582999
R9455 VSS.n76 VSS.n75 0.582999
R9456 VSS.n72 VSS.n71 0.582999
R9457 VSS.n69 VSS.n68 0.582999
R9458 VSS.n65 VSS.n64 0.582999
R9459 VSS.n88 VSS.n87 0.582999
R9460 VSS.n11211 VSS.n11210 0.582999
R9461 VSS.n11215 VSS.n11214 0.582999
R9462 VSS.n11218 VSS.n11217 0.582999
R9463 VSS.n11222 VSS.n11221 0.582999
R9464 VSS.n88 VSS.n86 0.582999
R9465 VSS.n11211 VSS.n11208 0.582999
R9466 VSS.n11215 VSS.n11207 0.582999
R9467 VSS.n11218 VSS.n11206 0.582999
R9468 VSS.n11222 VSS.n11205 0.582999
R9469 VSS.n10973 VSS.n10972 0.582999
R9470 VSS.n10969 VSS.n10968 0.582999
R9471 VSS.n10964 VSS.n10963 0.582999
R9472 VSS.n10960 VSS.n10959 0.582999
R9473 VSS.n10955 VSS.n10954 0.582999
R9474 VSS.n10973 VSS.n10971 0.582999
R9475 VSS.n10969 VSS.n10967 0.582999
R9476 VSS.n10964 VSS.n10962 0.582999
R9477 VSS.n10960 VSS.n10958 0.582999
R9478 VSS.n10955 VSS.n10953 0.582999
R9479 VSS.n212 VSS.n211 0.582999
R9480 VSS.n713 VSS.n712 0.582999
R9481 VSS.n717 VSS.n716 0.582999
R9482 VSS.n720 VSS.n719 0.582999
R9483 VSS.n724 VSS.n723 0.582999
R9484 VSS.n212 VSS.n210 0.582999
R9485 VSS.n713 VSS.n710 0.582999
R9486 VSS.n717 VSS.n709 0.582999
R9487 VSS.n720 VSS.n708 0.582999
R9488 VSS.n724 VSS.n707 0.582999
R9489 VSS.n1198 VSS.n1197 0.582999
R9490 VSS.n1194 VSS.n1193 0.582999
R9491 VSS.n1189 VSS.n1188 0.582999
R9492 VSS.n1173 VSS.n1172 0.582999
R9493 VSS.n768 VSS.n767 0.582999
R9494 VSS.n1198 VSS.n1196 0.582999
R9495 VSS.n1194 VSS.n1192 0.582999
R9496 VSS.n1189 VSS.n1187 0.582999
R9497 VSS.n1173 VSS.n1171 0.582999
R9498 VSS.n768 VSS.n766 0.582999
R9499 VSS.n9550 VSS.n9549 0.582999
R9500 VSS.n9553 VSS.n9552 0.582999
R9501 VSS.n9557 VSS.n9556 0.582999
R9502 VSS.n1158 VSS.n1157 0.582999
R9503 VSS.n793 VSS.n792 0.582999
R9504 VSS.n9550 VSS.n1161 0.582999
R9505 VSS.n9553 VSS.n1160 0.582999
R9506 VSS.n9557 VSS.n1159 0.582999
R9507 VSS.n1158 VSS.n1156 0.582999
R9508 VSS.n793 VSS.n791 0.582999
R9509 VSS.n1219 VSS.n1218 0.582999
R9510 VSS.n1227 VSS.n1226 0.582999
R9511 VSS.n1231 VSS.n1230 0.582999
R9512 VSS.n1433 VSS.n1432 0.582999
R9513 VSS.n1437 VSS.n1436 0.582999
R9514 VSS.n1219 VSS.n1217 0.582999
R9515 VSS.n1227 VSS.n1224 0.582999
R9516 VSS.n1231 VSS.n1223 0.582999
R9517 VSS.n1433 VSS.n1431 0.582999
R9518 VSS.n1437 VSS.n1430 0.582999
R9519 VSS.n9413 VSS.n9412 0.582999
R9520 VSS.n9409 VSS.n9408 0.582999
R9521 VSS.n9404 VSS.n9403 0.582999
R9522 VSS.n9400 VSS.n9399 0.582999
R9523 VSS.n9395 VSS.n9394 0.582999
R9524 VSS.n9391 VSS.n9390 0.582999
R9525 VSS.n9413 VSS.n9411 0.582999
R9526 VSS.n9409 VSS.n9407 0.582999
R9527 VSS.n9404 VSS.n9402 0.582999
R9528 VSS.n9400 VSS.n9398 0.582999
R9529 VSS.n9395 VSS.n9393 0.582999
R9530 VSS.n9391 VSS.n9389 0.582999
R9531 VSS.n9357 VSS.n9356 0.582999
R9532 VSS.n9360 VSS.n9359 0.582999
R9533 VSS.n9364 VSS.n9363 0.582999
R9534 VSS.n9367 VSS.n9366 0.582999
R9535 VSS.n9371 VSS.n9370 0.582999
R9536 VSS.n9374 VSS.n9373 0.582999
R9537 VSS.n9357 VSS.n1485 0.582999
R9538 VSS.n9360 VSS.n1484 0.582999
R9539 VSS.n9364 VSS.n1483 0.582999
R9540 VSS.n9367 VSS.n1481 0.582999
R9541 VSS.n9371 VSS.n1480 0.582999
R9542 VSS.n9374 VSS.n1479 0.582999
R9543 VSS.n9290 VSS.n9289 0.582999
R9544 VSS.n9286 VSS.n9285 0.582999
R9545 VSS.n9281 VSS.n9280 0.582999
R9546 VSS.n9277 VSS.n9276 0.582999
R9547 VSS.n9272 VSS.n9271 0.582999
R9548 VSS.n1503 VSS.n1502 0.582999
R9549 VSS.n9290 VSS.n9288 0.582999
R9550 VSS.n9286 VSS.n9284 0.582999
R9551 VSS.n9281 VSS.n9279 0.582999
R9552 VSS.n9277 VSS.n9275 0.582999
R9553 VSS.n9272 VSS.n9270 0.582999
R9554 VSS.n1503 VSS.n1501 0.582999
R9555 VSS.n1511 VSS.n1510 0.582999
R9556 VSS.n9225 VSS.n9224 0.582999
R9557 VSS.n9229 VSS.n9228 0.582999
R9558 VSS.n9232 VSS.n9231 0.582999
R9559 VSS.n9236 VSS.n9235 0.582999
R9560 VSS.n9239 VSS.n9238 0.582999
R9561 VSS.n1511 VSS.n1509 0.582999
R9562 VSS.n9225 VSS.n9222 0.582999
R9563 VSS.n9229 VSS.n9221 0.582999
R9564 VSS.n9232 VSS.n9220 0.582999
R9565 VSS.n9236 VSS.n9219 0.582999
R9566 VSS.n9239 VSS.n9218 0.582999
R9567 VSS.n9168 VSS.n9167 0.582999
R9568 VSS.n9164 VSS.n9163 0.582999
R9569 VSS.n9159 VSS.n9158 0.582999
R9570 VSS.n9155 VSS.n9154 0.582999
R9571 VSS.n9150 VSS.n9149 0.582999
R9572 VSS.n1521 VSS.n1520 0.582999
R9573 VSS.n9168 VSS.n9166 0.582999
R9574 VSS.n9164 VSS.n9162 0.582999
R9575 VSS.n9159 VSS.n9157 0.582999
R9576 VSS.n9155 VSS.n9153 0.582999
R9577 VSS.n9150 VSS.n9148 0.582999
R9578 VSS.n1521 VSS.n1519 0.582999
R9579 VSS.n9130 VSS.n9129 0.582999
R9580 VSS.n9126 VSS.n9125 0.582999
R9581 VSS.n9121 VSS.n9120 0.582999
R9582 VSS.n1530 VSS.n1529 0.582999
R9583 VSS.n9053 VSS.n9052 0.582999
R9584 VSS.n9056 VSS.n9055 0.582999
R9585 VSS.n9130 VSS.n9128 0.582999
R9586 VSS.n9126 VSS.n9124 0.582999
R9587 VSS.n9121 VSS.n9119 0.582999
R9588 VSS.n1530 VSS.n1528 0.582999
R9589 VSS.n9053 VSS.n9049 0.582999
R9590 VSS.n9056 VSS.n9048 0.582999
R9591 VSS.n11292 VSS.t733 0.558372
R9592 VSS.n819 VSS.n817 0.489579
R9593 VSS.n675 VSS.n652 0.489579
R9594 VSS.n9858 VSS.n9856 0.489579
R9595 VSS.n9876 VSS.n9874 0.489579
R9596 VSS.n11415 VSS.n11413 0.489579
R9597 VSS.n11448 VSS.n11446 0.489579
R9598 VSS.n9516 VSS.n9515 0.489579
R9599 VSS.n1251 VSS.n1249 0.489579
R9600 VSS.n9899 VSS.n9897 0.489579
R9601 VSS.n9912 VSS.n9910 0.489579
R9602 VSS.n9924 VSS.n9922 0.489579
R9603 VSS.n9615 VSS.n9614 0.489579
R9604 VSS.n821 VSS.n819 0.486026
R9605 VSS.n677 VSS.n675 0.486026
R9606 VSS.n9856 VSS.n656 0.486026
R9607 VSS.n9877 VSS.n9876 0.486026
R9608 VSS.n11416 VSS.n11415 0.486026
R9609 VSS.n11449 VSS.n11448 0.486026
R9610 VSS.n9515 VSS.n9513 0.486026
R9611 VSS.n1253 VSS.n1251 0.486026
R9612 VSS.n9901 VSS.n9899 0.486026
R9613 VSS.n9913 VSS.n9912 0.486026
R9614 VSS.n9922 VSS.n9920 0.486026
R9615 VSS.n9614 VSS.n9612 0.486026
R9616 VSS.n11314 VSS.n121 0.465835
R9617 VSS.n60 VSS.n59 0.46265
R9618 VSS.n11391 VSS.n11390 0.458898
R9619 VSS.n11317 VSS.n34 0.3755
R9620 VSS.n11319 VSS.n11318 0.3755
R9621 VSS.n11393 VSS.n11392 0.3755
R9622 VSS.n11390 VSS.n11389 0.3755
R9623 VSS.n11316 VSS.n11315 0.3755
R9624 VSS.n11314 VSS.n11313 0.3755
R9625 VSS.n10866 VSS.n10865 0.3755
R9626 VSS.n4804 VSS.n121 0.347815
R9627 VSS.n9461 VSS.n9460 0.240145
R9628 VSS.n9459 VSS.n1379 0.240145
R9629 VSS.n10398 VSS.n10391 0.236091
R9630 VSS.n9460 VSS.n9459 0.207127
R9631 VSS.n10863 VSS.n10862 0.186214
R9632 VSS.n10862 VSS.n10861 0.186214
R9633 VSS.n10858 VSS.n10857 0.186214
R9634 VSS.n10859 VSS.n10858 0.186214
R9635 VSS.n10333 VSS.n10332 0.177184
R9636 VSS.n9142 VSS.n9141 0.174974
R9637 VSS.n1490 VSS.n1489 0.174974
R9638 VSS.n1210 VSS.n1209 0.174974
R9639 VSS.n10948 VSS.n10947 0.174974
R9640 VSS.n10994 VSS.n10993 0.174974
R9641 VSS.n8975 VSS.n8974 0.174974
R9642 VSS.n980 VSS.n979 0.174974
R9643 VSS.n1038 VSS.n1037 0.174974
R9644 VSS.n1087 VSS.n1086 0.174974
R9645 VSS.n873 VSS.n872 0.174974
R9646 VSS.n10765 VSS.n242 0.163
R9647 VSS.n10860 VSS.n242 0.163
R9648 VSS.n10758 VSS.n243 0.163
R9649 VSS.n10860 VSS.n243 0.163
R9650 VSS.n9462 VSS.n9461 0.160263
R9651 VSS.n9468 VSS.n1379 0.160263
R9652 VSS.n9196 VSS.n9193 0.157683
R9653 VSS.n9191 VSS.n9188 0.157683
R9654 VSS.n9332 VSS.n9329 0.157683
R9655 VSS.n9327 VSS.n9324 0.157683
R9656 VSS.n170 VSS.n167 0.157683
R9657 VSS.n165 VSS.n162 0.157683
R9658 VSS.n9578 VSS.n9575 0.157683
R9659 VSS.n9573 VSS.n9570 0.157683
R9660 VSS.n193 VSS.n190 0.157683
R9661 VSS.n198 VSS.n195 0.157683
R9662 VSS.n471 VSS.n468 0.157683
R9663 VSS.n476 VSS.n473 0.157683
R9664 VSS.n9029 VSS.n9026 0.157683
R9665 VSS.n9024 VSS.n9021 0.157683
R9666 VSS.n264 VSS.n261 0.157683
R9667 VSS.n269 VSS.n266 0.157683
R9668 VSS.n336 VSS.n333 0.157683
R9669 VSS.n341 VSS.n338 0.157683
R9670 VSS.n408 VSS.n405 0.157683
R9671 VSS.n413 VSS.n410 0.157683
R9672 VSS.n10864 VSS.n240 0.14444
R9673 VSS.n10853 VSS.n10852 0.141041
R9674 VSS.n10852 VSS.n245 0.141041
R9675 VSS.n10793 VSS.n249 0.141041
R9676 VSS.n10849 VSS.n249 0.141041
R9677 VSS.n10796 VSS.n10795 0.14
R9678 VSS.n10801 VSS.n10795 0.14
R9679 VSS.n10802 VSS.n10794 0.14
R9680 VSS.n10807 VSS.n10794 0.14
R9681 VSS.n10374 VSS.n10372 0.14
R9682 VSS.n10377 VSS.n10372 0.14
R9683 VSS.n10378 VSS.n10371 0.14
R9684 VSS.n10382 VSS.n10371 0.14
R9685 VSS.n10383 VSS.n10370 0.14
R9686 VSS.n10386 VSS.n10370 0.14
R9687 VSS.n10614 VSS.n10369 0.14
R9688 VSS.n10618 VSS.n10369 0.14
R9689 VSS.n10619 VSS.n10368 0.14
R9690 VSS.n10622 VSS.n10368 0.14
R9691 VSS.n10623 VSS.n10367 0.14
R9692 VSS.n10627 VSS.n10367 0.14
R9693 VSS.n10628 VSS.n10366 0.14
R9694 VSS.n10631 VSS.n10366 0.14
R9695 VSS.n10685 VSS.n10293 0.14
R9696 VSS.n10683 VSS.n10293 0.14
R9697 VSS.n10682 VSS.n10295 0.14
R9698 VSS.n10680 VSS.n10295 0.14
R9699 VSS.n10303 VSS.n10298 0.14
R9700 VSS.n10301 VSS.n10298 0.14
R9701 VSS.n10762 VSS.n10739 0.132207
R9702 VSS.n9142 VSS.n9140 0.130788
R9703 VSS.n1490 VSS.n1488 0.130788
R9704 VSS.n1210 VSS.n1208 0.130788
R9705 VSS.n10948 VSS.n10946 0.130788
R9706 VSS.n10994 VSS.n10992 0.130788
R9707 VSS.n8975 VSS.n8973 0.130788
R9708 VSS.n980 VSS.n978 0.130788
R9709 VSS.n1038 VSS.n1036 0.130788
R9710 VSS.n1087 VSS.n1085 0.130788
R9711 VSS.n873 VSS.n871 0.130788
R9712 VSS.n6908 VSS.n6907 0.109625
R9713 VSS.n8233 VSS.n1822 0.109625
R9714 VSS.n6906 VSS.n2263 0.109625
R9715 VSS.n8232 VSS.n8231 0.109625
R9716 VSS.n5469 VSS.n5468 0.10925
R9717 VSS.n4140 VSS.n3184 0.10925
R9718 VSS.n4142 VSS.n4141 0.10925
R9719 VSS.n5470 VSS.n2743 0.10925
R9720 VSS.n10782 VSS.n248 0.108833
R9721 VSS.n10850 VSS.n248 0.108833
R9722 VSS.n10851 VSS.n250 0.108833
R9723 VSS.n10851 VSS.n10850 0.108833
R9724 VSS.n10452 VSS.n10451 0.105988
R9725 VSS.n10478 VSS.n10477 0.105988
R9726 VSS.n10561 VSS.n10560 0.105988
R9727 VSS.n10690 VSS.n10689 0.105988
R9728 VSS.n10640 VSS.n10639 0.105988
R9729 VSS.n10656 VSS.n10655 0.102012
R9730 VSS.n10593 VSS.n10592 0.102012
R9731 VSS.n10613 VSS.n10386 0.10175
R9732 VSS.n10762 VSS.n10759 0.100659
R9733 VSS.n10864 VSS.n10863 0.0996408
R9734 VSS.n11303 VSS.n11302 0.0986132
R9735 VSS.n11302 VSS.n11301 0.0986132
R9736 VSS.n10845 VSS.n10844 0.0986132
R9737 VSS.n10846 VSS.n10845 0.0986132
R9738 VSS.n9440 VSS.n1381 0.0933571
R9739 VSS.n9303 VSS.n1381 0.0933571
R9740 VSS.n1382 VSS.n1344 0.0917281
R9741 VSS.n1392 VSS.n1382 0.0917281
R9742 VSS.n9156 VSS.n1525 0.0886356
R9743 VSS.n9179 VSS.n1525 0.0886356
R9744 VSS.n9176 VSS.n9175 0.0886356
R9745 VSS.n9177 VSS.n9176 0.0886356
R9746 VSS.n9156 VSS.n1514 0.0886356
R9747 VSS.n9178 VSS.n1514 0.0886356
R9748 VSS.n9230 VSS.n1515 0.0886356
R9749 VSS.n1517 VSS.n1515 0.0886356
R9750 VSS.n9251 VSS.n9250 0.0886356
R9751 VSS.n9250 VSS.n9249 0.0886356
R9752 VSS.n9230 VSS.n1506 0.0886356
R9753 VSS.n1516 VSS.n1506 0.0886356
R9754 VSS.n9278 VSS.n1507 0.0886356
R9755 VSS.n9306 VSS.n1507 0.0886356
R9756 VSS.n9298 VSS.n9297 0.0886356
R9757 VSS.n9299 VSS.n9298 0.0886356
R9758 VSS.n9278 VSS.n1497 0.0886356
R9759 VSS.n9305 VSS.n1497 0.0886356
R9760 VSS.n8955 VSS.n1562 0.0886356
R9761 VSS.n1564 VSS.n1562 0.0886356
R9762 VSS.n8989 VSS.n1563 0.0886356
R9763 VSS.n9012 VSS.n1563 0.0886356
R9764 VSS.n9009 VSS.n9008 0.0886356
R9765 VSS.n9010 VSS.n9009 0.0886356
R9766 VSS.n8989 VSS.n1555 0.0886356
R9767 VSS.n9011 VSS.n1555 0.0886356
R9768 VSS.n9110 VSS.n1537 0.0886356
R9769 VSS.n1537 VSS.n1533 0.0886356
R9770 VSS.n9094 VSS.n9093 0.0886356
R9771 VSS.n9093 VSS.n9092 0.0886356
R9772 VSS.n9111 VSS.n9110 0.0886356
R9773 VSS.n9112 VSS.n9111 0.0886356
R9774 VSS.n9118 VSS.n9117 0.0886356
R9775 VSS.n9117 VSS.n9116 0.0886356
R9776 VSS.n1547 VSS.n1532 0.0886356
R9777 VSS.n9113 VSS.n1532 0.0886356
R9778 VSS.n9118 VSS.n1524 0.0886356
R9779 VSS.n9115 VSS.n1524 0.0886356
R9780 VSS.n969 VSS.n251 0.0886356
R9781 VSS.n279 VSS.n251 0.0886356
R9782 VSS.n10285 VSS.n10284 0.0886356
R9783 VSS.n10286 VSS.n10285 0.0886356
R9784 VSS.n10248 VSS.n276 0.0886356
R9785 VSS.n281 VSS.n276 0.0886356
R9786 VSS.n985 VSS.n277 0.0886356
R9787 VSS.n10245 VSS.n277 0.0886356
R9788 VSS.n10248 VSS.n10247 0.0886356
R9789 VSS.n10247 VSS.n10246 0.0886356
R9790 VSS.n10242 VSS.n10241 0.0886356
R9791 VSS.n10243 VSS.n10242 0.0886356
R9792 VSS.n1006 VSS.n289 0.0886356
R9793 VSS.n320 VSS.n289 0.0886356
R9794 VSS.n10241 VSS.n10240 0.0886356
R9795 VSS.n10240 VSS.n282 0.0886356
R9796 VSS.n10234 VSS.n290 0.0886356
R9797 VSS.n10237 VSS.n290 0.0886356
R9798 VSS.n10235 VSS.n10234 0.0886356
R9799 VSS.n10236 VSS.n10235 0.0886356
R9800 VSS.n1018 VSS.n321 0.0886356
R9801 VSS.n351 VSS.n321 0.0886356
R9802 VSS.n10188 VSS.n348 0.0886356
R9803 VSS.n353 VSS.n348 0.0886356
R9804 VSS.n1043 VSS.n349 0.0886356
R9805 VSS.n10185 VSS.n349 0.0886356
R9806 VSS.n10188 VSS.n10187 0.0886356
R9807 VSS.n10187 VSS.n10186 0.0886356
R9808 VSS.n10182 VSS.n10181 0.0886356
R9809 VSS.n10183 VSS.n10182 0.0886356
R9810 VSS.n1055 VSS.n361 0.0886356
R9811 VSS.n392 VSS.n361 0.0886356
R9812 VSS.n10181 VSS.n10180 0.0886356
R9813 VSS.n10180 VSS.n354 0.0886356
R9814 VSS.n10174 VSS.n362 0.0886356
R9815 VSS.n10177 VSS.n362 0.0886356
R9816 VSS.n10175 VSS.n10174 0.0886356
R9817 VSS.n10176 VSS.n10175 0.0886356
R9818 VSS.n1076 VSS.n393 0.0886356
R9819 VSS.n9301 VSS.n393 0.0886356
R9820 VSS.n10128 VSS.n420 0.0886356
R9821 VSS.n423 VSS.n420 0.0886356
R9822 VSS.n1092 VSS.n421 0.0886356
R9823 VSS.n10125 VSS.n421 0.0886356
R9824 VSS.n10128 VSS.n10127 0.0886356
R9825 VSS.n10127 VSS.n10126 0.0886356
R9826 VSS.n10122 VSS.n10121 0.0886356
R9827 VSS.n10123 VSS.n10122 0.0886356
R9828 VSS.n10121 VSS.n10120 0.0886356
R9829 VSS.n10120 VSS.n424 0.0886356
R9830 VSS.n9365 VSS.n1482 0.0886356
R9831 VSS.n1499 VSS.n1482 0.0886356
R9832 VSS.n9349 VSS.n9348 0.0886356
R9833 VSS.n9348 VSS.n9347 0.0886356
R9834 VSS.n9365 VSS.n1384 0.0886356
R9835 VSS.n1498 VSS.n1384 0.0886356
R9836 VSS.n9401 VSS.n1395 0.0886356
R9837 VSS.n1395 VSS.n1394 0.0886356
R9838 VSS.n9421 VSS.n9420 0.0886356
R9839 VSS.n9422 VSS.n9421 0.0886356
R9840 VSS.n9401 VSS.n1222 0.0886356
R9841 VSS.n1393 VSS.n1222 0.0886356
R9842 VSS.n9527 VSS.n1232 0.0886356
R9843 VSS.n9527 VSS.n9526 0.0886356
R9844 VSS.n9529 VSS.n9528 0.0886356
R9845 VSS.n9528 VSS.n434 0.0886356
R9846 VSS.n1232 VSS.n831 0.0886356
R9847 VSS.n9525 VSS.n831 0.0886356
R9848 VSS.n9558 VSS.n832 0.0886356
R9849 VSS.n9561 VSS.n832 0.0886356
R9850 VSS.n9542 VSS.n9541 0.0886356
R9851 VSS.n9541 VSS.n833 0.0886356
R9852 VSS.n9559 VSS.n9558 0.0886356
R9853 VSS.n9560 VSS.n9559 0.0886356
R9854 VSS.n1186 VSS.n1185 0.0886356
R9855 VSS.n1185 VSS.n1184 0.0886356
R9856 VSS.n1205 VSS.n1153 0.0886356
R9857 VSS.n1153 VSS.n506 0.0886356
R9858 VSS.n1186 VSS.n215 0.0886356
R9859 VSS.n1183 VSS.n215 0.0886356
R9860 VSS.n718 VSS.n216 0.0886356
R9861 VSS.n566 VSS.n216 0.0886356
R9862 VSS.n10931 VSS.n10930 0.0886356
R9863 VSS.n10930 VSS.n10929 0.0886356
R9864 VSS.n718 VSS.n179 0.0886356
R9865 VSS.n565 VSS.n179 0.0886356
R9866 VSS.n10961 VSS.n180 0.0886356
R9867 VSS.n180 VSS.n148 0.0886356
R9868 VSS.n10981 VSS.n10980 0.0886356
R9869 VSS.n10982 VSS.n10981 0.0886356
R9870 VSS.n10961 VSS.n91 0.0886356
R9871 VSS.n11279 VSS.n91 0.0886356
R9872 VSS.n11216 VSS.n92 0.0886356
R9873 VSS.n11288 VSS.n92 0.0886356
R9874 VSS.n11363 VSS.n11362 0.0886356
R9875 VSS.n11362 VSS.n11361 0.0886356
R9876 VSS.n11216 VSS.n4 0.0886356
R9877 VSS.n11287 VSS.n4 0.0886356
R9878 VSS.n70 VSS.n5 0.0886356
R9879 VSS.n11298 VSS.n5 0.0886356
R9880 VSS.n11376 VSS.n11375 0.0886356
R9881 VSS.n11375 VSS.n6 0.0886356
R9882 VSS.n1113 VSS.n431 0.0886356
R9883 VSS.n434 VSS.n431 0.0886356
R9884 VSS.n891 VSS.n432 0.0886356
R9885 VSS.n9526 VSS.n432 0.0886356
R9886 VSS.n1125 VSS.n835 0.0886356
R9887 VSS.n835 VSS.n833 0.0886356
R9888 VSS.n891 VSS.n834 0.0886356
R9889 VSS.n9525 VSS.n834 0.0886356
R9890 VSS.n9562 VSS.n1152 0.0886356
R9891 VSS.n9562 VSS.n9561 0.0886356
R9892 VSS.n868 VSS.n867 0.0886356
R9893 VSS.n867 VSS.n506 0.0886356
R9894 VSS.n1152 VSS.n504 0.0886356
R9895 VSS.n9560 VSS.n504 0.0886356
R9896 VSS.n851 VSS.n505 0.0886356
R9897 VSS.n1184 VSS.n505 0.0886356
R9898 VSS.n10928 VSS.n10927 0.0886356
R9899 VSS.n10929 VSS.n10928 0.0886356
R9900 VSS.n851 VSS.n219 0.0886356
R9901 VSS.n1183 VSS.n219 0.0886356
R9902 VSS.n10902 VSS.n220 0.0886356
R9903 VSS.n566 VSS.n220 0.0886356
R9904 VSS.n10984 VSS.n10983 0.0886356
R9905 VSS.n10983 VSS.n10982 0.0886356
R9906 VSS.n10902 VSS.n182 0.0886356
R9907 VSS.n565 VSS.n182 0.0886356
R9908 VSS.n11012 VSS.n183 0.0886356
R9909 VSS.n183 VSS.n148 0.0886356
R9910 VSS.n11360 VSS.n11359 0.0886356
R9911 VSS.n11361 VSS.n11360 0.0886356
R9912 VSS.n11012 VSS.n94 0.0886356
R9913 VSS.n11279 VSS.n94 0.0886356
R9914 VSS.n11069 VSS.n95 0.0886356
R9915 VSS.n11288 VSS.n95 0.0886356
R9916 VSS.n11347 VSS.n11346 0.0886356
R9917 VSS.n11346 VSS.n6 0.0886356
R9918 VSS.n11069 VSS.n7 0.0886356
R9919 VSS.n11287 VSS.n7 0.0886356
R9920 VSS.n11330 VSS.n8 0.0886356
R9921 VSS.n11298 VSS.n8 0.0886356
R9922 VSS.n9182 VSS.n9181 0.0871667
R9923 VSS.n9181 VSS.n9180 0.0871667
R9924 VSS.n9247 VSS.n9246 0.0871667
R9925 VSS.n9248 VSS.n9247 0.0871667
R9926 VSS.n9309 VSS.n9308 0.0871667
R9927 VSS.n9308 VSS.n9307 0.0871667
R9928 VSS.n9015 VSS.n9014 0.0871667
R9929 VSS.n9014 VSS.n9013 0.0871667
R9930 VSS.n9090 VSS.n9089 0.0871667
R9931 VSS.n9091 VSS.n9090 0.0871667
R9932 VSS.n9068 VSS.n1531 0.0871667
R9933 VSS.n9114 VSS.n1531 0.0871667
R9934 VSS.n10272 VSS.n252 0.0871667
R9935 VSS.n280 VSS.n252 0.0871667
R9936 VSS.n307 VSS.n278 0.0871667
R9937 VSS.n10244 VSS.n278 0.0871667
R9938 VSS.n10239 VSS.n319 0.0871667
R9939 VSS.n10239 VSS.n10238 0.0871667
R9940 VSS.n10212 VSS.n322 0.0871667
R9941 VSS.n352 VSS.n322 0.0871667
R9942 VSS.n370 VSS.n350 0.0871667
R9943 VSS.n10184 VSS.n350 0.0871667
R9944 VSS.n10179 VSS.n391 0.0871667
R9945 VSS.n10179 VSS.n10178 0.0871667
R9946 VSS.n10152 VSS.n394 0.0871667
R9947 VSS.n9300 VSS.n394 0.0871667
R9948 VSS.n1289 VSS.n422 0.0871667
R9949 VSS.n10124 VSS.n422 0.0871667
R9950 VSS.n9345 VSS.n9344 0.0871667
R9951 VSS.n9346 VSS.n9345 0.0871667
R9952 VSS.n9382 VSS.n9381 0.0871667
R9953 VSS.n9381 VSS.n1383 0.0871667
R9954 VSS.n1421 VSS.n435 0.0871667
R9955 VSS.n10118 VSS.n435 0.0871667
R9956 VSS.n9566 VSS.n9565 0.0871667
R9957 VSS.n9565 VSS.n9564 0.0871667
R9958 VSS.n9800 VSS.n507 0.0871667
R9959 VSS.n10067 VSS.n507 0.0871667
R9960 VSS.n694 VSS.n693 0.0871667
R9961 VSS.n693 VSS.n218 0.0871667
R9962 VSS.n11154 VSS.n11153 0.0871667
R9963 VSS.n11153 VSS.n11152 0.0871667
R9964 VSS.n11264 VSS.n11263 0.0871667
R9965 VSS.n11263 VSS.n93 0.0871667
R9966 VSS.n11470 VSS.n11469 0.0871667
R9967 VSS.n11469 VSS.n11468 0.0871667
R9968 VSS.n10119 VSS.n433 0.0871667
R9969 VSS.n10119 VSS.n10118 0.0871667
R9970 VSS.n9563 VSS.n458 0.0871667
R9971 VSS.n9564 VSS.n9563 0.0871667
R9972 VSS.n10069 VSS.n10068 0.0871667
R9973 VSS.n10068 VSS.n10067 0.0871667
R9974 VSS.n548 VSS.n547 0.0871667
R9975 VSS.n547 VSS.n218 0.0871667
R9976 VSS.n11151 VSS.n11150 0.0871667
R9977 VSS.n11152 VSS.n11151 0.0871667
R9978 VSS.n11038 VSS.n11037 0.0871667
R9979 VSS.n11037 VSS.n93 0.0871667
R9980 VSS.n11467 VSS.n11466 0.0871667
R9981 VSS.n11468 VSS.n11467 0.0871667
R9982 VSS.n1349 VSS.n438 0.08175
R9983 VSS.n10117 VSS.n438 0.08175
R9984 VSS.n1426 VSS.n437 0.08175
R9985 VSS.n10117 VSS.n437 0.08175
R9986 VSS.n9765 VSS.n9764 0.08175
R9987 VSS.n9766 VSS.n9765 0.08175
R9988 VSS.n9768 VSS.n9767 0.08175
R9989 VSS.n9767 VSS.n9766 0.08175
R9990 VSS.n9666 VSS.n510 0.08175
R9991 VSS.n10066 VSS.n510 0.08175
R9992 VSS.n9816 VSS.n509 0.08175
R9993 VSS.n10066 VSS.n509 0.08175
R9994 VSS.n10031 VSS.n10030 0.08175
R9995 VSS.n10032 VSS.n10031 0.08175
R9996 VSS.n750 VSS.n564 0.08175
R9997 VSS.n10032 VSS.n564 0.08175
R9998 VSS.n149 VSS.n147 0.08175
R9999 VSS.n11279 VSS.n149 0.08175
R10000 VSS.n11278 VSS.n11277 0.08175
R10001 VSS.n11279 VSS.n11278 0.08175
R10002 VSS.n11291 VSS.n138 0.08175
R10003 VSS.n11292 VSS.n11291 0.08175
R10004 VSS.n11226 VSS.n139 0.08175
R10005 VSS.n11292 VSS.n139 0.08175
R10006 VSS.n10116 VSS.n10115 0.08175
R10007 VSS.n10117 VSS.n10116 0.08175
R10008 VSS.n1349 VSS.n436 0.08175
R10009 VSS.n10117 VSS.n436 0.08175
R10010 VSS.n644 VSS.n487 0.08175
R10011 VSS.n9766 VSS.n644 0.08175
R10012 VSS.n9764 VSS.n645 0.08175
R10013 VSS.n9766 VSS.n645 0.08175
R10014 VSS.n10065 VSS.n10064 0.08175
R10015 VSS.n10066 VSS.n10065 0.08175
R10016 VSS.n9666 VSS.n508 0.08175
R10017 VSS.n10066 VSS.n508 0.08175
R10018 VSS.n10034 VSS.n10033 0.08175
R10019 VSS.n10033 VSS.n10032 0.08175
R10020 VSS.n10030 VSS.n563 0.08175
R10021 VSS.n10032 VSS.n563 0.08175
R10022 VSS.n11023 VSS.n145 0.08175
R10023 VSS.n11279 VSS.n145 0.08175
R10024 VSS.n11280 VSS.n147 0.08175
R10025 VSS.n11280 VSS.n11279 0.08175
R10026 VSS.n11081 VSS.n136 0.08175
R10027 VSS.n11292 VSS.n136 0.08175
R10028 VSS.n11293 VSS.n138 0.08175
R10029 VSS.n11293 VSS.n11292 0.08175
R10030 VSS.n10695 VSS.n10694 0.0769706
R10031 VSS.n10696 VSS.n10695 0.0769706
R10032 VSS.n10598 VSS.n10597 0.0769706
R10033 VSS.n10599 VSS.n10598 0.0769706
R10034 VSS.n10661 VSS.n10660 0.0769706
R10035 VSS.n10662 VSS.n10661 0.0769706
R10036 VSS.n10604 VSS.n10603 0.0769706
R10037 VSS.n10603 VSS.n10602 0.0769706
R10038 VSS.n10441 VSS.n10340 0.0769706
R10039 VSS.n10601 VSS.n10340 0.0769706
R10040 VSS.n10341 VSS.n240 0.0769706
R10041 VSS.n10341 VSS.n244 0.0769706
R10042 VSS.n10720 VSS.n131 0.0769706
R10043 VSS.n11300 VSS.n131 0.0769706
R10044 VSS.n10831 VSS.n130 0.0769706
R10045 VSS.n10848 VSS.n130 0.0769706
R10046 VSS.n10597 VSS.n10596 0.072814
R10047 VSS.n10694 VSS.n10693 0.072814
R10048 VSS.n9433 VSS.n9429 0.069264
R10049 VSS.n9431 VSS.n9429 0.069264
R10050 VSS.n9431 VSS.n9430 0.069264
R10051 VSS.n9430 VSS.n1380 0.069264
R10052 VSS.n9470 VSS.n9469 0.069264
R10053 VSS.n9471 VSS.n9470 0.069264
R10054 VSS.n9471 VSS.n1378 0.069264
R10055 VSS.n9473 VSS.n1378 0.069264
R10056 VSS.n10822 VSS.n129 0.0686515
R10057 VSS.n10842 VSS.n10698 0.0686515
R10058 VSS.n9449 VSS.n9448 0.0685756
R10059 VSS.n9450 VSS.n9449 0.0685756
R10060 VSS.n9450 VSS.n9423 0.0685756
R10061 VSS.n9452 VSS.n9423 0.0685756
R10062 VSS.n9458 VSS.n9453 0.0685756
R10063 VSS.n9456 VSS.n9453 0.0685756
R10064 VSS.n9456 VSS.n9455 0.0685756
R10065 VSS.n9455 VSS.n9454 0.0685756
R10066 VSS.n10660 VSS.n10345 0.0681047
R10067 VSS.n10660 VSS.n10659 0.0678953
R10068 VSS.n10844 VSS.n10843 0.0678497
R10069 VSS.n10586 VSS.n10288 0.0646975
R10070 VSS.n10442 VSS.n10288 0.0646975
R10071 VSS.n10464 VSS.n10343 0.0646975
R10072 VSS.n10600 VSS.n10343 0.0646975
R10073 VSS.n10665 VSS.n10664 0.0646975
R10074 VSS.n10664 VSS.n10663 0.0646975
R10075 VSS.n10428 VSS.n10289 0.0646975
R10076 VSS.n10442 VSS.n10289 0.0646975
R10077 VSS.n10349 VSS.n10342 0.0646975
R10078 VSS.n10663 VSS.n10342 0.0646975
R10079 VSS.n10531 VSS.n10344 0.0646975
R10080 VSS.n10600 VSS.n10344 0.0646975
R10081 VSS.n11304 VSS.n11303 0.0640412
R10082 VSS.n10597 VSS.n10481 0.063186
R10083 VSS.n10694 VSS.n10290 0.063186
R10084 VSS.n10841 VSS.n10734 0.0583997
R10085 VSS.n10609 VSS.n10608 0.0533671
R10086 VSS.n9464 VSS.n9463 0.0519852
R10087 VSS.n9465 VSS.n9464 0.0519852
R10088 VSS.n9467 VSS.n9466 0.0519852
R10089 VSS.n9466 VSS.n9465 0.0519852
R10090 VSS.n10534 VSS.n10497 0.0513741
R10091 VSS.n1389 VSS.n1388 0.0490981
R10092 VSS.n1390 VSS.n1389 0.0490981
R10093 VSS.n1235 VSS.n1234 0.0490981
R10094 VSS.n9524 VSS.n1235 0.0490981
R10095 VSS.n1234 VSS.n797 0.0490981
R10096 VSS.n9523 VSS.n797 0.0490981
R10097 VSS.n9887 VSS.n646 0.0490981
R10098 VSS.n9890 VSS.n646 0.0490981
R10099 VSS.n9888 VSS.n9887 0.0490981
R10100 VSS.n9889 VSS.n9888 0.0490981
R10101 VSS.n1181 VSS.n1180 0.0490981
R10102 VSS.n1182 VSS.n1181 0.0490981
R10103 VSS.n1176 VSS.n567 0.0490981
R10104 VSS.n567 VSS.n217 0.0490981
R10105 VSS.n671 VSS.n568 0.0490981
R10106 VSS.n568 VSS.n208 0.0490981
R10107 VSS.n671 VSS.n150 0.0490981
R10108 VSS.n181 VSS.n150 0.0490981
R10109 VSS.n144 VSS.n143 0.0490981
R10110 VSS.n11286 VSS.n144 0.0490981
R10111 VSS.n11290 VSS.n143 0.0490981
R10112 VSS.n11290 VSS.n11289 0.0490981
R10113 VSS.n135 VSS.n134 0.0490981
R10114 VSS.n11297 VSS.n135 0.0490981
R10115 VSS.n1330 VSS.n439 0.0490981
R10116 VSS.n1390 VSS.n439 0.0490981
R10117 VSS.n9521 VSS.n440 0.0490981
R10118 VSS.n9524 VSS.n440 0.0490981
R10119 VSS.n9522 VSS.n9521 0.0490981
R10120 VSS.n9523 VSS.n9522 0.0490981
R10121 VSS.n9892 VSS.n9891 0.0490981
R10122 VSS.n9891 VSS.n9890 0.0490981
R10123 VSS.n9892 VSS.n511 0.0490981
R10124 VSS.n9889 VSS.n511 0.0490981
R10125 VSS.n626 VSS.n512 0.0490981
R10126 VSS.n1182 VSS.n512 0.0490981
R10127 VSS.n623 VSS.n561 0.0490981
R10128 VSS.n561 VSS.n217 0.0490981
R10129 VSS.n9916 VSS.n562 0.0490981
R10130 VSS.n562 VSS.n208 0.0490981
R10131 VSS.n9916 VSS.n146 0.0490981
R10132 VSS.n181 VSS.n146 0.0490981
R10133 VSS.n11285 VSS.n11284 0.0490981
R10134 VSS.n11286 VSS.n11285 0.0490981
R10135 VSS.n11284 VSS.n137 0.0490981
R10136 VSS.n11289 VSS.n137 0.0490981
R10137 VSS.n11296 VSS.n11295 0.0490981
R10138 VSS.n11297 VSS.n11296 0.0490981
R10139 VSS.n9475 VSS.n9473 0.0456011
R10140 VSS.n9454 VSS.n1336 0.0451496
R10141 VSS.n10764 VSS.n10763 0.0431396
R10142 VSS.n10766 VSS.n10738 0.0431396
R10143 VSS.n10768 VSS.n10738 0.0431396
R10144 VSS.n10765 VSS.n10764 0.0420736
R10145 VSS.n1319 VSS.n1318 0.0414574
R10146 VSS.n10450 VSS.n10449 0.041314
R10147 VSS.n10480 VSS.n10479 0.041314
R10148 VSS.n10559 VSS.n10558 0.041314
R10149 VSS.n1416 VSS.n1415 0.0412447
R10150 VSS.n10658 VSS.n10657 0.0411047
R10151 VSS.n10595 VSS.n10594 0.0411047
R10152 VSS.n10692 VSS.n10691 0.0411047
R10153 VSS.n5469 VSS.n2742 0.04025
R10154 VSS.n5473 VSS.n2742 0.04025
R10155 VSS.n5474 VSS.n5473 0.04025
R10156 VSS.n5475 VSS.n5474 0.04025
R10157 VSS.n5475 VSS.n2740 0.04025
R10158 VSS.n5479 VSS.n2740 0.04025
R10159 VSS.n5480 VSS.n5479 0.04025
R10160 VSS.n5481 VSS.n5480 0.04025
R10161 VSS.n5481 VSS.n2738 0.04025
R10162 VSS.n5485 VSS.n2738 0.04025
R10163 VSS.n5486 VSS.n5485 0.04025
R10164 VSS.n5487 VSS.n5486 0.04025
R10165 VSS.n5487 VSS.n2736 0.04025
R10166 VSS.n5491 VSS.n2736 0.04025
R10167 VSS.n5492 VSS.n5491 0.04025
R10168 VSS.n5493 VSS.n5492 0.04025
R10169 VSS.n5493 VSS.n2734 0.04025
R10170 VSS.n5497 VSS.n2734 0.04025
R10171 VSS.n5498 VSS.n5497 0.04025
R10172 VSS.n5499 VSS.n5498 0.04025
R10173 VSS.n5499 VSS.n2732 0.04025
R10174 VSS.n5503 VSS.n2732 0.04025
R10175 VSS.n5504 VSS.n5503 0.04025
R10176 VSS.n5505 VSS.n5504 0.04025
R10177 VSS.n5505 VSS.n2730 0.04025
R10178 VSS.n5509 VSS.n2730 0.04025
R10179 VSS.n5510 VSS.n5509 0.04025
R10180 VSS.n5511 VSS.n5510 0.04025
R10181 VSS.n5511 VSS.n2728 0.04025
R10182 VSS.n5515 VSS.n2728 0.04025
R10183 VSS.n5516 VSS.n5515 0.04025
R10184 VSS.n5517 VSS.n5516 0.04025
R10185 VSS.n5517 VSS.n2726 0.04025
R10186 VSS.n5521 VSS.n2726 0.04025
R10187 VSS.n5522 VSS.n5521 0.04025
R10188 VSS.n5523 VSS.n5522 0.04025
R10189 VSS.n5523 VSS.n2724 0.04025
R10190 VSS.n5527 VSS.n2724 0.04025
R10191 VSS.n5528 VSS.n5527 0.04025
R10192 VSS.n5529 VSS.n5528 0.04025
R10193 VSS.n5529 VSS.n2722 0.04025
R10194 VSS.n5533 VSS.n2722 0.04025
R10195 VSS.n5534 VSS.n5533 0.04025
R10196 VSS.n5535 VSS.n5534 0.04025
R10197 VSS.n5535 VSS.n2720 0.04025
R10198 VSS.n5539 VSS.n2720 0.04025
R10199 VSS.n5540 VSS.n5539 0.04025
R10200 VSS.n5541 VSS.n5540 0.04025
R10201 VSS.n5541 VSS.n2718 0.04025
R10202 VSS.n5545 VSS.n2718 0.04025
R10203 VSS.n5546 VSS.n5545 0.04025
R10204 VSS.n5547 VSS.n5546 0.04025
R10205 VSS.n5547 VSS.n2716 0.04025
R10206 VSS.n5551 VSS.n2716 0.04025
R10207 VSS.n5552 VSS.n5551 0.04025
R10208 VSS.n5553 VSS.n5552 0.04025
R10209 VSS.n5553 VSS.n2714 0.04025
R10210 VSS.n5557 VSS.n2714 0.04025
R10211 VSS.n5558 VSS.n5557 0.04025
R10212 VSS.n5559 VSS.n5558 0.04025
R10213 VSS.n5559 VSS.n2712 0.04025
R10214 VSS.n5563 VSS.n2712 0.04025
R10215 VSS.n5564 VSS.n5563 0.04025
R10216 VSS.n5565 VSS.n5564 0.04025
R10217 VSS.n5565 VSS.n2710 0.04025
R10218 VSS.n5569 VSS.n2710 0.04025
R10219 VSS.n5570 VSS.n5569 0.04025
R10220 VSS.n5571 VSS.n5570 0.04025
R10221 VSS.n5571 VSS.n2708 0.04025
R10222 VSS.n5575 VSS.n2708 0.04025
R10223 VSS.n5576 VSS.n5575 0.04025
R10224 VSS.n5577 VSS.n5576 0.04025
R10225 VSS.n5577 VSS.n2706 0.04025
R10226 VSS.n5581 VSS.n2706 0.04025
R10227 VSS.n5582 VSS.n5581 0.04025
R10228 VSS.n5583 VSS.n5582 0.04025
R10229 VSS.n5583 VSS.n2704 0.04025
R10230 VSS.n5587 VSS.n2704 0.04025
R10231 VSS.n5588 VSS.n5587 0.04025
R10232 VSS.n5589 VSS.n5588 0.04025
R10233 VSS.n5589 VSS.n2702 0.04025
R10234 VSS.n5593 VSS.n2702 0.04025
R10235 VSS.n5594 VSS.n5593 0.04025
R10236 VSS.n5595 VSS.n5594 0.04025
R10237 VSS.n5595 VSS.n2700 0.04025
R10238 VSS.n5599 VSS.n2700 0.04025
R10239 VSS.n5600 VSS.n5599 0.04025
R10240 VSS.n5601 VSS.n5600 0.04025
R10241 VSS.n5601 VSS.n2698 0.04025
R10242 VSS.n5605 VSS.n2698 0.04025
R10243 VSS.n5606 VSS.n5605 0.04025
R10244 VSS.n5607 VSS.n5606 0.04025
R10245 VSS.n5607 VSS.n2696 0.04025
R10246 VSS.n5611 VSS.n2696 0.04025
R10247 VSS.n5612 VSS.n5611 0.04025
R10248 VSS.n5613 VSS.n5612 0.04025
R10249 VSS.n5613 VSS.n2694 0.04025
R10250 VSS.n5617 VSS.n2694 0.04025
R10251 VSS.n5618 VSS.n5617 0.04025
R10252 VSS.n5619 VSS.n5618 0.04025
R10253 VSS.n5619 VSS.n2692 0.04025
R10254 VSS.n5623 VSS.n2692 0.04025
R10255 VSS.n5624 VSS.n5623 0.04025
R10256 VSS.n5625 VSS.n5624 0.04025
R10257 VSS.n5625 VSS.n2690 0.04025
R10258 VSS.n5629 VSS.n2690 0.04025
R10259 VSS.n5630 VSS.n5629 0.04025
R10260 VSS.n5631 VSS.n5630 0.04025
R10261 VSS.n5631 VSS.n2688 0.04025
R10262 VSS.n5635 VSS.n2688 0.04025
R10263 VSS.n5636 VSS.n5635 0.04025
R10264 VSS.n5637 VSS.n5636 0.04025
R10265 VSS.n5637 VSS.n2686 0.04025
R10266 VSS.n5641 VSS.n2686 0.04025
R10267 VSS.n5642 VSS.n5641 0.04025
R10268 VSS.n5643 VSS.n5642 0.04025
R10269 VSS.n5643 VSS.n2684 0.04025
R10270 VSS.n5647 VSS.n2684 0.04025
R10271 VSS.n5648 VSS.n5647 0.04025
R10272 VSS.n5649 VSS.n5648 0.04025
R10273 VSS.n5649 VSS.n2682 0.04025
R10274 VSS.n5653 VSS.n2682 0.04025
R10275 VSS.n5654 VSS.n5653 0.04025
R10276 VSS.n5655 VSS.n5654 0.04025
R10277 VSS.n5655 VSS.n2680 0.04025
R10278 VSS.n5659 VSS.n2680 0.04025
R10279 VSS.n5660 VSS.n5659 0.04025
R10280 VSS.n5661 VSS.n5660 0.04025
R10281 VSS.n5661 VSS.n2678 0.04025
R10282 VSS.n5665 VSS.n2678 0.04025
R10283 VSS.n5666 VSS.n5665 0.04025
R10284 VSS.n5667 VSS.n5666 0.04025
R10285 VSS.n5667 VSS.n2676 0.04025
R10286 VSS.n5671 VSS.n2676 0.04025
R10287 VSS.n5672 VSS.n5671 0.04025
R10288 VSS.n5673 VSS.n5672 0.04025
R10289 VSS.n5673 VSS.n2674 0.04025
R10290 VSS.n5677 VSS.n2674 0.04025
R10291 VSS.n5678 VSS.n5677 0.04025
R10292 VSS.n5679 VSS.n5678 0.04025
R10293 VSS.n5679 VSS.n2672 0.04025
R10294 VSS.n5683 VSS.n2672 0.04025
R10295 VSS.n5684 VSS.n5683 0.04025
R10296 VSS.n5685 VSS.n5684 0.04025
R10297 VSS.n5685 VSS.n2670 0.04025
R10298 VSS.n5689 VSS.n2670 0.04025
R10299 VSS.n5690 VSS.n5689 0.04025
R10300 VSS.n5691 VSS.n5690 0.04025
R10301 VSS.n5691 VSS.n2668 0.04025
R10302 VSS.n5695 VSS.n2668 0.04025
R10303 VSS.n5696 VSS.n5695 0.04025
R10304 VSS.n5697 VSS.n5696 0.04025
R10305 VSS.n5697 VSS.n2666 0.04025
R10306 VSS.n5701 VSS.n2666 0.04025
R10307 VSS.n5702 VSS.n5701 0.04025
R10308 VSS.n5703 VSS.n5702 0.04025
R10309 VSS.n5703 VSS.n2664 0.04025
R10310 VSS.n5707 VSS.n2664 0.04025
R10311 VSS.n5708 VSS.n5707 0.04025
R10312 VSS.n5709 VSS.n5708 0.04025
R10313 VSS.n5709 VSS.n2662 0.04025
R10314 VSS.n5713 VSS.n2662 0.04025
R10315 VSS.n5714 VSS.n5713 0.04025
R10316 VSS.n5715 VSS.n5714 0.04025
R10317 VSS.n5715 VSS.n2660 0.04025
R10318 VSS.n5719 VSS.n2660 0.04025
R10319 VSS.n5720 VSS.n5719 0.04025
R10320 VSS.n5721 VSS.n5720 0.04025
R10321 VSS.n5721 VSS.n2658 0.04025
R10322 VSS.n5725 VSS.n2658 0.04025
R10323 VSS.n5726 VSS.n5725 0.04025
R10324 VSS.n5727 VSS.n5726 0.04025
R10325 VSS.n5727 VSS.n2656 0.04025
R10326 VSS.n5731 VSS.n2656 0.04025
R10327 VSS.n5732 VSS.n5731 0.04025
R10328 VSS.n5733 VSS.n5732 0.04025
R10329 VSS.n5733 VSS.n2654 0.04025
R10330 VSS.n5737 VSS.n2654 0.04025
R10331 VSS.n5738 VSS.n5737 0.04025
R10332 VSS.n5739 VSS.n5738 0.04025
R10333 VSS.n5739 VSS.n2652 0.04025
R10334 VSS.n5743 VSS.n2652 0.04025
R10335 VSS.n5744 VSS.n5743 0.04025
R10336 VSS.n5745 VSS.n5744 0.04025
R10337 VSS.n5745 VSS.n2650 0.04025
R10338 VSS.n5749 VSS.n2650 0.04025
R10339 VSS.n5750 VSS.n5749 0.04025
R10340 VSS.n5751 VSS.n5750 0.04025
R10341 VSS.n5751 VSS.n2648 0.04025
R10342 VSS.n5755 VSS.n2648 0.04025
R10343 VSS.n5756 VSS.n5755 0.04025
R10344 VSS.n5757 VSS.n5756 0.04025
R10345 VSS.n5757 VSS.n2646 0.04025
R10346 VSS.n5761 VSS.n2646 0.04025
R10347 VSS.n5762 VSS.n5761 0.04025
R10348 VSS.n5763 VSS.n5762 0.04025
R10349 VSS.n5763 VSS.n2644 0.04025
R10350 VSS.n5767 VSS.n2644 0.04025
R10351 VSS.n5768 VSS.n5767 0.04025
R10352 VSS.n5769 VSS.n5768 0.04025
R10353 VSS.n5769 VSS.n2642 0.04025
R10354 VSS.n5773 VSS.n2642 0.04025
R10355 VSS.n5774 VSS.n5773 0.04025
R10356 VSS.n5775 VSS.n5774 0.04025
R10357 VSS.n5775 VSS.n2640 0.04025
R10358 VSS.n5779 VSS.n2640 0.04025
R10359 VSS.n5780 VSS.n5779 0.04025
R10360 VSS.n5781 VSS.n5780 0.04025
R10361 VSS.n5781 VSS.n2638 0.04025
R10362 VSS.n5785 VSS.n2638 0.04025
R10363 VSS.n5786 VSS.n5785 0.04025
R10364 VSS.n5787 VSS.n5786 0.04025
R10365 VSS.n5787 VSS.n2636 0.04025
R10366 VSS.n5791 VSS.n2636 0.04025
R10367 VSS.n5792 VSS.n5791 0.04025
R10368 VSS.n5793 VSS.n5792 0.04025
R10369 VSS.n5793 VSS.n2634 0.04025
R10370 VSS.n5797 VSS.n2634 0.04025
R10371 VSS.n5798 VSS.n5797 0.04025
R10372 VSS.n5799 VSS.n5798 0.04025
R10373 VSS.n5799 VSS.n2632 0.04025
R10374 VSS.n5803 VSS.n2632 0.04025
R10375 VSS.n5804 VSS.n5803 0.04025
R10376 VSS.n5805 VSS.n5804 0.04025
R10377 VSS.n5805 VSS.n2630 0.04025
R10378 VSS.n5809 VSS.n2630 0.04025
R10379 VSS.n5810 VSS.n5809 0.04025
R10380 VSS.n5811 VSS.n5810 0.04025
R10381 VSS.n5811 VSS.n2628 0.04025
R10382 VSS.n5815 VSS.n2628 0.04025
R10383 VSS.n5816 VSS.n5815 0.04025
R10384 VSS.n5817 VSS.n5816 0.04025
R10385 VSS.n5817 VSS.n2626 0.04025
R10386 VSS.n5821 VSS.n2626 0.04025
R10387 VSS.n5822 VSS.n5821 0.04025
R10388 VSS.n5823 VSS.n5822 0.04025
R10389 VSS.n5823 VSS.n2624 0.04025
R10390 VSS.n5827 VSS.n2624 0.04025
R10391 VSS.n5828 VSS.n5827 0.04025
R10392 VSS.n5829 VSS.n5828 0.04025
R10393 VSS.n5829 VSS.n2622 0.04025
R10394 VSS.n5833 VSS.n2622 0.04025
R10395 VSS.n5834 VSS.n5833 0.04025
R10396 VSS.n5835 VSS.n5834 0.04025
R10397 VSS.n5835 VSS.n2620 0.04025
R10398 VSS.n5839 VSS.n2620 0.04025
R10399 VSS.n5840 VSS.n5839 0.04025
R10400 VSS.n5841 VSS.n5840 0.04025
R10401 VSS.n5841 VSS.n2618 0.04025
R10402 VSS.n5845 VSS.n2618 0.04025
R10403 VSS.n5846 VSS.n5845 0.04025
R10404 VSS.n5847 VSS.n5846 0.04025
R10405 VSS.n5847 VSS.n2616 0.04025
R10406 VSS.n5851 VSS.n2616 0.04025
R10407 VSS.n5852 VSS.n5851 0.04025
R10408 VSS.n5853 VSS.n5852 0.04025
R10409 VSS.n5853 VSS.n2614 0.04025
R10410 VSS.n5857 VSS.n2614 0.04025
R10411 VSS.n5858 VSS.n5857 0.04025
R10412 VSS.n5859 VSS.n5858 0.04025
R10413 VSS.n5859 VSS.n2612 0.04025
R10414 VSS.n5863 VSS.n2612 0.04025
R10415 VSS.n5864 VSS.n5863 0.04025
R10416 VSS.n5865 VSS.n5864 0.04025
R10417 VSS.n5865 VSS.n2610 0.04025
R10418 VSS.n5869 VSS.n2610 0.04025
R10419 VSS.n5870 VSS.n5869 0.04025
R10420 VSS.n5871 VSS.n5870 0.04025
R10421 VSS.n5871 VSS.n2608 0.04025
R10422 VSS.n5875 VSS.n2608 0.04025
R10423 VSS.n5876 VSS.n5875 0.04025
R10424 VSS.n5877 VSS.n5876 0.04025
R10425 VSS.n5877 VSS.n2606 0.04025
R10426 VSS.n5881 VSS.n2606 0.04025
R10427 VSS.n5882 VSS.n5881 0.04025
R10428 VSS.n5883 VSS.n5882 0.04025
R10429 VSS.n5883 VSS.n2604 0.04025
R10430 VSS.n5887 VSS.n2604 0.04025
R10431 VSS.n5888 VSS.n5887 0.04025
R10432 VSS.n5889 VSS.n5888 0.04025
R10433 VSS.n5889 VSS.n2602 0.04025
R10434 VSS.n5893 VSS.n2602 0.04025
R10435 VSS.n5894 VSS.n5893 0.04025
R10436 VSS.n5895 VSS.n5894 0.04025
R10437 VSS.n5895 VSS.n2600 0.04025
R10438 VSS.n5899 VSS.n2600 0.04025
R10439 VSS.n5900 VSS.n5899 0.04025
R10440 VSS.n5901 VSS.n5900 0.04025
R10441 VSS.n5901 VSS.n2598 0.04025
R10442 VSS.n5905 VSS.n2598 0.04025
R10443 VSS.n5906 VSS.n5905 0.04025
R10444 VSS.n5907 VSS.n5906 0.04025
R10445 VSS.n5907 VSS.n2596 0.04025
R10446 VSS.n5911 VSS.n2596 0.04025
R10447 VSS.n5912 VSS.n5911 0.04025
R10448 VSS.n5913 VSS.n5912 0.04025
R10449 VSS.n5913 VSS.n2594 0.04025
R10450 VSS.n5917 VSS.n2594 0.04025
R10451 VSS.n5918 VSS.n5917 0.04025
R10452 VSS.n5919 VSS.n5918 0.04025
R10453 VSS.n5919 VSS.n2592 0.04025
R10454 VSS.n5923 VSS.n2592 0.04025
R10455 VSS.n5924 VSS.n5923 0.04025
R10456 VSS.n5925 VSS.n5924 0.04025
R10457 VSS.n5925 VSS.n2590 0.04025
R10458 VSS.n5929 VSS.n2590 0.04025
R10459 VSS.n5930 VSS.n5929 0.04025
R10460 VSS.n5931 VSS.n5930 0.04025
R10461 VSS.n5931 VSS.n2588 0.04025
R10462 VSS.n5935 VSS.n2588 0.04025
R10463 VSS.n5936 VSS.n5935 0.04025
R10464 VSS.n5937 VSS.n5936 0.04025
R10465 VSS.n5937 VSS.n2586 0.04025
R10466 VSS.n5941 VSS.n2586 0.04025
R10467 VSS.n5942 VSS.n5941 0.04025
R10468 VSS.n5943 VSS.n5942 0.04025
R10469 VSS.n5943 VSS.n2584 0.04025
R10470 VSS.n5947 VSS.n2584 0.04025
R10471 VSS.n5948 VSS.n5947 0.04025
R10472 VSS.n5949 VSS.n5948 0.04025
R10473 VSS.n5949 VSS.n2582 0.04025
R10474 VSS.n5953 VSS.n2582 0.04025
R10475 VSS.n5954 VSS.n5953 0.04025
R10476 VSS.n5955 VSS.n5954 0.04025
R10477 VSS.n5955 VSS.n2580 0.04025
R10478 VSS.n5959 VSS.n2580 0.04025
R10479 VSS.n5960 VSS.n5959 0.04025
R10480 VSS.n5961 VSS.n5960 0.04025
R10481 VSS.n5961 VSS.n2578 0.04025
R10482 VSS.n5965 VSS.n2578 0.04025
R10483 VSS.n5966 VSS.n5965 0.04025
R10484 VSS.n5967 VSS.n5966 0.04025
R10485 VSS.n5967 VSS.n2576 0.04025
R10486 VSS.n5971 VSS.n2576 0.04025
R10487 VSS.n5972 VSS.n5971 0.04025
R10488 VSS.n5973 VSS.n5972 0.04025
R10489 VSS.n5973 VSS.n2574 0.04025
R10490 VSS.n5977 VSS.n2574 0.04025
R10491 VSS.n5978 VSS.n5977 0.04025
R10492 VSS.n5979 VSS.n5978 0.04025
R10493 VSS.n5979 VSS.n2572 0.04025
R10494 VSS.n5983 VSS.n2572 0.04025
R10495 VSS.n5984 VSS.n5983 0.04025
R10496 VSS.n5985 VSS.n5984 0.04025
R10497 VSS.n5985 VSS.n2570 0.04025
R10498 VSS.n5989 VSS.n2570 0.04025
R10499 VSS.n5990 VSS.n5989 0.04025
R10500 VSS.n5991 VSS.n5990 0.04025
R10501 VSS.n5991 VSS.n2568 0.04025
R10502 VSS.n5995 VSS.n2568 0.04025
R10503 VSS.n5996 VSS.n5995 0.04025
R10504 VSS.n5997 VSS.n5996 0.04025
R10505 VSS.n5997 VSS.n2566 0.04025
R10506 VSS.n6001 VSS.n2566 0.04025
R10507 VSS.n6002 VSS.n6001 0.04025
R10508 VSS.n6003 VSS.n6002 0.04025
R10509 VSS.n6003 VSS.n2564 0.04025
R10510 VSS.n6007 VSS.n2564 0.04025
R10511 VSS.n6008 VSS.n6007 0.04025
R10512 VSS.n6009 VSS.n6008 0.04025
R10513 VSS.n6009 VSS.n2562 0.04025
R10514 VSS.n6013 VSS.n2562 0.04025
R10515 VSS.n6014 VSS.n6013 0.04025
R10516 VSS.n6015 VSS.n6014 0.04025
R10517 VSS.n6015 VSS.n2560 0.04025
R10518 VSS.n6019 VSS.n2560 0.04025
R10519 VSS.n6020 VSS.n6019 0.04025
R10520 VSS.n6021 VSS.n6020 0.04025
R10521 VSS.n6021 VSS.n2558 0.04025
R10522 VSS.n6025 VSS.n2558 0.04025
R10523 VSS.n6026 VSS.n6025 0.04025
R10524 VSS.n6027 VSS.n6026 0.04025
R10525 VSS.n6027 VSS.n2556 0.04025
R10526 VSS.n6031 VSS.n2556 0.04025
R10527 VSS.n6032 VSS.n6031 0.04025
R10528 VSS.n6033 VSS.n6032 0.04025
R10529 VSS.n6033 VSS.n2554 0.04025
R10530 VSS.n6037 VSS.n2554 0.04025
R10531 VSS.n6038 VSS.n6037 0.04025
R10532 VSS.n6039 VSS.n6038 0.04025
R10533 VSS.n6039 VSS.n2552 0.04025
R10534 VSS.n6043 VSS.n2552 0.04025
R10535 VSS.n6044 VSS.n6043 0.04025
R10536 VSS.n6045 VSS.n6044 0.04025
R10537 VSS.n6045 VSS.n2550 0.04025
R10538 VSS.n6049 VSS.n2550 0.04025
R10539 VSS.n6050 VSS.n6049 0.04025
R10540 VSS.n6051 VSS.n6050 0.04025
R10541 VSS.n6051 VSS.n2548 0.04025
R10542 VSS.n6055 VSS.n2548 0.04025
R10543 VSS.n6056 VSS.n6055 0.04025
R10544 VSS.n6057 VSS.n6056 0.04025
R10545 VSS.n6057 VSS.n2546 0.04025
R10546 VSS.n6061 VSS.n2546 0.04025
R10547 VSS.n6062 VSS.n6061 0.04025
R10548 VSS.n6063 VSS.n6062 0.04025
R10549 VSS.n6063 VSS.n2544 0.04025
R10550 VSS.n6067 VSS.n2544 0.04025
R10551 VSS.n6068 VSS.n6067 0.04025
R10552 VSS.n6069 VSS.n6068 0.04025
R10553 VSS.n6069 VSS.n2542 0.04025
R10554 VSS.n6073 VSS.n2542 0.04025
R10555 VSS.n6074 VSS.n6073 0.04025
R10556 VSS.n6075 VSS.n6074 0.04025
R10557 VSS.n6075 VSS.n2540 0.04025
R10558 VSS.n6079 VSS.n2540 0.04025
R10559 VSS.n6080 VSS.n6079 0.04025
R10560 VSS.n6081 VSS.n6080 0.04025
R10561 VSS.n6081 VSS.n2538 0.04025
R10562 VSS.n6085 VSS.n2538 0.04025
R10563 VSS.n6086 VSS.n6085 0.04025
R10564 VSS.n6087 VSS.n6086 0.04025
R10565 VSS.n6087 VSS.n2536 0.04025
R10566 VSS.n6091 VSS.n2536 0.04025
R10567 VSS.n6092 VSS.n6091 0.04025
R10568 VSS.n6093 VSS.n6092 0.04025
R10569 VSS.n6093 VSS.n2534 0.04025
R10570 VSS.n6097 VSS.n2534 0.04025
R10571 VSS.n6098 VSS.n6097 0.04025
R10572 VSS.n6099 VSS.n6098 0.04025
R10573 VSS.n6099 VSS.n2532 0.04025
R10574 VSS.n6103 VSS.n2532 0.04025
R10575 VSS.n6104 VSS.n6103 0.04025
R10576 VSS.n6105 VSS.n6104 0.04025
R10577 VSS.n6105 VSS.n2530 0.04025
R10578 VSS.n6109 VSS.n2530 0.04025
R10579 VSS.n6110 VSS.n6109 0.04025
R10580 VSS.n6111 VSS.n6110 0.04025
R10581 VSS.n6111 VSS.n2528 0.04025
R10582 VSS.n6115 VSS.n2528 0.04025
R10583 VSS.n6116 VSS.n6115 0.04025
R10584 VSS.n6117 VSS.n6116 0.04025
R10585 VSS.n6117 VSS.n2526 0.04025
R10586 VSS.n6121 VSS.n2526 0.04025
R10587 VSS.n6122 VSS.n6121 0.04025
R10588 VSS.n6123 VSS.n6122 0.04025
R10589 VSS.n6123 VSS.n2524 0.04025
R10590 VSS.n6127 VSS.n2524 0.04025
R10591 VSS.n6128 VSS.n6127 0.04025
R10592 VSS.n6129 VSS.n6128 0.04025
R10593 VSS.n6129 VSS.n2522 0.04025
R10594 VSS.n6133 VSS.n2522 0.04025
R10595 VSS.n6134 VSS.n6133 0.04025
R10596 VSS.n6135 VSS.n6134 0.04025
R10597 VSS.n6135 VSS.n2520 0.04025
R10598 VSS.n6139 VSS.n2520 0.04025
R10599 VSS.n6140 VSS.n6139 0.04025
R10600 VSS.n6141 VSS.n6140 0.04025
R10601 VSS.n6141 VSS.n2518 0.04025
R10602 VSS.n6145 VSS.n2518 0.04025
R10603 VSS.n6146 VSS.n6145 0.04025
R10604 VSS.n6147 VSS.n6146 0.04025
R10605 VSS.n6147 VSS.n2516 0.04025
R10606 VSS.n6151 VSS.n2516 0.04025
R10607 VSS.n6152 VSS.n6151 0.04025
R10608 VSS.n6153 VSS.n6152 0.04025
R10609 VSS.n6153 VSS.n2514 0.04025
R10610 VSS.n6157 VSS.n2514 0.04025
R10611 VSS.n6158 VSS.n6157 0.04025
R10612 VSS.n6159 VSS.n6158 0.04025
R10613 VSS.n6159 VSS.n2512 0.04025
R10614 VSS.n6163 VSS.n2512 0.04025
R10615 VSS.n6164 VSS.n6163 0.04025
R10616 VSS.n6165 VSS.n6164 0.04025
R10617 VSS.n6165 VSS.n2510 0.04025
R10618 VSS.n6169 VSS.n2510 0.04025
R10619 VSS.n6170 VSS.n6169 0.04025
R10620 VSS.n6171 VSS.n6170 0.04025
R10621 VSS.n6171 VSS.n2508 0.04025
R10622 VSS.n6175 VSS.n2508 0.04025
R10623 VSS.n6176 VSS.n6175 0.04025
R10624 VSS.n6177 VSS.n6176 0.04025
R10625 VSS.n6177 VSS.n2506 0.04025
R10626 VSS.n6181 VSS.n2506 0.04025
R10627 VSS.n6182 VSS.n6181 0.04025
R10628 VSS.n6183 VSS.n6182 0.04025
R10629 VSS.n6183 VSS.n2504 0.04025
R10630 VSS.n6187 VSS.n2504 0.04025
R10631 VSS.n6188 VSS.n6187 0.04025
R10632 VSS.n6189 VSS.n6188 0.04025
R10633 VSS.n6189 VSS.n2502 0.04025
R10634 VSS.n6193 VSS.n2502 0.04025
R10635 VSS.n6194 VSS.n6193 0.04025
R10636 VSS.n6195 VSS.n6194 0.04025
R10637 VSS.n6195 VSS.n2500 0.04025
R10638 VSS.n6199 VSS.n2500 0.04025
R10639 VSS.n6200 VSS.n6199 0.04025
R10640 VSS.n6201 VSS.n6200 0.04025
R10641 VSS.n6201 VSS.n2498 0.04025
R10642 VSS.n6205 VSS.n2498 0.04025
R10643 VSS.n6206 VSS.n6205 0.04025
R10644 VSS.n6207 VSS.n6206 0.04025
R10645 VSS.n6207 VSS.n2496 0.04025
R10646 VSS.n6211 VSS.n2496 0.04025
R10647 VSS.n6212 VSS.n6211 0.04025
R10648 VSS.n6213 VSS.n6212 0.04025
R10649 VSS.n6213 VSS.n2494 0.04025
R10650 VSS.n6217 VSS.n2494 0.04025
R10651 VSS.n6218 VSS.n6217 0.04025
R10652 VSS.n6219 VSS.n6218 0.04025
R10653 VSS.n6219 VSS.n2492 0.04025
R10654 VSS.n6223 VSS.n2492 0.04025
R10655 VSS.n6224 VSS.n6223 0.04025
R10656 VSS.n6225 VSS.n6224 0.04025
R10657 VSS.n6225 VSS.n2490 0.04025
R10658 VSS.n6229 VSS.n2490 0.04025
R10659 VSS.n6230 VSS.n6229 0.04025
R10660 VSS.n6231 VSS.n6230 0.04025
R10661 VSS.n6231 VSS.n2488 0.04025
R10662 VSS.n6235 VSS.n2488 0.04025
R10663 VSS.n6236 VSS.n6235 0.04025
R10664 VSS.n6237 VSS.n6236 0.04025
R10665 VSS.n6237 VSS.n2486 0.04025
R10666 VSS.n6241 VSS.n2486 0.04025
R10667 VSS.n6242 VSS.n6241 0.04025
R10668 VSS.n6243 VSS.n6242 0.04025
R10669 VSS.n6243 VSS.n2484 0.04025
R10670 VSS.n6247 VSS.n2484 0.04025
R10671 VSS.n6248 VSS.n6247 0.04025
R10672 VSS.n6249 VSS.n6248 0.04025
R10673 VSS.n6249 VSS.n2482 0.04025
R10674 VSS.n6253 VSS.n2482 0.04025
R10675 VSS.n6254 VSS.n6253 0.04025
R10676 VSS.n6255 VSS.n6254 0.04025
R10677 VSS.n6255 VSS.n2480 0.04025
R10678 VSS.n6259 VSS.n2480 0.04025
R10679 VSS.n6260 VSS.n6259 0.04025
R10680 VSS.n6261 VSS.n6260 0.04025
R10681 VSS.n6261 VSS.n2478 0.04025
R10682 VSS.n6265 VSS.n2478 0.04025
R10683 VSS.n6266 VSS.n6265 0.04025
R10684 VSS.n6267 VSS.n6266 0.04025
R10685 VSS.n6267 VSS.n2476 0.04025
R10686 VSS.n6271 VSS.n2476 0.04025
R10687 VSS.n6272 VSS.n6271 0.04025
R10688 VSS.n6273 VSS.n6272 0.04025
R10689 VSS.n6273 VSS.n2474 0.04025
R10690 VSS.n6277 VSS.n2474 0.04025
R10691 VSS.n6278 VSS.n6277 0.04025
R10692 VSS.n6279 VSS.n6278 0.04025
R10693 VSS.n6279 VSS.n2472 0.04025
R10694 VSS.n6283 VSS.n2472 0.04025
R10695 VSS.n6284 VSS.n6283 0.04025
R10696 VSS.n6285 VSS.n6284 0.04025
R10697 VSS.n6285 VSS.n2470 0.04025
R10698 VSS.n6289 VSS.n2470 0.04025
R10699 VSS.n6290 VSS.n6289 0.04025
R10700 VSS.n6291 VSS.n6290 0.04025
R10701 VSS.n6291 VSS.n2468 0.04025
R10702 VSS.n6295 VSS.n2468 0.04025
R10703 VSS.n6296 VSS.n6295 0.04025
R10704 VSS.n6297 VSS.n6296 0.04025
R10705 VSS.n6297 VSS.n2466 0.04025
R10706 VSS.n6301 VSS.n2466 0.04025
R10707 VSS.n6302 VSS.n6301 0.04025
R10708 VSS.n6303 VSS.n6302 0.04025
R10709 VSS.n6303 VSS.n2464 0.04025
R10710 VSS.n6307 VSS.n2464 0.04025
R10711 VSS.n6308 VSS.n6307 0.04025
R10712 VSS.n6309 VSS.n6308 0.04025
R10713 VSS.n6309 VSS.n2462 0.04025
R10714 VSS.n6313 VSS.n2462 0.04025
R10715 VSS.n6314 VSS.n6313 0.04025
R10716 VSS.n6315 VSS.n6314 0.04025
R10717 VSS.n6315 VSS.n2460 0.04025
R10718 VSS.n6319 VSS.n2460 0.04025
R10719 VSS.n6320 VSS.n6319 0.04025
R10720 VSS.n6321 VSS.n6320 0.04025
R10721 VSS.n6321 VSS.n2458 0.04025
R10722 VSS.n6325 VSS.n2458 0.04025
R10723 VSS.n6326 VSS.n6325 0.04025
R10724 VSS.n6327 VSS.n6326 0.04025
R10725 VSS.n6327 VSS.n2456 0.04025
R10726 VSS.n6331 VSS.n2456 0.04025
R10727 VSS.n6332 VSS.n6331 0.04025
R10728 VSS.n6333 VSS.n6332 0.04025
R10729 VSS.n6333 VSS.n2454 0.04025
R10730 VSS.n6337 VSS.n2454 0.04025
R10731 VSS.n6338 VSS.n6337 0.04025
R10732 VSS.n6339 VSS.n6338 0.04025
R10733 VSS.n6339 VSS.n2452 0.04025
R10734 VSS.n6343 VSS.n2452 0.04025
R10735 VSS.n6344 VSS.n6343 0.04025
R10736 VSS.n6345 VSS.n6344 0.04025
R10737 VSS.n6345 VSS.n2450 0.04025
R10738 VSS.n6349 VSS.n2450 0.04025
R10739 VSS.n6350 VSS.n6349 0.04025
R10740 VSS.n6351 VSS.n6350 0.04025
R10741 VSS.n6351 VSS.n2448 0.04025
R10742 VSS.n6355 VSS.n2448 0.04025
R10743 VSS.n6356 VSS.n6355 0.04025
R10744 VSS.n6357 VSS.n6356 0.04025
R10745 VSS.n6357 VSS.n2446 0.04025
R10746 VSS.n6361 VSS.n2446 0.04025
R10747 VSS.n6362 VSS.n6361 0.04025
R10748 VSS.n6363 VSS.n6362 0.04025
R10749 VSS.n6363 VSS.n2444 0.04025
R10750 VSS.n6367 VSS.n2444 0.04025
R10751 VSS.n6368 VSS.n6367 0.04025
R10752 VSS.n6369 VSS.n6368 0.04025
R10753 VSS.n6369 VSS.n2442 0.04025
R10754 VSS.n6373 VSS.n2442 0.04025
R10755 VSS.n6374 VSS.n6373 0.04025
R10756 VSS.n6375 VSS.n6374 0.04025
R10757 VSS.n6375 VSS.n2440 0.04025
R10758 VSS.n6379 VSS.n2440 0.04025
R10759 VSS.n6380 VSS.n6379 0.04025
R10760 VSS.n6381 VSS.n6380 0.04025
R10761 VSS.n6381 VSS.n2438 0.04025
R10762 VSS.n6385 VSS.n2438 0.04025
R10763 VSS.n6386 VSS.n6385 0.04025
R10764 VSS.n6387 VSS.n6386 0.04025
R10765 VSS.n6387 VSS.n2436 0.04025
R10766 VSS.n6391 VSS.n2436 0.04025
R10767 VSS.n6392 VSS.n6391 0.04025
R10768 VSS.n6393 VSS.n6392 0.04025
R10769 VSS.n6393 VSS.n2434 0.04025
R10770 VSS.n6397 VSS.n2434 0.04025
R10771 VSS.n6398 VSS.n6397 0.04025
R10772 VSS.n6399 VSS.n6398 0.04025
R10773 VSS.n6399 VSS.n2432 0.04025
R10774 VSS.n6403 VSS.n2432 0.04025
R10775 VSS.n6404 VSS.n6403 0.04025
R10776 VSS.n6405 VSS.n6404 0.04025
R10777 VSS.n6405 VSS.n2430 0.04025
R10778 VSS.n6409 VSS.n2430 0.04025
R10779 VSS.n6410 VSS.n6409 0.04025
R10780 VSS.n6411 VSS.n6410 0.04025
R10781 VSS.n6411 VSS.n2428 0.04025
R10782 VSS.n6415 VSS.n2428 0.04025
R10783 VSS.n6416 VSS.n6415 0.04025
R10784 VSS.n6417 VSS.n6416 0.04025
R10785 VSS.n6417 VSS.n2426 0.04025
R10786 VSS.n6421 VSS.n2426 0.04025
R10787 VSS.n6422 VSS.n6421 0.04025
R10788 VSS.n6423 VSS.n6422 0.04025
R10789 VSS.n6423 VSS.n2424 0.04025
R10790 VSS.n6427 VSS.n2424 0.04025
R10791 VSS.n6428 VSS.n6427 0.04025
R10792 VSS.n6429 VSS.n6428 0.04025
R10793 VSS.n6429 VSS.n2422 0.04025
R10794 VSS.n6433 VSS.n2422 0.04025
R10795 VSS.n6434 VSS.n6433 0.04025
R10796 VSS.n6435 VSS.n6434 0.04025
R10797 VSS.n6435 VSS.n2420 0.04025
R10798 VSS.n6439 VSS.n2420 0.04025
R10799 VSS.n6440 VSS.n6439 0.04025
R10800 VSS.n6441 VSS.n6440 0.04025
R10801 VSS.n6441 VSS.n2418 0.04025
R10802 VSS.n6445 VSS.n2418 0.04025
R10803 VSS.n6446 VSS.n6445 0.04025
R10804 VSS.n6447 VSS.n6446 0.04025
R10805 VSS.n6447 VSS.n2416 0.04025
R10806 VSS.n6451 VSS.n2416 0.04025
R10807 VSS.n6452 VSS.n6451 0.04025
R10808 VSS.n6453 VSS.n6452 0.04025
R10809 VSS.n6453 VSS.n2414 0.04025
R10810 VSS.n6457 VSS.n2414 0.04025
R10811 VSS.n6458 VSS.n6457 0.04025
R10812 VSS.n6459 VSS.n6458 0.04025
R10813 VSS.n6459 VSS.n2412 0.04025
R10814 VSS.n6463 VSS.n2412 0.04025
R10815 VSS.n6464 VSS.n6463 0.04025
R10816 VSS.n6465 VSS.n6464 0.04025
R10817 VSS.n6465 VSS.n2410 0.04025
R10818 VSS.n6469 VSS.n2410 0.04025
R10819 VSS.n6470 VSS.n6469 0.04025
R10820 VSS.n6471 VSS.n6470 0.04025
R10821 VSS.n6471 VSS.n2408 0.04025
R10822 VSS.n6475 VSS.n2408 0.04025
R10823 VSS.n6476 VSS.n6475 0.04025
R10824 VSS.n6477 VSS.n6476 0.04025
R10825 VSS.n6477 VSS.n2406 0.04025
R10826 VSS.n6481 VSS.n2406 0.04025
R10827 VSS.n6482 VSS.n6481 0.04025
R10828 VSS.n6483 VSS.n6482 0.04025
R10829 VSS.n6483 VSS.n2404 0.04025
R10830 VSS.n6487 VSS.n2404 0.04025
R10831 VSS.n6488 VSS.n6487 0.04025
R10832 VSS.n6489 VSS.n6488 0.04025
R10833 VSS.n6489 VSS.n2402 0.04025
R10834 VSS.n6493 VSS.n2402 0.04025
R10835 VSS.n6494 VSS.n6493 0.04025
R10836 VSS.n6495 VSS.n6494 0.04025
R10837 VSS.n6495 VSS.n2400 0.04025
R10838 VSS.n6499 VSS.n2400 0.04025
R10839 VSS.n6500 VSS.n6499 0.04025
R10840 VSS.n6501 VSS.n6500 0.04025
R10841 VSS.n6501 VSS.n2398 0.04025
R10842 VSS.n6505 VSS.n2398 0.04025
R10843 VSS.n6506 VSS.n6505 0.04025
R10844 VSS.n6507 VSS.n6506 0.04025
R10845 VSS.n6507 VSS.n2396 0.04025
R10846 VSS.n6511 VSS.n2396 0.04025
R10847 VSS.n6512 VSS.n6511 0.04025
R10848 VSS.n6513 VSS.n6512 0.04025
R10849 VSS.n6513 VSS.n2394 0.04025
R10850 VSS.n6517 VSS.n2394 0.04025
R10851 VSS.n6518 VSS.n6517 0.04025
R10852 VSS.n6519 VSS.n6518 0.04025
R10853 VSS.n6519 VSS.n2392 0.04025
R10854 VSS.n6523 VSS.n2392 0.04025
R10855 VSS.n6524 VSS.n6523 0.04025
R10856 VSS.n6525 VSS.n6524 0.04025
R10857 VSS.n6525 VSS.n2390 0.04025
R10858 VSS.n6529 VSS.n2390 0.04025
R10859 VSS.n6530 VSS.n6529 0.04025
R10860 VSS.n6531 VSS.n6530 0.04025
R10861 VSS.n6531 VSS.n2388 0.04025
R10862 VSS.n6535 VSS.n2388 0.04025
R10863 VSS.n6536 VSS.n6535 0.04025
R10864 VSS.n6537 VSS.n6536 0.04025
R10865 VSS.n6537 VSS.n2386 0.04025
R10866 VSS.n6541 VSS.n2386 0.04025
R10867 VSS.n6542 VSS.n6541 0.04025
R10868 VSS.n6543 VSS.n6542 0.04025
R10869 VSS.n6543 VSS.n2384 0.04025
R10870 VSS.n6547 VSS.n2384 0.04025
R10871 VSS.n6548 VSS.n6547 0.04025
R10872 VSS.n6549 VSS.n6548 0.04025
R10873 VSS.n6549 VSS.n2382 0.04025
R10874 VSS.n6553 VSS.n2382 0.04025
R10875 VSS.n6554 VSS.n6553 0.04025
R10876 VSS.n6555 VSS.n6554 0.04025
R10877 VSS.n6555 VSS.n2380 0.04025
R10878 VSS.n6559 VSS.n2380 0.04025
R10879 VSS.n6560 VSS.n6559 0.04025
R10880 VSS.n6561 VSS.n6560 0.04025
R10881 VSS.n6561 VSS.n2378 0.04025
R10882 VSS.n6565 VSS.n2378 0.04025
R10883 VSS.n6566 VSS.n6565 0.04025
R10884 VSS.n6567 VSS.n6566 0.04025
R10885 VSS.n6567 VSS.n2376 0.04025
R10886 VSS.n6571 VSS.n2376 0.04025
R10887 VSS.n6572 VSS.n6571 0.04025
R10888 VSS.n6573 VSS.n6572 0.04025
R10889 VSS.n6573 VSS.n2374 0.04025
R10890 VSS.n6577 VSS.n2374 0.04025
R10891 VSS.n6578 VSS.n6577 0.04025
R10892 VSS.n6579 VSS.n6578 0.04025
R10893 VSS.n6579 VSS.n2372 0.04025
R10894 VSS.n6583 VSS.n2372 0.04025
R10895 VSS.n6584 VSS.n6583 0.04025
R10896 VSS.n6585 VSS.n6584 0.04025
R10897 VSS.n6585 VSS.n2370 0.04025
R10898 VSS.n6589 VSS.n2370 0.04025
R10899 VSS.n6590 VSS.n6589 0.04025
R10900 VSS.n6591 VSS.n6590 0.04025
R10901 VSS.n6591 VSS.n2368 0.04025
R10902 VSS.n6595 VSS.n2368 0.04025
R10903 VSS.n6596 VSS.n6595 0.04025
R10904 VSS.n6597 VSS.n6596 0.04025
R10905 VSS.n6597 VSS.n2366 0.04025
R10906 VSS.n6601 VSS.n2366 0.04025
R10907 VSS.n6602 VSS.n6601 0.04025
R10908 VSS.n6603 VSS.n6602 0.04025
R10909 VSS.n6603 VSS.n2364 0.04025
R10910 VSS.n6607 VSS.n2364 0.04025
R10911 VSS.n6608 VSS.n6607 0.04025
R10912 VSS.n6609 VSS.n6608 0.04025
R10913 VSS.n6609 VSS.n2362 0.04025
R10914 VSS.n6613 VSS.n2362 0.04025
R10915 VSS.n6614 VSS.n6613 0.04025
R10916 VSS.n6615 VSS.n6614 0.04025
R10917 VSS.n6615 VSS.n2360 0.04025
R10918 VSS.n6619 VSS.n2360 0.04025
R10919 VSS.n6620 VSS.n6619 0.04025
R10920 VSS.n6621 VSS.n6620 0.04025
R10921 VSS.n6621 VSS.n2358 0.04025
R10922 VSS.n6625 VSS.n2358 0.04025
R10923 VSS.n6626 VSS.n6625 0.04025
R10924 VSS.n6627 VSS.n6626 0.04025
R10925 VSS.n6627 VSS.n2356 0.04025
R10926 VSS.n6631 VSS.n2356 0.04025
R10927 VSS.n6632 VSS.n6631 0.04025
R10928 VSS.n6633 VSS.n6632 0.04025
R10929 VSS.n6633 VSS.n2354 0.04025
R10930 VSS.n6637 VSS.n2354 0.04025
R10931 VSS.n6638 VSS.n6637 0.04025
R10932 VSS.n6639 VSS.n6638 0.04025
R10933 VSS.n6639 VSS.n2352 0.04025
R10934 VSS.n6643 VSS.n2352 0.04025
R10935 VSS.n6644 VSS.n6643 0.04025
R10936 VSS.n6645 VSS.n6644 0.04025
R10937 VSS.n6645 VSS.n2350 0.04025
R10938 VSS.n6649 VSS.n2350 0.04025
R10939 VSS.n6650 VSS.n6649 0.04025
R10940 VSS.n6651 VSS.n6650 0.04025
R10941 VSS.n6651 VSS.n2348 0.04025
R10942 VSS.n6655 VSS.n2348 0.04025
R10943 VSS.n6656 VSS.n6655 0.04025
R10944 VSS.n6657 VSS.n6656 0.04025
R10945 VSS.n6657 VSS.n2346 0.04025
R10946 VSS.n6661 VSS.n2346 0.04025
R10947 VSS.n6662 VSS.n6661 0.04025
R10948 VSS.n6663 VSS.n6662 0.04025
R10949 VSS.n6663 VSS.n2344 0.04025
R10950 VSS.n6667 VSS.n2344 0.04025
R10951 VSS.n6668 VSS.n6667 0.04025
R10952 VSS.n6669 VSS.n6668 0.04025
R10953 VSS.n6669 VSS.n2342 0.04025
R10954 VSS.n6673 VSS.n2342 0.04025
R10955 VSS.n6674 VSS.n6673 0.04025
R10956 VSS.n6675 VSS.n6674 0.04025
R10957 VSS.n6675 VSS.n2340 0.04025
R10958 VSS.n6679 VSS.n2340 0.04025
R10959 VSS.n6680 VSS.n6679 0.04025
R10960 VSS.n6681 VSS.n6680 0.04025
R10961 VSS.n6681 VSS.n2338 0.04025
R10962 VSS.n6685 VSS.n2338 0.04025
R10963 VSS.n6686 VSS.n6685 0.04025
R10964 VSS.n6687 VSS.n6686 0.04025
R10965 VSS.n6687 VSS.n2336 0.04025
R10966 VSS.n6691 VSS.n2336 0.04025
R10967 VSS.n6692 VSS.n6691 0.04025
R10968 VSS.n6693 VSS.n6692 0.04025
R10969 VSS.n6693 VSS.n2334 0.04025
R10970 VSS.n6697 VSS.n2334 0.04025
R10971 VSS.n6698 VSS.n6697 0.04025
R10972 VSS.n6699 VSS.n6698 0.04025
R10973 VSS.n6699 VSS.n2332 0.04025
R10974 VSS.n6703 VSS.n2332 0.04025
R10975 VSS.n6704 VSS.n6703 0.04025
R10976 VSS.n6705 VSS.n6704 0.04025
R10977 VSS.n6705 VSS.n2330 0.04025
R10978 VSS.n6709 VSS.n2330 0.04025
R10979 VSS.n6710 VSS.n6709 0.04025
R10980 VSS.n6711 VSS.n6710 0.04025
R10981 VSS.n6711 VSS.n2328 0.04025
R10982 VSS.n6715 VSS.n2328 0.04025
R10983 VSS.n6716 VSS.n6715 0.04025
R10984 VSS.n6717 VSS.n6716 0.04025
R10985 VSS.n6717 VSS.n2326 0.04025
R10986 VSS.n6721 VSS.n2326 0.04025
R10987 VSS.n6722 VSS.n6721 0.04025
R10988 VSS.n6723 VSS.n6722 0.04025
R10989 VSS.n6723 VSS.n2324 0.04025
R10990 VSS.n6727 VSS.n2324 0.04025
R10991 VSS.n6728 VSS.n6727 0.04025
R10992 VSS.n6729 VSS.n6728 0.04025
R10993 VSS.n6729 VSS.n2322 0.04025
R10994 VSS.n6733 VSS.n2322 0.04025
R10995 VSS.n6734 VSS.n6733 0.04025
R10996 VSS.n6735 VSS.n6734 0.04025
R10997 VSS.n6735 VSS.n2320 0.04025
R10998 VSS.n6739 VSS.n2320 0.04025
R10999 VSS.n6740 VSS.n6739 0.04025
R11000 VSS.n6741 VSS.n6740 0.04025
R11001 VSS.n6741 VSS.n2318 0.04025
R11002 VSS.n6745 VSS.n2318 0.04025
R11003 VSS.n6746 VSS.n6745 0.04025
R11004 VSS.n6747 VSS.n6746 0.04025
R11005 VSS.n6747 VSS.n2316 0.04025
R11006 VSS.n6751 VSS.n2316 0.04025
R11007 VSS.n6752 VSS.n6751 0.04025
R11008 VSS.n6753 VSS.n6752 0.04025
R11009 VSS.n6753 VSS.n2314 0.04025
R11010 VSS.n6757 VSS.n2314 0.04025
R11011 VSS.n6758 VSS.n6757 0.04025
R11012 VSS.n6759 VSS.n6758 0.04025
R11013 VSS.n6759 VSS.n2312 0.04025
R11014 VSS.n6763 VSS.n2312 0.04025
R11015 VSS.n6764 VSS.n6763 0.04025
R11016 VSS.n6765 VSS.n6764 0.04025
R11017 VSS.n6765 VSS.n2310 0.04025
R11018 VSS.n6769 VSS.n2310 0.04025
R11019 VSS.n6770 VSS.n6769 0.04025
R11020 VSS.n6771 VSS.n6770 0.04025
R11021 VSS.n6771 VSS.n2308 0.04025
R11022 VSS.n6775 VSS.n2308 0.04025
R11023 VSS.n6776 VSS.n6775 0.04025
R11024 VSS.n6777 VSS.n6776 0.04025
R11025 VSS.n6777 VSS.n2306 0.04025
R11026 VSS.n6781 VSS.n2306 0.04025
R11027 VSS.n6782 VSS.n6781 0.04025
R11028 VSS.n6783 VSS.n6782 0.04025
R11029 VSS.n6783 VSS.n2304 0.04025
R11030 VSS.n6787 VSS.n2304 0.04025
R11031 VSS.n6788 VSS.n6787 0.04025
R11032 VSS.n6789 VSS.n6788 0.04025
R11033 VSS.n6789 VSS.n2302 0.04025
R11034 VSS.n6793 VSS.n2302 0.04025
R11035 VSS.n6794 VSS.n6793 0.04025
R11036 VSS.n6795 VSS.n6794 0.04025
R11037 VSS.n6795 VSS.n2300 0.04025
R11038 VSS.n6799 VSS.n2300 0.04025
R11039 VSS.n6800 VSS.n6799 0.04025
R11040 VSS.n6801 VSS.n6800 0.04025
R11041 VSS.n6801 VSS.n2298 0.04025
R11042 VSS.n6805 VSS.n2298 0.04025
R11043 VSS.n6806 VSS.n6805 0.04025
R11044 VSS.n6807 VSS.n6806 0.04025
R11045 VSS.n6807 VSS.n2296 0.04025
R11046 VSS.n6811 VSS.n2296 0.04025
R11047 VSS.n6812 VSS.n6811 0.04025
R11048 VSS.n6813 VSS.n6812 0.04025
R11049 VSS.n6813 VSS.n2294 0.04025
R11050 VSS.n6817 VSS.n2294 0.04025
R11051 VSS.n6818 VSS.n6817 0.04025
R11052 VSS.n6819 VSS.n6818 0.04025
R11053 VSS.n6819 VSS.n2292 0.04025
R11054 VSS.n6823 VSS.n2292 0.04025
R11055 VSS.n6824 VSS.n6823 0.04025
R11056 VSS.n6825 VSS.n6824 0.04025
R11057 VSS.n6825 VSS.n2290 0.04025
R11058 VSS.n6829 VSS.n2290 0.04025
R11059 VSS.n6830 VSS.n6829 0.04025
R11060 VSS.n6831 VSS.n6830 0.04025
R11061 VSS.n6831 VSS.n2288 0.04025
R11062 VSS.n6835 VSS.n2288 0.04025
R11063 VSS.n6836 VSS.n6835 0.04025
R11064 VSS.n6837 VSS.n6836 0.04025
R11065 VSS.n6837 VSS.n2286 0.04025
R11066 VSS.n6841 VSS.n2286 0.04025
R11067 VSS.n6842 VSS.n6841 0.04025
R11068 VSS.n6843 VSS.n6842 0.04025
R11069 VSS.n6843 VSS.n2284 0.04025
R11070 VSS.n6847 VSS.n2284 0.04025
R11071 VSS.n6848 VSS.n6847 0.04025
R11072 VSS.n6849 VSS.n6848 0.04025
R11073 VSS.n6849 VSS.n2282 0.04025
R11074 VSS.n6853 VSS.n2282 0.04025
R11075 VSS.n6854 VSS.n6853 0.04025
R11076 VSS.n6855 VSS.n6854 0.04025
R11077 VSS.n6855 VSS.n2280 0.04025
R11078 VSS.n6859 VSS.n2280 0.04025
R11079 VSS.n6860 VSS.n6859 0.04025
R11080 VSS.n6861 VSS.n6860 0.04025
R11081 VSS.n6861 VSS.n2278 0.04025
R11082 VSS.n6865 VSS.n2278 0.04025
R11083 VSS.n6866 VSS.n6865 0.04025
R11084 VSS.n6867 VSS.n6866 0.04025
R11085 VSS.n6867 VSS.n2276 0.04025
R11086 VSS.n6871 VSS.n2276 0.04025
R11087 VSS.n6872 VSS.n6871 0.04025
R11088 VSS.n6873 VSS.n6872 0.04025
R11089 VSS.n6873 VSS.n2274 0.04025
R11090 VSS.n6877 VSS.n2274 0.04025
R11091 VSS.n6878 VSS.n6877 0.04025
R11092 VSS.n6879 VSS.n6878 0.04025
R11093 VSS.n6879 VSS.n2272 0.04025
R11094 VSS.n6883 VSS.n2272 0.04025
R11095 VSS.n6884 VSS.n6883 0.04025
R11096 VSS.n6885 VSS.n6884 0.04025
R11097 VSS.n6885 VSS.n2270 0.04025
R11098 VSS.n6889 VSS.n2270 0.04025
R11099 VSS.n6890 VSS.n6889 0.04025
R11100 VSS.n6891 VSS.n6890 0.04025
R11101 VSS.n6891 VSS.n2268 0.04025
R11102 VSS.n6895 VSS.n2268 0.04025
R11103 VSS.n6896 VSS.n6895 0.04025
R11104 VSS.n6897 VSS.n6896 0.04025
R11105 VSS.n6897 VSS.n2266 0.04025
R11106 VSS.n6901 VSS.n2266 0.04025
R11107 VSS.n6902 VSS.n6901 0.04025
R11108 VSS.n6903 VSS.n6902 0.04025
R11109 VSS.n6903 VSS.n2264 0.04025
R11110 VSS.n6907 VSS.n2264 0.04025
R11111 VSS.n8229 VSS.n1822 0.04025
R11112 VSS.n8229 VSS.n8228 0.04025
R11113 VSS.n8228 VSS.n8227 0.04025
R11114 VSS.n8227 VSS.n1824 0.04025
R11115 VSS.n8223 VSS.n1824 0.04025
R11116 VSS.n8223 VSS.n8222 0.04025
R11117 VSS.n8222 VSS.n8221 0.04025
R11118 VSS.n8221 VSS.n1826 0.04025
R11119 VSS.n8217 VSS.n1826 0.04025
R11120 VSS.n8217 VSS.n8216 0.04025
R11121 VSS.n8216 VSS.n8215 0.04025
R11122 VSS.n8215 VSS.n1828 0.04025
R11123 VSS.n8211 VSS.n1828 0.04025
R11124 VSS.n8211 VSS.n8210 0.04025
R11125 VSS.n8210 VSS.n8209 0.04025
R11126 VSS.n8209 VSS.n1830 0.04025
R11127 VSS.n8205 VSS.n1830 0.04025
R11128 VSS.n8205 VSS.n8204 0.04025
R11129 VSS.n8204 VSS.n8203 0.04025
R11130 VSS.n8203 VSS.n1832 0.04025
R11131 VSS.n8199 VSS.n1832 0.04025
R11132 VSS.n8199 VSS.n8198 0.04025
R11133 VSS.n8198 VSS.n8197 0.04025
R11134 VSS.n8197 VSS.n1834 0.04025
R11135 VSS.n8193 VSS.n1834 0.04025
R11136 VSS.n8193 VSS.n8192 0.04025
R11137 VSS.n8192 VSS.n8191 0.04025
R11138 VSS.n8191 VSS.n1836 0.04025
R11139 VSS.n8187 VSS.n1836 0.04025
R11140 VSS.n8187 VSS.n8186 0.04025
R11141 VSS.n8186 VSS.n8185 0.04025
R11142 VSS.n8185 VSS.n1838 0.04025
R11143 VSS.n8181 VSS.n1838 0.04025
R11144 VSS.n8181 VSS.n8180 0.04025
R11145 VSS.n8180 VSS.n8179 0.04025
R11146 VSS.n8179 VSS.n1840 0.04025
R11147 VSS.n8175 VSS.n1840 0.04025
R11148 VSS.n8175 VSS.n8174 0.04025
R11149 VSS.n8174 VSS.n8173 0.04025
R11150 VSS.n8173 VSS.n1842 0.04025
R11151 VSS.n8169 VSS.n1842 0.04025
R11152 VSS.n8169 VSS.n8168 0.04025
R11153 VSS.n8168 VSS.n8167 0.04025
R11154 VSS.n8167 VSS.n1844 0.04025
R11155 VSS.n8163 VSS.n1844 0.04025
R11156 VSS.n8163 VSS.n8162 0.04025
R11157 VSS.n8162 VSS.n8161 0.04025
R11158 VSS.n8161 VSS.n1846 0.04025
R11159 VSS.n8157 VSS.n1846 0.04025
R11160 VSS.n8157 VSS.n8156 0.04025
R11161 VSS.n8156 VSS.n8155 0.04025
R11162 VSS.n8155 VSS.n1848 0.04025
R11163 VSS.n8151 VSS.n1848 0.04025
R11164 VSS.n8151 VSS.n8150 0.04025
R11165 VSS.n8150 VSS.n8149 0.04025
R11166 VSS.n8149 VSS.n1850 0.04025
R11167 VSS.n8145 VSS.n1850 0.04025
R11168 VSS.n8145 VSS.n8144 0.04025
R11169 VSS.n8144 VSS.n8143 0.04025
R11170 VSS.n8143 VSS.n1852 0.04025
R11171 VSS.n8139 VSS.n1852 0.04025
R11172 VSS.n8139 VSS.n8138 0.04025
R11173 VSS.n8138 VSS.n8137 0.04025
R11174 VSS.n8137 VSS.n1854 0.04025
R11175 VSS.n8133 VSS.n1854 0.04025
R11176 VSS.n8133 VSS.n8132 0.04025
R11177 VSS.n8132 VSS.n8131 0.04025
R11178 VSS.n8131 VSS.n1856 0.04025
R11179 VSS.n8127 VSS.n1856 0.04025
R11180 VSS.n8127 VSS.n8126 0.04025
R11181 VSS.n8126 VSS.n8125 0.04025
R11182 VSS.n8125 VSS.n1858 0.04025
R11183 VSS.n8121 VSS.n1858 0.04025
R11184 VSS.n8121 VSS.n8120 0.04025
R11185 VSS.n8120 VSS.n8119 0.04025
R11186 VSS.n8119 VSS.n1860 0.04025
R11187 VSS.n8115 VSS.n1860 0.04025
R11188 VSS.n8115 VSS.n8114 0.04025
R11189 VSS.n8114 VSS.n8113 0.04025
R11190 VSS.n8113 VSS.n1862 0.04025
R11191 VSS.n8109 VSS.n1862 0.04025
R11192 VSS.n8109 VSS.n8108 0.04025
R11193 VSS.n8108 VSS.n8107 0.04025
R11194 VSS.n8107 VSS.n1864 0.04025
R11195 VSS.n8103 VSS.n1864 0.04025
R11196 VSS.n8103 VSS.n8102 0.04025
R11197 VSS.n8102 VSS.n8101 0.04025
R11198 VSS.n8101 VSS.n1866 0.04025
R11199 VSS.n8097 VSS.n1866 0.04025
R11200 VSS.n8097 VSS.n8096 0.04025
R11201 VSS.n8096 VSS.n8095 0.04025
R11202 VSS.n8095 VSS.n1868 0.04025
R11203 VSS.n8091 VSS.n1868 0.04025
R11204 VSS.n8091 VSS.n8090 0.04025
R11205 VSS.n8090 VSS.n8089 0.04025
R11206 VSS.n8089 VSS.n1870 0.04025
R11207 VSS.n8085 VSS.n1870 0.04025
R11208 VSS.n8085 VSS.n8084 0.04025
R11209 VSS.n8084 VSS.n8083 0.04025
R11210 VSS.n8083 VSS.n1872 0.04025
R11211 VSS.n8079 VSS.n1872 0.04025
R11212 VSS.n8079 VSS.n8078 0.04025
R11213 VSS.n8078 VSS.n8077 0.04025
R11214 VSS.n8077 VSS.n1874 0.04025
R11215 VSS.n8073 VSS.n1874 0.04025
R11216 VSS.n8073 VSS.n8072 0.04025
R11217 VSS.n8072 VSS.n8071 0.04025
R11218 VSS.n8071 VSS.n1876 0.04025
R11219 VSS.n8067 VSS.n1876 0.04025
R11220 VSS.n8067 VSS.n8066 0.04025
R11221 VSS.n8066 VSS.n8065 0.04025
R11222 VSS.n8065 VSS.n1878 0.04025
R11223 VSS.n8061 VSS.n1878 0.04025
R11224 VSS.n8061 VSS.n8060 0.04025
R11225 VSS.n8060 VSS.n8059 0.04025
R11226 VSS.n8059 VSS.n1880 0.04025
R11227 VSS.n8055 VSS.n1880 0.04025
R11228 VSS.n8055 VSS.n8054 0.04025
R11229 VSS.n8054 VSS.n8053 0.04025
R11230 VSS.n8053 VSS.n1882 0.04025
R11231 VSS.n8049 VSS.n1882 0.04025
R11232 VSS.n8049 VSS.n8048 0.04025
R11233 VSS.n8048 VSS.n8047 0.04025
R11234 VSS.n8047 VSS.n1884 0.04025
R11235 VSS.n8043 VSS.n1884 0.04025
R11236 VSS.n8043 VSS.n8042 0.04025
R11237 VSS.n8042 VSS.n8041 0.04025
R11238 VSS.n8041 VSS.n1886 0.04025
R11239 VSS.n8037 VSS.n1886 0.04025
R11240 VSS.n8037 VSS.n8036 0.04025
R11241 VSS.n8036 VSS.n8035 0.04025
R11242 VSS.n8035 VSS.n1888 0.04025
R11243 VSS.n8031 VSS.n1888 0.04025
R11244 VSS.n8031 VSS.n8030 0.04025
R11245 VSS.n8030 VSS.n8029 0.04025
R11246 VSS.n8029 VSS.n1890 0.04025
R11247 VSS.n8025 VSS.n1890 0.04025
R11248 VSS.n8025 VSS.n8024 0.04025
R11249 VSS.n8024 VSS.n8023 0.04025
R11250 VSS.n8023 VSS.n1892 0.04025
R11251 VSS.n8019 VSS.n1892 0.04025
R11252 VSS.n8019 VSS.n8018 0.04025
R11253 VSS.n8018 VSS.n8017 0.04025
R11254 VSS.n8017 VSS.n1894 0.04025
R11255 VSS.n8013 VSS.n1894 0.04025
R11256 VSS.n8013 VSS.n8012 0.04025
R11257 VSS.n8012 VSS.n8011 0.04025
R11258 VSS.n8011 VSS.n1896 0.04025
R11259 VSS.n8007 VSS.n1896 0.04025
R11260 VSS.n8007 VSS.n8006 0.04025
R11261 VSS.n8006 VSS.n8005 0.04025
R11262 VSS.n8005 VSS.n1898 0.04025
R11263 VSS.n8001 VSS.n1898 0.04025
R11264 VSS.n8001 VSS.n8000 0.04025
R11265 VSS.n8000 VSS.n7999 0.04025
R11266 VSS.n7999 VSS.n1900 0.04025
R11267 VSS.n7995 VSS.n1900 0.04025
R11268 VSS.n7995 VSS.n7994 0.04025
R11269 VSS.n7994 VSS.n7993 0.04025
R11270 VSS.n7993 VSS.n1902 0.04025
R11271 VSS.n7989 VSS.n1902 0.04025
R11272 VSS.n7989 VSS.n7988 0.04025
R11273 VSS.n7988 VSS.n7987 0.04025
R11274 VSS.n7987 VSS.n1904 0.04025
R11275 VSS.n7983 VSS.n1904 0.04025
R11276 VSS.n7983 VSS.n7982 0.04025
R11277 VSS.n7982 VSS.n7981 0.04025
R11278 VSS.n7981 VSS.n1906 0.04025
R11279 VSS.n7977 VSS.n1906 0.04025
R11280 VSS.n7977 VSS.n7976 0.04025
R11281 VSS.n7976 VSS.n7975 0.04025
R11282 VSS.n7975 VSS.n1908 0.04025
R11283 VSS.n7971 VSS.n1908 0.04025
R11284 VSS.n7971 VSS.n7970 0.04025
R11285 VSS.n7970 VSS.n7969 0.04025
R11286 VSS.n7969 VSS.n1910 0.04025
R11287 VSS.n7965 VSS.n1910 0.04025
R11288 VSS.n7965 VSS.n7964 0.04025
R11289 VSS.n7964 VSS.n7963 0.04025
R11290 VSS.n7963 VSS.n1912 0.04025
R11291 VSS.n7959 VSS.n1912 0.04025
R11292 VSS.n7959 VSS.n7958 0.04025
R11293 VSS.n7958 VSS.n7957 0.04025
R11294 VSS.n7957 VSS.n1914 0.04025
R11295 VSS.n7953 VSS.n1914 0.04025
R11296 VSS.n7953 VSS.n7952 0.04025
R11297 VSS.n7952 VSS.n7951 0.04025
R11298 VSS.n7951 VSS.n1916 0.04025
R11299 VSS.n7947 VSS.n1916 0.04025
R11300 VSS.n7947 VSS.n7946 0.04025
R11301 VSS.n7946 VSS.n7945 0.04025
R11302 VSS.n7945 VSS.n1918 0.04025
R11303 VSS.n7941 VSS.n1918 0.04025
R11304 VSS.n7941 VSS.n7940 0.04025
R11305 VSS.n7940 VSS.n7939 0.04025
R11306 VSS.n7939 VSS.n1920 0.04025
R11307 VSS.n7935 VSS.n1920 0.04025
R11308 VSS.n7935 VSS.n7934 0.04025
R11309 VSS.n7934 VSS.n7933 0.04025
R11310 VSS.n7933 VSS.n1922 0.04025
R11311 VSS.n7929 VSS.n1922 0.04025
R11312 VSS.n7929 VSS.n7928 0.04025
R11313 VSS.n7928 VSS.n7927 0.04025
R11314 VSS.n7927 VSS.n1924 0.04025
R11315 VSS.n7923 VSS.n1924 0.04025
R11316 VSS.n7923 VSS.n7922 0.04025
R11317 VSS.n7922 VSS.n7921 0.04025
R11318 VSS.n7921 VSS.n1926 0.04025
R11319 VSS.n7917 VSS.n1926 0.04025
R11320 VSS.n7917 VSS.n7916 0.04025
R11321 VSS.n7916 VSS.n7915 0.04025
R11322 VSS.n7915 VSS.n1928 0.04025
R11323 VSS.n7911 VSS.n1928 0.04025
R11324 VSS.n7911 VSS.n7910 0.04025
R11325 VSS.n7910 VSS.n7909 0.04025
R11326 VSS.n7909 VSS.n1930 0.04025
R11327 VSS.n7905 VSS.n1930 0.04025
R11328 VSS.n7905 VSS.n7904 0.04025
R11329 VSS.n7904 VSS.n7903 0.04025
R11330 VSS.n7903 VSS.n1932 0.04025
R11331 VSS.n7899 VSS.n1932 0.04025
R11332 VSS.n7899 VSS.n7898 0.04025
R11333 VSS.n7898 VSS.n7897 0.04025
R11334 VSS.n7897 VSS.n1934 0.04025
R11335 VSS.n7893 VSS.n1934 0.04025
R11336 VSS.n7893 VSS.n7892 0.04025
R11337 VSS.n7892 VSS.n7891 0.04025
R11338 VSS.n7891 VSS.n1936 0.04025
R11339 VSS.n7887 VSS.n1936 0.04025
R11340 VSS.n7887 VSS.n7886 0.04025
R11341 VSS.n7886 VSS.n7885 0.04025
R11342 VSS.n7885 VSS.n1938 0.04025
R11343 VSS.n7881 VSS.n1938 0.04025
R11344 VSS.n7881 VSS.n7880 0.04025
R11345 VSS.n7880 VSS.n7879 0.04025
R11346 VSS.n7879 VSS.n1940 0.04025
R11347 VSS.n7875 VSS.n1940 0.04025
R11348 VSS.n7875 VSS.n7874 0.04025
R11349 VSS.n7874 VSS.n7873 0.04025
R11350 VSS.n7873 VSS.n1942 0.04025
R11351 VSS.n7869 VSS.n1942 0.04025
R11352 VSS.n7869 VSS.n7868 0.04025
R11353 VSS.n7868 VSS.n7867 0.04025
R11354 VSS.n7867 VSS.n1944 0.04025
R11355 VSS.n7863 VSS.n1944 0.04025
R11356 VSS.n7863 VSS.n7862 0.04025
R11357 VSS.n7862 VSS.n7861 0.04025
R11358 VSS.n7861 VSS.n1946 0.04025
R11359 VSS.n7857 VSS.n1946 0.04025
R11360 VSS.n7857 VSS.n7856 0.04025
R11361 VSS.n7856 VSS.n7855 0.04025
R11362 VSS.n7855 VSS.n1948 0.04025
R11363 VSS.n7851 VSS.n1948 0.04025
R11364 VSS.n7851 VSS.n7850 0.04025
R11365 VSS.n7850 VSS.n7849 0.04025
R11366 VSS.n7849 VSS.n1950 0.04025
R11367 VSS.n7845 VSS.n1950 0.04025
R11368 VSS.n7845 VSS.n7844 0.04025
R11369 VSS.n7844 VSS.n7843 0.04025
R11370 VSS.n7843 VSS.n1952 0.04025
R11371 VSS.n7839 VSS.n1952 0.04025
R11372 VSS.n7839 VSS.n7838 0.04025
R11373 VSS.n7838 VSS.n7837 0.04025
R11374 VSS.n7837 VSS.n1954 0.04025
R11375 VSS.n7833 VSS.n1954 0.04025
R11376 VSS.n7833 VSS.n7832 0.04025
R11377 VSS.n7832 VSS.n7831 0.04025
R11378 VSS.n7831 VSS.n1956 0.04025
R11379 VSS.n7827 VSS.n1956 0.04025
R11380 VSS.n7827 VSS.n7826 0.04025
R11381 VSS.n7826 VSS.n7825 0.04025
R11382 VSS.n7825 VSS.n1958 0.04025
R11383 VSS.n7821 VSS.n1958 0.04025
R11384 VSS.n7821 VSS.n7820 0.04025
R11385 VSS.n7820 VSS.n7819 0.04025
R11386 VSS.n7819 VSS.n1960 0.04025
R11387 VSS.n7815 VSS.n1960 0.04025
R11388 VSS.n7815 VSS.n7814 0.04025
R11389 VSS.n7814 VSS.n7813 0.04025
R11390 VSS.n7813 VSS.n1962 0.04025
R11391 VSS.n7809 VSS.n1962 0.04025
R11392 VSS.n7809 VSS.n7808 0.04025
R11393 VSS.n7808 VSS.n7807 0.04025
R11394 VSS.n7807 VSS.n1964 0.04025
R11395 VSS.n7803 VSS.n1964 0.04025
R11396 VSS.n7803 VSS.n7802 0.04025
R11397 VSS.n7802 VSS.n7801 0.04025
R11398 VSS.n7801 VSS.n1966 0.04025
R11399 VSS.n7797 VSS.n1966 0.04025
R11400 VSS.n7797 VSS.n7796 0.04025
R11401 VSS.n7796 VSS.n7795 0.04025
R11402 VSS.n7795 VSS.n1968 0.04025
R11403 VSS.n7791 VSS.n1968 0.04025
R11404 VSS.n7791 VSS.n7790 0.04025
R11405 VSS.n7790 VSS.n7789 0.04025
R11406 VSS.n7789 VSS.n1970 0.04025
R11407 VSS.n7785 VSS.n1970 0.04025
R11408 VSS.n7785 VSS.n7784 0.04025
R11409 VSS.n7784 VSS.n7783 0.04025
R11410 VSS.n7783 VSS.n1972 0.04025
R11411 VSS.n7779 VSS.n1972 0.04025
R11412 VSS.n7779 VSS.n7778 0.04025
R11413 VSS.n7778 VSS.n7777 0.04025
R11414 VSS.n7777 VSS.n1974 0.04025
R11415 VSS.n7773 VSS.n1974 0.04025
R11416 VSS.n7773 VSS.n7772 0.04025
R11417 VSS.n7772 VSS.n7771 0.04025
R11418 VSS.n7771 VSS.n1976 0.04025
R11419 VSS.n7767 VSS.n1976 0.04025
R11420 VSS.n7767 VSS.n7766 0.04025
R11421 VSS.n7766 VSS.n7765 0.04025
R11422 VSS.n7765 VSS.n1978 0.04025
R11423 VSS.n7761 VSS.n1978 0.04025
R11424 VSS.n7761 VSS.n7760 0.04025
R11425 VSS.n7760 VSS.n7759 0.04025
R11426 VSS.n7759 VSS.n1980 0.04025
R11427 VSS.n7755 VSS.n1980 0.04025
R11428 VSS.n7755 VSS.n7754 0.04025
R11429 VSS.n7754 VSS.n7753 0.04025
R11430 VSS.n7753 VSS.n1982 0.04025
R11431 VSS.n7749 VSS.n1982 0.04025
R11432 VSS.n7749 VSS.n7748 0.04025
R11433 VSS.n7748 VSS.n7747 0.04025
R11434 VSS.n7747 VSS.n1984 0.04025
R11435 VSS.n7743 VSS.n1984 0.04025
R11436 VSS.n7743 VSS.n7742 0.04025
R11437 VSS.n7742 VSS.n7741 0.04025
R11438 VSS.n7741 VSS.n1986 0.04025
R11439 VSS.n7737 VSS.n1986 0.04025
R11440 VSS.n7737 VSS.n7736 0.04025
R11441 VSS.n7736 VSS.n7735 0.04025
R11442 VSS.n7735 VSS.n1988 0.04025
R11443 VSS.n7731 VSS.n1988 0.04025
R11444 VSS.n7731 VSS.n7730 0.04025
R11445 VSS.n7730 VSS.n7729 0.04025
R11446 VSS.n7729 VSS.n1990 0.04025
R11447 VSS.n7725 VSS.n1990 0.04025
R11448 VSS.n7725 VSS.n7724 0.04025
R11449 VSS.n7724 VSS.n7723 0.04025
R11450 VSS.n7723 VSS.n1992 0.04025
R11451 VSS.n7719 VSS.n1992 0.04025
R11452 VSS.n7719 VSS.n7718 0.04025
R11453 VSS.n7718 VSS.n7717 0.04025
R11454 VSS.n7717 VSS.n1994 0.04025
R11455 VSS.n7713 VSS.n1994 0.04025
R11456 VSS.n7713 VSS.n7712 0.04025
R11457 VSS.n7712 VSS.n7711 0.04025
R11458 VSS.n7711 VSS.n1996 0.04025
R11459 VSS.n7707 VSS.n1996 0.04025
R11460 VSS.n7707 VSS.n7706 0.04025
R11461 VSS.n7706 VSS.n7705 0.04025
R11462 VSS.n7705 VSS.n1998 0.04025
R11463 VSS.n7701 VSS.n1998 0.04025
R11464 VSS.n7701 VSS.n7700 0.04025
R11465 VSS.n7700 VSS.n7699 0.04025
R11466 VSS.n7699 VSS.n2000 0.04025
R11467 VSS.n7695 VSS.n2000 0.04025
R11468 VSS.n7695 VSS.n7694 0.04025
R11469 VSS.n7694 VSS.n7693 0.04025
R11470 VSS.n7693 VSS.n2002 0.04025
R11471 VSS.n7689 VSS.n2002 0.04025
R11472 VSS.n7689 VSS.n7688 0.04025
R11473 VSS.n7688 VSS.n7687 0.04025
R11474 VSS.n7687 VSS.n2004 0.04025
R11475 VSS.n7683 VSS.n2004 0.04025
R11476 VSS.n7683 VSS.n7682 0.04025
R11477 VSS.n7682 VSS.n7681 0.04025
R11478 VSS.n7681 VSS.n2006 0.04025
R11479 VSS.n7677 VSS.n2006 0.04025
R11480 VSS.n7677 VSS.n7676 0.04025
R11481 VSS.n7676 VSS.n7675 0.04025
R11482 VSS.n7675 VSS.n2008 0.04025
R11483 VSS.n7671 VSS.n2008 0.04025
R11484 VSS.n7671 VSS.n7670 0.04025
R11485 VSS.n7670 VSS.n7669 0.04025
R11486 VSS.n7669 VSS.n2010 0.04025
R11487 VSS.n7665 VSS.n2010 0.04025
R11488 VSS.n7665 VSS.n7664 0.04025
R11489 VSS.n7664 VSS.n7663 0.04025
R11490 VSS.n7663 VSS.n2012 0.04025
R11491 VSS.n7659 VSS.n2012 0.04025
R11492 VSS.n7659 VSS.n7658 0.04025
R11493 VSS.n7658 VSS.n7657 0.04025
R11494 VSS.n7657 VSS.n2014 0.04025
R11495 VSS.n7653 VSS.n2014 0.04025
R11496 VSS.n7653 VSS.n7652 0.04025
R11497 VSS.n7652 VSS.n7651 0.04025
R11498 VSS.n7651 VSS.n2016 0.04025
R11499 VSS.n7647 VSS.n2016 0.04025
R11500 VSS.n7647 VSS.n7646 0.04025
R11501 VSS.n7646 VSS.n7645 0.04025
R11502 VSS.n7645 VSS.n2018 0.04025
R11503 VSS.n7641 VSS.n2018 0.04025
R11504 VSS.n7641 VSS.n7640 0.04025
R11505 VSS.n7640 VSS.n7639 0.04025
R11506 VSS.n7639 VSS.n2020 0.04025
R11507 VSS.n7635 VSS.n2020 0.04025
R11508 VSS.n7635 VSS.n7634 0.04025
R11509 VSS.n7634 VSS.n7633 0.04025
R11510 VSS.n7633 VSS.n2022 0.04025
R11511 VSS.n7629 VSS.n2022 0.04025
R11512 VSS.n7629 VSS.n7628 0.04025
R11513 VSS.n7628 VSS.n7627 0.04025
R11514 VSS.n7627 VSS.n2024 0.04025
R11515 VSS.n7623 VSS.n2024 0.04025
R11516 VSS.n7623 VSS.n7622 0.04025
R11517 VSS.n7622 VSS.n7621 0.04025
R11518 VSS.n7621 VSS.n2026 0.04025
R11519 VSS.n7617 VSS.n2026 0.04025
R11520 VSS.n7617 VSS.n7616 0.04025
R11521 VSS.n7616 VSS.n7615 0.04025
R11522 VSS.n7615 VSS.n2028 0.04025
R11523 VSS.n7611 VSS.n2028 0.04025
R11524 VSS.n7611 VSS.n7610 0.04025
R11525 VSS.n7610 VSS.n7609 0.04025
R11526 VSS.n7609 VSS.n2030 0.04025
R11527 VSS.n7605 VSS.n2030 0.04025
R11528 VSS.n7605 VSS.n7604 0.04025
R11529 VSS.n7604 VSS.n7603 0.04025
R11530 VSS.n7603 VSS.n2032 0.04025
R11531 VSS.n7599 VSS.n2032 0.04025
R11532 VSS.n7599 VSS.n7598 0.04025
R11533 VSS.n7598 VSS.n7597 0.04025
R11534 VSS.n7597 VSS.n2034 0.04025
R11535 VSS.n7593 VSS.n2034 0.04025
R11536 VSS.n7593 VSS.n7592 0.04025
R11537 VSS.n7592 VSS.n7591 0.04025
R11538 VSS.n7591 VSS.n2036 0.04025
R11539 VSS.n7587 VSS.n2036 0.04025
R11540 VSS.n7587 VSS.n7586 0.04025
R11541 VSS.n7586 VSS.n7585 0.04025
R11542 VSS.n7585 VSS.n2038 0.04025
R11543 VSS.n7581 VSS.n2038 0.04025
R11544 VSS.n7581 VSS.n7580 0.04025
R11545 VSS.n7580 VSS.n7579 0.04025
R11546 VSS.n7579 VSS.n2040 0.04025
R11547 VSS.n7575 VSS.n2040 0.04025
R11548 VSS.n7575 VSS.n7574 0.04025
R11549 VSS.n7574 VSS.n7573 0.04025
R11550 VSS.n7573 VSS.n2042 0.04025
R11551 VSS.n7569 VSS.n2042 0.04025
R11552 VSS.n7569 VSS.n7568 0.04025
R11553 VSS.n7568 VSS.n7567 0.04025
R11554 VSS.n7567 VSS.n2044 0.04025
R11555 VSS.n7563 VSS.n2044 0.04025
R11556 VSS.n7563 VSS.n7562 0.04025
R11557 VSS.n7562 VSS.n7561 0.04025
R11558 VSS.n7561 VSS.n2046 0.04025
R11559 VSS.n7557 VSS.n2046 0.04025
R11560 VSS.n7557 VSS.n7556 0.04025
R11561 VSS.n7556 VSS.n7555 0.04025
R11562 VSS.n7555 VSS.n2048 0.04025
R11563 VSS.n7551 VSS.n2048 0.04025
R11564 VSS.n7551 VSS.n7550 0.04025
R11565 VSS.n7550 VSS.n7549 0.04025
R11566 VSS.n7549 VSS.n2050 0.04025
R11567 VSS.n7545 VSS.n2050 0.04025
R11568 VSS.n7545 VSS.n7544 0.04025
R11569 VSS.n7544 VSS.n7543 0.04025
R11570 VSS.n7543 VSS.n2052 0.04025
R11571 VSS.n7539 VSS.n2052 0.04025
R11572 VSS.n7539 VSS.n7538 0.04025
R11573 VSS.n7538 VSS.n7537 0.04025
R11574 VSS.n7537 VSS.n2054 0.04025
R11575 VSS.n7533 VSS.n2054 0.04025
R11576 VSS.n7533 VSS.n7532 0.04025
R11577 VSS.n7532 VSS.n7531 0.04025
R11578 VSS.n7531 VSS.n2056 0.04025
R11579 VSS.n7527 VSS.n2056 0.04025
R11580 VSS.n7527 VSS.n7526 0.04025
R11581 VSS.n7526 VSS.n7525 0.04025
R11582 VSS.n7525 VSS.n2058 0.04025
R11583 VSS.n7521 VSS.n2058 0.04025
R11584 VSS.n7521 VSS.n7520 0.04025
R11585 VSS.n7520 VSS.n7519 0.04025
R11586 VSS.n7519 VSS.n2060 0.04025
R11587 VSS.n7515 VSS.n2060 0.04025
R11588 VSS.n7515 VSS.n7514 0.04025
R11589 VSS.n7514 VSS.n7513 0.04025
R11590 VSS.n7513 VSS.n2062 0.04025
R11591 VSS.n7509 VSS.n2062 0.04025
R11592 VSS.n7509 VSS.n7508 0.04025
R11593 VSS.n7508 VSS.n7507 0.04025
R11594 VSS.n7507 VSS.n2064 0.04025
R11595 VSS.n7503 VSS.n2064 0.04025
R11596 VSS.n7503 VSS.n7502 0.04025
R11597 VSS.n7502 VSS.n7501 0.04025
R11598 VSS.n7501 VSS.n2066 0.04025
R11599 VSS.n7497 VSS.n2066 0.04025
R11600 VSS.n7497 VSS.n7496 0.04025
R11601 VSS.n7496 VSS.n7495 0.04025
R11602 VSS.n7495 VSS.n2068 0.04025
R11603 VSS.n7491 VSS.n2068 0.04025
R11604 VSS.n7491 VSS.n7490 0.04025
R11605 VSS.n7490 VSS.n7489 0.04025
R11606 VSS.n7489 VSS.n2070 0.04025
R11607 VSS.n7485 VSS.n2070 0.04025
R11608 VSS.n7485 VSS.n7484 0.04025
R11609 VSS.n7484 VSS.n7483 0.04025
R11610 VSS.n7483 VSS.n2072 0.04025
R11611 VSS.n7479 VSS.n2072 0.04025
R11612 VSS.n7479 VSS.n7478 0.04025
R11613 VSS.n7478 VSS.n7477 0.04025
R11614 VSS.n7477 VSS.n2074 0.04025
R11615 VSS.n7473 VSS.n2074 0.04025
R11616 VSS.n7473 VSS.n7472 0.04025
R11617 VSS.n7472 VSS.n7471 0.04025
R11618 VSS.n7471 VSS.n2076 0.04025
R11619 VSS.n7467 VSS.n2076 0.04025
R11620 VSS.n7467 VSS.n7466 0.04025
R11621 VSS.n7466 VSS.n7465 0.04025
R11622 VSS.n7465 VSS.n2078 0.04025
R11623 VSS.n7461 VSS.n2078 0.04025
R11624 VSS.n7461 VSS.n7460 0.04025
R11625 VSS.n7460 VSS.n7459 0.04025
R11626 VSS.n7459 VSS.n2080 0.04025
R11627 VSS.n7455 VSS.n2080 0.04025
R11628 VSS.n7455 VSS.n7454 0.04025
R11629 VSS.n7454 VSS.n7453 0.04025
R11630 VSS.n7453 VSS.n2082 0.04025
R11631 VSS.n7449 VSS.n2082 0.04025
R11632 VSS.n7449 VSS.n7448 0.04025
R11633 VSS.n7448 VSS.n7447 0.04025
R11634 VSS.n7447 VSS.n2084 0.04025
R11635 VSS.n7443 VSS.n2084 0.04025
R11636 VSS.n7443 VSS.n7442 0.04025
R11637 VSS.n7442 VSS.n7441 0.04025
R11638 VSS.n7441 VSS.n2086 0.04025
R11639 VSS.n7437 VSS.n2086 0.04025
R11640 VSS.n7437 VSS.n7436 0.04025
R11641 VSS.n7436 VSS.n7435 0.04025
R11642 VSS.n7435 VSS.n2088 0.04025
R11643 VSS.n7431 VSS.n2088 0.04025
R11644 VSS.n7431 VSS.n7430 0.04025
R11645 VSS.n7430 VSS.n7429 0.04025
R11646 VSS.n7429 VSS.n2090 0.04025
R11647 VSS.n7425 VSS.n2090 0.04025
R11648 VSS.n7425 VSS.n7424 0.04025
R11649 VSS.n7424 VSS.n7423 0.04025
R11650 VSS.n7423 VSS.n2092 0.04025
R11651 VSS.n7419 VSS.n2092 0.04025
R11652 VSS.n7419 VSS.n7418 0.04025
R11653 VSS.n7418 VSS.n7417 0.04025
R11654 VSS.n7417 VSS.n2094 0.04025
R11655 VSS.n7413 VSS.n2094 0.04025
R11656 VSS.n7413 VSS.n7412 0.04025
R11657 VSS.n7412 VSS.n7411 0.04025
R11658 VSS.n7411 VSS.n2096 0.04025
R11659 VSS.n7407 VSS.n2096 0.04025
R11660 VSS.n7407 VSS.n7406 0.04025
R11661 VSS.n7406 VSS.n7405 0.04025
R11662 VSS.n7405 VSS.n2098 0.04025
R11663 VSS.n7401 VSS.n2098 0.04025
R11664 VSS.n7401 VSS.n7400 0.04025
R11665 VSS.n7400 VSS.n7399 0.04025
R11666 VSS.n7399 VSS.n2100 0.04025
R11667 VSS.n7395 VSS.n2100 0.04025
R11668 VSS.n7395 VSS.n7394 0.04025
R11669 VSS.n7394 VSS.n7393 0.04025
R11670 VSS.n7393 VSS.n2102 0.04025
R11671 VSS.n7389 VSS.n2102 0.04025
R11672 VSS.n7389 VSS.n7388 0.04025
R11673 VSS.n7388 VSS.n7387 0.04025
R11674 VSS.n7387 VSS.n2104 0.04025
R11675 VSS.n7383 VSS.n2104 0.04025
R11676 VSS.n7383 VSS.n7382 0.04025
R11677 VSS.n7382 VSS.n7381 0.04025
R11678 VSS.n7381 VSS.n2106 0.04025
R11679 VSS.n7377 VSS.n2106 0.04025
R11680 VSS.n7377 VSS.n7376 0.04025
R11681 VSS.n7376 VSS.n7375 0.04025
R11682 VSS.n7375 VSS.n2108 0.04025
R11683 VSS.n7371 VSS.n2108 0.04025
R11684 VSS.n7371 VSS.n7370 0.04025
R11685 VSS.n7370 VSS.n7369 0.04025
R11686 VSS.n7369 VSS.n2110 0.04025
R11687 VSS.n7365 VSS.n2110 0.04025
R11688 VSS.n7365 VSS.n7364 0.04025
R11689 VSS.n7364 VSS.n7363 0.04025
R11690 VSS.n7363 VSS.n2112 0.04025
R11691 VSS.n7359 VSS.n2112 0.04025
R11692 VSS.n7359 VSS.n7358 0.04025
R11693 VSS.n7358 VSS.n7357 0.04025
R11694 VSS.n7357 VSS.n2114 0.04025
R11695 VSS.n7353 VSS.n2114 0.04025
R11696 VSS.n7353 VSS.n7352 0.04025
R11697 VSS.n7352 VSS.n7351 0.04025
R11698 VSS.n7351 VSS.n2116 0.04025
R11699 VSS.n7347 VSS.n2116 0.04025
R11700 VSS.n7347 VSS.n7346 0.04025
R11701 VSS.n7346 VSS.n7345 0.04025
R11702 VSS.n7345 VSS.n2118 0.04025
R11703 VSS.n7341 VSS.n2118 0.04025
R11704 VSS.n7341 VSS.n7340 0.04025
R11705 VSS.n7340 VSS.n7339 0.04025
R11706 VSS.n7339 VSS.n2120 0.04025
R11707 VSS.n7335 VSS.n2120 0.04025
R11708 VSS.n7335 VSS.n7334 0.04025
R11709 VSS.n7334 VSS.n7333 0.04025
R11710 VSS.n7333 VSS.n2122 0.04025
R11711 VSS.n7329 VSS.n2122 0.04025
R11712 VSS.n7329 VSS.n7328 0.04025
R11713 VSS.n7328 VSS.n7327 0.04025
R11714 VSS.n7327 VSS.n2124 0.04025
R11715 VSS.n7323 VSS.n2124 0.04025
R11716 VSS.n7323 VSS.n7322 0.04025
R11717 VSS.n7322 VSS.n7321 0.04025
R11718 VSS.n7321 VSS.n2126 0.04025
R11719 VSS.n7317 VSS.n2126 0.04025
R11720 VSS.n7317 VSS.n7316 0.04025
R11721 VSS.n7316 VSS.n7315 0.04025
R11722 VSS.n7315 VSS.n2128 0.04025
R11723 VSS.n7311 VSS.n2128 0.04025
R11724 VSS.n7311 VSS.n7310 0.04025
R11725 VSS.n7310 VSS.n7309 0.04025
R11726 VSS.n7309 VSS.n2130 0.04025
R11727 VSS.n7305 VSS.n2130 0.04025
R11728 VSS.n7305 VSS.n7304 0.04025
R11729 VSS.n7304 VSS.n7303 0.04025
R11730 VSS.n7303 VSS.n2132 0.04025
R11731 VSS.n7299 VSS.n2132 0.04025
R11732 VSS.n7299 VSS.n7298 0.04025
R11733 VSS.n7298 VSS.n7297 0.04025
R11734 VSS.n7297 VSS.n2134 0.04025
R11735 VSS.n7293 VSS.n2134 0.04025
R11736 VSS.n7293 VSS.n7292 0.04025
R11737 VSS.n7292 VSS.n7291 0.04025
R11738 VSS.n7291 VSS.n2136 0.04025
R11739 VSS.n7287 VSS.n2136 0.04025
R11740 VSS.n7287 VSS.n7286 0.04025
R11741 VSS.n7286 VSS.n7285 0.04025
R11742 VSS.n7285 VSS.n2138 0.04025
R11743 VSS.n7281 VSS.n2138 0.04025
R11744 VSS.n7281 VSS.n7280 0.04025
R11745 VSS.n7280 VSS.n7279 0.04025
R11746 VSS.n7279 VSS.n2140 0.04025
R11747 VSS.n7275 VSS.n2140 0.04025
R11748 VSS.n7275 VSS.n7274 0.04025
R11749 VSS.n7274 VSS.n7273 0.04025
R11750 VSS.n7273 VSS.n2142 0.04025
R11751 VSS.n7269 VSS.n2142 0.04025
R11752 VSS.n7269 VSS.n7268 0.04025
R11753 VSS.n7268 VSS.n7267 0.04025
R11754 VSS.n7267 VSS.n2144 0.04025
R11755 VSS.n7263 VSS.n2144 0.04025
R11756 VSS.n7263 VSS.n7262 0.04025
R11757 VSS.n7262 VSS.n7261 0.04025
R11758 VSS.n7261 VSS.n2146 0.04025
R11759 VSS.n7257 VSS.n2146 0.04025
R11760 VSS.n7257 VSS.n7256 0.04025
R11761 VSS.n7256 VSS.n7255 0.04025
R11762 VSS.n7255 VSS.n2148 0.04025
R11763 VSS.n7251 VSS.n2148 0.04025
R11764 VSS.n7251 VSS.n7250 0.04025
R11765 VSS.n7250 VSS.n7249 0.04025
R11766 VSS.n7249 VSS.n2150 0.04025
R11767 VSS.n7245 VSS.n2150 0.04025
R11768 VSS.n7245 VSS.n7244 0.04025
R11769 VSS.n7244 VSS.n7243 0.04025
R11770 VSS.n7243 VSS.n2152 0.04025
R11771 VSS.n7239 VSS.n2152 0.04025
R11772 VSS.n7239 VSS.n7238 0.04025
R11773 VSS.n7238 VSS.n7237 0.04025
R11774 VSS.n7237 VSS.n2154 0.04025
R11775 VSS.n7233 VSS.n2154 0.04025
R11776 VSS.n7233 VSS.n7232 0.04025
R11777 VSS.n7232 VSS.n7231 0.04025
R11778 VSS.n7231 VSS.n2156 0.04025
R11779 VSS.n7227 VSS.n2156 0.04025
R11780 VSS.n7227 VSS.n7226 0.04025
R11781 VSS.n7226 VSS.n7225 0.04025
R11782 VSS.n7225 VSS.n2158 0.04025
R11783 VSS.n7221 VSS.n2158 0.04025
R11784 VSS.n7221 VSS.n7220 0.04025
R11785 VSS.n7220 VSS.n7219 0.04025
R11786 VSS.n7219 VSS.n2160 0.04025
R11787 VSS.n7215 VSS.n2160 0.04025
R11788 VSS.n7215 VSS.n7214 0.04025
R11789 VSS.n7214 VSS.n7213 0.04025
R11790 VSS.n7213 VSS.n2162 0.04025
R11791 VSS.n7209 VSS.n2162 0.04025
R11792 VSS.n7209 VSS.n7208 0.04025
R11793 VSS.n7208 VSS.n7207 0.04025
R11794 VSS.n7207 VSS.n2164 0.04025
R11795 VSS.n7203 VSS.n2164 0.04025
R11796 VSS.n7203 VSS.n7202 0.04025
R11797 VSS.n7202 VSS.n7201 0.04025
R11798 VSS.n7201 VSS.n2166 0.04025
R11799 VSS.n7197 VSS.n2166 0.04025
R11800 VSS.n7197 VSS.n7196 0.04025
R11801 VSS.n7196 VSS.n7195 0.04025
R11802 VSS.n7195 VSS.n2168 0.04025
R11803 VSS.n7191 VSS.n2168 0.04025
R11804 VSS.n7191 VSS.n7190 0.04025
R11805 VSS.n7190 VSS.n7189 0.04025
R11806 VSS.n7189 VSS.n2170 0.04025
R11807 VSS.n7185 VSS.n2170 0.04025
R11808 VSS.n7185 VSS.n7184 0.04025
R11809 VSS.n7184 VSS.n7183 0.04025
R11810 VSS.n7183 VSS.n2172 0.04025
R11811 VSS.n7179 VSS.n2172 0.04025
R11812 VSS.n7179 VSS.n7178 0.04025
R11813 VSS.n7178 VSS.n7177 0.04025
R11814 VSS.n7177 VSS.n2174 0.04025
R11815 VSS.n7173 VSS.n2174 0.04025
R11816 VSS.n7173 VSS.n7172 0.04025
R11817 VSS.n7172 VSS.n7171 0.04025
R11818 VSS.n7171 VSS.n2176 0.04025
R11819 VSS.n7167 VSS.n2176 0.04025
R11820 VSS.n7167 VSS.n7166 0.04025
R11821 VSS.n7166 VSS.n7165 0.04025
R11822 VSS.n7165 VSS.n2178 0.04025
R11823 VSS.n7161 VSS.n2178 0.04025
R11824 VSS.n7161 VSS.n7160 0.04025
R11825 VSS.n7160 VSS.n7159 0.04025
R11826 VSS.n7159 VSS.n2180 0.04025
R11827 VSS.n7155 VSS.n2180 0.04025
R11828 VSS.n7155 VSS.n7154 0.04025
R11829 VSS.n7154 VSS.n7153 0.04025
R11830 VSS.n7153 VSS.n2182 0.04025
R11831 VSS.n7149 VSS.n2182 0.04025
R11832 VSS.n7149 VSS.n7148 0.04025
R11833 VSS.n7148 VSS.n7147 0.04025
R11834 VSS.n7147 VSS.n2184 0.04025
R11835 VSS.n7143 VSS.n2184 0.04025
R11836 VSS.n7143 VSS.n7142 0.04025
R11837 VSS.n7142 VSS.n7141 0.04025
R11838 VSS.n7141 VSS.n2186 0.04025
R11839 VSS.n7137 VSS.n2186 0.04025
R11840 VSS.n7137 VSS.n7136 0.04025
R11841 VSS.n7136 VSS.n7135 0.04025
R11842 VSS.n7135 VSS.n2188 0.04025
R11843 VSS.n7131 VSS.n2188 0.04025
R11844 VSS.n7131 VSS.n7130 0.04025
R11845 VSS.n7130 VSS.n7129 0.04025
R11846 VSS.n7129 VSS.n2190 0.04025
R11847 VSS.n7125 VSS.n2190 0.04025
R11848 VSS.n7125 VSS.n7124 0.04025
R11849 VSS.n7124 VSS.n7123 0.04025
R11850 VSS.n7123 VSS.n2192 0.04025
R11851 VSS.n7119 VSS.n2192 0.04025
R11852 VSS.n7119 VSS.n7118 0.04025
R11853 VSS.n7118 VSS.n7117 0.04025
R11854 VSS.n7117 VSS.n2194 0.04025
R11855 VSS.n7113 VSS.n2194 0.04025
R11856 VSS.n7113 VSS.n7112 0.04025
R11857 VSS.n7112 VSS.n7111 0.04025
R11858 VSS.n7111 VSS.n2196 0.04025
R11859 VSS.n7107 VSS.n2196 0.04025
R11860 VSS.n7107 VSS.n7106 0.04025
R11861 VSS.n7106 VSS.n7105 0.04025
R11862 VSS.n7105 VSS.n2198 0.04025
R11863 VSS.n7101 VSS.n2198 0.04025
R11864 VSS.n7101 VSS.n7100 0.04025
R11865 VSS.n7100 VSS.n7099 0.04025
R11866 VSS.n7099 VSS.n2200 0.04025
R11867 VSS.n7095 VSS.n2200 0.04025
R11868 VSS.n7095 VSS.n7094 0.04025
R11869 VSS.n7094 VSS.n7093 0.04025
R11870 VSS.n7093 VSS.n2202 0.04025
R11871 VSS.n7089 VSS.n2202 0.04025
R11872 VSS.n7089 VSS.n7088 0.04025
R11873 VSS.n7088 VSS.n7087 0.04025
R11874 VSS.n7087 VSS.n2204 0.04025
R11875 VSS.n7083 VSS.n2204 0.04025
R11876 VSS.n7083 VSS.n7082 0.04025
R11877 VSS.n7082 VSS.n7081 0.04025
R11878 VSS.n7081 VSS.n2206 0.04025
R11879 VSS.n7077 VSS.n2206 0.04025
R11880 VSS.n7077 VSS.n7076 0.04025
R11881 VSS.n7076 VSS.n7075 0.04025
R11882 VSS.n7075 VSS.n2208 0.04025
R11883 VSS.n7071 VSS.n2208 0.04025
R11884 VSS.n7071 VSS.n7070 0.04025
R11885 VSS.n7070 VSS.n7069 0.04025
R11886 VSS.n7069 VSS.n2210 0.04025
R11887 VSS.n7065 VSS.n2210 0.04025
R11888 VSS.n7065 VSS.n7064 0.04025
R11889 VSS.n7064 VSS.n7063 0.04025
R11890 VSS.n7063 VSS.n2212 0.04025
R11891 VSS.n7059 VSS.n2212 0.04025
R11892 VSS.n7059 VSS.n7058 0.04025
R11893 VSS.n7058 VSS.n7057 0.04025
R11894 VSS.n7057 VSS.n2214 0.04025
R11895 VSS.n7053 VSS.n2214 0.04025
R11896 VSS.n7053 VSS.n7052 0.04025
R11897 VSS.n7052 VSS.n7051 0.04025
R11898 VSS.n7051 VSS.n2216 0.04025
R11899 VSS.n7047 VSS.n2216 0.04025
R11900 VSS.n7047 VSS.n7046 0.04025
R11901 VSS.n7046 VSS.n7045 0.04025
R11902 VSS.n7045 VSS.n2218 0.04025
R11903 VSS.n7041 VSS.n2218 0.04025
R11904 VSS.n7041 VSS.n7040 0.04025
R11905 VSS.n7040 VSS.n7039 0.04025
R11906 VSS.n7039 VSS.n2220 0.04025
R11907 VSS.n7035 VSS.n2220 0.04025
R11908 VSS.n7035 VSS.n7034 0.04025
R11909 VSS.n7034 VSS.n7033 0.04025
R11910 VSS.n7033 VSS.n2222 0.04025
R11911 VSS.n7029 VSS.n2222 0.04025
R11912 VSS.n7029 VSS.n7028 0.04025
R11913 VSS.n7028 VSS.n7027 0.04025
R11914 VSS.n7027 VSS.n2224 0.04025
R11915 VSS.n7023 VSS.n2224 0.04025
R11916 VSS.n7023 VSS.n7022 0.04025
R11917 VSS.n7022 VSS.n7021 0.04025
R11918 VSS.n7021 VSS.n2226 0.04025
R11919 VSS.n7017 VSS.n2226 0.04025
R11920 VSS.n7017 VSS.n7016 0.04025
R11921 VSS.n7016 VSS.n7015 0.04025
R11922 VSS.n7015 VSS.n2228 0.04025
R11923 VSS.n7011 VSS.n2228 0.04025
R11924 VSS.n7011 VSS.n7010 0.04025
R11925 VSS.n7010 VSS.n7009 0.04025
R11926 VSS.n7009 VSS.n2230 0.04025
R11927 VSS.n7005 VSS.n2230 0.04025
R11928 VSS.n7005 VSS.n7004 0.04025
R11929 VSS.n7004 VSS.n7003 0.04025
R11930 VSS.n7003 VSS.n2232 0.04025
R11931 VSS.n6999 VSS.n2232 0.04025
R11932 VSS.n6999 VSS.n6998 0.04025
R11933 VSS.n6998 VSS.n6997 0.04025
R11934 VSS.n6997 VSS.n2234 0.04025
R11935 VSS.n6993 VSS.n2234 0.04025
R11936 VSS.n6993 VSS.n6992 0.04025
R11937 VSS.n6992 VSS.n6991 0.04025
R11938 VSS.n6991 VSS.n2236 0.04025
R11939 VSS.n6987 VSS.n2236 0.04025
R11940 VSS.n6987 VSS.n6986 0.04025
R11941 VSS.n6986 VSS.n6985 0.04025
R11942 VSS.n6985 VSS.n2238 0.04025
R11943 VSS.n6981 VSS.n2238 0.04025
R11944 VSS.n6981 VSS.n6980 0.04025
R11945 VSS.n6980 VSS.n6979 0.04025
R11946 VSS.n6979 VSS.n2240 0.04025
R11947 VSS.n6975 VSS.n2240 0.04025
R11948 VSS.n6975 VSS.n6974 0.04025
R11949 VSS.n6974 VSS.n6973 0.04025
R11950 VSS.n6973 VSS.n2242 0.04025
R11951 VSS.n6969 VSS.n2242 0.04025
R11952 VSS.n6969 VSS.n6968 0.04025
R11953 VSS.n6968 VSS.n6967 0.04025
R11954 VSS.n6967 VSS.n2244 0.04025
R11955 VSS.n6963 VSS.n2244 0.04025
R11956 VSS.n6963 VSS.n6962 0.04025
R11957 VSS.n6962 VSS.n6961 0.04025
R11958 VSS.n6961 VSS.n2246 0.04025
R11959 VSS.n6957 VSS.n2246 0.04025
R11960 VSS.n6957 VSS.n6956 0.04025
R11961 VSS.n6956 VSS.n6955 0.04025
R11962 VSS.n6955 VSS.n2248 0.04025
R11963 VSS.n6951 VSS.n2248 0.04025
R11964 VSS.n6951 VSS.n6950 0.04025
R11965 VSS.n6950 VSS.n6949 0.04025
R11966 VSS.n6949 VSS.n2250 0.04025
R11967 VSS.n6945 VSS.n2250 0.04025
R11968 VSS.n6945 VSS.n6944 0.04025
R11969 VSS.n6944 VSS.n6943 0.04025
R11970 VSS.n6943 VSS.n2252 0.04025
R11971 VSS.n6939 VSS.n2252 0.04025
R11972 VSS.n6939 VSS.n6938 0.04025
R11973 VSS.n6938 VSS.n6937 0.04025
R11974 VSS.n6937 VSS.n2254 0.04025
R11975 VSS.n6933 VSS.n2254 0.04025
R11976 VSS.n6933 VSS.n6932 0.04025
R11977 VSS.n6932 VSS.n6931 0.04025
R11978 VSS.n6931 VSS.n2256 0.04025
R11979 VSS.n6927 VSS.n2256 0.04025
R11980 VSS.n6927 VSS.n6926 0.04025
R11981 VSS.n6926 VSS.n6925 0.04025
R11982 VSS.n6925 VSS.n2258 0.04025
R11983 VSS.n6921 VSS.n2258 0.04025
R11984 VSS.n6921 VSS.n6920 0.04025
R11985 VSS.n6920 VSS.n6919 0.04025
R11986 VSS.n6919 VSS.n2260 0.04025
R11987 VSS.n6915 VSS.n2260 0.04025
R11988 VSS.n6915 VSS.n6914 0.04025
R11989 VSS.n6914 VSS.n6913 0.04025
R11990 VSS.n6913 VSS.n2262 0.04025
R11991 VSS.n6909 VSS.n2262 0.04025
R11992 VSS.n6909 VSS.n6908 0.04025
R11993 VSS.n4140 VSS.n4139 0.04025
R11994 VSS.n4139 VSS.n4138 0.04025
R11995 VSS.n4138 VSS.n3186 0.04025
R11996 VSS.n4134 VSS.n3186 0.04025
R11997 VSS.n4134 VSS.n4133 0.04025
R11998 VSS.n4133 VSS.n4132 0.04025
R11999 VSS.n4132 VSS.n3188 0.04025
R12000 VSS.n4128 VSS.n3188 0.04025
R12001 VSS.n4128 VSS.n4127 0.04025
R12002 VSS.n4127 VSS.n4126 0.04025
R12003 VSS.n4126 VSS.n3190 0.04025
R12004 VSS.n4122 VSS.n3190 0.04025
R12005 VSS.n4122 VSS.n4121 0.04025
R12006 VSS.n4121 VSS.n4120 0.04025
R12007 VSS.n4120 VSS.n3192 0.04025
R12008 VSS.n4116 VSS.n3192 0.04025
R12009 VSS.n4116 VSS.n4115 0.04025
R12010 VSS.n4115 VSS.n4114 0.04025
R12011 VSS.n4114 VSS.n3194 0.04025
R12012 VSS.n4110 VSS.n3194 0.04025
R12013 VSS.n4110 VSS.n4109 0.04025
R12014 VSS.n4109 VSS.n4108 0.04025
R12015 VSS.n4108 VSS.n3196 0.04025
R12016 VSS.n4104 VSS.n3196 0.04025
R12017 VSS.n4104 VSS.n4103 0.04025
R12018 VSS.n4103 VSS.n4102 0.04025
R12019 VSS.n4102 VSS.n3198 0.04025
R12020 VSS.n4098 VSS.n3198 0.04025
R12021 VSS.n4098 VSS.n4097 0.04025
R12022 VSS.n4097 VSS.n4096 0.04025
R12023 VSS.n4096 VSS.n3200 0.04025
R12024 VSS.n4092 VSS.n3200 0.04025
R12025 VSS.n4092 VSS.n4091 0.04025
R12026 VSS.n4091 VSS.n4090 0.04025
R12027 VSS.n4090 VSS.n3202 0.04025
R12028 VSS.n4086 VSS.n3202 0.04025
R12029 VSS.n4086 VSS.n4085 0.04025
R12030 VSS.n4085 VSS.n4084 0.04025
R12031 VSS.n4084 VSS.n3204 0.04025
R12032 VSS.n4080 VSS.n3204 0.04025
R12033 VSS.n4080 VSS.n4079 0.04025
R12034 VSS.n4079 VSS.n4078 0.04025
R12035 VSS.n4078 VSS.n3206 0.04025
R12036 VSS.n4074 VSS.n3206 0.04025
R12037 VSS.n4074 VSS.n4073 0.04025
R12038 VSS.n4073 VSS.n4072 0.04025
R12039 VSS.n4072 VSS.n3208 0.04025
R12040 VSS.n4068 VSS.n3208 0.04025
R12041 VSS.n4068 VSS.n4067 0.04025
R12042 VSS.n4067 VSS.n4066 0.04025
R12043 VSS.n4066 VSS.n3210 0.04025
R12044 VSS.n4062 VSS.n3210 0.04025
R12045 VSS.n4062 VSS.n4061 0.04025
R12046 VSS.n4061 VSS.n4060 0.04025
R12047 VSS.n4060 VSS.n3212 0.04025
R12048 VSS.n4056 VSS.n3212 0.04025
R12049 VSS.n4056 VSS.n4055 0.04025
R12050 VSS.n4055 VSS.n4054 0.04025
R12051 VSS.n4054 VSS.n3214 0.04025
R12052 VSS.n4050 VSS.n3214 0.04025
R12053 VSS.n4050 VSS.n4049 0.04025
R12054 VSS.n4049 VSS.n4048 0.04025
R12055 VSS.n4048 VSS.n3216 0.04025
R12056 VSS.n4044 VSS.n3216 0.04025
R12057 VSS.n4044 VSS.n4043 0.04025
R12058 VSS.n4043 VSS.n4042 0.04025
R12059 VSS.n4042 VSS.n3218 0.04025
R12060 VSS.n4038 VSS.n3218 0.04025
R12061 VSS.n4038 VSS.n4037 0.04025
R12062 VSS.n4037 VSS.n4036 0.04025
R12063 VSS.n4036 VSS.n3220 0.04025
R12064 VSS.n4032 VSS.n3220 0.04025
R12065 VSS.n4032 VSS.n4031 0.04025
R12066 VSS.n4031 VSS.n4030 0.04025
R12067 VSS.n4030 VSS.n3222 0.04025
R12068 VSS.n4026 VSS.n3222 0.04025
R12069 VSS.n4026 VSS.n4025 0.04025
R12070 VSS.n4025 VSS.n4024 0.04025
R12071 VSS.n4024 VSS.n3224 0.04025
R12072 VSS.n4020 VSS.n3224 0.04025
R12073 VSS.n4020 VSS.n4019 0.04025
R12074 VSS.n4019 VSS.n4018 0.04025
R12075 VSS.n4018 VSS.n3226 0.04025
R12076 VSS.n4014 VSS.n3226 0.04025
R12077 VSS.n4014 VSS.n4013 0.04025
R12078 VSS.n4013 VSS.n4012 0.04025
R12079 VSS.n4012 VSS.n3228 0.04025
R12080 VSS.n4008 VSS.n3228 0.04025
R12081 VSS.n4008 VSS.n4007 0.04025
R12082 VSS.n4007 VSS.n4006 0.04025
R12083 VSS.n4006 VSS.n3230 0.04025
R12084 VSS.n4002 VSS.n3230 0.04025
R12085 VSS.n4002 VSS.n4001 0.04025
R12086 VSS.n4001 VSS.n4000 0.04025
R12087 VSS.n4000 VSS.n3232 0.04025
R12088 VSS.n3996 VSS.n3232 0.04025
R12089 VSS.n3996 VSS.n3995 0.04025
R12090 VSS.n3995 VSS.n3994 0.04025
R12091 VSS.n3994 VSS.n3234 0.04025
R12092 VSS.n3990 VSS.n3234 0.04025
R12093 VSS.n3990 VSS.n3989 0.04025
R12094 VSS.n3989 VSS.n3988 0.04025
R12095 VSS.n3988 VSS.n3236 0.04025
R12096 VSS.n3984 VSS.n3236 0.04025
R12097 VSS.n3984 VSS.n3983 0.04025
R12098 VSS.n3983 VSS.n3982 0.04025
R12099 VSS.n3982 VSS.n3238 0.04025
R12100 VSS.n3978 VSS.n3238 0.04025
R12101 VSS.n3978 VSS.n3977 0.04025
R12102 VSS.n3977 VSS.n3976 0.04025
R12103 VSS.n3976 VSS.n3240 0.04025
R12104 VSS.n3972 VSS.n3240 0.04025
R12105 VSS.n3972 VSS.n3971 0.04025
R12106 VSS.n3971 VSS.n3970 0.04025
R12107 VSS.n3970 VSS.n3242 0.04025
R12108 VSS.n3966 VSS.n3242 0.04025
R12109 VSS.n3966 VSS.n3965 0.04025
R12110 VSS.n3965 VSS.n3964 0.04025
R12111 VSS.n3964 VSS.n3244 0.04025
R12112 VSS.n3960 VSS.n3244 0.04025
R12113 VSS.n3960 VSS.n3959 0.04025
R12114 VSS.n3959 VSS.n3958 0.04025
R12115 VSS.n3958 VSS.n3246 0.04025
R12116 VSS.n3954 VSS.n3246 0.04025
R12117 VSS.n3954 VSS.n3953 0.04025
R12118 VSS.n3953 VSS.n3952 0.04025
R12119 VSS.n3952 VSS.n3248 0.04025
R12120 VSS.n3948 VSS.n3248 0.04025
R12121 VSS.n3948 VSS.n3947 0.04025
R12122 VSS.n3947 VSS.n3946 0.04025
R12123 VSS.n3946 VSS.n3250 0.04025
R12124 VSS.n3942 VSS.n3250 0.04025
R12125 VSS.n3942 VSS.n3941 0.04025
R12126 VSS.n3941 VSS.n3940 0.04025
R12127 VSS.n3940 VSS.n3252 0.04025
R12128 VSS.n3936 VSS.n3252 0.04025
R12129 VSS.n3936 VSS.n3935 0.04025
R12130 VSS.n3935 VSS.n3934 0.04025
R12131 VSS.n3934 VSS.n3254 0.04025
R12132 VSS.n3930 VSS.n3254 0.04025
R12133 VSS.n3930 VSS.n3929 0.04025
R12134 VSS.n3929 VSS.n3928 0.04025
R12135 VSS.n3928 VSS.n3256 0.04025
R12136 VSS.n3924 VSS.n3256 0.04025
R12137 VSS.n3924 VSS.n3923 0.04025
R12138 VSS.n3923 VSS.n3922 0.04025
R12139 VSS.n3922 VSS.n3258 0.04025
R12140 VSS.n3918 VSS.n3258 0.04025
R12141 VSS.n3918 VSS.n3917 0.04025
R12142 VSS.n3917 VSS.n3916 0.04025
R12143 VSS.n3916 VSS.n3260 0.04025
R12144 VSS.n3912 VSS.n3260 0.04025
R12145 VSS.n3912 VSS.n3911 0.04025
R12146 VSS.n3911 VSS.n3910 0.04025
R12147 VSS.n3910 VSS.n3262 0.04025
R12148 VSS.n3906 VSS.n3262 0.04025
R12149 VSS.n3906 VSS.n3905 0.04025
R12150 VSS.n3905 VSS.n3904 0.04025
R12151 VSS.n3904 VSS.n3264 0.04025
R12152 VSS.n3900 VSS.n3264 0.04025
R12153 VSS.n3900 VSS.n3899 0.04025
R12154 VSS.n3899 VSS.n3898 0.04025
R12155 VSS.n3898 VSS.n3266 0.04025
R12156 VSS.n3894 VSS.n3266 0.04025
R12157 VSS.n3894 VSS.n3893 0.04025
R12158 VSS.n3893 VSS.n3892 0.04025
R12159 VSS.n3892 VSS.n3268 0.04025
R12160 VSS.n3888 VSS.n3268 0.04025
R12161 VSS.n3888 VSS.n3887 0.04025
R12162 VSS.n3887 VSS.n3886 0.04025
R12163 VSS.n3886 VSS.n3270 0.04025
R12164 VSS.n3882 VSS.n3270 0.04025
R12165 VSS.n3882 VSS.n3881 0.04025
R12166 VSS.n3881 VSS.n3880 0.04025
R12167 VSS.n3880 VSS.n3272 0.04025
R12168 VSS.n3876 VSS.n3272 0.04025
R12169 VSS.n3876 VSS.n3875 0.04025
R12170 VSS.n3875 VSS.n3874 0.04025
R12171 VSS.n3874 VSS.n3274 0.04025
R12172 VSS.n3870 VSS.n3274 0.04025
R12173 VSS.n3870 VSS.n3869 0.04025
R12174 VSS.n3869 VSS.n3868 0.04025
R12175 VSS.n3868 VSS.n3276 0.04025
R12176 VSS.n3864 VSS.n3276 0.04025
R12177 VSS.n3864 VSS.n3863 0.04025
R12178 VSS.n3863 VSS.n3862 0.04025
R12179 VSS.n3862 VSS.n3278 0.04025
R12180 VSS.n3858 VSS.n3278 0.04025
R12181 VSS.n3858 VSS.n3857 0.04025
R12182 VSS.n3857 VSS.n3856 0.04025
R12183 VSS.n3856 VSS.n3280 0.04025
R12184 VSS.n3852 VSS.n3280 0.04025
R12185 VSS.n3852 VSS.n3851 0.04025
R12186 VSS.n3851 VSS.n3850 0.04025
R12187 VSS.n3850 VSS.n3282 0.04025
R12188 VSS.n3846 VSS.n3282 0.04025
R12189 VSS.n3846 VSS.n3845 0.04025
R12190 VSS.n3845 VSS.n3844 0.04025
R12191 VSS.n3844 VSS.n3284 0.04025
R12192 VSS.n3840 VSS.n3284 0.04025
R12193 VSS.n3840 VSS.n3839 0.04025
R12194 VSS.n3839 VSS.n3838 0.04025
R12195 VSS.n3838 VSS.n3286 0.04025
R12196 VSS.n3834 VSS.n3286 0.04025
R12197 VSS.n3834 VSS.n3833 0.04025
R12198 VSS.n3833 VSS.n3832 0.04025
R12199 VSS.n3832 VSS.n3288 0.04025
R12200 VSS.n3828 VSS.n3288 0.04025
R12201 VSS.n3828 VSS.n3827 0.04025
R12202 VSS.n3827 VSS.n3826 0.04025
R12203 VSS.n3826 VSS.n3290 0.04025
R12204 VSS.n3822 VSS.n3290 0.04025
R12205 VSS.n3822 VSS.n3821 0.04025
R12206 VSS.n3821 VSS.n3820 0.04025
R12207 VSS.n3820 VSS.n3292 0.04025
R12208 VSS.n3816 VSS.n3292 0.04025
R12209 VSS.n3816 VSS.n3815 0.04025
R12210 VSS.n3815 VSS.n3814 0.04025
R12211 VSS.n3814 VSS.n3294 0.04025
R12212 VSS.n3810 VSS.n3294 0.04025
R12213 VSS.n3810 VSS.n3809 0.04025
R12214 VSS.n3809 VSS.n3808 0.04025
R12215 VSS.n3808 VSS.n3296 0.04025
R12216 VSS.n3804 VSS.n3296 0.04025
R12217 VSS.n3804 VSS.n3803 0.04025
R12218 VSS.n3803 VSS.n3802 0.04025
R12219 VSS.n3802 VSS.n3298 0.04025
R12220 VSS.n3798 VSS.n3298 0.04025
R12221 VSS.n3798 VSS.n3797 0.04025
R12222 VSS.n3797 VSS.n3796 0.04025
R12223 VSS.n3796 VSS.n3300 0.04025
R12224 VSS.n3792 VSS.n3300 0.04025
R12225 VSS.n3792 VSS.n3791 0.04025
R12226 VSS.n3791 VSS.n3790 0.04025
R12227 VSS.n3790 VSS.n3302 0.04025
R12228 VSS.n3786 VSS.n3302 0.04025
R12229 VSS.n3786 VSS.n3785 0.04025
R12230 VSS.n3785 VSS.n3784 0.04025
R12231 VSS.n3784 VSS.n3304 0.04025
R12232 VSS.n3780 VSS.n3304 0.04025
R12233 VSS.n3780 VSS.n3779 0.04025
R12234 VSS.n3779 VSS.n3778 0.04025
R12235 VSS.n3778 VSS.n3306 0.04025
R12236 VSS.n3774 VSS.n3306 0.04025
R12237 VSS.n3774 VSS.n3773 0.04025
R12238 VSS.n3773 VSS.n3772 0.04025
R12239 VSS.n3772 VSS.n3308 0.04025
R12240 VSS.n3768 VSS.n3308 0.04025
R12241 VSS.n3768 VSS.n3767 0.04025
R12242 VSS.n3767 VSS.n3766 0.04025
R12243 VSS.n3766 VSS.n3310 0.04025
R12244 VSS.n3762 VSS.n3310 0.04025
R12245 VSS.n3762 VSS.n3761 0.04025
R12246 VSS.n3761 VSS.n3760 0.04025
R12247 VSS.n3760 VSS.n3312 0.04025
R12248 VSS.n3756 VSS.n3312 0.04025
R12249 VSS.n3756 VSS.n3755 0.04025
R12250 VSS.n3755 VSS.n3754 0.04025
R12251 VSS.n3754 VSS.n3314 0.04025
R12252 VSS.n3750 VSS.n3314 0.04025
R12253 VSS.n3750 VSS.n3749 0.04025
R12254 VSS.n3749 VSS.n3748 0.04025
R12255 VSS.n3748 VSS.n3316 0.04025
R12256 VSS.n3744 VSS.n3316 0.04025
R12257 VSS.n3744 VSS.n3743 0.04025
R12258 VSS.n3743 VSS.n3742 0.04025
R12259 VSS.n3742 VSS.n3318 0.04025
R12260 VSS.n3738 VSS.n3318 0.04025
R12261 VSS.n3738 VSS.n3737 0.04025
R12262 VSS.n3737 VSS.n3736 0.04025
R12263 VSS.n3736 VSS.n3320 0.04025
R12264 VSS.n3732 VSS.n3320 0.04025
R12265 VSS.n3732 VSS.n3731 0.04025
R12266 VSS.n3731 VSS.n3730 0.04025
R12267 VSS.n3730 VSS.n3322 0.04025
R12268 VSS.n3726 VSS.n3322 0.04025
R12269 VSS.n3726 VSS.n3725 0.04025
R12270 VSS.n3725 VSS.n3724 0.04025
R12271 VSS.n3724 VSS.n3324 0.04025
R12272 VSS.n3720 VSS.n3324 0.04025
R12273 VSS.n3720 VSS.n3719 0.04025
R12274 VSS.n3719 VSS.n3718 0.04025
R12275 VSS.n3718 VSS.n3326 0.04025
R12276 VSS.n3714 VSS.n3326 0.04025
R12277 VSS.n3714 VSS.n3713 0.04025
R12278 VSS.n3713 VSS.n3712 0.04025
R12279 VSS.n3712 VSS.n3328 0.04025
R12280 VSS.n3708 VSS.n3328 0.04025
R12281 VSS.n3708 VSS.n3707 0.04025
R12282 VSS.n3707 VSS.n3706 0.04025
R12283 VSS.n3706 VSS.n3330 0.04025
R12284 VSS.n3702 VSS.n3330 0.04025
R12285 VSS.n3702 VSS.n3701 0.04025
R12286 VSS.n3701 VSS.n3700 0.04025
R12287 VSS.n3700 VSS.n3332 0.04025
R12288 VSS.n3696 VSS.n3332 0.04025
R12289 VSS.n3696 VSS.n3695 0.04025
R12290 VSS.n3695 VSS.n3694 0.04025
R12291 VSS.n3694 VSS.n3334 0.04025
R12292 VSS.n3690 VSS.n3334 0.04025
R12293 VSS.n3690 VSS.n3689 0.04025
R12294 VSS.n3689 VSS.n3688 0.04025
R12295 VSS.n3688 VSS.n3336 0.04025
R12296 VSS.n3684 VSS.n3336 0.04025
R12297 VSS.n3684 VSS.n3683 0.04025
R12298 VSS.n3683 VSS.n3682 0.04025
R12299 VSS.n3682 VSS.n3338 0.04025
R12300 VSS.n3678 VSS.n3338 0.04025
R12301 VSS.n3678 VSS.n3677 0.04025
R12302 VSS.n3677 VSS.n3676 0.04025
R12303 VSS.n3676 VSS.n3340 0.04025
R12304 VSS.n3672 VSS.n3340 0.04025
R12305 VSS.n3672 VSS.n3671 0.04025
R12306 VSS.n3671 VSS.n3670 0.04025
R12307 VSS.n3670 VSS.n3342 0.04025
R12308 VSS.n3666 VSS.n3342 0.04025
R12309 VSS.n3666 VSS.n3665 0.04025
R12310 VSS.n3665 VSS.n3664 0.04025
R12311 VSS.n3664 VSS.n3344 0.04025
R12312 VSS.n3660 VSS.n3344 0.04025
R12313 VSS.n3660 VSS.n3659 0.04025
R12314 VSS.n3659 VSS.n3658 0.04025
R12315 VSS.n3658 VSS.n3346 0.04025
R12316 VSS.n3654 VSS.n3346 0.04025
R12317 VSS.n3654 VSS.n3653 0.04025
R12318 VSS.n3653 VSS.n3652 0.04025
R12319 VSS.n3652 VSS.n3348 0.04025
R12320 VSS.n3648 VSS.n3348 0.04025
R12321 VSS.n3648 VSS.n3647 0.04025
R12322 VSS.n3647 VSS.n3646 0.04025
R12323 VSS.n3646 VSS.n3350 0.04025
R12324 VSS.n3642 VSS.n3350 0.04025
R12325 VSS.n3642 VSS.n3641 0.04025
R12326 VSS.n3641 VSS.n3640 0.04025
R12327 VSS.n3640 VSS.n3352 0.04025
R12328 VSS.n3636 VSS.n3352 0.04025
R12329 VSS.n3636 VSS.n3635 0.04025
R12330 VSS.n3635 VSS.n3634 0.04025
R12331 VSS.n3634 VSS.n3354 0.04025
R12332 VSS.n3630 VSS.n3354 0.04025
R12333 VSS.n3630 VSS.n3629 0.04025
R12334 VSS.n3629 VSS.n3628 0.04025
R12335 VSS.n3628 VSS.n3356 0.04025
R12336 VSS.n3624 VSS.n3356 0.04025
R12337 VSS.n3624 VSS.n3623 0.04025
R12338 VSS.n3623 VSS.n3622 0.04025
R12339 VSS.n3622 VSS.n3358 0.04025
R12340 VSS.n3618 VSS.n3358 0.04025
R12341 VSS.n3618 VSS.n3617 0.04025
R12342 VSS.n3617 VSS.n3616 0.04025
R12343 VSS.n3616 VSS.n3360 0.04025
R12344 VSS.n3612 VSS.n3360 0.04025
R12345 VSS.n3612 VSS.n3611 0.04025
R12346 VSS.n3611 VSS.n3610 0.04025
R12347 VSS.n3610 VSS.n3362 0.04025
R12348 VSS.n3606 VSS.n3362 0.04025
R12349 VSS.n3606 VSS.n3605 0.04025
R12350 VSS.n3605 VSS.n3604 0.04025
R12351 VSS.n3604 VSS.n3364 0.04025
R12352 VSS.n3600 VSS.n3364 0.04025
R12353 VSS.n3600 VSS.n3599 0.04025
R12354 VSS.n3599 VSS.n3598 0.04025
R12355 VSS.n3598 VSS.n3366 0.04025
R12356 VSS.n3594 VSS.n3366 0.04025
R12357 VSS.n3594 VSS.n3593 0.04025
R12358 VSS.n3593 VSS.n3592 0.04025
R12359 VSS.n3592 VSS.n3368 0.04025
R12360 VSS.n3588 VSS.n3368 0.04025
R12361 VSS.n3588 VSS.n3587 0.04025
R12362 VSS.n3587 VSS.n3586 0.04025
R12363 VSS.n3586 VSS.n3370 0.04025
R12364 VSS.n3582 VSS.n3370 0.04025
R12365 VSS.n3582 VSS.n3581 0.04025
R12366 VSS.n3581 VSS.n3580 0.04025
R12367 VSS.n3580 VSS.n3372 0.04025
R12368 VSS.n3576 VSS.n3372 0.04025
R12369 VSS.n3576 VSS.n3575 0.04025
R12370 VSS.n3575 VSS.n3574 0.04025
R12371 VSS.n3574 VSS.n3374 0.04025
R12372 VSS.n3570 VSS.n3374 0.04025
R12373 VSS.n3570 VSS.n3569 0.04025
R12374 VSS.n3569 VSS.n3568 0.04025
R12375 VSS.n3568 VSS.n3376 0.04025
R12376 VSS.n3564 VSS.n3376 0.04025
R12377 VSS.n3564 VSS.n3563 0.04025
R12378 VSS.n3563 VSS.n3562 0.04025
R12379 VSS.n3562 VSS.n3378 0.04025
R12380 VSS.n3558 VSS.n3378 0.04025
R12381 VSS.n3558 VSS.n3557 0.04025
R12382 VSS.n3557 VSS.n3556 0.04025
R12383 VSS.n3556 VSS.n3380 0.04025
R12384 VSS.n3552 VSS.n3380 0.04025
R12385 VSS.n3552 VSS.n3551 0.04025
R12386 VSS.n3551 VSS.n3550 0.04025
R12387 VSS.n3550 VSS.n3382 0.04025
R12388 VSS.n3546 VSS.n3382 0.04025
R12389 VSS.n3546 VSS.n3545 0.04025
R12390 VSS.n3545 VSS.n3544 0.04025
R12391 VSS.n3544 VSS.n3384 0.04025
R12392 VSS.n3540 VSS.n3384 0.04025
R12393 VSS.n3540 VSS.n3539 0.04025
R12394 VSS.n3539 VSS.n3538 0.04025
R12395 VSS.n3538 VSS.n3386 0.04025
R12396 VSS.n3534 VSS.n3386 0.04025
R12397 VSS.n3534 VSS.n3533 0.04025
R12398 VSS.n3533 VSS.n3532 0.04025
R12399 VSS.n3532 VSS.n3388 0.04025
R12400 VSS.n3528 VSS.n3388 0.04025
R12401 VSS.n3528 VSS.n3527 0.04025
R12402 VSS.n3527 VSS.n3526 0.04025
R12403 VSS.n3526 VSS.n3390 0.04025
R12404 VSS.n3522 VSS.n3390 0.04025
R12405 VSS.n3522 VSS.n3521 0.04025
R12406 VSS.n3521 VSS.n3520 0.04025
R12407 VSS.n3520 VSS.n3392 0.04025
R12408 VSS.n3516 VSS.n3392 0.04025
R12409 VSS.n3516 VSS.n3515 0.04025
R12410 VSS.n3515 VSS.n3514 0.04025
R12411 VSS.n3514 VSS.n3394 0.04025
R12412 VSS.n3510 VSS.n3394 0.04025
R12413 VSS.n3510 VSS.n3509 0.04025
R12414 VSS.n3509 VSS.n3508 0.04025
R12415 VSS.n3508 VSS.n3396 0.04025
R12416 VSS.n3504 VSS.n3396 0.04025
R12417 VSS.n3504 VSS.n3503 0.04025
R12418 VSS.n3503 VSS.n3502 0.04025
R12419 VSS.n3502 VSS.n3398 0.04025
R12420 VSS.n3498 VSS.n3398 0.04025
R12421 VSS.n3498 VSS.n3497 0.04025
R12422 VSS.n3497 VSS.n3496 0.04025
R12423 VSS.n3496 VSS.n3400 0.04025
R12424 VSS.n3492 VSS.n3400 0.04025
R12425 VSS.n3492 VSS.n3491 0.04025
R12426 VSS.n3491 VSS.n3490 0.04025
R12427 VSS.n3490 VSS.n3402 0.04025
R12428 VSS.n3486 VSS.n3402 0.04025
R12429 VSS.n3486 VSS.n3485 0.04025
R12430 VSS.n3485 VSS.n3484 0.04025
R12431 VSS.n3484 VSS.n3404 0.04025
R12432 VSS.n3480 VSS.n3404 0.04025
R12433 VSS.n3480 VSS.n3479 0.04025
R12434 VSS.n3479 VSS.n3478 0.04025
R12435 VSS.n3478 VSS.n3406 0.04025
R12436 VSS.n3474 VSS.n3406 0.04025
R12437 VSS.n3474 VSS.n3473 0.04025
R12438 VSS.n3473 VSS.n3472 0.04025
R12439 VSS.n3472 VSS.n3408 0.04025
R12440 VSS.n3468 VSS.n3408 0.04025
R12441 VSS.n3468 VSS.n3467 0.04025
R12442 VSS.n3467 VSS.n3466 0.04025
R12443 VSS.n3466 VSS.n3410 0.04025
R12444 VSS.n3462 VSS.n3410 0.04025
R12445 VSS.n3462 VSS.n3461 0.04025
R12446 VSS.n3461 VSS.n3460 0.04025
R12447 VSS.n3460 VSS.n3412 0.04025
R12448 VSS.n3456 VSS.n3412 0.04025
R12449 VSS.n3456 VSS.n3455 0.04025
R12450 VSS.n3455 VSS.n3454 0.04025
R12451 VSS.n3454 VSS.n3414 0.04025
R12452 VSS.n3450 VSS.n3414 0.04025
R12453 VSS.n3450 VSS.n3449 0.04025
R12454 VSS.n3449 VSS.n3448 0.04025
R12455 VSS.n3448 VSS.n3416 0.04025
R12456 VSS.n3444 VSS.n3416 0.04025
R12457 VSS.n3444 VSS.n3443 0.04025
R12458 VSS.n3443 VSS.n3442 0.04025
R12459 VSS.n3442 VSS.n3418 0.04025
R12460 VSS.n3438 VSS.n3418 0.04025
R12461 VSS.n3438 VSS.n3437 0.04025
R12462 VSS.n3437 VSS.n3436 0.04025
R12463 VSS.n3436 VSS.n3420 0.04025
R12464 VSS.n3432 VSS.n3420 0.04025
R12465 VSS.n3432 VSS.n3431 0.04025
R12466 VSS.n3431 VSS.n3430 0.04025
R12467 VSS.n3430 VSS.n3422 0.04025
R12468 VSS.n3426 VSS.n3422 0.04025
R12469 VSS.n3426 VSS.n3425 0.04025
R12470 VSS.n3425 VSS.n3424 0.04025
R12471 VSS.n3424 VSS.n1582 0.04025
R12472 VSS.n8949 VSS.n1582 0.04025
R12473 VSS.n8949 VSS.n8948 0.04025
R12474 VSS.n8948 VSS.n8947 0.04025
R12475 VSS.n8947 VSS.n1584 0.04025
R12476 VSS.n8943 VSS.n1584 0.04025
R12477 VSS.n8943 VSS.n8942 0.04025
R12478 VSS.n8942 VSS.n8941 0.04025
R12479 VSS.n8941 VSS.n1586 0.04025
R12480 VSS.n8937 VSS.n1586 0.04025
R12481 VSS.n8937 VSS.n8936 0.04025
R12482 VSS.n8936 VSS.n8935 0.04025
R12483 VSS.n8935 VSS.n1588 0.04025
R12484 VSS.n8931 VSS.n1588 0.04025
R12485 VSS.n8931 VSS.n8930 0.04025
R12486 VSS.n8930 VSS.n8929 0.04025
R12487 VSS.n8929 VSS.n1590 0.04025
R12488 VSS.n8925 VSS.n1590 0.04025
R12489 VSS.n8925 VSS.n8924 0.04025
R12490 VSS.n8924 VSS.n8923 0.04025
R12491 VSS.n8923 VSS.n1592 0.04025
R12492 VSS.n8919 VSS.n1592 0.04025
R12493 VSS.n8919 VSS.n8918 0.04025
R12494 VSS.n8918 VSS.n8917 0.04025
R12495 VSS.n8917 VSS.n1594 0.04025
R12496 VSS.n8913 VSS.n1594 0.04025
R12497 VSS.n8913 VSS.n8912 0.04025
R12498 VSS.n8912 VSS.n8911 0.04025
R12499 VSS.n8911 VSS.n1596 0.04025
R12500 VSS.n8907 VSS.n1596 0.04025
R12501 VSS.n8907 VSS.n8906 0.04025
R12502 VSS.n8906 VSS.n8905 0.04025
R12503 VSS.n8905 VSS.n1598 0.04025
R12504 VSS.n8901 VSS.n1598 0.04025
R12505 VSS.n8901 VSS.n8900 0.04025
R12506 VSS.n8900 VSS.n8899 0.04025
R12507 VSS.n8899 VSS.n1600 0.04025
R12508 VSS.n8895 VSS.n1600 0.04025
R12509 VSS.n8895 VSS.n8894 0.04025
R12510 VSS.n8894 VSS.n8893 0.04025
R12511 VSS.n8893 VSS.n1602 0.04025
R12512 VSS.n8889 VSS.n1602 0.04025
R12513 VSS.n8889 VSS.n8888 0.04025
R12514 VSS.n8888 VSS.n8887 0.04025
R12515 VSS.n8887 VSS.n1604 0.04025
R12516 VSS.n8883 VSS.n1604 0.04025
R12517 VSS.n8883 VSS.n8882 0.04025
R12518 VSS.n8882 VSS.n8881 0.04025
R12519 VSS.n8881 VSS.n1606 0.04025
R12520 VSS.n8877 VSS.n1606 0.04025
R12521 VSS.n8877 VSS.n8876 0.04025
R12522 VSS.n8876 VSS.n8875 0.04025
R12523 VSS.n8875 VSS.n1608 0.04025
R12524 VSS.n8871 VSS.n1608 0.04025
R12525 VSS.n8871 VSS.n8870 0.04025
R12526 VSS.n8870 VSS.n8869 0.04025
R12527 VSS.n8869 VSS.n1610 0.04025
R12528 VSS.n8865 VSS.n1610 0.04025
R12529 VSS.n8865 VSS.n8864 0.04025
R12530 VSS.n8864 VSS.n8863 0.04025
R12531 VSS.n8863 VSS.n1612 0.04025
R12532 VSS.n8859 VSS.n1612 0.04025
R12533 VSS.n8859 VSS.n8858 0.04025
R12534 VSS.n8858 VSS.n8857 0.04025
R12535 VSS.n8857 VSS.n1614 0.04025
R12536 VSS.n8853 VSS.n1614 0.04025
R12537 VSS.n8853 VSS.n8852 0.04025
R12538 VSS.n8852 VSS.n8851 0.04025
R12539 VSS.n8851 VSS.n1616 0.04025
R12540 VSS.n8847 VSS.n1616 0.04025
R12541 VSS.n8847 VSS.n8846 0.04025
R12542 VSS.n8846 VSS.n8845 0.04025
R12543 VSS.n8845 VSS.n1618 0.04025
R12544 VSS.n8841 VSS.n1618 0.04025
R12545 VSS.n8841 VSS.n8840 0.04025
R12546 VSS.n8840 VSS.n8839 0.04025
R12547 VSS.n8839 VSS.n1620 0.04025
R12548 VSS.n8835 VSS.n1620 0.04025
R12549 VSS.n8835 VSS.n8834 0.04025
R12550 VSS.n8834 VSS.n8833 0.04025
R12551 VSS.n8833 VSS.n1622 0.04025
R12552 VSS.n8829 VSS.n1622 0.04025
R12553 VSS.n8829 VSS.n8828 0.04025
R12554 VSS.n8828 VSS.n8827 0.04025
R12555 VSS.n8827 VSS.n1624 0.04025
R12556 VSS.n8823 VSS.n1624 0.04025
R12557 VSS.n8823 VSS.n8822 0.04025
R12558 VSS.n8822 VSS.n8821 0.04025
R12559 VSS.n8821 VSS.n1626 0.04025
R12560 VSS.n8817 VSS.n1626 0.04025
R12561 VSS.n8817 VSS.n8816 0.04025
R12562 VSS.n8816 VSS.n8815 0.04025
R12563 VSS.n8815 VSS.n1628 0.04025
R12564 VSS.n8811 VSS.n1628 0.04025
R12565 VSS.n8811 VSS.n8810 0.04025
R12566 VSS.n8810 VSS.n8809 0.04025
R12567 VSS.n8809 VSS.n1630 0.04025
R12568 VSS.n8805 VSS.n1630 0.04025
R12569 VSS.n8805 VSS.n8804 0.04025
R12570 VSS.n8804 VSS.n8803 0.04025
R12571 VSS.n8803 VSS.n1632 0.04025
R12572 VSS.n8799 VSS.n1632 0.04025
R12573 VSS.n8799 VSS.n8798 0.04025
R12574 VSS.n8798 VSS.n8797 0.04025
R12575 VSS.n8797 VSS.n1634 0.04025
R12576 VSS.n8793 VSS.n1634 0.04025
R12577 VSS.n8793 VSS.n8792 0.04025
R12578 VSS.n8792 VSS.n8791 0.04025
R12579 VSS.n8791 VSS.n1636 0.04025
R12580 VSS.n8787 VSS.n1636 0.04025
R12581 VSS.n8787 VSS.n8786 0.04025
R12582 VSS.n8786 VSS.n8785 0.04025
R12583 VSS.n8785 VSS.n1638 0.04025
R12584 VSS.n8781 VSS.n1638 0.04025
R12585 VSS.n8781 VSS.n8780 0.04025
R12586 VSS.n8780 VSS.n8779 0.04025
R12587 VSS.n8779 VSS.n1640 0.04025
R12588 VSS.n8775 VSS.n1640 0.04025
R12589 VSS.n8775 VSS.n8774 0.04025
R12590 VSS.n8774 VSS.n8773 0.04025
R12591 VSS.n8773 VSS.n1642 0.04025
R12592 VSS.n8769 VSS.n1642 0.04025
R12593 VSS.n8769 VSS.n8768 0.04025
R12594 VSS.n8768 VSS.n8767 0.04025
R12595 VSS.n8767 VSS.n1644 0.04025
R12596 VSS.n8763 VSS.n1644 0.04025
R12597 VSS.n8763 VSS.n8762 0.04025
R12598 VSS.n8762 VSS.n8761 0.04025
R12599 VSS.n8761 VSS.n1646 0.04025
R12600 VSS.n8757 VSS.n1646 0.04025
R12601 VSS.n8757 VSS.n8756 0.04025
R12602 VSS.n8756 VSS.n8755 0.04025
R12603 VSS.n8755 VSS.n1648 0.04025
R12604 VSS.n8751 VSS.n1648 0.04025
R12605 VSS.n8751 VSS.n8750 0.04025
R12606 VSS.n8750 VSS.n8749 0.04025
R12607 VSS.n8749 VSS.n1650 0.04025
R12608 VSS.n8745 VSS.n1650 0.04025
R12609 VSS.n8745 VSS.n8744 0.04025
R12610 VSS.n8744 VSS.n8743 0.04025
R12611 VSS.n8743 VSS.n1652 0.04025
R12612 VSS.n8739 VSS.n1652 0.04025
R12613 VSS.n8739 VSS.n8738 0.04025
R12614 VSS.n8738 VSS.n8737 0.04025
R12615 VSS.n8737 VSS.n1654 0.04025
R12616 VSS.n8733 VSS.n1654 0.04025
R12617 VSS.n8733 VSS.n8732 0.04025
R12618 VSS.n8732 VSS.n8731 0.04025
R12619 VSS.n8731 VSS.n1656 0.04025
R12620 VSS.n8727 VSS.n1656 0.04025
R12621 VSS.n8727 VSS.n8726 0.04025
R12622 VSS.n8726 VSS.n8725 0.04025
R12623 VSS.n8725 VSS.n1658 0.04025
R12624 VSS.n8721 VSS.n1658 0.04025
R12625 VSS.n8721 VSS.n8720 0.04025
R12626 VSS.n8720 VSS.n8719 0.04025
R12627 VSS.n8719 VSS.n1660 0.04025
R12628 VSS.n8715 VSS.n1660 0.04025
R12629 VSS.n8715 VSS.n8714 0.04025
R12630 VSS.n8714 VSS.n8713 0.04025
R12631 VSS.n8713 VSS.n1662 0.04025
R12632 VSS.n8709 VSS.n1662 0.04025
R12633 VSS.n8709 VSS.n8708 0.04025
R12634 VSS.n8708 VSS.n8707 0.04025
R12635 VSS.n8707 VSS.n1664 0.04025
R12636 VSS.n8703 VSS.n1664 0.04025
R12637 VSS.n8703 VSS.n8702 0.04025
R12638 VSS.n8702 VSS.n8701 0.04025
R12639 VSS.n8701 VSS.n1666 0.04025
R12640 VSS.n8697 VSS.n1666 0.04025
R12641 VSS.n8697 VSS.n8696 0.04025
R12642 VSS.n8696 VSS.n8695 0.04025
R12643 VSS.n8695 VSS.n1668 0.04025
R12644 VSS.n8691 VSS.n1668 0.04025
R12645 VSS.n8691 VSS.n8690 0.04025
R12646 VSS.n8690 VSS.n8689 0.04025
R12647 VSS.n8689 VSS.n1670 0.04025
R12648 VSS.n8685 VSS.n1670 0.04025
R12649 VSS.n8685 VSS.n8684 0.04025
R12650 VSS.n8684 VSS.n8683 0.04025
R12651 VSS.n8683 VSS.n1672 0.04025
R12652 VSS.n8679 VSS.n1672 0.04025
R12653 VSS.n8679 VSS.n8678 0.04025
R12654 VSS.n8678 VSS.n8677 0.04025
R12655 VSS.n8677 VSS.n1674 0.04025
R12656 VSS.n8673 VSS.n1674 0.04025
R12657 VSS.n8673 VSS.n8672 0.04025
R12658 VSS.n8672 VSS.n8671 0.04025
R12659 VSS.n8671 VSS.n1676 0.04025
R12660 VSS.n8667 VSS.n1676 0.04025
R12661 VSS.n8667 VSS.n8666 0.04025
R12662 VSS.n8666 VSS.n8665 0.04025
R12663 VSS.n8665 VSS.n1678 0.04025
R12664 VSS.n8661 VSS.n1678 0.04025
R12665 VSS.n8661 VSS.n8660 0.04025
R12666 VSS.n8660 VSS.n8659 0.04025
R12667 VSS.n8659 VSS.n1680 0.04025
R12668 VSS.n8655 VSS.n1680 0.04025
R12669 VSS.n8655 VSS.n8654 0.04025
R12670 VSS.n8654 VSS.n8653 0.04025
R12671 VSS.n8653 VSS.n1682 0.04025
R12672 VSS.n8649 VSS.n1682 0.04025
R12673 VSS.n8649 VSS.n8648 0.04025
R12674 VSS.n8648 VSS.n8647 0.04025
R12675 VSS.n8647 VSS.n1684 0.04025
R12676 VSS.n8643 VSS.n1684 0.04025
R12677 VSS.n8643 VSS.n8642 0.04025
R12678 VSS.n8642 VSS.n8641 0.04025
R12679 VSS.n8641 VSS.n1686 0.04025
R12680 VSS.n8637 VSS.n1686 0.04025
R12681 VSS.n8637 VSS.n8636 0.04025
R12682 VSS.n8636 VSS.n8635 0.04025
R12683 VSS.n8635 VSS.n1688 0.04025
R12684 VSS.n8631 VSS.n1688 0.04025
R12685 VSS.n8631 VSS.n8630 0.04025
R12686 VSS.n8630 VSS.n8629 0.04025
R12687 VSS.n8629 VSS.n1690 0.04025
R12688 VSS.n8625 VSS.n1690 0.04025
R12689 VSS.n8625 VSS.n8624 0.04025
R12690 VSS.n8624 VSS.n8623 0.04025
R12691 VSS.n8623 VSS.n1692 0.04025
R12692 VSS.n8619 VSS.n1692 0.04025
R12693 VSS.n8619 VSS.n8618 0.04025
R12694 VSS.n8618 VSS.n8617 0.04025
R12695 VSS.n8617 VSS.n1694 0.04025
R12696 VSS.n8613 VSS.n1694 0.04025
R12697 VSS.n8613 VSS.n8612 0.04025
R12698 VSS.n8612 VSS.n8611 0.04025
R12699 VSS.n8611 VSS.n1696 0.04025
R12700 VSS.n8607 VSS.n1696 0.04025
R12701 VSS.n8607 VSS.n8606 0.04025
R12702 VSS.n8606 VSS.n8605 0.04025
R12703 VSS.n8605 VSS.n1698 0.04025
R12704 VSS.n8601 VSS.n1698 0.04025
R12705 VSS.n8601 VSS.n8600 0.04025
R12706 VSS.n8600 VSS.n8599 0.04025
R12707 VSS.n8599 VSS.n1700 0.04025
R12708 VSS.n8595 VSS.n1700 0.04025
R12709 VSS.n8595 VSS.n8594 0.04025
R12710 VSS.n8594 VSS.n8593 0.04025
R12711 VSS.n8593 VSS.n1702 0.04025
R12712 VSS.n8589 VSS.n1702 0.04025
R12713 VSS.n8589 VSS.n8588 0.04025
R12714 VSS.n8588 VSS.n8587 0.04025
R12715 VSS.n8587 VSS.n1704 0.04025
R12716 VSS.n8583 VSS.n1704 0.04025
R12717 VSS.n8583 VSS.n8582 0.04025
R12718 VSS.n8582 VSS.n8581 0.04025
R12719 VSS.n8581 VSS.n1706 0.04025
R12720 VSS.n8577 VSS.n1706 0.04025
R12721 VSS.n8577 VSS.n8576 0.04025
R12722 VSS.n8576 VSS.n8575 0.04025
R12723 VSS.n8575 VSS.n1708 0.04025
R12724 VSS.n8571 VSS.n1708 0.04025
R12725 VSS.n8571 VSS.n8570 0.04025
R12726 VSS.n8570 VSS.n8569 0.04025
R12727 VSS.n8569 VSS.n1710 0.04025
R12728 VSS.n8565 VSS.n1710 0.04025
R12729 VSS.n8565 VSS.n8564 0.04025
R12730 VSS.n8564 VSS.n8563 0.04025
R12731 VSS.n8563 VSS.n1712 0.04025
R12732 VSS.n8559 VSS.n1712 0.04025
R12733 VSS.n8559 VSS.n8558 0.04025
R12734 VSS.n8558 VSS.n8557 0.04025
R12735 VSS.n8557 VSS.n1714 0.04025
R12736 VSS.n8553 VSS.n1714 0.04025
R12737 VSS.n8553 VSS.n8552 0.04025
R12738 VSS.n8552 VSS.n8551 0.04025
R12739 VSS.n8551 VSS.n1716 0.04025
R12740 VSS.n8547 VSS.n1716 0.04025
R12741 VSS.n8547 VSS.n8546 0.04025
R12742 VSS.n8546 VSS.n8545 0.04025
R12743 VSS.n8545 VSS.n1718 0.04025
R12744 VSS.n8541 VSS.n1718 0.04025
R12745 VSS.n8541 VSS.n8540 0.04025
R12746 VSS.n8540 VSS.n8539 0.04025
R12747 VSS.n8539 VSS.n1720 0.04025
R12748 VSS.n8535 VSS.n1720 0.04025
R12749 VSS.n8535 VSS.n8534 0.04025
R12750 VSS.n8534 VSS.n8533 0.04025
R12751 VSS.n8533 VSS.n1722 0.04025
R12752 VSS.n8529 VSS.n1722 0.04025
R12753 VSS.n8529 VSS.n8528 0.04025
R12754 VSS.n8528 VSS.n8527 0.04025
R12755 VSS.n8527 VSS.n1724 0.04025
R12756 VSS.n8523 VSS.n1724 0.04025
R12757 VSS.n8523 VSS.n8522 0.04025
R12758 VSS.n8522 VSS.n8521 0.04025
R12759 VSS.n8521 VSS.n1726 0.04025
R12760 VSS.n8517 VSS.n1726 0.04025
R12761 VSS.n8517 VSS.n8516 0.04025
R12762 VSS.n8516 VSS.n8515 0.04025
R12763 VSS.n8515 VSS.n1728 0.04025
R12764 VSS.n8511 VSS.n1728 0.04025
R12765 VSS.n8511 VSS.n8510 0.04025
R12766 VSS.n8510 VSS.n8509 0.04025
R12767 VSS.n8509 VSS.n1730 0.04025
R12768 VSS.n8505 VSS.n1730 0.04025
R12769 VSS.n8505 VSS.n8504 0.04025
R12770 VSS.n8504 VSS.n8503 0.04025
R12771 VSS.n8503 VSS.n1732 0.04025
R12772 VSS.n8499 VSS.n1732 0.04025
R12773 VSS.n8499 VSS.n8498 0.04025
R12774 VSS.n8498 VSS.n8497 0.04025
R12775 VSS.n8497 VSS.n1734 0.04025
R12776 VSS.n8493 VSS.n1734 0.04025
R12777 VSS.n8493 VSS.n8492 0.04025
R12778 VSS.n8492 VSS.n8491 0.04025
R12779 VSS.n8491 VSS.n1736 0.04025
R12780 VSS.n8487 VSS.n1736 0.04025
R12781 VSS.n8487 VSS.n8486 0.04025
R12782 VSS.n8486 VSS.n8485 0.04025
R12783 VSS.n8485 VSS.n1738 0.04025
R12784 VSS.n8481 VSS.n1738 0.04025
R12785 VSS.n8481 VSS.n8480 0.04025
R12786 VSS.n8480 VSS.n8479 0.04025
R12787 VSS.n8479 VSS.n1740 0.04025
R12788 VSS.n8475 VSS.n1740 0.04025
R12789 VSS.n8475 VSS.n8474 0.04025
R12790 VSS.n8474 VSS.n8473 0.04025
R12791 VSS.n8473 VSS.n1742 0.04025
R12792 VSS.n8469 VSS.n1742 0.04025
R12793 VSS.n8469 VSS.n8468 0.04025
R12794 VSS.n8468 VSS.n8467 0.04025
R12795 VSS.n8467 VSS.n1744 0.04025
R12796 VSS.n8463 VSS.n1744 0.04025
R12797 VSS.n8463 VSS.n8462 0.04025
R12798 VSS.n8462 VSS.n8461 0.04025
R12799 VSS.n8461 VSS.n1746 0.04025
R12800 VSS.n8457 VSS.n1746 0.04025
R12801 VSS.n8457 VSS.n8456 0.04025
R12802 VSS.n8456 VSS.n8455 0.04025
R12803 VSS.n8455 VSS.n1748 0.04025
R12804 VSS.n8451 VSS.n1748 0.04025
R12805 VSS.n8451 VSS.n8450 0.04025
R12806 VSS.n8450 VSS.n8449 0.04025
R12807 VSS.n8449 VSS.n1750 0.04025
R12808 VSS.n8445 VSS.n1750 0.04025
R12809 VSS.n8445 VSS.n8444 0.04025
R12810 VSS.n8444 VSS.n8443 0.04025
R12811 VSS.n8443 VSS.n1752 0.04025
R12812 VSS.n8439 VSS.n1752 0.04025
R12813 VSS.n8439 VSS.n8438 0.04025
R12814 VSS.n8438 VSS.n8437 0.04025
R12815 VSS.n8437 VSS.n1754 0.04025
R12816 VSS.n8433 VSS.n1754 0.04025
R12817 VSS.n8433 VSS.n8432 0.04025
R12818 VSS.n8432 VSS.n8431 0.04025
R12819 VSS.n8431 VSS.n1756 0.04025
R12820 VSS.n8427 VSS.n1756 0.04025
R12821 VSS.n8427 VSS.n8426 0.04025
R12822 VSS.n8426 VSS.n8425 0.04025
R12823 VSS.n8425 VSS.n1758 0.04025
R12824 VSS.n8421 VSS.n1758 0.04025
R12825 VSS.n8421 VSS.n8420 0.04025
R12826 VSS.n8420 VSS.n8419 0.04025
R12827 VSS.n8419 VSS.n1760 0.04025
R12828 VSS.n8415 VSS.n1760 0.04025
R12829 VSS.n8415 VSS.n8414 0.04025
R12830 VSS.n8414 VSS.n8413 0.04025
R12831 VSS.n8413 VSS.n1762 0.04025
R12832 VSS.n8409 VSS.n1762 0.04025
R12833 VSS.n8409 VSS.n8408 0.04025
R12834 VSS.n8408 VSS.n8407 0.04025
R12835 VSS.n8407 VSS.n1764 0.04025
R12836 VSS.n8403 VSS.n1764 0.04025
R12837 VSS.n8403 VSS.n8402 0.04025
R12838 VSS.n8402 VSS.n8401 0.04025
R12839 VSS.n8401 VSS.n1766 0.04025
R12840 VSS.n8397 VSS.n1766 0.04025
R12841 VSS.n8397 VSS.n8396 0.04025
R12842 VSS.n8396 VSS.n8395 0.04025
R12843 VSS.n8395 VSS.n1768 0.04025
R12844 VSS.n8391 VSS.n1768 0.04025
R12845 VSS.n8391 VSS.n8390 0.04025
R12846 VSS.n8390 VSS.n8389 0.04025
R12847 VSS.n8389 VSS.n1770 0.04025
R12848 VSS.n8385 VSS.n1770 0.04025
R12849 VSS.n8385 VSS.n8384 0.04025
R12850 VSS.n8384 VSS.n8383 0.04025
R12851 VSS.n8383 VSS.n1772 0.04025
R12852 VSS.n8379 VSS.n1772 0.04025
R12853 VSS.n8379 VSS.n8378 0.04025
R12854 VSS.n8378 VSS.n8377 0.04025
R12855 VSS.n8377 VSS.n1774 0.04025
R12856 VSS.n8373 VSS.n1774 0.04025
R12857 VSS.n8373 VSS.n8372 0.04025
R12858 VSS.n8372 VSS.n8371 0.04025
R12859 VSS.n8371 VSS.n1776 0.04025
R12860 VSS.n8367 VSS.n1776 0.04025
R12861 VSS.n8367 VSS.n8366 0.04025
R12862 VSS.n8366 VSS.n8365 0.04025
R12863 VSS.n8365 VSS.n1778 0.04025
R12864 VSS.n8361 VSS.n1778 0.04025
R12865 VSS.n8361 VSS.n8360 0.04025
R12866 VSS.n8360 VSS.n8359 0.04025
R12867 VSS.n8359 VSS.n1780 0.04025
R12868 VSS.n8355 VSS.n1780 0.04025
R12869 VSS.n8355 VSS.n8354 0.04025
R12870 VSS.n8354 VSS.n8353 0.04025
R12871 VSS.n8353 VSS.n1782 0.04025
R12872 VSS.n8349 VSS.n1782 0.04025
R12873 VSS.n8349 VSS.n8348 0.04025
R12874 VSS.n8348 VSS.n8347 0.04025
R12875 VSS.n8347 VSS.n1784 0.04025
R12876 VSS.n8343 VSS.n1784 0.04025
R12877 VSS.n8343 VSS.n8342 0.04025
R12878 VSS.n8342 VSS.n8341 0.04025
R12879 VSS.n8341 VSS.n1786 0.04025
R12880 VSS.n8337 VSS.n1786 0.04025
R12881 VSS.n8337 VSS.n8336 0.04025
R12882 VSS.n8336 VSS.n8335 0.04025
R12883 VSS.n8335 VSS.n1788 0.04025
R12884 VSS.n8331 VSS.n1788 0.04025
R12885 VSS.n8331 VSS.n8330 0.04025
R12886 VSS.n8330 VSS.n8329 0.04025
R12887 VSS.n8329 VSS.n1790 0.04025
R12888 VSS.n8325 VSS.n1790 0.04025
R12889 VSS.n8325 VSS.n8324 0.04025
R12890 VSS.n8324 VSS.n8323 0.04025
R12891 VSS.n8323 VSS.n1792 0.04025
R12892 VSS.n8319 VSS.n1792 0.04025
R12893 VSS.n8319 VSS.n8318 0.04025
R12894 VSS.n8318 VSS.n8317 0.04025
R12895 VSS.n8317 VSS.n1794 0.04025
R12896 VSS.n8313 VSS.n1794 0.04025
R12897 VSS.n8313 VSS.n8312 0.04025
R12898 VSS.n8312 VSS.n8311 0.04025
R12899 VSS.n8311 VSS.n1796 0.04025
R12900 VSS.n8307 VSS.n1796 0.04025
R12901 VSS.n8307 VSS.n8306 0.04025
R12902 VSS.n8306 VSS.n8305 0.04025
R12903 VSS.n8305 VSS.n1798 0.04025
R12904 VSS.n8301 VSS.n1798 0.04025
R12905 VSS.n8301 VSS.n8300 0.04025
R12906 VSS.n8300 VSS.n8299 0.04025
R12907 VSS.n8299 VSS.n1800 0.04025
R12908 VSS.n8295 VSS.n1800 0.04025
R12909 VSS.n8295 VSS.n8294 0.04025
R12910 VSS.n8294 VSS.n8293 0.04025
R12911 VSS.n8293 VSS.n1802 0.04025
R12912 VSS.n8289 VSS.n1802 0.04025
R12913 VSS.n8289 VSS.n8288 0.04025
R12914 VSS.n8288 VSS.n8287 0.04025
R12915 VSS.n8287 VSS.n1804 0.04025
R12916 VSS.n8283 VSS.n1804 0.04025
R12917 VSS.n8283 VSS.n8282 0.04025
R12918 VSS.n8282 VSS.n8281 0.04025
R12919 VSS.n8281 VSS.n1806 0.04025
R12920 VSS.n8277 VSS.n1806 0.04025
R12921 VSS.n8277 VSS.n8276 0.04025
R12922 VSS.n8276 VSS.n8275 0.04025
R12923 VSS.n8275 VSS.n1808 0.04025
R12924 VSS.n8271 VSS.n1808 0.04025
R12925 VSS.n8271 VSS.n8270 0.04025
R12926 VSS.n8270 VSS.n8269 0.04025
R12927 VSS.n8269 VSS.n1810 0.04025
R12928 VSS.n8265 VSS.n1810 0.04025
R12929 VSS.n8265 VSS.n8264 0.04025
R12930 VSS.n8264 VSS.n8263 0.04025
R12931 VSS.n8263 VSS.n1812 0.04025
R12932 VSS.n8259 VSS.n1812 0.04025
R12933 VSS.n8259 VSS.n8258 0.04025
R12934 VSS.n8258 VSS.n8257 0.04025
R12935 VSS.n8257 VSS.n1814 0.04025
R12936 VSS.n8253 VSS.n1814 0.04025
R12937 VSS.n8253 VSS.n8252 0.04025
R12938 VSS.n8252 VSS.n8251 0.04025
R12939 VSS.n8251 VSS.n1816 0.04025
R12940 VSS.n8247 VSS.n1816 0.04025
R12941 VSS.n8247 VSS.n8246 0.04025
R12942 VSS.n8246 VSS.n8245 0.04025
R12943 VSS.n8245 VSS.n1818 0.04025
R12944 VSS.n8241 VSS.n1818 0.04025
R12945 VSS.n8241 VSS.n8240 0.04025
R12946 VSS.n8240 VSS.n8239 0.04025
R12947 VSS.n8239 VSS.n1820 0.04025
R12948 VSS.n8235 VSS.n1820 0.04025
R12949 VSS.n8235 VSS.n8234 0.04025
R12950 VSS.n8234 VSS.n8233 0.04025
R12951 VSS.n4144 VSS.n3184 0.04025
R12952 VSS.n4145 VSS.n4144 0.04025
R12953 VSS.n4146 VSS.n4145 0.04025
R12954 VSS.n4146 VSS.n3182 0.04025
R12955 VSS.n4150 VSS.n3182 0.04025
R12956 VSS.n4151 VSS.n4150 0.04025
R12957 VSS.n4152 VSS.n4151 0.04025
R12958 VSS.n4152 VSS.n3180 0.04025
R12959 VSS.n4156 VSS.n3180 0.04025
R12960 VSS.n4157 VSS.n4156 0.04025
R12961 VSS.n4158 VSS.n4157 0.04025
R12962 VSS.n4158 VSS.n3178 0.04025
R12963 VSS.n4162 VSS.n3178 0.04025
R12964 VSS.n4163 VSS.n4162 0.04025
R12965 VSS.n4164 VSS.n4163 0.04025
R12966 VSS.n4164 VSS.n3176 0.04025
R12967 VSS.n4168 VSS.n3176 0.04025
R12968 VSS.n4169 VSS.n4168 0.04025
R12969 VSS.n4170 VSS.n4169 0.04025
R12970 VSS.n4170 VSS.n3174 0.04025
R12971 VSS.n4174 VSS.n3174 0.04025
R12972 VSS.n4175 VSS.n4174 0.04025
R12973 VSS.n4176 VSS.n4175 0.04025
R12974 VSS.n4176 VSS.n3172 0.04025
R12975 VSS.n4180 VSS.n3172 0.04025
R12976 VSS.n4181 VSS.n4180 0.04025
R12977 VSS.n4182 VSS.n4181 0.04025
R12978 VSS.n4182 VSS.n3170 0.04025
R12979 VSS.n4186 VSS.n3170 0.04025
R12980 VSS.n4187 VSS.n4186 0.04025
R12981 VSS.n4188 VSS.n4187 0.04025
R12982 VSS.n4188 VSS.n3168 0.04025
R12983 VSS.n4192 VSS.n3168 0.04025
R12984 VSS.n4193 VSS.n4192 0.04025
R12985 VSS.n4194 VSS.n4193 0.04025
R12986 VSS.n4194 VSS.n3166 0.04025
R12987 VSS.n4198 VSS.n3166 0.04025
R12988 VSS.n4199 VSS.n4198 0.04025
R12989 VSS.n4200 VSS.n4199 0.04025
R12990 VSS.n4200 VSS.n3164 0.04025
R12991 VSS.n4204 VSS.n3164 0.04025
R12992 VSS.n4205 VSS.n4204 0.04025
R12993 VSS.n4206 VSS.n4205 0.04025
R12994 VSS.n4206 VSS.n3162 0.04025
R12995 VSS.n4210 VSS.n3162 0.04025
R12996 VSS.n4211 VSS.n4210 0.04025
R12997 VSS.n4212 VSS.n4211 0.04025
R12998 VSS.n4212 VSS.n3160 0.04025
R12999 VSS.n4216 VSS.n3160 0.04025
R13000 VSS.n4217 VSS.n4216 0.04025
R13001 VSS.n4218 VSS.n4217 0.04025
R13002 VSS.n4218 VSS.n3158 0.04025
R13003 VSS.n4222 VSS.n3158 0.04025
R13004 VSS.n4223 VSS.n4222 0.04025
R13005 VSS.n4224 VSS.n4223 0.04025
R13006 VSS.n4224 VSS.n3156 0.04025
R13007 VSS.n4228 VSS.n3156 0.04025
R13008 VSS.n4229 VSS.n4228 0.04025
R13009 VSS.n4230 VSS.n4229 0.04025
R13010 VSS.n4230 VSS.n3154 0.04025
R13011 VSS.n4234 VSS.n3154 0.04025
R13012 VSS.n4235 VSS.n4234 0.04025
R13013 VSS.n4236 VSS.n4235 0.04025
R13014 VSS.n4236 VSS.n3152 0.04025
R13015 VSS.n4240 VSS.n3152 0.04025
R13016 VSS.n4241 VSS.n4240 0.04025
R13017 VSS.n4242 VSS.n4241 0.04025
R13018 VSS.n4242 VSS.n3150 0.04025
R13019 VSS.n4246 VSS.n3150 0.04025
R13020 VSS.n4247 VSS.n4246 0.04025
R13021 VSS.n4248 VSS.n4247 0.04025
R13022 VSS.n4248 VSS.n3148 0.04025
R13023 VSS.n4252 VSS.n3148 0.04025
R13024 VSS.n4253 VSS.n4252 0.04025
R13025 VSS.n4254 VSS.n4253 0.04025
R13026 VSS.n4254 VSS.n3146 0.04025
R13027 VSS.n4258 VSS.n3146 0.04025
R13028 VSS.n4259 VSS.n4258 0.04025
R13029 VSS.n4260 VSS.n4259 0.04025
R13030 VSS.n4260 VSS.n3144 0.04025
R13031 VSS.n4264 VSS.n3144 0.04025
R13032 VSS.n4265 VSS.n4264 0.04025
R13033 VSS.n4266 VSS.n4265 0.04025
R13034 VSS.n4266 VSS.n3142 0.04025
R13035 VSS.n4270 VSS.n3142 0.04025
R13036 VSS.n4271 VSS.n4270 0.04025
R13037 VSS.n4272 VSS.n4271 0.04025
R13038 VSS.n4272 VSS.n3140 0.04025
R13039 VSS.n4276 VSS.n3140 0.04025
R13040 VSS.n4277 VSS.n4276 0.04025
R13041 VSS.n4278 VSS.n4277 0.04025
R13042 VSS.n4278 VSS.n3138 0.04025
R13043 VSS.n4282 VSS.n3138 0.04025
R13044 VSS.n4283 VSS.n4282 0.04025
R13045 VSS.n4284 VSS.n4283 0.04025
R13046 VSS.n4284 VSS.n3136 0.04025
R13047 VSS.n4288 VSS.n3136 0.04025
R13048 VSS.n4289 VSS.n4288 0.04025
R13049 VSS.n4290 VSS.n4289 0.04025
R13050 VSS.n4290 VSS.n3134 0.04025
R13051 VSS.n4294 VSS.n3134 0.04025
R13052 VSS.n4295 VSS.n4294 0.04025
R13053 VSS.n4296 VSS.n4295 0.04025
R13054 VSS.n4296 VSS.n3132 0.04025
R13055 VSS.n4300 VSS.n3132 0.04025
R13056 VSS.n4301 VSS.n4300 0.04025
R13057 VSS.n4302 VSS.n4301 0.04025
R13058 VSS.n4302 VSS.n3130 0.04025
R13059 VSS.n4306 VSS.n3130 0.04025
R13060 VSS.n4307 VSS.n4306 0.04025
R13061 VSS.n4308 VSS.n4307 0.04025
R13062 VSS.n4308 VSS.n3128 0.04025
R13063 VSS.n4312 VSS.n3128 0.04025
R13064 VSS.n4313 VSS.n4312 0.04025
R13065 VSS.n4314 VSS.n4313 0.04025
R13066 VSS.n4314 VSS.n3126 0.04025
R13067 VSS.n4318 VSS.n3126 0.04025
R13068 VSS.n4319 VSS.n4318 0.04025
R13069 VSS.n4320 VSS.n4319 0.04025
R13070 VSS.n4320 VSS.n3124 0.04025
R13071 VSS.n4324 VSS.n3124 0.04025
R13072 VSS.n4325 VSS.n4324 0.04025
R13073 VSS.n4326 VSS.n4325 0.04025
R13074 VSS.n4326 VSS.n3122 0.04025
R13075 VSS.n4330 VSS.n3122 0.04025
R13076 VSS.n4331 VSS.n4330 0.04025
R13077 VSS.n4332 VSS.n4331 0.04025
R13078 VSS.n4332 VSS.n3120 0.04025
R13079 VSS.n4336 VSS.n3120 0.04025
R13080 VSS.n4337 VSS.n4336 0.04025
R13081 VSS.n4338 VSS.n4337 0.04025
R13082 VSS.n4338 VSS.n3118 0.04025
R13083 VSS.n4342 VSS.n3118 0.04025
R13084 VSS.n4343 VSS.n4342 0.04025
R13085 VSS.n4344 VSS.n4343 0.04025
R13086 VSS.n4344 VSS.n3116 0.04025
R13087 VSS.n4348 VSS.n3116 0.04025
R13088 VSS.n4349 VSS.n4348 0.04025
R13089 VSS.n4350 VSS.n4349 0.04025
R13090 VSS.n4350 VSS.n3114 0.04025
R13091 VSS.n4354 VSS.n3114 0.04025
R13092 VSS.n4355 VSS.n4354 0.04025
R13093 VSS.n4356 VSS.n4355 0.04025
R13094 VSS.n4356 VSS.n3112 0.04025
R13095 VSS.n4360 VSS.n3112 0.04025
R13096 VSS.n4361 VSS.n4360 0.04025
R13097 VSS.n4362 VSS.n4361 0.04025
R13098 VSS.n4362 VSS.n3110 0.04025
R13099 VSS.n4366 VSS.n3110 0.04025
R13100 VSS.n4367 VSS.n4366 0.04025
R13101 VSS.n4368 VSS.n4367 0.04025
R13102 VSS.n4368 VSS.n3108 0.04025
R13103 VSS.n4372 VSS.n3108 0.04025
R13104 VSS.n4373 VSS.n4372 0.04025
R13105 VSS.n4374 VSS.n4373 0.04025
R13106 VSS.n4374 VSS.n3106 0.04025
R13107 VSS.n4378 VSS.n3106 0.04025
R13108 VSS.n4379 VSS.n4378 0.04025
R13109 VSS.n4380 VSS.n4379 0.04025
R13110 VSS.n4380 VSS.n3104 0.04025
R13111 VSS.n4384 VSS.n3104 0.04025
R13112 VSS.n4385 VSS.n4384 0.04025
R13113 VSS.n4386 VSS.n4385 0.04025
R13114 VSS.n4386 VSS.n3102 0.04025
R13115 VSS.n4390 VSS.n3102 0.04025
R13116 VSS.n4391 VSS.n4390 0.04025
R13117 VSS.n4392 VSS.n4391 0.04025
R13118 VSS.n4392 VSS.n3100 0.04025
R13119 VSS.n4396 VSS.n3100 0.04025
R13120 VSS.n4397 VSS.n4396 0.04025
R13121 VSS.n4398 VSS.n4397 0.04025
R13122 VSS.n4398 VSS.n3098 0.04025
R13123 VSS.n4402 VSS.n3098 0.04025
R13124 VSS.n4403 VSS.n4402 0.04025
R13125 VSS.n4404 VSS.n4403 0.04025
R13126 VSS.n4404 VSS.n3096 0.04025
R13127 VSS.n4408 VSS.n3096 0.04025
R13128 VSS.n4409 VSS.n4408 0.04025
R13129 VSS.n4410 VSS.n4409 0.04025
R13130 VSS.n4410 VSS.n3094 0.04025
R13131 VSS.n4414 VSS.n3094 0.04025
R13132 VSS.n4415 VSS.n4414 0.04025
R13133 VSS.n4416 VSS.n4415 0.04025
R13134 VSS.n4416 VSS.n3092 0.04025
R13135 VSS.n4420 VSS.n3092 0.04025
R13136 VSS.n4421 VSS.n4420 0.04025
R13137 VSS.n4422 VSS.n4421 0.04025
R13138 VSS.n4422 VSS.n3090 0.04025
R13139 VSS.n4426 VSS.n3090 0.04025
R13140 VSS.n4427 VSS.n4426 0.04025
R13141 VSS.n4428 VSS.n4427 0.04025
R13142 VSS.n4428 VSS.n3088 0.04025
R13143 VSS.n4432 VSS.n3088 0.04025
R13144 VSS.n4433 VSS.n4432 0.04025
R13145 VSS.n4434 VSS.n4433 0.04025
R13146 VSS.n4434 VSS.n3086 0.04025
R13147 VSS.n4438 VSS.n3086 0.04025
R13148 VSS.n4439 VSS.n4438 0.04025
R13149 VSS.n4440 VSS.n4439 0.04025
R13150 VSS.n4440 VSS.n3084 0.04025
R13151 VSS.n4444 VSS.n3084 0.04025
R13152 VSS.n4445 VSS.n4444 0.04025
R13153 VSS.n4446 VSS.n4445 0.04025
R13154 VSS.n4446 VSS.n3082 0.04025
R13155 VSS.n4450 VSS.n3082 0.04025
R13156 VSS.n4451 VSS.n4450 0.04025
R13157 VSS.n4452 VSS.n4451 0.04025
R13158 VSS.n4452 VSS.n3080 0.04025
R13159 VSS.n4456 VSS.n3080 0.04025
R13160 VSS.n4457 VSS.n4456 0.04025
R13161 VSS.n4458 VSS.n4457 0.04025
R13162 VSS.n4458 VSS.n3078 0.04025
R13163 VSS.n4462 VSS.n3078 0.04025
R13164 VSS.n4463 VSS.n4462 0.04025
R13165 VSS.n4464 VSS.n4463 0.04025
R13166 VSS.n4464 VSS.n3076 0.04025
R13167 VSS.n4468 VSS.n3076 0.04025
R13168 VSS.n4469 VSS.n4468 0.04025
R13169 VSS.n4470 VSS.n4469 0.04025
R13170 VSS.n4470 VSS.n3074 0.04025
R13171 VSS.n4474 VSS.n3074 0.04025
R13172 VSS.n4475 VSS.n4474 0.04025
R13173 VSS.n4476 VSS.n4475 0.04025
R13174 VSS.n4476 VSS.n3072 0.04025
R13175 VSS.n4480 VSS.n3072 0.04025
R13176 VSS.n4481 VSS.n4480 0.04025
R13177 VSS.n4482 VSS.n4481 0.04025
R13178 VSS.n4482 VSS.n3070 0.04025
R13179 VSS.n4486 VSS.n3070 0.04025
R13180 VSS.n4487 VSS.n4486 0.04025
R13181 VSS.n4488 VSS.n4487 0.04025
R13182 VSS.n4488 VSS.n3068 0.04025
R13183 VSS.n4492 VSS.n3068 0.04025
R13184 VSS.n4493 VSS.n4492 0.04025
R13185 VSS.n4494 VSS.n4493 0.04025
R13186 VSS.n4494 VSS.n3066 0.04025
R13187 VSS.n4498 VSS.n3066 0.04025
R13188 VSS.n4499 VSS.n4498 0.04025
R13189 VSS.n4500 VSS.n4499 0.04025
R13190 VSS.n4500 VSS.n3064 0.04025
R13191 VSS.n4504 VSS.n3064 0.04025
R13192 VSS.n4505 VSS.n4504 0.04025
R13193 VSS.n4506 VSS.n4505 0.04025
R13194 VSS.n4506 VSS.n3062 0.04025
R13195 VSS.n4510 VSS.n3062 0.04025
R13196 VSS.n4511 VSS.n4510 0.04025
R13197 VSS.n4512 VSS.n4511 0.04025
R13198 VSS.n4512 VSS.n3060 0.04025
R13199 VSS.n4516 VSS.n3060 0.04025
R13200 VSS.n4517 VSS.n4516 0.04025
R13201 VSS.n4518 VSS.n4517 0.04025
R13202 VSS.n4518 VSS.n3058 0.04025
R13203 VSS.n4522 VSS.n3058 0.04025
R13204 VSS.n4523 VSS.n4522 0.04025
R13205 VSS.n4524 VSS.n4523 0.04025
R13206 VSS.n4524 VSS.n3056 0.04025
R13207 VSS.n4528 VSS.n3056 0.04025
R13208 VSS.n4529 VSS.n4528 0.04025
R13209 VSS.n4530 VSS.n4529 0.04025
R13210 VSS.n4530 VSS.n3054 0.04025
R13211 VSS.n4534 VSS.n3054 0.04025
R13212 VSS.n4535 VSS.n4534 0.04025
R13213 VSS.n4536 VSS.n4535 0.04025
R13214 VSS.n4536 VSS.n3052 0.04025
R13215 VSS.n4540 VSS.n3052 0.04025
R13216 VSS.n4541 VSS.n4540 0.04025
R13217 VSS.n4542 VSS.n4541 0.04025
R13218 VSS.n4542 VSS.n3050 0.04025
R13219 VSS.n4546 VSS.n3050 0.04025
R13220 VSS.n4547 VSS.n4546 0.04025
R13221 VSS.n4548 VSS.n4547 0.04025
R13222 VSS.n4548 VSS.n3048 0.04025
R13223 VSS.n4552 VSS.n3048 0.04025
R13224 VSS.n4553 VSS.n4552 0.04025
R13225 VSS.n4554 VSS.n4553 0.04025
R13226 VSS.n4554 VSS.n3046 0.04025
R13227 VSS.n4558 VSS.n3046 0.04025
R13228 VSS.n4559 VSS.n4558 0.04025
R13229 VSS.n4560 VSS.n4559 0.04025
R13230 VSS.n4560 VSS.n3044 0.04025
R13231 VSS.n4564 VSS.n3044 0.04025
R13232 VSS.n4565 VSS.n4564 0.04025
R13233 VSS.n4566 VSS.n4565 0.04025
R13234 VSS.n4566 VSS.n3042 0.04025
R13235 VSS.n4570 VSS.n3042 0.04025
R13236 VSS.n4571 VSS.n4570 0.04025
R13237 VSS.n4572 VSS.n4571 0.04025
R13238 VSS.n4572 VSS.n3040 0.04025
R13239 VSS.n4576 VSS.n3040 0.04025
R13240 VSS.n4577 VSS.n4576 0.04025
R13241 VSS.n4578 VSS.n4577 0.04025
R13242 VSS.n4578 VSS.n3038 0.04025
R13243 VSS.n4582 VSS.n3038 0.04025
R13244 VSS.n4583 VSS.n4582 0.04025
R13245 VSS.n4584 VSS.n4583 0.04025
R13246 VSS.n4584 VSS.n3036 0.04025
R13247 VSS.n4588 VSS.n3036 0.04025
R13248 VSS.n4589 VSS.n4588 0.04025
R13249 VSS.n4590 VSS.n4589 0.04025
R13250 VSS.n4590 VSS.n3034 0.04025
R13251 VSS.n4594 VSS.n3034 0.04025
R13252 VSS.n4595 VSS.n4594 0.04025
R13253 VSS.n4596 VSS.n4595 0.04025
R13254 VSS.n4596 VSS.n3032 0.04025
R13255 VSS.n4600 VSS.n3032 0.04025
R13256 VSS.n4601 VSS.n4600 0.04025
R13257 VSS.n4602 VSS.n4601 0.04025
R13258 VSS.n4602 VSS.n3030 0.04025
R13259 VSS.n4606 VSS.n3030 0.04025
R13260 VSS.n4607 VSS.n4606 0.04025
R13261 VSS.n4608 VSS.n4607 0.04025
R13262 VSS.n4608 VSS.n3028 0.04025
R13263 VSS.n4612 VSS.n3028 0.04025
R13264 VSS.n4613 VSS.n4612 0.04025
R13265 VSS.n4614 VSS.n4613 0.04025
R13266 VSS.n4614 VSS.n3026 0.04025
R13267 VSS.n4618 VSS.n3026 0.04025
R13268 VSS.n4619 VSS.n4618 0.04025
R13269 VSS.n4620 VSS.n4619 0.04025
R13270 VSS.n4620 VSS.n3024 0.04025
R13271 VSS.n4624 VSS.n3024 0.04025
R13272 VSS.n4625 VSS.n4624 0.04025
R13273 VSS.n4626 VSS.n4625 0.04025
R13274 VSS.n4626 VSS.n3022 0.04025
R13275 VSS.n4630 VSS.n3022 0.04025
R13276 VSS.n4631 VSS.n4630 0.04025
R13277 VSS.n4632 VSS.n4631 0.04025
R13278 VSS.n4632 VSS.n3020 0.04025
R13279 VSS.n4636 VSS.n3020 0.04025
R13280 VSS.n4637 VSS.n4636 0.04025
R13281 VSS.n4638 VSS.n4637 0.04025
R13282 VSS.n4638 VSS.n3018 0.04025
R13283 VSS.n4642 VSS.n3018 0.04025
R13284 VSS.n4643 VSS.n4642 0.04025
R13285 VSS.n4644 VSS.n4643 0.04025
R13286 VSS.n4644 VSS.n3016 0.04025
R13287 VSS.n4648 VSS.n3016 0.04025
R13288 VSS.n4649 VSS.n4648 0.04025
R13289 VSS.n4650 VSS.n4649 0.04025
R13290 VSS.n4650 VSS.n3014 0.04025
R13291 VSS.n4654 VSS.n3014 0.04025
R13292 VSS.n4655 VSS.n4654 0.04025
R13293 VSS.n4656 VSS.n4655 0.04025
R13294 VSS.n4656 VSS.n3012 0.04025
R13295 VSS.n4660 VSS.n3012 0.04025
R13296 VSS.n4661 VSS.n4660 0.04025
R13297 VSS.n4662 VSS.n4661 0.04025
R13298 VSS.n4662 VSS.n3010 0.04025
R13299 VSS.n4666 VSS.n3010 0.04025
R13300 VSS.n4667 VSS.n4666 0.04025
R13301 VSS.n4668 VSS.n4667 0.04025
R13302 VSS.n4668 VSS.n3008 0.04025
R13303 VSS.n4672 VSS.n3008 0.04025
R13304 VSS.n4673 VSS.n4672 0.04025
R13305 VSS.n4674 VSS.n4673 0.04025
R13306 VSS.n4674 VSS.n3006 0.04025
R13307 VSS.n4678 VSS.n3006 0.04025
R13308 VSS.n4679 VSS.n4678 0.04025
R13309 VSS.n4680 VSS.n4679 0.04025
R13310 VSS.n4680 VSS.n3004 0.04025
R13311 VSS.n4684 VSS.n3004 0.04025
R13312 VSS.n4685 VSS.n4684 0.04025
R13313 VSS.n4686 VSS.n4685 0.04025
R13314 VSS.n4686 VSS.n3002 0.04025
R13315 VSS.n4690 VSS.n3002 0.04025
R13316 VSS.n4691 VSS.n4690 0.04025
R13317 VSS.n4692 VSS.n4691 0.04025
R13318 VSS.n4692 VSS.n3000 0.04025
R13319 VSS.n4696 VSS.n3000 0.04025
R13320 VSS.n4697 VSS.n4696 0.04025
R13321 VSS.n4698 VSS.n4697 0.04025
R13322 VSS.n4698 VSS.n2998 0.04025
R13323 VSS.n4702 VSS.n2998 0.04025
R13324 VSS.n4703 VSS.n4702 0.04025
R13325 VSS.n4704 VSS.n4703 0.04025
R13326 VSS.n4704 VSS.n2996 0.04025
R13327 VSS.n4708 VSS.n2996 0.04025
R13328 VSS.n4709 VSS.n4708 0.04025
R13329 VSS.n4710 VSS.n4709 0.04025
R13330 VSS.n4710 VSS.n2994 0.04025
R13331 VSS.n4714 VSS.n2994 0.04025
R13332 VSS.n4715 VSS.n4714 0.04025
R13333 VSS.n4716 VSS.n4715 0.04025
R13334 VSS.n4716 VSS.n2992 0.04025
R13335 VSS.n4720 VSS.n2992 0.04025
R13336 VSS.n4721 VSS.n4720 0.04025
R13337 VSS.n4722 VSS.n4721 0.04025
R13338 VSS.n4722 VSS.n2990 0.04025
R13339 VSS.n4726 VSS.n2990 0.04025
R13340 VSS.n4727 VSS.n4726 0.04025
R13341 VSS.n4728 VSS.n4727 0.04025
R13342 VSS.n4728 VSS.n2988 0.04025
R13343 VSS.n4732 VSS.n2988 0.04025
R13344 VSS.n4733 VSS.n4732 0.04025
R13345 VSS.n4734 VSS.n4733 0.04025
R13346 VSS.n4734 VSS.n2986 0.04025
R13347 VSS.n4738 VSS.n2986 0.04025
R13348 VSS.n4739 VSS.n4738 0.04025
R13349 VSS.n4740 VSS.n4739 0.04025
R13350 VSS.n4740 VSS.n2984 0.04025
R13351 VSS.n4744 VSS.n2984 0.04025
R13352 VSS.n4745 VSS.n4744 0.04025
R13353 VSS.n4746 VSS.n4745 0.04025
R13354 VSS.n4746 VSS.n2982 0.04025
R13355 VSS.n4750 VSS.n2982 0.04025
R13356 VSS.n4751 VSS.n4750 0.04025
R13357 VSS.n4752 VSS.n4751 0.04025
R13358 VSS.n4752 VSS.n2980 0.04025
R13359 VSS.n4756 VSS.n2980 0.04025
R13360 VSS.n4757 VSS.n4756 0.04025
R13361 VSS.n4758 VSS.n4757 0.04025
R13362 VSS.n4758 VSS.n2978 0.04025
R13363 VSS.n4762 VSS.n2978 0.04025
R13364 VSS.n4763 VSS.n4762 0.04025
R13365 VSS.n4764 VSS.n4763 0.04025
R13366 VSS.n4764 VSS.n2976 0.04025
R13367 VSS.n4768 VSS.n2976 0.04025
R13368 VSS.n4769 VSS.n4768 0.04025
R13369 VSS.n4770 VSS.n4769 0.04025
R13370 VSS.n4770 VSS.n2974 0.04025
R13371 VSS.n4774 VSS.n2974 0.04025
R13372 VSS.n4775 VSS.n4774 0.04025
R13373 VSS.n4776 VSS.n4775 0.04025
R13374 VSS.n4776 VSS.n2972 0.04025
R13375 VSS.n4780 VSS.n2972 0.04025
R13376 VSS.n4781 VSS.n4780 0.04025
R13377 VSS.n4782 VSS.n4781 0.04025
R13378 VSS.n4782 VSS.n2970 0.04025
R13379 VSS.n4786 VSS.n2970 0.04025
R13380 VSS.n4787 VSS.n4786 0.04025
R13381 VSS.n4788 VSS.n4787 0.04025
R13382 VSS.n4788 VSS.n2968 0.04025
R13383 VSS.n4792 VSS.n2968 0.04025
R13384 VSS.n4793 VSS.n4792 0.04025
R13385 VSS.n4794 VSS.n4793 0.04025
R13386 VSS.n4794 VSS.n2966 0.04025
R13387 VSS.n4798 VSS.n2966 0.04025
R13388 VSS.n4799 VSS.n4798 0.04025
R13389 VSS.n4800 VSS.n4799 0.04025
R13390 VSS.n4800 VSS.n2964 0.04025
R13391 VSS.n4807 VSS.n2964 0.04025
R13392 VSS.n4808 VSS.n4807 0.04025
R13393 VSS.n4809 VSS.n4808 0.04025
R13394 VSS.n4809 VSS.n2962 0.04025
R13395 VSS.n4813 VSS.n2962 0.04025
R13396 VSS.n4814 VSS.n4813 0.04025
R13397 VSS.n4815 VSS.n4814 0.04025
R13398 VSS.n4815 VSS.n2960 0.04025
R13399 VSS.n4819 VSS.n2960 0.04025
R13400 VSS.n4820 VSS.n4819 0.04025
R13401 VSS.n4821 VSS.n4820 0.04025
R13402 VSS.n4821 VSS.n2958 0.04025
R13403 VSS.n4825 VSS.n2958 0.04025
R13404 VSS.n4826 VSS.n4825 0.04025
R13405 VSS.n4827 VSS.n4826 0.04025
R13406 VSS.n4827 VSS.n2956 0.04025
R13407 VSS.n4831 VSS.n2956 0.04025
R13408 VSS.n4832 VSS.n4831 0.04025
R13409 VSS.n4833 VSS.n4832 0.04025
R13410 VSS.n4833 VSS.n2954 0.04025
R13411 VSS.n4837 VSS.n2954 0.04025
R13412 VSS.n4838 VSS.n4837 0.04025
R13413 VSS.n4839 VSS.n4838 0.04025
R13414 VSS.n4839 VSS.n2952 0.04025
R13415 VSS.n4843 VSS.n2952 0.04025
R13416 VSS.n4844 VSS.n4843 0.04025
R13417 VSS.n4845 VSS.n4844 0.04025
R13418 VSS.n4845 VSS.n2950 0.04025
R13419 VSS.n4849 VSS.n2950 0.04025
R13420 VSS.n4850 VSS.n4849 0.04025
R13421 VSS.n4851 VSS.n4850 0.04025
R13422 VSS.n4851 VSS.n2948 0.04025
R13423 VSS.n4855 VSS.n2948 0.04025
R13424 VSS.n4856 VSS.n4855 0.04025
R13425 VSS.n4857 VSS.n4856 0.04025
R13426 VSS.n4857 VSS.n2946 0.04025
R13427 VSS.n4861 VSS.n2946 0.04025
R13428 VSS.n4862 VSS.n4861 0.04025
R13429 VSS.n4863 VSS.n4862 0.04025
R13430 VSS.n4863 VSS.n2944 0.04025
R13431 VSS.n4867 VSS.n2944 0.04025
R13432 VSS.n4868 VSS.n4867 0.04025
R13433 VSS.n4869 VSS.n4868 0.04025
R13434 VSS.n4869 VSS.n2942 0.04025
R13435 VSS.n4873 VSS.n2942 0.04025
R13436 VSS.n4874 VSS.n4873 0.04025
R13437 VSS.n4875 VSS.n4874 0.04025
R13438 VSS.n4875 VSS.n2940 0.04025
R13439 VSS.n4879 VSS.n2940 0.04025
R13440 VSS.n4880 VSS.n4879 0.04025
R13441 VSS.n4881 VSS.n4880 0.04025
R13442 VSS.n4881 VSS.n2938 0.04025
R13443 VSS.n4885 VSS.n2938 0.04025
R13444 VSS.n4886 VSS.n4885 0.04025
R13445 VSS.n4887 VSS.n4886 0.04025
R13446 VSS.n4887 VSS.n2936 0.04025
R13447 VSS.n4891 VSS.n2936 0.04025
R13448 VSS.n4892 VSS.n4891 0.04025
R13449 VSS.n4893 VSS.n4892 0.04025
R13450 VSS.n4893 VSS.n2934 0.04025
R13451 VSS.n4897 VSS.n2934 0.04025
R13452 VSS.n4898 VSS.n4897 0.04025
R13453 VSS.n4899 VSS.n4898 0.04025
R13454 VSS.n4899 VSS.n2932 0.04025
R13455 VSS.n4903 VSS.n2932 0.04025
R13456 VSS.n4904 VSS.n4903 0.04025
R13457 VSS.n4905 VSS.n4904 0.04025
R13458 VSS.n4905 VSS.n2930 0.04025
R13459 VSS.n4909 VSS.n2930 0.04025
R13460 VSS.n4910 VSS.n4909 0.04025
R13461 VSS.n4911 VSS.n4910 0.04025
R13462 VSS.n4911 VSS.n2928 0.04025
R13463 VSS.n4915 VSS.n2928 0.04025
R13464 VSS.n4916 VSS.n4915 0.04025
R13465 VSS.n4917 VSS.n4916 0.04025
R13466 VSS.n4917 VSS.n2926 0.04025
R13467 VSS.n4921 VSS.n2926 0.04025
R13468 VSS.n4922 VSS.n4921 0.04025
R13469 VSS.n4923 VSS.n4922 0.04025
R13470 VSS.n4923 VSS.n2924 0.04025
R13471 VSS.n4927 VSS.n2924 0.04025
R13472 VSS.n4928 VSS.n4927 0.04025
R13473 VSS.n4929 VSS.n4928 0.04025
R13474 VSS.n4929 VSS.n2922 0.04025
R13475 VSS.n4933 VSS.n2922 0.04025
R13476 VSS.n4934 VSS.n4933 0.04025
R13477 VSS.n4935 VSS.n4934 0.04025
R13478 VSS.n4935 VSS.n2920 0.04025
R13479 VSS.n4939 VSS.n2920 0.04025
R13480 VSS.n4940 VSS.n4939 0.04025
R13481 VSS.n4941 VSS.n4940 0.04025
R13482 VSS.n4941 VSS.n2918 0.04025
R13483 VSS.n4945 VSS.n2918 0.04025
R13484 VSS.n4946 VSS.n4945 0.04025
R13485 VSS.n4947 VSS.n4946 0.04025
R13486 VSS.n4947 VSS.n2916 0.04025
R13487 VSS.n4951 VSS.n2916 0.04025
R13488 VSS.n4952 VSS.n4951 0.04025
R13489 VSS.n4953 VSS.n4952 0.04025
R13490 VSS.n4953 VSS.n2914 0.04025
R13491 VSS.n4957 VSS.n2914 0.04025
R13492 VSS.n4958 VSS.n4957 0.04025
R13493 VSS.n4959 VSS.n4958 0.04025
R13494 VSS.n4959 VSS.n2912 0.04025
R13495 VSS.n4963 VSS.n2912 0.04025
R13496 VSS.n4964 VSS.n4963 0.04025
R13497 VSS.n4965 VSS.n4964 0.04025
R13498 VSS.n4965 VSS.n2910 0.04025
R13499 VSS.n4969 VSS.n2910 0.04025
R13500 VSS.n4970 VSS.n4969 0.04025
R13501 VSS.n4971 VSS.n4970 0.04025
R13502 VSS.n4971 VSS.n2908 0.04025
R13503 VSS.n4975 VSS.n2908 0.04025
R13504 VSS.n4976 VSS.n4975 0.04025
R13505 VSS.n4977 VSS.n4976 0.04025
R13506 VSS.n4977 VSS.n2906 0.04025
R13507 VSS.n4981 VSS.n2906 0.04025
R13508 VSS.n4982 VSS.n4981 0.04025
R13509 VSS.n4983 VSS.n4982 0.04025
R13510 VSS.n4983 VSS.n2904 0.04025
R13511 VSS.n4987 VSS.n2904 0.04025
R13512 VSS.n4988 VSS.n4987 0.04025
R13513 VSS.n4989 VSS.n4988 0.04025
R13514 VSS.n4989 VSS.n2902 0.04025
R13515 VSS.n4993 VSS.n2902 0.04025
R13516 VSS.n4994 VSS.n4993 0.04025
R13517 VSS.n4995 VSS.n4994 0.04025
R13518 VSS.n4995 VSS.n2900 0.04025
R13519 VSS.n4999 VSS.n2900 0.04025
R13520 VSS.n5000 VSS.n4999 0.04025
R13521 VSS.n5001 VSS.n5000 0.04025
R13522 VSS.n5001 VSS.n2898 0.04025
R13523 VSS.n5005 VSS.n2898 0.04025
R13524 VSS.n5006 VSS.n5005 0.04025
R13525 VSS.n5007 VSS.n5006 0.04025
R13526 VSS.n5007 VSS.n2896 0.04025
R13527 VSS.n5011 VSS.n2896 0.04025
R13528 VSS.n5012 VSS.n5011 0.04025
R13529 VSS.n5013 VSS.n5012 0.04025
R13530 VSS.n5013 VSS.n2894 0.04025
R13531 VSS.n5017 VSS.n2894 0.04025
R13532 VSS.n5018 VSS.n5017 0.04025
R13533 VSS.n5019 VSS.n5018 0.04025
R13534 VSS.n5019 VSS.n2892 0.04025
R13535 VSS.n5023 VSS.n2892 0.04025
R13536 VSS.n5024 VSS.n5023 0.04025
R13537 VSS.n5025 VSS.n5024 0.04025
R13538 VSS.n5025 VSS.n2890 0.04025
R13539 VSS.n5029 VSS.n2890 0.04025
R13540 VSS.n5030 VSS.n5029 0.04025
R13541 VSS.n5031 VSS.n5030 0.04025
R13542 VSS.n5031 VSS.n2888 0.04025
R13543 VSS.n5035 VSS.n2888 0.04025
R13544 VSS.n5036 VSS.n5035 0.04025
R13545 VSS.n5037 VSS.n5036 0.04025
R13546 VSS.n5037 VSS.n2886 0.04025
R13547 VSS.n5041 VSS.n2886 0.04025
R13548 VSS.n5042 VSS.n5041 0.04025
R13549 VSS.n5043 VSS.n5042 0.04025
R13550 VSS.n5043 VSS.n2884 0.04025
R13551 VSS.n5047 VSS.n2884 0.04025
R13552 VSS.n5048 VSS.n5047 0.04025
R13553 VSS.n5049 VSS.n5048 0.04025
R13554 VSS.n5049 VSS.n2882 0.04025
R13555 VSS.n5053 VSS.n2882 0.04025
R13556 VSS.n5054 VSS.n5053 0.04025
R13557 VSS.n5055 VSS.n5054 0.04025
R13558 VSS.n5055 VSS.n2880 0.04025
R13559 VSS.n5059 VSS.n2880 0.04025
R13560 VSS.n5060 VSS.n5059 0.04025
R13561 VSS.n5061 VSS.n5060 0.04025
R13562 VSS.n5061 VSS.n2878 0.04025
R13563 VSS.n5065 VSS.n2878 0.04025
R13564 VSS.n5066 VSS.n5065 0.04025
R13565 VSS.n5067 VSS.n5066 0.04025
R13566 VSS.n5067 VSS.n2876 0.04025
R13567 VSS.n5071 VSS.n2876 0.04025
R13568 VSS.n5072 VSS.n5071 0.04025
R13569 VSS.n5073 VSS.n5072 0.04025
R13570 VSS.n5073 VSS.n2874 0.04025
R13571 VSS.n5077 VSS.n2874 0.04025
R13572 VSS.n5078 VSS.n5077 0.04025
R13573 VSS.n5079 VSS.n5078 0.04025
R13574 VSS.n5079 VSS.n2872 0.04025
R13575 VSS.n5083 VSS.n2872 0.04025
R13576 VSS.n5084 VSS.n5083 0.04025
R13577 VSS.n5085 VSS.n5084 0.04025
R13578 VSS.n5085 VSS.n2870 0.04025
R13579 VSS.n5089 VSS.n2870 0.04025
R13580 VSS.n5090 VSS.n5089 0.04025
R13581 VSS.n5091 VSS.n5090 0.04025
R13582 VSS.n5091 VSS.n2868 0.04025
R13583 VSS.n5095 VSS.n2868 0.04025
R13584 VSS.n5096 VSS.n5095 0.04025
R13585 VSS.n5097 VSS.n5096 0.04025
R13586 VSS.n5097 VSS.n2866 0.04025
R13587 VSS.n5101 VSS.n2866 0.04025
R13588 VSS.n5102 VSS.n5101 0.04025
R13589 VSS.n5103 VSS.n5102 0.04025
R13590 VSS.n5103 VSS.n2864 0.04025
R13591 VSS.n5107 VSS.n2864 0.04025
R13592 VSS.n5108 VSS.n5107 0.04025
R13593 VSS.n5109 VSS.n5108 0.04025
R13594 VSS.n5109 VSS.n2862 0.04025
R13595 VSS.n5113 VSS.n2862 0.04025
R13596 VSS.n5114 VSS.n5113 0.04025
R13597 VSS.n5115 VSS.n5114 0.04025
R13598 VSS.n5115 VSS.n2860 0.04025
R13599 VSS.n5119 VSS.n2860 0.04025
R13600 VSS.n5120 VSS.n5119 0.04025
R13601 VSS.n5121 VSS.n5120 0.04025
R13602 VSS.n5121 VSS.n2858 0.04025
R13603 VSS.n5125 VSS.n2858 0.04025
R13604 VSS.n5126 VSS.n5125 0.04025
R13605 VSS.n5127 VSS.n5126 0.04025
R13606 VSS.n5127 VSS.n2856 0.04025
R13607 VSS.n5131 VSS.n2856 0.04025
R13608 VSS.n5132 VSS.n5131 0.04025
R13609 VSS.n5133 VSS.n5132 0.04025
R13610 VSS.n5133 VSS.n2854 0.04025
R13611 VSS.n5137 VSS.n2854 0.04025
R13612 VSS.n5138 VSS.n5137 0.04025
R13613 VSS.n5139 VSS.n5138 0.04025
R13614 VSS.n5139 VSS.n2852 0.04025
R13615 VSS.n5143 VSS.n2852 0.04025
R13616 VSS.n5144 VSS.n5143 0.04025
R13617 VSS.n5145 VSS.n5144 0.04025
R13618 VSS.n5145 VSS.n2850 0.04025
R13619 VSS.n5149 VSS.n2850 0.04025
R13620 VSS.n5150 VSS.n5149 0.04025
R13621 VSS.n5151 VSS.n5150 0.04025
R13622 VSS.n5151 VSS.n2848 0.04025
R13623 VSS.n5155 VSS.n2848 0.04025
R13624 VSS.n5156 VSS.n5155 0.04025
R13625 VSS.n5157 VSS.n5156 0.04025
R13626 VSS.n5157 VSS.n2846 0.04025
R13627 VSS.n5161 VSS.n2846 0.04025
R13628 VSS.n5162 VSS.n5161 0.04025
R13629 VSS.n5163 VSS.n5162 0.04025
R13630 VSS.n5163 VSS.n2844 0.04025
R13631 VSS.n5167 VSS.n2844 0.04025
R13632 VSS.n5168 VSS.n5167 0.04025
R13633 VSS.n5169 VSS.n5168 0.04025
R13634 VSS.n5169 VSS.n2842 0.04025
R13635 VSS.n5173 VSS.n2842 0.04025
R13636 VSS.n5174 VSS.n5173 0.04025
R13637 VSS.n5175 VSS.n5174 0.04025
R13638 VSS.n5175 VSS.n2840 0.04025
R13639 VSS.n5179 VSS.n2840 0.04025
R13640 VSS.n5180 VSS.n5179 0.04025
R13641 VSS.n5181 VSS.n5180 0.04025
R13642 VSS.n5181 VSS.n2838 0.04025
R13643 VSS.n5185 VSS.n2838 0.04025
R13644 VSS.n5186 VSS.n5185 0.04025
R13645 VSS.n5187 VSS.n5186 0.04025
R13646 VSS.n5187 VSS.n2836 0.04025
R13647 VSS.n5191 VSS.n2836 0.04025
R13648 VSS.n5192 VSS.n5191 0.04025
R13649 VSS.n5193 VSS.n5192 0.04025
R13650 VSS.n5193 VSS.n2834 0.04025
R13651 VSS.n5197 VSS.n2834 0.04025
R13652 VSS.n5198 VSS.n5197 0.04025
R13653 VSS.n5199 VSS.n5198 0.04025
R13654 VSS.n5199 VSS.n2832 0.04025
R13655 VSS.n5203 VSS.n2832 0.04025
R13656 VSS.n5204 VSS.n5203 0.04025
R13657 VSS.n5205 VSS.n5204 0.04025
R13658 VSS.n5205 VSS.n2830 0.04025
R13659 VSS.n5209 VSS.n2830 0.04025
R13660 VSS.n5210 VSS.n5209 0.04025
R13661 VSS.n5211 VSS.n5210 0.04025
R13662 VSS.n5211 VSS.n2828 0.04025
R13663 VSS.n5215 VSS.n2828 0.04025
R13664 VSS.n5216 VSS.n5215 0.04025
R13665 VSS.n5217 VSS.n5216 0.04025
R13666 VSS.n5217 VSS.n2826 0.04025
R13667 VSS.n5221 VSS.n2826 0.04025
R13668 VSS.n5222 VSS.n5221 0.04025
R13669 VSS.n5223 VSS.n5222 0.04025
R13670 VSS.n5223 VSS.n2824 0.04025
R13671 VSS.n5227 VSS.n2824 0.04025
R13672 VSS.n5228 VSS.n5227 0.04025
R13673 VSS.n5229 VSS.n5228 0.04025
R13674 VSS.n5229 VSS.n2822 0.04025
R13675 VSS.n5233 VSS.n2822 0.04025
R13676 VSS.n5234 VSS.n5233 0.04025
R13677 VSS.n5235 VSS.n5234 0.04025
R13678 VSS.n5235 VSS.n2820 0.04025
R13679 VSS.n5239 VSS.n2820 0.04025
R13680 VSS.n5240 VSS.n5239 0.04025
R13681 VSS.n5241 VSS.n5240 0.04025
R13682 VSS.n5241 VSS.n2818 0.04025
R13683 VSS.n5245 VSS.n2818 0.04025
R13684 VSS.n5246 VSS.n5245 0.04025
R13685 VSS.n5247 VSS.n5246 0.04025
R13686 VSS.n5247 VSS.n2816 0.04025
R13687 VSS.n5251 VSS.n2816 0.04025
R13688 VSS.n5252 VSS.n5251 0.04025
R13689 VSS.n5253 VSS.n5252 0.04025
R13690 VSS.n5253 VSS.n2814 0.04025
R13691 VSS.n5257 VSS.n2814 0.04025
R13692 VSS.n5258 VSS.n5257 0.04025
R13693 VSS.n5259 VSS.n5258 0.04025
R13694 VSS.n5259 VSS.n2812 0.04025
R13695 VSS.n5263 VSS.n2812 0.04025
R13696 VSS.n5264 VSS.n5263 0.04025
R13697 VSS.n5265 VSS.n5264 0.04025
R13698 VSS.n5265 VSS.n2810 0.04025
R13699 VSS.n5269 VSS.n2810 0.04025
R13700 VSS.n5270 VSS.n5269 0.04025
R13701 VSS.n5271 VSS.n5270 0.04025
R13702 VSS.n5271 VSS.n2808 0.04025
R13703 VSS.n5275 VSS.n2808 0.04025
R13704 VSS.n5276 VSS.n5275 0.04025
R13705 VSS.n5277 VSS.n5276 0.04025
R13706 VSS.n5277 VSS.n2806 0.04025
R13707 VSS.n5281 VSS.n2806 0.04025
R13708 VSS.n5282 VSS.n5281 0.04025
R13709 VSS.n5283 VSS.n5282 0.04025
R13710 VSS.n5283 VSS.n2804 0.04025
R13711 VSS.n5287 VSS.n2804 0.04025
R13712 VSS.n5288 VSS.n5287 0.04025
R13713 VSS.n5289 VSS.n5288 0.04025
R13714 VSS.n5289 VSS.n2802 0.04025
R13715 VSS.n5293 VSS.n2802 0.04025
R13716 VSS.n5294 VSS.n5293 0.04025
R13717 VSS.n5295 VSS.n5294 0.04025
R13718 VSS.n5295 VSS.n2800 0.04025
R13719 VSS.n5299 VSS.n2800 0.04025
R13720 VSS.n5300 VSS.n5299 0.04025
R13721 VSS.n5301 VSS.n5300 0.04025
R13722 VSS.n5301 VSS.n2798 0.04025
R13723 VSS.n5305 VSS.n2798 0.04025
R13724 VSS.n5306 VSS.n5305 0.04025
R13725 VSS.n5307 VSS.n5306 0.04025
R13726 VSS.n5307 VSS.n2796 0.04025
R13727 VSS.n5311 VSS.n2796 0.04025
R13728 VSS.n5312 VSS.n5311 0.04025
R13729 VSS.n5313 VSS.n5312 0.04025
R13730 VSS.n5313 VSS.n2794 0.04025
R13731 VSS.n5317 VSS.n2794 0.04025
R13732 VSS.n5318 VSS.n5317 0.04025
R13733 VSS.n5319 VSS.n5318 0.04025
R13734 VSS.n5319 VSS.n2792 0.04025
R13735 VSS.n5323 VSS.n2792 0.04025
R13736 VSS.n5324 VSS.n5323 0.04025
R13737 VSS.n5325 VSS.n5324 0.04025
R13738 VSS.n5325 VSS.n2790 0.04025
R13739 VSS.n5329 VSS.n2790 0.04025
R13740 VSS.n5330 VSS.n5329 0.04025
R13741 VSS.n5331 VSS.n5330 0.04025
R13742 VSS.n5331 VSS.n2788 0.04025
R13743 VSS.n5335 VSS.n2788 0.04025
R13744 VSS.n5336 VSS.n5335 0.04025
R13745 VSS.n5337 VSS.n5336 0.04025
R13746 VSS.n5337 VSS.n2786 0.04025
R13747 VSS.n5341 VSS.n2786 0.04025
R13748 VSS.n5342 VSS.n5341 0.04025
R13749 VSS.n5343 VSS.n5342 0.04025
R13750 VSS.n5343 VSS.n2784 0.04025
R13751 VSS.n5347 VSS.n2784 0.04025
R13752 VSS.n5348 VSS.n5347 0.04025
R13753 VSS.n5349 VSS.n5348 0.04025
R13754 VSS.n5349 VSS.n2782 0.04025
R13755 VSS.n5353 VSS.n2782 0.04025
R13756 VSS.n5354 VSS.n5353 0.04025
R13757 VSS.n5355 VSS.n5354 0.04025
R13758 VSS.n5355 VSS.n2780 0.04025
R13759 VSS.n5359 VSS.n2780 0.04025
R13760 VSS.n5360 VSS.n5359 0.04025
R13761 VSS.n5361 VSS.n5360 0.04025
R13762 VSS.n5361 VSS.n2778 0.04025
R13763 VSS.n5365 VSS.n2778 0.04025
R13764 VSS.n5366 VSS.n5365 0.04025
R13765 VSS.n5367 VSS.n5366 0.04025
R13766 VSS.n5367 VSS.n2776 0.04025
R13767 VSS.n5371 VSS.n2776 0.04025
R13768 VSS.n5372 VSS.n5371 0.04025
R13769 VSS.n5373 VSS.n5372 0.04025
R13770 VSS.n5373 VSS.n2774 0.04025
R13771 VSS.n5377 VSS.n2774 0.04025
R13772 VSS.n5378 VSS.n5377 0.04025
R13773 VSS.n5379 VSS.n5378 0.04025
R13774 VSS.n5379 VSS.n2772 0.04025
R13775 VSS.n5383 VSS.n2772 0.04025
R13776 VSS.n5384 VSS.n5383 0.04025
R13777 VSS.n5385 VSS.n5384 0.04025
R13778 VSS.n5385 VSS.n2770 0.04025
R13779 VSS.n5389 VSS.n2770 0.04025
R13780 VSS.n5390 VSS.n5389 0.04025
R13781 VSS.n5391 VSS.n5390 0.04025
R13782 VSS.n5391 VSS.n2768 0.04025
R13783 VSS.n5395 VSS.n2768 0.04025
R13784 VSS.n5396 VSS.n5395 0.04025
R13785 VSS.n5397 VSS.n5396 0.04025
R13786 VSS.n5397 VSS.n2766 0.04025
R13787 VSS.n5401 VSS.n2766 0.04025
R13788 VSS.n5402 VSS.n5401 0.04025
R13789 VSS.n5403 VSS.n5402 0.04025
R13790 VSS.n5403 VSS.n2764 0.04025
R13791 VSS.n5407 VSS.n2764 0.04025
R13792 VSS.n5408 VSS.n5407 0.04025
R13793 VSS.n5409 VSS.n5408 0.04025
R13794 VSS.n5409 VSS.n2762 0.04025
R13795 VSS.n5413 VSS.n2762 0.04025
R13796 VSS.n5414 VSS.n5413 0.04025
R13797 VSS.n5415 VSS.n5414 0.04025
R13798 VSS.n5415 VSS.n2760 0.04025
R13799 VSS.n5419 VSS.n2760 0.04025
R13800 VSS.n5420 VSS.n5419 0.04025
R13801 VSS.n5421 VSS.n5420 0.04025
R13802 VSS.n5421 VSS.n2758 0.04025
R13803 VSS.n5425 VSS.n2758 0.04025
R13804 VSS.n5426 VSS.n5425 0.04025
R13805 VSS.n5427 VSS.n5426 0.04025
R13806 VSS.n5427 VSS.n2756 0.04025
R13807 VSS.n5431 VSS.n2756 0.04025
R13808 VSS.n5432 VSS.n5431 0.04025
R13809 VSS.n5433 VSS.n5432 0.04025
R13810 VSS.n5433 VSS.n2754 0.04025
R13811 VSS.n5437 VSS.n2754 0.04025
R13812 VSS.n5438 VSS.n5437 0.04025
R13813 VSS.n5439 VSS.n5438 0.04025
R13814 VSS.n5439 VSS.n2752 0.04025
R13815 VSS.n5443 VSS.n2752 0.04025
R13816 VSS.n5444 VSS.n5443 0.04025
R13817 VSS.n5445 VSS.n5444 0.04025
R13818 VSS.n5445 VSS.n2750 0.04025
R13819 VSS.n5449 VSS.n2750 0.04025
R13820 VSS.n5450 VSS.n5449 0.04025
R13821 VSS.n5451 VSS.n5450 0.04025
R13822 VSS.n5451 VSS.n2748 0.04025
R13823 VSS.n5455 VSS.n2748 0.04025
R13824 VSS.n5456 VSS.n5455 0.04025
R13825 VSS.n5457 VSS.n5456 0.04025
R13826 VSS.n5457 VSS.n2746 0.04025
R13827 VSS.n5461 VSS.n2746 0.04025
R13828 VSS.n5462 VSS.n5461 0.04025
R13829 VSS.n5463 VSS.n5462 0.04025
R13830 VSS.n5463 VSS.n2744 0.04025
R13831 VSS.n5467 VSS.n2744 0.04025
R13832 VSS.n5468 VSS.n5467 0.04025
R13833 VSS.n4143 VSS.n4142 0.04025
R13834 VSS.n4143 VSS.n3183 0.04025
R13835 VSS.n4147 VSS.n3183 0.04025
R13836 VSS.n4148 VSS.n4147 0.04025
R13837 VSS.n4149 VSS.n4148 0.04025
R13838 VSS.n4149 VSS.n3181 0.04025
R13839 VSS.n4153 VSS.n3181 0.04025
R13840 VSS.n4154 VSS.n4153 0.04025
R13841 VSS.n4155 VSS.n4154 0.04025
R13842 VSS.n4155 VSS.n3179 0.04025
R13843 VSS.n4159 VSS.n3179 0.04025
R13844 VSS.n4160 VSS.n4159 0.04025
R13845 VSS.n4161 VSS.n4160 0.04025
R13846 VSS.n4161 VSS.n3177 0.04025
R13847 VSS.n4165 VSS.n3177 0.04025
R13848 VSS.n4166 VSS.n4165 0.04025
R13849 VSS.n4167 VSS.n4166 0.04025
R13850 VSS.n4167 VSS.n3175 0.04025
R13851 VSS.n4171 VSS.n3175 0.04025
R13852 VSS.n4172 VSS.n4171 0.04025
R13853 VSS.n4173 VSS.n4172 0.04025
R13854 VSS.n4173 VSS.n3173 0.04025
R13855 VSS.n4177 VSS.n3173 0.04025
R13856 VSS.n4178 VSS.n4177 0.04025
R13857 VSS.n4179 VSS.n4178 0.04025
R13858 VSS.n4179 VSS.n3171 0.04025
R13859 VSS.n4183 VSS.n3171 0.04025
R13860 VSS.n4184 VSS.n4183 0.04025
R13861 VSS.n4185 VSS.n4184 0.04025
R13862 VSS.n4185 VSS.n3169 0.04025
R13863 VSS.n4189 VSS.n3169 0.04025
R13864 VSS.n4190 VSS.n4189 0.04025
R13865 VSS.n4191 VSS.n4190 0.04025
R13866 VSS.n4191 VSS.n3167 0.04025
R13867 VSS.n4195 VSS.n3167 0.04025
R13868 VSS.n4196 VSS.n4195 0.04025
R13869 VSS.n4197 VSS.n4196 0.04025
R13870 VSS.n4197 VSS.n3165 0.04025
R13871 VSS.n4201 VSS.n3165 0.04025
R13872 VSS.n4202 VSS.n4201 0.04025
R13873 VSS.n4203 VSS.n4202 0.04025
R13874 VSS.n4203 VSS.n3163 0.04025
R13875 VSS.n4207 VSS.n3163 0.04025
R13876 VSS.n4208 VSS.n4207 0.04025
R13877 VSS.n4209 VSS.n4208 0.04025
R13878 VSS.n4209 VSS.n3161 0.04025
R13879 VSS.n4213 VSS.n3161 0.04025
R13880 VSS.n4214 VSS.n4213 0.04025
R13881 VSS.n4215 VSS.n4214 0.04025
R13882 VSS.n4215 VSS.n3159 0.04025
R13883 VSS.n4219 VSS.n3159 0.04025
R13884 VSS.n4220 VSS.n4219 0.04025
R13885 VSS.n4221 VSS.n4220 0.04025
R13886 VSS.n4221 VSS.n3157 0.04025
R13887 VSS.n4225 VSS.n3157 0.04025
R13888 VSS.n4226 VSS.n4225 0.04025
R13889 VSS.n4227 VSS.n4226 0.04025
R13890 VSS.n4227 VSS.n3155 0.04025
R13891 VSS.n4231 VSS.n3155 0.04025
R13892 VSS.n4232 VSS.n4231 0.04025
R13893 VSS.n4233 VSS.n4232 0.04025
R13894 VSS.n4233 VSS.n3153 0.04025
R13895 VSS.n4237 VSS.n3153 0.04025
R13896 VSS.n4238 VSS.n4237 0.04025
R13897 VSS.n4239 VSS.n4238 0.04025
R13898 VSS.n4239 VSS.n3151 0.04025
R13899 VSS.n4243 VSS.n3151 0.04025
R13900 VSS.n4244 VSS.n4243 0.04025
R13901 VSS.n4245 VSS.n4244 0.04025
R13902 VSS.n4245 VSS.n3149 0.04025
R13903 VSS.n4249 VSS.n3149 0.04025
R13904 VSS.n4250 VSS.n4249 0.04025
R13905 VSS.n4251 VSS.n4250 0.04025
R13906 VSS.n4251 VSS.n3147 0.04025
R13907 VSS.n4255 VSS.n3147 0.04025
R13908 VSS.n4256 VSS.n4255 0.04025
R13909 VSS.n4257 VSS.n4256 0.04025
R13910 VSS.n4257 VSS.n3145 0.04025
R13911 VSS.n4261 VSS.n3145 0.04025
R13912 VSS.n4262 VSS.n4261 0.04025
R13913 VSS.n4263 VSS.n4262 0.04025
R13914 VSS.n4263 VSS.n3143 0.04025
R13915 VSS.n4267 VSS.n3143 0.04025
R13916 VSS.n4268 VSS.n4267 0.04025
R13917 VSS.n4269 VSS.n4268 0.04025
R13918 VSS.n4269 VSS.n3141 0.04025
R13919 VSS.n4273 VSS.n3141 0.04025
R13920 VSS.n4274 VSS.n4273 0.04025
R13921 VSS.n4275 VSS.n4274 0.04025
R13922 VSS.n4275 VSS.n3139 0.04025
R13923 VSS.n4279 VSS.n3139 0.04025
R13924 VSS.n4280 VSS.n4279 0.04025
R13925 VSS.n4281 VSS.n4280 0.04025
R13926 VSS.n4281 VSS.n3137 0.04025
R13927 VSS.n4285 VSS.n3137 0.04025
R13928 VSS.n4286 VSS.n4285 0.04025
R13929 VSS.n4287 VSS.n4286 0.04025
R13930 VSS.n4287 VSS.n3135 0.04025
R13931 VSS.n4291 VSS.n3135 0.04025
R13932 VSS.n4292 VSS.n4291 0.04025
R13933 VSS.n4293 VSS.n4292 0.04025
R13934 VSS.n4293 VSS.n3133 0.04025
R13935 VSS.n4297 VSS.n3133 0.04025
R13936 VSS.n4298 VSS.n4297 0.04025
R13937 VSS.n4299 VSS.n4298 0.04025
R13938 VSS.n4299 VSS.n3131 0.04025
R13939 VSS.n4303 VSS.n3131 0.04025
R13940 VSS.n4304 VSS.n4303 0.04025
R13941 VSS.n4305 VSS.n4304 0.04025
R13942 VSS.n4305 VSS.n3129 0.04025
R13943 VSS.n4309 VSS.n3129 0.04025
R13944 VSS.n4310 VSS.n4309 0.04025
R13945 VSS.n4311 VSS.n4310 0.04025
R13946 VSS.n4311 VSS.n3127 0.04025
R13947 VSS.n4315 VSS.n3127 0.04025
R13948 VSS.n4316 VSS.n4315 0.04025
R13949 VSS.n4317 VSS.n4316 0.04025
R13950 VSS.n4317 VSS.n3125 0.04025
R13951 VSS.n4321 VSS.n3125 0.04025
R13952 VSS.n4322 VSS.n4321 0.04025
R13953 VSS.n4323 VSS.n4322 0.04025
R13954 VSS.n4323 VSS.n3123 0.04025
R13955 VSS.n4327 VSS.n3123 0.04025
R13956 VSS.n4328 VSS.n4327 0.04025
R13957 VSS.n4329 VSS.n4328 0.04025
R13958 VSS.n4329 VSS.n3121 0.04025
R13959 VSS.n4333 VSS.n3121 0.04025
R13960 VSS.n4334 VSS.n4333 0.04025
R13961 VSS.n4335 VSS.n4334 0.04025
R13962 VSS.n4335 VSS.n3119 0.04025
R13963 VSS.n4339 VSS.n3119 0.04025
R13964 VSS.n4340 VSS.n4339 0.04025
R13965 VSS.n4341 VSS.n4340 0.04025
R13966 VSS.n4341 VSS.n3117 0.04025
R13967 VSS.n4345 VSS.n3117 0.04025
R13968 VSS.n4346 VSS.n4345 0.04025
R13969 VSS.n4347 VSS.n4346 0.04025
R13970 VSS.n4347 VSS.n3115 0.04025
R13971 VSS.n4351 VSS.n3115 0.04025
R13972 VSS.n4352 VSS.n4351 0.04025
R13973 VSS.n4353 VSS.n4352 0.04025
R13974 VSS.n4353 VSS.n3113 0.04025
R13975 VSS.n4357 VSS.n3113 0.04025
R13976 VSS.n4358 VSS.n4357 0.04025
R13977 VSS.n4359 VSS.n4358 0.04025
R13978 VSS.n4359 VSS.n3111 0.04025
R13979 VSS.n4363 VSS.n3111 0.04025
R13980 VSS.n4364 VSS.n4363 0.04025
R13981 VSS.n4365 VSS.n4364 0.04025
R13982 VSS.n4365 VSS.n3109 0.04025
R13983 VSS.n4369 VSS.n3109 0.04025
R13984 VSS.n4370 VSS.n4369 0.04025
R13985 VSS.n4371 VSS.n4370 0.04025
R13986 VSS.n4371 VSS.n3107 0.04025
R13987 VSS.n4375 VSS.n3107 0.04025
R13988 VSS.n4376 VSS.n4375 0.04025
R13989 VSS.n4377 VSS.n4376 0.04025
R13990 VSS.n4377 VSS.n3105 0.04025
R13991 VSS.n4381 VSS.n3105 0.04025
R13992 VSS.n4382 VSS.n4381 0.04025
R13993 VSS.n4383 VSS.n4382 0.04025
R13994 VSS.n4383 VSS.n3103 0.04025
R13995 VSS.n4387 VSS.n3103 0.04025
R13996 VSS.n4388 VSS.n4387 0.04025
R13997 VSS.n4389 VSS.n4388 0.04025
R13998 VSS.n4389 VSS.n3101 0.04025
R13999 VSS.n4393 VSS.n3101 0.04025
R14000 VSS.n4394 VSS.n4393 0.04025
R14001 VSS.n4395 VSS.n4394 0.04025
R14002 VSS.n4395 VSS.n3099 0.04025
R14003 VSS.n4399 VSS.n3099 0.04025
R14004 VSS.n4400 VSS.n4399 0.04025
R14005 VSS.n4401 VSS.n4400 0.04025
R14006 VSS.n4401 VSS.n3097 0.04025
R14007 VSS.n4405 VSS.n3097 0.04025
R14008 VSS.n4406 VSS.n4405 0.04025
R14009 VSS.n4407 VSS.n4406 0.04025
R14010 VSS.n4407 VSS.n3095 0.04025
R14011 VSS.n4411 VSS.n3095 0.04025
R14012 VSS.n4412 VSS.n4411 0.04025
R14013 VSS.n4413 VSS.n4412 0.04025
R14014 VSS.n4413 VSS.n3093 0.04025
R14015 VSS.n4417 VSS.n3093 0.04025
R14016 VSS.n4418 VSS.n4417 0.04025
R14017 VSS.n4419 VSS.n4418 0.04025
R14018 VSS.n4419 VSS.n3091 0.04025
R14019 VSS.n4423 VSS.n3091 0.04025
R14020 VSS.n4424 VSS.n4423 0.04025
R14021 VSS.n4425 VSS.n4424 0.04025
R14022 VSS.n4425 VSS.n3089 0.04025
R14023 VSS.n4429 VSS.n3089 0.04025
R14024 VSS.n4430 VSS.n4429 0.04025
R14025 VSS.n4431 VSS.n4430 0.04025
R14026 VSS.n4431 VSS.n3087 0.04025
R14027 VSS.n4435 VSS.n3087 0.04025
R14028 VSS.n4436 VSS.n4435 0.04025
R14029 VSS.n4437 VSS.n4436 0.04025
R14030 VSS.n4437 VSS.n3085 0.04025
R14031 VSS.n4441 VSS.n3085 0.04025
R14032 VSS.n4442 VSS.n4441 0.04025
R14033 VSS.n4443 VSS.n4442 0.04025
R14034 VSS.n4443 VSS.n3083 0.04025
R14035 VSS.n4447 VSS.n3083 0.04025
R14036 VSS.n4448 VSS.n4447 0.04025
R14037 VSS.n4449 VSS.n4448 0.04025
R14038 VSS.n4449 VSS.n3081 0.04025
R14039 VSS.n4453 VSS.n3081 0.04025
R14040 VSS.n4454 VSS.n4453 0.04025
R14041 VSS.n4455 VSS.n4454 0.04025
R14042 VSS.n4455 VSS.n3079 0.04025
R14043 VSS.n4459 VSS.n3079 0.04025
R14044 VSS.n4460 VSS.n4459 0.04025
R14045 VSS.n4461 VSS.n4460 0.04025
R14046 VSS.n4461 VSS.n3077 0.04025
R14047 VSS.n4465 VSS.n3077 0.04025
R14048 VSS.n4466 VSS.n4465 0.04025
R14049 VSS.n4467 VSS.n4466 0.04025
R14050 VSS.n4467 VSS.n3075 0.04025
R14051 VSS.n4471 VSS.n3075 0.04025
R14052 VSS.n4472 VSS.n4471 0.04025
R14053 VSS.n4473 VSS.n4472 0.04025
R14054 VSS.n4473 VSS.n3073 0.04025
R14055 VSS.n4477 VSS.n3073 0.04025
R14056 VSS.n4478 VSS.n4477 0.04025
R14057 VSS.n4479 VSS.n4478 0.04025
R14058 VSS.n4479 VSS.n3071 0.04025
R14059 VSS.n4483 VSS.n3071 0.04025
R14060 VSS.n4484 VSS.n4483 0.04025
R14061 VSS.n4485 VSS.n4484 0.04025
R14062 VSS.n4485 VSS.n3069 0.04025
R14063 VSS.n4489 VSS.n3069 0.04025
R14064 VSS.n4490 VSS.n4489 0.04025
R14065 VSS.n4491 VSS.n4490 0.04025
R14066 VSS.n4491 VSS.n3067 0.04025
R14067 VSS.n4495 VSS.n3067 0.04025
R14068 VSS.n4496 VSS.n4495 0.04025
R14069 VSS.n4497 VSS.n4496 0.04025
R14070 VSS.n4497 VSS.n3065 0.04025
R14071 VSS.n4501 VSS.n3065 0.04025
R14072 VSS.n4502 VSS.n4501 0.04025
R14073 VSS.n4503 VSS.n4502 0.04025
R14074 VSS.n4503 VSS.n3063 0.04025
R14075 VSS.n4507 VSS.n3063 0.04025
R14076 VSS.n4508 VSS.n4507 0.04025
R14077 VSS.n4509 VSS.n4508 0.04025
R14078 VSS.n4509 VSS.n3061 0.04025
R14079 VSS.n4513 VSS.n3061 0.04025
R14080 VSS.n4514 VSS.n4513 0.04025
R14081 VSS.n4515 VSS.n4514 0.04025
R14082 VSS.n4515 VSS.n3059 0.04025
R14083 VSS.n4519 VSS.n3059 0.04025
R14084 VSS.n4520 VSS.n4519 0.04025
R14085 VSS.n4521 VSS.n4520 0.04025
R14086 VSS.n4521 VSS.n3057 0.04025
R14087 VSS.n4525 VSS.n3057 0.04025
R14088 VSS.n4526 VSS.n4525 0.04025
R14089 VSS.n4527 VSS.n4526 0.04025
R14090 VSS.n4527 VSS.n3055 0.04025
R14091 VSS.n4531 VSS.n3055 0.04025
R14092 VSS.n4532 VSS.n4531 0.04025
R14093 VSS.n4533 VSS.n4532 0.04025
R14094 VSS.n4533 VSS.n3053 0.04025
R14095 VSS.n4537 VSS.n3053 0.04025
R14096 VSS.n4538 VSS.n4537 0.04025
R14097 VSS.n4539 VSS.n4538 0.04025
R14098 VSS.n4539 VSS.n3051 0.04025
R14099 VSS.n4543 VSS.n3051 0.04025
R14100 VSS.n4544 VSS.n4543 0.04025
R14101 VSS.n4545 VSS.n4544 0.04025
R14102 VSS.n4545 VSS.n3049 0.04025
R14103 VSS.n4549 VSS.n3049 0.04025
R14104 VSS.n4550 VSS.n4549 0.04025
R14105 VSS.n4551 VSS.n4550 0.04025
R14106 VSS.n4551 VSS.n3047 0.04025
R14107 VSS.n4555 VSS.n3047 0.04025
R14108 VSS.n4556 VSS.n4555 0.04025
R14109 VSS.n4557 VSS.n4556 0.04025
R14110 VSS.n4557 VSS.n3045 0.04025
R14111 VSS.n4561 VSS.n3045 0.04025
R14112 VSS.n4562 VSS.n4561 0.04025
R14113 VSS.n4563 VSS.n4562 0.04025
R14114 VSS.n4563 VSS.n3043 0.04025
R14115 VSS.n4567 VSS.n3043 0.04025
R14116 VSS.n4568 VSS.n4567 0.04025
R14117 VSS.n4569 VSS.n4568 0.04025
R14118 VSS.n4569 VSS.n3041 0.04025
R14119 VSS.n4573 VSS.n3041 0.04025
R14120 VSS.n4574 VSS.n4573 0.04025
R14121 VSS.n4575 VSS.n4574 0.04025
R14122 VSS.n4575 VSS.n3039 0.04025
R14123 VSS.n4579 VSS.n3039 0.04025
R14124 VSS.n4580 VSS.n4579 0.04025
R14125 VSS.n4581 VSS.n4580 0.04025
R14126 VSS.n4581 VSS.n3037 0.04025
R14127 VSS.n4585 VSS.n3037 0.04025
R14128 VSS.n4586 VSS.n4585 0.04025
R14129 VSS.n4587 VSS.n4586 0.04025
R14130 VSS.n4587 VSS.n3035 0.04025
R14131 VSS.n4591 VSS.n3035 0.04025
R14132 VSS.n4592 VSS.n4591 0.04025
R14133 VSS.n4593 VSS.n4592 0.04025
R14134 VSS.n4593 VSS.n3033 0.04025
R14135 VSS.n4597 VSS.n3033 0.04025
R14136 VSS.n4598 VSS.n4597 0.04025
R14137 VSS.n4599 VSS.n4598 0.04025
R14138 VSS.n4599 VSS.n3031 0.04025
R14139 VSS.n4603 VSS.n3031 0.04025
R14140 VSS.n4604 VSS.n4603 0.04025
R14141 VSS.n4605 VSS.n4604 0.04025
R14142 VSS.n4605 VSS.n3029 0.04025
R14143 VSS.n4609 VSS.n3029 0.04025
R14144 VSS.n4610 VSS.n4609 0.04025
R14145 VSS.n4611 VSS.n4610 0.04025
R14146 VSS.n4611 VSS.n3027 0.04025
R14147 VSS.n4615 VSS.n3027 0.04025
R14148 VSS.n4616 VSS.n4615 0.04025
R14149 VSS.n4617 VSS.n4616 0.04025
R14150 VSS.n4617 VSS.n3025 0.04025
R14151 VSS.n4621 VSS.n3025 0.04025
R14152 VSS.n4622 VSS.n4621 0.04025
R14153 VSS.n4623 VSS.n4622 0.04025
R14154 VSS.n4623 VSS.n3023 0.04025
R14155 VSS.n4627 VSS.n3023 0.04025
R14156 VSS.n4628 VSS.n4627 0.04025
R14157 VSS.n4629 VSS.n4628 0.04025
R14158 VSS.n4629 VSS.n3021 0.04025
R14159 VSS.n4633 VSS.n3021 0.04025
R14160 VSS.n4634 VSS.n4633 0.04025
R14161 VSS.n4635 VSS.n4634 0.04025
R14162 VSS.n4635 VSS.n3019 0.04025
R14163 VSS.n4639 VSS.n3019 0.04025
R14164 VSS.n4640 VSS.n4639 0.04025
R14165 VSS.n4641 VSS.n4640 0.04025
R14166 VSS.n4641 VSS.n3017 0.04025
R14167 VSS.n4645 VSS.n3017 0.04025
R14168 VSS.n4646 VSS.n4645 0.04025
R14169 VSS.n4647 VSS.n4646 0.04025
R14170 VSS.n4647 VSS.n3015 0.04025
R14171 VSS.n4651 VSS.n3015 0.04025
R14172 VSS.n4652 VSS.n4651 0.04025
R14173 VSS.n4653 VSS.n4652 0.04025
R14174 VSS.n4653 VSS.n3013 0.04025
R14175 VSS.n4657 VSS.n3013 0.04025
R14176 VSS.n4658 VSS.n4657 0.04025
R14177 VSS.n4659 VSS.n4658 0.04025
R14178 VSS.n4659 VSS.n3011 0.04025
R14179 VSS.n4663 VSS.n3011 0.04025
R14180 VSS.n4664 VSS.n4663 0.04025
R14181 VSS.n4665 VSS.n4664 0.04025
R14182 VSS.n4665 VSS.n3009 0.04025
R14183 VSS.n4669 VSS.n3009 0.04025
R14184 VSS.n4670 VSS.n4669 0.04025
R14185 VSS.n4671 VSS.n4670 0.04025
R14186 VSS.n4671 VSS.n3007 0.04025
R14187 VSS.n4675 VSS.n3007 0.04025
R14188 VSS.n4676 VSS.n4675 0.04025
R14189 VSS.n4677 VSS.n4676 0.04025
R14190 VSS.n4677 VSS.n3005 0.04025
R14191 VSS.n4681 VSS.n3005 0.04025
R14192 VSS.n4682 VSS.n4681 0.04025
R14193 VSS.n4683 VSS.n4682 0.04025
R14194 VSS.n4683 VSS.n3003 0.04025
R14195 VSS.n4687 VSS.n3003 0.04025
R14196 VSS.n4688 VSS.n4687 0.04025
R14197 VSS.n4689 VSS.n4688 0.04025
R14198 VSS.n4689 VSS.n3001 0.04025
R14199 VSS.n4693 VSS.n3001 0.04025
R14200 VSS.n4694 VSS.n4693 0.04025
R14201 VSS.n4695 VSS.n4694 0.04025
R14202 VSS.n4695 VSS.n2999 0.04025
R14203 VSS.n4699 VSS.n2999 0.04025
R14204 VSS.n4700 VSS.n4699 0.04025
R14205 VSS.n4701 VSS.n4700 0.04025
R14206 VSS.n4701 VSS.n2997 0.04025
R14207 VSS.n4705 VSS.n2997 0.04025
R14208 VSS.n4706 VSS.n4705 0.04025
R14209 VSS.n4707 VSS.n4706 0.04025
R14210 VSS.n4707 VSS.n2995 0.04025
R14211 VSS.n4711 VSS.n2995 0.04025
R14212 VSS.n4712 VSS.n4711 0.04025
R14213 VSS.n4713 VSS.n4712 0.04025
R14214 VSS.n4713 VSS.n2993 0.04025
R14215 VSS.n4717 VSS.n2993 0.04025
R14216 VSS.n4718 VSS.n4717 0.04025
R14217 VSS.n4719 VSS.n4718 0.04025
R14218 VSS.n4719 VSS.n2991 0.04025
R14219 VSS.n4723 VSS.n2991 0.04025
R14220 VSS.n4724 VSS.n4723 0.04025
R14221 VSS.n4725 VSS.n4724 0.04025
R14222 VSS.n4725 VSS.n2989 0.04025
R14223 VSS.n4729 VSS.n2989 0.04025
R14224 VSS.n4730 VSS.n4729 0.04025
R14225 VSS.n4731 VSS.n4730 0.04025
R14226 VSS.n4731 VSS.n2987 0.04025
R14227 VSS.n4735 VSS.n2987 0.04025
R14228 VSS.n4736 VSS.n4735 0.04025
R14229 VSS.n4737 VSS.n4736 0.04025
R14230 VSS.n4737 VSS.n2985 0.04025
R14231 VSS.n4741 VSS.n2985 0.04025
R14232 VSS.n4742 VSS.n4741 0.04025
R14233 VSS.n4743 VSS.n4742 0.04025
R14234 VSS.n4743 VSS.n2983 0.04025
R14235 VSS.n4747 VSS.n2983 0.04025
R14236 VSS.n4748 VSS.n4747 0.04025
R14237 VSS.n4749 VSS.n4748 0.04025
R14238 VSS.n4749 VSS.n2981 0.04025
R14239 VSS.n4753 VSS.n2981 0.04025
R14240 VSS.n4754 VSS.n4753 0.04025
R14241 VSS.n4755 VSS.n4754 0.04025
R14242 VSS.n4755 VSS.n2979 0.04025
R14243 VSS.n4759 VSS.n2979 0.04025
R14244 VSS.n4760 VSS.n4759 0.04025
R14245 VSS.n4761 VSS.n4760 0.04025
R14246 VSS.n4761 VSS.n2977 0.04025
R14247 VSS.n4765 VSS.n2977 0.04025
R14248 VSS.n4766 VSS.n4765 0.04025
R14249 VSS.n4767 VSS.n4766 0.04025
R14250 VSS.n4767 VSS.n2975 0.04025
R14251 VSS.n4771 VSS.n2975 0.04025
R14252 VSS.n4772 VSS.n4771 0.04025
R14253 VSS.n4773 VSS.n4772 0.04025
R14254 VSS.n4773 VSS.n2973 0.04025
R14255 VSS.n4777 VSS.n2973 0.04025
R14256 VSS.n4778 VSS.n4777 0.04025
R14257 VSS.n4779 VSS.n4778 0.04025
R14258 VSS.n4779 VSS.n2971 0.04025
R14259 VSS.n4783 VSS.n2971 0.04025
R14260 VSS.n4784 VSS.n4783 0.04025
R14261 VSS.n4785 VSS.n4784 0.04025
R14262 VSS.n4785 VSS.n2969 0.04025
R14263 VSS.n4789 VSS.n2969 0.04025
R14264 VSS.n4790 VSS.n4789 0.04025
R14265 VSS.n4791 VSS.n4790 0.04025
R14266 VSS.n4791 VSS.n2967 0.04025
R14267 VSS.n4795 VSS.n2967 0.04025
R14268 VSS.n4796 VSS.n4795 0.04025
R14269 VSS.n4797 VSS.n4796 0.04025
R14270 VSS.n4797 VSS.n2965 0.04025
R14271 VSS.n4801 VSS.n2965 0.04025
R14272 VSS.n4802 VSS.n4801 0.04025
R14273 VSS.n4806 VSS.n4802 0.04025
R14274 VSS.n4806 VSS.n2963 0.04025
R14275 VSS.n4810 VSS.n2963 0.04025
R14276 VSS.n4811 VSS.n4810 0.04025
R14277 VSS.n4812 VSS.n4811 0.04025
R14278 VSS.n4812 VSS.n2961 0.04025
R14279 VSS.n4816 VSS.n2961 0.04025
R14280 VSS.n4817 VSS.n4816 0.04025
R14281 VSS.n4818 VSS.n4817 0.04025
R14282 VSS.n4818 VSS.n2959 0.04025
R14283 VSS.n4822 VSS.n2959 0.04025
R14284 VSS.n4823 VSS.n4822 0.04025
R14285 VSS.n4824 VSS.n4823 0.04025
R14286 VSS.n4824 VSS.n2957 0.04025
R14287 VSS.n4828 VSS.n2957 0.04025
R14288 VSS.n4829 VSS.n4828 0.04025
R14289 VSS.n4830 VSS.n4829 0.04025
R14290 VSS.n4830 VSS.n2955 0.04025
R14291 VSS.n4834 VSS.n2955 0.04025
R14292 VSS.n4835 VSS.n4834 0.04025
R14293 VSS.n4836 VSS.n4835 0.04025
R14294 VSS.n4836 VSS.n2953 0.04025
R14295 VSS.n4840 VSS.n2953 0.04025
R14296 VSS.n4841 VSS.n4840 0.04025
R14297 VSS.n4842 VSS.n4841 0.04025
R14298 VSS.n4842 VSS.n2951 0.04025
R14299 VSS.n4846 VSS.n2951 0.04025
R14300 VSS.n4847 VSS.n4846 0.04025
R14301 VSS.n4848 VSS.n4847 0.04025
R14302 VSS.n4848 VSS.n2949 0.04025
R14303 VSS.n4852 VSS.n2949 0.04025
R14304 VSS.n4853 VSS.n4852 0.04025
R14305 VSS.n4854 VSS.n4853 0.04025
R14306 VSS.n4854 VSS.n2947 0.04025
R14307 VSS.n4858 VSS.n2947 0.04025
R14308 VSS.n4859 VSS.n4858 0.04025
R14309 VSS.n4860 VSS.n4859 0.04025
R14310 VSS.n4860 VSS.n2945 0.04025
R14311 VSS.n4864 VSS.n2945 0.04025
R14312 VSS.n4865 VSS.n4864 0.04025
R14313 VSS.n4866 VSS.n4865 0.04025
R14314 VSS.n4866 VSS.n2943 0.04025
R14315 VSS.n4870 VSS.n2943 0.04025
R14316 VSS.n4871 VSS.n4870 0.04025
R14317 VSS.n4872 VSS.n4871 0.04025
R14318 VSS.n4872 VSS.n2941 0.04025
R14319 VSS.n4876 VSS.n2941 0.04025
R14320 VSS.n4877 VSS.n4876 0.04025
R14321 VSS.n4878 VSS.n4877 0.04025
R14322 VSS.n4878 VSS.n2939 0.04025
R14323 VSS.n4882 VSS.n2939 0.04025
R14324 VSS.n4883 VSS.n4882 0.04025
R14325 VSS.n4884 VSS.n4883 0.04025
R14326 VSS.n4884 VSS.n2937 0.04025
R14327 VSS.n4888 VSS.n2937 0.04025
R14328 VSS.n4889 VSS.n4888 0.04025
R14329 VSS.n4890 VSS.n4889 0.04025
R14330 VSS.n4890 VSS.n2935 0.04025
R14331 VSS.n4894 VSS.n2935 0.04025
R14332 VSS.n4895 VSS.n4894 0.04025
R14333 VSS.n4896 VSS.n4895 0.04025
R14334 VSS.n4896 VSS.n2933 0.04025
R14335 VSS.n4900 VSS.n2933 0.04025
R14336 VSS.n4901 VSS.n4900 0.04025
R14337 VSS.n4902 VSS.n4901 0.04025
R14338 VSS.n4902 VSS.n2931 0.04025
R14339 VSS.n4906 VSS.n2931 0.04025
R14340 VSS.n4907 VSS.n4906 0.04025
R14341 VSS.n4908 VSS.n4907 0.04025
R14342 VSS.n4908 VSS.n2929 0.04025
R14343 VSS.n4912 VSS.n2929 0.04025
R14344 VSS.n4913 VSS.n4912 0.04025
R14345 VSS.n4914 VSS.n4913 0.04025
R14346 VSS.n4914 VSS.n2927 0.04025
R14347 VSS.n4918 VSS.n2927 0.04025
R14348 VSS.n4919 VSS.n4918 0.04025
R14349 VSS.n4920 VSS.n4919 0.04025
R14350 VSS.n4920 VSS.n2925 0.04025
R14351 VSS.n4924 VSS.n2925 0.04025
R14352 VSS.n4925 VSS.n4924 0.04025
R14353 VSS.n4926 VSS.n4925 0.04025
R14354 VSS.n4926 VSS.n2923 0.04025
R14355 VSS.n4930 VSS.n2923 0.04025
R14356 VSS.n4931 VSS.n4930 0.04025
R14357 VSS.n4932 VSS.n4931 0.04025
R14358 VSS.n4932 VSS.n2921 0.04025
R14359 VSS.n4936 VSS.n2921 0.04025
R14360 VSS.n4937 VSS.n4936 0.04025
R14361 VSS.n4938 VSS.n4937 0.04025
R14362 VSS.n4938 VSS.n2919 0.04025
R14363 VSS.n4942 VSS.n2919 0.04025
R14364 VSS.n4943 VSS.n4942 0.04025
R14365 VSS.n4944 VSS.n4943 0.04025
R14366 VSS.n4944 VSS.n2917 0.04025
R14367 VSS.n4948 VSS.n2917 0.04025
R14368 VSS.n4949 VSS.n4948 0.04025
R14369 VSS.n4950 VSS.n4949 0.04025
R14370 VSS.n4950 VSS.n2915 0.04025
R14371 VSS.n4954 VSS.n2915 0.04025
R14372 VSS.n4955 VSS.n4954 0.04025
R14373 VSS.n4956 VSS.n4955 0.04025
R14374 VSS.n4956 VSS.n2913 0.04025
R14375 VSS.n4960 VSS.n2913 0.04025
R14376 VSS.n4961 VSS.n4960 0.04025
R14377 VSS.n4962 VSS.n4961 0.04025
R14378 VSS.n4962 VSS.n2911 0.04025
R14379 VSS.n4966 VSS.n2911 0.04025
R14380 VSS.n4967 VSS.n4966 0.04025
R14381 VSS.n4968 VSS.n4967 0.04025
R14382 VSS.n4968 VSS.n2909 0.04025
R14383 VSS.n4972 VSS.n2909 0.04025
R14384 VSS.n4973 VSS.n4972 0.04025
R14385 VSS.n4974 VSS.n4973 0.04025
R14386 VSS.n4974 VSS.n2907 0.04025
R14387 VSS.n4978 VSS.n2907 0.04025
R14388 VSS.n4979 VSS.n4978 0.04025
R14389 VSS.n4980 VSS.n4979 0.04025
R14390 VSS.n4980 VSS.n2905 0.04025
R14391 VSS.n4984 VSS.n2905 0.04025
R14392 VSS.n4985 VSS.n4984 0.04025
R14393 VSS.n4986 VSS.n4985 0.04025
R14394 VSS.n4986 VSS.n2903 0.04025
R14395 VSS.n4990 VSS.n2903 0.04025
R14396 VSS.n4991 VSS.n4990 0.04025
R14397 VSS.n4992 VSS.n4991 0.04025
R14398 VSS.n4992 VSS.n2901 0.04025
R14399 VSS.n4996 VSS.n2901 0.04025
R14400 VSS.n4997 VSS.n4996 0.04025
R14401 VSS.n4998 VSS.n4997 0.04025
R14402 VSS.n4998 VSS.n2899 0.04025
R14403 VSS.n5002 VSS.n2899 0.04025
R14404 VSS.n5003 VSS.n5002 0.04025
R14405 VSS.n5004 VSS.n5003 0.04025
R14406 VSS.n5004 VSS.n2897 0.04025
R14407 VSS.n5008 VSS.n2897 0.04025
R14408 VSS.n5009 VSS.n5008 0.04025
R14409 VSS.n5010 VSS.n5009 0.04025
R14410 VSS.n5010 VSS.n2895 0.04025
R14411 VSS.n5014 VSS.n2895 0.04025
R14412 VSS.n5015 VSS.n5014 0.04025
R14413 VSS.n5016 VSS.n5015 0.04025
R14414 VSS.n5016 VSS.n2893 0.04025
R14415 VSS.n5020 VSS.n2893 0.04025
R14416 VSS.n5021 VSS.n5020 0.04025
R14417 VSS.n5022 VSS.n5021 0.04025
R14418 VSS.n5022 VSS.n2891 0.04025
R14419 VSS.n5026 VSS.n2891 0.04025
R14420 VSS.n5027 VSS.n5026 0.04025
R14421 VSS.n5028 VSS.n5027 0.04025
R14422 VSS.n5028 VSS.n2889 0.04025
R14423 VSS.n5032 VSS.n2889 0.04025
R14424 VSS.n5033 VSS.n5032 0.04025
R14425 VSS.n5034 VSS.n5033 0.04025
R14426 VSS.n5034 VSS.n2887 0.04025
R14427 VSS.n5038 VSS.n2887 0.04025
R14428 VSS.n5039 VSS.n5038 0.04025
R14429 VSS.n5040 VSS.n5039 0.04025
R14430 VSS.n5040 VSS.n2885 0.04025
R14431 VSS.n5044 VSS.n2885 0.04025
R14432 VSS.n5045 VSS.n5044 0.04025
R14433 VSS.n5046 VSS.n5045 0.04025
R14434 VSS.n5046 VSS.n2883 0.04025
R14435 VSS.n5050 VSS.n2883 0.04025
R14436 VSS.n5051 VSS.n5050 0.04025
R14437 VSS.n5052 VSS.n5051 0.04025
R14438 VSS.n5052 VSS.n2881 0.04025
R14439 VSS.n5056 VSS.n2881 0.04025
R14440 VSS.n5057 VSS.n5056 0.04025
R14441 VSS.n5058 VSS.n5057 0.04025
R14442 VSS.n5058 VSS.n2879 0.04025
R14443 VSS.n5062 VSS.n2879 0.04025
R14444 VSS.n5063 VSS.n5062 0.04025
R14445 VSS.n5064 VSS.n5063 0.04025
R14446 VSS.n5064 VSS.n2877 0.04025
R14447 VSS.n5068 VSS.n2877 0.04025
R14448 VSS.n5069 VSS.n5068 0.04025
R14449 VSS.n5070 VSS.n5069 0.04025
R14450 VSS.n5070 VSS.n2875 0.04025
R14451 VSS.n5074 VSS.n2875 0.04025
R14452 VSS.n5075 VSS.n5074 0.04025
R14453 VSS.n5076 VSS.n5075 0.04025
R14454 VSS.n5076 VSS.n2873 0.04025
R14455 VSS.n5080 VSS.n2873 0.04025
R14456 VSS.n5081 VSS.n5080 0.04025
R14457 VSS.n5082 VSS.n5081 0.04025
R14458 VSS.n5082 VSS.n2871 0.04025
R14459 VSS.n5086 VSS.n2871 0.04025
R14460 VSS.n5087 VSS.n5086 0.04025
R14461 VSS.n5088 VSS.n5087 0.04025
R14462 VSS.n5088 VSS.n2869 0.04025
R14463 VSS.n5092 VSS.n2869 0.04025
R14464 VSS.n5093 VSS.n5092 0.04025
R14465 VSS.n5094 VSS.n5093 0.04025
R14466 VSS.n5094 VSS.n2867 0.04025
R14467 VSS.n5098 VSS.n2867 0.04025
R14468 VSS.n5099 VSS.n5098 0.04025
R14469 VSS.n5100 VSS.n5099 0.04025
R14470 VSS.n5100 VSS.n2865 0.04025
R14471 VSS.n5104 VSS.n2865 0.04025
R14472 VSS.n5105 VSS.n5104 0.04025
R14473 VSS.n5106 VSS.n5105 0.04025
R14474 VSS.n5106 VSS.n2863 0.04025
R14475 VSS.n5110 VSS.n2863 0.04025
R14476 VSS.n5111 VSS.n5110 0.04025
R14477 VSS.n5112 VSS.n5111 0.04025
R14478 VSS.n5112 VSS.n2861 0.04025
R14479 VSS.n5116 VSS.n2861 0.04025
R14480 VSS.n5117 VSS.n5116 0.04025
R14481 VSS.n5118 VSS.n5117 0.04025
R14482 VSS.n5118 VSS.n2859 0.04025
R14483 VSS.n5122 VSS.n2859 0.04025
R14484 VSS.n5123 VSS.n5122 0.04025
R14485 VSS.n5124 VSS.n5123 0.04025
R14486 VSS.n5124 VSS.n2857 0.04025
R14487 VSS.n5128 VSS.n2857 0.04025
R14488 VSS.n5129 VSS.n5128 0.04025
R14489 VSS.n5130 VSS.n5129 0.04025
R14490 VSS.n5130 VSS.n2855 0.04025
R14491 VSS.n5134 VSS.n2855 0.04025
R14492 VSS.n5135 VSS.n5134 0.04025
R14493 VSS.n5136 VSS.n5135 0.04025
R14494 VSS.n5136 VSS.n2853 0.04025
R14495 VSS.n5140 VSS.n2853 0.04025
R14496 VSS.n5141 VSS.n5140 0.04025
R14497 VSS.n5142 VSS.n5141 0.04025
R14498 VSS.n5142 VSS.n2851 0.04025
R14499 VSS.n5146 VSS.n2851 0.04025
R14500 VSS.n5147 VSS.n5146 0.04025
R14501 VSS.n5148 VSS.n5147 0.04025
R14502 VSS.n5148 VSS.n2849 0.04025
R14503 VSS.n5152 VSS.n2849 0.04025
R14504 VSS.n5153 VSS.n5152 0.04025
R14505 VSS.n5154 VSS.n5153 0.04025
R14506 VSS.n5154 VSS.n2847 0.04025
R14507 VSS.n5158 VSS.n2847 0.04025
R14508 VSS.n5159 VSS.n5158 0.04025
R14509 VSS.n5160 VSS.n5159 0.04025
R14510 VSS.n5160 VSS.n2845 0.04025
R14511 VSS.n5164 VSS.n2845 0.04025
R14512 VSS.n5165 VSS.n5164 0.04025
R14513 VSS.n5166 VSS.n5165 0.04025
R14514 VSS.n5166 VSS.n2843 0.04025
R14515 VSS.n5170 VSS.n2843 0.04025
R14516 VSS.n5171 VSS.n5170 0.04025
R14517 VSS.n5172 VSS.n5171 0.04025
R14518 VSS.n5172 VSS.n2841 0.04025
R14519 VSS.n5176 VSS.n2841 0.04025
R14520 VSS.n5177 VSS.n5176 0.04025
R14521 VSS.n5178 VSS.n5177 0.04025
R14522 VSS.n5178 VSS.n2839 0.04025
R14523 VSS.n5182 VSS.n2839 0.04025
R14524 VSS.n5183 VSS.n5182 0.04025
R14525 VSS.n5184 VSS.n5183 0.04025
R14526 VSS.n5184 VSS.n2837 0.04025
R14527 VSS.n5188 VSS.n2837 0.04025
R14528 VSS.n5189 VSS.n5188 0.04025
R14529 VSS.n5190 VSS.n5189 0.04025
R14530 VSS.n5190 VSS.n2835 0.04025
R14531 VSS.n5194 VSS.n2835 0.04025
R14532 VSS.n5195 VSS.n5194 0.04025
R14533 VSS.n5196 VSS.n5195 0.04025
R14534 VSS.n5196 VSS.n2833 0.04025
R14535 VSS.n5200 VSS.n2833 0.04025
R14536 VSS.n5201 VSS.n5200 0.04025
R14537 VSS.n5202 VSS.n5201 0.04025
R14538 VSS.n5202 VSS.n2831 0.04025
R14539 VSS.n5206 VSS.n2831 0.04025
R14540 VSS.n5207 VSS.n5206 0.04025
R14541 VSS.n5208 VSS.n5207 0.04025
R14542 VSS.n5208 VSS.n2829 0.04025
R14543 VSS.n5212 VSS.n2829 0.04025
R14544 VSS.n5213 VSS.n5212 0.04025
R14545 VSS.n5214 VSS.n5213 0.04025
R14546 VSS.n5214 VSS.n2827 0.04025
R14547 VSS.n5218 VSS.n2827 0.04025
R14548 VSS.n5219 VSS.n5218 0.04025
R14549 VSS.n5220 VSS.n5219 0.04025
R14550 VSS.n5220 VSS.n2825 0.04025
R14551 VSS.n5224 VSS.n2825 0.04025
R14552 VSS.n5225 VSS.n5224 0.04025
R14553 VSS.n5226 VSS.n5225 0.04025
R14554 VSS.n5226 VSS.n2823 0.04025
R14555 VSS.n5230 VSS.n2823 0.04025
R14556 VSS.n5231 VSS.n5230 0.04025
R14557 VSS.n5232 VSS.n5231 0.04025
R14558 VSS.n5232 VSS.n2821 0.04025
R14559 VSS.n5236 VSS.n2821 0.04025
R14560 VSS.n5237 VSS.n5236 0.04025
R14561 VSS.n5238 VSS.n5237 0.04025
R14562 VSS.n5238 VSS.n2819 0.04025
R14563 VSS.n5242 VSS.n2819 0.04025
R14564 VSS.n5243 VSS.n5242 0.04025
R14565 VSS.n5244 VSS.n5243 0.04025
R14566 VSS.n5244 VSS.n2817 0.04025
R14567 VSS.n5248 VSS.n2817 0.04025
R14568 VSS.n5249 VSS.n5248 0.04025
R14569 VSS.n5250 VSS.n5249 0.04025
R14570 VSS.n5250 VSS.n2815 0.04025
R14571 VSS.n5254 VSS.n2815 0.04025
R14572 VSS.n5255 VSS.n5254 0.04025
R14573 VSS.n5256 VSS.n5255 0.04025
R14574 VSS.n5256 VSS.n2813 0.04025
R14575 VSS.n5260 VSS.n2813 0.04025
R14576 VSS.n5261 VSS.n5260 0.04025
R14577 VSS.n5262 VSS.n5261 0.04025
R14578 VSS.n5262 VSS.n2811 0.04025
R14579 VSS.n5266 VSS.n2811 0.04025
R14580 VSS.n5267 VSS.n5266 0.04025
R14581 VSS.n5268 VSS.n5267 0.04025
R14582 VSS.n5268 VSS.n2809 0.04025
R14583 VSS.n5272 VSS.n2809 0.04025
R14584 VSS.n5273 VSS.n5272 0.04025
R14585 VSS.n5274 VSS.n5273 0.04025
R14586 VSS.n5274 VSS.n2807 0.04025
R14587 VSS.n5278 VSS.n2807 0.04025
R14588 VSS.n5279 VSS.n5278 0.04025
R14589 VSS.n5280 VSS.n5279 0.04025
R14590 VSS.n5280 VSS.n2805 0.04025
R14591 VSS.n5284 VSS.n2805 0.04025
R14592 VSS.n5285 VSS.n5284 0.04025
R14593 VSS.n5286 VSS.n5285 0.04025
R14594 VSS.n5286 VSS.n2803 0.04025
R14595 VSS.n5290 VSS.n2803 0.04025
R14596 VSS.n5291 VSS.n5290 0.04025
R14597 VSS.n5292 VSS.n5291 0.04025
R14598 VSS.n5292 VSS.n2801 0.04025
R14599 VSS.n5296 VSS.n2801 0.04025
R14600 VSS.n5297 VSS.n5296 0.04025
R14601 VSS.n5298 VSS.n5297 0.04025
R14602 VSS.n5298 VSS.n2799 0.04025
R14603 VSS.n5302 VSS.n2799 0.04025
R14604 VSS.n5303 VSS.n5302 0.04025
R14605 VSS.n5304 VSS.n5303 0.04025
R14606 VSS.n5304 VSS.n2797 0.04025
R14607 VSS.n5308 VSS.n2797 0.04025
R14608 VSS.n5309 VSS.n5308 0.04025
R14609 VSS.n5310 VSS.n5309 0.04025
R14610 VSS.n5310 VSS.n2795 0.04025
R14611 VSS.n5314 VSS.n2795 0.04025
R14612 VSS.n5315 VSS.n5314 0.04025
R14613 VSS.n5316 VSS.n5315 0.04025
R14614 VSS.n5316 VSS.n2793 0.04025
R14615 VSS.n5320 VSS.n2793 0.04025
R14616 VSS.n5321 VSS.n5320 0.04025
R14617 VSS.n5322 VSS.n5321 0.04025
R14618 VSS.n5322 VSS.n2791 0.04025
R14619 VSS.n5326 VSS.n2791 0.04025
R14620 VSS.n5327 VSS.n5326 0.04025
R14621 VSS.n5328 VSS.n5327 0.04025
R14622 VSS.n5328 VSS.n2789 0.04025
R14623 VSS.n5332 VSS.n2789 0.04025
R14624 VSS.n5333 VSS.n5332 0.04025
R14625 VSS.n5334 VSS.n5333 0.04025
R14626 VSS.n5334 VSS.n2787 0.04025
R14627 VSS.n5338 VSS.n2787 0.04025
R14628 VSS.n5339 VSS.n5338 0.04025
R14629 VSS.n5340 VSS.n5339 0.04025
R14630 VSS.n5340 VSS.n2785 0.04025
R14631 VSS.n5344 VSS.n2785 0.04025
R14632 VSS.n5345 VSS.n5344 0.04025
R14633 VSS.n5346 VSS.n5345 0.04025
R14634 VSS.n5346 VSS.n2783 0.04025
R14635 VSS.n5350 VSS.n2783 0.04025
R14636 VSS.n5351 VSS.n5350 0.04025
R14637 VSS.n5352 VSS.n5351 0.04025
R14638 VSS.n5352 VSS.n2781 0.04025
R14639 VSS.n5356 VSS.n2781 0.04025
R14640 VSS.n5357 VSS.n5356 0.04025
R14641 VSS.n5358 VSS.n5357 0.04025
R14642 VSS.n5358 VSS.n2779 0.04025
R14643 VSS.n5362 VSS.n2779 0.04025
R14644 VSS.n5363 VSS.n5362 0.04025
R14645 VSS.n5364 VSS.n5363 0.04025
R14646 VSS.n5364 VSS.n2777 0.04025
R14647 VSS.n5368 VSS.n2777 0.04025
R14648 VSS.n5369 VSS.n5368 0.04025
R14649 VSS.n5370 VSS.n5369 0.04025
R14650 VSS.n5370 VSS.n2775 0.04025
R14651 VSS.n5374 VSS.n2775 0.04025
R14652 VSS.n5375 VSS.n5374 0.04025
R14653 VSS.n5376 VSS.n5375 0.04025
R14654 VSS.n5376 VSS.n2773 0.04025
R14655 VSS.n5380 VSS.n2773 0.04025
R14656 VSS.n5381 VSS.n5380 0.04025
R14657 VSS.n5382 VSS.n5381 0.04025
R14658 VSS.n5382 VSS.n2771 0.04025
R14659 VSS.n5386 VSS.n2771 0.04025
R14660 VSS.n5387 VSS.n5386 0.04025
R14661 VSS.n5388 VSS.n5387 0.04025
R14662 VSS.n5388 VSS.n2769 0.04025
R14663 VSS.n5392 VSS.n2769 0.04025
R14664 VSS.n5393 VSS.n5392 0.04025
R14665 VSS.n5394 VSS.n5393 0.04025
R14666 VSS.n5394 VSS.n2767 0.04025
R14667 VSS.n5398 VSS.n2767 0.04025
R14668 VSS.n5399 VSS.n5398 0.04025
R14669 VSS.n5400 VSS.n5399 0.04025
R14670 VSS.n5400 VSS.n2765 0.04025
R14671 VSS.n5404 VSS.n2765 0.04025
R14672 VSS.n5405 VSS.n5404 0.04025
R14673 VSS.n5406 VSS.n5405 0.04025
R14674 VSS.n5406 VSS.n2763 0.04025
R14675 VSS.n5410 VSS.n2763 0.04025
R14676 VSS.n5411 VSS.n5410 0.04025
R14677 VSS.n5412 VSS.n5411 0.04025
R14678 VSS.n5412 VSS.n2761 0.04025
R14679 VSS.n5416 VSS.n2761 0.04025
R14680 VSS.n5417 VSS.n5416 0.04025
R14681 VSS.n5418 VSS.n5417 0.04025
R14682 VSS.n5418 VSS.n2759 0.04025
R14683 VSS.n5422 VSS.n2759 0.04025
R14684 VSS.n5423 VSS.n5422 0.04025
R14685 VSS.n5424 VSS.n5423 0.04025
R14686 VSS.n5424 VSS.n2757 0.04025
R14687 VSS.n5428 VSS.n2757 0.04025
R14688 VSS.n5429 VSS.n5428 0.04025
R14689 VSS.n5430 VSS.n5429 0.04025
R14690 VSS.n5430 VSS.n2755 0.04025
R14691 VSS.n5434 VSS.n2755 0.04025
R14692 VSS.n5435 VSS.n5434 0.04025
R14693 VSS.n5436 VSS.n5435 0.04025
R14694 VSS.n5436 VSS.n2753 0.04025
R14695 VSS.n5440 VSS.n2753 0.04025
R14696 VSS.n5441 VSS.n5440 0.04025
R14697 VSS.n5442 VSS.n5441 0.04025
R14698 VSS.n5442 VSS.n2751 0.04025
R14699 VSS.n5446 VSS.n2751 0.04025
R14700 VSS.n5447 VSS.n5446 0.04025
R14701 VSS.n5448 VSS.n5447 0.04025
R14702 VSS.n5448 VSS.n2749 0.04025
R14703 VSS.n5452 VSS.n2749 0.04025
R14704 VSS.n5453 VSS.n5452 0.04025
R14705 VSS.n5454 VSS.n5453 0.04025
R14706 VSS.n5454 VSS.n2747 0.04025
R14707 VSS.n5458 VSS.n2747 0.04025
R14708 VSS.n5459 VSS.n5458 0.04025
R14709 VSS.n5460 VSS.n5459 0.04025
R14710 VSS.n5460 VSS.n2745 0.04025
R14711 VSS.n5464 VSS.n2745 0.04025
R14712 VSS.n5465 VSS.n5464 0.04025
R14713 VSS.n5466 VSS.n5465 0.04025
R14714 VSS.n5466 VSS.n2743 0.04025
R14715 VSS.n5471 VSS.n5470 0.04025
R14716 VSS.n5472 VSS.n5471 0.04025
R14717 VSS.n5472 VSS.n2741 0.04025
R14718 VSS.n5476 VSS.n2741 0.04025
R14719 VSS.n5477 VSS.n5476 0.04025
R14720 VSS.n5478 VSS.n5477 0.04025
R14721 VSS.n5478 VSS.n2739 0.04025
R14722 VSS.n5482 VSS.n2739 0.04025
R14723 VSS.n5483 VSS.n5482 0.04025
R14724 VSS.n5484 VSS.n5483 0.04025
R14725 VSS.n5484 VSS.n2737 0.04025
R14726 VSS.n5488 VSS.n2737 0.04025
R14727 VSS.n5489 VSS.n5488 0.04025
R14728 VSS.n5490 VSS.n5489 0.04025
R14729 VSS.n5490 VSS.n2735 0.04025
R14730 VSS.n5494 VSS.n2735 0.04025
R14731 VSS.n5495 VSS.n5494 0.04025
R14732 VSS.n5496 VSS.n5495 0.04025
R14733 VSS.n5496 VSS.n2733 0.04025
R14734 VSS.n5500 VSS.n2733 0.04025
R14735 VSS.n5501 VSS.n5500 0.04025
R14736 VSS.n5502 VSS.n5501 0.04025
R14737 VSS.n5502 VSS.n2731 0.04025
R14738 VSS.n5506 VSS.n2731 0.04025
R14739 VSS.n5507 VSS.n5506 0.04025
R14740 VSS.n5508 VSS.n5507 0.04025
R14741 VSS.n5508 VSS.n2729 0.04025
R14742 VSS.n5512 VSS.n2729 0.04025
R14743 VSS.n5513 VSS.n5512 0.04025
R14744 VSS.n5514 VSS.n5513 0.04025
R14745 VSS.n5514 VSS.n2727 0.04025
R14746 VSS.n5518 VSS.n2727 0.04025
R14747 VSS.n5519 VSS.n5518 0.04025
R14748 VSS.n5520 VSS.n5519 0.04025
R14749 VSS.n5520 VSS.n2725 0.04025
R14750 VSS.n5524 VSS.n2725 0.04025
R14751 VSS.n5525 VSS.n5524 0.04025
R14752 VSS.n5526 VSS.n5525 0.04025
R14753 VSS.n5526 VSS.n2723 0.04025
R14754 VSS.n5530 VSS.n2723 0.04025
R14755 VSS.n5531 VSS.n5530 0.04025
R14756 VSS.n5532 VSS.n5531 0.04025
R14757 VSS.n5532 VSS.n2721 0.04025
R14758 VSS.n5536 VSS.n2721 0.04025
R14759 VSS.n5537 VSS.n5536 0.04025
R14760 VSS.n5538 VSS.n5537 0.04025
R14761 VSS.n5538 VSS.n2719 0.04025
R14762 VSS.n5542 VSS.n2719 0.04025
R14763 VSS.n5543 VSS.n5542 0.04025
R14764 VSS.n5544 VSS.n5543 0.04025
R14765 VSS.n5544 VSS.n2717 0.04025
R14766 VSS.n5548 VSS.n2717 0.04025
R14767 VSS.n5549 VSS.n5548 0.04025
R14768 VSS.n5550 VSS.n5549 0.04025
R14769 VSS.n5550 VSS.n2715 0.04025
R14770 VSS.n5554 VSS.n2715 0.04025
R14771 VSS.n5555 VSS.n5554 0.04025
R14772 VSS.n5556 VSS.n5555 0.04025
R14773 VSS.n5556 VSS.n2713 0.04025
R14774 VSS.n5560 VSS.n2713 0.04025
R14775 VSS.n5561 VSS.n5560 0.04025
R14776 VSS.n5562 VSS.n5561 0.04025
R14777 VSS.n5562 VSS.n2711 0.04025
R14778 VSS.n5566 VSS.n2711 0.04025
R14779 VSS.n5567 VSS.n5566 0.04025
R14780 VSS.n5568 VSS.n5567 0.04025
R14781 VSS.n5568 VSS.n2709 0.04025
R14782 VSS.n5572 VSS.n2709 0.04025
R14783 VSS.n5573 VSS.n5572 0.04025
R14784 VSS.n5574 VSS.n5573 0.04025
R14785 VSS.n5574 VSS.n2707 0.04025
R14786 VSS.n5578 VSS.n2707 0.04025
R14787 VSS.n5579 VSS.n5578 0.04025
R14788 VSS.n5580 VSS.n5579 0.04025
R14789 VSS.n5580 VSS.n2705 0.04025
R14790 VSS.n5584 VSS.n2705 0.04025
R14791 VSS.n5585 VSS.n5584 0.04025
R14792 VSS.n5586 VSS.n5585 0.04025
R14793 VSS.n5586 VSS.n2703 0.04025
R14794 VSS.n5590 VSS.n2703 0.04025
R14795 VSS.n5591 VSS.n5590 0.04025
R14796 VSS.n5592 VSS.n5591 0.04025
R14797 VSS.n5592 VSS.n2701 0.04025
R14798 VSS.n5596 VSS.n2701 0.04025
R14799 VSS.n5597 VSS.n5596 0.04025
R14800 VSS.n5598 VSS.n5597 0.04025
R14801 VSS.n5598 VSS.n2699 0.04025
R14802 VSS.n5602 VSS.n2699 0.04025
R14803 VSS.n5603 VSS.n5602 0.04025
R14804 VSS.n5604 VSS.n5603 0.04025
R14805 VSS.n5604 VSS.n2697 0.04025
R14806 VSS.n5608 VSS.n2697 0.04025
R14807 VSS.n5609 VSS.n5608 0.04025
R14808 VSS.n5610 VSS.n5609 0.04025
R14809 VSS.n5610 VSS.n2695 0.04025
R14810 VSS.n5614 VSS.n2695 0.04025
R14811 VSS.n5615 VSS.n5614 0.04025
R14812 VSS.n5616 VSS.n5615 0.04025
R14813 VSS.n5616 VSS.n2693 0.04025
R14814 VSS.n5620 VSS.n2693 0.04025
R14815 VSS.n5621 VSS.n5620 0.04025
R14816 VSS.n5622 VSS.n5621 0.04025
R14817 VSS.n5622 VSS.n2691 0.04025
R14818 VSS.n5626 VSS.n2691 0.04025
R14819 VSS.n5627 VSS.n5626 0.04025
R14820 VSS.n5628 VSS.n5627 0.04025
R14821 VSS.n5628 VSS.n2689 0.04025
R14822 VSS.n5632 VSS.n2689 0.04025
R14823 VSS.n5633 VSS.n5632 0.04025
R14824 VSS.n5634 VSS.n5633 0.04025
R14825 VSS.n5634 VSS.n2687 0.04025
R14826 VSS.n5638 VSS.n2687 0.04025
R14827 VSS.n5639 VSS.n5638 0.04025
R14828 VSS.n5640 VSS.n5639 0.04025
R14829 VSS.n5640 VSS.n2685 0.04025
R14830 VSS.n5644 VSS.n2685 0.04025
R14831 VSS.n5645 VSS.n5644 0.04025
R14832 VSS.n5646 VSS.n5645 0.04025
R14833 VSS.n5646 VSS.n2683 0.04025
R14834 VSS.n5650 VSS.n2683 0.04025
R14835 VSS.n5651 VSS.n5650 0.04025
R14836 VSS.n5652 VSS.n5651 0.04025
R14837 VSS.n5652 VSS.n2681 0.04025
R14838 VSS.n5656 VSS.n2681 0.04025
R14839 VSS.n5657 VSS.n5656 0.04025
R14840 VSS.n5658 VSS.n5657 0.04025
R14841 VSS.n5658 VSS.n2679 0.04025
R14842 VSS.n5662 VSS.n2679 0.04025
R14843 VSS.n5663 VSS.n5662 0.04025
R14844 VSS.n5664 VSS.n5663 0.04025
R14845 VSS.n5664 VSS.n2677 0.04025
R14846 VSS.n5668 VSS.n2677 0.04025
R14847 VSS.n5669 VSS.n5668 0.04025
R14848 VSS.n5670 VSS.n5669 0.04025
R14849 VSS.n5670 VSS.n2675 0.04025
R14850 VSS.n5674 VSS.n2675 0.04025
R14851 VSS.n5675 VSS.n5674 0.04025
R14852 VSS.n5676 VSS.n5675 0.04025
R14853 VSS.n5676 VSS.n2673 0.04025
R14854 VSS.n5680 VSS.n2673 0.04025
R14855 VSS.n5681 VSS.n5680 0.04025
R14856 VSS.n5682 VSS.n5681 0.04025
R14857 VSS.n5682 VSS.n2671 0.04025
R14858 VSS.n5686 VSS.n2671 0.04025
R14859 VSS.n5687 VSS.n5686 0.04025
R14860 VSS.n5688 VSS.n5687 0.04025
R14861 VSS.n5688 VSS.n2669 0.04025
R14862 VSS.n5692 VSS.n2669 0.04025
R14863 VSS.n5693 VSS.n5692 0.04025
R14864 VSS.n5694 VSS.n5693 0.04025
R14865 VSS.n5694 VSS.n2667 0.04025
R14866 VSS.n5698 VSS.n2667 0.04025
R14867 VSS.n5699 VSS.n5698 0.04025
R14868 VSS.n5700 VSS.n5699 0.04025
R14869 VSS.n5700 VSS.n2665 0.04025
R14870 VSS.n5704 VSS.n2665 0.04025
R14871 VSS.n5705 VSS.n5704 0.04025
R14872 VSS.n5706 VSS.n5705 0.04025
R14873 VSS.n5706 VSS.n2663 0.04025
R14874 VSS.n5710 VSS.n2663 0.04025
R14875 VSS.n5711 VSS.n5710 0.04025
R14876 VSS.n5712 VSS.n5711 0.04025
R14877 VSS.n5712 VSS.n2661 0.04025
R14878 VSS.n5716 VSS.n2661 0.04025
R14879 VSS.n5717 VSS.n5716 0.04025
R14880 VSS.n5718 VSS.n5717 0.04025
R14881 VSS.n5718 VSS.n2659 0.04025
R14882 VSS.n5722 VSS.n2659 0.04025
R14883 VSS.n5723 VSS.n5722 0.04025
R14884 VSS.n5724 VSS.n5723 0.04025
R14885 VSS.n5724 VSS.n2657 0.04025
R14886 VSS.n5728 VSS.n2657 0.04025
R14887 VSS.n5729 VSS.n5728 0.04025
R14888 VSS.n5730 VSS.n5729 0.04025
R14889 VSS.n5730 VSS.n2655 0.04025
R14890 VSS.n5734 VSS.n2655 0.04025
R14891 VSS.n5735 VSS.n5734 0.04025
R14892 VSS.n5736 VSS.n5735 0.04025
R14893 VSS.n5736 VSS.n2653 0.04025
R14894 VSS.n5740 VSS.n2653 0.04025
R14895 VSS.n5741 VSS.n5740 0.04025
R14896 VSS.n5742 VSS.n5741 0.04025
R14897 VSS.n5742 VSS.n2651 0.04025
R14898 VSS.n5746 VSS.n2651 0.04025
R14899 VSS.n5747 VSS.n5746 0.04025
R14900 VSS.n5748 VSS.n5747 0.04025
R14901 VSS.n5748 VSS.n2649 0.04025
R14902 VSS.n5752 VSS.n2649 0.04025
R14903 VSS.n5753 VSS.n5752 0.04025
R14904 VSS.n5754 VSS.n5753 0.04025
R14905 VSS.n5754 VSS.n2647 0.04025
R14906 VSS.n5758 VSS.n2647 0.04025
R14907 VSS.n5759 VSS.n5758 0.04025
R14908 VSS.n5760 VSS.n5759 0.04025
R14909 VSS.n5760 VSS.n2645 0.04025
R14910 VSS.n5764 VSS.n2645 0.04025
R14911 VSS.n5765 VSS.n5764 0.04025
R14912 VSS.n5766 VSS.n5765 0.04025
R14913 VSS.n5766 VSS.n2643 0.04025
R14914 VSS.n5770 VSS.n2643 0.04025
R14915 VSS.n5771 VSS.n5770 0.04025
R14916 VSS.n5772 VSS.n5771 0.04025
R14917 VSS.n5772 VSS.n2641 0.04025
R14918 VSS.n5776 VSS.n2641 0.04025
R14919 VSS.n5777 VSS.n5776 0.04025
R14920 VSS.n5778 VSS.n5777 0.04025
R14921 VSS.n5778 VSS.n2639 0.04025
R14922 VSS.n5782 VSS.n2639 0.04025
R14923 VSS.n5783 VSS.n5782 0.04025
R14924 VSS.n5784 VSS.n5783 0.04025
R14925 VSS.n5784 VSS.n2637 0.04025
R14926 VSS.n5788 VSS.n2637 0.04025
R14927 VSS.n5789 VSS.n5788 0.04025
R14928 VSS.n5790 VSS.n5789 0.04025
R14929 VSS.n5790 VSS.n2635 0.04025
R14930 VSS.n5794 VSS.n2635 0.04025
R14931 VSS.n5795 VSS.n5794 0.04025
R14932 VSS.n5796 VSS.n5795 0.04025
R14933 VSS.n5796 VSS.n2633 0.04025
R14934 VSS.n5800 VSS.n2633 0.04025
R14935 VSS.n5801 VSS.n5800 0.04025
R14936 VSS.n5802 VSS.n5801 0.04025
R14937 VSS.n5802 VSS.n2631 0.04025
R14938 VSS.n5806 VSS.n2631 0.04025
R14939 VSS.n5807 VSS.n5806 0.04025
R14940 VSS.n5808 VSS.n5807 0.04025
R14941 VSS.n5808 VSS.n2629 0.04025
R14942 VSS.n5812 VSS.n2629 0.04025
R14943 VSS.n5813 VSS.n5812 0.04025
R14944 VSS.n5814 VSS.n5813 0.04025
R14945 VSS.n5814 VSS.n2627 0.04025
R14946 VSS.n5818 VSS.n2627 0.04025
R14947 VSS.n5819 VSS.n5818 0.04025
R14948 VSS.n5820 VSS.n5819 0.04025
R14949 VSS.n5820 VSS.n2625 0.04025
R14950 VSS.n5824 VSS.n2625 0.04025
R14951 VSS.n5825 VSS.n5824 0.04025
R14952 VSS.n5826 VSS.n5825 0.04025
R14953 VSS.n5826 VSS.n2623 0.04025
R14954 VSS.n5830 VSS.n2623 0.04025
R14955 VSS.n5831 VSS.n5830 0.04025
R14956 VSS.n5832 VSS.n5831 0.04025
R14957 VSS.n5832 VSS.n2621 0.04025
R14958 VSS.n5836 VSS.n2621 0.04025
R14959 VSS.n5837 VSS.n5836 0.04025
R14960 VSS.n5838 VSS.n5837 0.04025
R14961 VSS.n5838 VSS.n2619 0.04025
R14962 VSS.n5842 VSS.n2619 0.04025
R14963 VSS.n5843 VSS.n5842 0.04025
R14964 VSS.n5844 VSS.n5843 0.04025
R14965 VSS.n5844 VSS.n2617 0.04025
R14966 VSS.n5848 VSS.n2617 0.04025
R14967 VSS.n5849 VSS.n5848 0.04025
R14968 VSS.n5850 VSS.n5849 0.04025
R14969 VSS.n5850 VSS.n2615 0.04025
R14970 VSS.n5854 VSS.n2615 0.04025
R14971 VSS.n5855 VSS.n5854 0.04025
R14972 VSS.n5856 VSS.n5855 0.04025
R14973 VSS.n5856 VSS.n2613 0.04025
R14974 VSS.n5860 VSS.n2613 0.04025
R14975 VSS.n5861 VSS.n5860 0.04025
R14976 VSS.n5862 VSS.n5861 0.04025
R14977 VSS.n5862 VSS.n2611 0.04025
R14978 VSS.n5866 VSS.n2611 0.04025
R14979 VSS.n5867 VSS.n5866 0.04025
R14980 VSS.n5868 VSS.n5867 0.04025
R14981 VSS.n5868 VSS.n2609 0.04025
R14982 VSS.n5872 VSS.n2609 0.04025
R14983 VSS.n5873 VSS.n5872 0.04025
R14984 VSS.n5874 VSS.n5873 0.04025
R14985 VSS.n5874 VSS.n2607 0.04025
R14986 VSS.n5878 VSS.n2607 0.04025
R14987 VSS.n5879 VSS.n5878 0.04025
R14988 VSS.n5880 VSS.n5879 0.04025
R14989 VSS.n5880 VSS.n2605 0.04025
R14990 VSS.n5884 VSS.n2605 0.04025
R14991 VSS.n5885 VSS.n5884 0.04025
R14992 VSS.n5886 VSS.n5885 0.04025
R14993 VSS.n5886 VSS.n2603 0.04025
R14994 VSS.n5890 VSS.n2603 0.04025
R14995 VSS.n5891 VSS.n5890 0.04025
R14996 VSS.n5892 VSS.n5891 0.04025
R14997 VSS.n5892 VSS.n2601 0.04025
R14998 VSS.n5896 VSS.n2601 0.04025
R14999 VSS.n5897 VSS.n5896 0.04025
R15000 VSS.n5898 VSS.n5897 0.04025
R15001 VSS.n5898 VSS.n2599 0.04025
R15002 VSS.n5902 VSS.n2599 0.04025
R15003 VSS.n5903 VSS.n5902 0.04025
R15004 VSS.n5904 VSS.n5903 0.04025
R15005 VSS.n5904 VSS.n2597 0.04025
R15006 VSS.n5908 VSS.n2597 0.04025
R15007 VSS.n5909 VSS.n5908 0.04025
R15008 VSS.n5910 VSS.n5909 0.04025
R15009 VSS.n5910 VSS.n2595 0.04025
R15010 VSS.n5914 VSS.n2595 0.04025
R15011 VSS.n5915 VSS.n5914 0.04025
R15012 VSS.n5916 VSS.n5915 0.04025
R15013 VSS.n5916 VSS.n2593 0.04025
R15014 VSS.n5920 VSS.n2593 0.04025
R15015 VSS.n5921 VSS.n5920 0.04025
R15016 VSS.n5922 VSS.n5921 0.04025
R15017 VSS.n5922 VSS.n2591 0.04025
R15018 VSS.n5926 VSS.n2591 0.04025
R15019 VSS.n5927 VSS.n5926 0.04025
R15020 VSS.n5928 VSS.n5927 0.04025
R15021 VSS.n5928 VSS.n2589 0.04025
R15022 VSS.n5932 VSS.n2589 0.04025
R15023 VSS.n5933 VSS.n5932 0.04025
R15024 VSS.n5934 VSS.n5933 0.04025
R15025 VSS.n5934 VSS.n2587 0.04025
R15026 VSS.n5938 VSS.n2587 0.04025
R15027 VSS.n5939 VSS.n5938 0.04025
R15028 VSS.n5940 VSS.n5939 0.04025
R15029 VSS.n5940 VSS.n2585 0.04025
R15030 VSS.n5944 VSS.n2585 0.04025
R15031 VSS.n5945 VSS.n5944 0.04025
R15032 VSS.n5946 VSS.n5945 0.04025
R15033 VSS.n5946 VSS.n2583 0.04025
R15034 VSS.n5950 VSS.n2583 0.04025
R15035 VSS.n5951 VSS.n5950 0.04025
R15036 VSS.n5952 VSS.n5951 0.04025
R15037 VSS.n5952 VSS.n2581 0.04025
R15038 VSS.n5956 VSS.n2581 0.04025
R15039 VSS.n5957 VSS.n5956 0.04025
R15040 VSS.n5958 VSS.n5957 0.04025
R15041 VSS.n5958 VSS.n2579 0.04025
R15042 VSS.n5962 VSS.n2579 0.04025
R15043 VSS.n5963 VSS.n5962 0.04025
R15044 VSS.n5964 VSS.n5963 0.04025
R15045 VSS.n5964 VSS.n2577 0.04025
R15046 VSS.n5968 VSS.n2577 0.04025
R15047 VSS.n5969 VSS.n5968 0.04025
R15048 VSS.n5970 VSS.n5969 0.04025
R15049 VSS.n5970 VSS.n2575 0.04025
R15050 VSS.n5974 VSS.n2575 0.04025
R15051 VSS.n5975 VSS.n5974 0.04025
R15052 VSS.n5976 VSS.n5975 0.04025
R15053 VSS.n5976 VSS.n2573 0.04025
R15054 VSS.n5980 VSS.n2573 0.04025
R15055 VSS.n5981 VSS.n5980 0.04025
R15056 VSS.n5982 VSS.n5981 0.04025
R15057 VSS.n5982 VSS.n2571 0.04025
R15058 VSS.n5986 VSS.n2571 0.04025
R15059 VSS.n5987 VSS.n5986 0.04025
R15060 VSS.n5988 VSS.n5987 0.04025
R15061 VSS.n5988 VSS.n2569 0.04025
R15062 VSS.n5992 VSS.n2569 0.04025
R15063 VSS.n5993 VSS.n5992 0.04025
R15064 VSS.n5994 VSS.n5993 0.04025
R15065 VSS.n5994 VSS.n2567 0.04025
R15066 VSS.n5998 VSS.n2567 0.04025
R15067 VSS.n5999 VSS.n5998 0.04025
R15068 VSS.n6000 VSS.n5999 0.04025
R15069 VSS.n6000 VSS.n2565 0.04025
R15070 VSS.n6004 VSS.n2565 0.04025
R15071 VSS.n6005 VSS.n6004 0.04025
R15072 VSS.n6006 VSS.n6005 0.04025
R15073 VSS.n6006 VSS.n2563 0.04025
R15074 VSS.n6010 VSS.n2563 0.04025
R15075 VSS.n6011 VSS.n6010 0.04025
R15076 VSS.n6012 VSS.n6011 0.04025
R15077 VSS.n6012 VSS.n2561 0.04025
R15078 VSS.n6016 VSS.n2561 0.04025
R15079 VSS.n6017 VSS.n6016 0.04025
R15080 VSS.n6018 VSS.n6017 0.04025
R15081 VSS.n6018 VSS.n2559 0.04025
R15082 VSS.n6022 VSS.n2559 0.04025
R15083 VSS.n6023 VSS.n6022 0.04025
R15084 VSS.n6024 VSS.n6023 0.04025
R15085 VSS.n6024 VSS.n2557 0.04025
R15086 VSS.n6028 VSS.n2557 0.04025
R15087 VSS.n6029 VSS.n6028 0.04025
R15088 VSS.n6030 VSS.n6029 0.04025
R15089 VSS.n6030 VSS.n2555 0.04025
R15090 VSS.n6034 VSS.n2555 0.04025
R15091 VSS.n6035 VSS.n6034 0.04025
R15092 VSS.n6036 VSS.n6035 0.04025
R15093 VSS.n6036 VSS.n2553 0.04025
R15094 VSS.n6040 VSS.n2553 0.04025
R15095 VSS.n6041 VSS.n6040 0.04025
R15096 VSS.n6042 VSS.n6041 0.04025
R15097 VSS.n6042 VSS.n2551 0.04025
R15098 VSS.n6046 VSS.n2551 0.04025
R15099 VSS.n6047 VSS.n6046 0.04025
R15100 VSS.n6048 VSS.n6047 0.04025
R15101 VSS.n6048 VSS.n2549 0.04025
R15102 VSS.n6052 VSS.n2549 0.04025
R15103 VSS.n6053 VSS.n6052 0.04025
R15104 VSS.n6054 VSS.n6053 0.04025
R15105 VSS.n6054 VSS.n2547 0.04025
R15106 VSS.n6058 VSS.n2547 0.04025
R15107 VSS.n6059 VSS.n6058 0.04025
R15108 VSS.n6060 VSS.n6059 0.04025
R15109 VSS.n6060 VSS.n2545 0.04025
R15110 VSS.n6064 VSS.n2545 0.04025
R15111 VSS.n6065 VSS.n6064 0.04025
R15112 VSS.n6066 VSS.n6065 0.04025
R15113 VSS.n6066 VSS.n2543 0.04025
R15114 VSS.n6070 VSS.n2543 0.04025
R15115 VSS.n6071 VSS.n6070 0.04025
R15116 VSS.n6072 VSS.n6071 0.04025
R15117 VSS.n6072 VSS.n2541 0.04025
R15118 VSS.n6076 VSS.n2541 0.04025
R15119 VSS.n6077 VSS.n6076 0.04025
R15120 VSS.n6078 VSS.n6077 0.04025
R15121 VSS.n6078 VSS.n2539 0.04025
R15122 VSS.n6082 VSS.n2539 0.04025
R15123 VSS.n6083 VSS.n6082 0.04025
R15124 VSS.n6084 VSS.n6083 0.04025
R15125 VSS.n6084 VSS.n2537 0.04025
R15126 VSS.n6088 VSS.n2537 0.04025
R15127 VSS.n6089 VSS.n6088 0.04025
R15128 VSS.n6090 VSS.n6089 0.04025
R15129 VSS.n6090 VSS.n2535 0.04025
R15130 VSS.n6094 VSS.n2535 0.04025
R15131 VSS.n6095 VSS.n6094 0.04025
R15132 VSS.n6096 VSS.n6095 0.04025
R15133 VSS.n6096 VSS.n2533 0.04025
R15134 VSS.n6100 VSS.n2533 0.04025
R15135 VSS.n6101 VSS.n6100 0.04025
R15136 VSS.n6102 VSS.n6101 0.04025
R15137 VSS.n6102 VSS.n2531 0.04025
R15138 VSS.n6106 VSS.n2531 0.04025
R15139 VSS.n6107 VSS.n6106 0.04025
R15140 VSS.n6108 VSS.n6107 0.04025
R15141 VSS.n6108 VSS.n2529 0.04025
R15142 VSS.n6112 VSS.n2529 0.04025
R15143 VSS.n6113 VSS.n6112 0.04025
R15144 VSS.n6114 VSS.n6113 0.04025
R15145 VSS.n6114 VSS.n2527 0.04025
R15146 VSS.n6118 VSS.n2527 0.04025
R15147 VSS.n6119 VSS.n6118 0.04025
R15148 VSS.n6120 VSS.n6119 0.04025
R15149 VSS.n6120 VSS.n2525 0.04025
R15150 VSS.n6124 VSS.n2525 0.04025
R15151 VSS.n6125 VSS.n6124 0.04025
R15152 VSS.n6126 VSS.n6125 0.04025
R15153 VSS.n6126 VSS.n2523 0.04025
R15154 VSS.n6130 VSS.n2523 0.04025
R15155 VSS.n6131 VSS.n6130 0.04025
R15156 VSS.n6132 VSS.n6131 0.04025
R15157 VSS.n6132 VSS.n2521 0.04025
R15158 VSS.n6136 VSS.n2521 0.04025
R15159 VSS.n6137 VSS.n6136 0.04025
R15160 VSS.n6138 VSS.n6137 0.04025
R15161 VSS.n6138 VSS.n2519 0.04025
R15162 VSS.n6142 VSS.n2519 0.04025
R15163 VSS.n6143 VSS.n6142 0.04025
R15164 VSS.n6144 VSS.n6143 0.04025
R15165 VSS.n6144 VSS.n2517 0.04025
R15166 VSS.n6148 VSS.n2517 0.04025
R15167 VSS.n6149 VSS.n6148 0.04025
R15168 VSS.n6150 VSS.n6149 0.04025
R15169 VSS.n6150 VSS.n2515 0.04025
R15170 VSS.n6154 VSS.n2515 0.04025
R15171 VSS.n6155 VSS.n6154 0.04025
R15172 VSS.n6156 VSS.n6155 0.04025
R15173 VSS.n6156 VSS.n2513 0.04025
R15174 VSS.n6160 VSS.n2513 0.04025
R15175 VSS.n6161 VSS.n6160 0.04025
R15176 VSS.n6162 VSS.n6161 0.04025
R15177 VSS.n6162 VSS.n2511 0.04025
R15178 VSS.n6166 VSS.n2511 0.04025
R15179 VSS.n6167 VSS.n6166 0.04025
R15180 VSS.n6168 VSS.n6167 0.04025
R15181 VSS.n6168 VSS.n2509 0.04025
R15182 VSS.n6172 VSS.n2509 0.04025
R15183 VSS.n6173 VSS.n6172 0.04025
R15184 VSS.n6174 VSS.n6173 0.04025
R15185 VSS.n6174 VSS.n2507 0.04025
R15186 VSS.n6178 VSS.n2507 0.04025
R15187 VSS.n6179 VSS.n6178 0.04025
R15188 VSS.n6180 VSS.n6179 0.04025
R15189 VSS.n6180 VSS.n2505 0.04025
R15190 VSS.n6184 VSS.n2505 0.04025
R15191 VSS.n6185 VSS.n6184 0.04025
R15192 VSS.n6186 VSS.n6185 0.04025
R15193 VSS.n6186 VSS.n2503 0.04025
R15194 VSS.n6190 VSS.n2503 0.04025
R15195 VSS.n6191 VSS.n6190 0.04025
R15196 VSS.n6192 VSS.n6191 0.04025
R15197 VSS.n6192 VSS.n2501 0.04025
R15198 VSS.n6196 VSS.n2501 0.04025
R15199 VSS.n6197 VSS.n6196 0.04025
R15200 VSS.n6198 VSS.n6197 0.04025
R15201 VSS.n6198 VSS.n2499 0.04025
R15202 VSS.n6202 VSS.n2499 0.04025
R15203 VSS.n6203 VSS.n6202 0.04025
R15204 VSS.n6204 VSS.n6203 0.04025
R15205 VSS.n6204 VSS.n2497 0.04025
R15206 VSS.n6208 VSS.n2497 0.04025
R15207 VSS.n6209 VSS.n6208 0.04025
R15208 VSS.n6210 VSS.n6209 0.04025
R15209 VSS.n6210 VSS.n2495 0.04025
R15210 VSS.n6214 VSS.n2495 0.04025
R15211 VSS.n6215 VSS.n6214 0.04025
R15212 VSS.n6216 VSS.n6215 0.04025
R15213 VSS.n6216 VSS.n2493 0.04025
R15214 VSS.n6220 VSS.n2493 0.04025
R15215 VSS.n6221 VSS.n6220 0.04025
R15216 VSS.n6222 VSS.n6221 0.04025
R15217 VSS.n6222 VSS.n2491 0.04025
R15218 VSS.n6226 VSS.n2491 0.04025
R15219 VSS.n6227 VSS.n6226 0.04025
R15220 VSS.n6228 VSS.n6227 0.04025
R15221 VSS.n6228 VSS.n2489 0.04025
R15222 VSS.n6232 VSS.n2489 0.04025
R15223 VSS.n6233 VSS.n6232 0.04025
R15224 VSS.n6234 VSS.n6233 0.04025
R15225 VSS.n6234 VSS.n2487 0.04025
R15226 VSS.n6238 VSS.n2487 0.04025
R15227 VSS.n6239 VSS.n6238 0.04025
R15228 VSS.n6240 VSS.n6239 0.04025
R15229 VSS.n6240 VSS.n2485 0.04025
R15230 VSS.n6244 VSS.n2485 0.04025
R15231 VSS.n6245 VSS.n6244 0.04025
R15232 VSS.n6246 VSS.n6245 0.04025
R15233 VSS.n6246 VSS.n2483 0.04025
R15234 VSS.n6250 VSS.n2483 0.04025
R15235 VSS.n6251 VSS.n6250 0.04025
R15236 VSS.n6252 VSS.n6251 0.04025
R15237 VSS.n6252 VSS.n2481 0.04025
R15238 VSS.n6256 VSS.n2481 0.04025
R15239 VSS.n6257 VSS.n6256 0.04025
R15240 VSS.n6258 VSS.n6257 0.04025
R15241 VSS.n6258 VSS.n2479 0.04025
R15242 VSS.n6262 VSS.n2479 0.04025
R15243 VSS.n6263 VSS.n6262 0.04025
R15244 VSS.n6264 VSS.n6263 0.04025
R15245 VSS.n6264 VSS.n2477 0.04025
R15246 VSS.n6268 VSS.n2477 0.04025
R15247 VSS.n6269 VSS.n6268 0.04025
R15248 VSS.n6270 VSS.n6269 0.04025
R15249 VSS.n6270 VSS.n2475 0.04025
R15250 VSS.n6274 VSS.n2475 0.04025
R15251 VSS.n6275 VSS.n6274 0.04025
R15252 VSS.n6276 VSS.n6275 0.04025
R15253 VSS.n6276 VSS.n2473 0.04025
R15254 VSS.n6280 VSS.n2473 0.04025
R15255 VSS.n6281 VSS.n6280 0.04025
R15256 VSS.n6282 VSS.n6281 0.04025
R15257 VSS.n6282 VSS.n2471 0.04025
R15258 VSS.n6286 VSS.n2471 0.04025
R15259 VSS.n6287 VSS.n6286 0.04025
R15260 VSS.n6288 VSS.n6287 0.04025
R15261 VSS.n6288 VSS.n2469 0.04025
R15262 VSS.n6292 VSS.n2469 0.04025
R15263 VSS.n6293 VSS.n6292 0.04025
R15264 VSS.n6294 VSS.n6293 0.04025
R15265 VSS.n6294 VSS.n2467 0.04025
R15266 VSS.n6298 VSS.n2467 0.04025
R15267 VSS.n6299 VSS.n6298 0.04025
R15268 VSS.n6300 VSS.n6299 0.04025
R15269 VSS.n6300 VSS.n2465 0.04025
R15270 VSS.n6304 VSS.n2465 0.04025
R15271 VSS.n6305 VSS.n6304 0.04025
R15272 VSS.n6306 VSS.n6305 0.04025
R15273 VSS.n6306 VSS.n2463 0.04025
R15274 VSS.n6310 VSS.n2463 0.04025
R15275 VSS.n6311 VSS.n6310 0.04025
R15276 VSS.n6312 VSS.n6311 0.04025
R15277 VSS.n6312 VSS.n2461 0.04025
R15278 VSS.n6316 VSS.n2461 0.04025
R15279 VSS.n6317 VSS.n6316 0.04025
R15280 VSS.n6318 VSS.n6317 0.04025
R15281 VSS.n6318 VSS.n2459 0.04025
R15282 VSS.n6322 VSS.n2459 0.04025
R15283 VSS.n6323 VSS.n6322 0.04025
R15284 VSS.n6324 VSS.n6323 0.04025
R15285 VSS.n6324 VSS.n2457 0.04025
R15286 VSS.n6328 VSS.n2457 0.04025
R15287 VSS.n6329 VSS.n6328 0.04025
R15288 VSS.n6330 VSS.n6329 0.04025
R15289 VSS.n6330 VSS.n2455 0.04025
R15290 VSS.n6334 VSS.n2455 0.04025
R15291 VSS.n6335 VSS.n6334 0.04025
R15292 VSS.n6336 VSS.n6335 0.04025
R15293 VSS.n6336 VSS.n2453 0.04025
R15294 VSS.n6340 VSS.n2453 0.04025
R15295 VSS.n6341 VSS.n6340 0.04025
R15296 VSS.n6342 VSS.n6341 0.04025
R15297 VSS.n6342 VSS.n2451 0.04025
R15298 VSS.n6346 VSS.n2451 0.04025
R15299 VSS.n6347 VSS.n6346 0.04025
R15300 VSS.n6348 VSS.n6347 0.04025
R15301 VSS.n6348 VSS.n2449 0.04025
R15302 VSS.n6352 VSS.n2449 0.04025
R15303 VSS.n6353 VSS.n6352 0.04025
R15304 VSS.n6354 VSS.n6353 0.04025
R15305 VSS.n6354 VSS.n2447 0.04025
R15306 VSS.n6358 VSS.n2447 0.04025
R15307 VSS.n6359 VSS.n6358 0.04025
R15308 VSS.n6360 VSS.n6359 0.04025
R15309 VSS.n6360 VSS.n2445 0.04025
R15310 VSS.n6364 VSS.n2445 0.04025
R15311 VSS.n6365 VSS.n6364 0.04025
R15312 VSS.n6366 VSS.n6365 0.04025
R15313 VSS.n6366 VSS.n2443 0.04025
R15314 VSS.n6370 VSS.n2443 0.04025
R15315 VSS.n6371 VSS.n6370 0.04025
R15316 VSS.n6372 VSS.n6371 0.04025
R15317 VSS.n6372 VSS.n2441 0.04025
R15318 VSS.n6376 VSS.n2441 0.04025
R15319 VSS.n6377 VSS.n6376 0.04025
R15320 VSS.n6378 VSS.n6377 0.04025
R15321 VSS.n6378 VSS.n2439 0.04025
R15322 VSS.n6382 VSS.n2439 0.04025
R15323 VSS.n6383 VSS.n6382 0.04025
R15324 VSS.n6384 VSS.n6383 0.04025
R15325 VSS.n6384 VSS.n2437 0.04025
R15326 VSS.n6388 VSS.n2437 0.04025
R15327 VSS.n6389 VSS.n6388 0.04025
R15328 VSS.n6390 VSS.n6389 0.04025
R15329 VSS.n6390 VSS.n2435 0.04025
R15330 VSS.n6394 VSS.n2435 0.04025
R15331 VSS.n6395 VSS.n6394 0.04025
R15332 VSS.n6396 VSS.n6395 0.04025
R15333 VSS.n6396 VSS.n2433 0.04025
R15334 VSS.n6400 VSS.n2433 0.04025
R15335 VSS.n6401 VSS.n6400 0.04025
R15336 VSS.n6402 VSS.n6401 0.04025
R15337 VSS.n6402 VSS.n2431 0.04025
R15338 VSS.n6406 VSS.n2431 0.04025
R15339 VSS.n6407 VSS.n6406 0.04025
R15340 VSS.n6408 VSS.n6407 0.04025
R15341 VSS.n6408 VSS.n2429 0.04025
R15342 VSS.n6412 VSS.n2429 0.04025
R15343 VSS.n6413 VSS.n6412 0.04025
R15344 VSS.n6414 VSS.n6413 0.04025
R15345 VSS.n6414 VSS.n2427 0.04025
R15346 VSS.n6418 VSS.n2427 0.04025
R15347 VSS.n6419 VSS.n6418 0.04025
R15348 VSS.n6420 VSS.n6419 0.04025
R15349 VSS.n6420 VSS.n2425 0.04025
R15350 VSS.n6424 VSS.n2425 0.04025
R15351 VSS.n6425 VSS.n6424 0.04025
R15352 VSS.n6426 VSS.n6425 0.04025
R15353 VSS.n6426 VSS.n2423 0.04025
R15354 VSS.n6430 VSS.n2423 0.04025
R15355 VSS.n6431 VSS.n6430 0.04025
R15356 VSS.n6432 VSS.n6431 0.04025
R15357 VSS.n6432 VSS.n2421 0.04025
R15358 VSS.n6436 VSS.n2421 0.04025
R15359 VSS.n6437 VSS.n6436 0.04025
R15360 VSS.n6438 VSS.n6437 0.04025
R15361 VSS.n6438 VSS.n2419 0.04025
R15362 VSS.n6442 VSS.n2419 0.04025
R15363 VSS.n6443 VSS.n6442 0.04025
R15364 VSS.n6444 VSS.n6443 0.04025
R15365 VSS.n6444 VSS.n2417 0.04025
R15366 VSS.n6448 VSS.n2417 0.04025
R15367 VSS.n6449 VSS.n6448 0.04025
R15368 VSS.n6450 VSS.n6449 0.04025
R15369 VSS.n6450 VSS.n2415 0.04025
R15370 VSS.n6454 VSS.n2415 0.04025
R15371 VSS.n6455 VSS.n6454 0.04025
R15372 VSS.n6456 VSS.n6455 0.04025
R15373 VSS.n6456 VSS.n2413 0.04025
R15374 VSS.n6460 VSS.n2413 0.04025
R15375 VSS.n6461 VSS.n6460 0.04025
R15376 VSS.n6462 VSS.n6461 0.04025
R15377 VSS.n6462 VSS.n2411 0.04025
R15378 VSS.n6466 VSS.n2411 0.04025
R15379 VSS.n6467 VSS.n6466 0.04025
R15380 VSS.n6468 VSS.n6467 0.04025
R15381 VSS.n6468 VSS.n2409 0.04025
R15382 VSS.n6472 VSS.n2409 0.04025
R15383 VSS.n6473 VSS.n6472 0.04025
R15384 VSS.n6474 VSS.n6473 0.04025
R15385 VSS.n6474 VSS.n2407 0.04025
R15386 VSS.n6478 VSS.n2407 0.04025
R15387 VSS.n6479 VSS.n6478 0.04025
R15388 VSS.n6480 VSS.n6479 0.04025
R15389 VSS.n6480 VSS.n2405 0.04025
R15390 VSS.n6484 VSS.n2405 0.04025
R15391 VSS.n6485 VSS.n6484 0.04025
R15392 VSS.n6486 VSS.n6485 0.04025
R15393 VSS.n6486 VSS.n2403 0.04025
R15394 VSS.n6490 VSS.n2403 0.04025
R15395 VSS.n6491 VSS.n6490 0.04025
R15396 VSS.n6492 VSS.n6491 0.04025
R15397 VSS.n6492 VSS.n2401 0.04025
R15398 VSS.n6496 VSS.n2401 0.04025
R15399 VSS.n6497 VSS.n6496 0.04025
R15400 VSS.n6498 VSS.n6497 0.04025
R15401 VSS.n6498 VSS.n2399 0.04025
R15402 VSS.n6502 VSS.n2399 0.04025
R15403 VSS.n6503 VSS.n6502 0.04025
R15404 VSS.n6504 VSS.n6503 0.04025
R15405 VSS.n6504 VSS.n2397 0.04025
R15406 VSS.n6508 VSS.n2397 0.04025
R15407 VSS.n6509 VSS.n6508 0.04025
R15408 VSS.n6510 VSS.n6509 0.04025
R15409 VSS.n6510 VSS.n2395 0.04025
R15410 VSS.n6514 VSS.n2395 0.04025
R15411 VSS.n6515 VSS.n6514 0.04025
R15412 VSS.n6516 VSS.n6515 0.04025
R15413 VSS.n6516 VSS.n2393 0.04025
R15414 VSS.n6520 VSS.n2393 0.04025
R15415 VSS.n6521 VSS.n6520 0.04025
R15416 VSS.n6522 VSS.n6521 0.04025
R15417 VSS.n6522 VSS.n2391 0.04025
R15418 VSS.n6526 VSS.n2391 0.04025
R15419 VSS.n6527 VSS.n6526 0.04025
R15420 VSS.n6528 VSS.n6527 0.04025
R15421 VSS.n6528 VSS.n2389 0.04025
R15422 VSS.n6532 VSS.n2389 0.04025
R15423 VSS.n6533 VSS.n6532 0.04025
R15424 VSS.n6534 VSS.n6533 0.04025
R15425 VSS.n6534 VSS.n2387 0.04025
R15426 VSS.n6538 VSS.n2387 0.04025
R15427 VSS.n6539 VSS.n6538 0.04025
R15428 VSS.n6540 VSS.n6539 0.04025
R15429 VSS.n6540 VSS.n2385 0.04025
R15430 VSS.n6544 VSS.n2385 0.04025
R15431 VSS.n6545 VSS.n6544 0.04025
R15432 VSS.n6546 VSS.n6545 0.04025
R15433 VSS.n6546 VSS.n2383 0.04025
R15434 VSS.n6550 VSS.n2383 0.04025
R15435 VSS.n6551 VSS.n6550 0.04025
R15436 VSS.n6552 VSS.n6551 0.04025
R15437 VSS.n6552 VSS.n2381 0.04025
R15438 VSS.n6556 VSS.n2381 0.04025
R15439 VSS.n6557 VSS.n6556 0.04025
R15440 VSS.n6558 VSS.n6557 0.04025
R15441 VSS.n6558 VSS.n2379 0.04025
R15442 VSS.n6562 VSS.n2379 0.04025
R15443 VSS.n6563 VSS.n6562 0.04025
R15444 VSS.n6564 VSS.n6563 0.04025
R15445 VSS.n6564 VSS.n2377 0.04025
R15446 VSS.n6568 VSS.n2377 0.04025
R15447 VSS.n6569 VSS.n6568 0.04025
R15448 VSS.n6570 VSS.n6569 0.04025
R15449 VSS.n6570 VSS.n2375 0.04025
R15450 VSS.n6574 VSS.n2375 0.04025
R15451 VSS.n6575 VSS.n6574 0.04025
R15452 VSS.n6576 VSS.n6575 0.04025
R15453 VSS.n6576 VSS.n2373 0.04025
R15454 VSS.n6580 VSS.n2373 0.04025
R15455 VSS.n6581 VSS.n6580 0.04025
R15456 VSS.n6582 VSS.n6581 0.04025
R15457 VSS.n6582 VSS.n2371 0.04025
R15458 VSS.n6586 VSS.n2371 0.04025
R15459 VSS.n6587 VSS.n6586 0.04025
R15460 VSS.n6588 VSS.n6587 0.04025
R15461 VSS.n6588 VSS.n2369 0.04025
R15462 VSS.n6592 VSS.n2369 0.04025
R15463 VSS.n6593 VSS.n6592 0.04025
R15464 VSS.n6594 VSS.n6593 0.04025
R15465 VSS.n6594 VSS.n2367 0.04025
R15466 VSS.n6598 VSS.n2367 0.04025
R15467 VSS.n6599 VSS.n6598 0.04025
R15468 VSS.n6600 VSS.n6599 0.04025
R15469 VSS.n6600 VSS.n2365 0.04025
R15470 VSS.n6604 VSS.n2365 0.04025
R15471 VSS.n6605 VSS.n6604 0.04025
R15472 VSS.n6606 VSS.n6605 0.04025
R15473 VSS.n6606 VSS.n2363 0.04025
R15474 VSS.n6610 VSS.n2363 0.04025
R15475 VSS.n6611 VSS.n6610 0.04025
R15476 VSS.n6612 VSS.n6611 0.04025
R15477 VSS.n6612 VSS.n2361 0.04025
R15478 VSS.n6616 VSS.n2361 0.04025
R15479 VSS.n6617 VSS.n6616 0.04025
R15480 VSS.n6618 VSS.n6617 0.04025
R15481 VSS.n6618 VSS.n2359 0.04025
R15482 VSS.n6622 VSS.n2359 0.04025
R15483 VSS.n6623 VSS.n6622 0.04025
R15484 VSS.n6624 VSS.n6623 0.04025
R15485 VSS.n6624 VSS.n2357 0.04025
R15486 VSS.n6628 VSS.n2357 0.04025
R15487 VSS.n6629 VSS.n6628 0.04025
R15488 VSS.n6630 VSS.n6629 0.04025
R15489 VSS.n6630 VSS.n2355 0.04025
R15490 VSS.n6634 VSS.n2355 0.04025
R15491 VSS.n6635 VSS.n6634 0.04025
R15492 VSS.n6636 VSS.n6635 0.04025
R15493 VSS.n6636 VSS.n2353 0.04025
R15494 VSS.n6640 VSS.n2353 0.04025
R15495 VSS.n6641 VSS.n6640 0.04025
R15496 VSS.n6642 VSS.n6641 0.04025
R15497 VSS.n6642 VSS.n2351 0.04025
R15498 VSS.n6646 VSS.n2351 0.04025
R15499 VSS.n6647 VSS.n6646 0.04025
R15500 VSS.n6648 VSS.n6647 0.04025
R15501 VSS.n6648 VSS.n2349 0.04025
R15502 VSS.n6652 VSS.n2349 0.04025
R15503 VSS.n6653 VSS.n6652 0.04025
R15504 VSS.n6654 VSS.n6653 0.04025
R15505 VSS.n6654 VSS.n2347 0.04025
R15506 VSS.n6658 VSS.n2347 0.04025
R15507 VSS.n6659 VSS.n6658 0.04025
R15508 VSS.n6660 VSS.n6659 0.04025
R15509 VSS.n6660 VSS.n2345 0.04025
R15510 VSS.n6664 VSS.n2345 0.04025
R15511 VSS.n6665 VSS.n6664 0.04025
R15512 VSS.n6666 VSS.n6665 0.04025
R15513 VSS.n6666 VSS.n2343 0.04025
R15514 VSS.n6670 VSS.n2343 0.04025
R15515 VSS.n6671 VSS.n6670 0.04025
R15516 VSS.n6672 VSS.n6671 0.04025
R15517 VSS.n6672 VSS.n2341 0.04025
R15518 VSS.n6676 VSS.n2341 0.04025
R15519 VSS.n6677 VSS.n6676 0.04025
R15520 VSS.n6678 VSS.n6677 0.04025
R15521 VSS.n6678 VSS.n2339 0.04025
R15522 VSS.n6682 VSS.n2339 0.04025
R15523 VSS.n6683 VSS.n6682 0.04025
R15524 VSS.n6684 VSS.n6683 0.04025
R15525 VSS.n6684 VSS.n2337 0.04025
R15526 VSS.n6688 VSS.n2337 0.04025
R15527 VSS.n6689 VSS.n6688 0.04025
R15528 VSS.n6690 VSS.n6689 0.04025
R15529 VSS.n6690 VSS.n2335 0.04025
R15530 VSS.n6694 VSS.n2335 0.04025
R15531 VSS.n6695 VSS.n6694 0.04025
R15532 VSS.n6696 VSS.n6695 0.04025
R15533 VSS.n6696 VSS.n2333 0.04025
R15534 VSS.n6700 VSS.n2333 0.04025
R15535 VSS.n6701 VSS.n6700 0.04025
R15536 VSS.n6702 VSS.n6701 0.04025
R15537 VSS.n6702 VSS.n2331 0.04025
R15538 VSS.n6706 VSS.n2331 0.04025
R15539 VSS.n6707 VSS.n6706 0.04025
R15540 VSS.n6708 VSS.n6707 0.04025
R15541 VSS.n6708 VSS.n2329 0.04025
R15542 VSS.n6712 VSS.n2329 0.04025
R15543 VSS.n6713 VSS.n6712 0.04025
R15544 VSS.n6714 VSS.n6713 0.04025
R15545 VSS.n6714 VSS.n2327 0.04025
R15546 VSS.n6718 VSS.n2327 0.04025
R15547 VSS.n6719 VSS.n6718 0.04025
R15548 VSS.n6720 VSS.n6719 0.04025
R15549 VSS.n6720 VSS.n2325 0.04025
R15550 VSS.n6724 VSS.n2325 0.04025
R15551 VSS.n6725 VSS.n6724 0.04025
R15552 VSS.n6726 VSS.n6725 0.04025
R15553 VSS.n6726 VSS.n2323 0.04025
R15554 VSS.n6730 VSS.n2323 0.04025
R15555 VSS.n6731 VSS.n6730 0.04025
R15556 VSS.n6732 VSS.n6731 0.04025
R15557 VSS.n6732 VSS.n2321 0.04025
R15558 VSS.n6736 VSS.n2321 0.04025
R15559 VSS.n6737 VSS.n6736 0.04025
R15560 VSS.n6738 VSS.n6737 0.04025
R15561 VSS.n6738 VSS.n2319 0.04025
R15562 VSS.n6742 VSS.n2319 0.04025
R15563 VSS.n6743 VSS.n6742 0.04025
R15564 VSS.n6744 VSS.n6743 0.04025
R15565 VSS.n6744 VSS.n2317 0.04025
R15566 VSS.n6748 VSS.n2317 0.04025
R15567 VSS.n6749 VSS.n6748 0.04025
R15568 VSS.n6750 VSS.n6749 0.04025
R15569 VSS.n6750 VSS.n2315 0.04025
R15570 VSS.n6754 VSS.n2315 0.04025
R15571 VSS.n6755 VSS.n6754 0.04025
R15572 VSS.n6756 VSS.n6755 0.04025
R15573 VSS.n6756 VSS.n2313 0.04025
R15574 VSS.n6760 VSS.n2313 0.04025
R15575 VSS.n6761 VSS.n6760 0.04025
R15576 VSS.n6762 VSS.n6761 0.04025
R15577 VSS.n6762 VSS.n2311 0.04025
R15578 VSS.n6766 VSS.n2311 0.04025
R15579 VSS.n6767 VSS.n6766 0.04025
R15580 VSS.n6768 VSS.n6767 0.04025
R15581 VSS.n6768 VSS.n2309 0.04025
R15582 VSS.n6772 VSS.n2309 0.04025
R15583 VSS.n6773 VSS.n6772 0.04025
R15584 VSS.n6774 VSS.n6773 0.04025
R15585 VSS.n6774 VSS.n2307 0.04025
R15586 VSS.n6778 VSS.n2307 0.04025
R15587 VSS.n6779 VSS.n6778 0.04025
R15588 VSS.n6780 VSS.n6779 0.04025
R15589 VSS.n6780 VSS.n2305 0.04025
R15590 VSS.n6784 VSS.n2305 0.04025
R15591 VSS.n6785 VSS.n6784 0.04025
R15592 VSS.n6786 VSS.n6785 0.04025
R15593 VSS.n6786 VSS.n2303 0.04025
R15594 VSS.n6790 VSS.n2303 0.04025
R15595 VSS.n6791 VSS.n6790 0.04025
R15596 VSS.n6792 VSS.n6791 0.04025
R15597 VSS.n6792 VSS.n2301 0.04025
R15598 VSS.n6796 VSS.n2301 0.04025
R15599 VSS.n6797 VSS.n6796 0.04025
R15600 VSS.n6798 VSS.n6797 0.04025
R15601 VSS.n6798 VSS.n2299 0.04025
R15602 VSS.n6802 VSS.n2299 0.04025
R15603 VSS.n6803 VSS.n6802 0.04025
R15604 VSS.n6804 VSS.n6803 0.04025
R15605 VSS.n6804 VSS.n2297 0.04025
R15606 VSS.n6808 VSS.n2297 0.04025
R15607 VSS.n6809 VSS.n6808 0.04025
R15608 VSS.n6810 VSS.n6809 0.04025
R15609 VSS.n6810 VSS.n2295 0.04025
R15610 VSS.n6814 VSS.n2295 0.04025
R15611 VSS.n6815 VSS.n6814 0.04025
R15612 VSS.n6816 VSS.n6815 0.04025
R15613 VSS.n6816 VSS.n2293 0.04025
R15614 VSS.n6820 VSS.n2293 0.04025
R15615 VSS.n6821 VSS.n6820 0.04025
R15616 VSS.n6822 VSS.n6821 0.04025
R15617 VSS.n6822 VSS.n2291 0.04025
R15618 VSS.n6826 VSS.n2291 0.04025
R15619 VSS.n6827 VSS.n6826 0.04025
R15620 VSS.n6828 VSS.n6827 0.04025
R15621 VSS.n6828 VSS.n2289 0.04025
R15622 VSS.n6832 VSS.n2289 0.04025
R15623 VSS.n6833 VSS.n6832 0.04025
R15624 VSS.n6834 VSS.n6833 0.04025
R15625 VSS.n6834 VSS.n2287 0.04025
R15626 VSS.n6838 VSS.n2287 0.04025
R15627 VSS.n6839 VSS.n6838 0.04025
R15628 VSS.n6840 VSS.n6839 0.04025
R15629 VSS.n6840 VSS.n2285 0.04025
R15630 VSS.n6844 VSS.n2285 0.04025
R15631 VSS.n6845 VSS.n6844 0.04025
R15632 VSS.n6846 VSS.n6845 0.04025
R15633 VSS.n6846 VSS.n2283 0.04025
R15634 VSS.n6850 VSS.n2283 0.04025
R15635 VSS.n6851 VSS.n6850 0.04025
R15636 VSS.n6852 VSS.n6851 0.04025
R15637 VSS.n6852 VSS.n2281 0.04025
R15638 VSS.n6856 VSS.n2281 0.04025
R15639 VSS.n6857 VSS.n6856 0.04025
R15640 VSS.n6858 VSS.n6857 0.04025
R15641 VSS.n6858 VSS.n2279 0.04025
R15642 VSS.n6862 VSS.n2279 0.04025
R15643 VSS.n6863 VSS.n6862 0.04025
R15644 VSS.n6864 VSS.n6863 0.04025
R15645 VSS.n6864 VSS.n2277 0.04025
R15646 VSS.n6868 VSS.n2277 0.04025
R15647 VSS.n6869 VSS.n6868 0.04025
R15648 VSS.n6870 VSS.n6869 0.04025
R15649 VSS.n6870 VSS.n2275 0.04025
R15650 VSS.n6874 VSS.n2275 0.04025
R15651 VSS.n6875 VSS.n6874 0.04025
R15652 VSS.n6876 VSS.n6875 0.04025
R15653 VSS.n6876 VSS.n2273 0.04025
R15654 VSS.n6880 VSS.n2273 0.04025
R15655 VSS.n6881 VSS.n6880 0.04025
R15656 VSS.n6882 VSS.n6881 0.04025
R15657 VSS.n6882 VSS.n2271 0.04025
R15658 VSS.n6886 VSS.n2271 0.04025
R15659 VSS.n6887 VSS.n6886 0.04025
R15660 VSS.n6888 VSS.n6887 0.04025
R15661 VSS.n6888 VSS.n2269 0.04025
R15662 VSS.n6892 VSS.n2269 0.04025
R15663 VSS.n6893 VSS.n6892 0.04025
R15664 VSS.n6894 VSS.n6893 0.04025
R15665 VSS.n6894 VSS.n2267 0.04025
R15666 VSS.n6898 VSS.n2267 0.04025
R15667 VSS.n6899 VSS.n6898 0.04025
R15668 VSS.n6900 VSS.n6899 0.04025
R15669 VSS.n6900 VSS.n2265 0.04025
R15670 VSS.n6904 VSS.n2265 0.04025
R15671 VSS.n6905 VSS.n6904 0.04025
R15672 VSS.n6906 VSS.n6905 0.04025
R15673 VSS.n8231 VSS.n8230 0.04025
R15674 VSS.n8230 VSS.n1823 0.04025
R15675 VSS.n8226 VSS.n1823 0.04025
R15676 VSS.n8226 VSS.n8225 0.04025
R15677 VSS.n8225 VSS.n8224 0.04025
R15678 VSS.n8224 VSS.n1825 0.04025
R15679 VSS.n8220 VSS.n1825 0.04025
R15680 VSS.n8220 VSS.n8219 0.04025
R15681 VSS.n8219 VSS.n8218 0.04025
R15682 VSS.n8218 VSS.n1827 0.04025
R15683 VSS.n8214 VSS.n1827 0.04025
R15684 VSS.n8214 VSS.n8213 0.04025
R15685 VSS.n8213 VSS.n8212 0.04025
R15686 VSS.n8212 VSS.n1829 0.04025
R15687 VSS.n8208 VSS.n1829 0.04025
R15688 VSS.n8208 VSS.n8207 0.04025
R15689 VSS.n8207 VSS.n8206 0.04025
R15690 VSS.n8206 VSS.n1831 0.04025
R15691 VSS.n8202 VSS.n1831 0.04025
R15692 VSS.n8202 VSS.n8201 0.04025
R15693 VSS.n8201 VSS.n8200 0.04025
R15694 VSS.n8200 VSS.n1833 0.04025
R15695 VSS.n8196 VSS.n1833 0.04025
R15696 VSS.n8196 VSS.n8195 0.04025
R15697 VSS.n8195 VSS.n8194 0.04025
R15698 VSS.n8194 VSS.n1835 0.04025
R15699 VSS.n8190 VSS.n1835 0.04025
R15700 VSS.n8190 VSS.n8189 0.04025
R15701 VSS.n8189 VSS.n8188 0.04025
R15702 VSS.n8188 VSS.n1837 0.04025
R15703 VSS.n8184 VSS.n1837 0.04025
R15704 VSS.n8184 VSS.n8183 0.04025
R15705 VSS.n8183 VSS.n8182 0.04025
R15706 VSS.n8182 VSS.n1839 0.04025
R15707 VSS.n8178 VSS.n1839 0.04025
R15708 VSS.n8178 VSS.n8177 0.04025
R15709 VSS.n8177 VSS.n8176 0.04025
R15710 VSS.n8176 VSS.n1841 0.04025
R15711 VSS.n8172 VSS.n1841 0.04025
R15712 VSS.n8172 VSS.n8171 0.04025
R15713 VSS.n8171 VSS.n8170 0.04025
R15714 VSS.n8170 VSS.n1843 0.04025
R15715 VSS.n8166 VSS.n1843 0.04025
R15716 VSS.n8166 VSS.n8165 0.04025
R15717 VSS.n8165 VSS.n8164 0.04025
R15718 VSS.n8164 VSS.n1845 0.04025
R15719 VSS.n8160 VSS.n1845 0.04025
R15720 VSS.n8160 VSS.n8159 0.04025
R15721 VSS.n8159 VSS.n8158 0.04025
R15722 VSS.n8158 VSS.n1847 0.04025
R15723 VSS.n8154 VSS.n1847 0.04025
R15724 VSS.n8154 VSS.n8153 0.04025
R15725 VSS.n8153 VSS.n8152 0.04025
R15726 VSS.n8152 VSS.n1849 0.04025
R15727 VSS.n8148 VSS.n1849 0.04025
R15728 VSS.n8148 VSS.n8147 0.04025
R15729 VSS.n8147 VSS.n8146 0.04025
R15730 VSS.n8146 VSS.n1851 0.04025
R15731 VSS.n8142 VSS.n1851 0.04025
R15732 VSS.n8142 VSS.n8141 0.04025
R15733 VSS.n8141 VSS.n8140 0.04025
R15734 VSS.n8140 VSS.n1853 0.04025
R15735 VSS.n8136 VSS.n1853 0.04025
R15736 VSS.n8136 VSS.n8135 0.04025
R15737 VSS.n8135 VSS.n8134 0.04025
R15738 VSS.n8134 VSS.n1855 0.04025
R15739 VSS.n8130 VSS.n1855 0.04025
R15740 VSS.n8130 VSS.n8129 0.04025
R15741 VSS.n8129 VSS.n8128 0.04025
R15742 VSS.n8128 VSS.n1857 0.04025
R15743 VSS.n8124 VSS.n1857 0.04025
R15744 VSS.n8124 VSS.n8123 0.04025
R15745 VSS.n8123 VSS.n8122 0.04025
R15746 VSS.n8122 VSS.n1859 0.04025
R15747 VSS.n8118 VSS.n1859 0.04025
R15748 VSS.n8118 VSS.n8117 0.04025
R15749 VSS.n8117 VSS.n8116 0.04025
R15750 VSS.n8116 VSS.n1861 0.04025
R15751 VSS.n8112 VSS.n1861 0.04025
R15752 VSS.n8112 VSS.n8111 0.04025
R15753 VSS.n8111 VSS.n8110 0.04025
R15754 VSS.n8110 VSS.n1863 0.04025
R15755 VSS.n8106 VSS.n1863 0.04025
R15756 VSS.n8106 VSS.n8105 0.04025
R15757 VSS.n8105 VSS.n8104 0.04025
R15758 VSS.n8104 VSS.n1865 0.04025
R15759 VSS.n8100 VSS.n1865 0.04025
R15760 VSS.n8100 VSS.n8099 0.04025
R15761 VSS.n8099 VSS.n8098 0.04025
R15762 VSS.n8098 VSS.n1867 0.04025
R15763 VSS.n8094 VSS.n1867 0.04025
R15764 VSS.n8094 VSS.n8093 0.04025
R15765 VSS.n8093 VSS.n8092 0.04025
R15766 VSS.n8092 VSS.n1869 0.04025
R15767 VSS.n8088 VSS.n1869 0.04025
R15768 VSS.n8088 VSS.n8087 0.04025
R15769 VSS.n8087 VSS.n8086 0.04025
R15770 VSS.n8086 VSS.n1871 0.04025
R15771 VSS.n8082 VSS.n1871 0.04025
R15772 VSS.n8082 VSS.n8081 0.04025
R15773 VSS.n8081 VSS.n8080 0.04025
R15774 VSS.n8080 VSS.n1873 0.04025
R15775 VSS.n8076 VSS.n1873 0.04025
R15776 VSS.n8076 VSS.n8075 0.04025
R15777 VSS.n8075 VSS.n8074 0.04025
R15778 VSS.n8074 VSS.n1875 0.04025
R15779 VSS.n8070 VSS.n1875 0.04025
R15780 VSS.n8070 VSS.n8069 0.04025
R15781 VSS.n8069 VSS.n8068 0.04025
R15782 VSS.n8068 VSS.n1877 0.04025
R15783 VSS.n8064 VSS.n1877 0.04025
R15784 VSS.n8064 VSS.n8063 0.04025
R15785 VSS.n8063 VSS.n8062 0.04025
R15786 VSS.n8062 VSS.n1879 0.04025
R15787 VSS.n8058 VSS.n1879 0.04025
R15788 VSS.n8058 VSS.n8057 0.04025
R15789 VSS.n8057 VSS.n8056 0.04025
R15790 VSS.n8056 VSS.n1881 0.04025
R15791 VSS.n8052 VSS.n1881 0.04025
R15792 VSS.n8052 VSS.n8051 0.04025
R15793 VSS.n8051 VSS.n8050 0.04025
R15794 VSS.n8050 VSS.n1883 0.04025
R15795 VSS.n8046 VSS.n1883 0.04025
R15796 VSS.n8046 VSS.n8045 0.04025
R15797 VSS.n8045 VSS.n8044 0.04025
R15798 VSS.n8044 VSS.n1885 0.04025
R15799 VSS.n8040 VSS.n1885 0.04025
R15800 VSS.n8040 VSS.n8039 0.04025
R15801 VSS.n8039 VSS.n8038 0.04025
R15802 VSS.n8038 VSS.n1887 0.04025
R15803 VSS.n8034 VSS.n1887 0.04025
R15804 VSS.n8034 VSS.n8033 0.04025
R15805 VSS.n8033 VSS.n8032 0.04025
R15806 VSS.n8032 VSS.n1889 0.04025
R15807 VSS.n8028 VSS.n1889 0.04025
R15808 VSS.n8028 VSS.n8027 0.04025
R15809 VSS.n8027 VSS.n8026 0.04025
R15810 VSS.n8026 VSS.n1891 0.04025
R15811 VSS.n8022 VSS.n1891 0.04025
R15812 VSS.n8022 VSS.n8021 0.04025
R15813 VSS.n8021 VSS.n8020 0.04025
R15814 VSS.n8020 VSS.n1893 0.04025
R15815 VSS.n8016 VSS.n1893 0.04025
R15816 VSS.n8016 VSS.n8015 0.04025
R15817 VSS.n8015 VSS.n8014 0.04025
R15818 VSS.n8014 VSS.n1895 0.04025
R15819 VSS.n8010 VSS.n1895 0.04025
R15820 VSS.n8010 VSS.n8009 0.04025
R15821 VSS.n8009 VSS.n8008 0.04025
R15822 VSS.n8008 VSS.n1897 0.04025
R15823 VSS.n8004 VSS.n1897 0.04025
R15824 VSS.n8004 VSS.n8003 0.04025
R15825 VSS.n8003 VSS.n8002 0.04025
R15826 VSS.n8002 VSS.n1899 0.04025
R15827 VSS.n7998 VSS.n1899 0.04025
R15828 VSS.n7998 VSS.n7997 0.04025
R15829 VSS.n7997 VSS.n7996 0.04025
R15830 VSS.n7996 VSS.n1901 0.04025
R15831 VSS.n7992 VSS.n1901 0.04025
R15832 VSS.n7992 VSS.n7991 0.04025
R15833 VSS.n7991 VSS.n7990 0.04025
R15834 VSS.n7990 VSS.n1903 0.04025
R15835 VSS.n7986 VSS.n1903 0.04025
R15836 VSS.n7986 VSS.n7985 0.04025
R15837 VSS.n7985 VSS.n7984 0.04025
R15838 VSS.n7984 VSS.n1905 0.04025
R15839 VSS.n7980 VSS.n1905 0.04025
R15840 VSS.n7980 VSS.n7979 0.04025
R15841 VSS.n7979 VSS.n7978 0.04025
R15842 VSS.n7978 VSS.n1907 0.04025
R15843 VSS.n7974 VSS.n1907 0.04025
R15844 VSS.n7974 VSS.n7973 0.04025
R15845 VSS.n7973 VSS.n7972 0.04025
R15846 VSS.n7972 VSS.n1909 0.04025
R15847 VSS.n7968 VSS.n1909 0.04025
R15848 VSS.n7968 VSS.n7967 0.04025
R15849 VSS.n7967 VSS.n7966 0.04025
R15850 VSS.n7966 VSS.n1911 0.04025
R15851 VSS.n7962 VSS.n1911 0.04025
R15852 VSS.n7962 VSS.n7961 0.04025
R15853 VSS.n7961 VSS.n7960 0.04025
R15854 VSS.n7960 VSS.n1913 0.04025
R15855 VSS.n7956 VSS.n1913 0.04025
R15856 VSS.n7956 VSS.n7955 0.04025
R15857 VSS.n7955 VSS.n7954 0.04025
R15858 VSS.n7954 VSS.n1915 0.04025
R15859 VSS.n7950 VSS.n1915 0.04025
R15860 VSS.n7950 VSS.n7949 0.04025
R15861 VSS.n7949 VSS.n7948 0.04025
R15862 VSS.n7948 VSS.n1917 0.04025
R15863 VSS.n7944 VSS.n1917 0.04025
R15864 VSS.n7944 VSS.n7943 0.04025
R15865 VSS.n7943 VSS.n7942 0.04025
R15866 VSS.n7942 VSS.n1919 0.04025
R15867 VSS.n7938 VSS.n1919 0.04025
R15868 VSS.n7938 VSS.n7937 0.04025
R15869 VSS.n7937 VSS.n7936 0.04025
R15870 VSS.n7936 VSS.n1921 0.04025
R15871 VSS.n7932 VSS.n1921 0.04025
R15872 VSS.n7932 VSS.n7931 0.04025
R15873 VSS.n7931 VSS.n7930 0.04025
R15874 VSS.n7930 VSS.n1923 0.04025
R15875 VSS.n7926 VSS.n1923 0.04025
R15876 VSS.n7926 VSS.n7925 0.04025
R15877 VSS.n7925 VSS.n7924 0.04025
R15878 VSS.n7924 VSS.n1925 0.04025
R15879 VSS.n7920 VSS.n1925 0.04025
R15880 VSS.n7920 VSS.n7919 0.04025
R15881 VSS.n7919 VSS.n7918 0.04025
R15882 VSS.n7918 VSS.n1927 0.04025
R15883 VSS.n7914 VSS.n1927 0.04025
R15884 VSS.n7914 VSS.n7913 0.04025
R15885 VSS.n7913 VSS.n7912 0.04025
R15886 VSS.n7912 VSS.n1929 0.04025
R15887 VSS.n7908 VSS.n1929 0.04025
R15888 VSS.n7908 VSS.n7907 0.04025
R15889 VSS.n7907 VSS.n7906 0.04025
R15890 VSS.n7906 VSS.n1931 0.04025
R15891 VSS.n7902 VSS.n1931 0.04025
R15892 VSS.n7902 VSS.n7901 0.04025
R15893 VSS.n7901 VSS.n7900 0.04025
R15894 VSS.n7900 VSS.n1933 0.04025
R15895 VSS.n7896 VSS.n1933 0.04025
R15896 VSS.n7896 VSS.n7895 0.04025
R15897 VSS.n7895 VSS.n7894 0.04025
R15898 VSS.n7894 VSS.n1935 0.04025
R15899 VSS.n7890 VSS.n1935 0.04025
R15900 VSS.n7890 VSS.n7889 0.04025
R15901 VSS.n7889 VSS.n7888 0.04025
R15902 VSS.n7888 VSS.n1937 0.04025
R15903 VSS.n7884 VSS.n1937 0.04025
R15904 VSS.n7884 VSS.n7883 0.04025
R15905 VSS.n7883 VSS.n7882 0.04025
R15906 VSS.n7882 VSS.n1939 0.04025
R15907 VSS.n7878 VSS.n1939 0.04025
R15908 VSS.n7878 VSS.n7877 0.04025
R15909 VSS.n7877 VSS.n7876 0.04025
R15910 VSS.n7876 VSS.n1941 0.04025
R15911 VSS.n7872 VSS.n1941 0.04025
R15912 VSS.n7872 VSS.n7871 0.04025
R15913 VSS.n7871 VSS.n7870 0.04025
R15914 VSS.n7870 VSS.n1943 0.04025
R15915 VSS.n7866 VSS.n1943 0.04025
R15916 VSS.n7866 VSS.n7865 0.04025
R15917 VSS.n7865 VSS.n7864 0.04025
R15918 VSS.n7864 VSS.n1945 0.04025
R15919 VSS.n7860 VSS.n1945 0.04025
R15920 VSS.n7860 VSS.n7859 0.04025
R15921 VSS.n7859 VSS.n7858 0.04025
R15922 VSS.n7858 VSS.n1947 0.04025
R15923 VSS.n7854 VSS.n1947 0.04025
R15924 VSS.n7854 VSS.n7853 0.04025
R15925 VSS.n7853 VSS.n7852 0.04025
R15926 VSS.n7852 VSS.n1949 0.04025
R15927 VSS.n7848 VSS.n1949 0.04025
R15928 VSS.n7848 VSS.n7847 0.04025
R15929 VSS.n7847 VSS.n7846 0.04025
R15930 VSS.n7846 VSS.n1951 0.04025
R15931 VSS.n7842 VSS.n1951 0.04025
R15932 VSS.n7842 VSS.n7841 0.04025
R15933 VSS.n7841 VSS.n7840 0.04025
R15934 VSS.n7840 VSS.n1953 0.04025
R15935 VSS.n7836 VSS.n1953 0.04025
R15936 VSS.n7836 VSS.n7835 0.04025
R15937 VSS.n7835 VSS.n7834 0.04025
R15938 VSS.n7834 VSS.n1955 0.04025
R15939 VSS.n7830 VSS.n1955 0.04025
R15940 VSS.n7830 VSS.n7829 0.04025
R15941 VSS.n7829 VSS.n7828 0.04025
R15942 VSS.n7828 VSS.n1957 0.04025
R15943 VSS.n7824 VSS.n1957 0.04025
R15944 VSS.n7824 VSS.n7823 0.04025
R15945 VSS.n7823 VSS.n7822 0.04025
R15946 VSS.n7822 VSS.n1959 0.04025
R15947 VSS.n7818 VSS.n1959 0.04025
R15948 VSS.n7818 VSS.n7817 0.04025
R15949 VSS.n7817 VSS.n7816 0.04025
R15950 VSS.n7816 VSS.n1961 0.04025
R15951 VSS.n7812 VSS.n1961 0.04025
R15952 VSS.n7812 VSS.n7811 0.04025
R15953 VSS.n7811 VSS.n7810 0.04025
R15954 VSS.n7810 VSS.n1963 0.04025
R15955 VSS.n7806 VSS.n1963 0.04025
R15956 VSS.n7806 VSS.n7805 0.04025
R15957 VSS.n7805 VSS.n7804 0.04025
R15958 VSS.n7804 VSS.n1965 0.04025
R15959 VSS.n7800 VSS.n1965 0.04025
R15960 VSS.n7800 VSS.n7799 0.04025
R15961 VSS.n7799 VSS.n7798 0.04025
R15962 VSS.n7798 VSS.n1967 0.04025
R15963 VSS.n7794 VSS.n1967 0.04025
R15964 VSS.n7794 VSS.n7793 0.04025
R15965 VSS.n7793 VSS.n7792 0.04025
R15966 VSS.n7792 VSS.n1969 0.04025
R15967 VSS.n7788 VSS.n1969 0.04025
R15968 VSS.n7788 VSS.n7787 0.04025
R15969 VSS.n7787 VSS.n7786 0.04025
R15970 VSS.n7786 VSS.n1971 0.04025
R15971 VSS.n7782 VSS.n1971 0.04025
R15972 VSS.n7782 VSS.n7781 0.04025
R15973 VSS.n7781 VSS.n7780 0.04025
R15974 VSS.n7780 VSS.n1973 0.04025
R15975 VSS.n7776 VSS.n1973 0.04025
R15976 VSS.n7776 VSS.n7775 0.04025
R15977 VSS.n7775 VSS.n7774 0.04025
R15978 VSS.n7774 VSS.n1975 0.04025
R15979 VSS.n7770 VSS.n1975 0.04025
R15980 VSS.n7770 VSS.n7769 0.04025
R15981 VSS.n7769 VSS.n7768 0.04025
R15982 VSS.n7768 VSS.n1977 0.04025
R15983 VSS.n7764 VSS.n1977 0.04025
R15984 VSS.n7764 VSS.n7763 0.04025
R15985 VSS.n7763 VSS.n7762 0.04025
R15986 VSS.n7762 VSS.n1979 0.04025
R15987 VSS.n7758 VSS.n1979 0.04025
R15988 VSS.n7758 VSS.n7757 0.04025
R15989 VSS.n7757 VSS.n7756 0.04025
R15990 VSS.n7756 VSS.n1981 0.04025
R15991 VSS.n7752 VSS.n1981 0.04025
R15992 VSS.n7752 VSS.n7751 0.04025
R15993 VSS.n7751 VSS.n7750 0.04025
R15994 VSS.n7750 VSS.n1983 0.04025
R15995 VSS.n7746 VSS.n1983 0.04025
R15996 VSS.n7746 VSS.n7745 0.04025
R15997 VSS.n7745 VSS.n7744 0.04025
R15998 VSS.n7744 VSS.n1985 0.04025
R15999 VSS.n7740 VSS.n1985 0.04025
R16000 VSS.n7740 VSS.n7739 0.04025
R16001 VSS.n7739 VSS.n7738 0.04025
R16002 VSS.n7738 VSS.n1987 0.04025
R16003 VSS.n7734 VSS.n1987 0.04025
R16004 VSS.n7734 VSS.n7733 0.04025
R16005 VSS.n7733 VSS.n7732 0.04025
R16006 VSS.n7732 VSS.n1989 0.04025
R16007 VSS.n7728 VSS.n1989 0.04025
R16008 VSS.n7728 VSS.n7727 0.04025
R16009 VSS.n7727 VSS.n7726 0.04025
R16010 VSS.n7726 VSS.n1991 0.04025
R16011 VSS.n7722 VSS.n1991 0.04025
R16012 VSS.n7722 VSS.n7721 0.04025
R16013 VSS.n7721 VSS.n7720 0.04025
R16014 VSS.n7720 VSS.n1993 0.04025
R16015 VSS.n7716 VSS.n1993 0.04025
R16016 VSS.n7716 VSS.n7715 0.04025
R16017 VSS.n7715 VSS.n7714 0.04025
R16018 VSS.n7714 VSS.n1995 0.04025
R16019 VSS.n7710 VSS.n1995 0.04025
R16020 VSS.n7710 VSS.n7709 0.04025
R16021 VSS.n7709 VSS.n7708 0.04025
R16022 VSS.n7708 VSS.n1997 0.04025
R16023 VSS.n7704 VSS.n1997 0.04025
R16024 VSS.n7704 VSS.n7703 0.04025
R16025 VSS.n7703 VSS.n7702 0.04025
R16026 VSS.n7702 VSS.n1999 0.04025
R16027 VSS.n7698 VSS.n1999 0.04025
R16028 VSS.n7698 VSS.n7697 0.04025
R16029 VSS.n7697 VSS.n7696 0.04025
R16030 VSS.n7696 VSS.n2001 0.04025
R16031 VSS.n7692 VSS.n2001 0.04025
R16032 VSS.n7692 VSS.n7691 0.04025
R16033 VSS.n7691 VSS.n7690 0.04025
R16034 VSS.n7690 VSS.n2003 0.04025
R16035 VSS.n7686 VSS.n2003 0.04025
R16036 VSS.n7686 VSS.n7685 0.04025
R16037 VSS.n7685 VSS.n7684 0.04025
R16038 VSS.n7684 VSS.n2005 0.04025
R16039 VSS.n7680 VSS.n2005 0.04025
R16040 VSS.n7680 VSS.n7679 0.04025
R16041 VSS.n7679 VSS.n7678 0.04025
R16042 VSS.n7678 VSS.n2007 0.04025
R16043 VSS.n7674 VSS.n2007 0.04025
R16044 VSS.n7674 VSS.n7673 0.04025
R16045 VSS.n7673 VSS.n7672 0.04025
R16046 VSS.n7672 VSS.n2009 0.04025
R16047 VSS.n7668 VSS.n2009 0.04025
R16048 VSS.n7668 VSS.n7667 0.04025
R16049 VSS.n7667 VSS.n7666 0.04025
R16050 VSS.n7666 VSS.n2011 0.04025
R16051 VSS.n7662 VSS.n2011 0.04025
R16052 VSS.n7662 VSS.n7661 0.04025
R16053 VSS.n7661 VSS.n7660 0.04025
R16054 VSS.n7660 VSS.n2013 0.04025
R16055 VSS.n7656 VSS.n2013 0.04025
R16056 VSS.n7656 VSS.n7655 0.04025
R16057 VSS.n7655 VSS.n7654 0.04025
R16058 VSS.n7654 VSS.n2015 0.04025
R16059 VSS.n7650 VSS.n2015 0.04025
R16060 VSS.n7650 VSS.n7649 0.04025
R16061 VSS.n7649 VSS.n7648 0.04025
R16062 VSS.n7648 VSS.n2017 0.04025
R16063 VSS.n7644 VSS.n2017 0.04025
R16064 VSS.n7644 VSS.n7643 0.04025
R16065 VSS.n7643 VSS.n7642 0.04025
R16066 VSS.n7642 VSS.n2019 0.04025
R16067 VSS.n7638 VSS.n2019 0.04025
R16068 VSS.n7638 VSS.n7637 0.04025
R16069 VSS.n7637 VSS.n7636 0.04025
R16070 VSS.n7636 VSS.n2021 0.04025
R16071 VSS.n7632 VSS.n2021 0.04025
R16072 VSS.n7632 VSS.n7631 0.04025
R16073 VSS.n7631 VSS.n7630 0.04025
R16074 VSS.n7630 VSS.n2023 0.04025
R16075 VSS.n7626 VSS.n2023 0.04025
R16076 VSS.n7626 VSS.n7625 0.04025
R16077 VSS.n7625 VSS.n7624 0.04025
R16078 VSS.n7624 VSS.n2025 0.04025
R16079 VSS.n7620 VSS.n2025 0.04025
R16080 VSS.n7620 VSS.n7619 0.04025
R16081 VSS.n7619 VSS.n7618 0.04025
R16082 VSS.n7618 VSS.n2027 0.04025
R16083 VSS.n7614 VSS.n2027 0.04025
R16084 VSS.n7614 VSS.n7613 0.04025
R16085 VSS.n7613 VSS.n7612 0.04025
R16086 VSS.n7612 VSS.n2029 0.04025
R16087 VSS.n7608 VSS.n2029 0.04025
R16088 VSS.n7608 VSS.n7607 0.04025
R16089 VSS.n7607 VSS.n7606 0.04025
R16090 VSS.n7606 VSS.n2031 0.04025
R16091 VSS.n7602 VSS.n2031 0.04025
R16092 VSS.n7602 VSS.n7601 0.04025
R16093 VSS.n7601 VSS.n7600 0.04025
R16094 VSS.n7600 VSS.n2033 0.04025
R16095 VSS.n7596 VSS.n2033 0.04025
R16096 VSS.n7596 VSS.n7595 0.04025
R16097 VSS.n7595 VSS.n7594 0.04025
R16098 VSS.n7594 VSS.n2035 0.04025
R16099 VSS.n7590 VSS.n2035 0.04025
R16100 VSS.n7590 VSS.n7589 0.04025
R16101 VSS.n7589 VSS.n7588 0.04025
R16102 VSS.n7588 VSS.n2037 0.04025
R16103 VSS.n7584 VSS.n2037 0.04025
R16104 VSS.n7584 VSS.n7583 0.04025
R16105 VSS.n7583 VSS.n7582 0.04025
R16106 VSS.n7582 VSS.n2039 0.04025
R16107 VSS.n7578 VSS.n2039 0.04025
R16108 VSS.n7578 VSS.n7577 0.04025
R16109 VSS.n7577 VSS.n7576 0.04025
R16110 VSS.n7576 VSS.n2041 0.04025
R16111 VSS.n7572 VSS.n2041 0.04025
R16112 VSS.n7572 VSS.n7571 0.04025
R16113 VSS.n7571 VSS.n7570 0.04025
R16114 VSS.n7570 VSS.n2043 0.04025
R16115 VSS.n7566 VSS.n2043 0.04025
R16116 VSS.n7566 VSS.n7565 0.04025
R16117 VSS.n7565 VSS.n7564 0.04025
R16118 VSS.n7564 VSS.n2045 0.04025
R16119 VSS.n7560 VSS.n2045 0.04025
R16120 VSS.n7560 VSS.n7559 0.04025
R16121 VSS.n7559 VSS.n7558 0.04025
R16122 VSS.n7558 VSS.n2047 0.04025
R16123 VSS.n7554 VSS.n2047 0.04025
R16124 VSS.n7554 VSS.n7553 0.04025
R16125 VSS.n7553 VSS.n7552 0.04025
R16126 VSS.n7552 VSS.n2049 0.04025
R16127 VSS.n7548 VSS.n2049 0.04025
R16128 VSS.n7548 VSS.n7547 0.04025
R16129 VSS.n7547 VSS.n7546 0.04025
R16130 VSS.n7546 VSS.n2051 0.04025
R16131 VSS.n7542 VSS.n2051 0.04025
R16132 VSS.n7542 VSS.n7541 0.04025
R16133 VSS.n7541 VSS.n7540 0.04025
R16134 VSS.n7540 VSS.n2053 0.04025
R16135 VSS.n7536 VSS.n2053 0.04025
R16136 VSS.n7536 VSS.n7535 0.04025
R16137 VSS.n7535 VSS.n7534 0.04025
R16138 VSS.n7534 VSS.n2055 0.04025
R16139 VSS.n7530 VSS.n2055 0.04025
R16140 VSS.n7530 VSS.n7529 0.04025
R16141 VSS.n7529 VSS.n7528 0.04025
R16142 VSS.n7528 VSS.n2057 0.04025
R16143 VSS.n7524 VSS.n2057 0.04025
R16144 VSS.n7524 VSS.n7523 0.04025
R16145 VSS.n7523 VSS.n7522 0.04025
R16146 VSS.n7522 VSS.n2059 0.04025
R16147 VSS.n7518 VSS.n2059 0.04025
R16148 VSS.n7518 VSS.n7517 0.04025
R16149 VSS.n7517 VSS.n7516 0.04025
R16150 VSS.n7516 VSS.n2061 0.04025
R16151 VSS.n7512 VSS.n2061 0.04025
R16152 VSS.n7512 VSS.n7511 0.04025
R16153 VSS.n7511 VSS.n7510 0.04025
R16154 VSS.n7510 VSS.n2063 0.04025
R16155 VSS.n7506 VSS.n2063 0.04025
R16156 VSS.n7506 VSS.n7505 0.04025
R16157 VSS.n7505 VSS.n7504 0.04025
R16158 VSS.n7504 VSS.n2065 0.04025
R16159 VSS.n7500 VSS.n2065 0.04025
R16160 VSS.n7500 VSS.n7499 0.04025
R16161 VSS.n7499 VSS.n7498 0.04025
R16162 VSS.n7498 VSS.n2067 0.04025
R16163 VSS.n7494 VSS.n2067 0.04025
R16164 VSS.n7494 VSS.n7493 0.04025
R16165 VSS.n7493 VSS.n7492 0.04025
R16166 VSS.n7492 VSS.n2069 0.04025
R16167 VSS.n7488 VSS.n2069 0.04025
R16168 VSS.n7488 VSS.n7487 0.04025
R16169 VSS.n7487 VSS.n7486 0.04025
R16170 VSS.n7486 VSS.n2071 0.04025
R16171 VSS.n7482 VSS.n2071 0.04025
R16172 VSS.n7482 VSS.n7481 0.04025
R16173 VSS.n7481 VSS.n7480 0.04025
R16174 VSS.n7480 VSS.n2073 0.04025
R16175 VSS.n7476 VSS.n2073 0.04025
R16176 VSS.n7476 VSS.n7475 0.04025
R16177 VSS.n7475 VSS.n7474 0.04025
R16178 VSS.n7474 VSS.n2075 0.04025
R16179 VSS.n7470 VSS.n2075 0.04025
R16180 VSS.n7470 VSS.n7469 0.04025
R16181 VSS.n7469 VSS.n7468 0.04025
R16182 VSS.n7468 VSS.n2077 0.04025
R16183 VSS.n7464 VSS.n2077 0.04025
R16184 VSS.n7464 VSS.n7463 0.04025
R16185 VSS.n7463 VSS.n7462 0.04025
R16186 VSS.n7462 VSS.n2079 0.04025
R16187 VSS.n7458 VSS.n2079 0.04025
R16188 VSS.n7458 VSS.n7457 0.04025
R16189 VSS.n7457 VSS.n7456 0.04025
R16190 VSS.n7456 VSS.n2081 0.04025
R16191 VSS.n7452 VSS.n2081 0.04025
R16192 VSS.n7452 VSS.n7451 0.04025
R16193 VSS.n7451 VSS.n7450 0.04025
R16194 VSS.n7450 VSS.n2083 0.04025
R16195 VSS.n7446 VSS.n2083 0.04025
R16196 VSS.n7446 VSS.n7445 0.04025
R16197 VSS.n7445 VSS.n7444 0.04025
R16198 VSS.n7444 VSS.n2085 0.04025
R16199 VSS.n7440 VSS.n2085 0.04025
R16200 VSS.n7440 VSS.n7439 0.04025
R16201 VSS.n7439 VSS.n7438 0.04025
R16202 VSS.n7438 VSS.n2087 0.04025
R16203 VSS.n7434 VSS.n2087 0.04025
R16204 VSS.n7434 VSS.n7433 0.04025
R16205 VSS.n7433 VSS.n7432 0.04025
R16206 VSS.n7432 VSS.n2089 0.04025
R16207 VSS.n7428 VSS.n2089 0.04025
R16208 VSS.n7428 VSS.n7427 0.04025
R16209 VSS.n7427 VSS.n7426 0.04025
R16210 VSS.n7426 VSS.n2091 0.04025
R16211 VSS.n7422 VSS.n2091 0.04025
R16212 VSS.n7422 VSS.n7421 0.04025
R16213 VSS.n7421 VSS.n7420 0.04025
R16214 VSS.n7420 VSS.n2093 0.04025
R16215 VSS.n7416 VSS.n2093 0.04025
R16216 VSS.n7416 VSS.n7415 0.04025
R16217 VSS.n7415 VSS.n7414 0.04025
R16218 VSS.n7414 VSS.n2095 0.04025
R16219 VSS.n7410 VSS.n2095 0.04025
R16220 VSS.n7410 VSS.n7409 0.04025
R16221 VSS.n7409 VSS.n7408 0.04025
R16222 VSS.n7408 VSS.n2097 0.04025
R16223 VSS.n7404 VSS.n2097 0.04025
R16224 VSS.n7404 VSS.n7403 0.04025
R16225 VSS.n7403 VSS.n7402 0.04025
R16226 VSS.n7402 VSS.n2099 0.04025
R16227 VSS.n7398 VSS.n2099 0.04025
R16228 VSS.n7398 VSS.n7397 0.04025
R16229 VSS.n7397 VSS.n7396 0.04025
R16230 VSS.n7396 VSS.n2101 0.04025
R16231 VSS.n7392 VSS.n2101 0.04025
R16232 VSS.n7392 VSS.n7391 0.04025
R16233 VSS.n7391 VSS.n7390 0.04025
R16234 VSS.n7390 VSS.n2103 0.04025
R16235 VSS.n7386 VSS.n2103 0.04025
R16236 VSS.n7386 VSS.n7385 0.04025
R16237 VSS.n7385 VSS.n7384 0.04025
R16238 VSS.n7384 VSS.n2105 0.04025
R16239 VSS.n7380 VSS.n2105 0.04025
R16240 VSS.n7380 VSS.n7379 0.04025
R16241 VSS.n7379 VSS.n7378 0.04025
R16242 VSS.n7378 VSS.n2107 0.04025
R16243 VSS.n7374 VSS.n2107 0.04025
R16244 VSS.n7374 VSS.n7373 0.04025
R16245 VSS.n7373 VSS.n7372 0.04025
R16246 VSS.n7372 VSS.n2109 0.04025
R16247 VSS.n7368 VSS.n2109 0.04025
R16248 VSS.n7368 VSS.n7367 0.04025
R16249 VSS.n7367 VSS.n7366 0.04025
R16250 VSS.n7366 VSS.n2111 0.04025
R16251 VSS.n7362 VSS.n2111 0.04025
R16252 VSS.n7362 VSS.n7361 0.04025
R16253 VSS.n7361 VSS.n7360 0.04025
R16254 VSS.n7360 VSS.n2113 0.04025
R16255 VSS.n7356 VSS.n2113 0.04025
R16256 VSS.n7356 VSS.n7355 0.04025
R16257 VSS.n7355 VSS.n7354 0.04025
R16258 VSS.n7354 VSS.n2115 0.04025
R16259 VSS.n7350 VSS.n2115 0.04025
R16260 VSS.n7350 VSS.n7349 0.04025
R16261 VSS.n7349 VSS.n7348 0.04025
R16262 VSS.n7348 VSS.n2117 0.04025
R16263 VSS.n7344 VSS.n2117 0.04025
R16264 VSS.n7344 VSS.n7343 0.04025
R16265 VSS.n7343 VSS.n7342 0.04025
R16266 VSS.n7342 VSS.n2119 0.04025
R16267 VSS.n7338 VSS.n2119 0.04025
R16268 VSS.n7338 VSS.n7337 0.04025
R16269 VSS.n7337 VSS.n7336 0.04025
R16270 VSS.n7336 VSS.n2121 0.04025
R16271 VSS.n7332 VSS.n2121 0.04025
R16272 VSS.n7332 VSS.n7331 0.04025
R16273 VSS.n7331 VSS.n7330 0.04025
R16274 VSS.n7330 VSS.n2123 0.04025
R16275 VSS.n7326 VSS.n2123 0.04025
R16276 VSS.n7326 VSS.n7325 0.04025
R16277 VSS.n7325 VSS.n7324 0.04025
R16278 VSS.n7324 VSS.n2125 0.04025
R16279 VSS.n7320 VSS.n2125 0.04025
R16280 VSS.n7320 VSS.n7319 0.04025
R16281 VSS.n7319 VSS.n7318 0.04025
R16282 VSS.n7318 VSS.n2127 0.04025
R16283 VSS.n7314 VSS.n2127 0.04025
R16284 VSS.n7314 VSS.n7313 0.04025
R16285 VSS.n7313 VSS.n7312 0.04025
R16286 VSS.n7312 VSS.n2129 0.04025
R16287 VSS.n7308 VSS.n2129 0.04025
R16288 VSS.n7308 VSS.n7307 0.04025
R16289 VSS.n7307 VSS.n7306 0.04025
R16290 VSS.n7306 VSS.n2131 0.04025
R16291 VSS.n7302 VSS.n2131 0.04025
R16292 VSS.n7302 VSS.n7301 0.04025
R16293 VSS.n7301 VSS.n7300 0.04025
R16294 VSS.n7300 VSS.n2133 0.04025
R16295 VSS.n7296 VSS.n2133 0.04025
R16296 VSS.n7296 VSS.n7295 0.04025
R16297 VSS.n7295 VSS.n7294 0.04025
R16298 VSS.n7294 VSS.n2135 0.04025
R16299 VSS.n7290 VSS.n2135 0.04025
R16300 VSS.n7290 VSS.n7289 0.04025
R16301 VSS.n7289 VSS.n7288 0.04025
R16302 VSS.n7288 VSS.n2137 0.04025
R16303 VSS.n7284 VSS.n2137 0.04025
R16304 VSS.n7284 VSS.n7283 0.04025
R16305 VSS.n7283 VSS.n7282 0.04025
R16306 VSS.n7282 VSS.n2139 0.04025
R16307 VSS.n7278 VSS.n2139 0.04025
R16308 VSS.n7278 VSS.n7277 0.04025
R16309 VSS.n7277 VSS.n7276 0.04025
R16310 VSS.n7276 VSS.n2141 0.04025
R16311 VSS.n7272 VSS.n2141 0.04025
R16312 VSS.n7272 VSS.n7271 0.04025
R16313 VSS.n7271 VSS.n7270 0.04025
R16314 VSS.n7270 VSS.n2143 0.04025
R16315 VSS.n7266 VSS.n2143 0.04025
R16316 VSS.n7266 VSS.n7265 0.04025
R16317 VSS.n7265 VSS.n7264 0.04025
R16318 VSS.n7264 VSS.n2145 0.04025
R16319 VSS.n7260 VSS.n2145 0.04025
R16320 VSS.n7260 VSS.n7259 0.04025
R16321 VSS.n7259 VSS.n7258 0.04025
R16322 VSS.n7258 VSS.n2147 0.04025
R16323 VSS.n7254 VSS.n2147 0.04025
R16324 VSS.n7254 VSS.n7253 0.04025
R16325 VSS.n7253 VSS.n7252 0.04025
R16326 VSS.n7252 VSS.n2149 0.04025
R16327 VSS.n7248 VSS.n2149 0.04025
R16328 VSS.n7248 VSS.n7247 0.04025
R16329 VSS.n7247 VSS.n7246 0.04025
R16330 VSS.n7246 VSS.n2151 0.04025
R16331 VSS.n7242 VSS.n2151 0.04025
R16332 VSS.n7242 VSS.n7241 0.04025
R16333 VSS.n7241 VSS.n7240 0.04025
R16334 VSS.n7240 VSS.n2153 0.04025
R16335 VSS.n7236 VSS.n2153 0.04025
R16336 VSS.n7236 VSS.n7235 0.04025
R16337 VSS.n7235 VSS.n7234 0.04025
R16338 VSS.n7234 VSS.n2155 0.04025
R16339 VSS.n7230 VSS.n2155 0.04025
R16340 VSS.n7230 VSS.n7229 0.04025
R16341 VSS.n7229 VSS.n7228 0.04025
R16342 VSS.n7228 VSS.n2157 0.04025
R16343 VSS.n7224 VSS.n2157 0.04025
R16344 VSS.n7224 VSS.n7223 0.04025
R16345 VSS.n7223 VSS.n7222 0.04025
R16346 VSS.n7222 VSS.n2159 0.04025
R16347 VSS.n7218 VSS.n2159 0.04025
R16348 VSS.n7218 VSS.n7217 0.04025
R16349 VSS.n7217 VSS.n7216 0.04025
R16350 VSS.n7216 VSS.n2161 0.04025
R16351 VSS.n7212 VSS.n2161 0.04025
R16352 VSS.n7212 VSS.n7211 0.04025
R16353 VSS.n7211 VSS.n7210 0.04025
R16354 VSS.n7210 VSS.n2163 0.04025
R16355 VSS.n7206 VSS.n2163 0.04025
R16356 VSS.n7206 VSS.n7205 0.04025
R16357 VSS.n7205 VSS.n7204 0.04025
R16358 VSS.n7204 VSS.n2165 0.04025
R16359 VSS.n7200 VSS.n2165 0.04025
R16360 VSS.n7200 VSS.n7199 0.04025
R16361 VSS.n7199 VSS.n7198 0.04025
R16362 VSS.n7198 VSS.n2167 0.04025
R16363 VSS.n7194 VSS.n2167 0.04025
R16364 VSS.n7194 VSS.n7193 0.04025
R16365 VSS.n7193 VSS.n7192 0.04025
R16366 VSS.n7192 VSS.n2169 0.04025
R16367 VSS.n7188 VSS.n2169 0.04025
R16368 VSS.n7188 VSS.n7187 0.04025
R16369 VSS.n7187 VSS.n7186 0.04025
R16370 VSS.n7186 VSS.n2171 0.04025
R16371 VSS.n7182 VSS.n2171 0.04025
R16372 VSS.n7182 VSS.n7181 0.04025
R16373 VSS.n7181 VSS.n7180 0.04025
R16374 VSS.n7180 VSS.n2173 0.04025
R16375 VSS.n7176 VSS.n2173 0.04025
R16376 VSS.n7176 VSS.n7175 0.04025
R16377 VSS.n7175 VSS.n7174 0.04025
R16378 VSS.n7174 VSS.n2175 0.04025
R16379 VSS.n7170 VSS.n2175 0.04025
R16380 VSS.n7170 VSS.n7169 0.04025
R16381 VSS.n7169 VSS.n7168 0.04025
R16382 VSS.n7168 VSS.n2177 0.04025
R16383 VSS.n7164 VSS.n2177 0.04025
R16384 VSS.n7164 VSS.n7163 0.04025
R16385 VSS.n7163 VSS.n7162 0.04025
R16386 VSS.n7162 VSS.n2179 0.04025
R16387 VSS.n7158 VSS.n2179 0.04025
R16388 VSS.n7158 VSS.n7157 0.04025
R16389 VSS.n7157 VSS.n7156 0.04025
R16390 VSS.n7156 VSS.n2181 0.04025
R16391 VSS.n7152 VSS.n2181 0.04025
R16392 VSS.n7152 VSS.n7151 0.04025
R16393 VSS.n7151 VSS.n7150 0.04025
R16394 VSS.n7150 VSS.n2183 0.04025
R16395 VSS.n7146 VSS.n2183 0.04025
R16396 VSS.n7146 VSS.n7145 0.04025
R16397 VSS.n7145 VSS.n7144 0.04025
R16398 VSS.n7144 VSS.n2185 0.04025
R16399 VSS.n7140 VSS.n2185 0.04025
R16400 VSS.n7140 VSS.n7139 0.04025
R16401 VSS.n7139 VSS.n7138 0.04025
R16402 VSS.n7138 VSS.n2187 0.04025
R16403 VSS.n7134 VSS.n2187 0.04025
R16404 VSS.n7134 VSS.n7133 0.04025
R16405 VSS.n7133 VSS.n7132 0.04025
R16406 VSS.n7132 VSS.n2189 0.04025
R16407 VSS.n7128 VSS.n2189 0.04025
R16408 VSS.n7128 VSS.n7127 0.04025
R16409 VSS.n7127 VSS.n7126 0.04025
R16410 VSS.n7126 VSS.n2191 0.04025
R16411 VSS.n7122 VSS.n2191 0.04025
R16412 VSS.n7122 VSS.n7121 0.04025
R16413 VSS.n7121 VSS.n7120 0.04025
R16414 VSS.n7120 VSS.n2193 0.04025
R16415 VSS.n7116 VSS.n2193 0.04025
R16416 VSS.n7116 VSS.n7115 0.04025
R16417 VSS.n7115 VSS.n7114 0.04025
R16418 VSS.n7114 VSS.n2195 0.04025
R16419 VSS.n7110 VSS.n2195 0.04025
R16420 VSS.n7110 VSS.n7109 0.04025
R16421 VSS.n7109 VSS.n7108 0.04025
R16422 VSS.n7108 VSS.n2197 0.04025
R16423 VSS.n7104 VSS.n2197 0.04025
R16424 VSS.n7104 VSS.n7103 0.04025
R16425 VSS.n7103 VSS.n7102 0.04025
R16426 VSS.n7102 VSS.n2199 0.04025
R16427 VSS.n7098 VSS.n2199 0.04025
R16428 VSS.n7098 VSS.n7097 0.04025
R16429 VSS.n7097 VSS.n7096 0.04025
R16430 VSS.n7096 VSS.n2201 0.04025
R16431 VSS.n7092 VSS.n2201 0.04025
R16432 VSS.n7092 VSS.n7091 0.04025
R16433 VSS.n7091 VSS.n7090 0.04025
R16434 VSS.n7090 VSS.n2203 0.04025
R16435 VSS.n7086 VSS.n2203 0.04025
R16436 VSS.n7086 VSS.n7085 0.04025
R16437 VSS.n7085 VSS.n7084 0.04025
R16438 VSS.n7084 VSS.n2205 0.04025
R16439 VSS.n7080 VSS.n2205 0.04025
R16440 VSS.n7080 VSS.n7079 0.04025
R16441 VSS.n7079 VSS.n7078 0.04025
R16442 VSS.n7078 VSS.n2207 0.04025
R16443 VSS.n7074 VSS.n2207 0.04025
R16444 VSS.n7074 VSS.n7073 0.04025
R16445 VSS.n7073 VSS.n7072 0.04025
R16446 VSS.n7072 VSS.n2209 0.04025
R16447 VSS.n7068 VSS.n2209 0.04025
R16448 VSS.n7068 VSS.n7067 0.04025
R16449 VSS.n7067 VSS.n7066 0.04025
R16450 VSS.n7066 VSS.n2211 0.04025
R16451 VSS.n7062 VSS.n2211 0.04025
R16452 VSS.n7062 VSS.n7061 0.04025
R16453 VSS.n7061 VSS.n7060 0.04025
R16454 VSS.n7060 VSS.n2213 0.04025
R16455 VSS.n7056 VSS.n2213 0.04025
R16456 VSS.n7056 VSS.n7055 0.04025
R16457 VSS.n7055 VSS.n7054 0.04025
R16458 VSS.n7054 VSS.n2215 0.04025
R16459 VSS.n7050 VSS.n2215 0.04025
R16460 VSS.n7050 VSS.n7049 0.04025
R16461 VSS.n7049 VSS.n7048 0.04025
R16462 VSS.n7048 VSS.n2217 0.04025
R16463 VSS.n7044 VSS.n2217 0.04025
R16464 VSS.n7044 VSS.n7043 0.04025
R16465 VSS.n7043 VSS.n7042 0.04025
R16466 VSS.n7042 VSS.n2219 0.04025
R16467 VSS.n7038 VSS.n2219 0.04025
R16468 VSS.n7038 VSS.n7037 0.04025
R16469 VSS.n7037 VSS.n7036 0.04025
R16470 VSS.n7036 VSS.n2221 0.04025
R16471 VSS.n7032 VSS.n2221 0.04025
R16472 VSS.n7032 VSS.n7031 0.04025
R16473 VSS.n7031 VSS.n7030 0.04025
R16474 VSS.n7030 VSS.n2223 0.04025
R16475 VSS.n7026 VSS.n2223 0.04025
R16476 VSS.n7026 VSS.n7025 0.04025
R16477 VSS.n7025 VSS.n7024 0.04025
R16478 VSS.n7024 VSS.n2225 0.04025
R16479 VSS.n7020 VSS.n2225 0.04025
R16480 VSS.n7020 VSS.n7019 0.04025
R16481 VSS.n7019 VSS.n7018 0.04025
R16482 VSS.n7018 VSS.n2227 0.04025
R16483 VSS.n7014 VSS.n2227 0.04025
R16484 VSS.n7014 VSS.n7013 0.04025
R16485 VSS.n7013 VSS.n7012 0.04025
R16486 VSS.n7012 VSS.n2229 0.04025
R16487 VSS.n7008 VSS.n2229 0.04025
R16488 VSS.n7008 VSS.n7007 0.04025
R16489 VSS.n7007 VSS.n7006 0.04025
R16490 VSS.n7006 VSS.n2231 0.04025
R16491 VSS.n7002 VSS.n2231 0.04025
R16492 VSS.n7002 VSS.n7001 0.04025
R16493 VSS.n7001 VSS.n7000 0.04025
R16494 VSS.n7000 VSS.n2233 0.04025
R16495 VSS.n6996 VSS.n2233 0.04025
R16496 VSS.n6996 VSS.n6995 0.04025
R16497 VSS.n6995 VSS.n6994 0.04025
R16498 VSS.n6994 VSS.n2235 0.04025
R16499 VSS.n6990 VSS.n2235 0.04025
R16500 VSS.n6990 VSS.n6989 0.04025
R16501 VSS.n6989 VSS.n6988 0.04025
R16502 VSS.n6988 VSS.n2237 0.04025
R16503 VSS.n6984 VSS.n2237 0.04025
R16504 VSS.n6984 VSS.n6983 0.04025
R16505 VSS.n6983 VSS.n6982 0.04025
R16506 VSS.n6982 VSS.n2239 0.04025
R16507 VSS.n6978 VSS.n2239 0.04025
R16508 VSS.n6978 VSS.n6977 0.04025
R16509 VSS.n6977 VSS.n6976 0.04025
R16510 VSS.n6976 VSS.n2241 0.04025
R16511 VSS.n6972 VSS.n2241 0.04025
R16512 VSS.n6972 VSS.n6971 0.04025
R16513 VSS.n6971 VSS.n6970 0.04025
R16514 VSS.n6970 VSS.n2243 0.04025
R16515 VSS.n6966 VSS.n2243 0.04025
R16516 VSS.n6966 VSS.n6965 0.04025
R16517 VSS.n6965 VSS.n6964 0.04025
R16518 VSS.n6964 VSS.n2245 0.04025
R16519 VSS.n6960 VSS.n2245 0.04025
R16520 VSS.n6960 VSS.n6959 0.04025
R16521 VSS.n6959 VSS.n6958 0.04025
R16522 VSS.n6958 VSS.n2247 0.04025
R16523 VSS.n6954 VSS.n2247 0.04025
R16524 VSS.n6954 VSS.n6953 0.04025
R16525 VSS.n6953 VSS.n6952 0.04025
R16526 VSS.n6952 VSS.n2249 0.04025
R16527 VSS.n6948 VSS.n2249 0.04025
R16528 VSS.n6948 VSS.n6947 0.04025
R16529 VSS.n6947 VSS.n6946 0.04025
R16530 VSS.n6946 VSS.n2251 0.04025
R16531 VSS.n6942 VSS.n2251 0.04025
R16532 VSS.n6942 VSS.n6941 0.04025
R16533 VSS.n6941 VSS.n6940 0.04025
R16534 VSS.n6940 VSS.n2253 0.04025
R16535 VSS.n6936 VSS.n6935 0.04025
R16536 VSS.n6935 VSS.n6934 0.04025
R16537 VSS.n6934 VSS.n2255 0.04025
R16538 VSS.n6930 VSS.n2255 0.04025
R16539 VSS.n6930 VSS.n6929 0.04025
R16540 VSS.n6929 VSS.n6928 0.04025
R16541 VSS.n6928 VSS.n2257 0.04025
R16542 VSS.n6924 VSS.n2257 0.04025
R16543 VSS.n6924 VSS.n6923 0.04025
R16544 VSS.n6923 VSS.n6922 0.04025
R16545 VSS.n6922 VSS.n2259 0.04025
R16546 VSS.n6918 VSS.n2259 0.04025
R16547 VSS.n6918 VSS.n6917 0.04025
R16548 VSS.n6917 VSS.n6916 0.04025
R16549 VSS.n6916 VSS.n2261 0.04025
R16550 VSS.n6912 VSS.n2261 0.04025
R16551 VSS.n6912 VSS.n6911 0.04025
R16552 VSS.n6911 VSS.n6910 0.04025
R16553 VSS.n6910 VSS.n2263 0.04025
R16554 VSS.n4141 VSS.n3185 0.04025
R16555 VSS.n4137 VSS.n3185 0.04025
R16556 VSS.n4137 VSS.n4136 0.04025
R16557 VSS.n4136 VSS.n4135 0.04025
R16558 VSS.n4135 VSS.n3187 0.04025
R16559 VSS.n4131 VSS.n3187 0.04025
R16560 VSS.n4131 VSS.n4130 0.04025
R16561 VSS.n4130 VSS.n4129 0.04025
R16562 VSS.n4129 VSS.n3189 0.04025
R16563 VSS.n4125 VSS.n3189 0.04025
R16564 VSS.n4125 VSS.n4124 0.04025
R16565 VSS.n4124 VSS.n4123 0.04025
R16566 VSS.n4123 VSS.n3191 0.04025
R16567 VSS.n4119 VSS.n3191 0.04025
R16568 VSS.n4119 VSS.n4118 0.04025
R16569 VSS.n4118 VSS.n4117 0.04025
R16570 VSS.n4117 VSS.n3193 0.04025
R16571 VSS.n4113 VSS.n3193 0.04025
R16572 VSS.n4113 VSS.n4112 0.04025
R16573 VSS.n4112 VSS.n4111 0.04025
R16574 VSS.n4111 VSS.n3195 0.04025
R16575 VSS.n4107 VSS.n3195 0.04025
R16576 VSS.n4107 VSS.n4106 0.04025
R16577 VSS.n4106 VSS.n4105 0.04025
R16578 VSS.n4105 VSS.n3197 0.04025
R16579 VSS.n4101 VSS.n3197 0.04025
R16580 VSS.n4101 VSS.n4100 0.04025
R16581 VSS.n4100 VSS.n4099 0.04025
R16582 VSS.n4099 VSS.n3199 0.04025
R16583 VSS.n4095 VSS.n3199 0.04025
R16584 VSS.n4095 VSS.n4094 0.04025
R16585 VSS.n4094 VSS.n4093 0.04025
R16586 VSS.n4093 VSS.n3201 0.04025
R16587 VSS.n4089 VSS.n3201 0.04025
R16588 VSS.n4089 VSS.n4088 0.04025
R16589 VSS.n4088 VSS.n4087 0.04025
R16590 VSS.n4087 VSS.n3203 0.04025
R16591 VSS.n4083 VSS.n3203 0.04025
R16592 VSS.n4083 VSS.n4082 0.04025
R16593 VSS.n4082 VSS.n4081 0.04025
R16594 VSS.n4081 VSS.n3205 0.04025
R16595 VSS.n4077 VSS.n3205 0.04025
R16596 VSS.n4077 VSS.n4076 0.04025
R16597 VSS.n4076 VSS.n4075 0.04025
R16598 VSS.n4075 VSS.n3207 0.04025
R16599 VSS.n4071 VSS.n3207 0.04025
R16600 VSS.n4071 VSS.n4070 0.04025
R16601 VSS.n4070 VSS.n4069 0.04025
R16602 VSS.n4069 VSS.n3209 0.04025
R16603 VSS.n4065 VSS.n3209 0.04025
R16604 VSS.n4065 VSS.n4064 0.04025
R16605 VSS.n4064 VSS.n4063 0.04025
R16606 VSS.n4063 VSS.n3211 0.04025
R16607 VSS.n4059 VSS.n3211 0.04025
R16608 VSS.n4059 VSS.n4058 0.04025
R16609 VSS.n4058 VSS.n4057 0.04025
R16610 VSS.n4057 VSS.n3213 0.04025
R16611 VSS.n4053 VSS.n3213 0.04025
R16612 VSS.n4053 VSS.n4052 0.04025
R16613 VSS.n4052 VSS.n4051 0.04025
R16614 VSS.n4051 VSS.n3215 0.04025
R16615 VSS.n4047 VSS.n3215 0.04025
R16616 VSS.n4047 VSS.n4046 0.04025
R16617 VSS.n4046 VSS.n4045 0.04025
R16618 VSS.n4045 VSS.n3217 0.04025
R16619 VSS.n4041 VSS.n3217 0.04025
R16620 VSS.n4041 VSS.n4040 0.04025
R16621 VSS.n4040 VSS.n4039 0.04025
R16622 VSS.n4039 VSS.n3219 0.04025
R16623 VSS.n4035 VSS.n3219 0.04025
R16624 VSS.n4035 VSS.n4034 0.04025
R16625 VSS.n4034 VSS.n4033 0.04025
R16626 VSS.n4033 VSS.n3221 0.04025
R16627 VSS.n4029 VSS.n3221 0.04025
R16628 VSS.n4029 VSS.n4028 0.04025
R16629 VSS.n4028 VSS.n4027 0.04025
R16630 VSS.n4027 VSS.n3223 0.04025
R16631 VSS.n4023 VSS.n3223 0.04025
R16632 VSS.n4023 VSS.n4022 0.04025
R16633 VSS.n4022 VSS.n4021 0.04025
R16634 VSS.n4021 VSS.n3225 0.04025
R16635 VSS.n4017 VSS.n3225 0.04025
R16636 VSS.n4017 VSS.n4016 0.04025
R16637 VSS.n4016 VSS.n4015 0.04025
R16638 VSS.n4015 VSS.n3227 0.04025
R16639 VSS.n4011 VSS.n3227 0.04025
R16640 VSS.n4011 VSS.n4010 0.04025
R16641 VSS.n4010 VSS.n4009 0.04025
R16642 VSS.n4009 VSS.n3229 0.04025
R16643 VSS.n4005 VSS.n3229 0.04025
R16644 VSS.n4005 VSS.n4004 0.04025
R16645 VSS.n4004 VSS.n4003 0.04025
R16646 VSS.n4003 VSS.n3231 0.04025
R16647 VSS.n3999 VSS.n3231 0.04025
R16648 VSS.n3999 VSS.n3998 0.04025
R16649 VSS.n3998 VSS.n3997 0.04025
R16650 VSS.n3997 VSS.n3233 0.04025
R16651 VSS.n3993 VSS.n3233 0.04025
R16652 VSS.n3993 VSS.n3992 0.04025
R16653 VSS.n3992 VSS.n3991 0.04025
R16654 VSS.n3991 VSS.n3235 0.04025
R16655 VSS.n3987 VSS.n3235 0.04025
R16656 VSS.n3987 VSS.n3986 0.04025
R16657 VSS.n3986 VSS.n3985 0.04025
R16658 VSS.n3985 VSS.n3237 0.04025
R16659 VSS.n3981 VSS.n3237 0.04025
R16660 VSS.n3981 VSS.n3980 0.04025
R16661 VSS.n3980 VSS.n3979 0.04025
R16662 VSS.n3979 VSS.n3239 0.04025
R16663 VSS.n3975 VSS.n3239 0.04025
R16664 VSS.n3975 VSS.n3974 0.04025
R16665 VSS.n3974 VSS.n3973 0.04025
R16666 VSS.n3973 VSS.n3241 0.04025
R16667 VSS.n3969 VSS.n3241 0.04025
R16668 VSS.n3969 VSS.n3968 0.04025
R16669 VSS.n3968 VSS.n3967 0.04025
R16670 VSS.n3967 VSS.n3243 0.04025
R16671 VSS.n3963 VSS.n3243 0.04025
R16672 VSS.n3963 VSS.n3962 0.04025
R16673 VSS.n3962 VSS.n3961 0.04025
R16674 VSS.n3961 VSS.n3245 0.04025
R16675 VSS.n3957 VSS.n3245 0.04025
R16676 VSS.n3957 VSS.n3956 0.04025
R16677 VSS.n3956 VSS.n3955 0.04025
R16678 VSS.n3955 VSS.n3247 0.04025
R16679 VSS.n3951 VSS.n3247 0.04025
R16680 VSS.n3951 VSS.n3950 0.04025
R16681 VSS.n3950 VSS.n3949 0.04025
R16682 VSS.n3949 VSS.n3249 0.04025
R16683 VSS.n3945 VSS.n3249 0.04025
R16684 VSS.n3945 VSS.n3944 0.04025
R16685 VSS.n3944 VSS.n3943 0.04025
R16686 VSS.n3943 VSS.n3251 0.04025
R16687 VSS.n3939 VSS.n3251 0.04025
R16688 VSS.n3939 VSS.n3938 0.04025
R16689 VSS.n3938 VSS.n3937 0.04025
R16690 VSS.n3937 VSS.n3253 0.04025
R16691 VSS.n3933 VSS.n3253 0.04025
R16692 VSS.n3933 VSS.n3932 0.04025
R16693 VSS.n3932 VSS.n3931 0.04025
R16694 VSS.n3931 VSS.n3255 0.04025
R16695 VSS.n3927 VSS.n3255 0.04025
R16696 VSS.n3927 VSS.n3926 0.04025
R16697 VSS.n3926 VSS.n3925 0.04025
R16698 VSS.n3925 VSS.n3257 0.04025
R16699 VSS.n3921 VSS.n3257 0.04025
R16700 VSS.n3921 VSS.n3920 0.04025
R16701 VSS.n3920 VSS.n3919 0.04025
R16702 VSS.n3919 VSS.n3259 0.04025
R16703 VSS.n3915 VSS.n3259 0.04025
R16704 VSS.n3915 VSS.n3914 0.04025
R16705 VSS.n3914 VSS.n3913 0.04025
R16706 VSS.n3913 VSS.n3261 0.04025
R16707 VSS.n3909 VSS.n3261 0.04025
R16708 VSS.n3909 VSS.n3908 0.04025
R16709 VSS.n3908 VSS.n3907 0.04025
R16710 VSS.n3907 VSS.n3263 0.04025
R16711 VSS.n3903 VSS.n3263 0.04025
R16712 VSS.n3903 VSS.n3902 0.04025
R16713 VSS.n3902 VSS.n3901 0.04025
R16714 VSS.n3901 VSS.n3265 0.04025
R16715 VSS.n3897 VSS.n3265 0.04025
R16716 VSS.n3897 VSS.n3896 0.04025
R16717 VSS.n3896 VSS.n3895 0.04025
R16718 VSS.n3895 VSS.n3267 0.04025
R16719 VSS.n3891 VSS.n3267 0.04025
R16720 VSS.n3891 VSS.n3890 0.04025
R16721 VSS.n3890 VSS.n3889 0.04025
R16722 VSS.n3889 VSS.n3269 0.04025
R16723 VSS.n3885 VSS.n3269 0.04025
R16724 VSS.n3885 VSS.n3884 0.04025
R16725 VSS.n3884 VSS.n3883 0.04025
R16726 VSS.n3883 VSS.n3271 0.04025
R16727 VSS.n3879 VSS.n3271 0.04025
R16728 VSS.n3879 VSS.n3878 0.04025
R16729 VSS.n3878 VSS.n3877 0.04025
R16730 VSS.n3877 VSS.n3273 0.04025
R16731 VSS.n3873 VSS.n3273 0.04025
R16732 VSS.n3873 VSS.n3872 0.04025
R16733 VSS.n3872 VSS.n3871 0.04025
R16734 VSS.n3871 VSS.n3275 0.04025
R16735 VSS.n3867 VSS.n3275 0.04025
R16736 VSS.n3867 VSS.n3866 0.04025
R16737 VSS.n3866 VSS.n3865 0.04025
R16738 VSS.n3865 VSS.n3277 0.04025
R16739 VSS.n3861 VSS.n3277 0.04025
R16740 VSS.n3861 VSS.n3860 0.04025
R16741 VSS.n3860 VSS.n3859 0.04025
R16742 VSS.n3859 VSS.n3279 0.04025
R16743 VSS.n3855 VSS.n3279 0.04025
R16744 VSS.n3855 VSS.n3854 0.04025
R16745 VSS.n3854 VSS.n3853 0.04025
R16746 VSS.n3853 VSS.n3281 0.04025
R16747 VSS.n3849 VSS.n3281 0.04025
R16748 VSS.n3849 VSS.n3848 0.04025
R16749 VSS.n3848 VSS.n3847 0.04025
R16750 VSS.n3847 VSS.n3283 0.04025
R16751 VSS.n3843 VSS.n3283 0.04025
R16752 VSS.n3843 VSS.n3842 0.04025
R16753 VSS.n3842 VSS.n3841 0.04025
R16754 VSS.n3841 VSS.n3285 0.04025
R16755 VSS.n3837 VSS.n3285 0.04025
R16756 VSS.n3837 VSS.n3836 0.04025
R16757 VSS.n3836 VSS.n3835 0.04025
R16758 VSS.n3835 VSS.n3287 0.04025
R16759 VSS.n3831 VSS.n3287 0.04025
R16760 VSS.n3831 VSS.n3830 0.04025
R16761 VSS.n3830 VSS.n3829 0.04025
R16762 VSS.n3829 VSS.n3289 0.04025
R16763 VSS.n3825 VSS.n3289 0.04025
R16764 VSS.n3825 VSS.n3824 0.04025
R16765 VSS.n3824 VSS.n3823 0.04025
R16766 VSS.n3823 VSS.n3291 0.04025
R16767 VSS.n3819 VSS.n3291 0.04025
R16768 VSS.n3819 VSS.n3818 0.04025
R16769 VSS.n3818 VSS.n3817 0.04025
R16770 VSS.n3817 VSS.n3293 0.04025
R16771 VSS.n3813 VSS.n3293 0.04025
R16772 VSS.n3813 VSS.n3812 0.04025
R16773 VSS.n3812 VSS.n3811 0.04025
R16774 VSS.n3811 VSS.n3295 0.04025
R16775 VSS.n3807 VSS.n3295 0.04025
R16776 VSS.n3807 VSS.n3806 0.04025
R16777 VSS.n3806 VSS.n3805 0.04025
R16778 VSS.n3805 VSS.n3297 0.04025
R16779 VSS.n3801 VSS.n3297 0.04025
R16780 VSS.n3801 VSS.n3800 0.04025
R16781 VSS.n3800 VSS.n3799 0.04025
R16782 VSS.n3799 VSS.n3299 0.04025
R16783 VSS.n3795 VSS.n3299 0.04025
R16784 VSS.n3795 VSS.n3794 0.04025
R16785 VSS.n3794 VSS.n3793 0.04025
R16786 VSS.n3793 VSS.n3301 0.04025
R16787 VSS.n3789 VSS.n3301 0.04025
R16788 VSS.n3789 VSS.n3788 0.04025
R16789 VSS.n3788 VSS.n3787 0.04025
R16790 VSS.n3787 VSS.n3303 0.04025
R16791 VSS.n3783 VSS.n3303 0.04025
R16792 VSS.n3783 VSS.n3782 0.04025
R16793 VSS.n3782 VSS.n3781 0.04025
R16794 VSS.n3781 VSS.n3305 0.04025
R16795 VSS.n3777 VSS.n3305 0.04025
R16796 VSS.n3777 VSS.n3776 0.04025
R16797 VSS.n3776 VSS.n3775 0.04025
R16798 VSS.n3775 VSS.n3307 0.04025
R16799 VSS.n3771 VSS.n3307 0.04025
R16800 VSS.n3771 VSS.n3770 0.04025
R16801 VSS.n3770 VSS.n3769 0.04025
R16802 VSS.n3769 VSS.n3309 0.04025
R16803 VSS.n3765 VSS.n3309 0.04025
R16804 VSS.n3765 VSS.n3764 0.04025
R16805 VSS.n3764 VSS.n3763 0.04025
R16806 VSS.n3763 VSS.n3311 0.04025
R16807 VSS.n3759 VSS.n3311 0.04025
R16808 VSS.n3759 VSS.n3758 0.04025
R16809 VSS.n3758 VSS.n3757 0.04025
R16810 VSS.n3757 VSS.n3313 0.04025
R16811 VSS.n3753 VSS.n3313 0.04025
R16812 VSS.n3753 VSS.n3752 0.04025
R16813 VSS.n3752 VSS.n3751 0.04025
R16814 VSS.n3751 VSS.n3315 0.04025
R16815 VSS.n3747 VSS.n3315 0.04025
R16816 VSS.n3747 VSS.n3746 0.04025
R16817 VSS.n3746 VSS.n3745 0.04025
R16818 VSS.n3745 VSS.n3317 0.04025
R16819 VSS.n3741 VSS.n3317 0.04025
R16820 VSS.n3741 VSS.n3740 0.04025
R16821 VSS.n3740 VSS.n3739 0.04025
R16822 VSS.n3739 VSS.n3319 0.04025
R16823 VSS.n3735 VSS.n3319 0.04025
R16824 VSS.n3735 VSS.n3734 0.04025
R16825 VSS.n3734 VSS.n3733 0.04025
R16826 VSS.n3733 VSS.n3321 0.04025
R16827 VSS.n3729 VSS.n3321 0.04025
R16828 VSS.n3729 VSS.n3728 0.04025
R16829 VSS.n3728 VSS.n3727 0.04025
R16830 VSS.n3727 VSS.n3323 0.04025
R16831 VSS.n3723 VSS.n3323 0.04025
R16832 VSS.n3723 VSS.n3722 0.04025
R16833 VSS.n3722 VSS.n3721 0.04025
R16834 VSS.n3721 VSS.n3325 0.04025
R16835 VSS.n3717 VSS.n3325 0.04025
R16836 VSS.n3717 VSS.n3716 0.04025
R16837 VSS.n3716 VSS.n3715 0.04025
R16838 VSS.n3715 VSS.n3327 0.04025
R16839 VSS.n3711 VSS.n3327 0.04025
R16840 VSS.n3711 VSS.n3710 0.04025
R16841 VSS.n3710 VSS.n3709 0.04025
R16842 VSS.n3709 VSS.n3329 0.04025
R16843 VSS.n3705 VSS.n3329 0.04025
R16844 VSS.n3705 VSS.n3704 0.04025
R16845 VSS.n3704 VSS.n3703 0.04025
R16846 VSS.n3703 VSS.n3331 0.04025
R16847 VSS.n3699 VSS.n3331 0.04025
R16848 VSS.n3699 VSS.n3698 0.04025
R16849 VSS.n3698 VSS.n3697 0.04025
R16850 VSS.n3697 VSS.n3333 0.04025
R16851 VSS.n3693 VSS.n3333 0.04025
R16852 VSS.n3693 VSS.n3692 0.04025
R16853 VSS.n3692 VSS.n3691 0.04025
R16854 VSS.n3691 VSS.n3335 0.04025
R16855 VSS.n3687 VSS.n3335 0.04025
R16856 VSS.n3687 VSS.n3686 0.04025
R16857 VSS.n3686 VSS.n3685 0.04025
R16858 VSS.n3685 VSS.n3337 0.04025
R16859 VSS.n3681 VSS.n3337 0.04025
R16860 VSS.n3681 VSS.n3680 0.04025
R16861 VSS.n3680 VSS.n3679 0.04025
R16862 VSS.n3679 VSS.n3339 0.04025
R16863 VSS.n3675 VSS.n3339 0.04025
R16864 VSS.n3675 VSS.n3674 0.04025
R16865 VSS.n3674 VSS.n3673 0.04025
R16866 VSS.n3673 VSS.n3341 0.04025
R16867 VSS.n3669 VSS.n3341 0.04025
R16868 VSS.n3669 VSS.n3668 0.04025
R16869 VSS.n3668 VSS.n3667 0.04025
R16870 VSS.n3667 VSS.n3343 0.04025
R16871 VSS.n3663 VSS.n3343 0.04025
R16872 VSS.n3663 VSS.n3662 0.04025
R16873 VSS.n3662 VSS.n3661 0.04025
R16874 VSS.n3661 VSS.n3345 0.04025
R16875 VSS.n3657 VSS.n3345 0.04025
R16876 VSS.n3657 VSS.n3656 0.04025
R16877 VSS.n3656 VSS.n3655 0.04025
R16878 VSS.n3655 VSS.n3347 0.04025
R16879 VSS.n3651 VSS.n3347 0.04025
R16880 VSS.n3651 VSS.n3650 0.04025
R16881 VSS.n3650 VSS.n3649 0.04025
R16882 VSS.n3649 VSS.n3349 0.04025
R16883 VSS.n3645 VSS.n3349 0.04025
R16884 VSS.n3645 VSS.n3644 0.04025
R16885 VSS.n3644 VSS.n3643 0.04025
R16886 VSS.n3643 VSS.n3351 0.04025
R16887 VSS.n3639 VSS.n3351 0.04025
R16888 VSS.n3639 VSS.n3638 0.04025
R16889 VSS.n3638 VSS.n3637 0.04025
R16890 VSS.n3637 VSS.n3353 0.04025
R16891 VSS.n3633 VSS.n3353 0.04025
R16892 VSS.n3633 VSS.n3632 0.04025
R16893 VSS.n3632 VSS.n3631 0.04025
R16894 VSS.n3631 VSS.n3355 0.04025
R16895 VSS.n3627 VSS.n3355 0.04025
R16896 VSS.n3627 VSS.n3626 0.04025
R16897 VSS.n3626 VSS.n3625 0.04025
R16898 VSS.n3625 VSS.n3357 0.04025
R16899 VSS.n3621 VSS.n3357 0.04025
R16900 VSS.n3621 VSS.n3620 0.04025
R16901 VSS.n3620 VSS.n3619 0.04025
R16902 VSS.n3619 VSS.n3359 0.04025
R16903 VSS.n3615 VSS.n3359 0.04025
R16904 VSS.n3615 VSS.n3614 0.04025
R16905 VSS.n3614 VSS.n3613 0.04025
R16906 VSS.n3613 VSS.n3361 0.04025
R16907 VSS.n3609 VSS.n3361 0.04025
R16908 VSS.n3609 VSS.n3608 0.04025
R16909 VSS.n3608 VSS.n3607 0.04025
R16910 VSS.n3607 VSS.n3363 0.04025
R16911 VSS.n3603 VSS.n3363 0.04025
R16912 VSS.n3603 VSS.n3602 0.04025
R16913 VSS.n3602 VSS.n3601 0.04025
R16914 VSS.n3601 VSS.n3365 0.04025
R16915 VSS.n3597 VSS.n3365 0.04025
R16916 VSS.n3597 VSS.n3596 0.04025
R16917 VSS.n3596 VSS.n3595 0.04025
R16918 VSS.n3595 VSS.n3367 0.04025
R16919 VSS.n3591 VSS.n3367 0.04025
R16920 VSS.n3591 VSS.n3590 0.04025
R16921 VSS.n3590 VSS.n3589 0.04025
R16922 VSS.n3589 VSS.n3369 0.04025
R16923 VSS.n3585 VSS.n3369 0.04025
R16924 VSS.n3585 VSS.n3584 0.04025
R16925 VSS.n3584 VSS.n3583 0.04025
R16926 VSS.n3583 VSS.n3371 0.04025
R16927 VSS.n3579 VSS.n3371 0.04025
R16928 VSS.n3579 VSS.n3578 0.04025
R16929 VSS.n3578 VSS.n3577 0.04025
R16930 VSS.n3577 VSS.n3373 0.04025
R16931 VSS.n3573 VSS.n3373 0.04025
R16932 VSS.n3573 VSS.n3572 0.04025
R16933 VSS.n3572 VSS.n3571 0.04025
R16934 VSS.n3571 VSS.n3375 0.04025
R16935 VSS.n3567 VSS.n3375 0.04025
R16936 VSS.n3567 VSS.n3566 0.04025
R16937 VSS.n3566 VSS.n3565 0.04025
R16938 VSS.n3565 VSS.n3377 0.04025
R16939 VSS.n3561 VSS.n3377 0.04025
R16940 VSS.n3561 VSS.n3560 0.04025
R16941 VSS.n3560 VSS.n3559 0.04025
R16942 VSS.n3559 VSS.n3379 0.04025
R16943 VSS.n3555 VSS.n3379 0.04025
R16944 VSS.n3555 VSS.n3554 0.04025
R16945 VSS.n3554 VSS.n3553 0.04025
R16946 VSS.n3553 VSS.n3381 0.04025
R16947 VSS.n3549 VSS.n3381 0.04025
R16948 VSS.n3549 VSS.n3548 0.04025
R16949 VSS.n3548 VSS.n3547 0.04025
R16950 VSS.n3547 VSS.n3383 0.04025
R16951 VSS.n3543 VSS.n3383 0.04025
R16952 VSS.n3543 VSS.n3542 0.04025
R16953 VSS.n3542 VSS.n3541 0.04025
R16954 VSS.n3541 VSS.n3385 0.04025
R16955 VSS.n3537 VSS.n3385 0.04025
R16956 VSS.n3537 VSS.n3536 0.04025
R16957 VSS.n3536 VSS.n3535 0.04025
R16958 VSS.n3535 VSS.n3387 0.04025
R16959 VSS.n3531 VSS.n3387 0.04025
R16960 VSS.n3531 VSS.n3530 0.04025
R16961 VSS.n3530 VSS.n3529 0.04025
R16962 VSS.n3529 VSS.n3389 0.04025
R16963 VSS.n3525 VSS.n3389 0.04025
R16964 VSS.n3525 VSS.n3524 0.04025
R16965 VSS.n3524 VSS.n3523 0.04025
R16966 VSS.n3523 VSS.n3391 0.04025
R16967 VSS.n3519 VSS.n3391 0.04025
R16968 VSS.n3519 VSS.n3518 0.04025
R16969 VSS.n3518 VSS.n3517 0.04025
R16970 VSS.n3517 VSS.n3393 0.04025
R16971 VSS.n3513 VSS.n3393 0.04025
R16972 VSS.n3513 VSS.n3512 0.04025
R16973 VSS.n3512 VSS.n3511 0.04025
R16974 VSS.n3511 VSS.n3395 0.04025
R16975 VSS.n3507 VSS.n3395 0.04025
R16976 VSS.n3507 VSS.n3506 0.04025
R16977 VSS.n3506 VSS.n3505 0.04025
R16978 VSS.n3505 VSS.n3397 0.04025
R16979 VSS.n3501 VSS.n3397 0.04025
R16980 VSS.n3501 VSS.n3500 0.04025
R16981 VSS.n3500 VSS.n3499 0.04025
R16982 VSS.n3499 VSS.n3399 0.04025
R16983 VSS.n3495 VSS.n3399 0.04025
R16984 VSS.n3495 VSS.n3494 0.04025
R16985 VSS.n3494 VSS.n3493 0.04025
R16986 VSS.n3493 VSS.n3401 0.04025
R16987 VSS.n3489 VSS.n3401 0.04025
R16988 VSS.n3489 VSS.n3488 0.04025
R16989 VSS.n3488 VSS.n3487 0.04025
R16990 VSS.n3487 VSS.n3403 0.04025
R16991 VSS.n3483 VSS.n3403 0.04025
R16992 VSS.n3483 VSS.n3482 0.04025
R16993 VSS.n3482 VSS.n3481 0.04025
R16994 VSS.n3481 VSS.n3405 0.04025
R16995 VSS.n3477 VSS.n3405 0.04025
R16996 VSS.n3477 VSS.n3476 0.04025
R16997 VSS.n3476 VSS.n3475 0.04025
R16998 VSS.n3475 VSS.n3407 0.04025
R16999 VSS.n3471 VSS.n3407 0.04025
R17000 VSS.n3471 VSS.n3470 0.04025
R17001 VSS.n3470 VSS.n3469 0.04025
R17002 VSS.n3469 VSS.n3409 0.04025
R17003 VSS.n3465 VSS.n3409 0.04025
R17004 VSS.n3465 VSS.n3464 0.04025
R17005 VSS.n3464 VSS.n3463 0.04025
R17006 VSS.n3463 VSS.n3411 0.04025
R17007 VSS.n3459 VSS.n3411 0.04025
R17008 VSS.n3459 VSS.n3458 0.04025
R17009 VSS.n3458 VSS.n3457 0.04025
R17010 VSS.n3457 VSS.n3413 0.04025
R17011 VSS.n3453 VSS.n3413 0.04025
R17012 VSS.n3453 VSS.n3452 0.04025
R17013 VSS.n3452 VSS.n3451 0.04025
R17014 VSS.n3451 VSS.n3415 0.04025
R17015 VSS.n3447 VSS.n3415 0.04025
R17016 VSS.n3447 VSS.n3446 0.04025
R17017 VSS.n3446 VSS.n3445 0.04025
R17018 VSS.n3445 VSS.n3417 0.04025
R17019 VSS.n3441 VSS.n3417 0.04025
R17020 VSS.n3441 VSS.n3440 0.04025
R17021 VSS.n3440 VSS.n3439 0.04025
R17022 VSS.n3439 VSS.n3419 0.04025
R17023 VSS.n3435 VSS.n3419 0.04025
R17024 VSS.n3435 VSS.n3434 0.04025
R17025 VSS.n3434 VSS.n3433 0.04025
R17026 VSS.n3433 VSS.n3421 0.04025
R17027 VSS.n3429 VSS.n3421 0.04025
R17028 VSS.n3429 VSS.n3428 0.04025
R17029 VSS.n3428 VSS.n3427 0.04025
R17030 VSS.n3427 VSS.n3423 0.04025
R17031 VSS.n3423 VSS.n1581 0.04025
R17032 VSS.n8951 VSS.n1581 0.04025
R17033 VSS.n8951 VSS.n8950 0.04025
R17034 VSS.n8950 VSS.n1583 0.04025
R17035 VSS.n8946 VSS.n1583 0.04025
R17036 VSS.n8946 VSS.n8945 0.04025
R17037 VSS.n8945 VSS.n8944 0.04025
R17038 VSS.n8944 VSS.n1585 0.04025
R17039 VSS.n8940 VSS.n1585 0.04025
R17040 VSS.n8940 VSS.n8939 0.04025
R17041 VSS.n8939 VSS.n8938 0.04025
R17042 VSS.n8938 VSS.n1587 0.04025
R17043 VSS.n8934 VSS.n1587 0.04025
R17044 VSS.n8934 VSS.n8933 0.04025
R17045 VSS.n8933 VSS.n8932 0.04025
R17046 VSS.n8932 VSS.n1589 0.04025
R17047 VSS.n8928 VSS.n1589 0.04025
R17048 VSS.n8928 VSS.n8927 0.04025
R17049 VSS.n8927 VSS.n8926 0.04025
R17050 VSS.n8926 VSS.n1591 0.04025
R17051 VSS.n8922 VSS.n1591 0.04025
R17052 VSS.n8922 VSS.n8921 0.04025
R17053 VSS.n8921 VSS.n8920 0.04025
R17054 VSS.n8920 VSS.n1593 0.04025
R17055 VSS.n8916 VSS.n1593 0.04025
R17056 VSS.n8916 VSS.n8915 0.04025
R17057 VSS.n8915 VSS.n8914 0.04025
R17058 VSS.n8914 VSS.n1595 0.04025
R17059 VSS.n8910 VSS.n1595 0.04025
R17060 VSS.n8910 VSS.n8909 0.04025
R17061 VSS.n8909 VSS.n8908 0.04025
R17062 VSS.n8908 VSS.n1597 0.04025
R17063 VSS.n8904 VSS.n1597 0.04025
R17064 VSS.n8904 VSS.n8903 0.04025
R17065 VSS.n8903 VSS.n8902 0.04025
R17066 VSS.n8902 VSS.n1599 0.04025
R17067 VSS.n8898 VSS.n1599 0.04025
R17068 VSS.n8898 VSS.n8897 0.04025
R17069 VSS.n8897 VSS.n8896 0.04025
R17070 VSS.n8896 VSS.n1601 0.04025
R17071 VSS.n8892 VSS.n1601 0.04025
R17072 VSS.n8892 VSS.n8891 0.04025
R17073 VSS.n8891 VSS.n8890 0.04025
R17074 VSS.n8890 VSS.n1603 0.04025
R17075 VSS.n8886 VSS.n1603 0.04025
R17076 VSS.n8886 VSS.n8885 0.04025
R17077 VSS.n8885 VSS.n8884 0.04025
R17078 VSS.n8884 VSS.n1605 0.04025
R17079 VSS.n8880 VSS.n1605 0.04025
R17080 VSS.n8880 VSS.n8879 0.04025
R17081 VSS.n8879 VSS.n8878 0.04025
R17082 VSS.n8878 VSS.n1607 0.04025
R17083 VSS.n8874 VSS.n1607 0.04025
R17084 VSS.n8874 VSS.n8873 0.04025
R17085 VSS.n8873 VSS.n8872 0.04025
R17086 VSS.n8872 VSS.n1609 0.04025
R17087 VSS.n8868 VSS.n1609 0.04025
R17088 VSS.n8868 VSS.n8867 0.04025
R17089 VSS.n8867 VSS.n8866 0.04025
R17090 VSS.n8866 VSS.n1611 0.04025
R17091 VSS.n8862 VSS.n1611 0.04025
R17092 VSS.n8862 VSS.n8861 0.04025
R17093 VSS.n8861 VSS.n8860 0.04025
R17094 VSS.n8860 VSS.n1613 0.04025
R17095 VSS.n8856 VSS.n1613 0.04025
R17096 VSS.n8856 VSS.n8855 0.04025
R17097 VSS.n8855 VSS.n8854 0.04025
R17098 VSS.n8854 VSS.n1615 0.04025
R17099 VSS.n8850 VSS.n1615 0.04025
R17100 VSS.n8850 VSS.n8849 0.04025
R17101 VSS.n8849 VSS.n8848 0.04025
R17102 VSS.n8848 VSS.n1617 0.04025
R17103 VSS.n8844 VSS.n1617 0.04025
R17104 VSS.n8844 VSS.n8843 0.04025
R17105 VSS.n8843 VSS.n8842 0.04025
R17106 VSS.n8842 VSS.n1619 0.04025
R17107 VSS.n8838 VSS.n1619 0.04025
R17108 VSS.n8838 VSS.n8837 0.04025
R17109 VSS.n8837 VSS.n8836 0.04025
R17110 VSS.n8836 VSS.n1621 0.04025
R17111 VSS.n8832 VSS.n1621 0.04025
R17112 VSS.n8832 VSS.n8831 0.04025
R17113 VSS.n8831 VSS.n8830 0.04025
R17114 VSS.n8830 VSS.n1623 0.04025
R17115 VSS.n8826 VSS.n1623 0.04025
R17116 VSS.n8826 VSS.n8825 0.04025
R17117 VSS.n8825 VSS.n8824 0.04025
R17118 VSS.n8824 VSS.n1625 0.04025
R17119 VSS.n8820 VSS.n1625 0.04025
R17120 VSS.n8820 VSS.n8819 0.04025
R17121 VSS.n8819 VSS.n8818 0.04025
R17122 VSS.n8818 VSS.n1627 0.04025
R17123 VSS.n8814 VSS.n1627 0.04025
R17124 VSS.n8814 VSS.n8813 0.04025
R17125 VSS.n8813 VSS.n8812 0.04025
R17126 VSS.n8812 VSS.n1629 0.04025
R17127 VSS.n8808 VSS.n1629 0.04025
R17128 VSS.n8808 VSS.n8807 0.04025
R17129 VSS.n8807 VSS.n8806 0.04025
R17130 VSS.n8806 VSS.n1631 0.04025
R17131 VSS.n8802 VSS.n1631 0.04025
R17132 VSS.n8802 VSS.n8801 0.04025
R17133 VSS.n8801 VSS.n8800 0.04025
R17134 VSS.n8800 VSS.n1633 0.04025
R17135 VSS.n8796 VSS.n1633 0.04025
R17136 VSS.n8796 VSS.n8795 0.04025
R17137 VSS.n8795 VSS.n8794 0.04025
R17138 VSS.n8794 VSS.n1635 0.04025
R17139 VSS.n8790 VSS.n1635 0.04025
R17140 VSS.n8790 VSS.n8789 0.04025
R17141 VSS.n8789 VSS.n8788 0.04025
R17142 VSS.n8788 VSS.n1637 0.04025
R17143 VSS.n8784 VSS.n1637 0.04025
R17144 VSS.n8784 VSS.n8783 0.04025
R17145 VSS.n8783 VSS.n8782 0.04025
R17146 VSS.n8782 VSS.n1639 0.04025
R17147 VSS.n8778 VSS.n1639 0.04025
R17148 VSS.n8778 VSS.n8777 0.04025
R17149 VSS.n8777 VSS.n8776 0.04025
R17150 VSS.n8776 VSS.n1641 0.04025
R17151 VSS.n8772 VSS.n1641 0.04025
R17152 VSS.n8772 VSS.n8771 0.04025
R17153 VSS.n8771 VSS.n8770 0.04025
R17154 VSS.n8770 VSS.n1643 0.04025
R17155 VSS.n8766 VSS.n1643 0.04025
R17156 VSS.n8766 VSS.n8765 0.04025
R17157 VSS.n8765 VSS.n8764 0.04025
R17158 VSS.n8764 VSS.n1645 0.04025
R17159 VSS.n8760 VSS.n1645 0.04025
R17160 VSS.n8760 VSS.n8759 0.04025
R17161 VSS.n8759 VSS.n8758 0.04025
R17162 VSS.n8758 VSS.n1647 0.04025
R17163 VSS.n8754 VSS.n1647 0.04025
R17164 VSS.n8754 VSS.n8753 0.04025
R17165 VSS.n8753 VSS.n8752 0.04025
R17166 VSS.n8752 VSS.n1649 0.04025
R17167 VSS.n8748 VSS.n1649 0.04025
R17168 VSS.n8748 VSS.n8747 0.04025
R17169 VSS.n8747 VSS.n8746 0.04025
R17170 VSS.n8746 VSS.n1651 0.04025
R17171 VSS.n8742 VSS.n1651 0.04025
R17172 VSS.n8742 VSS.n8741 0.04025
R17173 VSS.n8741 VSS.n8740 0.04025
R17174 VSS.n8740 VSS.n1653 0.04025
R17175 VSS.n8736 VSS.n1653 0.04025
R17176 VSS.n8736 VSS.n8735 0.04025
R17177 VSS.n8735 VSS.n8734 0.04025
R17178 VSS.n8734 VSS.n1655 0.04025
R17179 VSS.n8730 VSS.n1655 0.04025
R17180 VSS.n8730 VSS.n8729 0.04025
R17181 VSS.n8729 VSS.n8728 0.04025
R17182 VSS.n8728 VSS.n1657 0.04025
R17183 VSS.n8724 VSS.n1657 0.04025
R17184 VSS.n8724 VSS.n8723 0.04025
R17185 VSS.n8723 VSS.n8722 0.04025
R17186 VSS.n8722 VSS.n1659 0.04025
R17187 VSS.n8718 VSS.n1659 0.04025
R17188 VSS.n8718 VSS.n8717 0.04025
R17189 VSS.n8717 VSS.n8716 0.04025
R17190 VSS.n8716 VSS.n1661 0.04025
R17191 VSS.n8712 VSS.n1661 0.04025
R17192 VSS.n8712 VSS.n8711 0.04025
R17193 VSS.n8711 VSS.n8710 0.04025
R17194 VSS.n8710 VSS.n1663 0.04025
R17195 VSS.n8706 VSS.n1663 0.04025
R17196 VSS.n8706 VSS.n8705 0.04025
R17197 VSS.n8705 VSS.n8704 0.04025
R17198 VSS.n8704 VSS.n1665 0.04025
R17199 VSS.n8700 VSS.n1665 0.04025
R17200 VSS.n8700 VSS.n8699 0.04025
R17201 VSS.n8699 VSS.n8698 0.04025
R17202 VSS.n8698 VSS.n1667 0.04025
R17203 VSS.n8694 VSS.n1667 0.04025
R17204 VSS.n8694 VSS.n8693 0.04025
R17205 VSS.n8693 VSS.n8692 0.04025
R17206 VSS.n8692 VSS.n1669 0.04025
R17207 VSS.n8688 VSS.n1669 0.04025
R17208 VSS.n8688 VSS.n8687 0.04025
R17209 VSS.n8687 VSS.n8686 0.04025
R17210 VSS.n8686 VSS.n1671 0.04025
R17211 VSS.n8682 VSS.n1671 0.04025
R17212 VSS.n8682 VSS.n8681 0.04025
R17213 VSS.n8681 VSS.n8680 0.04025
R17214 VSS.n8680 VSS.n1673 0.04025
R17215 VSS.n8676 VSS.n1673 0.04025
R17216 VSS.n8676 VSS.n8675 0.04025
R17217 VSS.n8675 VSS.n8674 0.04025
R17218 VSS.n8674 VSS.n1675 0.04025
R17219 VSS.n8670 VSS.n1675 0.04025
R17220 VSS.n8670 VSS.n8669 0.04025
R17221 VSS.n8669 VSS.n8668 0.04025
R17222 VSS.n8668 VSS.n1677 0.04025
R17223 VSS.n8664 VSS.n1677 0.04025
R17224 VSS.n8664 VSS.n8663 0.04025
R17225 VSS.n8663 VSS.n8662 0.04025
R17226 VSS.n8662 VSS.n1679 0.04025
R17227 VSS.n8658 VSS.n1679 0.04025
R17228 VSS.n8658 VSS.n8657 0.04025
R17229 VSS.n8657 VSS.n8656 0.04025
R17230 VSS.n8656 VSS.n1681 0.04025
R17231 VSS.n8652 VSS.n1681 0.04025
R17232 VSS.n8652 VSS.n8651 0.04025
R17233 VSS.n8651 VSS.n8650 0.04025
R17234 VSS.n8650 VSS.n1683 0.04025
R17235 VSS.n8646 VSS.n1683 0.04025
R17236 VSS.n8646 VSS.n8645 0.04025
R17237 VSS.n8645 VSS.n8644 0.04025
R17238 VSS.n8644 VSS.n1685 0.04025
R17239 VSS.n8640 VSS.n1685 0.04025
R17240 VSS.n8640 VSS.n8639 0.04025
R17241 VSS.n8639 VSS.n8638 0.04025
R17242 VSS.n8638 VSS.n1687 0.04025
R17243 VSS.n8634 VSS.n1687 0.04025
R17244 VSS.n8634 VSS.n8633 0.04025
R17245 VSS.n8633 VSS.n8632 0.04025
R17246 VSS.n8632 VSS.n1689 0.04025
R17247 VSS.n8628 VSS.n1689 0.04025
R17248 VSS.n8628 VSS.n8627 0.04025
R17249 VSS.n8627 VSS.n8626 0.04025
R17250 VSS.n8626 VSS.n1691 0.04025
R17251 VSS.n8622 VSS.n1691 0.04025
R17252 VSS.n8622 VSS.n8621 0.04025
R17253 VSS.n8621 VSS.n8620 0.04025
R17254 VSS.n8620 VSS.n1693 0.04025
R17255 VSS.n8616 VSS.n1693 0.04025
R17256 VSS.n8616 VSS.n8615 0.04025
R17257 VSS.n8615 VSS.n8614 0.04025
R17258 VSS.n8614 VSS.n1695 0.04025
R17259 VSS.n8610 VSS.n1695 0.04025
R17260 VSS.n8610 VSS.n8609 0.04025
R17261 VSS.n8609 VSS.n8608 0.04025
R17262 VSS.n8608 VSS.n1697 0.04025
R17263 VSS.n8604 VSS.n1697 0.04025
R17264 VSS.n8604 VSS.n8603 0.04025
R17265 VSS.n8603 VSS.n8602 0.04025
R17266 VSS.n8602 VSS.n1699 0.04025
R17267 VSS.n8598 VSS.n1699 0.04025
R17268 VSS.n8598 VSS.n8597 0.04025
R17269 VSS.n8597 VSS.n8596 0.04025
R17270 VSS.n8596 VSS.n1701 0.04025
R17271 VSS.n8592 VSS.n1701 0.04025
R17272 VSS.n8592 VSS.n8591 0.04025
R17273 VSS.n8591 VSS.n8590 0.04025
R17274 VSS.n8590 VSS.n1703 0.04025
R17275 VSS.n8586 VSS.n1703 0.04025
R17276 VSS.n8586 VSS.n8585 0.04025
R17277 VSS.n8585 VSS.n8584 0.04025
R17278 VSS.n8584 VSS.n1705 0.04025
R17279 VSS.n8580 VSS.n1705 0.04025
R17280 VSS.n8580 VSS.n8579 0.04025
R17281 VSS.n8579 VSS.n8578 0.04025
R17282 VSS.n8578 VSS.n1707 0.04025
R17283 VSS.n8574 VSS.n1707 0.04025
R17284 VSS.n8574 VSS.n8573 0.04025
R17285 VSS.n8573 VSS.n8572 0.04025
R17286 VSS.n8572 VSS.n1709 0.04025
R17287 VSS.n8568 VSS.n1709 0.04025
R17288 VSS.n8568 VSS.n8567 0.04025
R17289 VSS.n8567 VSS.n8566 0.04025
R17290 VSS.n8566 VSS.n1711 0.04025
R17291 VSS.n8562 VSS.n1711 0.04025
R17292 VSS.n8562 VSS.n8561 0.04025
R17293 VSS.n8561 VSS.n8560 0.04025
R17294 VSS.n8560 VSS.n1713 0.04025
R17295 VSS.n8556 VSS.n1713 0.04025
R17296 VSS.n8556 VSS.n8555 0.04025
R17297 VSS.n8555 VSS.n8554 0.04025
R17298 VSS.n8554 VSS.n1715 0.04025
R17299 VSS.n8550 VSS.n1715 0.04025
R17300 VSS.n8550 VSS.n8549 0.04025
R17301 VSS.n8549 VSS.n8548 0.04025
R17302 VSS.n8548 VSS.n1717 0.04025
R17303 VSS.n8544 VSS.n1717 0.04025
R17304 VSS.n8544 VSS.n8543 0.04025
R17305 VSS.n8543 VSS.n8542 0.04025
R17306 VSS.n8542 VSS.n1719 0.04025
R17307 VSS.n8538 VSS.n1719 0.04025
R17308 VSS.n8538 VSS.n8537 0.04025
R17309 VSS.n8537 VSS.n8536 0.04025
R17310 VSS.n8536 VSS.n1721 0.04025
R17311 VSS.n8532 VSS.n1721 0.04025
R17312 VSS.n8532 VSS.n8531 0.04025
R17313 VSS.n8531 VSS.n8530 0.04025
R17314 VSS.n8530 VSS.n1723 0.04025
R17315 VSS.n8526 VSS.n1723 0.04025
R17316 VSS.n8526 VSS.n8525 0.04025
R17317 VSS.n8525 VSS.n8524 0.04025
R17318 VSS.n8524 VSS.n1725 0.04025
R17319 VSS.n8520 VSS.n1725 0.04025
R17320 VSS.n8520 VSS.n8519 0.04025
R17321 VSS.n8519 VSS.n8518 0.04025
R17322 VSS.n8518 VSS.n1727 0.04025
R17323 VSS.n8514 VSS.n1727 0.04025
R17324 VSS.n8514 VSS.n8513 0.04025
R17325 VSS.n8513 VSS.n8512 0.04025
R17326 VSS.n8512 VSS.n1729 0.04025
R17327 VSS.n8508 VSS.n1729 0.04025
R17328 VSS.n8508 VSS.n8507 0.04025
R17329 VSS.n8507 VSS.n8506 0.04025
R17330 VSS.n8506 VSS.n1731 0.04025
R17331 VSS.n8502 VSS.n1731 0.04025
R17332 VSS.n8502 VSS.n8501 0.04025
R17333 VSS.n8501 VSS.n8500 0.04025
R17334 VSS.n8500 VSS.n1733 0.04025
R17335 VSS.n8496 VSS.n1733 0.04025
R17336 VSS.n8496 VSS.n8495 0.04025
R17337 VSS.n8495 VSS.n8494 0.04025
R17338 VSS.n8494 VSS.n1735 0.04025
R17339 VSS.n8490 VSS.n1735 0.04025
R17340 VSS.n8490 VSS.n8489 0.04025
R17341 VSS.n8489 VSS.n8488 0.04025
R17342 VSS.n8488 VSS.n1737 0.04025
R17343 VSS.n8484 VSS.n1737 0.04025
R17344 VSS.n8484 VSS.n8483 0.04025
R17345 VSS.n8483 VSS.n8482 0.04025
R17346 VSS.n8482 VSS.n1739 0.04025
R17347 VSS.n8478 VSS.n1739 0.04025
R17348 VSS.n8478 VSS.n8477 0.04025
R17349 VSS.n8477 VSS.n8476 0.04025
R17350 VSS.n8476 VSS.n1741 0.04025
R17351 VSS.n8472 VSS.n1741 0.04025
R17352 VSS.n8472 VSS.n8471 0.04025
R17353 VSS.n8471 VSS.n8470 0.04025
R17354 VSS.n8470 VSS.n1743 0.04025
R17355 VSS.n8466 VSS.n1743 0.04025
R17356 VSS.n8466 VSS.n8465 0.04025
R17357 VSS.n8465 VSS.n8464 0.04025
R17358 VSS.n8464 VSS.n1745 0.04025
R17359 VSS.n8460 VSS.n1745 0.04025
R17360 VSS.n8460 VSS.n8459 0.04025
R17361 VSS.n8459 VSS.n8458 0.04025
R17362 VSS.n8458 VSS.n1747 0.04025
R17363 VSS.n8454 VSS.n1747 0.04025
R17364 VSS.n8454 VSS.n8453 0.04025
R17365 VSS.n8453 VSS.n8452 0.04025
R17366 VSS.n8452 VSS.n1749 0.04025
R17367 VSS.n8448 VSS.n1749 0.04025
R17368 VSS.n8448 VSS.n8447 0.04025
R17369 VSS.n8447 VSS.n8446 0.04025
R17370 VSS.n8446 VSS.n1751 0.04025
R17371 VSS.n8442 VSS.n1751 0.04025
R17372 VSS.n8442 VSS.n8441 0.04025
R17373 VSS.n8441 VSS.n8440 0.04025
R17374 VSS.n8440 VSS.n1753 0.04025
R17375 VSS.n8436 VSS.n1753 0.04025
R17376 VSS.n8436 VSS.n8435 0.04025
R17377 VSS.n8435 VSS.n8434 0.04025
R17378 VSS.n8434 VSS.n1755 0.04025
R17379 VSS.n8430 VSS.n1755 0.04025
R17380 VSS.n8430 VSS.n8429 0.04025
R17381 VSS.n8429 VSS.n8428 0.04025
R17382 VSS.n8428 VSS.n1757 0.04025
R17383 VSS.n8424 VSS.n1757 0.04025
R17384 VSS.n8424 VSS.n8423 0.04025
R17385 VSS.n8423 VSS.n8422 0.04025
R17386 VSS.n8422 VSS.n1759 0.04025
R17387 VSS.n8418 VSS.n1759 0.04025
R17388 VSS.n8418 VSS.n8417 0.04025
R17389 VSS.n8417 VSS.n8416 0.04025
R17390 VSS.n8416 VSS.n1761 0.04025
R17391 VSS.n8412 VSS.n1761 0.04025
R17392 VSS.n8412 VSS.n8411 0.04025
R17393 VSS.n8411 VSS.n8410 0.04025
R17394 VSS.n8410 VSS.n1763 0.04025
R17395 VSS.n8406 VSS.n1763 0.04025
R17396 VSS.n8406 VSS.n8405 0.04025
R17397 VSS.n8405 VSS.n8404 0.04025
R17398 VSS.n8404 VSS.n1765 0.04025
R17399 VSS.n8400 VSS.n1765 0.04025
R17400 VSS.n8400 VSS.n8399 0.04025
R17401 VSS.n8399 VSS.n8398 0.04025
R17402 VSS.n8398 VSS.n1767 0.04025
R17403 VSS.n8394 VSS.n1767 0.04025
R17404 VSS.n8394 VSS.n8393 0.04025
R17405 VSS.n8393 VSS.n8392 0.04025
R17406 VSS.n8392 VSS.n1769 0.04025
R17407 VSS.n8388 VSS.n1769 0.04025
R17408 VSS.n8388 VSS.n8387 0.04025
R17409 VSS.n8387 VSS.n8386 0.04025
R17410 VSS.n8386 VSS.n1771 0.04025
R17411 VSS.n8382 VSS.n1771 0.04025
R17412 VSS.n8382 VSS.n8381 0.04025
R17413 VSS.n8381 VSS.n8380 0.04025
R17414 VSS.n8380 VSS.n1773 0.04025
R17415 VSS.n8376 VSS.n1773 0.04025
R17416 VSS.n8376 VSS.n8375 0.04025
R17417 VSS.n8375 VSS.n8374 0.04025
R17418 VSS.n8374 VSS.n1775 0.04025
R17419 VSS.n8370 VSS.n1775 0.04025
R17420 VSS.n8370 VSS.n8369 0.04025
R17421 VSS.n8369 VSS.n8368 0.04025
R17422 VSS.n8368 VSS.n1777 0.04025
R17423 VSS.n8364 VSS.n1777 0.04025
R17424 VSS.n8364 VSS.n8363 0.04025
R17425 VSS.n8363 VSS.n8362 0.04025
R17426 VSS.n8362 VSS.n1779 0.04025
R17427 VSS.n8358 VSS.n1779 0.04025
R17428 VSS.n8358 VSS.n8357 0.04025
R17429 VSS.n8357 VSS.n8356 0.04025
R17430 VSS.n8356 VSS.n1781 0.04025
R17431 VSS.n8352 VSS.n1781 0.04025
R17432 VSS.n8352 VSS.n8351 0.04025
R17433 VSS.n8351 VSS.n8350 0.04025
R17434 VSS.n8350 VSS.n1783 0.04025
R17435 VSS.n8346 VSS.n1783 0.04025
R17436 VSS.n8346 VSS.n8345 0.04025
R17437 VSS.n8345 VSS.n8344 0.04025
R17438 VSS.n8344 VSS.n1785 0.04025
R17439 VSS.n8340 VSS.n1785 0.04025
R17440 VSS.n8340 VSS.n8339 0.04025
R17441 VSS.n8339 VSS.n8338 0.04025
R17442 VSS.n8338 VSS.n1787 0.04025
R17443 VSS.n8334 VSS.n1787 0.04025
R17444 VSS.n8334 VSS.n8333 0.04025
R17445 VSS.n8333 VSS.n8332 0.04025
R17446 VSS.n8332 VSS.n1789 0.04025
R17447 VSS.n8328 VSS.n1789 0.04025
R17448 VSS.n8328 VSS.n8327 0.04025
R17449 VSS.n8327 VSS.n8326 0.04025
R17450 VSS.n8326 VSS.n1791 0.04025
R17451 VSS.n8322 VSS.n1791 0.04025
R17452 VSS.n8322 VSS.n8321 0.04025
R17453 VSS.n8321 VSS.n8320 0.04025
R17454 VSS.n8320 VSS.n1793 0.04025
R17455 VSS.n8316 VSS.n1793 0.04025
R17456 VSS.n8316 VSS.n8315 0.04025
R17457 VSS.n8315 VSS.n8314 0.04025
R17458 VSS.n8314 VSS.n1795 0.04025
R17459 VSS.n8310 VSS.n1795 0.04025
R17460 VSS.n8310 VSS.n8309 0.04025
R17461 VSS.n8309 VSS.n8308 0.04025
R17462 VSS.n8308 VSS.n1797 0.04025
R17463 VSS.n8304 VSS.n1797 0.04025
R17464 VSS.n8304 VSS.n8303 0.04025
R17465 VSS.n8303 VSS.n8302 0.04025
R17466 VSS.n8302 VSS.n1799 0.04025
R17467 VSS.n8298 VSS.n1799 0.04025
R17468 VSS.n8298 VSS.n8297 0.04025
R17469 VSS.n8297 VSS.n8296 0.04025
R17470 VSS.n8296 VSS.n1801 0.04025
R17471 VSS.n8292 VSS.n1801 0.04025
R17472 VSS.n8292 VSS.n8291 0.04025
R17473 VSS.n8291 VSS.n8290 0.04025
R17474 VSS.n8290 VSS.n1803 0.04025
R17475 VSS.n8286 VSS.n1803 0.04025
R17476 VSS.n8286 VSS.n8285 0.04025
R17477 VSS.n8285 VSS.n8284 0.04025
R17478 VSS.n8284 VSS.n1805 0.04025
R17479 VSS.n8280 VSS.n1805 0.04025
R17480 VSS.n8280 VSS.n8279 0.04025
R17481 VSS.n8279 VSS.n8278 0.04025
R17482 VSS.n8278 VSS.n1807 0.04025
R17483 VSS.n8274 VSS.n1807 0.04025
R17484 VSS.n8274 VSS.n8273 0.04025
R17485 VSS.n8273 VSS.n8272 0.04025
R17486 VSS.n8272 VSS.n1809 0.04025
R17487 VSS.n8268 VSS.n1809 0.04025
R17488 VSS.n8268 VSS.n8267 0.04025
R17489 VSS.n8267 VSS.n8266 0.04025
R17490 VSS.n8266 VSS.n1811 0.04025
R17491 VSS.n8262 VSS.n1811 0.04025
R17492 VSS.n8262 VSS.n8261 0.04025
R17493 VSS.n8261 VSS.n8260 0.04025
R17494 VSS.n8260 VSS.n1813 0.04025
R17495 VSS.n8256 VSS.n1813 0.04025
R17496 VSS.n8256 VSS.n8255 0.04025
R17497 VSS.n8255 VSS.n8254 0.04025
R17498 VSS.n8254 VSS.n1815 0.04025
R17499 VSS.n8250 VSS.n1815 0.04025
R17500 VSS.n8250 VSS.n8249 0.04025
R17501 VSS.n8249 VSS.n8248 0.04025
R17502 VSS.n8248 VSS.n1817 0.04025
R17503 VSS.n8244 VSS.n1817 0.04025
R17504 VSS.n8244 VSS.n8243 0.04025
R17505 VSS.n8243 VSS.n8242 0.04025
R17506 VSS.n8242 VSS.n1819 0.04025
R17507 VSS.n8238 VSS.n1819 0.04025
R17508 VSS.n8238 VSS.n8237 0.04025
R17509 VSS.n8237 VSS.n8236 0.04025
R17510 VSS.n8236 VSS.n1821 0.04025
R17511 VSS.n8232 VSS.n1821 0.04025
R17512 VSS.n10642 VSS.n10641 0.039811
R17513 VSS.n11335 VSS.n11334 0.0390622
R17514 VSS.n77 VSS.n76 0.0390622
R17515 VSS.n11398 VSS.n0 0.0389239
R17516 VSS.n1575 VSS.n1573 0.0385696
R17517 VSS.n8962 VSS.n8961 0.0385696
R17518 VSS.n962 VSS.n961 0.0385696
R17519 VSS.n10280 VSS.n10279 0.0385696
R17520 VSS.n10454 VSS.n10453 0.0385295
R17521 VSS.n10476 VSS.n10475 0.0385295
R17522 VSS VSS.n0 0.0379215
R17523 VSS.n65 VSS.n63 0.0377578
R17524 VSS.n11333 VSS.n11332 0.0371211
R17525 VSS.n11328 VSS.n11327 0.0371211
R17526 VSS.n67 VSS.n66 0.0371211
R17527 VSS.n74 VSS.n73 0.0371211
R17528 VSS.n1577 VSS.n1576 0.0366533
R17529 VSS.n8959 VSS.n8958 0.0366533
R17530 VSS.n960 VSS.n959 0.0366533
R17531 VSS.n10282 VSS.n10281 0.0366533
R17532 VSS.n11326 VSS.n11325 0.0366035
R17533 VSS.n9434 VSS.n9433 0.0359944
R17534 VSS.n10868 VSS.n238 0.0359286
R17535 VSS.n11337 VSS.n111 0.0359286
R17536 VSS.n11399 VSS.n58 0.0359286
R17537 VSS.n10536 VSS.n10493 0.0359286
R17538 VSS VSS.n11470 0.0357042
R17539 VSS.n9448 VSS.n9447 0.035639
R17540 VSS.n10670 VSS.n10669 0.0354077
R17541 VSS.n10358 VSS.n10357 0.0354077
R17542 VSS.n10424 VSS.n10423 0.0354077
R17543 VSS.n10432 VSS.n10431 0.0354077
R17544 VSS.n10469 VSS.n10468 0.0353617
R17545 VSS.n10461 VSS.n10460 0.0353617
R17546 VSS.n10867 VSS.n239 0.0345
R17547 VSS.n11315 VSS.n106 0.0345
R17548 VSS.n11389 VSS.n11388 0.0345
R17549 VSS.n11394 VSS.n11393 0.0345
R17550 VSS.n11320 VSS.n11319 0.0345
R17551 VSS.n35 VSS.n34 0.0345
R17552 VSS.n10706 VSS.n10705 0.0345
R17553 VSS.n10529 VSS.n10499 0.0345
R17554 VSS.n11313 VSS.n11312 0.0345
R17555 VSS.n10566 VSS.n10565 0.0345
R17556 VSS.n10865 VSS.n225 0.0345
R17557 VSS.n10605 VSS.n10604 0.0342762
R17558 VSS.n10753 VSS.n10752 0.0342758
R17559 VSS.n8979 VSS.n8971 0.0341
R17560 VSS.n8977 VSS.n8971 0.0341
R17561 VSS.n8972 VSS.n1554 0.0341
R17562 VSS.n9096 VSS.n9095 0.0341
R17563 VSS.n9097 VSS.n9096 0.0341
R17564 VSS.n9097 VSS.n1553 0.0341
R17565 VSS.n9099 VSS.n1553 0.0341
R17566 VSS.n8966 VSS.n8965 0.0341
R17567 VSS.n8967 VSS.n8966 0.0341
R17568 VSS.n8967 VSS.n1565 0.0341
R17569 VSS.n8969 VSS.n1565 0.0341
R17570 VSS.n9007 VSS.n8970 0.0341
R17571 VSS.n9005 VSS.n8970 0.0341
R17572 VSS.n9005 VSS.n9004 0.0341
R17573 VSS.n9004 VSS.n9003 0.0341
R17574 VSS.n842 VSS.n838 0.0341
R17575 VSS.n840 VSS.n838 0.0341
R17576 VSS.n840 VSS.n839 0.0341
R17577 VSS.n839 VSS.n221 0.0341
R17578 VSS.n10926 VSS.n222 0.0341
R17579 VSS.n10924 VSS.n222 0.0341
R17580 VSS.n10924 VSS.n10923 0.0341
R17581 VSS.n10923 VSS.n10922 0.0341
R17582 VSS.n877 VSS.n836 0.0341
R17583 VSS.n875 VSS.n836 0.0341
R17584 VSS.n870 VSS.n869 0.0341
R17585 VSS.n866 VSS.n837 0.0341
R17586 VSS.n864 VSS.n837 0.0341
R17587 VSS.n864 VSS.n863 0.0341
R17588 VSS.n863 VSS.n862 0.0341
R17589 VSS.n1121 VSS.n1120 0.0341
R17590 VSS.n1122 VSS.n1121 0.0341
R17591 VSS.n1122 VSS.n879 0.0341
R17592 VSS.n1124 VSS.n879 0.0341
R17593 VSS.n1127 VSS.n1126 0.0341
R17594 VSS.n1128 VSS.n1127 0.0341
R17595 VSS.n1128 VSS.n878 0.0341
R17596 VSS.n1130 VSS.n878 0.0341
R17597 VSS.n1109 VSS.n1108 0.0341
R17598 VSS.n1110 VSS.n1109 0.0341
R17599 VSS.n1110 VSS.n902 0.0341
R17600 VSS.n1112 VSS.n902 0.0341
R17601 VSS.n1115 VSS.n1114 0.0341
R17602 VSS.n1116 VSS.n1115 0.0341
R17603 VSS.n1116 VSS.n901 0.0341
R17604 VSS.n1118 VSS.n901 0.0341
R17605 VSS.n1084 VSS.n1083 0.0341
R17606 VSS.n1089 VSS.n1084 0.0341
R17607 VSS.n1091 VSS.n904 0.0341
R17608 VSS.n1094 VSS.n1093 0.0341
R17609 VSS.n1095 VSS.n1094 0.0341
R17610 VSS.n1095 VSS.n903 0.0341
R17611 VSS.n1097 VSS.n903 0.0341
R17612 VSS.n1072 VSS.n1071 0.0341
R17613 VSS.n1073 VSS.n1072 0.0341
R17614 VSS.n1073 VSS.n915 0.0341
R17615 VSS.n1075 VSS.n915 0.0341
R17616 VSS.n1078 VSS.n1077 0.0341
R17617 VSS.n1079 VSS.n1078 0.0341
R17618 VSS.n1079 VSS.n914 0.0341
R17619 VSS.n1081 VSS.n914 0.0341
R17620 VSS.n1051 VSS.n1050 0.0341
R17621 VSS.n1052 VSS.n1051 0.0341
R17622 VSS.n1052 VSS.n917 0.0341
R17623 VSS.n1054 VSS.n917 0.0341
R17624 VSS.n1057 VSS.n1056 0.0341
R17625 VSS.n1058 VSS.n1057 0.0341
R17626 VSS.n1058 VSS.n916 0.0341
R17627 VSS.n1060 VSS.n916 0.0341
R17628 VSS.n1035 VSS.n1034 0.0341
R17629 VSS.n1040 VSS.n1035 0.0341
R17630 VSS.n1042 VSS.n928 0.0341
R17631 VSS.n1045 VSS.n1044 0.0341
R17632 VSS.n1046 VSS.n1045 0.0341
R17633 VSS.n1046 VSS.n927 0.0341
R17634 VSS.n1048 VSS.n927 0.0341
R17635 VSS.n1014 VSS.n1013 0.0341
R17636 VSS.n1015 VSS.n1014 0.0341
R17637 VSS.n1015 VSS.n930 0.0341
R17638 VSS.n1017 VSS.n930 0.0341
R17639 VSS.n1020 VSS.n1019 0.0341
R17640 VSS.n1021 VSS.n1020 0.0341
R17641 VSS.n1021 VSS.n929 0.0341
R17642 VSS.n1023 VSS.n929 0.0341
R17643 VSS.n1002 VSS.n1001 0.0341
R17644 VSS.n1003 VSS.n1002 0.0341
R17645 VSS.n1003 VSS.n941 0.0341
R17646 VSS.n1005 VSS.n941 0.0341
R17647 VSS.n1008 VSS.n1007 0.0341
R17648 VSS.n1009 VSS.n1008 0.0341
R17649 VSS.n1009 VSS.n940 0.0341
R17650 VSS.n1011 VSS.n940 0.0341
R17651 VSS.n977 VSS.n976 0.0341
R17652 VSS.n982 VSS.n977 0.0341
R17653 VSS.n984 VSS.n943 0.0341
R17654 VSS.n987 VSS.n986 0.0341
R17655 VSS.n988 VSS.n987 0.0341
R17656 VSS.n988 VSS.n942 0.0341
R17657 VSS.n990 VSS.n942 0.0341
R17658 VSS.n965 VSS.n964 0.0341
R17659 VSS.n966 VSS.n965 0.0341
R17660 VSS.n966 VSS.n954 0.0341
R17661 VSS.n968 VSS.n954 0.0341
R17662 VSS.n971 VSS.n970 0.0341
R17663 VSS.n972 VSS.n971 0.0341
R17664 VSS.n972 VSS.n953 0.0341
R17665 VSS.n974 VSS.n953 0.0341
R17666 VSS.n10920 VSS.n10916 0.0341
R17667 VSS.n10918 VSS.n10916 0.0341
R17668 VSS.n10918 VSS.n10917 0.0341
R17669 VSS.n10917 VSS.n207 0.0341
R17670 VSS.n10986 VSS.n10985 0.0341
R17671 VSS.n10987 VSS.n10986 0.0341
R17672 VSS.n10987 VSS.n206 0.0341
R17673 VSS.n10989 VSS.n206 0.0341
R17674 VSS.n10998 VSS.n10990 0.0341
R17675 VSS.n10996 VSS.n10990 0.0341
R17676 VSS.n10991 VSS.n96 0.0341
R17677 VSS.n11358 VSS.n97 0.0341
R17678 VSS.n11356 VSS.n97 0.0341
R17679 VSS.n11356 VSS.n11355 0.0341
R17680 VSS.n11355 VSS.n11354 0.0341
R17681 VSS.n11352 VSS.n101 0.0341
R17682 VSS.n11350 VSS.n101 0.0341
R17683 VSS.n11350 VSS.n11349 0.0341
R17684 VSS.n11349 VSS.n11348 0.0341
R17685 VSS.n11345 VSS.n102 0.0341
R17686 VSS.n11343 VSS.n102 0.0341
R17687 VSS.n11343 VSS.n11342 0.0341
R17688 VSS.n11342 VSS.n11341 0.0341
R17689 VSS.n11371 VSS.n11370 0.0341
R17690 VSS.n11372 VSS.n11371 0.0341
R17691 VSS.n11372 VSS.n85 0.0341
R17692 VSS.n11374 VSS.n85 0.0341
R17693 VSS.n11378 VSS.n11377 0.0341
R17694 VSS.n11379 VSS.n11378 0.0341
R17695 VSS.n11379 VSS.n84 0.0341
R17696 VSS.n11381 VSS.n84 0.0341
R17697 VSS.n10952 VSS.n10944 0.0341
R17698 VSS.n10950 VSS.n10944 0.0341
R17699 VSS.n10945 VSS.n90 0.0341
R17700 VSS.n11365 VSS.n11364 0.0341
R17701 VSS.n11366 VSS.n11365 0.0341
R17702 VSS.n11366 VSS.n89 0.0341
R17703 VSS.n11368 VSS.n89 0.0341
R17704 VSS.n10939 VSS.n10938 0.0341
R17705 VSS.n10940 VSS.n10939 0.0341
R17706 VSS.n10940 VSS.n209 0.0341
R17707 VSS.n10942 VSS.n209 0.0341
R17708 VSS.n10979 VSS.n10943 0.0341
R17709 VSS.n10977 VSS.n10943 0.0341
R17710 VSS.n10977 VSS.n10976 0.0341
R17711 VSS.n10976 VSS.n10975 0.0341
R17712 VSS.n1168 VSS.n1164 0.0341
R17713 VSS.n1166 VSS.n1164 0.0341
R17714 VSS.n1166 VSS.n1165 0.0341
R17715 VSS.n1165 VSS.n214 0.0341
R17716 VSS.n10933 VSS.n10932 0.0341
R17717 VSS.n10934 VSS.n10933 0.0341
R17718 VSS.n10934 VSS.n213 0.0341
R17719 VSS.n10936 VSS.n213 0.0341
R17720 VSS.n1214 VSS.n1162 0.0341
R17721 VSS.n1212 VSS.n1162 0.0341
R17722 VSS.n1207 VSS.n1206 0.0341
R17723 VSS.n1204 VSS.n1163 0.0341
R17724 VSS.n1202 VSS.n1163 0.0341
R17725 VSS.n1202 VSS.n1201 0.0341
R17726 VSS.n1201 VSS.n1200 0.0341
R17727 VSS.n9537 VSS.n9536 0.0341
R17728 VSS.n9538 VSS.n9537 0.0341
R17729 VSS.n9538 VSS.n1216 0.0341
R17730 VSS.n9540 VSS.n1216 0.0341
R17731 VSS.n9544 VSS.n9543 0.0341
R17732 VSS.n9545 VSS.n9544 0.0341
R17733 VSS.n9545 VSS.n1215 0.0341
R17734 VSS.n9547 VSS.n1215 0.0341
R17735 VSS.n1402 VSS.n1398 0.0341
R17736 VSS.n1400 VSS.n1398 0.0341
R17737 VSS.n1400 VSS.n1399 0.0341
R17738 VSS.n1399 VSS.n1221 0.0341
R17739 VSS.n9531 VSS.n9530 0.0341
R17740 VSS.n9532 VSS.n9531 0.0341
R17741 VSS.n9532 VSS.n1220 0.0341
R17742 VSS.n9534 VSS.n1220 0.0341
R17743 VSS.n1494 VSS.n1486 0.0341
R17744 VSS.n1492 VSS.n1486 0.0341
R17745 VSS.n1487 VSS.n1396 0.0341
R17746 VSS.n9419 VSS.n1397 0.0341
R17747 VSS.n9417 VSS.n1397 0.0341
R17748 VSS.n9417 VSS.n9416 0.0341
R17749 VSS.n9416 VSS.n9415 0.0341
R17750 VSS.n9268 VSS.n9264 0.0341
R17751 VSS.n9266 VSS.n9264 0.0341
R17752 VSS.n9266 VSS.n9265 0.0341
R17753 VSS.n9265 VSS.n1496 0.0341
R17754 VSS.n9351 VSS.n9350 0.0341
R17755 VSS.n9352 VSS.n9351 0.0341
R17756 VSS.n9352 VSS.n1495 0.0341
R17757 VSS.n9354 VSS.n1495 0.0341
R17758 VSS.n9259 VSS.n9258 0.0341
R17759 VSS.n9260 VSS.n9259 0.0341
R17760 VSS.n9260 VSS.n1508 0.0341
R17761 VSS.n9262 VSS.n1508 0.0341
R17762 VSS.n9296 VSS.n9263 0.0341
R17763 VSS.n9294 VSS.n9263 0.0341
R17764 VSS.n9294 VSS.n9293 0.0341
R17765 VSS.n9293 VSS.n9292 0.0341
R17766 VSS.n9146 VSS.n9138 0.0341
R17767 VSS.n9144 VSS.n9138 0.0341
R17768 VSS.n9139 VSS.n1513 0.0341
R17769 VSS.n9253 VSS.n9252 0.0341
R17770 VSS.n9254 VSS.n9253 0.0341
R17771 VSS.n9254 VSS.n1512 0.0341
R17772 VSS.n9256 VSS.n1512 0.0341
R17773 VSS.n9133 VSS.n9132 0.0341
R17774 VSS.n9134 VSS.n9133 0.0341
R17775 VSS.n9134 VSS.n1526 0.0341
R17776 VSS.n9136 VSS.n1526 0.0341
R17777 VSS.n9174 VSS.n9137 0.0341
R17778 VSS.n9172 VSS.n9137 0.0341
R17779 VSS.n9172 VSS.n9171 0.0341
R17780 VSS.n9171 VSS.n9170 0.0341
R17781 VSS.n1552 VSS.n1541 0.0341
R17782 VSS.n1550 VSS.n1541 0.0341
R17783 VSS.n1550 VSS.n1549 0.0341
R17784 VSS.n1549 VSS.n1548 0.0341
R17785 VSS.n1546 VSS.n1542 0.0341
R17786 VSS.n1544 VSS.n1542 0.0341
R17787 VSS.n1544 VSS.n1543 0.0341
R17788 VSS.n1543 VSS.n1527 0.0341
R17789 VSS.n11401 VSS.n11400 0.033821
R17790 VSS.n10676 VSS.n10336 0.0337454
R17791 VSS.n10674 VSS.n10336 0.0337454
R17792 VSS.n10674 VSS.n10673 0.0337454
R17793 VSS.n10673 VSS.n10672 0.0337454
R17794 VSS.n10672 VSS.n10337 0.0337454
R17795 VSS.n10670 VSS.n10337 0.0337454
R17796 VSS.n10669 VSS.n10338 0.0337454
R17797 VSS.n10667 VSS.n10338 0.0337454
R17798 VSS.n10667 VSS.n10666 0.0337454
R17799 VSS.n10355 VSS.n10339 0.0337454
R17800 VSS.n10357 VSS.n10355 0.0337454
R17801 VSS.n10358 VSS.n10354 0.0337454
R17802 VSS.n10360 VSS.n10354 0.0337454
R17803 VSS.n10361 VSS.n10360 0.0337454
R17804 VSS.n10362 VSS.n10361 0.0337454
R17805 VSS.n10362 VSS.n10353 0.0337454
R17806 VSS.n10364 VSS.n10353 0.0337454
R17807 VSS.n10417 VSS.n10291 0.0337454
R17808 VSS.n10419 VSS.n10417 0.0337454
R17809 VSS.n10420 VSS.n10419 0.0337454
R17810 VSS.n10421 VSS.n10420 0.0337454
R17811 VSS.n10421 VSS.n10416 0.0337454
R17812 VSS.n10423 VSS.n10416 0.0337454
R17813 VSS.n10424 VSS.n10415 0.0337454
R17814 VSS.n10426 VSS.n10415 0.0337454
R17815 VSS.n10427 VSS.n10426 0.0337454
R17816 VSS.n10429 VSS.n10414 0.0337454
R17817 VSS.n10431 VSS.n10414 0.0337454
R17818 VSS.n10432 VSS.n10413 0.0337454
R17819 VSS.n10434 VSS.n10413 0.0337454
R17820 VSS.n10435 VSS.n10434 0.0337454
R17821 VSS.n10436 VSS.n10435 0.0337454
R17822 VSS.n10436 VSS.n10412 0.0337454
R17823 VSS.n10438 VSS.n10412 0.0337454
R17824 VSS.n10475 VSS.n10443 0.0337016
R17825 VSS.n10473 VSS.n10443 0.0337016
R17826 VSS.n10473 VSS.n10472 0.0337016
R17827 VSS.n10472 VSS.n10471 0.0337016
R17828 VSS.n10471 VSS.n10444 0.0337016
R17829 VSS.n10469 VSS.n10444 0.0337016
R17830 VSS.n10468 VSS.n10445 0.0337016
R17831 VSS.n10466 VSS.n10445 0.0337016
R17832 VSS.n10466 VSS.n10465 0.0337016
R17833 VSS.n10463 VSS.n10446 0.0337016
R17834 VSS.n10461 VSS.n10446 0.0337016
R17835 VSS.n10460 VSS.n10447 0.0337016
R17836 VSS.n10458 VSS.n10447 0.0337016
R17837 VSS.n10458 VSS.n10457 0.0337016
R17838 VSS.n10457 VSS.n10456 0.0337016
R17839 VSS.n10456 VSS.n10448 0.0337016
R17840 VSS.n10454 VSS.n10448 0.0337016
R17841 VSS.n10665 VSS.n10339 0.033033
R17842 VSS.n10429 VSS.n10428 0.033033
R17843 VSS.n10464 VSS.n10463 0.0329901
R17844 VSS.n9486 VSS.n9485 0.0329468
R17845 VSS.n9484 VSS.n9483 0.0329468
R17846 VSS.n9482 VSS.n9481 0.0329468
R17847 VSS.n1410 VSS.n1409 0.0329468
R17848 VSS.n1412 VSS.n1411 0.0329468
R17849 VSS.n1414 VSS.n1413 0.0329468
R17850 VSS.n1321 VSS.n1320 0.0329468
R17851 VSS.n1323 VSS.n1322 0.0329468
R17852 VSS.n1325 VSS.n1324 0.0329468
R17853 VSS.n9509 VSS.n9508 0.0329468
R17854 VSS.n10819 VSS.n10818 0.032073
R17855 VSS.n10777 VSS.n10776 0.032073
R17856 VSS.n10788 VSS.n10787 0.032073
R17857 VSS.n9485 VSS.n9477 0.0319894
R17858 VSS.n9484 VSS.n9477 0.0319894
R17859 VSS.n9483 VSS.n9478 0.0319894
R17860 VSS.n9482 VSS.n9478 0.0319894
R17861 VSS.n9481 VSS.n9479 0.0319894
R17862 VSS.n9480 VSS.n9479 0.0319894
R17863 VSS.n1386 VSS.n1385 0.0319894
R17864 VSS.n1408 VSS.n1407 0.0319894
R17865 VSS.n1409 VSS.n1407 0.0319894
R17866 VSS.n1410 VSS.n1406 0.0319894
R17867 VSS.n1411 VSS.n1406 0.0319894
R17868 VSS.n1412 VSS.n1405 0.0319894
R17869 VSS.n1413 VSS.n1405 0.0319894
R17870 VSS.n1414 VSS.n1404 0.0319894
R17871 VSS.n1415 VSS.n1404 0.0319894
R17872 VSS.n1319 VSS.n1271 0.0319894
R17873 VSS.n1320 VSS.n1271 0.0319894
R17874 VSS.n1321 VSS.n1270 0.0319894
R17875 VSS.n1322 VSS.n1270 0.0319894
R17876 VSS.n1323 VSS.n1269 0.0319894
R17877 VSS.n1324 VSS.n1269 0.0319894
R17878 VSS.n1325 VSS.n1268 0.0319894
R17879 VSS.n1326 VSS.n1268 0.0319894
R17880 VSS.n1332 VSS.n1331 0.0319894
R17881 VSS.n9510 VSS.n1334 0.0319894
R17882 VSS.n9509 VSS.n1334 0.0319894
R17883 VSS.n10752 VSS.n10747 0.0319607
R17884 VSS.n10750 VSS.n10747 0.0319607
R17885 VSS.n10750 VSS.n10749 0.0319607
R17886 VSS.n10749 VSS.n10748 0.0319607
R17887 VSS.n10815 VSS.n10814 0.0319607
R17888 VSS.n10816 VSS.n10815 0.0319607
R17889 VSS.n10816 VSS.n10813 0.0319607
R17890 VSS.n10818 VSS.n10813 0.0319607
R17891 VSS.n10778 VSS.n10777 0.0319607
R17892 VSS.n10779 VSS.n10778 0.0319607
R17893 VSS.n10779 VSS.n10737 0.0319607
R17894 VSS.n10781 VSS.n10737 0.0319607
R17895 VSS.n10784 VSS.n10783 0.0319607
R17896 VSS.n10785 VSS.n10784 0.0319607
R17897 VSS.n10785 VSS.n10736 0.0319607
R17898 VSS.n10787 VSS.n10736 0.0319607
R17899 VSS.n10494 VSS.n10441 0.0319161
R17900 VSS.n10582 VSS.n10581 0.0315563
R17901 VSS.n10649 VSS.n10648 0.0315563
R17902 VSS.n10453 VSS.n10452 0.0314767
R17903 VSS.n10451 VSS.n10450 0.0314767
R17904 VSS.n10449 VSS.n10345 0.0314767
R17905 VSS.n10659 VSS.n10658 0.0314767
R17906 VSS.n10657 VSS.n10656 0.0314767
R17907 VSS.n10477 VSS.n10476 0.0314767
R17908 VSS.n10479 VSS.n10478 0.0314767
R17909 VSS.n10481 VSS.n10480 0.0314767
R17910 VSS.n10596 VSS.n10595 0.0314767
R17911 VSS.n10594 VSS.n10593 0.0314767
R17912 VSS.n10560 VSS.n10559 0.0314767
R17913 VSS.n10558 VSS.n10290 0.0314767
R17914 VSS.n10693 VSS.n10692 0.0314767
R17915 VSS.n10691 VSS.n10690 0.0314767
R17916 VSS.n10689 VSS.n10688 0.0314767
R17917 VSS.n10641 VSS.n10640 0.0314767
R17918 VSS.n10572 VSS.n10561 0.0313721
R17919 VSS.n1388 VSS.n1387 0.0311383
R17920 VSS.n1333 VSS.n1330 0.0311383
R17921 VSS.n11331 VSS.n11330 0.0301981
R17922 VSS.n72 VSS.n70 0.0301981
R17923 VSS.n10575 VSS.n10574 0.0301831
R17924 VSS.n10278 VSS.n10277 0.0301505
R17925 VSS.n1572 VSS.n1570 0.0300866
R17926 VSS.n10575 VSS.n10555 0.0300775
R17927 VSS.n10577 VSS.n10555 0.0300775
R17928 VSS.n10578 VSS.n10577 0.0300775
R17929 VSS.n10579 VSS.n10578 0.0300775
R17930 VSS.n10579 VSS.n10554 0.0300775
R17931 VSS.n10581 VSS.n10554 0.0300775
R17932 VSS.n10582 VSS.n10553 0.0300775
R17933 VSS.n10584 VSS.n10553 0.0300775
R17934 VSS.n10585 VSS.n10584 0.0300775
R17935 VSS.n10651 VSS.n10650 0.0300775
R17936 VSS.n10650 VSS.n10649 0.0300775
R17937 VSS.n10648 VSS.n10350 0.0300775
R17938 VSS.n10646 VSS.n10350 0.0300775
R17939 VSS.n10646 VSS.n10645 0.0300775
R17940 VSS.n10645 VSS.n10644 0.0300775
R17941 VSS.n10644 VSS.n10351 0.0300775
R17942 VSS.n10642 VSS.n10351 0.0300775
R17943 VSS.n8965 VSS.n8964 0.0299989
R17944 VSS.n964 VSS.n963 0.0299989
R17945 VSS.n8957 VSS.n8955 0.0298187
R17946 VSS.n9073 VSS.n9046 0.0294988
R17947 VSS.n9071 VSS.n9046 0.0294988
R17948 VSS.n9071 VSS.n9070 0.0294988
R17949 VSS.n9070 VSS.n9069 0.0294988
R17950 VSS.n9067 VSS.n9047 0.0294988
R17951 VSS.n9065 VSS.n9047 0.0294988
R17952 VSS.n9065 VSS.n9064 0.0294988
R17953 VSS.n9064 VSS.n9063 0.0294988
R17954 VSS.n9041 VSS.n9040 0.0294988
R17955 VSS.n9042 VSS.n9041 0.0294988
R17956 VSS.n9042 VSS.n1556 0.0294988
R17957 VSS.n9044 VSS.n1556 0.0294988
R17958 VSS.n9088 VSS.n9045 0.0294988
R17959 VSS.n9086 VSS.n9045 0.0294988
R17960 VSS.n9086 VSS.n9085 0.0294988
R17961 VSS.n9085 VSS.n9084 0.0294988
R17962 VSS.n1570 VSS.n1566 0.0294988
R17963 VSS.n1568 VSS.n1566 0.0294988
R17964 VSS.n1568 VSS.n1567 0.0294988
R17965 VSS.n1567 VSS.n1561 0.0294988
R17966 VSS.n9017 VSS.n9016 0.0294988
R17967 VSS.n9036 VSS.n9017 0.0294988
R17968 VSS.n9036 VSS.n9035 0.0294988
R17969 VSS.n1285 VSS.n416 0.0294988
R17970 VSS.n1286 VSS.n1285 0.0294988
R17971 VSS.n1286 VSS.n1284 0.0294988
R17972 VSS.n1288 VSS.n1284 0.0294988
R17973 VSS.n1291 VSS.n1290 0.0294988
R17974 VSS.n1292 VSS.n1291 0.0294988
R17975 VSS.n1292 VSS.n1283 0.0294988
R17976 VSS.n1294 VSS.n1283 0.0294988
R17977 VSS.n10157 VSS.n401 0.0294988
R17978 VSS.n10155 VSS.n401 0.0294988
R17979 VSS.n10155 VSS.n10154 0.0294988
R17980 VSS.n10154 VSS.n10153 0.0294988
R17981 VSS.n10151 VSS.n402 0.0294988
R17982 VSS.n10149 VSS.n402 0.0294988
R17983 VSS.n10149 VSS.n10148 0.0294988
R17984 VSS.n387 VSS.n386 0.0294988
R17985 VSS.n388 VSS.n387 0.0294988
R17986 VSS.n388 VSS.n363 0.0294988
R17987 VSS.n390 VSS.n363 0.0294988
R17988 VSS.n10160 VSS.n10159 0.0294988
R17989 VSS.n10161 VSS.n10160 0.0294988
R17990 VSS.n10161 VSS.n10158 0.0294988
R17991 VSS.n10163 VSS.n10158 0.0294988
R17992 VSS.n366 VSS.n344 0.0294988
R17993 VSS.n367 VSS.n366 0.0294988
R17994 VSS.n367 VSS.n365 0.0294988
R17995 VSS.n369 VSS.n365 0.0294988
R17996 VSS.n372 VSS.n371 0.0294988
R17997 VSS.n373 VSS.n372 0.0294988
R17998 VSS.n373 VSS.n364 0.0294988
R17999 VSS.n375 VSS.n364 0.0294988
R18000 VSS.n10217 VSS.n329 0.0294988
R18001 VSS.n10215 VSS.n329 0.0294988
R18002 VSS.n10215 VSS.n10214 0.0294988
R18003 VSS.n10214 VSS.n10213 0.0294988
R18004 VSS.n10211 VSS.n330 0.0294988
R18005 VSS.n10209 VSS.n330 0.0294988
R18006 VSS.n10209 VSS.n10208 0.0294988
R18007 VSS.n315 VSS.n314 0.0294988
R18008 VSS.n316 VSS.n315 0.0294988
R18009 VSS.n316 VSS.n291 0.0294988
R18010 VSS.n318 VSS.n291 0.0294988
R18011 VSS.n10220 VSS.n10219 0.0294988
R18012 VSS.n10221 VSS.n10220 0.0294988
R18013 VSS.n10221 VSS.n10218 0.0294988
R18014 VSS.n10223 VSS.n10218 0.0294988
R18015 VSS.n303 VSS.n272 0.0294988
R18016 VSS.n304 VSS.n303 0.0294988
R18017 VSS.n304 VSS.n302 0.0294988
R18018 VSS.n306 VSS.n302 0.0294988
R18019 VSS.n309 VSS.n308 0.0294988
R18020 VSS.n310 VSS.n309 0.0294988
R18021 VSS.n310 VSS.n301 0.0294988
R18022 VSS.n312 VSS.n301 0.0294988
R18023 VSS.n10277 VSS.n257 0.0294988
R18024 VSS.n10275 VSS.n257 0.0294988
R18025 VSS.n10275 VSS.n10274 0.0294988
R18026 VSS.n10274 VSS.n10273 0.0294988
R18027 VSS.n10271 VSS.n258 0.0294988
R18028 VSS.n10269 VSS.n258 0.0294988
R18029 VSS.n10269 VSS.n10268 0.0294988
R18030 VSS.n9377 VSS.n9376 0.0294988
R18031 VSS.n9378 VSS.n9377 0.0294988
R18032 VSS.n9378 VSS.n1477 0.0294988
R18033 VSS.n9380 VSS.n1477 0.0294988
R18034 VSS.n9384 VSS.n9383 0.0294988
R18035 VSS.n9385 VSS.n9384 0.0294988
R18036 VSS.n9385 VSS.n1476 0.0294988
R18037 VSS.n9387 VSS.n1476 0.0294988
R18038 VSS.n9317 VSS.n9316 0.0294988
R18039 VSS.n9318 VSS.n9317 0.0294988
R18040 VSS.n9318 VSS.n1500 0.0294988
R18041 VSS.n9320 VSS.n1500 0.0294988
R18042 VSS.n9343 VSS.n9321 0.0294988
R18043 VSS.n9341 VSS.n9321 0.0294988
R18044 VSS.n9341 VSS.n9340 0.0294988
R18045 VSS.n9217 VSS.n9213 0.0294988
R18046 VSS.n9215 VSS.n9213 0.0294988
R18047 VSS.n9215 VSS.n9214 0.0294988
R18048 VSS.n9214 VSS.n1505 0.0294988
R18049 VSS.n9311 VSS.n9310 0.0294988
R18050 VSS.n9312 VSS.n9311 0.0294988
R18051 VSS.n9312 VSS.n1504 0.0294988
R18052 VSS.n9314 VSS.n1504 0.0294988
R18053 VSS.n9208 VSS.n9207 0.0294988
R18054 VSS.n9209 VSS.n9208 0.0294988
R18055 VSS.n9209 VSS.n1518 0.0294988
R18056 VSS.n9211 VSS.n1518 0.0294988
R18057 VSS.n9245 VSS.n9212 0.0294988
R18058 VSS.n9243 VSS.n9212 0.0294988
R18059 VSS.n9243 VSS.n9242 0.0294988
R18060 VSS.n9242 VSS.n9241 0.0294988
R18061 VSS.n9061 VSS.n9057 0.0294988
R18062 VSS.n9059 VSS.n9057 0.0294988
R18063 VSS.n9059 VSS.n9058 0.0294988
R18064 VSS.n9058 VSS.n1523 0.0294988
R18065 VSS.n9184 VSS.n9183 0.0294988
R18066 VSS.n9203 VSS.n9184 0.0294988
R18067 VSS.n9203 VSS.n9202 0.0294988
R18068 VSS.n10825 VSS.n10821 0.029033
R18069 VSS.n9487 VSS.n9486 0.0286128
R18070 VSS.n10769 VSS.n10768 0.0280818
R18071 VSS.n10634 VSS.n10352 0.0277138
R18072 VSS.n9002 VSS.n8979 0.02738
R18073 VSS.n9100 VSS.n9099 0.02738
R18074 VSS.n9003 VSS.n9002 0.02738
R18075 VSS.n861 VSS.n842 0.02738
R18076 VSS.n10922 VSS.n10921 0.02738
R18077 VSS.n1131 VSS.n877 0.02738
R18078 VSS.n862 VSS.n861 0.02738
R18079 VSS.n1120 VSS.n1119 0.02738
R18080 VSS.n1131 VSS.n1130 0.02738
R18081 VSS.n1108 VSS.n1107 0.02738
R18082 VSS.n1119 VSS.n1118 0.02738
R18083 VSS.n1083 VSS.n1082 0.02738
R18084 VSS.n1107 VSS.n1097 0.02738
R18085 VSS.n1071 VSS.n1070 0.02738
R18086 VSS.n1082 VSS.n1081 0.02738
R18087 VSS.n1050 VSS.n1049 0.02738
R18088 VSS.n1070 VSS.n1060 0.02738
R18089 VSS.n1034 VSS.n1033 0.02738
R18090 VSS.n1049 VSS.n1048 0.02738
R18091 VSS.n1013 VSS.n1012 0.02738
R18092 VSS.n1033 VSS.n1023 0.02738
R18093 VSS.n1001 VSS.n1000 0.02738
R18094 VSS.n1012 VSS.n1011 0.02738
R18095 VSS.n976 VSS.n975 0.02738
R18096 VSS.n1000 VSS.n990 0.02738
R18097 VSS.n975 VSS.n974 0.02738
R18098 VSS.n10921 VSS.n10920 0.02738
R18099 VSS.n10999 VSS.n10989 0.02738
R18100 VSS.n10999 VSS.n10998 0.02738
R18101 VSS.n11354 VSS.n11353 0.02738
R18102 VSS.n11353 VSS.n11352 0.02738
R18103 VSS.n11341 VSS.n11340 0.02738
R18104 VSS.n11370 VSS.n11369 0.02738
R18105 VSS.n11382 VSS.n11381 0.02738
R18106 VSS.n10974 VSS.n10952 0.02738
R18107 VSS.n11369 VSS.n11368 0.02738
R18108 VSS.n10938 VSS.n10937 0.02738
R18109 VSS.n10975 VSS.n10974 0.02738
R18110 VSS.n1199 VSS.n1168 0.02738
R18111 VSS.n10937 VSS.n10936 0.02738
R18112 VSS.n9548 VSS.n1214 0.02738
R18113 VSS.n1200 VSS.n1199 0.02738
R18114 VSS.n9536 VSS.n9535 0.02738
R18115 VSS.n9548 VSS.n9547 0.02738
R18116 VSS.n9414 VSS.n1402 0.02738
R18117 VSS.n9535 VSS.n9534 0.02738
R18118 VSS.n9355 VSS.n1494 0.02738
R18119 VSS.n9415 VSS.n9414 0.02738
R18120 VSS.n9291 VSS.n9268 0.02738
R18121 VSS.n9355 VSS.n9354 0.02738
R18122 VSS.n9258 VSS.n9257 0.02738
R18123 VSS.n9292 VSS.n9291 0.02738
R18124 VSS.n9169 VSS.n9146 0.02738
R18125 VSS.n9257 VSS.n9256 0.02738
R18126 VSS.n9132 VSS.n9131 0.02738
R18127 VSS.n9170 VSS.n9169 0.02738
R18128 VSS.n9100 VSS.n1552 0.02738
R18129 VSS.n9131 VSS.n1527 0.02738
R18130 VSS.n10633 VSS.n10364 0.0271502
R18131 VSS.n10842 VSS.n10841 0.0261855
R18132 VSS.n10763 VSS.n10762 0.0259315
R18133 VSS.n10746 VSS.n10745 0.0255699
R18134 VSS.n9198 VSS.n9186 0.0255051
R18135 VSS.n9335 VSS.n9334 0.0255051
R18136 VSS.n172 VSS.n160 0.0255051
R18137 VSS.n9582 VSS.n9580 0.0255051
R18138 VSS.n11140 VSS.n200 0.0255051
R18139 VSS.n482 VSS.n481 0.0255051
R18140 VSS.n9031 VSS.n9019 0.0255051
R18141 VSS.n10263 VSS.n271 0.0255051
R18142 VSS.n10203 VSS.n343 0.0255051
R18143 VSS.n10143 VSS.n415 0.0255051
R18144 VSS.n10823 VSS.n10822 0.024829
R18145 VSS.n9083 VSS.n9073 0.0236991
R18146 VSS.n9063 VSS.n9062 0.0236991
R18147 VSS.n9040 VSS.n9039 0.0236991
R18148 VSS.n9084 VSS.n9083 0.0236991
R18149 VSS.n9039 VSS.n9038 0.0236991
R18150 VSS.n10141 VSS.n416 0.0236991
R18151 VSS.n1295 VSS.n1294 0.0236991
R18152 VSS.n10164 VSS.n10157 0.0236991
R18153 VSS.n10142 VSS.n10141 0.0236991
R18154 VSS.n386 VSS.n385 0.0236991
R18155 VSS.n10164 VSS.n10163 0.0236991
R18156 VSS.n10201 VSS.n344 0.0236991
R18157 VSS.n385 VSS.n375 0.0236991
R18158 VSS.n10224 VSS.n10217 0.0236991
R18159 VSS.n10202 VSS.n10201 0.0236991
R18160 VSS.n314 VSS.n313 0.0236991
R18161 VSS.n10224 VSS.n10223 0.0236991
R18162 VSS.n10261 VSS.n272 0.0236991
R18163 VSS.n313 VSS.n312 0.0236991
R18164 VSS.n10262 VSS.n10261 0.0236991
R18165 VSS.n9376 VSS.n9375 0.0236991
R18166 VSS.n9388 VSS.n9387 0.0236991
R18167 VSS.n9316 VSS.n9315 0.0236991
R18168 VSS.n9375 VSS.n1478 0.0236991
R18169 VSS.n9240 VSS.n9217 0.0236991
R18170 VSS.n9315 VSS.n9314 0.0236991
R18171 VSS.n9207 VSS.n9206 0.0236991
R18172 VSS.n9241 VSS.n9240 0.0236991
R18173 VSS.n9062 VSS.n9061 0.0236991
R18174 VSS.n9206 VSS.n9205 0.0236991
R18175 VSS.n10651 VSS.n10349 0.0231186
R18176 VSS.n6936 VSS.n61 0.023
R18177 VSS.n10843 VSS.n10733 0.0229499
R18178 VSS.n8977 VSS.n8976 0.022805
R18179 VSS.n875 VSS.n874 0.022805
R18180 VSS.n1089 VSS.n1088 0.022805
R18181 VSS.n1040 VSS.n1039 0.022805
R18182 VSS.n982 VSS.n981 0.022805
R18183 VSS.n10996 VSS.n10995 0.022805
R18184 VSS.n10950 VSS.n10949 0.022805
R18185 VSS.n1212 VSS.n1211 0.022805
R18186 VSS.n1492 VSS.n1491 0.022805
R18187 VSS.n9144 VSS.n9143 0.022805
R18188 VSS.n10639 VSS.n10638 0.0217442
R18189 VSS.n9200 VSS.n9198 0.0215309
R18190 VSS.n9338 VSS.n9334 0.0215309
R18191 VSS.n175 VSS.n172 0.0215309
R18192 VSS.n9585 VSS.n9580 0.0215309
R18193 VSS.n11143 VSS.n200 0.0215309
R18194 VSS.n481 VSS.n480 0.0215309
R18195 VSS.n9033 VSS.n9031 0.0215309
R18196 VSS.n10266 VSS.n271 0.0215309
R18197 VSS.n10206 VSS.n343 0.0215309
R18198 VSS.n10146 VSS.n415 0.0215309
R18199 VSS.n10688 VSS.n10687 0.0213083
R18200 VSS.n10496 VSS.n10495 0.0209545
R18201 VSS.n10607 VSS.n10606 0.0208496
R18202 VSS.n9752 VSS.n9649 0.0206923
R18203 VSS.n9864 VSS.n178 0.0206923
R18204 VSS.n1260 VSS.n455 0.0206923
R18205 VSS.n634 VSS.n499 0.0206923
R18206 VSS.n10015 VSS.n9934 0.0206923
R18207 VSS.n9993 VSS.n9954 0.0206923
R18208 VSS.n11195 VSS.n11194 0.0206923
R18209 VSS.n9626 VSS.n9625 0.0206923
R18210 VSS.n10677 VSS.n10676 0.0206172
R18211 VSS.n10687 VSS.n10291 0.0206172
R18212 VSS.n786 VSS.n785 0.0205874
R18213 VSS.n9730 VSS.n9693 0.0205874
R18214 VSS.n9842 VSS.n9841 0.0205874
R18215 VSS.n10015 VSS.n578 0.0205874
R18216 VSS.n9626 VSS.n804 0.0205874
R18217 VSS.n9752 VSS.n9661 0.0205874
R18218 VSS.n10048 VSS.n546 0.0205874
R18219 VSS.n9730 VSS.n9717 0.0205874
R18220 VSS.n590 VSS.n184 0.0205874
R18221 VSS.n11051 VSS.n11050 0.0205874
R18222 VSS.n9993 VSS.n9966 0.0205874
R18223 VSS.n9602 VSS.n9601 0.0205874
R18224 VSS.n10439 VSS.n10438 0.0204409
R18225 VSS.n11330 VSS.n11329 0.0203634
R18226 VSS.n70 VSS.n69 0.0203634
R18227 VSS.n10284 VSS.n10283 0.0201097
R18228 VSS.n9095 VSS.n9094 0.01994
R18229 VSS.n9008 VSS.n9007 0.01994
R18230 VSS.n10927 VSS.n10926 0.01994
R18231 VSS.n868 VSS.n866 0.01994
R18232 VSS.n1126 VSS.n1125 0.01994
R18233 VSS.n1114 VSS.n1113 0.01994
R18234 VSS.n1093 VSS.n1092 0.01994
R18235 VSS.n1077 VSS.n1076 0.01994
R18236 VSS.n1056 VSS.n1055 0.01994
R18237 VSS.n1044 VSS.n1043 0.01994
R18238 VSS.n1019 VSS.n1018 0.01994
R18239 VSS.n1007 VSS.n1006 0.01994
R18240 VSS.n986 VSS.n985 0.01994
R18241 VSS.n970 VSS.n969 0.01994
R18242 VSS.n10985 VSS.n10984 0.01994
R18243 VSS.n11359 VSS.n11358 0.01994
R18244 VSS.n11347 VSS.n11345 0.01994
R18245 VSS.n11377 VSS.n11376 0.01994
R18246 VSS.n11364 VSS.n11363 0.01994
R18247 VSS.n10980 VSS.n10979 0.01994
R18248 VSS.n10932 VSS.n10931 0.01994
R18249 VSS.n1205 VSS.n1204 0.01994
R18250 VSS.n9543 VSS.n9542 0.01994
R18251 VSS.n9530 VSS.n9529 0.01994
R18252 VSS.n9420 VSS.n9419 0.01994
R18253 VSS.n9350 VSS.n9349 0.01994
R18254 VSS.n9297 VSS.n9296 0.01994
R18255 VSS.n9252 VSS.n9251 0.01994
R18256 VSS.n9175 VSS.n9174 0.01994
R18257 VSS.n1547 VSS.n1546 0.01994
R18258 VSS.n11334 VSS.n11333 0.0196517
R18259 VSS.n11332 VSS.n11331 0.0196517
R18260 VSS.n11329 VSS.n11328 0.0196517
R18261 VSS.n11327 VSS.n11326 0.0196517
R18262 VSS.n66 VSS.n65 0.0196517
R18263 VSS.n69 VSS.n67 0.0196517
R18264 VSS.n73 VSS.n72 0.0196517
R18265 VSS.n76 VSS.n74 0.0196517
R18266 VSS.n9080 VSS.n9079 0.0194273
R18267 VSS.n9105 VSS.n9103 0.0194273
R18268 VSS.n858 VSS.n857 0.0194273
R18269 VSS.n1104 VSS.n1103 0.0194273
R18270 VSS.n1279 VSS.n1278 0.0194273
R18271 VSS.n924 VSS.n923 0.0194273
R18272 VSS.n381 VSS.n380 0.0194273
R18273 VSS.n997 VSS.n996 0.0194273
R18274 VSS.n297 VSS.n296 0.0194273
R18275 VSS.n11063 VSS.n11060 0.0194273
R18276 VSS.n11211 VSS.n11209 0.0194273
R18277 VSS.n1195 VSS.n1194 0.0194273
R18278 VSS.n9395 VSS.n9392 0.0194273
R18279 VSS.n9410 VSS.n9409 0.0194273
R18280 VSS.n9237 VSS.n9236 0.0194273
R18281 VSS.n9225 VSS.n9223 0.0194273
R18282 VSS.n1573 VSS.n1572 0.019407
R18283 VSS.n1576 VSS.n1575 0.019407
R18284 VSS.n1579 VSS.n1577 0.019407
R18285 VSS.n8958 VSS.n8957 0.019407
R18286 VSS.n8961 VSS.n8959 0.019407
R18287 VSS.n8964 VSS.n8962 0.019407
R18288 VSS.n963 VSS.n962 0.019407
R18289 VSS.n961 VSS.n960 0.019407
R18290 VSS.n959 VSS.n958 0.019407
R18291 VSS.n10283 VSS.n10282 0.019407
R18292 VSS.n10281 VSS.n10280 0.019407
R18293 VSS.n10279 VSS.n10278 0.019407
R18294 VSS.n9445 VSS.n9444 0.0192683
R18295 VSS.n9436 VSS.n9435 0.0192683
R18296 VSS.n8983 VSS.n8980 0.0189267
R18297 VSS.n8998 VSS.n8997 0.0189267
R18298 VSS.n1138 VSS.n1135 0.0189267
R18299 VSS.n911 VSS.n910 0.0189267
R18300 VSS.n10137 VSS.n10136 0.0189267
R18301 VSS.n1030 VSS.n1029 0.0189267
R18302 VSS.n10197 VSS.n10196 0.0189267
R18303 VSS.n950 VSS.n949 0.0189267
R18304 VSS.n10257 VSS.n10256 0.0189267
R18305 VSS.n11006 VSS.n11003 0.0189267
R18306 VSS.n10970 VSS.n10969 0.0189267
R18307 VSS.n9553 VSS.n9551 0.0189267
R18308 VSS.n9372 VSS.n9371 0.0189267
R18309 VSS.n9360 VSS.n9358 0.0189267
R18310 VSS.n9150 VSS.n9147 0.0189267
R18311 VSS.n9165 VSS.n9164 0.0189267
R18312 VSS VSS.n10823 0.0186978
R18313 VSS.n111 VSS.n110 0.0186448
R18314 VSS.n107 VSS.n106 0.0186448
R18315 VSS.n11385 VSS.n83 0.0186448
R18316 VSS.n83 VSS.n82 0.0186448
R18317 VSS.n11388 VSS.n79 0.0186448
R18318 VSS.n11397 VSS.n56 0.0186448
R18319 VSS.n11394 VSS.n55 0.0186448
R18320 VSS.n37 VSS.n30 0.0186448
R18321 VSS.n33 VSS.n30 0.0186448
R18322 VSS.n35 VSS.n29 0.0186448
R18323 VSS.n10704 VSS.n10702 0.0186448
R18324 VSS.n10704 VSS.n10699 0.0186448
R18325 VSS.n10705 VSS.n10700 0.0186448
R18326 VSS.n11307 VSS.n11306 0.0186448
R18327 VSS.n11307 VSS.n126 0.0186448
R18328 VSS.n11312 VSS.n11311 0.0186448
R18329 VSS.n10564 VSS.n10557 0.0186448
R18330 VSS.n10568 VSS.n10557 0.0186448
R18331 VSS.n10569 VSS.n10562 0.0186448
R18332 VSS.n10568 VSS.n10563 0.0186448
R18333 VSS.n10566 VSS.n10562 0.0186448
R18334 VSS.n10571 VSS.n10564 0.0186448
R18335 VSS.n230 VSS.n226 0.0186448
R18336 VSS.n10911 VSS.n225 0.0186448
R18337 VSS.n230 VSS.n229 0.0186448
R18338 VSS.n10912 VSS.n10911 0.0186448
R18339 VSS.n227 VSS.n226 0.0186448
R18340 VSS.n108 VSS.n107 0.0186448
R18341 VSS.n110 VSS.n109 0.0186448
R18342 VSS.n37 VSS.n32 0.0186448
R18343 VSS.n11432 VSS.n33 0.0186448
R18344 VSS.n11430 VSS.n29 0.0186448
R18345 VSS.n11396 VSS.n55 0.0186448
R18346 VSS.n11397 VSS.n58 0.0186448
R18347 VSS.n11386 VSS.n11385 0.0186448
R18348 VSS.n11383 VSS.n79 0.0186448
R18349 VSS.n82 VSS.n62 0.0186448
R18350 VSS.n11311 VSS.n124 0.0186448
R18351 VSS.n126 VSS.n122 0.0186448
R18352 VSS.n11309 VSS.n11306 0.0186448
R18353 VSS.n10729 VSS.n10700 0.0186448
R18354 VSS.n10707 VSS.n10699 0.0186448
R18355 VSS.n10731 VSS.n10702 0.0186448
R18356 VSS.n9077 VSS.n9076 0.0184746
R18357 VSS.n9107 VSS.n9106 0.0184746
R18358 VSS.n855 VSS.n854 0.0184746
R18359 VSS.n848 VSS.n847 0.0184746
R18360 VSS.n1101 VSS.n1100 0.0184746
R18361 VSS.n1275 VSS.n1274 0.0184746
R18362 VSS.n921 VSS.n920 0.0184746
R18363 VSS.n377 VSS.n376 0.0184746
R18364 VSS.n994 VSS.n993 0.0184746
R18365 VSS.n293 VSS.n292 0.0184746
R18366 VSS.n11065 VSS.n11064 0.0184746
R18367 VSS.n11074 VSS.n11073 0.0184746
R18368 VSS.n11220 VSS.n11219 0.0184746
R18369 VSS.n11213 VSS.n11212 0.0184746
R18370 VSS.n1170 VSS.n1169 0.0184746
R18371 VSS.n1191 VSS.n1190 0.0184746
R18372 VSS.n9397 VSS.n9396 0.0184746
R18373 VSS.n9406 VSS.n9405 0.0184746
R18374 VSS.n9234 VSS.n9233 0.0184746
R18375 VSS.n9227 VSS.n9226 0.0184746
R18376 VSS.n898 VSS.n897 0.0183443
R18377 VSS.n1067 VSS.n1066 0.0183443
R18378 VSS.n10169 VSS.n10167 0.0183443
R18379 VSS.n937 VSS.n936 0.0183443
R18380 VSS.n10229 VSS.n10227 0.0183443
R18381 VSS.n10909 VSS.n10908 0.0183443
R18382 VSS.n713 VSS.n711 0.0183443
R18383 VSS.n1227 VSS.n1225 0.0183443
R18384 VSS.n9272 VSS.n9269 0.0183443
R18385 VSS.n9287 VSS.n9286 0.0183443
R18386 VSS.n9054 VSS.n9053 0.0183443
R18387 VSS.n9127 VSS.n9126 0.0183443
R18388 VSS.n9069 VSS.n9068 0.0183136
R18389 VSS.n9089 VSS.n9044 0.0183136
R18390 VSS.n9015 VSS.n1561 0.0183136
R18391 VSS.n1289 VSS.n1288 0.0183136
R18392 VSS.n10153 VSS.n10152 0.0183136
R18393 VSS.n391 VSS.n390 0.0183136
R18394 VSS.n370 VSS.n369 0.0183136
R18395 VSS.n10213 VSS.n10212 0.0183136
R18396 VSS.n319 VSS.n318 0.0183136
R18397 VSS.n307 VSS.n306 0.0183136
R18398 VSS.n10273 VSS.n10272 0.0183136
R18399 VSS.n9382 VSS.n9380 0.0183136
R18400 VSS.n9344 VSS.n9320 0.0183136
R18401 VSS.n9309 VSS.n1505 0.0183136
R18402 VSS.n9246 VSS.n9211 0.0183136
R18403 VSS.n9182 VSS.n1523 0.0183136
R18404 VSS.n10060 VSS.n536 0.0182205
R18405 VSS.n11078 VSS.n11077 0.0182205
R18406 VSS.n11223 VSS.n11222 0.0182205
R18407 VSS.n9823 VSS.n768 0.0182205
R18408 VSS.n9467 VSS.n1380 0.0181966
R18409 VSS.n10771 VSS.n10770 0.0181748
R18410 VSS.n9463 VSS.n9452 0.0180195
R18411 VSS.n958 VSS.n253 0.0180018
R18412 VSS.n8985 VSS.n8984 0.0179991
R18413 VSS.n8994 VSS.n8993 0.0179991
R18414 VSS.n1140 VSS.n1139 0.0179991
R18415 VSS.n1149 VSS.n1148 0.0179991
R18416 VSS.n908 VSS.n907 0.0179991
R18417 VSS.n10133 VSS.n10132 0.0179991
R18418 VSS.n1027 VSS.n1026 0.0179991
R18419 VSS.n10193 VSS.n10192 0.0179991
R18420 VSS.n947 VSS.n946 0.0179991
R18421 VSS.n10253 VSS.n10252 0.0179991
R18422 VSS.n11008 VSS.n11007 0.0179991
R18423 VSS.n11017 VSS.n11016 0.0179991
R18424 VSS.n10957 VSS.n10956 0.0179991
R18425 VSS.n10966 VSS.n10965 0.0179991
R18426 VSS.n1155 VSS.n1154 0.0179991
R18427 VSS.n9555 VSS.n9554 0.0179991
R18428 VSS.n9369 VSS.n9368 0.0179991
R18429 VSS.n9362 VSS.n9361 0.0179991
R18430 VSS.n9152 VSS.n9151 0.0179991
R18431 VSS.n9161 VSS.n9160 0.0179991
R18432 VSS.n1147 VSS.n491 0.0177518
R18433 VSS.n11022 VSS.n11020 0.0177518
R18434 VSS.n10955 VSS.n151 0.0177518
R18435 VSS.n9781 VSS.n793 0.0177518
R18436 VSS.n2253 VSS.n61 0.01775
R18437 VSS.n895 VSS.n894 0.0174461
R18438 VSS.n888 VSS.n887 0.0174461
R18439 VSS.n1064 VSS.n1063 0.0174461
R18440 VSS.n10171 VSS.n10170 0.0174461
R18441 VSS.n934 VSS.n933 0.0174461
R18442 VSS.n10231 VSS.n10230 0.0174461
R18443 VSS.n10906 VSS.n10905 0.0174461
R18444 VSS.n10899 VSS.n10898 0.0174461
R18445 VSS.n722 VSS.n721 0.0174461
R18446 VSS.n715 VSS.n714 0.0174461
R18447 VSS.n1435 VSS.n1434 0.0174461
R18448 VSS.n1229 VSS.n1228 0.0174461
R18449 VSS.n9274 VSS.n9273 0.0174461
R18450 VSS.n9283 VSS.n9282 0.0174461
R18451 VSS.n9051 VSS.n9050 0.0174461
R18452 VSS.n9123 VSS.n9122 0.0174461
R18453 VSS.n9443 VSS.n9442 0.0174024
R18454 VSS.n9438 VSS.n9437 0.0174024
R18455 VSS.n10757 VSS.n10740 0.0173337
R18456 VSS.n10755 VSS.n10740 0.0173337
R18457 VSS.n886 VSS.n448 0.0172066
R18458 VSS.n10897 VSS.n10895 0.0172066
R18459 VSS.n725 VSS.n724 0.0172066
R18460 VSS.n1438 VSS.n1437 0.0172066
R18461 VSS.n1386 VSS.n811 0.0169894
R18462 VSS.n1332 VSS.n1327 0.0169894
R18463 VSS.n10759 VSS.n10758 0.0169128
R18464 VSS.n1408 VSS.n814 0.0167766
R18465 VSS.n9511 VSS.n9510 0.0167766
R18466 VSS.n9446 VSS.n9445 0.0167439
R18467 VSS.n9444 VSS.n9424 0.0167439
R18468 VSS.n9443 VSS.n9424 0.0167439
R18469 VSS.n9442 VSS.n9425 0.0167439
R18470 VSS.n9441 VSS.n9425 0.0167439
R18471 VSS.n9439 VSS.n9426 0.0167439
R18472 VSS.n9438 VSS.n9426 0.0167439
R18473 VSS.n9437 VSS.n9427 0.0167439
R18474 VSS.n9436 VSS.n9427 0.0167439
R18475 VSS.n9435 VSS.n9428 0.0167439
R18476 VSS.n10726 VSS.n10708 0.0167142
R18477 VSS.n10725 VSS.n10708 0.0167142
R18478 VSS.n10724 VSS.n10709 0.0167142
R18479 VSS.n10723 VSS.n10709 0.0167142
R18480 VSS.n10722 VSS.n10710 0.0167142
R18481 VSS.n10721 VSS.n10710 0.0167142
R18482 VSS.n10719 VSS.n10711 0.0167142
R18483 VSS.n10718 VSS.n10711 0.0167142
R18484 VSS.n1387 VSS.n814 0.0166702
R18485 VSS.n9511 VSS.n1333 0.0166702
R18486 VSS.n10677 VSS.n10335 0.016599
R18487 VSS.n9648 VSS.n9647 0.0164965
R18488 VSS.n9646 VSS.n9645 0.0164965
R18489 VSS.n9644 VSS.n9643 0.0164965
R18490 VSS.n780 VSS.n779 0.0164965
R18491 VSS.n782 VSS.n781 0.0164965
R18492 VSS.n784 VSS.n783 0.0164965
R18493 VSS.n662 VSS.n661 0.0164965
R18494 VSS.n664 VSS.n663 0.0164965
R18495 VSS.n666 VSS.n665 0.0164965
R18496 VSS.n9870 VSS.n9869 0.0164965
R18497 VSS.n9868 VSS.n9867 0.0164965
R18498 VSS.n9866 VSS.n9865 0.0164965
R18499 VSS.n1262 VSS.n1261 0.0164965
R18500 VSS.n1264 VSS.n1263 0.0164965
R18501 VSS.n1266 VSS.n1265 0.0164965
R18502 VSS.n1246 VSS.n1245 0.0164965
R18503 VSS.n1244 VSS.n1243 0.0164965
R18504 VSS.n1242 VSS.n1241 0.0164965
R18505 VSS.n636 VSS.n635 0.0164965
R18506 VSS.n638 VSS.n637 0.0164965
R18507 VSS.n640 VSS.n639 0.0164965
R18508 VSS.n9656 VSS.n9655 0.0164965
R18509 VSS.n9658 VSS.n9657 0.0164965
R18510 VSS.n9660 VSS.n9659 0.0164965
R18511 VSS.n592 VSS.n591 0.0164965
R18512 VSS.n594 VSS.n593 0.0164965
R18513 VSS.n596 VSS.n595 0.0164965
R18514 VSS.n9929 VSS.n9928 0.0164965
R18515 VSS.n9931 VSS.n9930 0.0164965
R18516 VSS.n9933 VSS.n9932 0.0164965
R18517 VSS.n11049 VSS.n11048 0.0164965
R18518 VSS.n11047 VSS.n11046 0.0164965
R18519 VSS.n11045 VSS.n11044 0.0164965
R18520 VSS.n9949 VSS.n9948 0.0164965
R18521 VSS.n9951 VSS.n9950 0.0164965
R18522 VSS.n9953 VSS.n9952 0.0164965
R18523 VSS.n9965 VSS.n9964 0.0164965
R18524 VSS.n9963 VSS.n9962 0.0164965
R18525 VSS.n9961 VSS.n9960 0.0164965
R18526 VSS.n11189 VSS.n11188 0.0164965
R18527 VSS.n11191 VSS.n11190 0.0164965
R18528 VSS.n11193 VSS.n11192 0.0164965
R18529 VSS.n9624 VSS.n9623 0.0164965
R18530 VSS.n9622 VSS.n9621 0.0164965
R18531 VSS.n9620 VSS.n9619 0.0164965
R18532 VSS.n9608 VSS.n9607 0.0164965
R18533 VSS.n9606 VSS.n9605 0.0164965
R18534 VSS.n9604 VSS.n9603 0.0164965
R18535 VSS.n9480 VSS.n811 0.0164574
R18536 VSS.n1327 VSS.n1326 0.0164574
R18537 VSS.n10754 VSS.n10753 0.0164441
R18538 VSS.n9691 VSS.n9690 0.0163916
R18539 VSS.n9688 VSS.n9687 0.0163916
R18540 VSS.n9685 VSS.n9684 0.0163916
R18541 VSS.n9851 VSS.n9850 0.0163916
R18542 VSS.n9848 VSS.n9847 0.0163916
R18543 VSS.n9845 VSS.n9844 0.0163916
R18544 VSS.n606 VSS.n605 0.0163916
R18545 VSS.n611 VSS.n610 0.0163916
R18546 VSS.n616 VSS.n615 0.0163916
R18547 VSS.n9703 VSS.n9702 0.0163916
R18548 VSS.n9708 VSS.n9707 0.0163916
R18549 VSS.n9713 VSS.n9712 0.0163916
R18550 VSS.n10743 VSS.n10742 0.0160769
R18551 VSS.n10497 VSS.n10496 0.0160245
R18552 VSS.n10495 VSS.n10494 0.0160245
R18553 VSS.n10606 VSS.n10605 0.0160245
R18554 VSS.n10608 VSS.n10607 0.0160245
R18555 VSS.n9649 VSS.n9639 0.0160245
R18556 VSS.n9648 VSS.n9639 0.0160245
R18557 VSS.n9647 VSS.n9640 0.0160245
R18558 VSS.n9646 VSS.n9640 0.0160245
R18559 VSS.n9645 VSS.n9641 0.0160245
R18560 VSS.n9644 VSS.n9641 0.0160245
R18561 VSS.n9643 VSS.n9642 0.0160245
R18562 VSS.n9642 VSS.n649 0.0160245
R18563 VSS.n9885 VSS.n647 0.0160245
R18564 VSS.n778 VSS.n777 0.0160245
R18565 VSS.n779 VSS.n777 0.0160245
R18566 VSS.n780 VSS.n776 0.0160245
R18567 VSS.n781 VSS.n776 0.0160245
R18568 VSS.n782 VSS.n775 0.0160245
R18569 VSS.n783 VSS.n775 0.0160245
R18570 VSS.n784 VSS.n774 0.0160245
R18571 VSS.n785 VSS.n774 0.0160245
R18572 VSS.n660 VSS.n578 0.0160245
R18573 VSS.n661 VSS.n660 0.0160245
R18574 VSS.n662 VSS.n659 0.0160245
R18575 VSS.n663 VSS.n659 0.0160245
R18576 VSS.n664 VSS.n658 0.0160245
R18577 VSS.n665 VSS.n658 0.0160245
R18578 VSS.n666 VSS.n657 0.0160245
R18579 VSS.n667 VSS.n657 0.0160245
R18580 VSS.n673 VSS.n672 0.0160245
R18581 VSS.n9871 VSS.n9860 0.0160245
R18582 VSS.n9870 VSS.n9860 0.0160245
R18583 VSS.n9869 VSS.n9861 0.0160245
R18584 VSS.n9868 VSS.n9861 0.0160245
R18585 VSS.n9867 VSS.n9862 0.0160245
R18586 VSS.n9866 VSS.n9862 0.0160245
R18587 VSS.n9865 VSS.n9863 0.0160245
R18588 VSS.n9864 VSS.n9863 0.0160245
R18589 VSS.n1260 VSS.n1259 0.0160245
R18590 VSS.n1261 VSS.n1259 0.0160245
R18591 VSS.n1262 VSS.n1258 0.0160245
R18592 VSS.n1263 VSS.n1258 0.0160245
R18593 VSS.n1264 VSS.n1257 0.0160245
R18594 VSS.n1265 VSS.n1257 0.0160245
R18595 VSS.n1266 VSS.n1256 0.0160245
R18596 VSS.n1267 VSS.n1256 0.0160245
R18597 VSS.n9519 VSS.n1236 0.0160245
R18598 VSS.n1247 VSS.n1237 0.0160245
R18599 VSS.n1246 VSS.n1237 0.0160245
R18600 VSS.n1245 VSS.n1238 0.0160245
R18601 VSS.n1244 VSS.n1238 0.0160245
R18602 VSS.n1243 VSS.n1239 0.0160245
R18603 VSS.n1242 VSS.n1239 0.0160245
R18604 VSS.n1241 VSS.n1240 0.0160245
R18605 VSS.n1240 VSS.n804 0.0160245
R18606 VSS.n634 VSS.n633 0.0160245
R18607 VSS.n635 VSS.n633 0.0160245
R18608 VSS.n636 VSS.n632 0.0160245
R18609 VSS.n637 VSS.n632 0.0160245
R18610 VSS.n638 VSS.n631 0.0160245
R18611 VSS.n639 VSS.n631 0.0160245
R18612 VSS.n640 VSS.n630 0.0160245
R18613 VSS.n641 VSS.n630 0.0160245
R18614 VSS.n9894 VSS.n643 0.0160245
R18615 VSS.n9654 VSS.n9653 0.0160245
R18616 VSS.n9655 VSS.n9653 0.0160245
R18617 VSS.n9656 VSS.n9652 0.0160245
R18618 VSS.n9657 VSS.n9652 0.0160245
R18619 VSS.n9658 VSS.n9651 0.0160245
R18620 VSS.n9659 VSS.n9651 0.0160245
R18621 VSS.n9660 VSS.n9650 0.0160245
R18622 VSS.n9661 VSS.n9650 0.0160245
R18623 VSS.n590 VSS.n589 0.0160245
R18624 VSS.n591 VSS.n589 0.0160245
R18625 VSS.n592 VSS.n588 0.0160245
R18626 VSS.n593 VSS.n588 0.0160245
R18627 VSS.n594 VSS.n587 0.0160245
R18628 VSS.n595 VSS.n587 0.0160245
R18629 VSS.n596 VSS.n586 0.0160245
R18630 VSS.n597 VSS.n586 0.0160245
R18631 VSS.n9915 VSS.n583 0.0160245
R18632 VSS.n9927 VSS.n582 0.0160245
R18633 VSS.n9928 VSS.n582 0.0160245
R18634 VSS.n9929 VSS.n581 0.0160245
R18635 VSS.n9930 VSS.n581 0.0160245
R18636 VSS.n9931 VSS.n580 0.0160245
R18637 VSS.n9932 VSS.n580 0.0160245
R18638 VSS.n9933 VSS.n579 0.0160245
R18639 VSS.n9934 VSS.n579 0.0160245
R18640 VSS.n11050 VSS.n11039 0.0160245
R18641 VSS.n11049 VSS.n11039 0.0160245
R18642 VSS.n11048 VSS.n11040 0.0160245
R18643 VSS.n11047 VSS.n11040 0.0160245
R18644 VSS.n11046 VSS.n11041 0.0160245
R18645 VSS.n11045 VSS.n11041 0.0160245
R18646 VSS.n11044 VSS.n11042 0.0160245
R18647 VSS.n11043 VSS.n11042 0.0160245
R18648 VSS.n11283 VSS.n11282 0.0160245
R18649 VSS.n9947 VSS.n9946 0.0160245
R18650 VSS.n9948 VSS.n9946 0.0160245
R18651 VSS.n9949 VSS.n9945 0.0160245
R18652 VSS.n9950 VSS.n9945 0.0160245
R18653 VSS.n9951 VSS.n9944 0.0160245
R18654 VSS.n9952 VSS.n9944 0.0160245
R18655 VSS.n9953 VSS.n9943 0.0160245
R18656 VSS.n9954 VSS.n9943 0.0160245
R18657 VSS.n9966 VSS.n9955 0.0160245
R18658 VSS.n9965 VSS.n9955 0.0160245
R18659 VSS.n9964 VSS.n9956 0.0160245
R18660 VSS.n9963 VSS.n9956 0.0160245
R18661 VSS.n9962 VSS.n9957 0.0160245
R18662 VSS.n9961 VSS.n9957 0.0160245
R18663 VSS.n9960 VSS.n9958 0.0160245
R18664 VSS.n9959 VSS.n9958 0.0160245
R18665 VSS.n142 VSS.n141 0.0160245
R18666 VSS.n11187 VSS.n11186 0.0160245
R18667 VSS.n11188 VSS.n11186 0.0160245
R18668 VSS.n11189 VSS.n11185 0.0160245
R18669 VSS.n11190 VSS.n11185 0.0160245
R18670 VSS.n11191 VSS.n11184 0.0160245
R18671 VSS.n11192 VSS.n11184 0.0160245
R18672 VSS.n11193 VSS.n11183 0.0160245
R18673 VSS.n11194 VSS.n11183 0.0160245
R18674 VSS.n9625 VSS.n806 0.0160245
R18675 VSS.n9624 VSS.n806 0.0160245
R18676 VSS.n9623 VSS.n807 0.0160245
R18677 VSS.n9622 VSS.n807 0.0160245
R18678 VSS.n9621 VSS.n808 0.0160245
R18679 VSS.n9620 VSS.n808 0.0160245
R18680 VSS.n9619 VSS.n809 0.0160245
R18681 VSS.n9618 VSS.n809 0.0160245
R18682 VSS.n1233 VSS.n810 0.0160245
R18683 VSS.n9609 VSS.n823 0.0160245
R18684 VSS.n9608 VSS.n823 0.0160245
R18685 VSS.n9607 VSS.n824 0.0160245
R18686 VSS.n9606 VSS.n824 0.0160245
R18687 VSS.n9605 VSS.n825 0.0160245
R18688 VSS.n9604 VSS.n825 0.0160245
R18689 VSS.n9603 VSS.n826 0.0160245
R18690 VSS.n9602 VSS.n826 0.0160245
R18691 VSS.n10824 VSS 0.0159286
R18692 VSS.n9672 VSS.n9671 0.0159196
R18693 VSS.n9692 VSS.n9673 0.0159196
R18694 VSS.n9675 VSS.n9674 0.0159196
R18695 VSS.n9689 VSS.n9676 0.0159196
R18696 VSS.n9678 VSS.n9677 0.0159196
R18697 VSS.n9686 VSS.n9679 0.0159196
R18698 VSS.n9681 VSS.n9680 0.0159196
R18699 VSS.n9683 VSS.n9682 0.0159196
R18700 VSS.n681 VSS.n680 0.0159196
R18701 VSS.n9852 VSS.n682 0.0159196
R18702 VSS.n684 VSS.n683 0.0159196
R18703 VSS.n9849 VSS.n685 0.0159196
R18704 VSS.n687 VSS.n686 0.0159196
R18705 VSS.n9846 VSS.n688 0.0159196
R18706 VSS.n690 VSS.n689 0.0159196
R18707 VSS.n9843 VSS.n691 0.0159196
R18708 VSS.n604 VSS.n603 0.0159196
R18709 VSS.n602 VSS.n601 0.0159196
R18710 VSS.n609 VSS.n608 0.0159196
R18711 VSS.n607 VSS.n600 0.0159196
R18712 VSS.n614 VSS.n613 0.0159196
R18713 VSS.n612 VSS.n599 0.0159196
R18714 VSS.n619 VSS.n618 0.0159196
R18715 VSS.n617 VSS.n598 0.0159196
R18716 VSS.n9701 VSS.n9700 0.0159196
R18717 VSS.n9699 VSS.n9697 0.0159196
R18718 VSS.n9706 VSS.n9705 0.0159196
R18719 VSS.n9704 VSS.n9696 0.0159196
R18720 VSS.n9711 VSS.n9710 0.0159196
R18721 VSS.n9709 VSS.n9695 0.0159196
R18722 VSS.n9716 VSS.n9715 0.0159196
R18723 VSS.n9714 VSS.n9694 0.0159196
R18724 VSS.n10439 VSS.n10335 0.0158871
R18725 VSS.n10587 VSS.n10586 0.0157873
R18726 VSS.n10814 VSS.n250 0.0156685
R18727 VSS.n10783 VSS.n10782 0.0156685
R18728 VSS.n10717 VSS.n10712 0.0156595
R18729 VSS.n9887 VSS.n9886 0.0156049
R18730 VSS.n671 VSS.n668 0.0156049
R18731 VSS.n9521 VSS.n9520 0.0156049
R18732 VSS.n9893 VSS.n9892 0.0156049
R18733 VSS.n9917 VSS.n9916 0.0156049
R18734 VSS.n11284 VSS.n11281 0.0156049
R18735 VSS.n143 VSS.n140 0.0156049
R18736 VSS.n1234 VSS.n815 0.0156049
R18737 VSS.n1177 VSS.n1176 0.0155
R18738 VSS.n1180 VSS.n1179 0.0155
R18739 VSS.n623 VSS.n622 0.0155
R18740 VSS.n9905 VSS.n626 0.0155
R18741 VSS.n11470 VSS.n3 0.0152621
R18742 VSS.n8955 VSS.n8954 0.0152551
R18743 VSS.n9094 VSS.n1554 0.01514
R18744 VSS.n9008 VSS.n8969 0.01514
R18745 VSS.n10927 VSS.n221 0.01514
R18746 VSS.n869 VSS.n868 0.01514
R18747 VSS.n1125 VSS.n1124 0.01514
R18748 VSS.n1113 VSS.n1112 0.01514
R18749 VSS.n1092 VSS.n1091 0.01514
R18750 VSS.n1076 VSS.n1075 0.01514
R18751 VSS.n1055 VSS.n1054 0.01514
R18752 VSS.n1043 VSS.n1042 0.01514
R18753 VSS.n1018 VSS.n1017 0.01514
R18754 VSS.n1006 VSS.n1005 0.01514
R18755 VSS.n985 VSS.n984 0.01514
R18756 VSS.n969 VSS.n968 0.01514
R18757 VSS.n10984 VSS.n207 0.01514
R18758 VSS.n11359 VSS.n96 0.01514
R18759 VSS.n11348 VSS.n11347 0.01514
R18760 VSS.n11376 VSS.n11374 0.01514
R18761 VSS.n11363 VSS.n90 0.01514
R18762 VSS.n10980 VSS.n10942 0.01514
R18763 VSS.n10931 VSS.n214 0.01514
R18764 VSS.n1206 VSS.n1205 0.01514
R18765 VSS.n9542 VSS.n9540 0.01514
R18766 VSS.n9529 VSS.n1221 0.01514
R18767 VSS.n9420 VSS.n1396 0.01514
R18768 VSS.n9349 VSS.n1496 0.01514
R18769 VSS.n9297 VSS.n9262 0.01514
R18770 VSS.n9251 VSS.n1513 0.01514
R18771 VSS.n9175 VSS.n9136 0.01514
R18772 VSS.n1548 VSS.n1547 0.01514
R18773 VSS.n9110 VSS.n9109 0.0150766
R18774 VSS.n853 VSS.n851 0.0150766
R18775 VSS.n10121 VSS.n427 0.0150766
R18776 VSS.n10181 VSS.n357 0.0150766
R18777 VSS.n10241 VSS.n285 0.0150766
R18778 VSS.n11069 VSS.n11068 0.0150766
R18779 VSS.n11216 VSS.n11215 0.0150766
R18780 VSS.n1189 VSS.n1186 0.0150766
R18781 VSS.n9404 VSS.n9401 0.0150766
R18782 VSS.n9230 VSS.n9229 0.0150766
R18783 VSS.n8992 VSS.n8989 0.014691
R18784 VSS.n1152 VSS.n1143 0.014691
R18785 VSS.n10128 VSS.n419 0.014691
R18786 VSS.n10188 VSS.n347 0.014691
R18787 VSS.n10248 VSS.n275 0.014691
R18788 VSS.n11012 VSS.n11011 0.014691
R18789 VSS.n10964 VSS.n10961 0.014691
R18790 VSS.n9558 VSS.n9557 0.014691
R18791 VSS.n9365 VSS.n9364 0.014691
R18792 VSS.n9159 VSS.n9156 0.014691
R18793 VSS.n78 VSS.n77 0.014605
R18794 VSS.n10716 VSS.n10712 0.0144843
R18795 VSS.n10715 VSS.n10713 0.0144843
R18796 VSS.n10714 VSS.n10713 0.0144843
R18797 VSS.n893 VSS.n891 0.0142425
R18798 VSS.n10174 VSS.n397 0.0142425
R18799 VSS.n10234 VSS.n325 0.0142425
R18800 VSS.n10904 VSS.n10902 0.0142425
R18801 VSS.n718 VSS.n717 0.0142425
R18802 VSS.n1232 VSS.n1231 0.0142425
R18803 VSS.n9281 VSS.n9278 0.0142425
R18804 VSS.n9121 VSS.n9118 0.0142425
R18805 VSS.n9038 VSS.n1560 0.0141709
R18806 VSS.n10144 VSS.n10142 0.0141709
R18807 VSS.n10204 VSS.n10202 0.0141709
R18808 VSS.n10264 VSS.n10262 0.0141709
R18809 VSS.n9336 VSS.n1478 0.0141709
R18810 VSS.n9205 VSS.n1522 0.0141709
R18811 VSS.n9629 VSS.n9628 0.0139852
R18812 VSS.n9755 VSS.n9754 0.0139852
R18813 VSS.n9750 VSS.n9749 0.0139852
R18814 VSS.n9733 VSS.n9732 0.0139852
R18815 VSS.n9728 VSS.n9727 0.0139852
R18816 VSS.n10013 VSS.n10012 0.0139852
R18817 VSS.n9996 VSS.n9995 0.0139852
R18818 VSS.n9991 VSS.n9990 0.0139852
R18819 VSS.n10634 VSS.n10633 0.0137679
R18820 VSS.n10748 VSS.n250 0.0136461
R18821 VSS.n10782 VSS.n10781 0.0136461
R18822 VSS.n11436 VSS.n11435 0.0133485
R18823 VSS.n11403 VSS.n11402 0.0133485
R18824 VSS.n11427 VSS.n11426 0.0132877
R18825 VSS.n9032 VSS.n9018 0.0132388
R18826 VSS.n10145 VSS.n403 0.0132388
R18827 VSS.n10205 VSS.n331 0.0132388
R18828 VSS.n10265 VSS.n259 0.0132388
R18829 VSS.n9337 VSS.n9322 0.0132388
R18830 VSS.n9199 VSS.n9185 0.0132388
R18831 VSS.n1363 VSS.n1362 0.013182
R18832 VSS.n9760 VSS.n9759 0.013182
R18833 VSS.n9738 VSS.n9737 0.013182
R18834 VSS.n10001 VSS.n10000 0.013182
R18835 VSS.n9979 VSS.n9978 0.013182
R18836 VSS.n8976 VSS.n8972 0.0127708
R18837 VSS.n874 VSS.n870 0.0127708
R18838 VSS.n1088 VSS.n904 0.0127708
R18839 VSS.n1039 VSS.n928 0.0127708
R18840 VSS.n981 VSS.n943 0.0127708
R18841 VSS.n10995 VSS.n10991 0.0127708
R18842 VSS.n10949 VSS.n10945 0.0127708
R18843 VSS.n1211 VSS.n1207 0.0127708
R18844 VSS.n1491 VSS.n1487 0.0127708
R18845 VSS.n9143 VSS.n9139 0.0127708
R18846 VSS.n9508 VSS.n1335 0.012534
R18847 VSS.n9493 VSS.n1374 0.0123788
R18848 VSS.n9974 VSS.n31 0.0123788
R18849 VSS.n1374 VSS.n1346 0.0123365
R18850 VSS.n1372 VSS.n1346 0.0123365
R18851 VSS.n1372 VSS.n1371 0.0123365
R18852 VSS.n1371 VSS.n1370 0.0123365
R18853 VSS.n1369 VSS.n1368 0.0123365
R18854 VSS.n1368 VSS.n1348 0.0123365
R18855 VSS.n1366 VSS.n1365 0.0123365
R18856 VSS.n1365 VSS.n1364 0.0123365
R18857 VSS.n1362 VSS.n1351 0.0123365
R18858 VSS.n1360 VSS.n1351 0.0123365
R18859 VSS.n1360 VSS.n1359 0.0123365
R18860 VSS.n1355 VSS.n1354 0.0123365
R18861 VSS.n1354 VSS.n805 0.0123365
R18862 VSS.n9627 VSS.n803 0.0123365
R18863 VSS.n9628 VSS.n803 0.0123365
R18864 VSS.n9629 VSS.n802 0.0123365
R18865 VSS.n9631 VSS.n802 0.0123365
R18866 VSS.n9631 VSS.n801 0.0123365
R18867 VSS.n9633 VSS.n801 0.0123365
R18868 VSS.n9635 VSS.n9634 0.0123365
R18869 VSS.n9635 VSS.n798 0.0123365
R18870 VSS.n9763 VSS.n800 0.0123365
R18871 VSS.n9761 VSS.n800 0.0123365
R18872 VSS.n9759 VSS.n9636 0.0123365
R18873 VSS.n9757 VSS.n9636 0.0123365
R18874 VSS.n9757 VSS.n9756 0.0123365
R18875 VSS.n9756 VSS.n9755 0.0123365
R18876 VSS.n9754 VSS.n9638 0.0123365
R18877 VSS.n9753 VSS.n9638 0.0123365
R18878 VSS.n9751 VSS.n9662 0.0123365
R18879 VSS.n9750 VSS.n9662 0.0123365
R18880 VSS.n9749 VSS.n9663 0.0123365
R18881 VSS.n9747 VSS.n9663 0.0123365
R18882 VSS.n9747 VSS.n9746 0.0123365
R18883 VSS.n9746 VSS.n9745 0.0123365
R18884 VSS.n9744 VSS.n9743 0.0123365
R18885 VSS.n9743 VSS.n9665 0.0123365
R18886 VSS.n9741 VSS.n9740 0.0123365
R18887 VSS.n9740 VSS.n9739 0.0123365
R18888 VSS.n9737 VSS.n9668 0.0123365
R18889 VSS.n9735 VSS.n9668 0.0123365
R18890 VSS.n9735 VSS.n9734 0.0123365
R18891 VSS.n9734 VSS.n9733 0.0123365
R18892 VSS.n9732 VSS.n9670 0.0123365
R18893 VSS.n9731 VSS.n9670 0.0123365
R18894 VSS.n9729 VSS.n9718 0.0123365
R18895 VSS.n9728 VSS.n9718 0.0123365
R18896 VSS.n9727 VSS.n9719 0.0123365
R18897 VSS.n9725 VSS.n9719 0.0123365
R18898 VSS.n9725 VSS.n9724 0.0123365
R18899 VSS.n9724 VSS.n9723 0.0123365
R18900 VSS.n9722 VSS.n9721 0.0123365
R18901 VSS.n9721 VSS.n569 0.0123365
R18902 VSS.n10029 VSS.n571 0.0123365
R18903 VSS.n10027 VSS.n571 0.0123365
R18904 VSS.n10022 VSS.n574 0.0123365
R18905 VSS.n10022 VSS.n10021 0.0123365
R18906 VSS.n10017 VSS.n577 0.0123365
R18907 VSS.n10016 VSS.n577 0.0123365
R18908 VSS.n10014 VSS.n9935 0.0123365
R18909 VSS.n10013 VSS.n9935 0.0123365
R18910 VSS.n10012 VSS.n9936 0.0123365
R18911 VSS.n10010 VSS.n9936 0.0123365
R18912 VSS.n10010 VSS.n10009 0.0123365
R18913 VSS.n10009 VSS.n10008 0.0123365
R18914 VSS.n10007 VSS.n10006 0.0123365
R18915 VSS.n10006 VSS.n9938 0.0123365
R18916 VSS.n10004 VSS.n10003 0.0123365
R18917 VSS.n10003 VSS.n10002 0.0123365
R18918 VSS.n10000 VSS.n9940 0.0123365
R18919 VSS.n9998 VSS.n9940 0.0123365
R18920 VSS.n9998 VSS.n9997 0.0123365
R18921 VSS.n9997 VSS.n9996 0.0123365
R18922 VSS.n9995 VSS.n9942 0.0123365
R18923 VSS.n9994 VSS.n9942 0.0123365
R18924 VSS.n9992 VSS.n9967 0.0123365
R18925 VSS.n9991 VSS.n9967 0.0123365
R18926 VSS.n9990 VSS.n9968 0.0123365
R18927 VSS.n9988 VSS.n9968 0.0123365
R18928 VSS.n9988 VSS.n9987 0.0123365
R18929 VSS.n9987 VSS.n9986 0.0123365
R18930 VSS.n9985 VSS.n9984 0.0123365
R18931 VSS.n9984 VSS.n9970 0.0123365
R18932 VSS.n9982 VSS.n9981 0.0123365
R18933 VSS.n9981 VSS.n9980 0.0123365
R18934 VSS.n9978 VSS.n9972 0.0123365
R18935 VSS.n9976 VSS.n9972 0.0123365
R18936 VSS.n9976 VSS.n9975 0.0123365
R18937 VSS.n9975 VSS.n9974 0.0123365
R18938 VSS.n10284 VSS.n253 0.0123169
R18939 VSS.n11460 VSS.n11459 0.0121335
R18940 VSS.n9068 VSS.n9067 0.0120995
R18941 VSS.n9089 VSS.n9088 0.0120995
R18942 VSS.n9016 VSS.n9015 0.0120995
R18943 VSS.n1290 VSS.n1289 0.0120995
R18944 VSS.n10152 VSS.n10151 0.0120995
R18945 VSS.n10159 VSS.n391 0.0120995
R18946 VSS.n371 VSS.n370 0.0120995
R18947 VSS.n10212 VSS.n10211 0.0120995
R18948 VSS.n10219 VSS.n319 0.0120995
R18949 VSS.n308 VSS.n307 0.0120995
R18950 VSS.n10272 VSS.n10271 0.0120995
R18951 VSS.n9383 VSS.n9382 0.0120995
R18952 VSS.n9344 VSS.n9343 0.0120995
R18953 VSS.n9310 VSS.n9309 0.0120995
R18954 VSS.n9246 VSS.n9245 0.0120995
R18955 VSS.n9183 VSS.n9182 0.0120995
R18956 VSS.n1349 VSS.n1348 0.0119138
R18957 VSS.n9764 VSS.n798 0.0119138
R18958 VSS.n9666 VSS.n9665 0.0119138
R18959 VSS.n10030 VSS.n569 0.0119138
R18960 VSS.n9938 VSS.n147 0.0119138
R18961 VSS.n9970 VSS.n138 0.0119138
R18962 VSS.n10727 VSS.n10726 0.0118938
R18963 VSS.n10725 VSS.n10724 0.0118938
R18964 VSS.n10723 VSS.n10722 0.0118938
R18965 VSS.n10718 VSS.n10717 0.0118938
R18966 VSS.n10772 VSS.n10771 0.0118287
R18967 VSS.n10774 VSS.n10773 0.011514
R18968 VSS.n9626 VSS.n805 0.0114911
R18969 VSS.n9627 VSS.n9626 0.0114911
R18970 VSS.n9753 VSS.n9752 0.0114911
R18971 VSS.n9752 VSS.n9751 0.0114911
R18972 VSS.n9731 VSS.n9730 0.0114911
R18973 VSS.n9730 VSS.n9729 0.0114911
R18974 VSS.n10016 VSS.n10015 0.0114911
R18975 VSS.n10015 VSS.n10014 0.0114911
R18976 VSS.n9994 VSS.n9993 0.0114911
R18977 VSS.n9993 VSS.n9992 0.0114911
R18978 VSS.n10638 VSS.n10352 0.0113855
R18979 VSS.n10610 VSS.n10440 0.0113305
R18980 VSS.n11336 VSS.n11335 0.0112405
R18981 VSS.n1356 VSS.n1355 0.0111529
R18982 VSS.n10018 VSS.n10017 0.0111529
R18983 VSS.n11434 VSS.n11433 0.0111311
R18984 VSS.n10745 VSS.n10744 0.0105699
R18985 VSS.n10755 VSS.n10754 0.0105401
R18986 VSS.n10026 VSS.n10025 0.0105188
R18987 VSS.n10728 VSS.n10727 0.0104148
R18988 VSS.n10716 VSS.n10715 0.0103268
R18989 VSS.n10714 VSS.n125 0.0103268
R18990 VSS.n9110 VSS.n1536 0.0102495
R18991 VSS.n851 VSS.n850 0.0102495
R18992 VSS.n10121 VSS.n430 0.0102495
R18993 VSS.n10181 VSS.n360 0.0102495
R18994 VSS.n10241 VSS.n288 0.0102495
R18995 VSS.n11072 VSS.n11069 0.0102495
R18996 VSS.n11218 VSS.n11216 0.0102495
R18997 VSS.n1186 VSS.n1173 0.0102495
R18998 VSS.n9401 VSS.n9400 0.0102495
R18999 VSS.n9232 VSS.n9230 0.0102495
R19000 VSS.n10574 VSS.n10573 0.0101279
R19001 VSS.n10857 VSS.n10856 0.00999301
R19002 VSS.n8989 VSS.n8988 0.00999158
R19003 VSS.n1152 VSS.n1151 0.00999158
R19004 VSS.n10131 VSS.n10128 0.00999158
R19005 VSS.n10191 VSS.n10188 0.00999158
R19006 VSS.n10251 VSS.n10248 0.00999158
R19007 VSS.n11015 VSS.n11012 0.00999158
R19008 VSS.n10961 VSS.n10960 0.00999158
R19009 VSS.n9558 VSS.n1158 0.00999158
R19010 VSS.n9367 VSS.n9365 0.00999158
R19011 VSS.n9156 VSS.n9155 0.00999158
R19012 VSS.n1359 VSS.n1358 0.00992696
R19013 VSS.n10021 VSS.n10020 0.00992696
R19014 VSS.n9082 VSS.n9080 0.00990014
R19015 VSS.n9079 VSS.n9077 0.00990014
R19016 VSS.n9076 VSS.n1536 0.00990014
R19017 VSS.n9109 VSS.n9107 0.00990014
R19018 VSS.n9106 VSS.n9105 0.00990014
R19019 VSS.n9103 VSS.n9102 0.00990014
R19020 VSS.n860 VSS.n858 0.00990014
R19021 VSS.n857 VSS.n855 0.00990014
R19022 VSS.n854 VSS.n853 0.00990014
R19023 VSS.n850 VSS.n848 0.00990014
R19024 VSS.n847 VSS.n536 0.00990014
R19025 VSS.n1106 VSS.n1104 0.00990014
R19026 VSS.n1103 VSS.n1101 0.00990014
R19027 VSS.n1100 VSS.n427 0.00990014
R19028 VSS.n1274 VSS.n430 0.00990014
R19029 VSS.n1278 VSS.n1275 0.00990014
R19030 VSS.n1282 VSS.n1279 0.00990014
R19031 VSS.n926 VSS.n924 0.00990014
R19032 VSS.n923 VSS.n921 0.00990014
R19033 VSS.n920 VSS.n357 0.00990014
R19034 VSS.n376 VSS.n360 0.00990014
R19035 VSS.n380 VSS.n377 0.00990014
R19036 VSS.n384 VSS.n381 0.00990014
R19037 VSS.n999 VSS.n997 0.00990014
R19038 VSS.n996 VSS.n994 0.00990014
R19039 VSS.n993 VSS.n285 0.00990014
R19040 VSS.n292 VSS.n288 0.00990014
R19041 VSS.n296 VSS.n293 0.00990014
R19042 VSS.n300 VSS.n297 0.00990014
R19043 VSS.n11060 VSS.n100 0.00990014
R19044 VSS.n11064 VSS.n11063 0.00990014
R19045 VSS.n11068 VSS.n11065 0.00990014
R19046 VSS.n11073 VSS.n11072 0.00990014
R19047 VSS.n11077 VSS.n11074 0.00990014
R19048 VSS.n11222 VSS.n11220 0.00990014
R19049 VSS.n11219 VSS.n11218 0.00990014
R19050 VSS.n11215 VSS.n11213 0.00990014
R19051 VSS.n11212 VSS.n11211 0.00990014
R19052 VSS.n11209 VSS.n88 0.00990014
R19053 VSS.n1169 VSS.n768 0.00990014
R19054 VSS.n1173 VSS.n1170 0.00990014
R19055 VSS.n1190 VSS.n1189 0.00990014
R19056 VSS.n1194 VSS.n1191 0.00990014
R19057 VSS.n1198 VSS.n1195 0.00990014
R19058 VSS.n9392 VSS.n9391 0.00990014
R19059 VSS.n9396 VSS.n9395 0.00990014
R19060 VSS.n9400 VSS.n9397 0.00990014
R19061 VSS.n9405 VSS.n9404 0.00990014
R19062 VSS.n9409 VSS.n9406 0.00990014
R19063 VSS.n9413 VSS.n9410 0.00990014
R19064 VSS.n9239 VSS.n9237 0.00990014
R19065 VSS.n9236 VSS.n9234 0.00990014
R19066 VSS.n9233 VSS.n9232 0.00990014
R19067 VSS.n9229 VSS.n9227 0.00990014
R19068 VSS.n9226 VSS.n9225 0.00990014
R19069 VSS.n9223 VSS.n1511 0.00990014
R19070 VSS.n11458 VSS.n11457 0.00976426
R19071 VSS.n11456 VSS.n11455 0.00976426
R19072 VSS.n11454 VSS.n11453 0.00976426
R19073 VSS.n11442 VSS.n11441 0.00976426
R19074 VSS.n11440 VSS.n11439 0.00976426
R19075 VSS.n11438 VSS.n11437 0.00976426
R19076 VSS.n11425 VSS.n11424 0.00976426
R19077 VSS.n11423 VSS.n11422 0.00976426
R19078 VSS.n11421 VSS.n11420 0.00976426
R19079 VSS.n11409 VSS.n11408 0.00976426
R19080 VSS.n11407 VSS.n11406 0.00976426
R19081 VSS.n11405 VSS.n11404 0.00976426
R19082 VSS.n574 VSS.n573 0.00975787
R19083 VSS.n891 VSS.n890 0.00969162
R19084 VSS.n10174 VSS.n10173 0.00969162
R19085 VSS.n10234 VSS.n10233 0.00969162
R19086 VSS.n10902 VSS.n10901 0.00969162
R19087 VSS.n720 VSS.n718 0.00969162
R19088 VSS.n1433 VSS.n1232 0.00969162
R19089 VSS.n9278 VSS.n9277 0.00969162
R19090 VSS.n9118 VSS.n1530 0.00969162
R19091 VSS.n8980 VSS.n1559 0.00965149
R19092 VSS.n8984 VSS.n8983 0.00965149
R19093 VSS.n8988 VSS.n8985 0.00965149
R19094 VSS.n8993 VSS.n8992 0.00965149
R19095 VSS.n8997 VSS.n8994 0.00965149
R19096 VSS.n9001 VSS.n8998 0.00965149
R19097 VSS.n1135 VSS.n1134 0.00965149
R19098 VSS.n1139 VSS.n1138 0.00965149
R19099 VSS.n1143 VSS.n1140 0.00965149
R19100 VSS.n1151 VSS.n1149 0.00965149
R19101 VSS.n1148 VSS.n1147 0.00965149
R19102 VSS.n913 VSS.n911 0.00965149
R19103 VSS.n910 VSS.n908 0.00965149
R19104 VSS.n907 VSS.n419 0.00965149
R19105 VSS.n10132 VSS.n10131 0.00965149
R19106 VSS.n10136 VSS.n10133 0.00965149
R19107 VSS.n10140 VSS.n10137 0.00965149
R19108 VSS.n1032 VSS.n1030 0.00965149
R19109 VSS.n1029 VSS.n1027 0.00965149
R19110 VSS.n1026 VSS.n347 0.00965149
R19111 VSS.n10192 VSS.n10191 0.00965149
R19112 VSS.n10196 VSS.n10193 0.00965149
R19113 VSS.n10200 VSS.n10197 0.00965149
R19114 VSS.n952 VSS.n950 0.00965149
R19115 VSS.n949 VSS.n947 0.00965149
R19116 VSS.n946 VSS.n275 0.00965149
R19117 VSS.n10252 VSS.n10251 0.00965149
R19118 VSS.n10256 VSS.n10253 0.00965149
R19119 VSS.n10260 VSS.n10257 0.00965149
R19120 VSS.n11003 VSS.n11002 0.00965149
R19121 VSS.n11007 VSS.n11006 0.00965149
R19122 VSS.n11011 VSS.n11008 0.00965149
R19123 VSS.n11016 VSS.n11015 0.00965149
R19124 VSS.n11020 VSS.n11017 0.00965149
R19125 VSS.n10956 VSS.n10955 0.00965149
R19126 VSS.n10960 VSS.n10957 0.00965149
R19127 VSS.n10965 VSS.n10964 0.00965149
R19128 VSS.n10969 VSS.n10966 0.00965149
R19129 VSS.n10973 VSS.n10970 0.00965149
R19130 VSS.n1154 VSS.n793 0.00965149
R19131 VSS.n1158 VSS.n1155 0.00965149
R19132 VSS.n9557 VSS.n9555 0.00965149
R19133 VSS.n9554 VSS.n9553 0.00965149
R19134 VSS.n9551 VSS.n9550 0.00965149
R19135 VSS.n9374 VSS.n9372 0.00965149
R19136 VSS.n9371 VSS.n9369 0.00965149
R19137 VSS.n9368 VSS.n9367 0.00965149
R19138 VSS.n9364 VSS.n9362 0.00965149
R19139 VSS.n9361 VSS.n9360 0.00965149
R19140 VSS.n9358 VSS.n9357 0.00965149
R19141 VSS.n9147 VSS.n1521 0.00965149
R19142 VSS.n9151 VSS.n9150 0.00965149
R19143 VSS.n9155 VSS.n9152 0.00965149
R19144 VSS.n9160 VSS.n9159 0.00965149
R19145 VSS.n9164 VSS.n9161 0.00965149
R19146 VSS.n9168 VSS.n9165 0.00965149
R19147 VSS.n11431 VSS.n11428 0.00958201
R19148 VSS.n11459 VSS.n14 0.00949089
R19149 VSS.n11458 VSS.n14 0.00949089
R19150 VSS.n11457 VSS.n15 0.00949089
R19151 VSS.n11456 VSS.n15 0.00949089
R19152 VSS.n11455 VSS.n16 0.00949089
R19153 VSS.n11454 VSS.n16 0.00949089
R19154 VSS.n11453 VSS.n17 0.00949089
R19155 VSS.n11452 VSS.n17 0.00949089
R19156 VSS.n11294 VSS.n23 0.00949089
R19157 VSS.n11443 VSS.n24 0.00949089
R19158 VSS.n11442 VSS.n24 0.00949089
R19159 VSS.n11441 VSS.n25 0.00949089
R19160 VSS.n11440 VSS.n25 0.00949089
R19161 VSS.n11439 VSS.n26 0.00949089
R19162 VSS.n11438 VSS.n26 0.00949089
R19163 VSS.n11437 VSS.n27 0.00949089
R19164 VSS.n11436 VSS.n27 0.00949089
R19165 VSS.n11435 VSS.n28 0.00949089
R19166 VSS.n11434 VSS.n28 0.00949089
R19167 VSS.n11428 VSS.n38 0.00949089
R19168 VSS.n11427 VSS.n38 0.00949089
R19169 VSS.n11426 VSS.n39 0.00949089
R19170 VSS.n11425 VSS.n39 0.00949089
R19171 VSS.n11424 VSS.n40 0.00949089
R19172 VSS.n11423 VSS.n40 0.00949089
R19173 VSS.n11422 VSS.n41 0.00949089
R19174 VSS.n11421 VSS.n41 0.00949089
R19175 VSS.n11420 VSS.n42 0.00949089
R19176 VSS.n11419 VSS.n42 0.00949089
R19177 VSS.n133 VSS.n48 0.00949089
R19178 VSS.n11410 VSS.n49 0.00949089
R19179 VSS.n11409 VSS.n49 0.00949089
R19180 VSS.n11408 VSS.n50 0.00949089
R19181 VSS.n11407 VSS.n50 0.00949089
R19182 VSS.n11406 VSS.n51 0.00949089
R19183 VSS.n11405 VSS.n51 0.00949089
R19184 VSS.n11404 VSS.n52 0.00949089
R19185 VSS.n11403 VSS.n52 0.00949089
R19186 VSS.n11402 VSS.n53 0.00949089
R19187 VSS.n11401 VSS.n53 0.00949089
R19188 VSS.n63 VSS.n3 0.00949089
R19189 VSS.n11310 VSS.n125 0.00947638
R19190 VSS.n900 VSS.n898 0.00936227
R19191 VSS.n897 VSS.n895 0.00936227
R19192 VSS.n894 VSS.n893 0.00936227
R19193 VSS.n890 VSS.n888 0.00936227
R19194 VSS.n887 VSS.n886 0.00936227
R19195 VSS.n1069 VSS.n1067 0.00936227
R19196 VSS.n1066 VSS.n1064 0.00936227
R19197 VSS.n1063 VSS.n397 0.00936227
R19198 VSS.n10173 VSS.n10171 0.00936227
R19199 VSS.n10170 VSS.n10169 0.00936227
R19200 VSS.n10167 VSS.n10166 0.00936227
R19201 VSS.n939 VSS.n937 0.00936227
R19202 VSS.n936 VSS.n934 0.00936227
R19203 VSS.n933 VSS.n325 0.00936227
R19204 VSS.n10233 VSS.n10231 0.00936227
R19205 VSS.n10230 VSS.n10229 0.00936227
R19206 VSS.n10227 VSS.n10226 0.00936227
R19207 VSS.n10908 VSS.n10906 0.00936227
R19208 VSS.n10905 VSS.n10904 0.00936227
R19209 VSS.n10901 VSS.n10899 0.00936227
R19210 VSS.n10898 VSS.n10897 0.00936227
R19211 VSS.n724 VSS.n722 0.00936227
R19212 VSS.n721 VSS.n720 0.00936227
R19213 VSS.n717 VSS.n715 0.00936227
R19214 VSS.n714 VSS.n713 0.00936227
R19215 VSS.n711 VSS.n212 0.00936227
R19216 VSS.n1437 VSS.n1435 0.00936227
R19217 VSS.n1434 VSS.n1433 0.00936227
R19218 VSS.n1231 VSS.n1229 0.00936227
R19219 VSS.n1228 VSS.n1227 0.00936227
R19220 VSS.n1225 VSS.n1219 0.00936227
R19221 VSS.n9269 VSS.n1503 0.00936227
R19222 VSS.n9273 VSS.n9272 0.00936227
R19223 VSS.n9277 VSS.n9274 0.00936227
R19224 VSS.n9282 VSS.n9281 0.00936227
R19225 VSS.n9286 VSS.n9283 0.00936227
R19226 VSS.n9290 VSS.n9287 0.00936227
R19227 VSS.n9056 VSS.n9054 0.00936227
R19228 VSS.n9053 VSS.n9051 0.00936227
R19229 VSS.n9050 VSS.n1530 0.00936227
R19230 VSS.n9122 VSS.n9121 0.00936227
R19231 VSS.n9126 VSS.n9123 0.00936227
R19232 VSS.n9130 VSS.n9127 0.00936227
R19233 VSS.n10840 VSS.n10734 0.0092701
R19234 VSS.n11295 VSS.n18 0.00924789
R19235 VSS.n134 VSS.n43 0.00924789
R19236 VSS.n9885 VSS.n9884 0.00862937
R19237 VSS.n9872 VSS.n673 0.00862937
R19238 VSS.n9519 VSS.n9518 0.00862937
R19239 VSS.n9895 VSS.n9894 0.00862937
R19240 VSS.n9926 VSS.n583 0.00862937
R19241 VSS.n11282 VSS.n22 0.00862937
R19242 VSS.n141 VSS.n47 0.00862937
R19243 VSS.n9617 VSS.n810 0.00862937
R19244 VSS.n778 VSS.n648 0.00852448
R19245 VSS.n9879 VSS.n667 0.00852448
R19246 VSS.n1255 VSS.n1247 0.00852448
R19247 VSS.n9654 VSS.n628 0.00852448
R19248 VSS.n9918 VSS.n597 0.00852448
R19249 VSS.n11043 VSS.n19 0.00852448
R19250 VSS.n9959 VSS.n44 0.00852448
R19251 VSS.n9610 VSS.n9609 0.00852448
R19252 VSS.n9496 VSS.n9493 0.00847863
R19253 VSS.n9886 VSS.n648 0.00847203
R19254 VSS.n9881 VSS.n654 0.00847203
R19255 VSS.n1178 VSS.n679 0.00847203
R19256 VSS.n9879 VSS.n668 0.00847203
R19257 VSS.n9520 VSS.n1255 0.00847203
R19258 VSS.n9893 VSS.n628 0.00847203
R19259 VSS.n9907 VSS.n9906 0.00847203
R19260 VSS.n9904 VSS.n9903 0.00847203
R19261 VSS.n9918 VSS.n9917 0.00847203
R19262 VSS.n11281 VSS.n19 0.00847203
R19263 VSS.n140 VSS.n44 0.00847203
R19264 VSS.n9610 VSS.n815 0.00847203
R19265 VSS.n9884 VSS.n649 0.00836713
R19266 VSS.n9882 VSS.n653 0.00836713
R19267 VSS.n9854 VSS.n9853 0.00836713
R19268 VSS.n9872 VSS.n9871 0.00836713
R19269 VSS.n9518 VSS.n1267 0.00836713
R19270 VSS.n9895 VSS.n641 0.00836713
R19271 VSS.n621 VSS.n620 0.00836713
R19272 VSS.n9698 VSS.n627 0.00836713
R19273 VSS.n9927 VSS.n9926 0.00836713
R19274 VSS.n9947 VSS.n22 0.00836713
R19275 VSS.n11187 VSS.n47 0.00836713
R19276 VSS.n9618 VSS.n9617 0.00836713
R19277 VSS.n9500 VSS.n9499 0.00819275
R19278 VSS.n9492 VSS.n1375 0.00819275
R19279 VSS.n10552 VSS.n10551 0.00799437
R19280 VSS.n10540 VSS.n10539 0.00799437
R19281 VSS.n9469 VSS.n9468 0.00788202
R19282 VSS.n9462 VSS.n9458 0.00780812
R19283 VSS.n9441 VSS.n9440 0.00779878
R19284 VSS.n10839 VSS.n10735 0.00773913
R19285 VSS.n10836 VSS.n10790 0.00773913
R19286 VSS.n10835 VSS.n10790 0.00773913
R19287 VSS.n10829 VSS.n10811 0.00773913
R19288 VSS.n10826 VSS.n10820 0.00773913
R19289 VSS.n9506 VSS.n9505 0.00767297
R19290 VSS.n1339 VSS.n1338 0.00767297
R19291 VSS.n10811 VSS.n10810 0.00761685
R19292 VSS.n10590 VSS.n10589 0.00752176
R19293 VSS.n10490 VSS.n10489 0.00752176
R19294 VSS.n10538 VSS.n10491 0.00752176
R19295 VSS.n10525 VSS.n10524 0.007488
R19296 VSS.n10513 VSS.n10512 0.007488
R19297 VSS.n10741 VSS.n247 0.00721329
R19298 VSS.n10636 VSS.n10635 0.00704376
R19299 VSS.n10760 VSS.n241 0.00704376
R19300 VSS.n10761 VSS.n10760 0.00704376
R19301 VSS.n11384 VSS.n11382 0.00703487
R19302 VSS.n10505 VSS.n10504 0.00701538
R19303 VSS.n10522 VSS.n10506 0.00701538
R19304 VSS.n10521 VSS.n10507 0.00701538
R19305 VSS.n10509 VSS.n10508 0.00701538
R19306 VSS.n10518 VSS.n10517 0.00701538
R19307 VSS.n10516 VSS.n10515 0.00701538
R19308 VSS.n9447 VSS.n9446 0.00681098
R19309 VSS.n10567 VSS.n10556 0.00674846
R19310 VSS.n10570 VSS.n10567 0.00674846
R19311 VSS.n9503 VSS.n9502 0.00671138
R19312 VSS.n1342 VSS.n1341 0.00671138
R19313 VSS.n10484 VSS.n10483 0.00667779
R19314 VSS.n10549 VSS.n10485 0.00667779
R19315 VSS.n10548 VSS.n10486 0.00667779
R19316 VSS.n10488 VSS.n10487 0.00667779
R19317 VSS.n10545 VSS.n10544 0.00667779
R19318 VSS.n10543 VSS.n10542 0.00667779
R19319 VSS.n9434 VSS.n9428 0.00659146
R19320 VSS.n10720 VSS.n10719 0.00658034
R19321 VSS.n10773 VSS.n10772 0.00653147
R19322 VSS.n9504 VSS.n1340 0.00647748
R19323 VSS.n9501 VSS.n1343 0.00639951
R19324 VSS.n10775 VSS.n10774 0.00632168
R19325 VSS.n10732 VSS.n10701 0.00625167
R19326 VSS.n10610 VSS.n10609 0.00619059
R19327 VSS.n10592 VSS.n10482 0.00617142
R19328 VSS.n10527 VSS.n10500 0.00617142
R19329 VSS.n10503 VSS.n10502 0.00617142
R19330 VSS.n10511 VSS.n10510 0.00617142
R19331 VSS.n10348 VSS.n10347 0.00617142
R19332 VSS.n9488 VSS.n9487 0.00616561
R19333 VSS.n10856 VSS.n10855 0.00611189
R19334 VSS.n9490 VSS.n9489 0.00582775
R19335 VSS.n9474 VSS.n1377 0.00582775
R19336 VSS.n10721 VSS.n10720 0.00581345
R19337 VSS.n10825 VSS.n10824 0.00559341
R19338 VSS.n81 VSS.n78 0.00554673
R19339 VSS.n10894 VSS.n10893 0.00554202
R19340 VSS.n11463 VSS.n11462 0.00554202
R19341 VSS.n11462 VSS.n11461 0.00554202
R19342 VSS.n11310 VSS.n127 0.00550787
R19343 VSS.n11102 VSS.n11101 0.005488
R19344 VSS.n11084 VSS.n11080 0.005488
R19345 VSS.n10910 VSS.n10909 0.00547006
R19346 VSS.n11082 VSS.n11081 0.00536194
R19347 VSS.n8954 VSS.n1579 0.00535451
R19348 VSS.n10827 VSS.n10812 0.00529348
R19349 VSS.n10873 VSS.n10872 0.00528992
R19350 VSS.n192 VSS.n191 0.00523684
R19351 VSS.n197 VSS.n196 0.00523684
R19352 VSS.n470 VSS.n469 0.00523684
R19353 VSS.n475 VSS.n474 0.00523684
R19354 VSS.n263 VSS.n262 0.00523684
R19355 VSS.n268 VSS.n267 0.00523684
R19356 VSS.n335 VSS.n334 0.00523684
R19357 VSS.n340 VSS.n339 0.00523684
R19358 VSS.n407 VSS.n406 0.00523684
R19359 VSS.n412 VSS.n411 0.00523684
R19360 VSS.n11099 VSS.n11086 0.00523589
R19361 VSS.n11444 VSS.n23 0.00520807
R19362 VSS.n11411 VSS.n48 0.00520807
R19363 VSS.n1337 VSS.n1336 0.00520401
R19364 VSS.n10060 VSS.n10059 0.00516387
R19365 VSS.n11083 VSS.n11078 0.00516387
R19366 VSS.n11452 VSS.n11451 0.00514732
R19367 VSS.n11419 VSS.n11418 0.00514732
R19368 VSS.n10108 VSS.n10107 0.00512785
R19369 VSS.n450 VSS.n449 0.00512785
R19370 VSS.n10105 VSS.n451 0.00512785
R19371 VSS.n11451 VSS.n18 0.00511694
R19372 VSS.n11418 VSS.n43 0.00511694
R19373 VSS.n538 VSS.n537 0.00507383
R19374 VSS.n10057 VSS.n539 0.00507383
R19375 VSS.n10056 VSS.n540 0.00507383
R19376 VSS.n542 VSS.n541 0.00507383
R19377 VSS.n11444 VSS.n11443 0.00505619
R19378 VSS.n11411 VSS.n11410 0.00505619
R19379 VSS.n1316 VSS.n1315 0.00496579
R19380 VSS.n1297 VSS.n1273 0.00496579
R19381 VSS.n10891 VSS.n10874 0.00492977
R19382 VSS.n10890 VSS.n10889 0.00492977
R19383 VSS.n10888 VSS.n10875 0.00492977
R19384 VSS.n10855 VSS.n10854 0.00490559
R19385 VSS.n10637 VSS.n240 0.00489366
R19386 VSS.n10863 VSS.n241 0.00489366
R19387 VSS.n1296 VSS.n1295 0.00487585
R19388 VSS.n9495 VSS.n9494 0.00486616
R19389 VSS.n9497 VSS.n1345 0.00486616
R19390 VSS.n10834 VSS.n10833 0.00485326
R19391 VSS.n551 VSS.n549 0.00483974
R19392 VSS.n10045 VSS.n10044 0.00483974
R19393 VSS.n11105 VSS.n11104 0.00483974
R19394 VSS.n10100 VSS.n457 0.00482173
R19395 VSS.n10099 VSS.n10098 0.00482173
R19396 VSS.n10097 VSS.n10096 0.00482173
R19397 VSS.n10054 VSS.n10053 0.0047497
R19398 VSS.n186 VSS.n185 0.00469568
R19399 VSS.n11147 VSS.n187 0.00469568
R19400 VSS.n11146 VSS.n11145 0.00469568
R19401 VSS.n10530 VSS.n10498 0.00465229
R19402 VSS.n531 VSS.n530 0.00464166
R19403 VSS.n529 VSS.n528 0.00464166
R19404 VSS.n515 VSS.n514 0.00464166
R19405 VSS.n10061 VSS.n533 0.00464166
R19406 VSS.n10809 VSS.n10808 0.00463315
R19407 VSS.n9491 VSS.n1376 0.00463225
R19408 VSS.n10877 VSS.n10876 0.00460564
R19409 VSS.n10886 VSS.n10885 0.00460564
R19410 VSS.n11336 VSS.n105 0.00455578
R19411 VSS.n11338 VSS.n105 0.00455578
R19412 VSS.n11098 VSS.n11087 0.00455162
R19413 VSS.n11089 VSS.n11088 0.00455162
R19414 VSS.n11096 VSS.n11095 0.00455162
R19415 VSS.n11091 VSS.n11090 0.00455162
R19416 VSS.n11093 VSS.n11092 0.00455162
R19417 VSS.n456 VSS.n455 0.00446158
R19418 VSS.n10064 VSS.n513 0.00446158
R19419 VSS.n10838 VSS.n10789 0.0044375
R19420 VSS.n10638 VSS.n10637 0.00442625
R19421 VSS.n10104 VSS.n452 0.00442557
R19422 VSS.n454 VSS.n453 0.00442557
R19423 VSS.n747 VSS.n726 0.0044234
R19424 VSS.n747 VSS.n746 0.0044234
R19425 VSS.n10838 VSS.n10837 0.00441304
R19426 VSS.n10048 VSS.n10047 0.00440756
R19427 VSS.n11246 VSS.n11245 0.00438136
R19428 VSS.n11229 VSS.n11225 0.00438136
R19429 VSS.n11243 VSS.n11230 0.00438136
R19430 VSS.n10895 VSS.n235 0.00437155
R19431 VSS.n119 VSS.n13 0.00436387
R19432 VSS.n1309 VSS.n1308 0.00433553
R19433 VSS.n1307 VSS.n1306 0.00433553
R19434 VSS.n10854 VSS.n10853 0.00432867
R19435 VSS.n11227 VSS.n11226 0.00428328
R19436 VSS.n10502 VSS.n10500 0.00428095
R19437 VSS.n10525 VSS.n10503 0.00428095
R19438 VSS.n10512 VSS.n10511 0.00428095
R19439 VSS.n10510 VSS.n10346 0.00428095
R19440 VSS.n10655 VSS.n10346 0.00428095
R19441 VSS.n10654 VSS.n10347 0.00428095
R19442 VSS.n1313 VSS.n1311 0.00426351
R19443 VSS.n10535 VSS.n10534 0.00424719
R19444 VSS.n10528 VSS.n10527 0.00424719
R19445 VSS.n10792 VSS.n10791 0.00424185
R19446 VSS.n11055 VSS.n11054 0.00422749
R19447 VSS.n11108 VSS.n11056 0.00422749
R19448 VSS.n11107 VSS.n11057 0.00422749
R19449 VSS.n11059 VSS.n11058 0.00422749
R19450 VSS.n461 VSS.n459 0.00419148
R19451 VSS.n10093 VSS.n10092 0.00419148
R19452 VSS.n478 VSS.n460 0.00419148
R19453 VSS.n553 VSS.n550 0.00413745
R19454 VSS.n10042 VSS.n554 0.00413745
R19455 VSS.n9826 VSS.n9823 0.00412915
R19456 VSS.n11228 VSS.n11223 0.00412915
R19457 VSS.n10103 VSS.n10102 0.00410144
R19458 VSS.n1450 VSS.n1449 0.00410112
R19459 VSS.n1440 VSS.n1439 0.00410112
R19460 VSS.n1447 VSS.n1441 0.00410112
R19461 VSS.n1376 VSS.n1375 0.0040605
R19462 VSS.n9491 VSS.n9490 0.0040605
R19463 VSS.n9825 VSS.n9824 0.00405908
R19464 VSS.n9828 VSS.n765 0.00405908
R19465 VSS.n9831 VSS.n9830 0.00405908
R19466 VSS.n9829 VSS.n764 0.00405908
R19467 VSS.n9195 VSS.n9194 0.00405263
R19468 VSS.n9190 VSS.n9189 0.00405263
R19469 VSS.n9331 VSS.n9330 0.00405263
R19470 VSS.n9326 VSS.n9325 0.00405263
R19471 VSS.n169 VSS.n168 0.00405263
R19472 VSS.n164 VSS.n163 0.00405263
R19473 VSS.n9577 VSS.n9576 0.00405263
R19474 VSS.n9572 VSS.n9571 0.00405263
R19475 VSS.n9028 VSS.n9027 0.00405263
R19476 VSS.n9023 VSS.n9022 0.00405263
R19477 VSS.n544 VSS.n543 0.00404742
R19478 VSS.n10051 VSS.n545 0.00404742
R19479 VSS.n10050 VSS.n10049 0.00404742
R19480 VSS.n10728 VSS.n10703 0.00401077
R19481 VSS.n10730 VSS.n10703 0.00401077
R19482 VSS.n4805 VSS.n1580 0.00400211
R19483 VSS.n10833 VSS.n10791 0.00399728
R19484 VSS.n9388 VSS.n1475 0.00399694
R19485 VSS.n11120 VSS.n11119 0.0039934
R19486 VSS.n11035 VSS.n11034 0.0039934
R19487 VSS.n1473 VSS.n1418 0.00397501
R19488 VSS.n1472 VSS.n1471 0.00397501
R19489 VSS.n448 VSS.n447 0.00395738
R19490 VSS.n745 VSS.n727 0.00394699
R19491 VSS.n729 VSS.n728 0.00394699
R19492 VSS.n743 VSS.n742 0.00394699
R19493 VSS.n11 VSS.n10 0.00392137
R19494 VSS.n11463 VSS.n12 0.00392137
R19495 VSS.n10884 VSS.n10878 0.00390336
R19496 VSS.n10880 VSS.n10879 0.00390336
R19497 VSS.n10883 VSS.n10882 0.00390336
R19498 VSS.n11111 VSS.n11110 0.00390336
R19499 VSS.n697 VSS.n695 0.00387693
R19500 VSS.n761 VSS.n760 0.00387693
R19501 VSS.n11249 VSS.n11248 0.00387693
R19502 VSS.n9599 VSS.n828 0.00386291
R19503 VSS.n830 VSS.n829 0.00386291
R19504 VSS.n9598 VSS.n9597 0.00386291
R19505 VSS.n10776 VSS.n10769 0.00385664
R19506 VSS.n9494 VSS.n1345 0.0038266
R19507 VSS.n9497 VSS.n9496 0.0038266
R19508 VSS.n10041 VSS.n555 0.00381333
R19509 VSS.n557 VSS.n556 0.00381333
R19510 VSS.n9834 VSS.n9833 0.00380687
R19511 VSS.n10074 VSS.n497 0.00379532
R19512 VSS.n11325 VSS.n11324 0.00377731
R19513 VSS.n10551 VSS.n10483 0.00377457
R19514 VSS.n10485 VSS.n10484 0.00377457
R19515 VSS.n10549 VSS.n10548 0.00377457
R19516 VSS.n10487 VSS.n10486 0.00377457
R19517 VSS.n10545 VSS.n10488 0.00377457
R19518 VSS.n10544 VSS.n10543 0.00377457
R19519 VSS.n10542 VSS.n10540 0.00377457
R19520 VSS.n11157 VSS.n11156 0.00376483
R19521 VSS.n11159 VSS.n158 0.00376483
R19522 VSS.n11158 VSS.n177 0.00376483
R19523 VSS.n1301 VSS.n1300 0.00372329
R19524 VSS.n1304 VSS.n1302 0.00372329
R19525 VSS.n9813 VSS.n9812 0.00372279
R19526 VSS.n9811 VSS.n770 0.00372279
R19527 VSS.n9818 VSS.n9817 0.00372279
R19528 VSS.n9821 VSS.n769 0.00372279
R19529 VSS.n1295 VSS.n1282 0.00370748
R19530 VSS.n385 VSS.n384 0.00370748
R19531 VSS.n313 VSS.n300 0.00370748
R19532 VSS.n517 VSS.n503 0.00370528
R19533 VSS.n519 VSS.n518 0.00370528
R19534 VSS.n524 VSS.n521 0.00370528
R19535 VSS.n523 VSS.n522 0.00370528
R19536 VSS.n526 VSS.n516 0.00370528
R19537 VSS.n740 VSS.n739 0.00369477
R19538 VSS.n731 VSS.n730 0.00369477
R19539 VSS.n11129 VSS.n11128 0.00368728
R19540 VSS.n11025 VSS.n11024 0.00368728
R19541 VSS.n119 VSS.n118 0.00367595
R19542 VSS.n9083 VSS.n9082 0.00367572
R19543 VSS.n9391 VSS.n9388 0.00367572
R19544 VSS.n9240 VSS.n9239 0.00367572
R19545 VSS.n11340 VSS.n103 0.00367038
R19546 VSS.n11138 VSS.n11137 0.00366927
R19547 VSS.n203 VSS.n202 0.00366927
R19548 VSS.n11135 VSS.n204 0.00366927
R19549 VSS.n11134 VSS.n11132 0.00366927
R19550 VSS.n11242 VSS.n11231 0.00365273
R19551 VSS.n11233 VSS.n11232 0.00365273
R19552 VSS.n11240 VSS.n11239 0.00365273
R19553 VSS.n11235 VSS.n11234 0.00365273
R19554 VSS.n11237 VSS.n11236 0.00365273
R19555 VSS.n1318 VSS.n1272 0.00365126
R19556 VSS.n10141 VSS.n10140 0.00362264
R19557 VSS.n10201 VSS.n10200 0.00362264
R19558 VSS.n10261 VSS.n10260 0.00362264
R19559 VSS.n11038 VSS.n11036 0.00359724
R19560 VSS.n11305 VSS.n123 0.00359693
R19561 VSS.n11308 VSS.n123 0.00359693
R19562 VSS.n9039 VSS.n1559 0.00359172
R19563 VSS.n9375 VSS.n9374 0.00359172
R19564 VSS.n9206 VSS.n1521 0.00359172
R19565 VSS.n9601 VSS.n9600 0.00358267
R19566 VSS.n9816 VSS.n9815 0.00358267
R19567 VSS.n11117 VSS.n11051 0.00356122
R19568 VSS.n10828 VSS.n10827 0.00355707
R19569 VSS.n1446 VSS.n1442 0.00355465
R19570 VSS.n1444 VSS.n1443 0.00355465
R19571 VSS.n9841 VSS.n9840 0.00354064
R19572 VSS.n10166 VSS.n10164 0.00352395
R19573 VSS.n10226 VSS.n10224 0.00352395
R19574 VSS.n749 VSS.n725 0.00351261
R19575 VSS.n9315 VSS.n1503 0.00349401
R19576 VSS.n9062 VSS.n9056 0.00349401
R19577 VSS.n1468 VSS.n1467 0.00348459
R19578 VSS.n1466 VSS.n1465 0.00348459
R19579 VSS.n1424 VSS.n1423 0.00348459
R19580 VSS.n496 VSS.n495 0.00347119
R19581 VSS.n10076 VSS.n10075 0.00347119
R19582 VSS.n10524 VSS.n10504 0.00343698
R19583 VSS.n10506 VSS.n10505 0.00343698
R19584 VSS.n10522 VSS.n10521 0.00343698
R19585 VSS.n10508 VSS.n10507 0.00343698
R19586 VSS.n10518 VSS.n10509 0.00343698
R19587 VSS.n10517 VSS.n10516 0.00343698
R19588 VSS.n10515 VSS.n10513 0.00343698
R19589 VSS.n499 VSS.n498 0.00343517
R19590 VSS.n11126 VSS.n11027 0.00343517
R19591 VSS.n1470 VSS.n1419 0.00342854
R19592 VSS.n11199 VSS.n11198 0.00340051
R19593 VSS.n11252 VSS.n11200 0.00340051
R19594 VSS.n11251 VSS.n11201 0.00340051
R19595 VSS.n11203 VSS.n11202 0.00340051
R19596 VSS.n1303 VSS.n441 0.00339916
R19597 VSS.n10114 VSS.n442 0.00339916
R19598 VSS.n444 VSS.n443 0.00339916
R19599 VSS.n10112 VSS.n10111 0.00339916
R19600 VSS.n10084 VSS.n10083 0.00339916
R19601 VSS.n9475 VSS.n9474 0.00338478
R19602 VSS.n11022 VSS.n11021 0.00338115
R19603 VSS.n9589 VSS.n9567 0.00337249
R19604 VSS.n9593 VSS.n9592 0.00337249
R19605 VSS.n9588 VSS.n9587 0.00337249
R19606 VSS.n10039 VSS.n10038 0.00334514
R19607 VSS.n1357 VSS.n1356 0.00333232
R19608 VSS.n10019 VSS.n10018 0.00333232
R19609 VSS.n699 VSS.n696 0.00333045
R19610 VSS.n758 VSS.n700 0.00333045
R19611 VSS.n1445 VSS.n827 0.00330243
R19612 VSS.n9440 VSS.n9439 0.00329878
R19613 VSS.n11122 VSS.n11031 0.00329112
R19614 VSS.n11033 VSS.n11032 0.00329112
R19615 VSS.n9476 VSS.n9475 0.00328083
R19616 VSS.n493 VSS.n492 0.00327311
R19617 VSS.n10081 VSS.n10080 0.00327311
R19618 VSS.n10079 VSS.n10078 0.00327311
R19619 VSS.n495 VSS.n494 0.00327311
R19620 VSS.n9836 VSS.n9835 0.00326039
R19621 VSS.n9838 VSS.n763 0.00326039
R19622 VSS.n9837 VSS.n692 0.00326039
R19623 VSS.n10111 VSS.n10110 0.0032551
R19624 VSS.n447 VSS.n446 0.0032551
R19625 VSS.n10089 VSS.n484 0.0032551
R19626 VSS.n486 VSS.n485 0.0032551
R19627 VSS.n10087 VSS.n10086 0.0032551
R19628 VSS.n489 VSS.n488 0.0032551
R19629 VSS.n10084 VSS.n490 0.0032551
R19630 VSS.n11267 VSS.n11180 0.00321836
R19631 VSS.n11182 VSS.n11181 0.00321836
R19632 VSS.n10831 VSS.n10830 0.00321467
R19633 VSS.n11053 VSS.n11052 0.00320108
R19634 VSS.n11115 VSS.n11114 0.00320108
R19635 VSS.n11113 VSS.n11112 0.00320108
R19636 VSS.n1438 VSS.n1429 0.00319033
R19637 VSS.n10533 VSS.n10532 0.00316692
R19638 VSS.n10025 VSS.n10024 0.00316322
R19639 VSS.n11340 VSS.n11339 0.00315277
R19640 VSS.n737 VSS.n732 0.0031483
R19641 VSS.n736 VSS.n735 0.0031483
R19642 VSS.n734 VSS.n733 0.0031483
R19643 VSS.n11255 VSS.n11254 0.0031483
R19644 VSS.n10832 VSS.n10809 0.0031413
R19645 VSS.n10638 VSS.n10635 0.0031175
R19646 VSS.n10535 VSS.n10492 0.0030994
R19647 VSS.n11433 VSS.n31 0.00308184
R19648 VSS.n10024 VSS.n573 0.00307868
R19649 VSS.n757 VSS.n701 0.00307823
R19650 VSS.n703 VSS.n702 0.00307823
R19651 VSS.n492 VSS.n491 0.00307503
R19652 VSS.n10072 VSS.n10071 0.00307503
R19653 VSS.n501 VSS.n500 0.00307503
R19654 VSS.n10070 VSS.n502 0.00307503
R19655 VSS.n11125 VSS.n11028 0.00307503
R19656 VSS.n11030 VSS.n11029 0.00307503
R19657 VSS.n9495 VSS.n1344 0.00307291
R19658 VSS.n9793 VSS.n9792 0.00306422
R19659 VSS.n11131 VSS.n205 0.00305702
R19660 VSS.n1463 VSS.n1425 0.00300817
R19661 VSS.n4806 VSS.n4805 0.00300278
R19662 VSS.n9803 VSS.n9802 0.00299416
R19663 VSS.n9801 VSS.n772 0.00299416
R19664 VSS.n9808 VSS.n9805 0.00299416
R19665 VSS.n9807 VSS.n9806 0.00299416
R19666 VSS.n9810 VSS.n771 0.00299416
R19667 VSS.n11132 VSS.n11131 0.00298499
R19668 VSS.n11021 VSS.n205 0.00298499
R19669 VSS.n11276 VSS.n152 0.00298015
R19670 VSS.n11173 VSS.n11172 0.00298015
R19671 VSS.n11274 VSS.n11273 0.00298015
R19672 VSS.n10083 VSS.n491 0.00296699
R19673 VSS.n10071 VSS.n500 0.00296699
R19674 VSS.n502 VSS.n501 0.00296699
R19675 VSS.n11126 VSS.n11125 0.00296699
R19676 VSS.n11029 VSS.n11028 0.00296699
R19677 VSS.n11123 VSS.n11030 0.00296699
R19678 VSS.n11163 VSS.n11162 0.00296614
R19679 VSS.n11165 VSS.n11164 0.00296614
R19680 VSS.n11168 VSS.n155 0.00296614
R19681 VSS.n10604 VSS.n10441 0.00296504
R19682 VSS.n1416 VSS.n1403 0.00295213
R19683 VSS.n10587 VSS.n10482 0.00293061
R19684 VSS.n10591 VSS.n10590 0.00293061
R19685 VSS.n10589 VSS.n10552 0.00293061
R19686 VSS.n10539 VSS.n10489 0.00293061
R19687 VSS.n10491 VSS.n10490 0.00293061
R19688 VSS.n11461 VSS.n11460 0.00291297
R19689 VSS.n11265 VSS.n11264 0.00291009
R19690 VSS.n1358 VSS.n1357 0.00290958
R19691 VSS.n10020 VSS.n10019 0.00290958
R19692 VSS.n11261 VSS.n11195 0.00288206
R19693 VSS.n9035 VSS.n9034 0.00288205
R19694 VSS.n10148 VSS.n10147 0.00288205
R19695 VSS.n10208 VSS.n10207 0.00288205
R19696 VSS.n10268 VSS.n10267 0.00288205
R19697 VSS.n9340 VSS.n9339 0.00288205
R19698 VSS.n9202 VSS.n9201 0.00288205
R19699 VSS.n10090 VSS.n483 0.00287695
R19700 VSS.n11141 VSS.n11139 0.00287695
R19701 VSS.n10832 VSS.n10831 0.00287228
R19702 VSS.n9489 VSS.n1377 0.002865
R19703 VSS.n10440 VSS.n10335 0.00286014
R19704 VSS.n11115 VSS.n11053 0.00284094
R19705 VSS.n11114 VSS.n11113 0.00284094
R19706 VSS.n11112 VSS.n11111 0.00284094
R19707 VSS.n10046 VSS.n548 0.00282293
R19708 VSS.n9791 VSS.n789 0.002812
R19709 VSS.n9790 VSS.n787 0.002812
R19710 VSS.n11460 VSS.n13 0.00280492
R19711 VSS.n8952 VSS.n8951 0.00280297
R19712 VSS.n4803 VSS.n2503 0.00280297
R19713 VSS.n10788 VSS.n10735 0.00279891
R19714 VSS.n10110 VSS.n446 0.00278691
R19715 VSS.n485 VSS.n484 0.00278691
R19716 VSS.n10086 VSS.n488 0.00278691
R19717 VSS.n490 VSS.n489 0.00278691
R19718 VSS.n788 VSS.n786 0.00278398
R19719 VSS.n10081 VSS.n493 0.00276891
R19720 VSS.n10080 VSS.n10079 0.00276891
R19721 VSS.n10078 VSS.n494 0.00276891
R19722 VSS.n1462 VSS.n1461 0.00275596
R19723 VSS.n1456 VSS.n1455 0.00275596
R19724 VSS.n1459 VSS.n1427 0.00275596
R19725 VSS.n9780 VSS.n9779 0.00275596
R19726 VSS.n11123 VSS.n11122 0.0027509
R19727 VSS.n11032 VSS.n11031 0.0027509
R19728 VSS.n11120 VSS.n11033 0.0027509
R19729 VSS.n154 VSS.n151 0.00274194
R19730 VSS.n9507 VSS.n1336 0.00273506
R19731 VSS.n11321 VSS.n117 0.00273289
R19732 VSS.n11178 VSS.n11177 0.00267188
R19733 VSS.n11268 VSS.n11179 0.00267188
R19734 VSS.n11431 VSS.n36 0.00266998
R19735 VSS.n57 VSS.n54 0.00266998
R19736 VSS.n11398 VSS.n11395 0.00266998
R19737 VSS.n11429 VSS.n36 0.00266998
R19738 VSS.n11400 VSS.n54 0.00266998
R19739 VSS.n11395 VSS.n57 0.00266998
R19740 VSS.n10035 VSS.n10034 0.00266086
R19741 VSS.n9783 VSS.n9782 0.00265787
R19742 VSS.n9785 VSS.n9784 0.00265787
R19743 VSS.n9788 VSS.n790 0.00265787
R19744 VSS.n9787 VSS.n789 0.00265787
R19745 VSS.n10776 VSS.n10775 0.00265035
R19746 VSS.n10742 VSS.n10741 0.00265035
R19747 VSS.n10910 VSS.n228 0.0026461
R19748 VSS.n10913 VSS.n228 0.0026461
R19749 VSS.n1453 VSS.n1452 0.00264386
R19750 VSS.n1429 VSS.n1428 0.00264386
R19751 VSS.n9772 VSS.n9771 0.00264386
R19752 VSS.n9770 VSS.n9769 0.00264386
R19753 VSS.n9777 VSS.n795 0.00264386
R19754 VSS.n9776 VSS.n9775 0.00264386
R19755 VSS.n443 VSS.n442 0.00264286
R19756 VSS.n10112 VSS.n444 0.00264286
R19757 VSS.n487 VSS.n486 0.00260684
R19758 VSS.n10072 VSS.n499 0.00260684
R19759 VSS.n754 VSS.n753 0.00260182
R19760 VSS.n705 VSS.n704 0.00260182
R19761 VSS.n751 VSS.n706 0.00260182
R19762 VSS.n11197 VSS.n11196 0.00260182
R19763 VSS.n11259 VSS.n11258 0.00260182
R19764 VSS.n11257 VSS.n11256 0.00260182
R19765 VSS.n10076 VSS.n496 0.00257083
R19766 VSS.n11387 VSS.n81 0.00257045
R19767 VSS.n1454 VSS.n1453 0.00255979
R19768 VSS.n10829 VSS.n10828 0.00252989
R19769 VSS.n9488 VSS.n9476 0.00252714
R19770 VSS.n1298 VSS.n433 0.00251681
R19771 VSS.n462 VSS.n458 0.00251681
R19772 VSS.n10069 VSS.n503 0.00251681
R19773 VSS.n552 VSS.n548 0.00251681
R19774 VSS.n11150 VSS.n11149 0.00251681
R19775 VSS.n11466 VSS.n11465 0.00251681
R19776 VSS.n9782 VSS.n9781 0.00250374
R19777 VSS.n9798 VSS.n9795 0.00250374
R19778 VSS.n9797 VSS.n9796 0.00250374
R19779 VSS.n9799 VSS.n773 0.00250374
R19780 VSS.n11175 VSS.n11174 0.00250374
R19781 VSS.n11271 VSS.n11176 0.00250374
R19782 VSS.n156 VSS.n153 0.00248972
R19783 VSS.n11171 VSS.n11170 0.00248972
R19784 VSS.n11023 VSS.n11022 0.00248079
R19785 VSS.n11052 VSS.n11051 0.00248079
R19786 VSS.n10115 VSS.n441 0.00246279
R19787 VSS.n10090 VSS.n10089 0.00246279
R19788 VSS.n9779 VSS.n794 0.00244769
R19789 VSS.n11171 VSS.n153 0.00243368
R19790 VSS.n11170 VSS.n154 0.00243368
R19791 VSS.n9781 VSS.n9780 0.00241966
R19792 VSS.n9798 VSS.n9797 0.00241966
R19793 VSS.n9796 VSS.n773 0.00241966
R19794 VSS.n11273 VSS.n11174 0.00241966
R19795 VSS.n11176 VSS.n11175 0.00241966
R19796 VSS.n11271 VSS.n11270 0.00241966
R19797 VSS.n10655 VSS.n10654 0.00239047
R19798 VSS.n11137 VSS.n202 0.00237275
R19799 VSS.n204 VSS.n203 0.00237275
R19800 VSS.n11135 VSS.n11134 0.00237275
R19801 VSS.n11128 VSS.n11024 0.00235474
R19802 VSS.n11026 VSS.n11025 0.00235474
R19803 VSS.n9583 VSS.n796 0.0023496
R19804 VSS.n11161 VSS.n157 0.0023496
R19805 VSS.n518 VSS.n517 0.00233673
R19806 VSS.n521 VSS.n519 0.00233673
R19807 VSS.n524 VSS.n523 0.00233673
R19808 VSS.n522 VSS.n516 0.00233673
R19809 VSS.n753 VSS.n704 0.00232158
R19810 VSS.n706 VSS.n705 0.00232158
R19811 VSS.n11259 VSS.n11197 0.00232158
R19812 VSS.n11258 VSS.n11257 0.00232158
R19813 VSS.n11256 VSS.n11255 0.00232158
R19814 VSS.n1312 VSS.n433 0.00231873
R19815 VSS.n1302 VSS.n1301 0.00231873
R19816 VSS.n1304 VSS.n1303 0.00231873
R19817 VSS.n11150 VSS.n184 0.00231873
R19818 VSS.n11322 VSS.n11321 0.00231873
R19819 VSS.n762 VSS.n694 0.00230757
R19820 VSS.n1343 VSS.n1342 0.00229324
R19821 VSS.n9501 VSS.n9500 0.00229324
R19822 VSS.n1452 VSS.n1428 0.00227954
R19823 VSS.n9771 VSS.n9770 0.00227954
R19824 VSS.n9777 VSS.n9776 0.00227954
R19825 VSS.n9775 VSS.n9774 0.00227954
R19826 VSS.n10574 VSS.n10556 0.00227907
R19827 VSS.n9785 VSS.n9783 0.00226553
R19828 VSS.n9784 VSS.n790 0.00226553
R19829 VSS.n9788 VSS.n9787 0.00226553
R19830 VSS.n10037 VSS.n236 0.00226471
R19831 VSS.n11270 VSS.n11177 0.00225152
R19832 VSS.n11179 VSS.n11178 0.00225152
R19833 VSS.n11268 VSS.n11267 0.00225152
R19834 VSS.n10075 VSS.n10074 0.0022467
R19835 VSS.n498 VSS.n497 0.0022467
R19836 VSS.n10857 VSS.n246 0.00223077
R19837 VSS.n556 VSS.n555 0.00222869
R19838 VSS.n10039 VSS.n557 0.00222869
R19839 VSS.n1340 VSS.n1339 0.00221528
R19840 VSS.n9504 VSS.n9503 0.00221528
R19841 VSS.n11093 VSS.n9 0.00219268
R19842 VSS.n751 VSS.n750 0.00218146
R19843 VSS.n10095 VSS.n458 0.00217467
R19844 VSS.n1455 VSS.n1427 0.00216745
R19845 VSS.n1459 VSS.n1458 0.00216745
R19846 VSS.n10870 VSS.n10869 0.00215666
R19847 VSS.n9769 VSS.n9768 0.00213942
R19848 VSS.n9795 VSS.n786 0.00213942
R19849 VSS.n10885 VSS.n10884 0.00213866
R19850 VSS.n10879 VSS.n10878 0.00213866
R19851 VSS.n10883 VSS.n10880 0.00213866
R19852 VSS.n10035 VSS.n560 0.00212065
R19853 VSS.n11118 VSS.n11117 0.00212065
R19854 VSS.n11465 VSS.n10 0.00212065
R19855 VSS.n12 VSS.n11 0.00212065
R19856 VSS.n9791 VSS.n9790 0.0021114
R19857 VSS.n10537 VSS.n10492 0.00208665
R19858 VSS.n10108 VSS.n448 0.00208463
R19859 VSS.n1422 VSS.n1421 0.00206936
R19860 VSS.n9590 VSS.n9566 0.00206936
R19861 VSS.n9803 VSS.n9800 0.00206936
R19862 VSS.n698 VSS.n694 0.00206936
R19863 VSS.n11155 VSS.n11154 0.00206936
R19864 VSS.n11139 VSS.n11138 0.00204862
R19865 VSS.n11119 VSS.n11034 0.00204862
R19866 VSS.n11036 VSS.n11035 0.00204862
R19867 VSS.n11277 VSS.n151 0.00204134
R19868 VSS.n11196 VSS.n11195 0.00204134
R19869 VSS.n1461 VSS.n1426 0.00202732
R19870 VSS.n9772 VSS.n796 0.00202732
R19871 VSS.n10053 VSS.n543 0.0019946
R19872 VSS.n545 VSS.n544 0.0019946
R19873 VSS.n10051 VSS.n10050 0.0019946
R19874 VSS.n9502 VSS.n1341 0.00198137
R19875 VSS.n10921 VSS.n223 0.00196707
R19876 VSS.n11165 VSS.n11163 0.00195726
R19877 VSS.n11164 VSS.n155 0.00195726
R19878 VSS.n11168 VSS.n11167 0.00195726
R19879 VSS.n9499 VSS.n9498 0.00195539
R19880 VSS.n11172 VSS.n152 0.00194325
R19881 VSS.n11274 VSS.n11173 0.00194325
R19882 VSS.n1370 VSS.n1369 0.00193729
R19883 VSS.n9634 VSS.n9633 0.00193729
R19884 VSS.n9745 VSS.n9744 0.00193729
R19885 VSS.n9723 VSS.n9722 0.00193729
R19886 VSS.n10008 VSS.n10007 0.00193729
R19887 VSS.n9986 VSS.n9985 0.00193729
R19888 VSS.n9802 VSS.n9801 0.00192924
R19889 VSS.n9805 VSS.n772 0.00192924
R19890 VSS.n9808 VSS.n9807 0.00192924
R19891 VSS.n9806 VSS.n771 0.00192924
R19892 VSS.n10868 VSS.n10867 0.00192857
R19893 VSS.n11315 VSS.n109 0.00192857
R19894 VSS.n11389 VSS.n62 0.00192857
R19895 VSS.n11393 VSS.n56 0.00192857
R19896 VSS.n11319 VSS.n120 0.00192857
R19897 VSS.n11432 VSS.n34 0.00192857
R19898 VSS.n10707 VSS.n10706 0.00192857
R19899 VSS.n10499 VSS.n10493 0.00192857
R19900 VSS.n11313 VSS.n122 0.00192857
R19901 VSS.n10565 VSS.n10563 0.00192857
R19902 VSS.n10865 VSS.n229 0.00192857
R19903 VSS.n10096 VSS.n10095 0.00192257
R19904 VSS.n10820 VSS.n10819 0.00191848
R19905 VSS.n9468 VSS.n9467 0.00191573
R19906 VSS.n1421 VSS.n1420 0.00191523
R19907 VSS.n1425 VSS.n1424 0.00191523
R19908 VSS.n1463 VSS.n1462 0.00191523
R19909 VSS.n11154 VSS.n178 0.00191523
R19910 VSS.n10044 VSS.n550 0.00190456
R19911 VSS.n554 VSS.n553 0.00190456
R19912 VSS.n10042 VSS.n10041 0.00190456
R19913 VSS.n11466 VSS.n9 0.00190456
R19914 VSS.n9463 VSS.n9462 0.00190156
R19915 VSS.n9793 VSS.n787 0.00185918
R19916 VSS.n9792 VSS.n788 0.00185918
R19917 VSS.n462 VSS.n461 0.00185054
R19918 VSS.n10093 VSS.n459 0.00185054
R19919 VSS.n10092 VSS.n460 0.00185054
R19920 VSS.n11325 VSS.n116 0.00185054
R19921 VSS.n10592 VSS.n10591 0.00185034
R19922 VSS.n702 VSS.n701 0.00184517
R19923 VSS.n755 VSS.n703 0.00184517
R19924 VSS.n10531 VSS.n10530 0.00181658
R19925 VSS.n1318 VSS.n1317 0.00181453
R19926 VSS.n11110 VSS.n11054 0.00181453
R19927 VSS.n11056 VSS.n11055 0.00181453
R19928 VSS.n11108 VSS.n11107 0.00181453
R19929 VSS.n11058 VSS.n11057 0.00181453
R19930 VSS.n11105 VSS.n11059 0.00181453
R19931 VSS.n9595 VSS.n9566 0.00180313
R19932 VSS.n9102 VSS.n9100 0.00180205
R19933 VSS.n861 VSS.n860 0.00180205
R19934 VSS.n1107 VSS.n1106 0.00180205
R19935 VSS.n1049 VSS.n926 0.00180205
R19936 VSS.n1000 VSS.n999 0.00180205
R19937 VSS.n11353 VSS.n100 0.00180205
R19938 VSS.n11369 VSS.n88 0.00180205
R19939 VSS.n1199 VSS.n1198 0.00180205
R19940 VSS.n9414 VSS.n9413 0.00180205
R19941 VSS.n9257 VSS.n1511 0.00180205
R19942 VSS.n11339 VSS.n11338 0.00179403
R19943 VSS.n1311 VSS.n1297 0.00177851
R19944 VSS.n1313 VSS.n1312 0.00177851
R19945 VSS.n10882 VSS.n184 0.00177851
R19946 VSS.n732 VSS.n731 0.00177511
R19947 VSS.n737 VSS.n736 0.00177511
R19948 VSS.n735 VSS.n734 0.00177511
R19949 VSS.n9002 VSS.n9001 0.00176761
R19950 VSS.n1134 VSS.n1131 0.00176761
R19951 VSS.n1082 VSS.n913 0.00176761
R19952 VSS.n1033 VSS.n1032 0.00176761
R19953 VSS.n975 VSS.n952 0.00176761
R19954 VSS.n11002 VSS.n10999 0.00176761
R19955 VSS.n10974 VSS.n10973 0.00176761
R19956 VSS.n9550 VSS.n9548 0.00176761
R19957 VSS.n9357 VSS.n9355 0.00176761
R19958 VSS.n9169 VSS.n9168 0.00176761
R19959 VSS.n11262 VSS.n11261 0.00176109
R19960 VSS.n10744 VSS.n10743 0.00175874
R19961 VSS.n1450 VSS.n1438 0.00173307
R19962 VSS.n1119 VSS.n900 0.00172754
R19963 VSS.n1070 VSS.n1069 0.00172754
R19964 VSS.n1012 VSS.n939 0.00172754
R19965 VSS.n10921 VSS.n10915 0.00172754
R19966 VSS.n10937 VSS.n212 0.00172754
R19967 VSS.n9535 VSS.n1219 0.00172754
R19968 VSS.n9291 VSS.n9290 0.00172754
R19969 VSS.n9131 VSS.n9130 0.00172754
R19970 VSS.n1309 VSS.n1298 0.00170648
R19971 VSS.n1308 VSS.n1307 0.00170648
R19972 VSS.n1306 VSS.n1299 0.00170648
R19973 VSS.n11162 VSS.n11161 0.00170504
R19974 VSS.n11181 VSS.n11180 0.00170504
R19975 VSS.n11265 VSS.n11182 0.00170504
R19976 VSS.n558 VSS.n237 0.00168848
R19977 VSS.n10806 VSS.n10804 0.00168421
R19978 VSS.n10800 VSS.n10798 0.00168421
R19979 VSS.n10630 VSS.n10629 0.00168421
R19980 VSS.n10626 VSS.n10625 0.00168421
R19981 VSS.n10621 VSS.n10620 0.00168421
R19982 VSS.n10617 VSS.n10616 0.00168421
R19983 VSS.n10385 VSS.n10384 0.00168421
R19984 VSS.n10381 VSS.n10380 0.00168421
R19985 VSS.n10376 VSS.n10375 0.00168421
R19986 VSS.n10302 VSS.n10299 0.00168421
R19987 VSS.n10681 VSS.n10297 0.00168421
R19988 VSS.n10684 VSS.n10294 0.00168421
R19989 VSS.n9813 VSS.n9810 0.00167702
R19990 VSS.n10837 VSS.n10836 0.00167391
R19991 VSS.n10826 VSS.n10825 0.00167391
R19992 VSS.n10895 VSS.n10894 0.00167047
R19993 VSS.n9836 VSS.n9834 0.00166301
R19994 VSS.n9835 VSS.n763 0.00166301
R19995 VSS.n9838 VSS.n9837 0.00166301
R19996 VSS.n559 VSS.n558 0.00165246
R19997 VSS.n10049 VSS.n10048 0.00163445
R19998 VSS.n10105 VSS.n10104 0.00161645
R19999 VSS.n453 VSS.n452 0.00161645
R20000 VSS.n10103 VSS.n454 0.00161645
R20001 VSS.n201 VSS.n188 0.00161645
R20002 VSS.n9597 VSS.n9595 0.00160696
R20003 VSS.n11142 VSS.n201 0.00159844
R20004 VSS.n760 VSS.n696 0.00159295
R20005 VSS.n700 VSS.n699 0.00159295
R20006 VSS.n758 VSS.n757 0.00159295
R20007 VSS.n10102 VSS.n455 0.00158043
R20008 VSS.n560 VSS.n559 0.00158043
R20009 VSS.n10766 VSS.n10765 0.00156599
R20010 VSS.n10762 VSS.n10761 0.00155167
R20011 VSS.n9590 VSS.n9589 0.00155091
R20012 VSS.n9593 VSS.n9567 0.00155091
R20013 VSS.n9592 VSS.n9588 0.00155091
R20014 VSS.n10869 VSS.n237 0.00154442
R20015 VSS.n10819 VSS.n10812 0.00152717
R20016 VSS.n1417 VSS.n1416 0.00152289
R20017 VSS.n11254 VSS.n11198 0.00152289
R20018 VSS.n11200 VSS.n11199 0.00152289
R20019 VSS.n11252 VSS.n11251 0.00152289
R20020 VSS.n11202 VSS.n11201 0.00152289
R20021 VSS.n9584 VSS.n9581 0.00150887
R20022 VSS.n10789 VSS.n10788 0.00150272
R20023 VSS.n1471 VSS.n1470 0.00149486
R20024 VSS.n1420 VSS.n1419 0.00149486
R20025 VSS.n733 VSS.n178 0.00149486
R20026 VSS.n11088 VSS.n11087 0.0014904
R20027 VSS.n11096 VSS.n11089 0.0014904
R20028 VSS.n11095 VSS.n11090 0.0014904
R20029 VSS.n11092 VSS.n11091 0.0014904
R20030 VSS.n118 VSS.n117 0.0014904
R20031 VSS.n1468 VSS.n1422 0.00143881
R20032 VSS.n1467 VSS.n1466 0.00143881
R20033 VSS.n1465 VSS.n1423 0.00143881
R20034 VSS.n10886 VSS.n10877 0.00143638
R20035 VSS.n466 VSS.n465 0.00141837
R20036 VSS.n726 VSS.n725 0.00141079
R20037 VSS.n531 VSS.n527 0.00140036
R20038 VSS.n530 VSS.n529 0.00140036
R20039 VSS.n528 VSS.n513 0.00140036
R20040 VSS.n10063 VSS.n514 0.00140036
R20041 VSS.n533 VSS.n515 0.00140036
R20042 VSS.n10754 VSS.n10746 0.00139161
R20043 VSS.n9841 VSS.n692 0.00138277
R20044 VSS.n1447 VSS.n1446 0.00136875
R20045 VSS.n1443 VSS.n1442 0.00136875
R20046 VSS.n1445 VSS.n1444 0.00136875
R20047 VSS.n173 VSS.n159 0.00136875
R20048 VSS.n174 VSS.n173 0.00135474
R20049 VSS.n1388 VSS.n1385 0.00135106
R20050 VSS.n1331 VSS.n1330 0.00135106
R20051 VSS.n11149 VSS.n185 0.00134634
R20052 VSS.n187 VSS.n186 0.00134634
R20053 VSS.n11147 VSS.n11146 0.00134634
R20054 VSS.n10538 VSS.n10537 0.00134396
R20055 VSS.n9601 VSS.n827 0.00134073
R20056 VSS.n11303 VSS.n129 0.00130178
R20057 VSS.n10844 VSS.n10698 0.00130178
R20058 VSS.n10853 VSS.n247 0.00128671
R20059 VSS.n11237 VSS.n0 0.00128468
R20060 VSS.n10047 VSS.n10046 0.00127431
R20061 VSS.n11232 VSS.n11231 0.00127067
R20062 VSS.n11240 VSS.n11233 0.00127067
R20063 VSS.n11239 VSS.n11234 0.00127067
R20064 VSS.n11236 VSS.n11235 0.00127067
R20065 VSS.n11429 VSS.n31 0.00125937
R20066 VSS.n1337 VSS.n1335 0.00125368
R20067 VSS.n9507 VSS.n9506 0.00125368
R20068 VSS.n9498 VSS.n1344 0.00125368
R20069 VSS.n10835 VSS.n10834 0.0012337
R20070 VSS.n739 VSS.n730 0.00122863
R20071 VSS.n457 VSS.n456 0.00122029
R20072 VSS.n10100 VSS.n10099 0.00122029
R20073 VSS.n10098 VSS.n10097 0.00122029
R20074 VSS.n9581 VSS.n9568 0.00121462
R20075 VSS.n10666 VSS.n10665 0.0012124
R20076 VSS.n10428 VSS.n10427 0.0012124
R20077 VSS.n10465 VSS.n10464 0.00121146
R20078 VSS.n552 VSS.n551 0.00120228
R20079 VSS.n10045 VSS.n549 0.00120228
R20080 VSS.n9812 VSS.n9811 0.00120061
R20081 VSS.n9815 VSS.n770 0.00120061
R20082 VSS.n9819 VSS.n9818 0.00120061
R20083 VSS.n9817 VSS.n769 0.00120061
R20084 VSS.n464 VSS.n463 0.00118427
R20085 VSS.n11099 VSS.n11098 0.00116627
R20086 VSS.n11157 VSS.n11155 0.00115857
R20087 VSS.n11156 VSS.n158 0.00115857
R20088 VSS.n11159 VSS.n11158 0.00115857
R20089 VSS.n10586 VSS.n10585 0.0011338
R20090 VSS.n1300 VSS.n1299 0.00111224
R20091 VSS.n465 VSS.n464 0.00111224
R20092 VSS.n527 VSS.n526 0.00111224
R20093 VSS.n10874 VSS.n10873 0.00111224
R20094 VSS.n10891 VSS.n10890 0.00111224
R20095 VSS.n10889 VSS.n10888 0.00111224
R20096 VSS.n10876 VSS.n10875 0.00111224
R20097 VSS.n9840 VSS.n762 0.00110252
R20098 VSS.n10915 VSS.n10913 0.0010988
R20099 VSS.n1364 VSS.n1363 0.00109183
R20100 VSS.n9761 VSS.n9760 0.00109183
R20101 VSS.n9739 VSS.n9738 0.00109183
R20102 VSS.n10027 VSS.n10026 0.00109183
R20103 VSS.n10002 VSS.n10001 0.00109183
R20104 VSS.n9980 VSS.n9979 0.00109183
R20105 VSS.n11387 VSS.n11382 0.00108231
R20106 VSS.n1296 VSS.n1272 0.00107623
R20107 VSS.n1317 VSS.n1316 0.00107623
R20108 VSS.n1315 VSS.n1273 0.00107623
R20109 VSS.n10870 VSS.n236 0.00107623
R20110 VSS.n9600 VSS.n9599 0.00106049
R20111 VSS.n829 VSS.n828 0.00106049
R20112 VSS.n9598 VSS.n830 0.00106049
R20113 VSS.n11317 VSS.n59 0.00104767
R20114 VSS.n698 VSS.n697 0.00104647
R20115 VSS.n761 VSS.n695 0.00104647
R20116 VSS.n11249 VSS.n11204 0.00104647
R20117 VSS.n10070 VSS.n10069 0.00102221
R20118 VSS.n10061 VSS.n10060 0.00102221
R20119 VSS.n9505 VSS.n1338 0.00101978
R20120 VSS.n11243 VSS.n11242 0.00101845
R20121 VSS.n10733 VSS.n10732 0.000993001
R20122 VSS.n755 VSS.n754 0.000976413
R20123 VSS.n746 VSS.n745 0.000976413
R20124 VSS.n728 VSS.n727 0.000976413
R20125 VSS.n743 VSS.n729 0.000976413
R20126 VSS.n742 VSS.n740 0.000976413
R20127 VSS.n11167 VSS.n156 0.000976413
R20128 VSS.n11204 VSS.n11203 0.000976413
R20129 VSS.n10059 VSS.n537 0.000968187
R20130 VSS.n539 VSS.n538 0.000968187
R20131 VSS.n10057 VSS.n10056 0.000968187
R20132 VSS.n541 VSS.n540 0.000968187
R20133 VSS.n10054 VSS.n542 0.000968187
R20134 VSS.n10038 VSS.n10037 0.000968187
R20135 VSS.n1475 VSS.n1403 0.000948389
R20136 VSS.n1418 VSS.n1417 0.000948389
R20137 VSS.n1473 VSS.n1472 0.000948389
R20138 VSS.n10534 VSS.n10533 0.00093886
R20139 VSS.n1366 VSS.n1349 0.000922734
R20140 VSS.n9764 VSS.n9763 0.000922734
R20141 VSS.n9741 VSS.n9666 0.000922734
R20142 VSS.n10030 VSS.n10029 0.000922734
R20143 VSS.n10004 VSS.n147 0.000922734
R20144 VSS.n9982 VSS.n138 0.000922734
R20145 VSS.n10758 VSS.n10757 0.000920842
R20146 VSS.n9887 VSS.n647 0.00091958
R20147 VSS.n1176 VSS.n1175 0.00091958
R20148 VSS.n1180 VSS.n1174 0.00091958
R20149 VSS.n672 VSS.n671 0.00091958
R20150 VSS.n9521 VSS.n1236 0.00091958
R20151 VSS.n9892 VSS.n643 0.00091958
R20152 VSS.n624 VSS.n623 0.00091958
R20153 VSS.n626 VSS.n625 0.00091958
R20154 VSS.n9916 VSS.n9915 0.00091958
R20155 VSS.n11284 VSS.n11283 0.00091958
R20156 VSS.n143 VSS.n142 0.00091958
R20157 VSS.n1234 VSS.n1233 0.00091958
R20158 VSS.n10107 VSS.n449 0.000914166
R20159 VSS.n451 VSS.n450 0.000914166
R20160 VSS.n479 VSS.n478 0.000914166
R20161 VSS.n11145 VSS.n11144 0.000914166
R20162 VSS.n11322 VSS.n116 0.000914166
R20163 VSS.n9800 VSS.n9799 0.000906352
R20164 VSS.n11118 VSS.n11038 0.000896158
R20165 VSS.n10808 VSS.n10793 0.000866848
R20166 VSS.n9826 VSS.n9825 0.000864316
R20167 VSS.n9824 VSS.n765 0.000864316
R20168 VSS.n9831 VSS.n9828 0.000864316
R20169 VSS.n9830 VSS.n9829 0.000864316
R20170 VSS.n9833 VSS.n764 0.000864316
R20171 VSS.n11104 VSS.n11078 0.00082413
R20172 VSS.n1449 VSS.n1439 0.000822279
R20173 VSS.n1441 VSS.n1440 0.000822279
R20174 VSS.n9587 VSS.n9586 0.000822279
R20175 VSS.n177 VSS.n176 0.000822279
R20176 VSS.n11264 VSS.n11262 0.000808267
R20177 VSS.n10730 VSS.n10701 0.000773889
R20178 VSS.n10840 VSS.n10839 0.000769022
R20179 VSS.n11248 VSS.n11223 0.000752219
R20180 VSS.n10893 VSS.n10872 0.000752101
R20181 VSS.n11027 VSS.n11026 0.000752101
R20182 VSS.n11086 VSS.n11085 0.000752101
R20183 VSS.n11295 VSS.n11294 0.000742997
R20184 VSS.n134 VSS.n133 0.000742997
R20185 VSS.n9823 VSS.n9822 0.000710182
R20186 VSS.n10532 VSS.n10531 0.000702551
R20187 VSS.n10349 VSS.n10348 0.000702551
R20188 VSS.n1458 VSS.n1454 0.00069617
R20189 VSS.n9774 VSS.n794 0.00069617
R20190 VSS.n9822 VSS.n9821 0.00069617
R20191 VSS.n11308 VSS.n127 0.000688976
R20192 VSS.n10115 VSS.n10114 0.000680072
R20193 VSS.n10087 VSS.n487 0.000680072
R20194 VSS.n10064 VSS.n10063 0.000680072
R20195 VSS.n10034 VSS.n235 0.000680072
R20196 VSS.n11129 VSS.n11023 0.000680072
R20197 VSS.n1456 VSS.n1426 0.000640121
R20198 VSS.n9768 VSS.n795 0.000640121
R20199 VSS.n9819 VSS.n9816 0.000640121
R20200 VSS.n750 VSS.n749 0.000640121
R20201 VSS.n11277 VSS.n11276 0.000640121
R20202 VSS.n11081 VSS.n11079 0.00062605
R20203 VSS.n10830 VSS.n10810 0.000622283
R20204 VSS.n10770 VSS.n246 0.000604895
R20205 VSS.n9693 VSS.n9671 0.000604895
R20206 VSS.n9673 VSS.n9672 0.000604895
R20207 VSS.n9692 VSS.n9691 0.000604895
R20208 VSS.n9690 VSS.n9674 0.000604895
R20209 VSS.n9676 VSS.n9675 0.000604895
R20210 VSS.n9689 VSS.n9688 0.000604895
R20211 VSS.n9687 VSS.n9677 0.000604895
R20212 VSS.n9679 VSS.n9678 0.000604895
R20213 VSS.n9686 VSS.n9685 0.000604895
R20214 VSS.n9684 VSS.n9680 0.000604895
R20215 VSS.n9682 VSS.n9681 0.000604895
R20216 VSS.n9683 VSS.n653 0.000604895
R20217 VSS.n1177 VSS.n654 0.000604895
R20218 VSS.n1175 VSS.n1174 0.000604895
R20219 VSS.n1179 VSS.n1178 0.000604895
R20220 VSS.n9853 VSS.n680 0.000604895
R20221 VSS.n682 VSS.n681 0.000604895
R20222 VSS.n9852 VSS.n9851 0.000604895
R20223 VSS.n9850 VSS.n683 0.000604895
R20224 VSS.n685 VSS.n684 0.000604895
R20225 VSS.n9849 VSS.n9848 0.000604895
R20226 VSS.n9847 VSS.n686 0.000604895
R20227 VSS.n688 VSS.n687 0.000604895
R20228 VSS.n9846 VSS.n9845 0.000604895
R20229 VSS.n9844 VSS.n689 0.000604895
R20230 VSS.n691 VSS.n690 0.000604895
R20231 VSS.n9843 VSS.n9842 0.000604895
R20232 VSS.n604 VSS.n546 0.000604895
R20233 VSS.n603 VSS.n602 0.000604895
R20234 VSS.n605 VSS.n601 0.000604895
R20235 VSS.n609 VSS.n606 0.000604895
R20236 VSS.n608 VSS.n607 0.000604895
R20237 VSS.n610 VSS.n600 0.000604895
R20238 VSS.n614 VSS.n611 0.000604895
R20239 VSS.n613 VSS.n612 0.000604895
R20240 VSS.n615 VSS.n599 0.000604895
R20241 VSS.n619 VSS.n616 0.000604895
R20242 VSS.n618 VSS.n617 0.000604895
R20243 VSS.n620 VSS.n598 0.000604895
R20244 VSS.n9906 VSS.n622 0.000604895
R20245 VSS.n625 VSS.n624 0.000604895
R20246 VSS.n9905 VSS.n9904 0.000604895
R20247 VSS.n9701 VSS.n9698 0.000604895
R20248 VSS.n9700 VSS.n9699 0.000604895
R20249 VSS.n9702 VSS.n9697 0.000604895
R20250 VSS.n9706 VSS.n9703 0.000604895
R20251 VSS.n9705 VSS.n9704 0.000604895
R20252 VSS.n9707 VSS.n9696 0.000604895
R20253 VSS.n9711 VSS.n9708 0.000604895
R20254 VSS.n9710 VSS.n9709 0.000604895
R20255 VSS.n9712 VSS.n9695 0.000604895
R20256 VSS.n9716 VSS.n9713 0.000604895
R20257 VSS.n9715 VSS.n9714 0.000604895
R20258 VSS.n9717 VSS.n9694 0.000604895
R20259 VSS.n10573 VSS.n10572 0.000604651
R20260 VSS.n9034 VSS.n9018 0.000603567
R20261 VSS.n9032 VSS.n1560 0.000603567
R20262 VSS.n10147 VSS.n403 0.000603567
R20263 VSS.n10145 VSS.n10144 0.000603567
R20264 VSS.n10207 VSS.n331 0.000603567
R20265 VSS.n10205 VSS.n10204 0.000603567
R20266 VSS.n10267 VSS.n259 0.000603567
R20267 VSS.n10265 VSS.n10264 0.000603567
R20268 VSS.n9339 VSS.n9322 0.000603567
R20269 VSS.n9337 VSS.n9336 0.000603567
R20270 VSS.n9201 VSS.n9185 0.000603567
R20271 VSS.n9199 VSS.n1522 0.000603567
R20272 VSS.n11226 VSS.n11224 0.000598085
R20273 VSS.n10793 VSS.n10792 0.000597826
R20274 VSS.n11083 VSS.n11082 0.000554022
R20275 VSS.n11102 VSS.n11079 0.000554022
R20276 VSS.n11101 VSS.n11080 0.000554022
R20277 VSS.n11085 VSS.n11084 0.000554022
R20278 VSS.n9882 VSS.n9881 0.000552448
R20279 VSS.n9854 VSS.n679 0.000552448
R20280 VSS.n9907 VSS.n621 0.000552448
R20281 VSS.n9903 VSS.n627 0.000552448
R20282 VSS.n11305 VSS.n11304 0.000547244
R20283 VSS.n11228 VSS.n11227 0.000542036
R20284 VSS.n11246 VSS.n11224 0.000542036
R20285 VSS.n11245 VSS.n11225 0.000542036
R20286 VSS.n11230 VSS.n11229 0.000542036
R20287 VSS.n10528 VSS.n10498 0.000533758
R20288 VSS.n9493 VSS.n9492 0.000525989
R20289 VSS.n479 VSS.n466 0.000518007
R20290 VSS.n483 VSS.n463 0.000518007
R20291 VSS.n11144 VSS.n188 0.000518007
R20292 VSS.n11142 VSS.n11141 0.000518007
R20293 VSS.n9586 VSS.n9568 0.000514012
R20294 VSS.n9584 VSS.n9583 0.000514012
R20295 VSS.n176 VSS.n159 0.000514012
R20296 VSS.n174 VSS.n157 0.000514012
R20297 a_52635_34067.t59 a_52635_34067.t62 9.46371
R20298 a_52635_34067.t12 a_52635_34067.t35 8.7152
R20299 a_52635_34067.t22 a_52635_34067.t39 8.7152
R20300 a_52635_34067.n7 a_52635_34067.t133 9.1601
R20301 a_52635_34067.n9 a_52635_34067.t234 9.1601
R20302 a_52635_34067.n13 a_52635_34067.t176 9.17607
R20303 a_52635_34067.n24 a_52635_34067.t121 9.17607
R20304 a_52635_34067.n109 a_52635_34067.t228 8.10567
R20305 a_52635_34067.n92 a_52635_34067.t159 8.10567
R20306 a_52635_34067.n92 a_52635_34067.t98 8.10567
R20307 a_52635_34067.n92 a_52635_34067.t233 8.10567
R20308 a_52635_34067.n92 a_52635_34067.t163 8.10567
R20309 a_52635_34067.n55 a_52635_34067.t169 8.10567
R20310 a_52635_34067.n55 a_52635_34067.t175 8.10567
R20311 a_52635_34067.n55 a_52635_34067.t114 8.10567
R20312 a_52635_34067.n55 a_52635_34067.t201 8.10567
R20313 a_52635_34067.n60 a_52635_34067.t177 8.10567
R20314 a_52635_34067.n60 a_52635_34067.t160 8.10567
R20315 a_52635_34067.n60 a_52635_34067.t99 8.10567
R20316 a_52635_34067.n60 a_52635_34067.t183 8.10567
R20317 a_52635_34067.n90 a_52635_34067.t209 8.10567
R20318 a_52635_34067.n90 a_52635_34067.t100 8.10567
R20319 a_52635_34067.n90 a_52635_34067.t223 8.10567
R20320 a_52635_34067.n58 a_52635_34067.t222 8.10567
R20321 a_52635_34067.n58 a_52635_34067.t118 8.10567
R20322 a_52635_34067.n58 a_52635_34067.t102 8.10567
R20323 a_52635_34067.n109 a_52635_34067.t198 8.10567
R20324 a_52635_34067.n109 a_52635_34067.t129 8.10567
R20325 a_52635_34067.n109 a_52635_34067.t197 8.10567
R20326 a_52635_34067.n116 a_52635_34067.t224 8.10567
R20327 a_52635_34067.n107 a_52635_34067.t149 8.10567
R20328 a_52635_34067.n107 a_52635_34067.t88 8.10567
R20329 a_52635_34067.n107 a_52635_34067.t232 8.10567
R20330 a_52635_34067.n107 a_52635_34067.t155 8.10567
R20331 a_52635_34067.n74 a_52635_34067.t161 8.10567
R20332 a_52635_34067.n74 a_52635_34067.t165 8.10567
R20333 a_52635_34067.n74 a_52635_34067.t106 8.10567
R20334 a_52635_34067.n74 a_52635_34067.t194 8.10567
R20335 a_52635_34067.n75 a_52635_34067.t168 8.10567
R20336 a_52635_34067.n75 a_52635_34067.t151 8.10567
R20337 a_52635_34067.n75 a_52635_34067.t93 8.10567
R20338 a_52635_34067.n75 a_52635_34067.t174 8.10567
R20339 a_52635_34067.n102 a_52635_34067.t162 8.10567
R20340 a_52635_34067.n102 a_52635_34067.t238 8.10567
R20341 a_52635_34067.n102 a_52635_34067.t189 8.10567
R20342 a_52635_34067.n100 a_52635_34067.t182 8.10567
R20343 a_52635_34067.n100 a_52635_34067.t79 8.10567
R20344 a_52635_34067.n100 a_52635_34067.t65 8.10567
R20345 a_52635_34067.n116 a_52635_34067.t187 8.10567
R20346 a_52635_34067.n116 a_52635_34067.t123 8.10567
R20347 a_52635_34067.n116 a_52635_34067.t185 8.10567
R20348 a_52635_34067.n111 a_52635_34067.t179 8.10567
R20349 a_52635_34067.n95 a_52635_34067.t105 8.10567
R20350 a_52635_34067.n95 a_52635_34067.t225 8.10567
R20351 a_52635_34067.n95 a_52635_34067.t195 8.10567
R20352 a_52635_34067.n95 a_52635_34067.t112 8.10567
R20353 a_52635_34067.n64 a_52635_34067.t116 8.10567
R20354 a_52635_34067.n64 a_52635_34067.t120 8.10567
R20355 a_52635_34067.n64 a_52635_34067.t235 8.10567
R20356 a_52635_34067.n64 a_52635_34067.t140 8.10567
R20357 a_52635_34067.n68 a_52635_34067.t122 8.10567
R20358 a_52635_34067.n68 a_52635_34067.t109 8.10567
R20359 a_52635_34067.n68 a_52635_34067.t226 8.10567
R20360 a_52635_34067.n68 a_52635_34067.t127 8.10567
R20361 a_52635_34067.n88 a_52635_34067.t146 8.10567
R20362 a_52635_34067.n88 a_52635_34067.t229 8.10567
R20363 a_52635_34067.n88 a_52635_34067.t171 8.10567
R20364 a_52635_34067.n86 a_52635_34067.t164 8.10567
R20365 a_52635_34067.n86 a_52635_34067.t66 8.10567
R20366 a_52635_34067.n86 a_52635_34067.t231 8.10567
R20367 a_52635_34067.n111 a_52635_34067.t137 8.10567
R20368 a_52635_34067.n111 a_52635_34067.t77 8.10567
R20369 a_52635_34067.n111 a_52635_34067.t136 8.10567
R20370 a_52635_34067.n112 a_52635_34067.t145 8.10567
R20371 a_52635_34067.n104 a_52635_34067.t72 8.10567
R20372 a_52635_34067.n104 a_52635_34067.t205 8.10567
R20373 a_52635_34067.n104 a_52635_34067.t158 8.10567
R20374 a_52635_34067.n104 a_52635_34067.t81 8.10567
R20375 a_52635_34067.n82 a_52635_34067.t83 8.10567
R20376 a_52635_34067.n82 a_52635_34067.t89 8.10567
R20377 a_52635_34067.n82 a_52635_34067.t217 8.10567
R20378 a_52635_34067.n82 a_52635_34067.t113 8.10567
R20379 a_52635_34067.n79 a_52635_34067.t92 8.10567
R20380 a_52635_34067.n79 a_52635_34067.t76 8.10567
R20381 a_52635_34067.n79 a_52635_34067.t206 8.10567
R20382 a_52635_34067.n79 a_52635_34067.t97 8.10567
R20383 a_52635_34067.n98 a_52635_34067.t86 8.10567
R20384 a_52635_34067.n98 a_52635_34067.t170 8.10567
R20385 a_52635_34067.n98 a_52635_34067.t111 8.10567
R20386 a_52635_34067.n96 a_52635_34067.t104 8.10567
R20387 a_52635_34067.n96 a_52635_34067.t191 8.10567
R20388 a_52635_34067.n96 a_52635_34067.t172 8.10567
R20389 a_52635_34067.n112 a_52635_34067.t110 8.10567
R20390 a_52635_34067.n112 a_52635_34067.t227 8.10567
R20391 a_52635_34067.n112 a_52635_34067.t108 8.10567
R20392 a_52635_34067.n19 a_52635_34067.t188 8.10567
R20393 a_52635_34067.n19 a_52635_34067.t196 8.10567
R20394 a_52635_34067.n19 a_52635_34067.t128 8.10567
R20395 a_52635_34067.n19 a_52635_34067.t216 8.10567
R20396 a_52635_34067.n11 a_52635_34067.t193 8.10567
R20397 a_52635_34067.n177 a_52635_34067.t84 8.10567
R20398 a_52635_34067.n176 a_52635_34067.t214 8.10567
R20399 a_52635_34067.n12 a_52635_34067.t115 8.10567
R20400 a_52635_34067.n12 a_52635_34067.t69 8.10567
R20401 a_52635_34067.n12 a_52635_34067.t181 8.10567
R20402 a_52635_34067.n1 a_52635_34067.t240 8.10567
R20403 a_52635_34067.n1 a_52635_34067.t213 8.10567
R20404 a_52635_34067.n1 a_52635_34067.t144 8.10567
R20405 a_52635_34067.n41 a_52635_34067.t210 8.10567
R20406 a_52635_34067.n175 a_52635_34067.t101 8.10567
R20407 a_52635_34067.n174 a_52635_34067.t85 8.10567
R20408 a_52635_34067.n16 a_52635_34067.t199 8.10567
R20409 a_52635_34067.n16 a_52635_34067.t178 8.10567
R20410 a_52635_34067.n42 a_52635_34067.t117 8.10567
R20411 a_52635_34067.n42 a_52635_34067.t203 8.10567
R20412 a_52635_34067.n36 a_52635_34067.t143 8.10567
R20413 a_52635_34067.n36 a_52635_34067.t148 8.10567
R20414 a_52635_34067.n36 a_52635_34067.t87 8.10567
R20415 a_52635_34067.n36 a_52635_34067.t173 8.10567
R20416 a_52635_34067.n5 a_52635_34067.t180 8.10567
R20417 a_52635_34067.n155 a_52635_34067.t78 8.10567
R20418 a_52635_34067.n154 a_52635_34067.t207 8.10567
R20419 a_52635_34067.n6 a_52635_34067.t70 8.10567
R20420 a_52635_34067.n6 a_52635_34067.t221 8.10567
R20421 a_52635_34067.n6 a_52635_34067.t139 8.10567
R20422 a_52635_34067.n27 a_52635_34067.t215 8.10567
R20423 a_52635_34067.n27 a_52635_34067.t167 8.10567
R20424 a_52635_34067.n27 a_52635_34067.t107 8.10567
R20425 a_52635_34067.n51 a_52635_34067.t202 8.10567
R20426 a_52635_34067.n153 a_52635_34067.t95 8.10567
R20427 a_52635_34067.n152 a_52635_34067.t80 8.10567
R20428 a_52635_34067.n43 a_52635_34067.t150 8.10567
R20429 a_52635_34067.n43 a_52635_34067.t134 8.10567
R20430 a_52635_34067.n47 a_52635_34067.t74 8.10567
R20431 a_52635_34067.n47 a_52635_34067.t156 8.10567
R20432 a_52635_34067.n21 a_52635_34067.t130 8.10567
R20433 a_52635_34067.n21 a_52635_34067.t135 8.10567
R20434 a_52635_34067.n21 a_52635_34067.t75 8.10567
R20435 a_52635_34067.n21 a_52635_34067.t157 8.10567
R20436 a_52635_34067.n157 a_52635_34067.t132 8.10567
R20437 a_52635_34067.n158 a_52635_34067.t219 8.10567
R20438 a_52635_34067.n20 a_52635_34067.t154 8.10567
R20439 a_52635_34067.n25 a_52635_34067.t236 8.10567
R20440 a_52635_34067.n25 a_52635_34067.t211 8.10567
R20441 a_52635_34067.n25 a_52635_34067.t126 8.10567
R20442 a_52635_34067.n4 a_52635_34067.t200 8.10567
R20443 a_52635_34067.n4 a_52635_34067.t153 8.10567
R20444 a_52635_34067.n4 a_52635_34067.t94 8.10567
R20445 a_52635_34067.n37 a_52635_34067.t147 8.10567
R20446 a_52635_34067.n151 a_52635_34067.t230 8.10567
R20447 a_52635_34067.n150 a_52635_34067.t220 8.10567
R20448 a_52635_34067.n38 a_52635_34067.t138 8.10567
R20449 a_52635_34067.n38 a_52635_34067.t124 8.10567
R20450 a_52635_34067.n39 a_52635_34067.t239 8.10567
R20451 a_52635_34067.n39 a_52635_34067.t142 8.10567
R20452 a_52635_34067.n33 a_52635_34067.t68 8.10567
R20453 a_52635_34067.n33 a_52635_34067.t71 8.10567
R20454 a_52635_34067.n33 a_52635_34067.t204 8.10567
R20455 a_52635_34067.n33 a_52635_34067.t96 8.10567
R20456 a_52635_34067.n162 a_52635_34067.t103 8.10567
R20457 a_52635_34067.n163 a_52635_34067.t190 8.10567
R20458 a_52635_34067.n31 a_52635_34067.t125 8.10567
R20459 a_52635_34067.n10 a_52635_34067.t184 8.10567
R20460 a_52635_34067.n10 a_52635_34067.t141 8.10567
R20461 a_52635_34067.n10 a_52635_34067.t67 8.10567
R20462 a_52635_34067.n30 a_52635_34067.t131 8.10567
R20463 a_52635_34067.n30 a_52635_34067.t91 8.10567
R20464 a_52635_34067.n30 a_52635_34067.t218 8.10567
R20465 a_52635_34067.n48 a_52635_34067.t119 8.10567
R20466 a_52635_34067.n161 a_52635_34067.t208 8.10567
R20467 a_52635_34067.n160 a_52635_34067.t192 8.10567
R20468 a_52635_34067.n45 a_52635_34067.t73 8.10567
R20469 a_52635_34067.n45 a_52635_34067.t237 8.10567
R20470 a_52635_34067.n49 a_52635_34067.t186 8.10567
R20471 a_52635_34067.n49 a_52635_34067.t82 8.10567
R20472 a_52635_34067.t12 a_52635_34067.n212 7.22198
R20473 a_52635_34067.t22 a_52635_34067.n195 7.22198
R20474 a_52635_34067.t57 a_52635_34067.t58 7.12006
R20475 a_52635_34067.n182 a_52635_34067.t5 6.77653
R20476 a_52635_34067.n142 a_52635_34067.t55 6.77653
R20477 a_52635_34067.n141 a_52635_34067.t44 6.7761
R20478 a_52635_34067.n205 a_52635_34067.t45 6.7761
R20479 a_52635_34067.n138 a_52635_34067.t61 6.86989
R20480 a_52635_34067.n127 a_52635_34067.t14 6.77231
R20481 a_52635_34067.n137 a_52635_34067.t23 6.77231
R20482 a_52635_34067.n188 a_52635_34067.t56 6.14835
R20483 a_52635_34067.n186 a_52635_34067.t64 6.14517
R20484 a_52635_34067.n140 a_52635_34067.t40 5.85898
R20485 a_52635_34067.t16 a_52635_34067.t13 5.70489
R20486 a_52635_34067.n195 a_52635_34067.t25 5.70489
R20487 a_52635_34067.t8 a_52635_34067.t34 5.70489
R20488 a_52635_34067.n212 a_52635_34067.t17 5.70489
R20489 a_52635_34067.n185 a_52635_34067.t63 5.61877
R20490 a_52635_34067.n143 a_52635_34067.t26 5.50607
R20491 a_52635_34067.n203 a_52635_34067.t48 5.50607
R20492 a_52635_34067.n183 a_52635_34067.t28 5.50607
R20493 a_52635_34067.n142 a_52635_34067.t43 5.50475
R20494 a_52635_34067.n141 a_52635_34067.t29 5.50475
R20495 a_52635_34067.n182 a_52635_34067.t6 5.50475
R20496 a_52635_34067.n199 a_52635_34067.t38 5.50475
R20497 a_52635_34067.n202 a_52635_34067.t42 5.50475
R20498 a_52635_34067.n205 a_52635_34067.t30 5.50475
R20499 a_52635_34067.n216 a_52635_34067.t37 5.50475
R20500 a_52635_34067.n139 a_52635_34067.t47 5.50475
R20501 a_52635_34067.n144 a_52635_34067.t50 5.50475
R20502 a_52635_34067.n204 a_52635_34067.t46 5.50475
R20503 a_52635_34067.n201 a_52635_34067.t10 5.50475
R20504 a_52635_34067.n200 a_52635_34067.t51 5.50475
R20505 a_52635_34067.n184 a_52635_34067.t54 5.50475
R20506 a_52635_34067.t0 a_52635_34067.n140 5.50475
R20507 a_52635_34067.n17 a_52635_34067.n16 0.595624
R20508 a_52635_34067.n85 a_52635_34067.n38 0.595624
R20509 a_52635_34067.n34 a_52635_34067.n43 0.607617
R20510 a_52635_34067.n46 a_52635_34067.n45 0.607617
R20511 a_52635_34067.n118 a_52635_34067.t32 5.5012
R20512 a_52635_34067.t52 a_52635_34067.n119 5.5012
R20513 a_52635_34067.t53 a_52635_34067.n120 5.5012
R20514 a_52635_34067.t1 a_52635_34067.n121 5.5012
R20515 a_52635_34067.t20 a_52635_34067.n122 5.5012
R20516 a_52635_34067.t2 a_52635_34067.n123 5.5012
R20517 a_52635_34067.t41 a_52635_34067.n124 5.5012
R20518 a_52635_34067.t7 a_52635_34067.n125 5.5012
R20519 a_52635_34067.t31 a_52635_34067.n126 5.5012
R20520 a_52635_34067.t15 a_52635_34067.n127 5.5012
R20521 a_52635_34067.n128 a_52635_34067.t36 5.5012
R20522 a_52635_34067.n129 a_52635_34067.t9 5.5012
R20523 a_52635_34067.n130 a_52635_34067.t11 5.5012
R20524 a_52635_34067.n131 a_52635_34067.t18 5.5012
R20525 a_52635_34067.n132 a_52635_34067.t27 5.5012
R20526 a_52635_34067.n133 a_52635_34067.t19 5.5012
R20527 a_52635_34067.n134 a_52635_34067.t4 5.5012
R20528 a_52635_34067.t21 a_52635_34067.n135 5.5012
R20529 a_52635_34067.t33 a_52635_34067.n136 5.5012
R20530 a_52635_34067.t24 a_52635_34067.n137 5.5012
R20531 a_52635_34067.t60 a_52635_34067.n138 5.66099
R20532 a_52635_34067.n107 a_52635_34067.n106 0.020246
R20533 a_52635_34067.n105 a_52635_34067.n104 0.020246
R20534 a_52635_34067.n74 a_52635_34067.n72 0.150783
R20535 a_52635_34067.n75 a_52635_34067.n71 0.150803
R20536 a_52635_34067.n116 a_52635_34067.n115 0.0676355
R20537 a_52635_34067.n82 a_52635_34067.n81 0.150803
R20538 a_52635_34067.n80 a_52635_34067.n79 0.150806
R20539 a_52635_34067.n113 a_52635_34067.n112 0.0676255
R20540 a_52635_34067.n60 a_52635_34067.n53 0.153625
R20541 a_52635_34067.n55 a_52635_34067.n54 0.153625
R20542 a_52635_34067.n93 a_52635_34067.n92 0.020088
R20543 a_52635_34067.n76 a_52635_34067.n75 0.246907
R20544 a_52635_34067.n74 a_52635_34067.n73 0.246877
R20545 a_52635_34067.n69 a_52635_34067.n68 0.153625
R20546 a_52635_34067.n65 a_52635_34067.n64 0.153625
R20547 a_52635_34067.n95 a_52635_34067.n94 0.020088
R20548 a_52635_34067.n111 a_52635_34067.n110 0.0201939
R20549 a_52635_34067.n68 a_52635_34067.n67 0.246907
R20550 a_52635_34067.n64 a_52635_34067.n63 0.246907
R20551 a_52635_34067.n79 a_52635_34067.n84 0.246907
R20552 a_52635_34067.n83 a_52635_34067.n82 0.246907
R20553 a_52635_34067.n109 a_52635_34067.n57 0.0201939
R20554 a_52635_34067.n61 a_52635_34067.n60 0.246907
R20555 a_52635_34067.n56 a_52635_34067.n55 0.246907
R20556 a_52635_34067.n27 a_52635_34067.n26 0.260442
R20557 a_52635_34067.n52 a_52635_34067.n47 0.591264
R20558 a_52635_34067.n36 a_52635_34067.n35 0.310971
R20559 a_52635_34067.n7 a_52635_34067.n6 0.258567
R20560 a_52635_34067.n4 a_52635_34067.n3 0.208479
R20561 a_52635_34067.n40 a_52635_34067.n39 0.591642
R20562 a_52635_34067.n22 a_52635_34067.n21 0.623337
R20563 a_52635_34067.n25 a_52635_34067.n24 0.259585
R20564 a_52635_34067.n30 a_52635_34067.n29 0.260442
R20565 a_52635_34067.n50 a_52635_34067.n49 0.591264
R20566 a_52635_34067.n33 a_52635_34067.n32 0.310971
R20567 a_52635_34067.n10 a_52635_34067.n9 0.258567
R20568 a_52635_34067.n1 a_52635_34067.n0 0.208479
R20569 a_52635_34067.n42 a_52635_34067.n15 0.591642
R20570 a_52635_34067.n19 a_52635_34067.n18 0.623337
R20571 a_52635_34067.n13 a_52635_34067.n12 0.259585
R20572 a_52635_34067.n191 a_52635_34067.n190 3.48654
R20573 a_52635_34067.n194 a_52635_34067.n190 3.42822
R20574 a_52635_34067.n147 a_52635_34067.n145 3.37173
R20575 a_52635_34067.t8 a_52635_34067.n211 3.23904
R20576 a_52635_34067.t16 a_52635_34067.n181 3.23904
R20577 a_52635_34067.n187 a_52635_34067.t57 3.23004
R20578 a_52635_34067.n201 a_52635_34067.n200 2.60203
R20579 a_52635_34067.n140 a_52635_34067.n139 2.60203
R20580 a_52635_34067.n184 a_52635_34067.n183 2.52436
R20581 a_52635_34067.n204 a_52635_34067.n203 2.52436
R20582 a_52635_34067.n144 a_52635_34067.n143 2.52436
R20583 a_52635_34067.n171 a_52635_34067.n170 2.40699
R20584 a_52635_34067.n159 a_52635_34067.n149 2.30989
R20585 a_52635_34067.n156 a_52635_34067.n44 2.30989
R20586 a_52635_34067.n187 a_52635_34067.n186 2.2807
R20587 a_52635_34067.n91 a_52635_34067.n90 0.427602
R20588 a_52635_34067.n59 a_52635_34067.n58 0.427602
R20589 a_52635_34067.n89 a_52635_34067.n88 0.427602
R20590 a_52635_34067.n87 a_52635_34067.n86 0.427602
R20591 a_52635_34067.n103 a_52635_34067.n102 0.420727
R20592 a_52635_34067.n101 a_52635_34067.n100 0.420727
R20593 a_52635_34067.n99 a_52635_34067.n98 0.420727
R20594 a_52635_34067.n97 a_52635_34067.n96 0.420727
R20595 a_52635_34067.n67 a_52635_34067.n66 2.96488
R20596 a_52635_34067.n62 a_52635_34067.n94 2.94096
R20597 a_52635_34067.n108 a_52635_34067.n61 2.96488
R20598 a_52635_34067.n93 a_52635_34067.n117 2.94096
R20599 a_52635_34067.n166 a_52635_34067.n114 2.07182
R20600 a_52635_34067.n167 a_52635_34067.n70 2.07182
R20601 a_52635_34067.n114 a_52635_34067.n71 2.75706
R20602 a_52635_34067.n106 a_52635_34067.n70 2.90773
R20603 a_52635_34067.n80 a_52635_34067.n78 2.75704
R20604 a_52635_34067.n77 a_52635_34067.n105 2.90773
R20605 a_52635_34067.n169 a_52635_34067.n147 1.80314
R20606 a_52635_34067.n180 a_52635_34067.n179 1.70908
R20607 a_52635_34067.n172 a_52635_34067.n171 1.68395
R20608 a_52635_34067.n179 a_52635_34067.n178 1.68395
R20609 a_52635_34067.n78 a_52635_34067.n165 1.5005
R20610 a_52635_34067.n66 a_52635_34067.n166 1.5005
R20611 a_52635_34067.n170 a_52635_34067.n108 1.5005
R20612 a_52635_34067.n117 a_52635_34067.n169 1.5005
R20613 a_52635_34067.n168 a_52635_34067.n77 1.5005
R20614 a_52635_34067.n167 a_52635_34067.n62 1.5005
R20615 a_52635_34067.n164 a_52635_34067.n28 1.5005
R20616 a_52635_34067.n159 a_52635_34067.n2 1.5005
R20617 a_52635_34067.n173 a_52635_34067.n172 1.5005
R20618 a_52635_34067.n178 a_52635_34067.n14 1.5005
R20619 a_52635_34067.n8 a_52635_34067.n148 1.5005
R20620 a_52635_34067.n23 a_52635_34067.n156 1.5005
R20621 a_52635_34067.n194 a_52635_34067.n193 1.5005
R20622 a_52635_34067.n196 a_52635_34067.t22 1.5005
R20623 a_52635_34067.n198 a_52635_34067.n197 1.5005
R20624 a_52635_34067.n208 a_52635_34067.n146 1.5005
R20625 a_52635_34067.n213 a_52635_34067.t12 1.5005
R20626 a_52635_34067.n189 a_52635_34067.n188 1.5005
R20627 a_52635_34067.n192 a_52635_34067.n191 1.5005
R20628 a_52635_34067.n207 a_52635_34067.n206 1.5005
R20629 a_52635_34067.n210 a_52635_34067.n209 1.5005
R20630 a_52635_34067.n180 a_52635_34067.t40 1.5005
R20631 a_52635_34067.n215 a_52635_34067.n214 1.5005
R20632 a_52635_34067.n166 a_52635_34067.n165 1.47516
R20633 a_52635_34067.n168 a_52635_34067.n167 1.47516
R20634 a_52635_34067.n190 a_52635_34067.n189 1.41182
R20635 a_52635_34067.n26 a_52635_34067.t166 9.17619
R20636 a_52635_34067.n29 a_52635_34067.t90 9.17619
R20637 a_52635_34067.n212 a_52635_34067.t8 1.27228
R20638 a_52635_34067.n200 a_52635_34067.n199 1.27228
R20639 a_52635_34067.n202 a_52635_34067.n201 1.27228
R20640 a_52635_34067.n195 a_52635_34067.t16 1.27228
R20641 a_52635_34067.n139 a_52635_34067.n216 1.27228
R20642 a_52635_34067.n183 a_52635_34067.n182 1.26756
R20643 a_52635_34067.n203 a_52635_34067.n202 1.26756
R20644 a_52635_34067.n143 a_52635_34067.n142 1.26756
R20645 a_52635_34067.n6 a_52635_34067.n5 1.24866
R20646 a_52635_34067.n47 a_52635_34067.n51 1.24866
R20647 a_52635_34067.n162 a_52635_34067.n10 1.24866
R20648 a_52635_34067.n49 a_52635_34067.n48 1.24866
R20649 a_52635_34067.n152 a_52635_34067.n27 1.24629
R20650 a_52635_34067.n160 a_52635_34067.n30 1.24629
R20651 a_52635_34067.n164 a_52635_34067.n159 1.23709
R20652 a_52635_34067.n156 a_52635_34067.n148 1.23709
R20653 a_52635_34067.n176 a_52635_34067.n19 1.22261
R20654 a_52635_34067.n174 a_52635_34067.n1 1.22261
R20655 a_52635_34067.n21 a_52635_34067.n20 1.22261
R20656 a_52635_34067.n150 a_52635_34067.n4 1.22261
R20657 a_52635_34067.n12 a_52635_34067.n11 1.21313
R20658 a_52635_34067.n42 a_52635_34067.n41 1.21313
R20659 a_52635_34067.n157 a_52635_34067.n25 1.21313
R20660 a_52635_34067.n39 a_52635_34067.n37 1.21313
R20661 a_52635_34067.n214 a_52635_34067.n145 1.10472
R20662 a_52635_34067.n172 a_52635_34067.n164 0.809892
R20663 a_52635_34067.n178 a_52635_34067.n148 0.809892
R20664 a_52635_34067.n198 a_52635_34067.n184 0.796291
R20665 a_52635_34067.n206 a_52635_34067.n204 0.796291
R20666 a_52635_34067.n215 a_52635_34067.n144 0.796291
R20667 a_52635_34067.n213 a_52635_34067.n146 0.780703
R20668 a_52635_34067.n196 a_52635_34067.n194 0.780703
R20669 a_52635_34067.n211 a_52635_34067.n210 0.780703
R20670 a_52635_34067.n191 a_52635_34067.n181 0.780703
R20671 a_52635_34067.n188 a_52635_34067.t59 0.769291
R20672 a_52635_34067.n186 a_52635_34067.n185 0.767125
R20673 a_52635_34067.n52 a_52635_34067.n149 1.14908
R20674 a_52635_34067.n44 a_52635_34067.n7 1.39299
R20675 a_52635_34067.n28 a_52635_34067.n50 1.14908
R20676 a_52635_34067.n9 a_52635_34067.n8 1.39299
R20677 a_52635_34067.n2 a_52635_34067.n40 1.11421
R20678 a_52635_34067.n24 a_52635_34067.n23 1.35707
R20679 a_52635_34067.n173 a_52635_34067.n15 1.11421
R20680 a_52635_34067.n14 a_52635_34067.n13 1.35707
R20681 a_52635_34067.n177 a_52635_34067.n176 0.673132
R20682 a_52635_34067.n11 a_52635_34067.n177 0.673132
R20683 a_52635_34067.n175 a_52635_34067.n174 0.673132
R20684 a_52635_34067.n41 a_52635_34067.n175 0.673132
R20685 a_52635_34067.n155 a_52635_34067.n154 0.673132
R20686 a_52635_34067.n5 a_52635_34067.n155 0.673132
R20687 a_52635_34067.n153 a_52635_34067.n152 0.673132
R20688 a_52635_34067.n51 a_52635_34067.n153 0.673132
R20689 a_52635_34067.n20 a_52635_34067.n158 0.673132
R20690 a_52635_34067.n158 a_52635_34067.n157 0.673132
R20691 a_52635_34067.n151 a_52635_34067.n150 0.673132
R20692 a_52635_34067.n37 a_52635_34067.n151 0.673132
R20693 a_52635_34067.n31 a_52635_34067.n163 0.673132
R20694 a_52635_34067.n163 a_52635_34067.n162 0.673132
R20695 a_52635_34067.n161 a_52635_34067.n160 0.673132
R20696 a_52635_34067.n48 a_52635_34067.n161 0.673132
R20697 a_52635_34067.n214 a_52635_34067.n213 0.638405
R20698 a_52635_34067.n197 a_52635_34067.n196 0.638405
R20699 a_52635_34067.n189 a_52635_34067.n187 0.638405
R20700 a_52635_34067.n211 a_52635_34067.n180 0.638405
R20701 a_52635_34067.n207 a_52635_34067.n181 0.638405
R20702 a_52635_34067.n197 a_52635_34067.n146 0.628372
R20703 a_52635_34067.n210 a_52635_34067.n207 0.628372
R20704 a_52635_34067.n179 a_52635_34067.n147 0.604355
R20705 a_52635_34067.n171 a_52635_34067.n145 0.603852
R20706 a_52635_34067.n170 a_52635_34067.n165 0.571818
R20707 a_52635_34067.n169 a_52635_34067.n168 0.571818
R20708 a_52635_34067.n199 a_52635_34067.n198 0.476484
R20709 a_52635_34067.n206 a_52635_34067.n205 0.476484
R20710 a_52635_34067.n216 a_52635_34067.n215 0.476484
R20711 a_52635_34067.t40 a_52635_34067.n141 0.476484
R20712 a_52635_34067.n52 a_52635_34067.n34 1.14166
R20713 a_52635_34067.n44 a_52635_34067.n35 2.75347
R20714 a_52635_34067.n46 a_52635_34067.n50 1.14166
R20715 a_52635_34067.n8 a_52635_34067.n32 2.75347
R20716 a_52635_34067.n124 a_52635_34067.n208 0.478684
R20717 a_52635_34067.n209 a_52635_34067.n118 0.478684
R20718 a_52635_34067.n193 a_52635_34067.n134 0.478684
R20719 a_52635_34067.n192 a_52635_34067.n128 0.478684
R20720 a_52635_34067.n59 a_52635_34067.n57 2.03311
R20721 a_52635_34067.n53 a_52635_34067.n59 2.04491
R20722 a_52635_34067.n54 a_52635_34067.n53 4.37762
R20723 a_52635_34067.n91 a_52635_34067.n54 1.87961
R20724 a_52635_34067.n91 a_52635_34067.n93 2.19836
R20725 a_52635_34067.n101 a_52635_34067.n115 2.03667
R20726 a_52635_34067.n76 a_52635_34067.n101 2.2172
R20727 a_52635_34067.n76 a_52635_34067.n73 4.49278
R20728 a_52635_34067.n103 a_52635_34067.n73 1.82125
R20729 a_52635_34067.n103 a_52635_34067.n106 2.19319
R20730 a_52635_34067.n115 a_52635_34067.n114 1.65342
R20731 a_52635_34067.n72 a_52635_34067.n71 4.34534
R20732 a_52635_34067.n72 a_52635_34067.n70 1.50598
R20733 a_52635_34067.n87 a_52635_34067.n110 2.03311
R20734 a_52635_34067.n69 a_52635_34067.n87 2.04491
R20735 a_52635_34067.n65 a_52635_34067.n69 4.37762
R20736 a_52635_34067.n89 a_52635_34067.n65 1.87961
R20737 a_52635_34067.n94 a_52635_34067.n89 2.19836
R20738 a_52635_34067.n66 a_52635_34067.n110 1.65903
R20739 a_52635_34067.n67 a_52635_34067.n63 4.49309
R20740 a_52635_34067.n63 a_52635_34067.n62 1.44546
R20741 a_52635_34067.n97 a_52635_34067.n113 2.03657
R20742 a_52635_34067.n97 a_52635_34067.n84 2.21715
R20743 a_52635_34067.n83 a_52635_34067.n84 4.49317
R20744 a_52635_34067.n99 a_52635_34067.n83 1.82113
R20745 a_52635_34067.n105 a_52635_34067.n99 2.19319
R20746 a_52635_34067.n78 a_52635_34067.n113 1.65366
R20747 a_52635_34067.n81 a_52635_34067.n80 4.34574
R20748 a_52635_34067.n81 a_52635_34067.n77 1.50586
R20749 a_52635_34067.n57 a_52635_34067.n108 1.65903
R20750 a_52635_34067.n61 a_52635_34067.n56 4.49309
R20751 a_52635_34067.n56 a_52635_34067.n117 1.44546
R20752 a_52635_34067.n149 a_52635_34067.n26 2.8103
R20753 a_52635_34067.n35 a_52635_34067.n34 4.38327
R20754 a_52635_34067.n3 a_52635_34067.n2 2.83621
R20755 a_52635_34067.n40 a_52635_34067.n85 1.15119
R20756 a_52635_34067.n85 a_52635_34067.n22 4.37089
R20757 a_52635_34067.n22 a_52635_34067.n23 2.6764
R20758 a_52635_34067.n29 a_52635_34067.n28 2.8103
R20759 a_52635_34067.n46 a_52635_34067.n32 4.38327
R20760 a_52635_34067.n173 a_52635_34067.n0 2.83621
R20761 a_52635_34067.n17 a_52635_34067.n15 1.15119
R20762 a_52635_34067.n18 a_52635_34067.n17 4.37089
R20763 a_52635_34067.n18 a_52635_34067.n14 2.6764
R20764 a_52635_34067.n126 a_52635_34067.n127 1.27228
R20765 a_52635_34067.n125 a_52635_34067.n126 2.51878
R20766 a_52635_34067.n208 a_52635_34067.n125 0.794091
R20767 a_52635_34067.n123 a_52635_34067.n124 1.27228
R20768 a_52635_34067.n122 a_52635_34067.n123 2.60203
R20769 a_52635_34067.n121 a_52635_34067.n122 1.27228
R20770 a_52635_34067.n120 a_52635_34067.n121 1.27228
R20771 a_52635_34067.n119 a_52635_34067.n120 2.51878
R20772 a_52635_34067.n209 a_52635_34067.n119 0.794091
R20773 a_52635_34067.t49 a_52635_34067.n118 6.77266
R20774 a_52635_34067.n136 a_52635_34067.n137 1.27228
R20775 a_52635_34067.n135 a_52635_34067.n136 2.51878
R20776 a_52635_34067.n193 a_52635_34067.n135 0.794091
R20777 a_52635_34067.n133 a_52635_34067.n134 1.27228
R20778 a_52635_34067.n132 a_52635_34067.n133 2.60203
R20779 a_52635_34067.n131 a_52635_34067.n132 1.27228
R20780 a_52635_34067.n130 a_52635_34067.n131 1.27228
R20781 a_52635_34067.n129 a_52635_34067.n130 2.51878
R20782 a_52635_34067.n192 a_52635_34067.n129 0.794091
R20783 a_52635_34067.t3 a_52635_34067.n128 6.77266
R20784 a_52635_34067.n185 a_52635_34067.n138 3.17898
R20785 a_52635_34067.n16 a_52635_34067.n42 2.16997
R20786 a_52635_34067.n39 a_52635_34067.n38 2.16997
R20787 a_52635_34067.n154 a_52635_34067.n36 2.13563
R20788 a_52635_34067.n33 a_52635_34067.n31 2.13563
R20789 a_52635_34067.n43 a_52635_34067.n47 2.13445
R20790 a_52635_34067.n49 a_52635_34067.n45 2.13445
R20791 a_52635_34067.t152 a_52635_34067.n3 9.16748
R20792 a_52635_34067.t212 a_52635_34067.n0 9.16748
R20793 VDD.n7996 VDD.n2188 714.056
R20794 VDD.n7994 VDD.n2188 712.232
R20795 VDD.n7996 VDD.n2187 707.59
R20796 VDD.n7994 VDD.n2187 705.766
R20797 VDD.n1743 VDD.n686 694.492
R20798 VDD.n1717 VDD.n710 694.492
R20799 VDD.n1351 VDD.n1350 694.492
R20800 VDD.n1427 VDD.n850 694.492
R20801 VDD.n1416 VDD.n845 694.492
R20802 VDD.n1720 VDD.n707 694.492
R20803 VDD.n1653 VDD.n758 694.492
R20804 VDD.n1344 VDD.n1343 694.492
R20805 VDD.n1357 VDD.n848 694.492
R20806 VDD.n1413 VDD.n875 694.492
R20807 VDD.n762 VDD.n760 694.492
R20808 VDD.n1741 VDD.n691 694.492
R20809 VDD.n688 VDD.n686 694.078
R20810 VDD.n711 VDD.n710 694.078
R20811 VDD.n1351 VDD.n1276 694.078
R20812 VDD.n1427 VDD.n849 694.078
R20813 VDD.n1416 VDD.n846 694.078
R20814 VDD.n1720 VDD.n708 694.078
R20815 VDD.n761 VDD.n758 694.078
R20816 VDD.n1348 VDD.n1344 694.078
R20817 VDD.n1355 VDD.n848 694.078
R20818 VDD.n1390 VDD.n875 694.078
R20819 VDD.n1651 VDD.n762 694.078
R20820 VDD.n691 VDD.n689 694.078
R20821 VDD.n1743 VDD.n687 692.172
R20822 VDD.n1717 VDD.n712 692.172
R20823 VDD.n1350 VDD.n1277 692.172
R20824 VDD.n1353 VDD.n850 692.172
R20825 VDD.n1430 VDD.n845 692.172
R20826 VDD.n859 VDD.n707 692.172
R20827 VDD.n1653 VDD.n759 692.172
R20828 VDD.n1347 VDD.n1343 692.172
R20829 VDD.n1357 VDD.n1083 692.172
R20830 VDD.n1413 VDD.n847 692.172
R20831 VDD.n764 VDD.n760 692.172
R20832 VDD.n1741 VDD.n692 692.172
R20833 VDD.n688 VDD.n687 691.758
R20834 VDD.n712 VDD.n711 691.758
R20835 VDD.n1277 VDD.n1276 691.758
R20836 VDD.n1353 VDD.n849 691.758
R20837 VDD.n1430 VDD.n846 691.758
R20838 VDD.n859 VDD.n708 691.758
R20839 VDD.n761 VDD.n759 691.758
R20840 VDD.n1348 VDD.n1347 691.758
R20841 VDD.n1355 VDD.n1083 691.758
R20842 VDD.n1390 VDD.n847 691.758
R20843 VDD.n1651 VDD.n764 691.758
R20844 VDD.n692 VDD.n689 691.758
R20845 VDD.n2331 VDD.n2235 647.574
R20846 VDD.n2351 VDD.n2321 647.574
R20847 VDD.n5276 VDD.n5221 647.574
R20848 VDD.n5305 VDD.n5304 647.574
R20849 VDD.n7042 VDD.n7041 647.574
R20850 VDD.n5277 VDD.n5264 647.574
R20851 VDD.n5312 VDD.n5306 647.574
R20852 VDD.n2332 VDD.n2236 647.574
R20853 VDD.n2367 VDD.n2352 647.574
R20854 VDD.n5278 VDD.n5266 647.574
R20855 VDD.n5378 VDD.n5307 647.574
R20856 VDD.n7835 VDD.n2234 647.574
R20857 VDD.n2353 VDD.n2312 647.574
R20858 VDD.n6578 VDD.n5270 647.574
R20859 VDD.n5942 VDD.n5308 647.574
R20860 VDD.n7833 VDD.n2238 647.574
R20861 VDD.n2331 VDD.n2318 642.269
R20862 VDD.n2369 VDD.n2351 642.269
R20863 VDD.n5282 VDD.n5276 642.269
R20864 VDD.n5305 VDD.n5303 642.269
R20865 VDD.n7041 VDD.n2349 642.269
R20866 VDD.n6371 VDD.n5277 642.269
R20867 VDD.n5311 VDD.n5306 642.269
R20868 VDD.n2332 VDD.n2319 642.269
R20869 VDD.n6634 VDD.n2352 642.269
R20870 VDD.n6369 VDD.n5278 642.269
R20871 VDD.n6310 VDD.n5307 642.269
R20872 VDD.n7134 VDD.n2234 642.269
R20873 VDD.n6632 VDD.n2353 642.269
R20874 VDD.n6578 VDD.n5275 642.269
R20875 VDD.n6312 VDD.n5308 642.269
R20876 VDD.n7132 VDD.n2238 642.269
R20877 VDD.n7087 VDD.n2235 640.197
R20878 VDD.n7039 VDD.n2321 640.197
R20879 VDD.n6576 VDD.n5221 640.197
R20880 VDD.n6397 VDD.n5304 640.197
R20881 VDD.n7042 VDD.n2348 640.197
R20882 VDD.n5281 VDD.n5264 640.197
R20883 VDD.n6395 VDD.n5312 640.197
R20884 VDD.n7085 VDD.n2236 640.197
R20885 VDD.n2368 VDD.n2367 640.197
R20886 VDD.n5280 VDD.n5266 640.197
R20887 VDD.n5378 VDD.n5310 640.197
R20888 VDD.n7835 VDD.n2210 640.197
R20889 VDD.n2357 VDD.n2312 640.197
R20890 VDD.n5279 VDD.n5270 640.197
R20891 VDD.n5942 VDD.n5309 640.197
R20892 VDD.n7833 VDD.n2237 640.197
R20893 VDD.n7087 VDD.n2318 634.891
R20894 VDD.n7039 VDD.n2369 634.891
R20895 VDD.n6576 VDD.n5282 634.891
R20896 VDD.n6397 VDD.n5303 634.891
R20897 VDD.n2349 VDD.n2348 634.891
R20898 VDD.n6371 VDD.n5281 634.891
R20899 VDD.n6395 VDD.n5311 634.891
R20900 VDD.n7085 VDD.n2319 634.891
R20901 VDD.n6634 VDD.n2368 634.891
R20902 VDD.n6369 VDD.n5280 634.891
R20903 VDD.n6310 VDD.n5310 634.891
R20904 VDD.n7134 VDD.n2210 634.891
R20905 VDD.n6632 VDD.n2357 634.891
R20906 VDD.n5279 VDD.n5275 634.891
R20907 VDD.n6312 VDD.n5309 634.891
R20908 VDD.n7132 VDD.n2237 634.891
R20909 VDD.n1550 VDD.n1521 614.001
R20910 VDD.n1550 VDD.n1549 613.338
R20911 VDD.n1552 VDD.n1521 607.537
R20912 VDD.n1552 VDD.n1549 606.872
R20913 VDD.n12614 VDD.n13 477.971
R20914 VDD.n12610 VDD.n16 477.971
R20915 VDD.n12529 VDD.n31 477.971
R20916 VDD.n12522 VDD.n43 477.971
R20917 VDD.n12516 VDD.n96 477.971
R20918 VDD.n12473 VDD.n111 477.971
R20919 VDD.n11027 VDD.n1771 477.971
R20920 VDD.n11006 VDD.n1785 477.971
R20921 VDD.n10999 VDD.n10998 477.971
R20922 VDD.n10994 VDD.n1833 477.971
R20923 VDD.n10951 VDD.n1848 477.971
R20924 VDD.n10944 VDD.n10943 477.971
R20925 VDD.n10939 VDD.n1898 477.971
R20926 VDD.n10896 VDD.n1913 477.971
R20927 VDD.n10889 VDD.n10888 477.971
R20928 VDD.n10884 VDD.n1925 477.971
R20929 VDD.n10841 VDD.n1940 477.971
R20930 VDD.n10834 VDD.n10833 477.971
R20931 VDD.n10829 VDD.n1990 477.971
R20932 VDD.n10783 VDD.n2013 477.971
R20933 VDD.n10776 VDD.n10775 477.971
R20934 VDD.n9157 VDD.n8473 477.971
R20935 VDD.n9033 VDD.n8491 477.971
R20936 VDD.n9014 VDD.n8500 477.971
R20937 VDD.n8936 VDD.n8508 477.971
R20938 VDD.n8883 VDD.n8519 477.971
R20939 VDD.n8805 VDD.n8527 477.971
R20940 VDD.n12460 VDD.n176 477.971
R20941 VDD.n12466 VDD.n123 477.971
R20942 VDD.n9178 VDD.n8460 477.971
R20943 VDD.n12592 VDD.n14 470.842
R20944 VDD.n30 VDD.n17 470.842
R20945 VDD.n12524 VDD.n32 470.842
R20946 VDD.n12521 VDD.n44 470.842
R20947 VDD.n110 VDD.n97 470.842
R20948 VDD.n12468 VDD.n112 470.842
R20949 VDD.n11030 VDD.n1772 470.842
R20950 VDD.n11001 VDD.n1784 470.842
R20951 VDD.n1795 VDD.n1794 470.842
R20952 VDD.n1846 VDD.n1832 470.842
R20953 VDD.n10946 VDD.n1847 470.842
R20954 VDD.n1860 VDD.n1859 470.842
R20955 VDD.n1911 VDD.n1897 470.842
R20956 VDD.n10891 VDD.n1912 470.842
R20957 VDD.n1921 VDD.n1920 470.842
R20958 VDD.n1938 VDD.n1924 470.842
R20959 VDD.n10836 VDD.n1939 470.842
R20960 VDD.n1952 VDD.n1951 470.842
R20961 VDD.n2011 VDD.n1989 470.842
R20962 VDD.n10778 VDD.n2012 470.842
R20963 VDD.n2025 VDD.n2024 470.842
R20964 VDD.n9160 VDD.n8466 470.842
R20965 VDD.n9036 VDD.n8480 470.842
R20966 VDD.n9009 VDD.n8501 470.842
R20967 VDD.n8939 VDD.n8509 470.842
R20968 VDD.n8878 VDD.n8520 470.842
R20969 VDD.n8808 VDD.n8528 470.842
R20970 VDD.n8539 VDD.n177 470.842
R20971 VDD.n12465 VDD.n124 470.842
R20972 VDD.n9182 VDD.n8461 470.842
R20973 VDD.n12614 VDD.n14 470.842
R20974 VDD.n30 VDD.n16 470.842
R20975 VDD.n12524 VDD.n31 470.842
R20976 VDD.n44 VDD.n43 470.842
R20977 VDD.n110 VDD.n96 470.842
R20978 VDD.n12468 VDD.n111 470.842
R20979 VDD.n11027 VDD.n1772 470.842
R20980 VDD.n11001 VDD.n1785 470.842
R20981 VDD.n10998 VDD.n1795 470.842
R20982 VDD.n1846 VDD.n1833 470.842
R20983 VDD.n10946 VDD.n1848 470.842
R20984 VDD.n10943 VDD.n1860 470.842
R20985 VDD.n1911 VDD.n1898 470.842
R20986 VDD.n10891 VDD.n1913 470.842
R20987 VDD.n10888 VDD.n1921 470.842
R20988 VDD.n1938 VDD.n1925 470.842
R20989 VDD.n10836 VDD.n1940 470.842
R20990 VDD.n10833 VDD.n1952 470.842
R20991 VDD.n2011 VDD.n1990 470.842
R20992 VDD.n10778 VDD.n2013 470.842
R20993 VDD.n10775 VDD.n2025 470.842
R20994 VDD.n9157 VDD.n8466 470.842
R20995 VDD.n9033 VDD.n8480 470.842
R20996 VDD.n9014 VDD.n8501 470.842
R20997 VDD.n8936 VDD.n8509 470.842
R20998 VDD.n8883 VDD.n8520 470.842
R20999 VDD.n8805 VDD.n8528 470.842
R21000 VDD.n8539 VDD.n176 470.842
R21001 VDD.n124 VDD.n123 470.842
R21002 VDD.n9182 VDD.n8460 470.842
R21003 VDD.n12592 VDD.n13 469.683
R21004 VDD.n12610 VDD.n17 469.683
R21005 VDD.n12529 VDD.n32 469.683
R21006 VDD.n12522 VDD.n12521 469.683
R21007 VDD.n12516 VDD.n97 469.683
R21008 VDD.n12473 VDD.n112 469.683
R21009 VDD.n11030 VDD.n1771 469.683
R21010 VDD.n11006 VDD.n1784 469.683
R21011 VDD.n10999 VDD.n1794 469.683
R21012 VDD.n10994 VDD.n1832 469.683
R21013 VDD.n10951 VDD.n1847 469.683
R21014 VDD.n10944 VDD.n1859 469.683
R21015 VDD.n10939 VDD.n1897 469.683
R21016 VDD.n10896 VDD.n1912 469.683
R21017 VDD.n10889 VDD.n1920 469.683
R21018 VDD.n10884 VDD.n1924 469.683
R21019 VDD.n10841 VDD.n1939 469.683
R21020 VDD.n10834 VDD.n1951 469.683
R21021 VDD.n10829 VDD.n1989 469.683
R21022 VDD.n10783 VDD.n2012 469.683
R21023 VDD.n10776 VDD.n2024 469.683
R21024 VDD.n9160 VDD.n8473 469.683
R21025 VDD.n9036 VDD.n8491 469.683
R21026 VDD.n9009 VDD.n8500 469.683
R21027 VDD.n8939 VDD.n8508 469.683
R21028 VDD.n8878 VDD.n8519 469.683
R21029 VDD.n8808 VDD.n8527 469.683
R21030 VDD.n12460 VDD.n177 469.683
R21031 VDD.n12466 VDD.n12465 469.683
R21032 VDD.n9178 VDD.n8461 469.683
R21033 VDD.n8078 VDD.n2123 351.805
R21034 VDD.n8078 VDD.n2124 351.639
R21035 VDD.n8076 VDD.n2123 350.479
R21036 VDD.n8076 VDD.n2124 350.313
R21037 VDD.t1665 VDD.t920 338.731
R21038 VDD.t994 VDD.t2299 338.731
R21039 VDD.t692 VDD.t1665 260.622
R21040 VDD.t1188 VDD.t994 260.622
R21041 VDD.t920 VDD.n1521 167.008
R21042 VDD.t2299 VDD.n1549 167.008
R21043 VDD.n1551 VDD.t692 156.792
R21044 VDD.n1551 VDD.t1188 155.268
R21045 VDD.t338 VDD.t1099 142.93
R21046 VDD.t1419 VDD.t337 142.93
R21047 VDD.t1747 VDD.t521 142.93
R21048 VDD.t522 VDD.t2231 142.93
R21049 VDD.t322 VDD.t2485 142.93
R21050 VDD.t321 VDD.t944 142.93
R21051 VDD.t500 VDD.t917 142.93
R21052 VDD.t2777 VDD.t497 142.93
R21053 VDD.t893 VDD.t553 142.93
R21054 VDD.t552 VDD.t697 142.93
R21055 VDD.t643 VDD.t801 142.93
R21056 VDD.t2774 VDD.t1049 142.93
R21057 VDD.t1841 VDD.t2118 142.93
R21058 VDD.t1183 VDD.t2924 142.93
R21059 VDD.t1365 VDD.t352 142.93
R21060 VDD.t351 VDD.t1799 142.93
R21061 VDD.t1378 VDD.t875 142.93
R21062 VDD.t2261 VDD.t1262 142.93
R21063 VDD.t1512 VDD.t638 142.93
R21064 VDD.t2573 VDD.t2542 142.93
R21065 VDD.t955 VDD.t3747 142.93
R21066 VDD.t3678 VDD.t1370 142.93
R21067 VDD.t496 VDD.t1549 142.93
R21068 VDD.t507 VDD.t648 142.93
R21069 VDD.t287 VDD.t1714 142.93
R21070 VDD.t1206 VDD.t288 142.93
R21071 VDD.t1177 VDD.t1494 142.93
R21072 VDD.t3423 VDD.t677 142.93
R21073 VDD.t305 VDD.t2349 142.93
R21074 VDD.t302 VDD.t1349 142.93
R21075 VDD.t538 VDD.t1481 142.93
R21076 VDD.t535 VDD.t1086 142.93
R21077 VDD.t1290 VDD.t1570 142.93
R21078 VDD.t1155 VDD.t1904 142.93
R21079 VDD.t1515 VDD.t532 142.93
R21080 VDD.t523 VDD.t1611 142.93
R21081 VDD.t1996 VDD.t625 142.93
R21082 VDD.t795 VDD.t748 142.93
R21083 VDD.t550 VDD.t1653 142.93
R21084 VDD.t828 VDD.t548 142.93
R21085 VDD.t725 VDD.t1486 142.93
R21086 VDD.t2729 VDD.t1821 142.93
R21087 VDD.t501 VDD.t1787 142.93
R21088 VDD.t2344 VDD.t610 142.93
R21089 VDD.t2058 VDD.t792 142.93
R21090 VDD.t1408 VDD.t2251 142.93
R21091 VDD.t898 VDD.t1 142.93
R21092 VDD.t0 VDD.t1489 142.93
R21093 VDD.t2464 VDD.t546 142.93
R21094 VDD.t543 VDD.t2099 142.93
R21095 VDD.t630 VDD.t297 142.93
R21096 VDD.t417 VDD.t667 142.93
R21097 VDD.t842 VDD.t2325 142.93
R21098 VDD.t2559 VDD.t836 142.93
R21099 VDD.t2079 VDD.t1796 142.93
R21100 VDD.t560 VDD.t2160 142.93
R21101 VDD.t2155 VDD.t1893 142.93
R21102 VDD.t680 VDD.t2254 142.93
R21103 VDD.t551 VDD.t2142 142.93
R21104 VDD.t2399 VDD.t622 142.93
R21105 VDD.t1099 VDD.t965 96.8792
R21106 VDD.t335 VDD.t338 96.8792
R21107 VDD.t337 VDD.t336 96.8792
R21108 VDD.t1642 VDD.t1419 96.8792
R21109 VDD.t1354 VDD.t1747 96.8792
R21110 VDD.t521 VDD.t520 96.8792
R21111 VDD.t519 VDD.t522 96.8792
R21112 VDD.t2231 VDD.t1112 96.8792
R21113 VDD.t2485 VDD.t852 96.8792
R21114 VDD.t298 VDD.t322 96.8792
R21115 VDD.t293 VDD.t321 96.8792
R21116 VDD.t944 VDD.t745 96.8792
R21117 VDD.t917 VDD.t789 96.8792
R21118 VDD.t499 VDD.t500 96.8792
R21119 VDD.t497 VDD.t498 96.8792
R21120 VDD.t1142 VDD.t2777 96.8792
R21121 VDD.t935 VDD.t893 96.8792
R21122 VDD.t553 VDD.t555 96.8792
R21123 VDD.t554 VDD.t552 96.8792
R21124 VDD.t697 VDD.t780 96.8792
R21125 VDD.t801 VDD.t1658 96.8792
R21126 VDD.t1442 VDD.t643 96.8792
R21127 VDD.t3354 VDD.t2774 96.8792
R21128 VDD.t1049 VDD.t2680 96.8792
R21129 VDD.t2118 VDD.t855 96.8792
R21130 VDD.t571 VDD.t1841 96.8792
R21131 VDD.t2924 VDD.t3570 96.8792
R21132 VDD.t905 VDD.t1183 96.8792
R21133 VDD.t2570 VDD.t1365 96.8792
R21134 VDD.t352 VDD.t363 96.8792
R21135 VDD.t353 VDD.t351 96.8792
R21136 VDD.t1799 VDD.t1957 96.8792
R21137 VDD.t875 VDD.t1936 96.8792
R21138 VDD.t866 VDD.t1378 96.8792
R21139 VDD.t1338 VDD.t2261 96.8792
R21140 VDD.t1262 VDD.t1209 96.8792
R21141 VDD.t638 VDD.t798 96.8792
R21142 VDD.t3013 VDD.t1512 96.8792
R21143 VDD.t2542 VDD.t664 96.8792
R21144 VDD.t1373 VDD.t2573 96.8792
R21145 VDD.t813 VDD.t955 96.8792
R21146 VDD.t3747 VDD.t2921 96.8792
R21147 VDD.t1405 VDD.t3678 96.8792
R21148 VDD.t1370 VDD.t1180 96.8792
R21149 VDD.t1549 VDD.t674 96.8792
R21150 VDD.t508 VDD.t496 96.8792
R21151 VDD.t510 VDD.t507 96.8792
R21152 VDD.t648 VDD.t1439 96.8792
R21153 VDD.t1714 VDD.t1164 96.8792
R21154 VDD.t290 VDD.t287 96.8792
R21155 VDD.t288 VDD.t289 96.8792
R21156 VDD.t1081 VDD.t1206 96.8792
R21157 VDD.t1322 VDD.t1177 96.8792
R21158 VDD.t1494 VDD.t1711 96.8792
R21159 VDD.t3613 VDD.t3423 96.8792
R21160 VDD.t677 VDD.t930 96.8792
R21161 VDD.t2349 VDD.t598 96.8792
R21162 VDD.t303 VDD.t305 96.8792
R21163 VDD.t326 VDD.t302 96.8792
R21164 VDD.t1349 VDD.t755 96.8792
R21165 VDD.t1481 VDD.t833 96.8792
R21166 VDD.t536 VDD.t538 96.8792
R21167 VDD.t537 VDD.t535 96.8792
R21168 VDD.t1086 VDD.t1780 96.8792
R21169 VDD.t1570 VDD.t1218 96.8792
R21170 VDD.t1540 VDD.t1290 96.8792
R21171 VDD.t1904 VDD.t845 96.8792
R21172 VDD.t1884 VDD.t1155 96.8792
R21173 VDD.t1299 VDD.t1515 96.8792
R21174 VDD.t532 VDD.t524 96.8792
R21175 VDD.t529 VDD.t523 96.8792
R21176 VDD.t1611 VDD.t686 96.8792
R21177 VDD.t625 VDD.t635 96.8792
R21178 VDD.t2240 VDD.t1996 96.8792
R21179 VDD.t2422 VDD.t795 96.8792
R21180 VDD.t748 VDD.t976 96.8792
R21181 VDD.t1653 VDD.t1424 96.8792
R21182 VDD.t549 VDD.t550 96.8792
R21183 VDD.t548 VDD.t547 96.8792
R21184 VDD.t619 VDD.t828 96.8792
R21185 VDD.t1505 VDD.t725 96.8792
R21186 VDD.t1486 VDD.t1708 96.8792
R21187 VDD.t1850 VDD.t2729 96.8792
R21188 VDD.t1821 VDD.t2076 96.8792
R21189 VDD.t1787 VDD.t1052 96.8792
R21190 VDD.t2382 VDD.t501 96.8792
R21191 VDD.t502 VDD.t2344 96.8792
R21192 VDD.t610 VDD.t823 96.8792
R21193 VDD.t792 VDD.t1127 96.8792
R21194 VDD.t2812 VDD.t2058 96.8792
R21195 VDD.t2251 VDD.t2021 96.8792
R21196 VDD.t810 VDD.t1408 96.8792
R21197 VDD.t1195 VDD.t898 96.8792
R21198 VDD.t1 VDD.t6 96.8792
R21199 VDD.t2 VDD.t0 96.8792
R21200 VDD.t1489 VDD.t1333 96.8792
R21201 VDD.t1265 VDD.t2464 96.8792
R21202 VDD.t546 VDD.t544 96.8792
R21203 VDD.t545 VDD.t543 96.8792
R21204 VDD.t2099 VDD.t1015 96.8792
R21205 VDD.t1818 VDD.t630 96.8792
R21206 VDD.t297 VDD.t367 96.8792
R21207 VDD.t301 VDD.t417 96.8792
R21208 VDD.t667 VDD.t979 96.8792
R21209 VDD.t1251 VDD.t842 96.8792
R21210 VDD.t2325 VDD.t707 96.8792
R21211 VDD.t2288 VDD.t2559 96.8792
R21212 VDD.t836 VDD.t1042 96.8792
R21213 VDD.t1824 VDD.t2079 96.8792
R21214 VDD.t1796 VDD.t2061 96.8792
R21215 VDD.t2189 VDD.t560 96.8792
R21216 VDD.t2160 VDD.t2447 96.8792
R21217 VDD.t1917 VDD.t2155 96.8792
R21218 VDD.t1893 VDD.t2127 96.8792
R21219 VDD.t2302 VDD.t680 96.8792
R21220 VDD.t2254 VDD.t603 96.8792
R21221 VDD.t2142 VDD.t1867 96.8792
R21222 VDD.t2088 VDD.t551 96.8792
R21223 VDD.t622 VDD.t2228 96.8792
R21224 VDD.t720 VDD.t2399 96.8792
R21225 VDD.t568 VDD.t405 85.1494
R21226 VDD.t12 VDD.t910 85.1494
R21227 VDD.t34 VDD.t925 85.1494
R21228 VDD.t390 VDD.t962 81.7244
R21229 VDD.t965 VDD.n1771 81.1238
R21230 VDD.t755 VDD.n2025 81.1238
R21231 VDD.t833 VDD.n13 81.1238
R21232 VDD.n9182 VDD.t720 81.1238
R21233 VDD.n1786 VDD.t1642 81.017
R21234 VDD.n11005 VDD.t1354 81.017
R21235 VDD.t1112 VDD.n11002 81.017
R21236 VDD.t852 VDD.n1787 81.017
R21237 VDD.t745 VDD.n10996 81.017
R21238 VDD.n10995 VDD.t789 81.017
R21239 VDD.n1851 VDD.t1142 81.017
R21240 VDD.n10950 VDD.t935 81.017
R21241 VDD.t780 VDD.n10947 81.017
R21242 VDD.t1658 VDD.n1852 81.017
R21243 VDD.t2680 VDD.n10941 81.017
R21244 VDD.n10940 VDD.t855 81.017
R21245 VDD.n1916 VDD.t905 81.017
R21246 VDD.n10895 VDD.t2570 81.017
R21247 VDD.t1957 VDD.n10892 81.017
R21248 VDD.t1936 VDD.n1917 81.017
R21249 VDD.t1209 VDD.n10886 81.017
R21250 VDD.n10885 VDD.t798 81.017
R21251 VDD.n1943 VDD.t1373 81.017
R21252 VDD.n10840 VDD.t813 81.017
R21253 VDD.t1180 VDD.n10837 81.017
R21254 VDD.t674 VDD.n1944 81.017
R21255 VDD.t1439 VDD.n10831 81.017
R21256 VDD.n10830 VDD.t1164 81.017
R21257 VDD.n2016 VDD.t1081 81.017
R21258 VDD.n10782 VDD.t1322 81.017
R21259 VDD.t930 VDD.n10779 81.017
R21260 VDD.t598 VDD.n2017 81.017
R21261 VDD.t1780 VDD.n12612 81.017
R21262 VDD.n12611 VDD.t1218 81.017
R21263 VDD.n35 VDD.t1884 81.017
R21264 VDD.n12528 VDD.t1299 81.017
R21265 VDD.t686 VDD.n12525 81.017
R21266 VDD.t635 VDD.n36 81.017
R21267 VDD.t976 VDD.n12518 81.017
R21268 VDD.n12517 VDD.t1424 81.017
R21269 VDD.n115 VDD.t619 81.017
R21270 VDD.n12472 VDD.t1505 81.017
R21271 VDD.t2076 VDD.n12469 81.017
R21272 VDD.t1052 VDD.n116 81.017
R21273 VDD.t823 VDD.n12462 81.017
R21274 VDD.n12461 VDD.t1127 81.017
R21275 VDD.n8538 VDD.t810 81.017
R21276 VDD.n8537 VDD.t1195 81.017
R21277 VDD.t1333 VDD.n8530 81.017
R21278 VDD.n8529 VDD.t1265 81.017
R21279 VDD.t1015 VDD.n8881 81.017
R21280 VDD.n8880 VDD.t1818 81.017
R21281 VDD.t979 VDD.n8511 81.017
R21282 VDD.n8510 VDD.t1251 81.017
R21283 VDD.t1042 VDD.n9012 81.017
R21284 VDD.n9011 VDD.t1824 81.017
R21285 VDD.t2447 VDD.n8493 81.017
R21286 VDD.n8492 VDD.t1917 81.017
R21287 VDD.t603 VDD.n8462 81.017
R21288 VDD.t1867 VDD.n9179 81.017
R21289 VDD.t16 VDD.t27 79.7265
R21290 VDD.t14 VDD.t32 79.7265
R21291 VDD.t407 VDD.t390 79.5362
R21292 VDD.n11029 VDD.t335 70.2717
R21293 VDD.t520 VDD.n11004 70.2717
R21294 VDD.n1831 VDD.t298 70.2717
R21295 VDD.n1849 VDD.t499 70.2717
R21296 VDD.t555 VDD.n10949 70.2717
R21297 VDD.n1896 VDD.t1442 70.2717
R21298 VDD.n1914 VDD.t571 70.2717
R21299 VDD.t363 VDD.n10894 70.2717
R21300 VDD.n1923 VDD.t866 70.2717
R21301 VDD.n1941 VDD.t3013 70.2717
R21302 VDD.t2921 VDD.n10839 70.2717
R21303 VDD.n1988 VDD.t508 70.2717
R21304 VDD.n2014 VDD.t290 70.2717
R21305 VDD.t1711 VDD.n10781 70.2717
R21306 VDD.n10773 VDD.t303 70.2717
R21307 VDD.n15 VDD.t536 70.2717
R21308 VDD.n33 VDD.t1540 70.2717
R21309 VDD.t524 VDD.n12527 70.2717
R21310 VDD.n12520 VDD.t2240 70.2717
R21311 VDD.n113 VDD.t549 70.2717
R21312 VDD.t1708 VDD.n12471 70.2717
R21313 VDD.n12464 VDD.t2382 70.2717
R21314 VDD.n8535 VDD.t2812 70.2717
R21315 VDD.n8807 VDD.t6 70.2717
R21316 VDD.n8879 VDD.t544 70.2717
R21317 VDD.n8938 VDD.t367 70.2717
R21318 VDD.n9010 VDD.t707 70.2717
R21319 VDD.n9035 VDD.t2061 70.2717
R21320 VDD.n9159 VDD.t2127 70.2717
R21321 VDD.n9180 VDD.t2088 70.2717
R21322 VDD.n11028 VDD.t336 64.1315
R21323 VDD.n11003 VDD.t519 64.1315
R21324 VDD.n10997 VDD.t293 64.1315
R21325 VDD.t498 VDD.n1850 64.1315
R21326 VDD.n10948 VDD.t554 64.1315
R21327 VDD.n10942 VDD.t3354 64.1315
R21328 VDD.t3570 VDD.n1915 64.1315
R21329 VDD.n10893 VDD.t353 64.1315
R21330 VDD.n10887 VDD.t1338 64.1315
R21331 VDD.t664 VDD.n1942 64.1315
R21332 VDD.n10838 VDD.t1405 64.1315
R21333 VDD.n10832 VDD.t510 64.1315
R21334 VDD.t289 VDD.n2015 64.1315
R21335 VDD.n10780 VDD.t3613 64.1315
R21336 VDD.n10774 VDD.t326 64.1315
R21337 VDD.n12613 VDD.t537 64.1315
R21338 VDD.t845 VDD.n34 64.1315
R21339 VDD.n12526 VDD.t529 64.1315
R21340 VDD.n12519 VDD.t2422 64.1315
R21341 VDD.t547 VDD.n114 64.1315
R21342 VDD.n12470 VDD.t1850 64.1315
R21343 VDD.n12463 VDD.t502 64.1315
R21344 VDD.t2021 VDD.n8536 64.1315
R21345 VDD.n8806 VDD.t2 64.1315
R21346 VDD.n8882 VDD.t545 64.1315
R21347 VDD.n8937 VDD.t301 64.1315
R21348 VDD.n9013 VDD.t2288 64.1315
R21349 VDD.n9034 VDD.t2189 64.1315
R21350 VDD.n9158 VDD.t2302 64.1315
R21351 VDD.t2228 VDD.n9181 64.1315
R21352 VDD.t405 VDD.t402 54.0391
R21353 VDD.t38 VDD.t12 54.0391
R21354 VDD.t18 VDD.t16 54.0391
R21355 VDD.t23 VDD.t14 54.0391
R21356 VDD.t32 VDD.t25 54.0391
R21357 VDD.t25 VDD.t20 54.0391
R21358 VDD.t20 VDD.t34 54.0391
R21359 VDD.n7995 VDD.t27 50.3287
R21360 VDD.n6633 VDD.n5268 46.8594
R21361 VDD.t962 VDD.n2123 45.4522
R21362 VDD.t925 VDD.n2188 45.3596
R21363 VDD.n2354 VDD.t568 45.2864
R21364 VDD.t910 VDD.n2355 45.2864
R21365 VDD.n2356 VDD.t18 42.0517
R21366 VDD.t683 VDD.t472 38.7904
R21367 VDD.t742 VDD.t470 38.7904
R21368 VDD.t689 VDD.t468 38.7904
R21369 VDD.t656 VDD.t471 38.7904
R21370 VDD.t878 VDD.t474 38.7904
R21371 VDD.t469 VDD.t557 38.7904
R21372 VDD.t316 VDD.t563 38.7904
R21373 VDD.t307 VDD.t818 38.7904
R21374 VDD.t315 VDD.t700 38.7904
R21375 VDD.t653 VDD.t306 38.7904
R21376 VDD.t661 VDD.t311 38.7904
R21377 VDD.t574 VDD.t310 38.7904
R21378 VDD.n8077 VDD.t402 37.9607
R21379 VDD.t472 VDD.t427 36.32
R21380 VDD.t470 VDD.t423 36.32
R21381 VDD.t468 VDD.t425 36.32
R21382 VDD.t471 VDD.t429 36.32
R21383 VDD.t474 VDD.t439 36.32
R21384 VDD.t434 VDD.t469 36.32
R21385 VDD.t314 VDD.t316 36.32
R21386 VDD.t317 VDD.t307 36.32
R21387 VDD.t341 VDD.t315 36.32
R21388 VDD.t306 VDD.t312 36.32
R21389 VDD.t311 VDD.t309 36.32
R21390 VDD.t310 VDD.t320 36.32
R21391 VDD.t586 VDD.t393 31.8205
R21392 VDD.t839 VDD.t395 31.8205
R21393 VDD.t616 VDD.t391 31.8205
R21394 VDD.t398 VDD.t613 31.8205
R21395 VDD.t886 VDD.t82 31.8205
R21396 VDD.t70 VDD.t583 31.8205
R21397 VDD.t49 VDD.t883 31.8205
R21398 VDD.t55 VDD.t593 31.8205
R21399 VDD.t406 VDD.t410 29.7939
R21400 VDD.t397 VDD.t401 29.7939
R21401 VDD.t403 VDD.t404 29.7939
R21402 VDD.t396 VDD.t400 29.7939
R21403 VDD.t60 VDD.t78 29.7939
R21404 VDD.t64 VDD.t47 29.7939
R21405 VDD.t76 VDD.t62 29.7939
R21406 VDD.t58 VDD.t120 29.7939
R21407 VDD.n10996 VDD.n10995 29.1665
R21408 VDD.n10941 VDD.n10940 29.1665
R21409 VDD.n10886 VDD.n10885 29.1665
R21410 VDD.n10831 VDD.n10830 29.1665
R21411 VDD.n12525 VDD.n36 29.1665
R21412 VDD.n12469 VDD.n116 29.1665
R21413 VDD.n8530 VDD.n8529 29.1665
R21414 VDD.n9012 VDD.n9011 29.1665
R21415 VDD.t427 VDD.t432 24.618
R21416 VDD.t425 VDD.t442 24.618
R21417 VDD.t439 VDD.t444 24.618
R21418 VDD.t318 VDD.t314 24.618
R21419 VDD.t319 VDD.t341 24.618
R21420 VDD.t309 VDD.t313 24.618
R21421 VDD.n11005 VDD.n1786 24.5613
R21422 VDD.n11002 VDD.n1787 24.5613
R21423 VDD.n10950 VDD.n1851 24.5613
R21424 VDD.n10947 VDD.n1852 24.5613
R21425 VDD.n10895 VDD.n1916 24.5613
R21426 VDD.n10892 VDD.n1917 24.5613
R21427 VDD.n10840 VDD.n1943 24.5613
R21428 VDD.n10837 VDD.n1944 24.5613
R21429 VDD.n10782 VDD.n2016 24.5613
R21430 VDD.n10779 VDD.n2017 24.5613
R21431 VDD.n12612 VDD.n12611 24.5613
R21432 VDD.n12528 VDD.n35 24.5613
R21433 VDD.n12518 VDD.n12517 24.5613
R21434 VDD.n12472 VDD.n115 24.5613
R21435 VDD.n12462 VDD.n12461 24.5613
R21436 VDD.n8538 VDD.n8537 24.5613
R21437 VDD.n8881 VDD.n8880 24.5613
R21438 VDD.n8511 VDD.n8510 24.5613
R21439 VDD.n8493 VDD.n8492 24.5613
R21440 VDD.n9179 VDD.n8462 24.5613
R21441 VDD.n1742 VDD.t423 24.0112
R21442 VDD.n1718 VDD.t429 24.0112
R21443 VDD.n1414 VDD.t434 24.0112
R21444 VDD.n1356 VDD.t317 24.0112
R21445 VDD.n1349 VDD.t312 24.0112
R21446 VDD.n1652 VDD.t320 24.0112
R21447 VDD.n690 VDD.t683 20.6307
R21448 VDD.n709 VDD.t742 20.6307
R21449 VDD.n1719 VDD.t689 20.6307
R21450 VDD.n874 VDD.t656 20.6307
R21451 VDD.n1415 VDD.t878 20.6307
R21452 VDD.n1429 VDD.t557 20.6307
R21453 VDD.n1428 VDD.t563 20.6307
R21454 VDD.t818 VDD.n1354 20.6307
R21455 VDD.t700 VDD.n1084 20.6307
R21456 VDD.n1346 VDD.t653 20.6307
R21457 VDD.n1345 VDD.t661 20.6307
R21458 VDD.n763 VDD.t574 20.6307
R21459 VDD.t393 VDD.t416 20.1946
R21460 VDD.t416 VDD.t394 20.1946
R21461 VDD.t394 VDD.t406 20.1946
R21462 VDD.t401 VDD.t413 20.1946
R21463 VDD.t412 VDD.t397 20.1946
R21464 VDD.t399 VDD.t412 20.1946
R21465 VDD.t395 VDD.t399 20.1946
R21466 VDD.t391 VDD.t415 20.1946
R21467 VDD.t415 VDD.t392 20.1946
R21468 VDD.t392 VDD.t403 20.1946
R21469 VDD.t409 VDD.t396 20.1946
R21470 VDD.t400 VDD.t408 20.1946
R21471 VDD.t408 VDD.t411 20.1946
R21472 VDD.t411 VDD.t398 20.1946
R21473 VDD.t82 VDD.t137 20.1946
R21474 VDD.t137 VDD.t68 20.1946
R21475 VDD.t68 VDD.t60 20.1946
R21476 VDD.t96 VDD.t64 20.1946
R21477 VDD.t47 VDD.t53 20.1946
R21478 VDD.t53 VDD.t115 20.1946
R21479 VDD.t115 VDD.t70 20.1946
R21480 VDD.t66 VDD.t49 20.1946
R21481 VDD.t134 VDD.t66 20.1946
R21482 VDD.t62 VDD.t134 20.1946
R21483 VDD.t73 VDD.t58 20.1946
R21484 VDD.t120 VDD.t51 20.1946
R21485 VDD.t51 VDD.t122 20.1946
R21486 VDD.t122 VDD.t55 20.1946
R21487 VDD.n6396 VDD.t410 19.0569
R21488 VDD.n6577 VDD.t404 19.0569
R21489 VDD.n7040 VDD.t78 19.0569
R21490 VDD.n7086 VDD.t76 19.0569
R21491 VDD.n6311 VDD.t586 16.9237
R21492 VDD.n5376 VDD.t839 16.9237
R21493 VDD.n6370 VDD.t616 16.9237
R21494 VDD.t613 VDD.n5268 16.9237
R21495 VDD.n6633 VDD.t886 16.9237
R21496 VDD.n7133 VDD.t883 16.9237
R21497 VDD.n7834 VDD.t593 16.9237
R21498 VDD.n8077 VDD.t407 16.0789
R21499 VDD.t583 VDD.n2356 15.3594
R21500 VDD.n2355 VDD.n2354 13.7004
R21501 VDD.n2356 VDD.t38 11.9879
R21502 VDD.n696 VDD.t487 10.8219
R21503 VDD.n949 VDD.t476 10.378
R21504 VDD.n1448 VDD.t386 9.30374
R21505 VDD.n11029 VDD.n11028 8.52856
R21506 VDD.n11004 VDD.n11003 8.52856
R21507 VDD.n10997 VDD.n1831 8.52856
R21508 VDD.n1850 VDD.n1849 8.52856
R21509 VDD.n10949 VDD.n10948 8.52856
R21510 VDD.n10942 VDD.n1896 8.52856
R21511 VDD.n1915 VDD.n1914 8.52856
R21512 VDD.n10894 VDD.n10893 8.52856
R21513 VDD.n10887 VDD.n1923 8.52856
R21514 VDD.n1942 VDD.n1941 8.52856
R21515 VDD.n10839 VDD.n10838 8.52856
R21516 VDD.n10832 VDD.n1988 8.52856
R21517 VDD.n2015 VDD.n2014 8.52856
R21518 VDD.n10781 VDD.n10780 8.52856
R21519 VDD.n10774 VDD.n10773 8.52856
R21520 VDD.n12613 VDD.n15 8.52856
R21521 VDD.n34 VDD.n33 8.52856
R21522 VDD.n12527 VDD.n12526 8.52856
R21523 VDD.n12520 VDD.n12519 8.52856
R21524 VDD.n114 VDD.n113 8.52856
R21525 VDD.n12471 VDD.n12470 8.52856
R21526 VDD.n12464 VDD.n12463 8.52856
R21527 VDD.n8536 VDD.n8535 8.52856
R21528 VDD.n8807 VDD.n8806 8.52856
R21529 VDD.n8882 VDD.n8879 8.52856
R21530 VDD.n8938 VDD.n8937 8.52856
R21531 VDD.n9013 VDD.n9010 8.52856
R21532 VDD.n9035 VDD.n9034 8.52856
R21533 VDD.n9159 VDD.n9158 8.52856
R21534 VDD.n9181 VDD.n9180 8.52856
R21535 VDD.n1442 VDD.t3073 8.19583
R21536 VDD.n1478 VDD.t2763 8.14522
R21537 VDD.t1066 VDD.n1611 8.14522
R21538 VDD.n1609 VDD.t3835 8.14522
R21539 VDD.n1477 VDD.t4069 8.14522
R21540 VDD.t1168 VDD.n1751 8.11081
R21541 VDD VDD.t3999 8.10685
R21542 VDD.n1752 VDD.t1168 8.10567
R21543 VDD.n969 VDD.t3580 8.10567
R21544 VDD.t3580 VDD.n682 8.10567
R21545 VDD.n971 VDD.t2544 8.10567
R21546 VDD.t2544 VDD.n970 8.10567
R21547 VDD.n973 VDD.t2667 8.10567
R21548 VDD.t2667 VDD.n972 8.10567
R21549 VDD.n975 VDD.t1430 8.10567
R21550 VDD.t1430 VDD.n974 8.10567
R21551 VDD.n977 VDD.t1559 8.10567
R21552 VDD.t1559 VDD.n976 8.10567
R21553 VDD.n987 VDD.t4609 8.10567
R21554 VDD.t4609 VDD.n986 8.10567
R21555 VDD.n989 VDD.t805 8.10567
R21556 VDD.t805 VDD.n988 8.10567
R21557 VDD.n991 VDD.t3845 8.10567
R21558 VDD.t3845 VDD.n990 8.10567
R21559 VDD.n993 VDD.t3977 8.10567
R21560 VDD.t3977 VDD.n992 8.10567
R21561 VDD.n995 VDD.t2930 8.10567
R21562 VDD.t2930 VDD.n994 8.10567
R21563 VDD.n997 VDD.t937 8.10567
R21564 VDD.t937 VDD.n996 8.10567
R21565 VDD.n1006 VDD.t682 8.10567
R21566 VDD.t682 VDD.n1005 8.10567
R21567 VDD.n1008 VDD.t3329 8.10567
R21568 VDD.t3329 VDD.n1007 8.10567
R21569 VDD.n1010 VDD.t2223 8.10567
R21570 VDD.t2223 VDD.n1009 8.10567
R21571 VDD.n1012 VDD.t2621 8.10567
R21572 VDD.t2621 VDD.n1011 8.10567
R21573 VDD.n1014 VDD.t2497 8.10567
R21574 VDD.t2497 VDD.n1013 8.10567
R21575 VDD.n1016 VDD.t2627 8.10567
R21576 VDD.t2627 VDD.n1015 8.10567
R21577 VDD.t1396 VDD.n1030 8.10567
R21578 VDD.n1031 VDD.t1396 8.10567
R21579 VDD.t1509 VDD.n1028 8.10567
R21580 VDD.n1029 VDD.t1509 8.10567
R21581 VDD.t4543 VDD.n1026 8.10567
R21582 VDD.n1027 VDD.t4543 8.10567
R21583 VDD.t2565 VDD.n1024 8.10567
R21584 VDD.n1025 VDD.t2565 8.10567
R21585 VDD.t1340 VDD.n1022 8.10567
R21586 VDD.n1023 VDD.t1340 8.10567
R21587 VDD.t3999 VDD.n12643 8.10567
R21588 VDD.n12563 VDD.t1480 8.10567
R21589 VDD.n12563 VDD.t832 8.10567
R21590 VDD.n12566 VDD.t1847 8.10567
R21591 VDD.n12566 VDD.t1161 8.10567
R21592 VDD.n12567 VDD.t2561 8.10567
R21593 VDD.n12567 VDD.t1765 8.10567
R21594 VDD.n12573 VDD.t1860 8.10567
R21595 VDD.n12573 VDD.t1172 8.10567
R21596 VDD.n12574 VDD.t2294 8.10567
R21597 VDD.n12574 VDD.t1535 8.10567
R21598 VDD.n12577 VDD.t3851 8.10567
R21599 VDD.n12577 VDD.t3217 8.10567
R21600 VDD.n8633 VDD.t1807 8.10567
R21601 VDD.n8634 VDD.t2639 8.10567
R21602 VDD.n12617 VDD.t1464 8.10567
R21603 VDD.n11 VDD.t2663 8.10567
R21604 VDD.n8630 VDD.t1569 8.10567
R21605 VDD.n8630 VDD.t3123 8.10567
R21606 VDD.n8627 VDD.t1938 8.10567
R21607 VDD.n8627 VDD.t3437 8.10567
R21608 VDD.n8626 VDD.t2651 8.10567
R21609 VDD.n8626 VDD.t4043 8.10567
R21610 VDD.n12606 VDD.t1965 8.10567
R21611 VDD.n12606 VDD.t3447 8.10567
R21612 VDD.n12605 VDD.t2413 8.10567
R21613 VDD.n12605 VDD.t3805 8.10567
R21614 VDD.n12602 VDD.t3943 8.10567
R21615 VDD.n12602 VDD.t1217 8.10567
R21616 VDD.n8630 VDD.t1779 8.10567
R21617 VDD.n8630 VDD.t2994 8.10567
R21618 VDD.n8627 VDD.t2180 8.10567
R21619 VDD.n8627 VDD.t3297 8.10567
R21620 VDD.n8626 VDD.t2862 8.10567
R21621 VDD.n8626 VDD.t3871 8.10567
R21622 VDD.n12606 VDD.t2203 8.10567
R21623 VDD.n12606 VDD.t3307 8.10567
R21624 VDD.n12605 VDD.t2643 8.10567
R21625 VDD.n12605 VDD.t3637 8.10567
R21626 VDD.n12602 VDD.t4171 8.10567
R21627 VDD.n12602 VDD.t1085 8.10567
R21628 VDD.n12555 VDD.t4187 8.10567
R21629 VDD.n12595 VDD.t752 8.10567
R21630 VDD.n12556 VDD.t3827 8.10567
R21631 VDD.n12588 VDD.t777 8.10567
R21632 VDD.n12545 VDD.t4265 8.10567
R21633 VDD.n25 VDD.t844 8.10567
R21634 VDD.n12551 VDD.t3915 8.10567
R21635 VDD.n24 VDD.t1289 8.10567
R21636 VDD.n8661 VDD.t3370 8.10567
R21637 VDD.n8661 VDD.t3207 8.10567
R21638 VDD.n8658 VDD.t3718 8.10567
R21639 VDD.n8658 VDD.t3507 8.10567
R21640 VDD.n8657 VDD.t4327 8.10567
R21641 VDD.n8657 VDD.t4133 8.10567
R21642 VDD.n12534 VDD.t3734 8.10567
R21643 VDD.n12534 VDD.t3527 8.10567
R21644 VDD.n12535 VDD.t4127 8.10567
R21645 VDD.n12535 VDD.t3891 8.10567
R21646 VDD.n12539 VDD.t1514 8.10567
R21647 VDD.n12539 VDD.t1298 8.10567
R21648 VDD.n8661 VDD.t1883 8.10567
R21649 VDD.n8661 VDD.t3063 8.10567
R21650 VDD.n8658 VDD.t2285 8.10567
R21651 VDD.n8658 VDD.t3356 8.10567
R21652 VDD.n8657 VDD.t2958 8.10567
R21653 VDD.n8657 VDD.t3973 8.10567
R21654 VDD.n12534 VDD.t2318 8.10567
R21655 VDD.n12534 VDD.t3372 8.10567
R21656 VDD.n12535 VDD.t2737 8.10567
R21657 VDD.n12535 VDD.t3740 8.10567
R21658 VDD.n12539 VDD.t4251 8.10567
R21659 VDD.n12539 VDD.t1154 8.10567
R21660 VDD.n8621 VDD.t1903 8.10567
R21661 VDD.n8651 VDD.t2733 8.10567
R21662 VDD.n8622 VDD.t1539 8.10567
R21663 VDD.n8645 VDD.t3189 8.10567
R21664 VDD.n8619 VDD.t3680 8.10567
R21665 VDD.n8672 VDD.t727 8.10567
R21666 VDD.n8620 VDD.t3345 8.10567
R21667 VDD.n8666 VDD.t763 8.10567
R21668 VDD.n8616 VDD.t4063 8.10567
R21669 VDD.n8616 VDD.t3841 8.10567
R21670 VDD.n8613 VDD.t4389 8.10567
R21671 VDD.n8613 VDD.t4211 8.10567
R21672 VDD.n8612 VDD.t890 8.10567
R21673 VDD.n8612 VDD.t634 8.10567
R21674 VDD.n80 VDD.t4403 8.10567
R21675 VDD.n80 VDD.t4229 8.10567
R21676 VDD.n81 VDD.t624 8.10567
R21677 VDD.n81 VDD.t4549 8.10567
R21678 VDD.n85 VDD.t2263 8.10567
R21679 VDD.n85 VDD.t2031 8.10567
R21680 VDD.n8616 VDD.t685 8.10567
R21681 VDD.n8616 VDD.t3467 8.10567
R21682 VDD.n8613 VDD.t1056 8.10567
R21683 VDD.n8613 VDD.t3799 8.10567
R21684 VDD.n8612 VDD.t1648 8.10567
R21685 VDD.n8612 VDD.t4399 8.10567
R21686 VDD.n80 VDD.t1074 8.10567
R21687 VDD.n80 VDD.t3819 8.10567
R21688 VDD.n81 VDD.t1414 8.10567
R21689 VDD.n81 VDD.t4219 8.10567
R21690 VDD.n85 VDD.t3103 8.10567
R21691 VDD.n85 VDD.t1610 8.10567
R21692 VDD.n73 VDD.t1852 8.10567
R21693 VDD.n54 VDD.t3127 8.10567
R21694 VDD.n47 VDD.t1491 8.10567
R21695 VDD.n48 VDD.t3151 8.10567
R21696 VDD.n12499 VDD.t794 8.10567
R21697 VDD.n12501 VDD.t2421 8.10567
R21698 VDD.n45 VDD.t2239 8.10567
R21699 VDD.n91 VDD.t1995 8.10567
R21700 VDD.n8694 VDD.t1652 8.10567
R21701 VDD.n8694 VDD.t1423 8.10567
R21702 VDD.n8691 VDD.t2033 8.10567
R21703 VDD.n8691 VDD.t1775 8.10567
R21704 VDD.n8690 VDD.t2722 8.10567
R21705 VDD.n8690 VDD.t2509 8.10567
R21706 VDD.n12512 VDD.t2053 8.10567
R21707 VDD.n12512 VDD.t1789 8.10567
R21708 VDD.n12511 VDD.t2499 8.10567
R21709 VDD.n12511 VDD.t2219 8.10567
R21710 VDD.n12508 VDD.t4015 8.10567
R21711 VDD.n12508 VDD.t3793 8.10567
R21712 VDD.n8694 VDD.t4353 8.10567
R21713 VDD.n8694 VDD.t4165 8.10567
R21714 VDD.n8691 VDD.t4703 8.10567
R21715 VDD.n8691 VDD.t4481 8.10567
R21716 VDD.n8690 VDD.t1152 8.10567
R21717 VDD.n8690 VDD.t983 8.10567
R21718 VDD.n12512 VDD.t4721 8.10567
R21719 VDD.n12512 VDD.t4489 8.10567
R21720 VDD.n12511 VDD.t975 8.10567
R21721 VDD.n12511 VDD.t747 8.10567
R21722 VDD.n12508 VDD.t2633 8.10567
R21723 VDD.n12508 VDD.t2407 8.10567
R21724 VDD.n8608 VDD.t2682 8.10567
R21725 VDD.n8684 VDD.t4181 8.10567
R21726 VDD.n8609 VDD.t4047 8.10567
R21727 VDD.n8678 VDD.t3817 8.10567
R21728 VDD.n8605 VDD.t2787 8.10567
R21729 VDD.n8710 VDD.t4259 8.10567
R21730 VDD.n8606 VDD.t1631 8.10567
R21731 VDD.n8704 VDD.t1402 8.10567
R21732 VDD.n8602 VDD.t4147 8.10567
R21733 VDD.n8602 VDD.t1504 8.10567
R21734 VDD.n8599 VDD.t4469 8.10567
R21735 VDD.n8599 VDD.t1873 8.10567
R21736 VDD.n8598 VDD.t967 8.10567
R21737 VDD.n8598 VDD.t2597 8.10567
R21738 VDD.n12478 VDD.t4483 8.10567
R21739 VDD.n12478 VDD.t1890 8.10567
R21740 VDD.n12479 VDD.t724 8.10567
R21741 VDD.n12479 VDD.t2346 8.10567
R21742 VDD.n12483 VDD.t2384 8.10567
R21743 VDD.n12483 VDD.t3877 8.10567
R21744 VDD.n8602 VDD.t4439 8.10567
R21745 VDD.n8602 VDD.t4245 8.10567
R21746 VDD.n8599 VDD.t618 8.10567
R21747 VDD.n8599 VDD.t4547 8.10567
R21748 VDD.n8598 VDD.t1232 8.10567
R21749 VDD.n8598 VDD.t1046 8.10567
R21750 VDD.n12478 VDD.t650 8.10567
R21751 VDD.n12478 VDD.t4573 8.10567
R21752 VDD.n12479 VDD.t1035 8.10567
R21753 VDD.n12479 VDD.t827 8.10567
R21754 VDD.n12483 VDD.t2712 8.10567
R21755 VDD.n12483 VDD.t2495 8.10567
R21756 VDD.n12489 VDD.t902 8.10567
R21757 VDD.n105 VDD.t2521 8.10567
R21758 VDD.n12495 VDD.t3995 8.10567
R21759 VDD.n104 VDD.t3771 8.10567
R21760 VDD.n162 VDD.t2728 8.10567
R21761 VDD.n143 VDD.t4227 8.10567
R21762 VDD.n136 VDD.t4077 8.10567
R21763 VDD.n137 VDD.t3857 8.10567
R21764 VDD.n8732 VDD.t3629 8.10567
R21765 VDD.n8732 VDD.t1051 8.10567
R21766 VDD.n8729 VDD.t4007 8.10567
R21767 VDD.n8729 VDD.t1382 8.10567
R21768 VDD.n8728 VDD.t4585 8.10567
R21769 VDD.n8728 VDD.t2012 8.10567
R21770 VDD.n126 VDD.t4029 8.10567
R21771 VDD.n126 VDD.t1392 8.10567
R21772 VDD.n127 VDD.t4375 8.10567
R21773 VDD.n127 VDD.t1763 8.10567
R21774 VDD.n131 VDD.t1786 8.10567
R21775 VDD.n131 VDD.t3392 8.10567
R21776 VDD.n8732 VDD.t2075 8.10567
R21777 VDD.n8732 VDD.t1820 8.10567
R21778 VDD.n8729 VDD.t2493 8.10567
R21779 VDD.n8729 VDD.t2217 8.10567
R21780 VDD.n8728 VDD.t3095 8.10567
R21781 VDD.n8728 VDD.t2890 8.10567
R21782 VDD.n126 VDD.t2513 8.10567
R21783 VDD.n126 VDD.t2235 8.10567
R21784 VDD.n127 VDD.t2878 8.10567
R21785 VDD.n127 VDD.t2671 8.10567
R21786 VDD.n131 VDD.t4381 8.10567
R21787 VDD.n131 VDD.t4195 8.10567
R21788 VDD.n8594 VDD.t4453 8.10567
R21789 VDD.n8722 VDD.t1849 8.10567
R21790 VDD.n8595 VDD.t1707 8.10567
R21791 VDD.n8716 VDD.t1485 8.10567
R21792 VDD.n8592 VDD.t2343 8.10567
R21793 VDD.n8743 VDD.t3849 8.10567
R21794 VDD.n8593 VDD.t2381 8.10567
R21795 VDD.n8737 VDD.t2096 8.10567
R21796 VDD.n8589 VDD.t4217 8.10567
R21797 VDD.n8589 VDD.t1126 8.10567
R21798 VDD.n8586 VDD.t4523 8.10567
R21799 VDD.n8586 VDD.t1458 8.10567
R21800 VDD.n8585 VDD.t1019 8.10567
R21801 VDD.n8585 VDD.t2105 8.10567
R21802 VDD.n12456 VDD.t4531 8.10567
R21803 VDD.n12456 VDD.t1474 8.10567
R21804 VDD.n12455 VDD.t791 8.10567
R21805 VDD.n12455 VDD.t1858 8.10567
R21806 VDD.n12452 VDD.t2453 8.10567
R21807 VDD.n12452 VDD.t3485 8.10567
R21808 VDD.n8589 VDD.t2714 8.10567
R21809 VDD.n8589 VDD.t3825 8.10567
R21810 VDD.n8586 VDD.t3057 8.10567
R21811 VDD.n8586 VDD.t4193 8.10567
R21812 VDD.n8585 VDD.t3600 8.10567
R21813 VDD.n8585 VDD.t609 8.10567
R21814 VDD.n12456 VDD.t3075 8.10567
R21815 VDD.n12456 VDD.t4215 8.10567
R21816 VDD.n12455 VDD.t3384 8.10567
R21817 VDD.n12455 VDD.t4533 8.10567
R21818 VDD.n12452 VDD.t822 8.10567
R21819 VDD.n12452 VDD.t2002 8.10567
R21820 VDD.n669 VDD.t3125 8.10567
R21821 VDD.n669 VDD.t1669 8.10567
R21822 VDD.n11063 VDD.t2797 8.10567
R21823 VDD.n11063 VDD.t1309 8.10567
R21824 VDD.n661 VDD.t1098 8.10567
R21825 VDD.n661 VDD.t3881 8.10567
R21826 VDD.n11097 VDD.t2789 8.10567
R21827 VDD.n11097 VDD.t1292 8.10567
R21828 VDD.n651 VDD.t2390 8.10567
R21829 VDD.n651 VDD.t964 8.10567
R21830 VDD.n11119 VDD.t2041 8.10567
R21831 VDD.n11119 VDD.t3941 8.10567
R21832 VDD.n5717 VDD.t4221 8.10567
R21833 VDD.n5718 VDD.t1753 8.10567
R21834 VDD.n11033 VDD.t1240 8.10567
R21835 VDD.n1769 VDD.t3590 8.10567
R21836 VDD.n5714 VDD.t2611 8.10567
R21837 VDD.n5714 VDD.t2124 8.10567
R21838 VDD.n5711 VDD.t2182 8.10567
R21839 VDD.n5711 VDD.t1738 8.10567
R21840 VDD.n5710 VDD.t4701 8.10567
R21841 VDD.n5710 VDD.t4305 8.10567
R21842 VDD.n11011 VDD.t2166 8.10567
R21843 VDD.n11011 VDD.t1728 8.10567
R21844 VDD.n11012 VDD.t1746 8.10567
R21845 VDD.n11012 VDD.t1353 8.10567
R21846 VDD.n11016 VDD.t2866 8.10567
R21847 VDD.n11016 VDD.t2067 8.10567
R21848 VDD.n5714 VDD.t2487 8.10567
R21849 VDD.n5714 VDD.t4705 8.10567
R21850 VDD.n5711 VDD.t2065 8.10567
R21851 VDD.n5711 VDD.t4357 8.10567
R21852 VDD.n5710 VDD.t4559 8.10567
R21853 VDD.n5710 VDD.t2834 8.10567
R21854 VDD.n11011 VDD.t2045 8.10567
R21855 VDD.n11011 VDD.t4347 8.10567
R21856 VDD.n11012 VDD.t1641 8.10567
R21857 VDD.n11012 VDD.t3981 8.10567
R21858 VDD.n11016 VDD.t2361 8.10567
R21859 VDD.n11016 VDD.t1418 8.10567
R21860 VDD.n11022 VDD.t3692 8.10567
R21861 VDD.n1779 VDD.t2613 8.10567
R21862 VDD.n1773 VDD.t580 8.10567
R21863 VDD.n1775 VDD.t3945 8.10567
R21864 VDD.n1806 VDD.t4451 8.10567
R21865 VDD.n1820 VDD.t3315 8.10567
R21866 VDD.n1807 VDD.t1356 8.10567
R21867 VDD.n1814 VDD.t1553 8.10567
R21868 VDD.n5740 VDD.t4355 8.10567
R21869 VDD.n5740 VDD.t1557 8.10567
R21870 VDD.n5737 VDD.t4019 8.10567
R21871 VDD.n5737 VDD.t1199 8.10567
R21872 VDD.n5736 VDD.t2484 8.10567
R21873 VDD.n5736 VDD.t3777 8.10567
R21874 VDD.n1797 VDD.t4001 8.10567
R21875 VDD.n1797 VDD.t1190 8.10567
R21876 VDD.n1798 VDD.t3619 8.10567
R21877 VDD.n1798 VDD.t851 8.10567
R21878 VDD.n1802 VDD.t4033 8.10567
R21879 VDD.n1802 VDD.t2884 8.10567
R21880 VDD.n5740 VDD.t1845 8.10567
R21881 VDD.n5740 VDD.t4189 8.10567
R21882 VDD.n5737 VDD.t1478 8.10567
R21883 VDD.n5737 VDD.t3823 8.10567
R21884 VDD.n5736 VDD.t4055 8.10567
R21885 VDD.n5736 VDD.t2233 8.10567
R21886 VDD.n1797 VDD.t1470 8.10567
R21887 VDD.n1797 VDD.t3809 8.10567
R21888 VDD.n1798 VDD.t1111 8.10567
R21889 VDD.n1798 VDD.t3449 8.10567
R21890 VDD.n1802 VDD.t3113 8.10567
R21891 VDD.n1802 VDD.t2230 8.10567
R21892 VDD.n5706 VDD.t3647 8.10567
R21893 VDD.n5730 VDD.t1224 8.10567
R21894 VDD.n5707 VDD.t729 8.10567
R21895 VDD.n5724 VDD.t1615 8.10567
R21896 VDD.n5753 VDD.t1315 8.10567
R21897 VDD.n5751 VDD.t1660 8.10567
R21898 VDD.n5705 VDD.t2655 8.10567
R21899 VDD.n5745 VDD.t3489 8.10567
R21900 VDD.n5701 VDD.t3947 8.10567
R21901 VDD.n5701 VDD.t1137 8.10567
R21902 VDD.n5698 VDD.t3584 8.10567
R21903 VDD.n5698 VDD.t803 8.10567
R21904 VDD.n5697 VDD.t1967 8.10567
R21905 VDD.n5697 VDD.t3351 8.10567
R21906 VDD.n10990 VDD.t3565 8.10567
R21907 VDD.n10990 VDD.t788 8.10567
R21908 VDD.n10989 VDD.t3245 8.10567
R21909 VDD.n10989 VDD.t4529 8.10567
R21910 VDD.n10986 VDD.t916 8.10567
R21911 VDD.n10986 VDD.t3843 8.10567
R21912 VDD.n5701 VDD.t744 8.10567
R21913 VDD.n5701 VDD.t943 8.10567
R21914 VDD.n5698 VDD.t4507 8.10567
R21915 VDD.n5698 VDD.t4711 8.10567
R21916 VDD.n5697 VDD.t3010 8.10567
R21917 VDD.n5697 VDD.t3167 8.10567
R21918 VDD.n10990 VDD.t4495 8.10567
R21919 VDD.n10990 VDD.t4697 8.10567
R21920 VDD.n10989 VDD.t4161 8.10567
R21921 VDD.n10989 VDD.t4325 8.10567
R21922 VDD.n10986 VDD.t4605 8.10567
R21923 VDD.n10986 VDD.t3139 8.10567
R21924 VDD.n10977 VDD.t1500 8.10567
R21925 VDD.n10979 VDD.t1384 8.10567
R21926 VDD.n1796 VDD.t2690 8.10567
R21927 VDD.n1826 VDD.t2886 8.10567
R21928 VDD.n10967 VDD.t1135 8.10567
R21929 VDD.n1841 VDD.t1328 8.10567
R21930 VDD.n10973 VDD.t3627 8.10567
R21931 VDD.n1840 VDD.t2517 8.10567
R21932 VDD.n5795 VDD.t1596 8.10567
R21933 VDD.n5795 VDD.t3067 8.10567
R21934 VDD.n5792 VDD.t1234 8.10567
R21935 VDD.n5792 VDD.t2726 8.10567
R21936 VDD.n5791 VDD.t3803 8.10567
R21937 VDD.n5791 VDD.t1029 8.10567
R21938 VDD.n10956 VDD.t1226 8.10567
R21939 VDD.n10956 VDD.t2704 8.10567
R21940 VDD.n10957 VDD.t892 8.10567
R21941 VDD.n10957 VDD.t2279 8.10567
R21942 VDD.n10961 VDD.t2122 8.10567
R21943 VDD.n10961 VDD.t934 8.10567
R21944 VDD.n5795 VDD.t3305 8.10567
R21945 VDD.n5795 VDD.t4641 8.10567
R21946 VDD.n5792 VDD.t3006 8.10567
R21947 VDD.n5792 VDD.t4291 8.10567
R21948 VDD.n5791 VDD.t1281 8.10567
R21949 VDD.n5791 VDD.t2776 8.10567
R21950 VDD.n10956 VDD.t2990 8.10567
R21951 VDD.n10956 VDD.t4279 8.10567
R21952 VDD.n10957 VDD.t2617 8.10567
R21953 VDD.n10957 VDD.t3909 8.10567
R21954 VDD.n10961 VDD.t1141 8.10567
R21955 VDD.n10961 VDD.t4125 8.10567
R21956 VDD.n5693 VDD.t1360 8.10567
R21957 VDD.n5785 VDD.t2363 8.10567
R21958 VDD.n5694 VDD.t2139 8.10567
R21959 VDD.n5779 VDD.t3523 8.10567
R21960 VDD.n5691 VDD.t868 8.10567
R21961 VDD.n5806 VDD.t1726 8.10567
R21962 VDD.n5692 VDD.t3983 8.10567
R21963 VDD.n5800 VDD.t1174 8.10567
R21964 VDD.n5688 VDD.t1517 8.10567
R21965 VDD.n5688 VDD.t2539 8.10567
R21966 VDD.n5685 VDD.t1170 8.10567
R21967 VDD.n5685 VDD.t2103 8.10567
R21968 VDD.n5684 VDD.t3736 8.10567
R21969 VDD.n5684 VDD.t4627 8.10567
R21970 VDD.n1880 VDD.t1157 8.10567
R21971 VDD.n1880 VDD.t2092 8.10567
R21972 VDD.n1881 VDD.t800 8.10567
R21973 VDD.n1881 VDD.t1685 8.10567
R21974 VDD.n1885 VDD.t1436 8.10567
R21975 VDD.n1885 VDD.t1657 8.10567
R21976 VDD.n5688 VDD.t2814 8.10567
R21977 VDD.n5688 VDD.t4129 8.10567
R21978 VDD.n5685 VDD.t2455 8.10567
R21979 VDD.n5685 VDD.t3759 8.10567
R21980 VDD.n5684 VDD.t779 8.10567
R21981 VDD.n5684 VDD.t2152 8.10567
R21982 VDD.n1880 VDD.t2442 8.10567
R21983 VDD.n1880 VDD.t3742 8.10567
R21984 VDD.n1881 VDD.t1981 8.10567
R21985 VDD.n1881 VDD.t3374 8.10567
R21986 VDD.n1885 VDD.t1901 8.10567
R21987 VDD.n1885 VDD.t696 8.10567
R21988 VDD.n1862 VDD.t1899 8.10567
R21989 VDD.n1876 VDD.t2115 8.10567
R21990 VDD.n1863 VDD.t702 8.10567
R21991 VDD.n1870 VDD.t3653 8.10567
R21992 VDD.n10922 VDD.t3199 8.10567
R21993 VDD.n10924 VDD.t3353 8.10567
R21994 VDD.n1861 VDD.t1441 8.10567
R21995 VDD.n1891 VDD.t4401 8.10567
R21996 VDD.n5850 VDD.t4103 8.10567
R21997 VDD.n5850 VDD.t854 8.10567
R21998 VDD.n5847 VDD.t3728 8.10567
R21999 VDD.n5847 VDD.t4621 8.10567
R22000 VDD.n5846 VDD.t2117 8.10567
R22001 VDD.n5846 VDD.t3093 8.10567
R22002 VDD.n10935 VDD.t3716 8.10567
R22003 VDD.n10935 VDD.t4601 8.10567
R22004 VDD.n10934 VDD.t3339 8.10567
R22005 VDD.n10934 VDD.t4253 8.10567
R22006 VDD.n10931 VDD.t2174 8.10567
R22007 VDD.n10931 VDD.t2440 8.10567
R22008 VDD.n5850 VDD.t4537 8.10567
R22009 VDD.n5850 VDD.t1767 8.10567
R22010 VDD.n5847 VDD.t4233 8.10567
R22011 VDD.n5847 VDD.t1410 8.10567
R22012 VDD.n5846 VDD.t2679 8.10567
R22013 VDD.n5846 VDD.t3991 8.10567
R22014 VDD.n10935 VDD.t4223 8.10567
R22015 VDD.n10935 VDD.t1398 8.10567
R22016 VDD.n10934 VDD.t3829 8.10567
R22017 VDD.n10934 VDD.t1048 8.10567
R22018 VDD.n10931 VDD.t3201 8.10567
R22019 VDD.n10931 VDD.t1923 8.10567
R22020 VDD.n5820 VDD.t2773 8.10567
R22021 VDD.n5818 VDD.t3592 8.10567
R22022 VDD.n5681 VDD.t3457 8.10567
R22023 VDD.n5812 VDD.t642 8.10567
R22024 VDD.n5678 VDD.t2923 8.10567
R22025 VDD.n5861 VDD.t3749 8.10567
R22026 VDD.n5679 VDD.t4625 8.10567
R22027 VDD.n5855 VDD.t1840 8.10567
R22028 VDD.n5675 VDD.t2137 8.10567
R22029 VDD.n5675 VDD.t4443 8.10567
R22030 VDD.n5672 VDD.t1751 8.10567
R22031 VDD.n5672 VDD.t4117 8.10567
R22032 VDD.n5671 VDD.t4319 8.10567
R22033 VDD.n5671 VDD.t2569 8.10567
R22034 VDD.n10901 VDD.t1736 8.10567
R22035 VDD.n10901 VDD.t4097 8.10567
R22036 VDD.n10902 VDD.t1364 8.10567
R22037 VDD.n10902 VDD.t3702 8.10567
R22038 VDD.n10906 VDD.t3975 8.10567
R22039 VDD.n10906 VDD.t3181 8.10567
R22040 VDD.n5675 VDD.t1600 8.10567
R22041 VDD.n5675 VDD.t1944 8.10567
R22042 VDD.n5672 VDD.t1238 8.10567
R22043 VDD.n5672 VDD.t1580 8.10567
R22044 VDD.n5671 VDD.t3813 8.10567
R22045 VDD.n5671 VDD.t4159 8.10567
R22046 VDD.n10901 VDD.t1228 8.10567
R22047 VDD.n10901 VDD.t1555 8.10567
R22048 VDD.n10902 VDD.t904 8.10567
R22049 VDD.n10902 VDD.t1182 8.10567
R22050 VDD.n10906 VDD.t2355 8.10567
R22051 VDD.n10906 VDD.t2172 8.10567
R22052 VDD.n10912 VDD.t3368 8.10567
R22053 VDD.n1906 VDD.t3569 8.10567
R22054 VDD.n10918 VDD.t570 8.10567
R22055 VDD.n1905 VDD.t3567 8.10567
R22056 VDD.n5510 VDD.t4561 8.10567
R22057 VDD.n5524 VDD.t3398 8.10567
R22058 VDD.n5511 VDD.t2972 8.10567
R22059 VDD.n5518 VDD.t607 8.10567
R22060 VDD.n5897 VDD.t1576 8.10567
R22061 VDD.n5897 VDD.t3921 8.10567
R22062 VDD.n5894 VDD.t1222 8.10567
R22063 VDD.n5894 VDD.t3563 8.10567
R22064 VDD.n5893 VDD.t3789 8.10567
R22065 VDD.n5893 VDD.t1935 8.10567
R22066 VDD.n5494 VDD.t1197 8.10567
R22067 VDD.n5494 VDD.t3545 8.10567
R22068 VDD.n5495 VDD.t874 8.10567
R22069 VDD.n5495 VDD.t3223 8.10567
R22070 VDD.n5499 VDD.t4709 8.10567
R22071 VDD.n5499 VDD.t3883 8.10567
R22072 VDD.n5897 VDD.t3939 8.10567
R22073 VDD.n5897 VDD.t3795 8.10567
R22074 VDD.n5894 VDD.t3578 8.10567
R22075 VDD.n5894 VDD.t3461 8.10567
R22076 VDD.n5893 VDD.t1956 8.10567
R22077 VDD.n5893 VDD.t1798 8.10567
R22078 VDD.n5494 VDD.t3555 8.10567
R22079 VDD.n5494 VDD.t3441 8.10567
R22080 VDD.n5495 VDD.t3239 8.10567
R22081 VDD.n5495 VDD.t3111 8.10567
R22082 VDD.n5499 VDD.t2111 8.10567
R22083 VDD.n5499 VDD.t3402 8.10567
R22084 VDD.n5667 VDD.t4675 8.10567
R22085 VDD.n5873 VDD.t1886 8.10567
R22086 VDD.n5668 VDD.t932 8.10567
R22087 VDD.n5867 VDD.t3696 8.10567
R22088 VDD.n5545 VDD.t2816 8.10567
R22089 VDD.n5543 VDD.t1337 8.10567
R22090 VDD.n5663 VDD.t865 8.10567
R22091 VDD.n5542 VDD.t3213 8.10567
R22092 VDD.n5633 VDD.t1027 8.10567
R22093 VDD.n5633 VDD.t2848 8.10567
R22094 VDD.n5630 VDD.t658 8.10567
R22095 VDD.n5630 VDD.t2491 8.10567
R22096 VDD.n5629 VDD.t3273 8.10567
R22097 VDD.n5629 VDD.t797 8.10567
R22098 VDD.n10880 VDD.t637 8.10567
R22099 VDD.n10880 VDD.t2482 8.10567
R22100 VDD.n10879 VDD.t4411 8.10567
R22101 VDD.n10879 VDD.t2023 8.10567
R22102 VDD.n10876 VDD.t4331 8.10567
R22103 VDD.n10876 VDD.t3215 8.10567
R22104 VDD.n5633 VDD.t1973 8.10567
R22105 VDD.n5633 VDD.t3293 8.10567
R22106 VDD.n5630 VDD.t1604 8.10567
R22107 VDD.n5630 VDD.t2986 8.10567
R22108 VDD.n5629 VDD.t4185 8.10567
R22109 VDD.n5629 VDD.t1261 8.10567
R22110 VDD.n10880 VDD.t1588 8.10567
R22111 VDD.n10880 VDD.t2964 8.10567
R22112 VDD.n10879 VDD.t1208 8.10567
R22113 VDD.n10879 VDD.t2595 8.10567
R22114 VDD.n10876 VDD.t3911 8.10567
R22115 VDD.n10876 VDD.t4167 8.10567
R22116 VDD.n10867 VDD.t2260 8.10567
R22117 VDD.n10869 VDD.t4163 8.10567
R22118 VDD.n5506 VDD.t2258 8.10567
R22119 VDD.n5504 VDD.t1377 8.10567
R22120 VDD.n10857 VDD.t2541 8.10567
R22121 VDD.n1933 VDD.t663 8.10567
R22122 VDD.n10863 VDD.t3012 8.10567
R22123 VDD.n1932 VDD.t2094 8.10567
R22124 VDD.n5612 VDD.t4623 8.10567
R22125 VDD.n5612 VDD.t825 8.10567
R22126 VDD.n5609 VDD.t4287 8.10567
R22127 VDD.n5609 VDD.t4599 8.10567
R22128 VDD.n5608 VDD.t2757 8.10567
R22129 VDD.n5608 VDD.t3079 8.10567
R22130 VDD.n10846 VDD.t4271 8.10567
R22131 VDD.n10846 VDD.t4575 8.10567
R22132 VDD.n10847 VDD.t3895 8.10567
R22133 VDD.n10847 VDD.t4239 8.10567
R22134 VDD.n10851 VDD.t954 8.10567
R22135 VDD.n10851 VDD.t812 8.10567
R22136 VDD.n5612 VDD.t2150 8.10567
R22137 VDD.n5612 VDD.t4447 8.10567
R22138 VDD.n5609 VDD.t1757 8.10567
R22139 VDD.n5609 VDD.t4121 8.10567
R22140 VDD.n5608 VDD.t4323 8.10567
R22141 VDD.n5608 VDD.t2572 8.10567
R22142 VDD.n10846 VDD.t1742 8.10567
R22143 VDD.n10846 VDD.t4099 8.10567
R22144 VDD.n10847 VDD.t1372 8.10567
R22145 VDD.n10847 VDD.t3708 8.10567
R22146 VDD.n10851 VDD.t4143 8.10567
R22147 VDD.n10851 VDD.t3319 8.10567
R22148 VDD.n5617 VDD.t2982 8.10567
R22149 VDD.n5548 VDD.t3905 8.10567
R22150 VDD.n5623 VDD.t3390 8.10567
R22151 VDD.n5547 VDD.t1511 8.10567
R22152 VDD.n5596 VDD.t4723 8.10567
R22153 VDD.n5550 VDD.t3364 8.10567
R22154 VDD.n5602 VDD.t2920 8.10567
R22155 VDD.n5549 VDD.t3746 8.10567
R22156 VDD.n5591 VDD.t2401 8.10567
R22157 VDD.n5591 VDD.t2747 8.10567
R22158 VDD.n5588 VDD.t1969 8.10567
R22159 VDD.n5588 VDD.t2373 8.10567
R22160 VDD.n5587 VDD.t4487 8.10567
R22161 VDD.n5587 VDD.t673 8.10567
R22162 VDD.n1972 VDD.t1942 8.10567
R22163 VDD.n1972 VDD.t2353 8.10567
R22164 VDD.n1973 VDD.t1548 8.10567
R22165 VDD.n1973 VDD.t1895 8.10567
R22166 VDD.n1977 VDD.t2178 8.10567
R22167 VDD.n1977 VDD.t2049 8.10567
R22168 VDD.n5591 VDD.t3987 8.10567
R22169 VDD.n5591 VDD.t2148 8.10567
R22170 VDD.n5588 VDD.t3623 8.10567
R22171 VDD.n5588 VDD.t1755 8.10567
R22172 VDD.n5587 VDD.t2010 8.10567
R22173 VDD.n5587 VDD.t4321 8.10567
R22174 VDD.n1972 VDD.t3608 8.10567
R22175 VDD.n1972 VDD.t1740 8.10567
R22176 VDD.n1973 VDD.t3283 8.10567
R22177 VDD.n1973 VDD.t1369 8.10567
R22178 VDD.n1977 VDD.t1179 8.10567
R22179 VDD.n1977 VDD.t4493 8.10567
R22180 VDD.n1954 VDD.t3677 8.10567
R22181 VDD.n1968 VDD.t1404 8.10567
R22182 VDD.n1955 VDD.t3675 8.10567
R22183 VDD.n1962 VDD.t3887 8.10567
R22184 VDD.n10809 VDD.t4435 8.10567
R22185 VDD.n10811 VDD.t3289 8.10567
R22186 VDD.n1953 VDD.t4431 8.10567
R22187 VDD.n1983 VDD.t4633 8.10567
R22188 VDD.n2116 VDD.t2567 8.10567
R22189 VDD.n2116 VDD.t3863 8.10567
R22190 VDD.n2113 VDD.t2133 8.10567
R22191 VDD.n2113 VDD.t3515 8.10567
R22192 VDD.n2112 VDD.t4665 8.10567
R22193 VDD.n2112 VDD.t1875 8.10567
R22194 VDD.n10825 VDD.t2113 8.10567
R22195 VDD.n10825 VDD.t3503 8.10567
R22196 VDD.n10824 VDD.t1713 8.10567
R22197 VDD.n10824 VDD.t3173 8.10567
R22198 VDD.n10821 VDD.t2468 8.10567
R22199 VDD.n10821 VDD.t1163 8.10567
R22200 VDD.n2116 VDD.t3463 8.10567
R22201 VDD.n2116 VDD.t647 8.10567
R22202 VDD.n2113 VDD.t3153 8.10567
R22203 VDD.n2113 VDD.t4455 8.10567
R22204 VDD.n2112 VDD.t1438 8.10567
R22205 VDD.n2112 VDD.t2932 8.10567
R22206 VDD.n10825 VDD.t3131 8.10567
R22207 VDD.n10825 VDD.t4429 8.10567
R22208 VDD.n10824 VDD.t2791 8.10567
R22209 VDD.n10824 VDD.t4073 8.10567
R22210 VDD.n10821 VDD.t1954 8.10567
R22211 VDD.n10821 VDD.t769 8.10567
R22212 VDD.n5554 VDD.t4209 8.10567
R22213 VDD.n5552 VDD.t1390 8.10567
R22214 VDD.n5581 VDD.t2377 8.10567
R22215 VDD.n5551 VDD.t3265 8.10567
R22216 VDD.n2102 VDD.t4105 8.10567
R22217 VDD.n8106 VDD.t861 8.10567
R22218 VDD.n2103 VDD.t671 8.10567
R22219 VDD.n8100 VDD.t2081 8.10567
R22220 VDD.n2099 VDD.t1929 8.10567
R22221 VDD.n2099 VDD.t3333 8.10567
R22222 VDD.n2096 VDD.t1563 8.10567
R22223 VDD.n2096 VDD.t3041 8.10567
R22224 VDD.n2095 VDD.t4151 8.10567
R22225 VDD.n2095 VDD.t1321 8.10567
R22226 VDD.n10788 VDD.t1542 8.10567
R22227 VDD.n10788 VDD.t3027 8.10567
R22228 VDD.n10789 VDD.t1176 8.10567
R22229 VDD.n10789 VDD.t2661 8.10567
R22230 VDD.n10793 VDD.t3203 8.10567
R22231 VDD.n10793 VDD.t1925 8.10567
R22232 VDD.n2099 VDD.t1793 8.10567
R22233 VDD.n2099 VDD.t3255 8.10567
R22234 VDD.n2096 VDD.t1432 8.10567
R22235 VDD.n2096 VDD.t2926 8.10567
R22236 VDD.n2095 VDD.t4027 8.10567
R22237 VDD.n2095 VDD.t1205 8.10567
R22238 VDD.n10788 VDD.t1421 8.10567
R22239 VDD.n10788 VDD.t2906 8.10567
R22240 VDD.n10789 VDD.t1080 8.10567
R22241 VDD.n10789 VDD.t2537 8.10567
R22242 VDD.n10793 VDD.t2741 8.10567
R22243 VDD.n10793 VDD.t1412 8.10567
R22244 VDD.n10799 VDD.t2739 8.10567
R22245 VDD.n2006 VDD.t2936 8.10567
R22246 VDD.n10805 VDD.t1000 8.10567
R22247 VDD.n2005 VDD.t3937 8.10567
R22248 VDD.n2036 VDD.t3422 8.10567
R22249 VDD.n2050 VDD.t3612 8.10567
R22250 VDD.n2037 VDD.t1710 8.10567
R22251 VDD.n2044 VDD.t4681 8.10567
R22252 VDD.n8128 VDD.t4257 8.10567
R22253 VDD.n8128 VDD.t1012 8.10567
R22254 VDD.n8125 VDD.t3901 8.10567
R22255 VDD.n8125 VDD.t632 8.10567
R22256 VDD.n8124 VDD.t2348 8.10567
R22257 VDD.n8124 VDD.t3249 8.10567
R22258 VDD.n2027 VDD.t3879 8.10567
R22259 VDD.n2027 VDD.t597 8.10567
R22260 VDD.n2028 VDD.t3511 8.10567
R22261 VDD.n2028 VDD.t4393 8.10567
R22262 VDD.n2032 VDD.t3037 8.10567
R22263 VDD.n2032 VDD.t3221 8.10567
R22264 VDD.n8128 VDD.t1259 8.10567
R22265 VDD.n8128 VDD.t2751 8.10567
R22266 VDD.n8125 VDD.t952 8.10567
R22267 VDD.n8125 VDD.t2379 8.10567
R22268 VDD.n8124 VDD.t3487 8.10567
R22269 VDD.n8124 VDD.t676 8.10567
R22270 VDD.n2027 VDD.t929 8.10567
R22271 VDD.n2027 VDD.t2359 8.10567
R22272 VDD.n2028 VDD.t4683 8.10567
R22273 VDD.n2028 VDD.t1897 8.10567
R22274 VDD.n2032 VDD.t3425 8.10567
R22275 VDD.n2032 VDD.t2225 8.10567
R22276 VDD.n2091 VDD.t3549 8.10567
R22277 VDD.n8118 VDD.t4449 8.10567
R22278 VDD.n2092 VDD.t4297 8.10567
R22279 VDD.n8112 VDD.t1493 8.10567
R22280 VDD.n8141 VDD.t1203 8.10567
R22281 VDD.n8139 VDD.t2146 8.10567
R22282 VDD.n2090 VDD.t1979 8.10567
R22283 VDD.n8133 VDD.t3366 8.10567
R22284 VDD.n8173 VDD.t754 8.10567
R22285 VDD.n8173 VDD.t2120 8.10567
R22286 VDD.n8188 VDD.t4517 8.10567
R22287 VDD.n8188 VDD.t1732 8.10567
R22288 VDD.n2078 VDD.t3019 8.10567
R22289 VDD.n2078 VDD.t4303 8.10567
R22290 VDD.n8222 VDD.t4503 8.10567
R22291 VDD.n8222 VDD.t1718 8.10567
R22292 VDD.n8229 VDD.t4173 8.10567
R22293 VDD.n8229 VDD.t1348 8.10567
R22294 VDD.n2064 VDD.t4183 8.10567
R22295 VDD.n2064 VDD.t3035 8.10567
R22296 VDD.n10768 VDD.t4615 8.10567
R22297 VDD.n2060 VDD.t669 8.10567
R22298 VDD.n2026 VDD.t3039 8.10567
R22299 VDD.n2056 VDD.t1730 8.10567
R22300 VDD.n2248 VDD.t3953 8.10567
R22301 VDD.n2250 VDD.t3586 8.10567
R22302 VDD.n7780 VDD.t1078 8.10567
R22303 VDD.n2272 VDD.t1090 8.10567
R22304 VDD.n7719 VDD.t2826 8.10567
R22305 VDD.n2282 VDD.t2451 8.10567
R22306 VDD.n2292 VDD.t2710 8.10567
R22307 VDD.n7825 VDD.t2051 8.10567
R22308 VDD.n7824 VDD.t1662 8.10567
R22309 VDD.n2240 VDD.t2329 8.10567
R22310 VDD.n7097 VDD.t3107 8.10567
R22311 VDD.n7093 VDD.t3963 8.10567
R22312 VDD.n7102 VDD.t1146 8.10567
R22313 VDD.n7090 VDD.t3969 8.10567
R22314 VDD.n7089 VDD.t3045 8.10567
R22315 VDD.n7109 VDD.t4699 8.10567
R22316 VDD.n2329 VDD.t1919 8.10567
R22317 VDD.n7115 VDD.t2424 8.10567
R22318 VDD.n2327 VDD.t3724 8.10567
R22319 VDD.n7120 VDD.t971 8.10567
R22320 VDD.n2324 VDD.t2246 8.10567
R22321 VDD.n2240 VDD.t4335 8.10567
R22322 VDD.n7097 VDD.t969 8.10567
R22323 VDD.n7093 VDD.t1830 8.10567
R22324 VDD.n7102 VDD.t3281 8.10567
R22325 VDD.n7090 VDD.t1838 8.10567
R22326 VDD.n7089 VDD.t900 8.10567
R22327 VDD.n7109 VDD.t2700 8.10567
R22328 VDD.n2329 VDD.t4003 8.10567
R22329 VDD.n7115 VDD.t4391 8.10567
R22330 VDD.n2327 VDD.t1613 8.10567
R22331 VDD.n7120 VDD.t3081 8.10567
R22332 VDD.n2324 VDD.t4283 8.10567
R22333 VDD.n2400 VDD.t2872 8.10567
R22334 VDD.n2398 VDD.t4425 8.10567
R22335 VDD.n2397 VDD.t4091 8.10567
R22336 VDD.n7129 VDD.t991 8.10567
R22337 VDD.n7128 VDD.t4741 8.10567
R22338 VDD.n7126 VDD.t2292 8.10567
R22339 VDD.n2400 VDD.t2525 8.10567
R22340 VDD.n2398 VDD.t4113 8.10567
R22341 VDD.n2397 VDD.t3732 8.10567
R22342 VDD.n7129 VDD.t582 8.10567
R22343 VDD.n7128 VDD.t4395 8.10567
R22344 VDD.n7126 VDD.t1888 8.10567
R22345 VDD.n2343 VDD.t4309 8.10567
R22346 VDD.n2345 VDD.t2016 8.10567
R22347 VDD.n2346 VDD.t1639 8.10567
R22348 VDD.n7045 VDD.t3929 8.10567
R22349 VDD.n7046 VDD.t3561 8.10567
R22350 VDD.n2343 VDD.t3979 8.10567
R22351 VDD.n2345 VDD.t1655 8.10567
R22352 VDD.n2346 VDD.t1283 8.10567
R22353 VDD.n7045 VDD.t3576 8.10567
R22354 VDD.n7046 VDD.t3267 8.10567
R22355 VDD.n7071 VDD.t1813 8.10567
R22356 VDD.n7069 VDD.t2830 8.10567
R22357 VDD.n7076 VDD.t4141 8.10567
R22358 VDD.n7066 VDD.t2838 8.10567
R22359 VDD.n2335 VDD.t1734 8.10567
R22360 VDD.n7083 VDD.t3519 8.10567
R22361 VDD.n7063 VDD.t731 8.10567
R22362 VDD.n2336 VDD.t1131 8.10567
R22363 VDD.n2337 VDD.t2615 8.10567
R22364 VDD.n2338 VDD.t3907 8.10567
R22365 VDD.n2339 VDD.t1021 8.10567
R22366 VDD.n2340 VDD.t1060 8.10567
R22367 VDD.n6655 VDD.t694 8.10567
R22368 VDD.n6658 VDD.t1434 8.10567
R22369 VDD.n6653 VDD.t2928 8.10567
R22370 VDD.n6663 VDD.t3755 8.10567
R22371 VDD.n6650 VDD.t1313 8.10567
R22372 VDD.n6649 VDD.t830 8.10567
R22373 VDD.n6648 VDD.t3191 8.10567
R22374 VDD.n6647 VDD.t4491 8.10567
R22375 VDD.n6676 VDD.t4011 8.10567
R22376 VDD.n6645 VDD.t1109 8.10567
R22377 VDD.n6681 VDD.t2575 8.10567
R22378 VDD.n6642 VDD.t3414 8.10567
R22379 VDD.n7071 VDD.t1832 8.10567
R22380 VDD.n7069 VDD.t2846 8.10567
R22381 VDD.n7076 VDD.t4157 8.10567
R22382 VDD.n7066 VDD.t2852 8.10567
R22383 VDD.n2335 VDD.t1749 8.10567
R22384 VDD.n7083 VDD.t3531 8.10567
R22385 VDD.n7063 VDD.t757 8.10567
R22386 VDD.n2336 VDD.t1144 8.10567
R22387 VDD.n2337 VDD.t2631 8.10567
R22388 VDD.n2338 VDD.t3925 8.10567
R22389 VDD.n2339 VDD.t1033 8.10567
R22390 VDD.n2340 VDD.t1070 8.10567
R22391 VDD.n6655 VDD.t715 8.10567
R22392 VDD.n6658 VDD.t1466 8.10567
R22393 VDD.n6653 VDD.t2956 8.10567
R22394 VDD.n6663 VDD.t3775 8.10567
R22395 VDD.n6650 VDD.t1326 8.10567
R22396 VDD.n6649 VDD.t857 8.10567
R22397 VDD.n6648 VDD.t3211 8.10567
R22398 VDD.n6647 VDD.t4505 8.10567
R22399 VDD.n6676 VDD.t4025 8.10567
R22400 VDD.n6645 VDD.t1120 8.10567
R22401 VDD.n6681 VDD.t2593 8.10567
R22402 VDD.n6642 VDD.t3429 8.10567
R22403 VDD.n6711 VDD.t2870 8.10567
R22404 VDD.n6709 VDD.t4423 8.10567
R22405 VDD.n6708 VDD.t4089 8.10567
R22406 VDD.n6704 VDD.t989 8.10567
R22407 VDD.n6703 VDD.t4739 8.10567
R22408 VDD.n6701 VDD.t2290 8.10567
R22409 VDD.n6711 VDD.t704 8.10567
R22410 VDD.n6709 VDD.t2444 8.10567
R22411 VDD.n6708 VDD.t1998 8.10567
R22412 VDD.n6704 VDD.t3109 8.10567
R22413 VDD.n6703 VDD.t2779 8.10567
R22414 VDD.n6701 VDD.t4329 8.10567
R22415 VDD.n6697 VDD.t4307 8.10567
R22416 VDD.n6695 VDD.t2014 8.10567
R22417 VDD.n6694 VDD.t1637 8.10567
R22418 VDD.n6690 VDD.t3927 8.10567
R22419 VDD.n6689 VDD.t3559 8.10567
R22420 VDD.n6687 VDD.t1058 8.10567
R22421 VDD.n6697 VDD.t2256 8.10567
R22422 VDD.n6695 VDD.t4111 8.10567
R22423 VDD.n6694 VDD.t3730 8.10567
R22424 VDD.n6690 VDD.t1815 8.10567
R22425 VDD.n6689 VDD.t1448 8.10567
R22426 VDD.n6687 VDD.t3187 8.10567
R22427 VDD.n6640 VDD.t1072 8.10567
R22428 VDD.n6638 VDD.t2805 8.10567
R22429 VDD.n6637 VDD.t2434 8.10567
R22430 VDD.n5434 VDD.t2688 8.10567
R22431 VDD.n5435 VDD.t2273 8.10567
R22432 VDD.n5437 VDD.t1952 8.10567
R22433 VDD.n6640 VDD.t3205 8.10567
R22434 VDD.n6638 VDD.t612 8.10567
R22435 VDD.n6637 VDD.t4409 8.10567
R22436 VDD.n5434 VDD.t4677 8.10567
R22437 VDD.n5435 VDD.t4315 8.10567
R22438 VDD.n5437 VDD.t4049 8.10567
R22439 VDD.n5442 VDD.t885 8.10567
R22440 VDD.n5440 VDD.t2603 8.10567
R22441 VDD.n5439 VDD.t2164 8.10567
R22442 VDD.n6629 VDD.t2215 8.10567
R22443 VDD.n6628 VDD.t1805 8.10567
R22444 VDD.n6626 VDD.t3684 8.10567
R22445 VDD.n5442 VDD.t3021 8.10567
R22446 VDD.n5440 VDD.t4557 8.10567
R22447 VDD.n5439 VDD.t4241 8.10567
R22448 VDD.n6629 VDD.t4273 8.10567
R22449 VDD.n6628 VDD.t3919 8.10567
R22450 VDD.n6626 VDD.t1592 8.10567
R22451 VDD.n2374 VDD.t3269 8.10567
R22452 VDD.n2373 VDD.t4553 8.10567
R22453 VDD.n7030 VDD.t1311 8.10567
R22454 VDD.n2372 VDD.t3149 8.10567
R22455 VDD.n2371 VDD.t2649 8.10567
R22456 VDD.n7037 VDD.t722 8.10567
R22457 VDD.n6716 VDD.t2101 8.10567
R22458 VDD.n6715 VDD.t1551 8.10567
R22459 VDD.n6722 VDD.t2944 8.10567
R22460 VDD.n2407 VDD.t4243 8.10567
R22461 VDD.n2406 VDD.t1004 8.10567
R22462 VDD.n2385 VDD.t3588 8.10567
R22463 VDD.n6872 VDD.t4473 8.10567
R22464 VDD.n2391 VDD.t1687 8.10567
R22465 VDD.n6867 VDD.t4477 8.10567
R22466 VDD.n2392 VDD.t3513 8.10567
R22467 VDD.n6862 VDD.t1092 8.10567
R22468 VDD.n2393 VDD.t2554 8.10567
R22469 VDD.n2394 VDD.t2974 8.10567
R22470 VDD.n6854 VDD.t4267 8.10567
R22471 VDD.n2395 VDD.t1460 8.10567
R22472 VDD.n2404 VDD.t2842 8.10567
R22473 VDD.n5236 VDD.t2761 8.10567
R22474 VDD.n5234 VDD.t4057 8.10567
R22475 VDD.n5241 VDD.t807 8.10567
R22476 VDD.n5231 VDD.t2635 8.10567
R22477 VDD.n5230 VDD.t2039 8.10567
R22478 VDD.n5248 VDD.t4339 8.10567
R22479 VDD.n5227 VDD.t1531 8.10567
R22480 VDD.n5254 VDD.t1044 8.10567
R22481 VDD.n5225 VDD.t2388 8.10567
R22482 VDD.n5259 VDD.t3690 8.10567
R22483 VDD.n5222 VDD.t4571 8.10567
R22484 VDD.n5236 VDD.t4725 8.10567
R22485 VDD.n5234 VDD.t1946 8.10567
R22486 VDD.n5241 VDD.t2954 8.10567
R22487 VDD.n5231 VDD.t4577 8.10567
R22488 VDD.n5230 VDD.t4101 8.10567
R22489 VDD.n5248 VDD.t2277 8.10567
R22490 VDD.n5227 VDD.t3621 8.10567
R22491 VDD.n5254 VDD.t3161 8.10567
R22492 VDD.n5225 VDD.t4363 8.10567
R22493 VDD.n5259 VDD.t1574 8.10567
R22494 VDD.n5222 VDD.t2591 8.10567
R22495 VDD.n5474 VDD.t4417 8.10567
R22496 VDD.n5475 VDD.t565 8.10567
R22497 VDD.n5476 VDD.t1985 8.10567
R22498 VDD.n5477 VDD.t4299 8.10567
R22499 VDD.n5478 VDD.t3787 8.10567
R22500 VDD.n5479 VDD.t1933 8.10567
R22501 VDD.n5480 VDD.t2333 8.10567
R22502 VDD.n5482 VDD.t3229 8.10567
R22503 VDD.n5483 VDD.t4087 8.10567
R22504 VDD.n5484 VDD.t1271 8.10567
R22505 VDD.n5485 VDD.t4095 8.10567
R22506 VDD.n5486 VDD.t4371 8.10567
R22507 VDD.n5474 VDD.t3337 8.10567
R22508 VDD.n5475 VDD.t3659 8.10567
R22509 VDD.n5476 VDD.t914 8.10567
R22510 VDD.n5477 VDD.t3263 8.10567
R22511 VDD.n5478 VDD.t2785 8.10567
R22512 VDD.n5479 VDD.t872 8.10567
R22513 VDD.n5480 VDD.t1166 8.10567
R22514 VDD.n5482 VDD.t2085 8.10567
R22515 VDD.n5483 VDD.t3051 8.10567
R22516 VDD.n5484 VDD.t4349 8.10567
R22517 VDD.n5485 VDD.t3055 8.10567
R22518 VDD.n5486 VDD.t3309 8.10567
R22519 VDD.n5446 VDD.t627 8.10567
R22520 VDD.n5391 VDD.t2037 8.10567
R22521 VDD.n5451 VDD.t3017 8.10567
R22522 VDD.n5388 VDD.t4667 8.10567
R22523 VDD.n5387 VDD.t4175 8.10567
R22524 VDD.n5458 VDD.t2386 8.10567
R22525 VDD.n5384 VDD.t3688 8.10567
R22526 VDD.n5464 VDD.t4541 8.10567
R22527 VDD.n5382 VDD.t4437 8.10567
R22528 VDD.n5469 VDD.t1650 8.10567
R22529 VDD.n5379 VDD.t3993 8.10567
R22530 VDD.n5446 VDD.t3700 8.10567
R22531 VDD.n5391 VDD.t948 8.10567
R22532 VDD.n5451 VDD.t1809 8.10567
R22533 VDD.n5388 VDD.t3582 8.10567
R22534 VDD.n5387 VDD.t3121 8.10567
R22535 VDD.n5458 VDD.t1192 8.10567
R22536 VDD.n5384 VDD.t2677 8.10567
R22537 VDD.n5464 VDD.t3499 8.10567
R22538 VDD.n5382 VDD.t3358 8.10567
R22539 VDD.n5469 VDD.t4713 8.10567
R22540 VDD.n5379 VDD.t2970 8.10567
R22541 VDD.n6264 VDD.t2478 8.10567
R22542 VDD.n6263 VDD.t2047 8.10567
R22543 VDD.n6366 VDD.t2341 8.10567
R22544 VDD.n6365 VDD.t1908 8.10567
R22545 VDD.n6363 VDD.t1621 8.10567
R22546 VDD.n6264 VDD.t3388 8.10567
R22547 VDD.n6263 VDD.t3089 8.10567
R22548 VDD.n6366 VDD.t3303 8.10567
R22549 VDD.n6365 VDD.t3000 8.10567
R22550 VDD.n6363 VDD.t2706 8.10567
R22551 VDD.n5937 VDD.t4689 8.10567
R22552 VDD.n5939 VDD.t2211 8.10567
R22553 VDD.n5940 VDD.t1801 8.10567
R22554 VDD.n5945 VDD.t1854 8.10567
R22555 VDD.n5946 VDD.t1483 8.10567
R22556 VDD.n5948 VDD.t3380 8.10567
R22557 VDD.n5937 VDD.t1498 8.10567
R22558 VDD.n5939 VDD.t3237 8.10567
R22559 VDD.n5940 VDD.t2896 8.10567
R22560 VDD.n5945 VDD.t2950 8.10567
R22561 VDD.n5946 VDD.t2583 8.10567
R22562 VDD.n5948 VDD.t4351 8.10567
R22563 VDD.n5271 VDD.t2457 8.10567
R22564 VDD.n6590 VDD.t3757 8.10567
R22565 VDD.n5272 VDD.t4647 8.10567
R22566 VDD.n6585 VDD.t2281 8.10567
R22567 VDD.n5273 VDD.t1699 8.10567
R22568 VDD.n6580 VDD.t4051 8.10567
R22569 VDD.n5924 VDD.t1242 8.10567
R22570 VDD.n5928 VDD.t2170 8.10567
R22571 VDD.n5923 VDD.t2027 8.10567
R22572 VDD.n5933 VDD.t3412 8.10567
R22573 VDD.n5922 VDD.t1527 8.10567
R22574 VDD.n6234 VDD.t3899 8.10567
R22575 VDD.n6232 VDD.t1114 8.10567
R22576 VDD.n6239 VDD.t2035 8.10567
R22577 VDD.n6229 VDD.t3769 8.10567
R22578 VDD.n6228 VDD.t3291 8.10567
R22579 VDD.n6246 VDD.t1388 8.10567
R22580 VDD.n6225 VDD.t2864 8.10567
R22581 VDD.n6252 VDD.t3663 8.10567
R22582 VDD.n6223 VDD.t3539 8.10567
R22583 VDD.n6257 VDD.t773 8.10567
R22584 VDD.n6220 VDD.t3141 8.10567
R22585 VDD.n6219 VDD.t733 8.10567
R22586 VDD.n6215 VDD.t1689 8.10567
R22587 VDD.n6270 VDD.t3533 8.10567
R22588 VDD.n6213 VDD.t3861 8.10567
R22589 VDD.n6275 VDD.t1083 8.10567
R22590 VDD.n6210 VDD.t3410 8.10567
R22591 VDD.n6209 VDD.t2962 8.10567
R22592 VDD.n6282 VDD.t1037 8.10567
R22593 VDD.n6206 VDD.t1346 8.10567
R22594 VDD.n6288 VDD.t2308 8.10567
R22595 VDD.n6204 VDD.t3227 8.10567
R22596 VDD.n6293 VDD.t4519 8.10567
R22597 VDD.n6201 VDD.t3233 8.10567
R22598 VDD.n6200 VDD.t3491 8.10567
R22599 VDD.n6234 VDD.t3917 8.10567
R22600 VDD.n6232 VDD.t1124 8.10567
R22601 VDD.n6239 VDD.t2055 8.10567
R22602 VDD.n6229 VDD.t3785 8.10567
R22603 VDD.n6228 VDD.t3299 8.10567
R22604 VDD.n6246 VDD.t1400 8.10567
R22605 VDD.n6225 VDD.t2876 8.10567
R22606 VDD.n6252 VDD.t3682 8.10567
R22607 VDD.n6223 VDD.t3551 8.10567
R22608 VDD.n6257 VDD.t784 8.10567
R22609 VDD.n6220 VDD.t3155 8.10567
R22610 VDD.n6219 VDD.t759 8.10567
R22611 VDD.n6215 VDD.t1705 8.10567
R22612 VDD.n6270 VDD.t3543 8.10567
R22613 VDD.n6213 VDD.t3875 8.10567
R22614 VDD.n6275 VDD.t1101 8.10567
R22615 VDD.n6210 VDD.t3431 8.10567
R22616 VDD.n6209 VDD.t2978 8.10567
R22617 VDD.n6282 VDD.t1062 8.10567
R22618 VDD.n6206 VDD.t1362 8.10567
R22619 VDD.n6288 VDD.t2331 8.10567
R22620 VDD.n6204 VDD.t3241 8.10567
R22621 VDD.n6293 VDD.t4525 8.10567
R22622 VDD.n6201 VDD.t3247 8.10567
R22623 VDD.n6200 VDD.t3501 8.10567
R22624 VDD.n6302 VDD.t1006 8.10567
R22625 VDD.n6303 VDD.t585 8.10567
R22626 VDD.n6307 VDD.t895 8.10567
R22627 VDD.n6306 VDD.t4651 8.10567
R22628 VDD.n5985 VDD.t786 8.10567
R22629 VDD.n5986 VDD.t4535 8.10567
R22630 VDD.n6315 VDD.t4593 8.10567
R22631 VDD.n6316 VDD.t4261 8.10567
R22632 VDD.n6318 VDD.t1948 8.10567
R22633 VDD.n5952 VDD.t2008 8.10567
R22634 VDD.n5921 VDD.t2415 8.10567
R22635 VDD.n5957 VDD.t3720 8.10567
R22636 VDD.n5920 VDD.t1862 8.10567
R22637 VDD.n5919 VDD.t1335 8.10567
R22638 VDD.n5964 VDD.t3673 8.10567
R22639 VDD.n5918 VDD.t4023 8.10567
R22640 VDD.n5970 VDD.t761 8.10567
R22641 VDD.n5917 VDD.t1635 8.10567
R22642 VDD.n5975 VDD.t3097 8.10567
R22643 VDD.n5916 VDD.t1644 8.10567
R22644 VDD.n6180 VDD.t1064 8.10567
R22645 VDD.n6182 VDD.t2795 8.10567
R22646 VDD.n6183 VDD.t2417 8.10567
R22647 VDD.n6187 VDD.t3404 8.10567
R22648 VDD.n6188 VDD.t3091 8.10567
R22649 VDD.n6192 VDD.t4419 8.10567
R22650 VDD.n6193 VDD.t4085 8.10567
R22651 VDD.n6197 VDD.t2205 8.10567
R22652 VDD.n6198 VDD.t1791 8.10567
R22653 VDD.n6381 VDD.t4719 8.10567
R22654 VDD.n5319 VDD.t927 8.10567
R22655 VDD.n6386 VDD.t2339 8.10567
R22656 VDD.n5316 VDD.t4569 8.10567
R22657 VDD.n5315 VDD.t4093 8.10567
R22658 VDD.n6393 VDD.t2269 8.10567
R22659 VDD.n5995 VDD.t2659 8.10567
R22660 VDD.n5999 VDD.t3481 8.10567
R22661 VDD.n5992 VDD.t4361 8.10567
R22662 VDD.n6004 VDD.t1565 8.10567
R22663 VDD.n5989 VDD.t4367 8.10567
R22664 VDD.n6010 VDD.t4671 8.10567
R22665 VDD.n6381 VDD.t2716 8.10567
R22666 VDD.n5319 VDD.t3043 8.10567
R22667 VDD.n6386 VDD.t4341 8.10567
R22668 VDD.n5316 VDD.t2589 8.10567
R22669 VDD.n5315 VDD.t1977 8.10567
R22670 VDD.n6393 VDD.t4295 8.10567
R22671 VDD.n5995 VDD.t4613 8.10567
R22672 VDD.n5999 VDD.t1342 8.10567
R22673 VDD.n5992 VDD.t2327 8.10567
R22674 VDD.n6004 VDD.t3639 8.10567
R22675 VDD.n5989 VDD.t2337 8.10567
R22676 VDD.n6010 VDD.t2665 8.10567
R22677 VDD.n5335 VDD.t959 8.10567
R22678 VDD.n5333 VDD.t2392 8.10567
R22679 VDD.n5340 VDD.t3277 8.10567
R22680 VDD.n5330 VDD.t820 8.10567
R22681 VDD.n5329 VDD.t4441 8.10567
R22682 VDD.n5347 VDD.t2694 8.10567
R22683 VDD.n5326 VDD.t3997 8.10567
R22684 VDD.n5353 VDD.t713 8.10567
R22685 VDD.n5324 VDD.t4731 8.10567
R22686 VDD.n5358 VDD.t1959 8.10567
R22687 VDD.n5321 VDD.t4277 8.10567
R22688 VDD.n5335 VDD.t3077 8.10567
R22689 VDD.n5333 VDD.t4369 8.10567
R22690 VDD.n5340 VDD.t1122 8.10567
R22691 VDD.n5330 VDD.t2960 8.10567
R22692 VDD.n5329 VDD.t2430 8.10567
R22693 VDD.n5347 VDD.t4661 8.10567
R22694 VDD.n5326 VDD.t1871 8.10567
R22695 VDD.n5353 VDD.t2860 8.10567
R22696 VDD.n5324 VDD.t2735 8.10567
R22697 VDD.n5358 VDD.t4039 8.10567
R22698 VDD.n5321 VDD.t2199 8.10567
R22699 VDD.n5363 VDD.t2556 8.10567
R22700 VDD.n5365 VDD.t4137 8.10567
R22701 VDD.n5366 VDD.t3763 8.10567
R22702 VDD.n5370 VDD.t615 8.10567
R22703 VDD.n5371 VDD.t4421 8.10567
R22704 VDD.n5373 VDD.t1921 8.10567
R22705 VDD.n5363 VDD.t3471 8.10567
R22706 VDD.n5365 VDD.t973 8.10567
R22707 VDD.n5366 VDD.t4733 8.10567
R22708 VDD.n5370 VDD.t1608 8.10567
R22709 VDD.n5371 VDD.t1248 8.10567
R22710 VDD.n5373 VDD.t3008 8.10567
R22711 VDD.n6377 VDD.t4005 8.10567
R22712 VDD.n6375 VDD.t1671 8.10567
R22713 VDD.n6374 VDD.t1305 8.10567
R22714 VDD.n6216 VDD.t3596 8.10567
R22715 VDD.n6217 VDD.t3287 8.10567
R22716 VDD.n6377 VDD.t838 8.10567
R22717 VDD.n6375 VDD.t2771 8.10567
R22718 VDD.n6374 VDD.t2394 8.10567
R22719 VDD.n6216 VDD.t4545 8.10567
R22720 VDD.n6217 VDD.t4237 8.10567
R22721 VDD.n5298 VDD.t1107 8.10567
R22722 VDD.n6409 VDD.t1416 8.10567
R22723 VDD.n5300 VDD.t2898 8.10567
R22724 VDD.n6404 VDD.t1002 8.10567
R22725 VDD.n5301 VDD.t4595 8.10567
R22726 VDD.n6399 VDD.t2858 8.10567
R22727 VDD.n6159 VDD.t3169 8.10567
R22728 VDD.n6163 VDD.t4013 8.10567
R22729 VDD.n6158 VDD.t767 8.10567
R22730 VDD.n6168 VDD.t2131 8.10567
R22731 VDD.n6018 VDD.t775 8.10567
R22732 VDD.n5287 VDD.t1450 8.10567
R22733 VDD.n5286 VDD.t2946 8.10567
R22734 VDD.n6567 VDD.t3767 8.10567
R22735 VDD.n5285 VDD.t1317 8.10567
R22736 VDD.n5284 VDD.t849 8.10567
R22737 VDD.n6574 VDD.t3209 8.10567
R22738 VDD.n6026 VDD.t4499 8.10567
R22739 VDD.n6025 VDD.t1230 8.10567
R22740 VDD.n6032 VDD.t1118 8.10567
R22741 VDD.n6023 VDD.t2581 8.10567
R22742 VDD.n6022 VDD.t645 8.10567
R22743 VDD.n8065 VDD.t1096 8.10567
R22744 VDD.n2159 VDD.t3751 8.10567
R22745 VDD.n2161 VDD.t2168 8.10567
R22746 VDD.n8014 VDD.t909 8.10567
R22747 VDD.n7861 VDD.t1380 8.10567
R22748 VDD.n7862 VDD.t3965 8.10567
R22749 VDD.n7911 VDD.t2304 8.10567
R22750 VDD.n7852 VDD.t2692 8.10567
R22751 VDD.n2207 VDD.t1213 8.10567
R22752 VDD.n2214 VDD.t4385 8.10567
R22753 VDD.n2232 VDD.t1991 8.10567
R22754 VDD.n2221 VDD.t3378 8.10567
R22755 VDD.n7987 VDD.t3791 8.10567
R22756 VDD.n2191 VDD.t1017 8.10567
R22757 VDD.n2195 VDD.t2470 8.10567
R22758 VDD.n2194 VDD.t3645 8.10567
R22759 VDD.n2198 VDD.t3686 8.10567
R22760 VDD.n2200 VDD.t3349 8.10567
R22761 VDD.n7961 VDD.t4131 8.10567
R22762 VDD.n6599 VDD.t1303 8.10567
R22763 VDD.n2205 VDD.t2783 8.10567
R22764 VDD.n2217 VDD.t4479 8.10567
R22765 VDD.n2213 VDD.t1691 8.10567
R22766 VDD.n2211 VDD.t3061 8.10567
R22767 VDD.n2220 VDD.t4359 8.10567
R22768 VDD.n7988 VDD.t1105 8.10567
R22769 VDD.n2190 VDD.t2006 8.10567
R22770 VDD.n2196 VDD.t3400 8.10567
R22771 VDD.n2197 VDD.t1428 8.10567
R22772 VDD.n7974 VDD.t2438 8.10567
R22773 VDD.n2201 VDD.t1010 8.10567
R22774 VDD.n7967 VDD.t1881 8.10567
R22775 VDD.n7962 VDD.t2755 8.10567
R22776 VDD.n6602 VDD.t2265 8.10567
R22777 VDD.n6598 VDD.t3989 8.10567
R22778 VDD.n6597 VDD.t3479 8.10567
R22779 VDD.n6609 VDD.t1602 8.10567
R22780 VDD.n6596 VDD.t3071 8.10567
R22781 VDD.n6615 VDD.t2563 8.10567
R22782 VDD.n6595 VDD.t3753 8.10567
R22783 VDD.n6620 VDD.t998 8.10567
R22784 VDD.n6594 VDD.t1864 8.10567
R22785 VDD.n2358 VDD.t2803 8.10567
R22786 VDD.n2359 VDD.t2432 8.10567
R22787 VDD.n2364 VDD.t2686 8.10567
R22788 VDD.n2363 VDD.t2271 8.10567
R22789 VDD.n2361 VDD.t1950 8.10567
R22790 VDD.n2358 VDD.t2449 8.10567
R22791 VDD.n2359 VDD.t2004 8.10567
R22792 VDD.n2364 VDD.t2306 8.10567
R22793 VDD.n2363 VDD.t1879 8.10567
R22794 VDD.n2361 VDD.t1594 8.10567
R22795 VDD.n7140 VDD.t882 8.10567
R22796 VDD.n7138 VDD.t2601 8.10567
R22797 VDD.n7137 VDD.t2162 8.10567
R22798 VDD.n2315 VDD.t2213 8.10567
R22799 VDD.n2314 VDD.t1803 8.10567
R22800 VDD.n7140 VDD.t4663 8.10567
R22801 VDD.n7138 VDD.t2176 8.10567
R22802 VDD.n7137 VDD.t1773 8.10567
R22803 VDD.n2315 VDD.t1826 8.10567
R22804 VDD.n2314 VDD.t1462 8.10567
R22805 VDD.n5407 VDD.t2459 8.10567
R22806 VDD.n5405 VDD.t3761 8.10567
R22807 VDD.n5412 VDD.t4649 8.10567
R22808 VDD.n5402 VDD.t2283 8.10567
R22809 VDD.n5401 VDD.t1701 8.10567
R22810 VDD.n5419 VDD.t4053 8.10567
R22811 VDD.n5398 VDD.t1244 8.10567
R22812 VDD.n5425 VDD.t765 8.10567
R22813 VDD.n5396 VDD.t2029 8.10567
R22814 VDD.n5430 VDD.t3416 8.10567
R22815 VDD.n5393 VDD.t4301 8.10567
R22816 VDD.n5407 VDD.t1257 8.10567
R22817 VDD.n5405 VDD.t2749 8.10567
R22818 VDD.n5412 VDD.t3574 8.10567
R22819 VDD.n5402 VDD.t1133 8.10567
R22820 VDD.n5401 VDD.t600 8.10567
R22821 VDD.n5419 VDD.t3025 8.10567
R22822 VDD.n5398 VDD.t4317 8.10567
R22823 VDD.n5425 VDD.t3807 8.10567
R22824 VDD.n5396 VDD.t946 8.10567
R22825 VDD.n5430 VDD.t2369 8.10567
R22826 VDD.n5393 VDD.t3261 8.10567
R22827 VDD.n2297 VDD.t1975 8.10567
R22828 VDD.n2298 VDD.t2832 8.10567
R22829 VDD.n2299 VDD.t3643 8.10567
R22830 VDD.n2300 VDD.t907 8.10567
R22831 VDD.n2301 VDD.t3651 8.10567
R22832 VDD.n2302 VDD.t2759 8.10567
R22833 VDD.n2303 VDD.t4397 8.10567
R22834 VDD.n2304 VDD.t1619 8.10567
R22835 VDD.n2306 VDD.t2073 8.10567
R22836 VDD.n2307 VDD.t3453 8.10567
R22837 VDD.n2308 VDD.t640 8.10567
R22838 VDD.n2309 VDD.t1914 8.10567
R22839 VDD.n2297 VDD.t912 8.10567
R22840 VDD.n2298 VDD.t1633 8.10567
R22841 VDD.n2299 VDD.t2641 8.10567
R22842 VDD.n2300 VDD.t3949 8.10567
R22843 VDD.n2301 VDD.t2653 8.10567
R22844 VDD.n2302 VDD.t1546 8.10567
R22845 VDD.n2303 VDD.t3331 8.10567
R22846 VDD.n2304 VDD.t4687 8.10567
R22847 VDD.n2306 VDD.t985 8.10567
R22848 VDD.n2307 VDD.t2411 8.10567
R22849 VDD.n2308 VDD.t3712 8.10567
R22850 VDD.n2309 VDD.t847 8.10567
R22851 VDD.n2295 VDD.t2625 8.10567
R22852 VDD.n2294 VDD.t2191 8.10567
R22853 VDD.n7838 VDD.t2242 8.10567
R22854 VDD.n7839 VDD.t1834 8.10567
R22855 VDD.n7841 VDD.t3710 8.10567
R22856 VDD.n7844 VDD.t4465 8.10567
R22857 VDD.n2208 VDD.t1201 8.10567
R22858 VDD.n7177 VDD.t2312 8.10567
R22859 VDD.n7945 VDD.t1394 8.10567
R22860 VDD.n7944 VDD.t3985 8.10567
R22861 VDD.n7854 VDD.t2335 8.10567
R22862 VDD.n2148 VDD.t1116 8.10567
R22863 VDD.n8050 VDD.t3779 8.10567
R22864 VDD.n8049 VDD.t2195 8.10567
R22865 VDD.n2149 VDD.t924 8.10567
R22866 VDD.n2174 VDD.t2801 8.10567
R22867 VDD.n2171 VDD.t4107 8.10567
R22868 VDD.n2179 VDD.t1185 8.10567
R22869 VDD.n2170 VDD.t2669 8.10567
R22870 VDD.n2169 VDD.t3493 8.10567
R22871 VDD.n2186 VDD.t4373 8.10567
R22872 VDD.n2168 VDD.t1584 8.10567
R22873 VDD.n8002 VDD.t3833 8.10567
R22874 VDD.n2167 VDD.t4727 8.10567
R22875 VDD.n8007 VDD.t3376 8.10567
R22876 VDD.n2166 VDD.t4275 8.10567
R22877 VDD.n2389 VDD.t2894 8.10567
R22878 VDD.n2387 VDD.t4457 8.10567
R22879 VDD.n2386 VDD.t4119 8.10567
R22880 VDD.n7830 VDD.t1008 8.10567
R22881 VDD.n7829 VDD.t592 8.10567
R22882 VDD.n9133 VDD.t3517 8.10567
R22883 VDD.n9128 VDD.t3321 8.10567
R22884 VDD.n9133 VDD.t2998 8.10567
R22885 VDD.n9128 VDD.t2793 8.10567
R22886 VDD.n9127 VDD.t3313 8.10567
R22887 VDD.n9127 VDD.t3133 8.10567
R22888 VDD.n9125 VDD.t719 8.10567
R22889 VDD.n9125 VDD.t4645 8.10567
R22890 VDD.n9137 VDD.t2629 8.10567
R22891 VDD.n9137 VDD.t2398 8.10567
R22892 VDD.n9135 VDD.t2976 8.10567
R22893 VDD.n9135 VDD.t2765 8.10567
R22894 VDD.n9140 VDD.t2546 8.10567
R22895 VDD.n9085 VDD.t4041 8.10567
R22896 VDD.n9146 VDD.t3897 8.10567
R22897 VDD.n9084 VDD.t3671 8.10567
R22898 VDD.n9081 VDD.t2141 8.10567
R22899 VDD.n9081 VDD.t3694 8.10567
R22900 VDD.n9078 VDD.t2579 8.10567
R22901 VDD.n9078 VDD.t4061 8.10567
R22902 VDD.n9077 VDD.t3165 8.10567
R22903 VDD.n9077 VDD.t4655 8.10567
R22904 VDD.n9174 VDD.t2599 8.10567
R22905 VDD.n9174 VDD.t4075 8.10567
R22906 VDD.n9173 VDD.t2968 8.10567
R22907 VDD.n9173 VDD.t4433 8.10567
R22908 VDD.n9170 VDD.t4463 8.10567
R22909 VDD.n9170 VDD.t1866 8.10567
R22910 VDD.n9081 VDD.t2535 8.10567
R22911 VDD.n9081 VDD.t2253 8.10567
R22912 VDD.n9078 VDD.t2880 8.10567
R22913 VDD.n9078 VDD.t2673 8.10567
R22914 VDD.n9077 VDD.t3439 8.10567
R22915 VDD.n9077 VDD.t3259 8.10567
R22916 VDD.n9174 VDD.t2902 8.10567
R22917 VDD.n9174 VDD.t2684 8.10567
R22918 VDD.n9173 VDD.t3253 8.10567
R22919 VDD.n9173 VDD.t3053 8.10567
R22920 VDD.n9170 VDD.t602 8.10567
R22921 VDD.n9170 VDD.t4539 8.10567
R22922 VDD.n8471 VDD.t3101 8.10567
R22923 VDD.n9163 VDD.t4567 8.10567
R22924 VDD.n8485 VDD.t4459 8.10567
R22925 VDD.n8484 VDD.t4255 8.10567
R22926 VDD.n8580 VDD.t4059 8.10567
R22927 VDD.n8760 VDD.t3839 8.10567
R22928 VDD.n8581 VDD.t4515 8.10567
R22929 VDD.n8754 VDD.t3859 8.10567
R22930 VDD.n8577 VDD.t4281 8.10567
R22931 VDD.n8577 VDD.t1194 8.10567
R22932 VDD.n8574 VDD.t4617 8.10567
R22933 VDD.n8574 VDD.t1537 8.10567
R22934 VDD.n8573 VDD.t1094 8.10567
R22935 VDD.n8573 VDD.t2207 8.10567
R22936 VDD.n8567 VDD.t4643 8.10567
R22937 VDD.n8567 VDD.t1561 8.10567
R22938 VDD.n8566 VDD.t897 8.10567
R22939 VDD.n8566 VDD.t1963 8.10567
R22940 VDD.n8563 VDD.t2548 8.10567
R22941 VDD.n8563 VDD.t3557 8.10567
R22942 VDD.n8577 VDD.t2702 8.10567
R22943 VDD.n8577 VDD.t1407 8.10567
R22944 VDD.n8574 VDD.t3047 8.10567
R22945 VDD.n8574 VDD.t1761 8.10567
R22946 VDD.n8573 VDD.t3594 8.10567
R22947 VDD.n8573 VDD.t2489 8.10567
R22948 VDD.n8567 VDD.t3065 8.10567
R22949 VDD.n8567 VDD.t1777 8.10567
R22950 VDD.n8566 VDD.t3382 8.10567
R22951 VDD.n8566 VDD.t2201 8.10567
R22952 VDD.n8563 VDD.t809 8.10567
R22953 VDD.n8563 VDD.t3781 8.10567
R22954 VDD.n8548 VDD.t2250 8.10567
R22955 VDD.n8556 VDD.t2020 8.10567
R22956 VDD.n8549 VDD.t2811 8.10567
R22957 VDD.n8550 VDD.t2057 8.10567
R22958 VDD.n8830 VDD.t2868 8.10567
R22959 VDD.n8811 VDD.t2107 8.10567
R22960 VDD.n8544 VDD.t1031 8.10567
R22961 VDD.n8543 VDD.t2129 8.10567
R22962 VDD.n8795 VDD.t2463 8.10567
R22963 VDD.n8795 VDD.t3163 8.10567
R22964 VDD.n8792 VDD.t2820 8.10567
R22965 VDD.n8792 VDD.t3475 8.10567
R22966 VDD.n8791 VDD.t3360 8.10567
R22967 VDD.n8791 VDD.t4083 8.10567
R22968 VDD.n8785 VDD.t2836 8.10567
R22969 VDD.n8785 VDD.t3495 8.10567
R22970 VDD.n8784 VDD.t3185 8.10567
R22971 VDD.n8784 VDD.t3853 8.10567
R22972 VDD.n8781 VDD.t4707 8.10567
R22973 VDD.n8781 VDD.t1264 8.10567
R22974 VDD.n8795 VDD.t3235 8.10567
R22975 VDD.n8795 VDD.t1488 8.10567
R22976 VDD.n8792 VDD.t3537 8.10567
R22977 VDD.n8792 VDD.t1856 8.10567
R22978 VDD.n8791 VDD.t4169 8.10567
R22979 VDD.n8791 VDD.t2577 8.10567
R22980 VDD.n8785 VDD.t3547 8.10567
R22981 VDD.n8785 VDD.t1877 8.10567
R22982 VDD.n8784 VDD.t3935 8.10567
R22983 VDD.n8784 VDD.t2316 8.10567
R22984 VDD.n8781 VDD.t1332 8.10567
R22985 VDD.n8781 VDD.t3865 8.10567
R22986 VDD.n8800 VDD.t4583 8.10567
R22987 VDD.n8770 VDD.t3933 8.10567
R22988 VDD.n8531 VDD.t2940 8.10567
R22989 VDD.n8766 VDD.t3957 8.10567
R22990 VDD.n8517 VDD.t2519 8.10567
R22991 VDD.n8886 VDD.t3445 8.10567
R22992 VDD.n8772 VDD.t2436 8.10567
R22993 VDD.n8771 VDD.t3469 8.10567
R22994 VDD.n8849 VDD.t2552 8.10567
R22995 VDD.n8849 VDD.t3649 8.10567
R22996 VDD.n8853 VDD.t2900 8.10567
R22997 VDD.n8853 VDD.t4031 8.10567
R22998 VDD.n8854 VDD.t3459 8.10567
R22999 VDD.n8854 VDD.t4611 8.10567
R23000 VDD.n8862 VDD.t2912 8.10567
R23001 VDD.n8862 VDD.t4045 8.10567
R23002 VDD.n8863 VDD.t3275 8.10567
R23003 VDD.n8863 VDD.t4387 8.10567
R23004 VDD.n8867 VDD.t629 8.10567
R23005 VDD.n8867 VDD.t1817 8.10567
R23006 VDD.n8849 VDD.t1014 8.10567
R23007 VDD.n8849 VDD.t2098 8.10567
R23008 VDD.n8853 VDD.t1330 8.10567
R23009 VDD.n8853 VDD.t2531 8.10567
R23010 VDD.n8854 VDD.t1971 8.10567
R23011 VDD.n8854 VDD.t3129 8.10567
R23012 VDD.n8862 VDD.t1351 8.10567
R23013 VDD.n8862 VDD.t2550 8.10567
R23014 VDD.n8863 VDD.t1724 8.10567
R23015 VDD.n8863 VDD.t2918 8.10567
R23016 VDD.n8867 VDD.t3347 8.10567
R23017 VDD.n8867 VDD.t4415 8.10567
R23018 VDD.n8873 VDD.t576 8.10567
R23019 VDD.n8843 VDD.t1590 8.10567
R23020 VDD.n8521 VDD.t4691 8.10567
R23021 VDD.n8839 VDD.t1617 8.10567
R23022 VDD.n8506 VDD.t2466 8.10567
R23023 VDD.n8942 VDD.t1675 8.10567
R23024 VDD.n8845 VDD.t595 8.10567
R23025 VDD.n8844 VDD.t2209 8.10567
R23026 VDD.n8926 VDD.t4249 8.10567
R23027 VDD.n8926 VDD.t1250 8.10567
R23028 VDD.n8923 VDD.t4555 8.10567
R23029 VDD.n8923 VDD.t1606 8.10567
R23030 VDD.n8922 VDD.t1054 8.10567
R23031 VDD.n8922 VDD.t2267 8.10567
R23032 VDD.n8916 VDD.t4579 8.10567
R23033 VDD.n8916 VDD.t1625 8.10567
R23034 VDD.n8915 VDD.t841 8.10567
R23035 VDD.n8915 VDD.t2018 8.10567
R23036 VDD.n8912 VDD.t2503 8.10567
R23037 VDD.n8912 VDD.t3610 8.10567
R23038 VDD.n8926 VDD.t2854 8.10567
R23039 VDD.n8926 VDD.t3867 8.10567
R23040 VDD.n8923 VDD.t3183 8.10567
R23041 VDD.n8923 VDD.t4235 8.10567
R23042 VDD.n8922 VDD.t3744 8.10567
R23043 VDD.n8922 VDD.t666 8.10567
R23044 VDD.n8916 VDD.t3197 8.10567
R23045 VDD.n8916 VDD.t4247 8.10567
R23046 VDD.n8915 VDD.t3529 8.10567
R23047 VDD.n8915 VDD.t4589 8.10567
R23048 VDD.n8912 VDD.t978 8.10567
R23049 VDD.n8912 VDD.t2063 8.10567
R23050 VDD.n8931 VDD.t4225 8.10567
R23051 VDD.n8901 VDD.t3525 8.10567
R23052 VDD.n8512 VDD.t2527 8.10567
R23053 VDD.n8897 VDD.t4017 8.10567
R23054 VDD.n8498 VDD.t4289 8.10567
R23055 VDD.n9017 VDD.t4081 8.10567
R23056 VDD.n8903 VDD.t2623 8.10567
R23057 VDD.n8902 VDD.t4109 8.10567
R23058 VDD.n8976 VDD.t2078 8.10567
R23059 VDD.n8976 VDD.t1823 8.10567
R23060 VDD.n8980 VDD.t2501 8.10567
R23061 VDD.n8980 VDD.t2221 8.10567
R23062 VDD.n8981 VDD.t3099 8.10567
R23063 VDD.n8981 VDD.t2892 8.10567
R23064 VDD.n8989 VDD.t2515 8.10567
R23065 VDD.n8989 VDD.t2237 8.10567
R23066 VDD.n8990 VDD.t2882 8.10567
R23067 VDD.n8990 VDD.t2675 8.10567
R23068 VDD.n8994 VDD.t4383 8.10567
R23069 VDD.n8994 VDD.t4201 8.10567
R23070 VDD.n8976 VDD.t2948 8.10567
R23071 VDD.n8976 VDD.t2731 8.10567
R23072 VDD.n8980 VDD.t3271 8.10567
R23073 VDD.n8980 VDD.t3069 8.10567
R23074 VDD.n8981 VDD.t3831 8.10567
R23075 VDD.n8981 VDD.t3615 8.10567
R23076 VDD.n8989 VDD.t3279 8.10567
R23077 VDD.n8989 VDD.t3083 8.10567
R23078 VDD.n8990 VDD.t3604 8.10567
R23079 VDD.n8990 VDD.t3406 8.10567
R23080 VDD.n8994 VDD.t1041 8.10567
R23081 VDD.n8994 VDD.t835 8.10567
R23082 VDD.n8970 VDD.t2558 8.10567
R23083 VDD.n8952 VDD.t2287 8.10567
R23084 VDD.n8502 VDD.t706 8.10567
R23085 VDD.n8948 VDD.t2324 8.10567
R23086 VDD.n8489 VDD.t3023 8.10567
R23087 VDD.n9039 VDD.t4485 8.10567
R23088 VDD.n8972 VDD.t4365 8.10567
R23089 VDD.n8971 VDD.t4177 8.10567
R23090 VDD.n9060 VDD.t2154 8.10567
R23091 VDD.n9060 VDD.t1916 8.10567
R23092 VDD.n9057 VDD.t2585 8.10567
R23093 VDD.n9057 VDD.t2351 8.10567
R23094 VDD.n9056 VDD.t3175 8.10567
R23095 VDD.n9056 VDD.t2988 8.10567
R23096 VDD.n9050 VDD.t2607 8.10567
R23097 VDD.n9050 VDD.t2371 8.10567
R23098 VDD.n9049 VDD.t2980 8.10567
R23099 VDD.n9049 VDD.t2767 8.10567
R23100 VDD.n9046 VDD.t4467 8.10567
R23101 VDD.n9046 VDD.t4269 8.10567
R23102 VDD.n9060 VDD.t2446 8.10567
R23103 VDD.n9060 VDD.t2159 8.10567
R23104 VDD.n9057 VDD.t2807 8.10567
R23105 VDD.n9057 VDD.t2587 8.10567
R23106 VDD.n9056 VDD.t3335 8.10567
R23107 VDD.n9056 VDD.t3177 8.10567
R23108 VDD.n9050 VDD.t2822 8.10567
R23109 VDD.n9050 VDD.t2609 8.10567
R23110 VDD.n9049 VDD.t3171 8.10567
R23111 VDD.n9049 VDD.t2984 8.10567
R23112 VDD.n9046 VDD.t4693 8.10567
R23113 VDD.n9046 VDD.t4471 8.10567
R23114 VDD.n9028 VDD.t559 8.10567
R23115 VDD.n9027 VDD.t2188 8.10567
R23116 VDD.n8494 VDD.t2060 8.10567
R23117 VDD.n9023 VDD.t1795 8.10567
R23118 VDD.n9152 VDD.t679 8.10567
R23119 VDD.n9074 VDD.t2301 8.10567
R23120 VDD.n8474 VDD.t2126 8.10567
R23121 VDD.n9070 VDD.t1892 8.10567
R23122 VDD.n185 VDD.t4603 8.10567
R23123 VDD.n187 VDD.t2043 8.10567
R23124 VDD.n125 VDD.t4629 8.10567
R23125 VDD.n171 VDD.t4405 8.10567
R23126 VDD.n9117 VDD.t621 8.10567
R23127 VDD.n9098 VDD.t2227 8.10567
R23128 VDD.n9091 VDD.t2087 8.10567
R23129 VDD.n9092 VDD.t1836 8.10567
R23130 VDD.n1155 VDD.t3606 8.10567
R23131 VDD.t3606 VDD.n1139 8.10567
R23132 VDD.t4263 VDD.n1153 8.10567
R23133 VDD.n1154 VDD.t4263 8.10567
R23134 VDD.t3195 VDD.n1151 8.10567
R23135 VDD.n1152 VDD.t3195 8.10567
R23136 VDD.t3301 VDD.n1149 8.10567
R23137 VDD.n1150 VDD.t3301 8.10567
R23138 VDD.t2157 VDD.n1147 8.10567
R23139 VDD.n1148 VDD.t2157 8.10567
R23140 VDD.t2320 VDD.n1145 8.10567
R23141 VDD.n1146 VDD.t2320 8.10567
R23142 VDD.n1723 VDD.t1139 8.10567
R23143 VDD.t1139 VDD.n1722 8.10567
R23144 VDD.n1725 VDD.t1456 8.10567
R23145 VDD.t1456 VDD.n1724 8.10567
R23146 VDD.n1727 VDD.t4501 8.10567
R23147 VDD.t4501 VDD.n1726 8.10567
R23148 VDD.n1729 VDD.t4635 8.10567
R23149 VDD.t4635 VDD.n1728 8.10567
R23150 VDD.n1731 VDD.t3535 8.10567
R23151 VDD.t3535 VDD.n1730 8.10567
R23152 VDD.n1155 VDD.t750 8.10567
R23153 VDD.t750 VDD.n1139 8.10567
R23154 VDD.n1153 VDD.t3913 8.10567
R23155 VDD.n1154 VDD.t3913 8.10567
R23156 VDD.n1151 VDD.t2874 8.10567
R23157 VDD.n1152 VDD.t2874 8.10567
R23158 VDD.n1149 VDD.t3004 8.10567
R23159 VDD.n1150 VDD.t3004 8.10567
R23160 VDD.n1147 VDD.t1771 8.10567
R23161 VDD.n1148 VDD.t1771 8.10567
R23162 VDD.n1145 VDD.t1912 8.10567
R23163 VDD.n1146 VDD.t1912 8.10567
R23164 VDD.n1723 VDD.t815 8.10567
R23165 VDD.n1722 VDD.t815 8.10567
R23166 VDD.n1725 VDD.t1129 8.10567
R23167 VDD.n1724 VDD.t1129 8.10567
R23168 VDD.n1727 VDD.t4191 8.10567
R23169 VDD.n1726 VDD.t4191 8.10567
R23170 VDD.n1729 VDD.t4293 8.10567
R23171 VDD.n1728 VDD.t4293 8.10567
R23172 VDD.n1731 VDD.t3243 8.10567
R23173 VDD.n1730 VDD.t3243 8.10567
R23174 VDD.n928 VDD.t688 8.10567
R23175 VDD.t688 VDD.n699 8.10567
R23176 VDD.n930 VDD.t3738 8.10567
R23177 VDD.t3738 VDD.n929 8.10567
R23178 VDD.n932 VDD.t4071 8.10567
R23179 VDD.t4071 VDD.n931 8.10567
R23180 VDD.n934 VDD.t3961 8.10567
R23181 VDD.t3961 VDD.n933 8.10567
R23182 VDD.n936 VDD.t4079 8.10567
R23183 VDD.t4079 VDD.n935 8.10567
R23184 VDD.n1048 VDD.t3033 8.10567
R23185 VDD.t3033 VDD.n1047 8.10567
R23186 VDD.n1050 VDD.t3143 8.10567
R23187 VDD.t3143 VDD.n1049 8.10567
R23188 VDD.n1052 VDD.t1961 8.10567
R23189 VDD.t1961 VDD.n1051 8.10567
R23190 VDD.n1054 VDD.t4035 8.10567
R23191 VDD.t4035 VDD.n1053 8.10567
R23192 VDD.n1056 VDD.t2992 8.10567
R23193 VDD.t2992 VDD.n1055 8.10567
R23194 VDD.n1058 VDD.t1344 8.10567
R23195 VDD.t1344 VDD.n1057 8.10567
R23196 VDD.n928 VDD.t4231 8.10567
R23197 VDD.t4231 VDD.n699 8.10567
R23198 VDD.n930 VDD.t3159 8.10567
R23199 VDD.n929 VDD.t3159 8.10567
R23200 VDD.n932 VDD.t3451 8.10567
R23201 VDD.n931 VDD.t3451 8.10567
R23202 VDD.n934 VDD.t3327 8.10567
R23203 VDD.n933 VDD.t3327 8.10567
R23204 VDD.n936 VDD.t3455 8.10567
R23205 VDD.n935 VDD.t3455 8.10567
R23206 VDD.n1048 VDD.t2396 8.10567
R23207 VDD.n1047 VDD.t2396 8.10567
R23208 VDD.n1050 VDD.t2523 8.10567
R23209 VDD.n1049 VDD.t2523 8.10567
R23210 VDD.n1052 VDD.t1296 8.10567
R23211 VDD.n1051 VDD.t1296 8.10567
R23212 VDD.n1054 VDD.t3396 8.10567
R23213 VDD.n1053 VDD.t3396 8.10567
R23214 VDD.n1056 VDD.t2314 8.10567
R23215 VDD.n1055 VDD.t2314 8.10567
R23216 VDD.n1058 VDD.t741 8.10567
R23217 VDD.n1057 VDD.t741 8.10567
R23218 VDD.t2144 VDD.n1706 8.10567
R23219 VDD.n1707 VDD.t2144 8.10567
R23220 VDD.t1025 VDD.n1704 8.10567
R23221 VDD.n1705 VDD.t1025 8.10567
R23222 VDD.t1319 VDD.n1702 8.10567
R23223 VDD.n1703 VDD.t1319 8.10567
R23224 VDD.t1211 VDD.n1700 8.10567
R23225 VDD.n1701 VDD.t1211 8.10567
R23226 VDD.t1324 VDD.n1698 8.10567
R23227 VDD.n1699 VDD.t1324 8.10567
R23228 VDD.n886 VDD.t4379 8.10567
R23229 VDD.t4379 VDD.n885 8.10567
R23230 VDD.n888 VDD.t4497 8.10567
R23231 VDD.t4497 VDD.n887 8.10567
R23232 VDD.n890 VDD.t3420 8.10567
R23233 VDD.t3420 VDD.n889 8.10567
R23234 VDD.n892 VDD.t1279 8.10567
R23235 VDD.t1279 VDD.n891 8.10567
R23236 VDD.n894 VDD.t4345 8.10567
R23237 VDD.t4345 VDD.n893 8.10567
R23238 VDD.n896 VDD.t2888 8.10567
R23239 VDD.t2888 VDD.n895 8.10567
R23240 VDD.n1706 VDD.t1472 8.10567
R23241 VDD.n1707 VDD.t1472 8.10567
R23242 VDD.n1704 VDD.t4513 8.10567
R23243 VDD.n1705 VDD.t4513 8.10567
R23244 VDD.n1702 VDD.t709 8.10567
R23245 VDD.n1703 VDD.t709 8.10567
R23246 VDD.n1700 VDD.t4735 8.10567
R23247 VDD.n1701 VDD.t4735 8.10567
R23248 VDD.n1698 VDD.t711 8.10567
R23249 VDD.n1699 VDD.t711 8.10567
R23250 VDD.n886 VDD.t3765 8.10567
R23251 VDD.n885 VDD.t3765 8.10567
R23252 VDD.n888 VDD.t3885 8.10567
R23253 VDD.n887 VDD.t3885 8.10567
R23254 VDD.n890 VDD.t2850 8.10567
R23255 VDD.n889 VDD.t2850 8.10567
R23256 VDD.n892 VDD.t655 8.10567
R23257 VDD.n891 VDD.t655 8.10567
R23258 VDD.n894 VDD.t3704 8.10567
R23259 VDD.n893 VDD.t3704 8.10567
R23260 VDD.n896 VDD.t2193 8.10567
R23261 VDD.n895 VDD.t2193 8.10567
R23262 VDD.t4213 VDD.n1475 8.10567
R23263 VDD.n1476 VDD.t4213 8.10567
R23264 VDD.t3147 VDD.n1473 8.10567
R23265 VDD.n1474 VDD.t3147 8.10567
R23266 VDD.t3427 VDD.n1471 8.10567
R23267 VDD.n1472 VDD.t3427 8.10567
R23268 VDD.t3323 VDD.n1469 8.10567
R23269 VDD.n1470 VDD.t3323 8.10567
R23270 VDD.t3435 VDD.n1467 8.10567
R23271 VDD.n1468 VDD.t3435 8.10567
R23272 VDD.n1293 VDD.t2367 8.10567
R23273 VDD.t2367 VDD.n742 8.10567
R23274 VDD.n1295 VDD.t2507 8.10567
R23275 VDD.t2507 VDD.n1294 8.10567
R23276 VDD.n1297 VDD.t1277 8.10567
R23277 VDD.t1277 VDD.n1296 8.10567
R23278 VDD.n1299 VDD.t3362 8.10567
R23279 VDD.t3362 VDD.n1298 8.10567
R23280 VDD.n1301 VDD.t2275 8.10567
R23281 VDD.t2275 VDD.n1300 8.10567
R23282 VDD.n1303 VDD.t699 8.10567
R23283 VDD.t699 VDD.n1302 8.10567
R23284 VDD.n1475 VDD.t817 8.10567
R23285 VDD.n1476 VDD.t817 8.10567
R23286 VDD.n1473 VDD.t3855 8.10567
R23287 VDD.n1474 VDD.t3855 8.10567
R23288 VDD.n1471 VDD.t4199 8.10567
R23289 VDD.n1472 VDD.t4199 8.10567
R23290 VDD.n1469 VDD.t4065 8.10567
R23291 VDD.n1470 VDD.t4065 8.10567
R23292 VDD.n1467 VDD.t4207 8.10567
R23293 VDD.n1468 VDD.t4207 8.10567
R23294 VDD.n1293 VDD.t3137 8.10567
R23295 VDD.t3137 VDD.n742 8.10567
R23296 VDD.n1295 VDD.t3251 8.10567
R23297 VDD.n1294 VDD.t3251 8.10567
R23298 VDD.n1297 VDD.t2090 8.10567
R23299 VDD.n1296 VDD.t2090 8.10567
R23300 VDD.n1299 VDD.t4153 8.10567
R23301 VDD.n1298 VDD.t4153 8.10567
R23302 VDD.n1301 VDD.t3087 8.10567
R23303 VDD.n1300 VDD.t3087 8.10567
R23304 VDD.n1303 VDD.t1454 8.10567
R23305 VDD.n1302 VDD.t1454 8.10567
R23306 VDD.n1234 VDD.t1784 8.10567
R23307 VDD.t1784 VDD.n1219 8.10567
R23308 VDD.t3669 VDD.n1232 8.10567
R23309 VDD.n1233 VDD.t3669 8.10567
R23310 VDD.t2647 VDD.n1230 8.10567
R23311 VDD.n1231 VDD.t2647 8.10567
R23312 VDD.t2781 VDD.n1228 8.10567
R23313 VDD.n1229 VDD.t2781 8.10567
R23314 VDD.t1533 VDD.n1226 8.10567
R23315 VDD.n1227 VDD.t1533 8.10567
R23316 VDD.t1667 VDD.n1085 8.10567
R23317 VDD.n1225 VDD.t1667 8.10567
R23318 VDD.t4717 VDD.n1099 8.10567
R23319 VDD.n1100 VDD.t4717 8.10567
R23320 VDD.t922 VDD.n1097 8.10567
R23321 VDD.n1098 VDD.t922 8.10567
R23322 VDD.t3955 VDD.n1095 8.10567
R23323 VDD.n1096 VDD.t3955 8.10567
R23324 VDD.t4069 VDD.n813 8.10567
R23325 VDD.n1234 VDD.t4203 8.10567
R23326 VDD.t4203 VDD.n1219 8.10567
R23327 VDD.n1232 VDD.t2357 8.10567
R23328 VDD.n1233 VDD.t2357 8.10567
R23329 VDD.n1230 VDD.t1148 8.10567
R23330 VDD.n1231 VDD.t1148 8.10567
R23331 VDD.n1228 VDD.t1267 8.10567
R23332 VDD.n1229 VDD.t1267 8.10567
R23333 VDD.n1226 VDD.t4333 8.10567
R23334 VDD.n1227 VDD.t4333 8.10567
R23335 VDD.t4445 VDD.n1085 8.10567
R23336 VDD.n1225 VDD.t4445 8.10567
R23337 VDD.n1099 VDD.t3343 8.10567
R23338 VDD.n1100 VDD.t3343 8.10567
R23339 VDD.n1097 VDD.t3655 8.10567
R23340 VDD.n1098 VDD.t3655 8.10567
R23341 VDD.n1095 VDD.t2637 8.10567
R23342 VDD.n1096 VDD.t2637 8.10567
R23343 VDD.t2763 VDD.n813 8.10567
R23344 VDD.n1267 VDD.t2904 8.10567
R23345 VDD.t2904 VDD.n1251 8.10567
R23346 VDD.t660 VDD.n1265 8.10567
R23347 VDD.n1266 VDD.t660 8.10567
R23348 VDD.t3714 VDD.n1263 8.10567
R23349 VDD.n1264 VDD.t3714 8.10567
R23350 VDD.t3837 VDD.n1261 8.10567
R23351 VDD.n1262 VDD.t3837 8.10567
R23352 VDD.t2809 VDD.n1259 8.10567
R23353 VDD.n1260 VDD.t2809 8.10567
R23354 VDD.t2916 VDD.n1257 8.10567
R23355 VDD.n1258 VDD.t2916 8.10567
R23356 VDD.t1695 VDD.n1617 8.10567
R23357 VDD.n1618 VDD.t1695 8.10567
R23358 VDD.t2069 VDD.n1615 8.10567
R23359 VDD.n1616 VDD.t2069 8.10567
R23360 VDD.t957 VDD.n1613 8.10567
R23361 VDD.n1614 VDD.t957 8.10567
R23362 VDD.n1267 VDD.t1039 8.10567
R23363 VDD.t1039 VDD.n1251 8.10567
R23364 VDD.n1265 VDD.t3465 8.10567
R23365 VDD.n1266 VDD.t3465 8.10567
R23366 VDD.n1263 VDD.t2403 8.10567
R23367 VDD.n1264 VDD.t2403 8.10567
R23368 VDD.n1261 VDD.t2529 8.10567
R23369 VDD.n1262 VDD.t2529 8.10567
R23370 VDD.n1259 VDD.t1301 8.10567
R23371 VDD.n1260 VDD.t1301 8.10567
R23372 VDD.n1257 VDD.t1426 8.10567
R23373 VDD.n1258 VDD.t1426 8.10567
R23374 VDD.n1617 VDD.t4475 8.10567
R23375 VDD.n1618 VDD.t4475 8.10567
R23376 VDD.n1615 VDD.t652 8.10567
R23377 VDD.n1616 VDD.t652 8.10567
R23378 VDD.n1613 VDD.t3698 8.10567
R23379 VDD.n1614 VDD.t3698 8.10567
R23380 VDD.n1612 VDD.t1066 8.10567
R23381 VDD.n1612 VDD.t3835 8.10567
R23382 VDD.t2461 VDD.n1590 8.10567
R23383 VDD.n1591 VDD.t2461 8.10567
R23384 VDD.t1236 VDD.n1588 8.10567
R23385 VDD.n1589 VDD.t1236 8.10567
R23386 VDD.t1567 VDD.n1586 8.10567
R23387 VDD.n1587 VDD.t1567 8.10567
R23388 VDD.t1444 VDD.n1584 8.10567
R23389 VDD.n1585 VDD.t1444 8.10567
R23390 VDD.t1578 VDD.n1582 8.10567
R23391 VDD.n1583 VDD.t1578 8.10567
R23392 VDD.t4619 VDD.n1670 8.10567
R23393 VDD.n1671 VDD.t4619 8.10567
R23394 VDD.t4743 VDD.n1668 8.10567
R23395 VDD.n1669 VDD.t4743 8.10567
R23396 VDD.t3631 VDD.n1666 8.10567
R23397 VDD.n1667 VDD.t3631 8.10567
R23398 VDD.n1576 VDD.t2753 8.10567
R23399 VDD.t2753 VDD.n1575 8.10567
R23400 VDD.n1570 VDD.t573 8.10567
R23401 VDD.t573 VDD.n1569 8.10567
R23402 VDD.n1572 VDD.t3641 8.10567
R23403 VDD.t3641 VDD.n1571 8.10567
R23404 VDD.n1574 VDD.t3783 8.10567
R23405 VDD.t3783 VDD.n1573 8.10567
R23406 VDD.t2322 VDD.n1637 8.10567
R23407 VDD.n1638 VDD.t2322 8.10567
R23408 VDD.n1634 VDD.t2480 8.10567
R23409 VDD.t2480 VDD.n774 8.10567
R23410 VDD.n1631 VDD.t1255 8.10567
R23411 VDD.t1255 VDD.n777 8.10567
R23412 VDD.n1628 VDD.t1386 8.10567
R23413 VDD.t1386 VDD.n779 8.10567
R23414 VDD.n1568 VDD.t4427 8.10567
R23415 VDD.t4427 VDD.n1567 8.10567
R23416 VDD.t3408 VDD.n1641 8.10567
R23417 VDD.n1642 VDD.t3408 8.10567
R23418 VDD.n1133 VDD.t950 8.10567
R23419 VDD.t950 VDD.n1118 8.10567
R23420 VDD.t3625 VDD.n1131 8.10567
R23421 VDD.n1132 VDD.t3625 8.10567
R23422 VDD.t2605 VDD.n1129 8.10567
R23423 VDD.n1130 VDD.t2605 8.10567
R23424 VDD.t2724 VDD.n1127 8.10567
R23425 VDD.n1128 VDD.t2724 8.10567
R23426 VDD.t1496 VDD.n1125 8.10567
R23427 VDD.n1126 VDD.t1496 8.10567
R23428 VDD.t1629 VDD.n852 8.10567
R23429 VDD.n1124 VDD.t1629 8.10567
R23430 VDD.t4679 VDD.n872 8.10567
R23431 VDD.n873 VDD.t4679 8.10567
R23432 VDD.t877 VDD.n870 8.10567
R23433 VDD.n871 VDD.t877 8.10567
R23434 VDD.t3903 VDD.n868 8.10567
R23435 VDD.n869 VDD.t3903 8.10567
R23436 VDD.t4037 VDD.n866 8.10567
R23437 VDD.n867 VDD.t4037 8.10567
R23438 VDD.t2996 VDD.n728 8.10567
R23439 VDD.n865 VDD.t2996 8.10567
R23440 VDD.n1133 VDD.t2244 8.10567
R23441 VDD.t2244 VDD.n1118 8.10567
R23442 VDD.n1131 VDD.t3317 8.10567
R23443 VDD.n1132 VDD.t3317 8.10567
R23444 VDD.n1129 VDD.t2186 8.10567
R23445 VDD.n1130 VDD.t2186 8.10567
R23446 VDD.n1127 VDD.t2365 8.10567
R23447 VDD.n1128 VDD.t2365 8.10567
R23448 VDD.n1125 VDD.t1159 8.10567
R23449 VDD.n1126 VDD.t1159 8.10567
R23450 VDD.t1273 VDD.n852 8.10567
R23451 VDD.n1124 VDD.t1273 8.10567
R23452 VDD.n872 VDD.t4337 8.10567
R23453 VDD.n873 VDD.t4337 8.10567
R23454 VDD.n870 VDD.t4657 8.10567
R23455 VDD.n871 VDD.t4657 8.10567
R23456 VDD.n868 VDD.t3553 8.10567
R23457 VDD.n869 VDD.t3553 8.10567
R23458 VDD.n866 VDD.t3665 8.10567
R23459 VDD.n867 VDD.t3665 8.10567
R23460 VDD.t2645 VDD.n728 8.10567
R23461 VDD.n865 VDD.t2645 8.10567
R23462 VDD.n1204 VDD.t4179 8.10567
R23463 VDD.t4179 VDD.n1189 8.10567
R23464 VDD.t3722 VDD.n1202 8.10567
R23465 VDD.n1203 VDD.t3722 8.10567
R23466 VDD.t2696 VDD.n1200 8.10567
R23467 VDD.n1201 VDD.t2696 8.10567
R23468 VDD.t2818 VDD.n1198 8.10567
R23469 VDD.n1199 VDD.t2818 8.10567
R23470 VDD.t1598 VDD.n1196 8.10567
R23471 VDD.n1197 VDD.t1598 8.10567
R23472 VDD.t1716 VDD.n851 8.10567
R23473 VDD.n1195 VDD.t1716 8.10567
R23474 VDD.n1433 VDD.t590 8.10567
R23475 VDD.t590 VDD.n1432 8.10567
R23476 VDD.n1435 VDD.t981 8.10567
R23477 VDD.t981 VDD.n1434 8.10567
R23478 VDD.n1437 VDD.t4009 8.10567
R23479 VDD.t4009 VDD.n1436 8.10567
R23480 VDD.n1439 VDD.t4135 8.10567
R23481 VDD.t4135 VDD.n1438 8.10567
R23482 VDD.n1204 VDD.t1269 8.10567
R23483 VDD.t1269 VDD.n1189 8.10567
R23484 VDD.n1202 VDD.t3386 8.10567
R23485 VDD.n1203 VDD.t3386 8.10567
R23486 VDD.n1200 VDD.t2310 8.10567
R23487 VDD.n1201 VDD.t2310 8.10567
R23488 VDD.n1198 VDD.t2474 8.10567
R23489 VDD.n1199 VDD.t2474 8.10567
R23490 VDD.n1196 VDD.t1253 8.10567
R23491 VDD.n1197 VDD.t1253 8.10567
R23492 VDD.t1375 VDD.n851 8.10567
R23493 VDD.n1195 VDD.t1375 8.10567
R23494 VDD.n1433 VDD.t4413 8.10567
R23495 VDD.n1432 VDD.t4413 8.10567
R23496 VDD.n1435 VDD.t556 8.10567
R23497 VDD.n1434 VDD.t556 8.10567
R23498 VDD.n1437 VDD.t3633 8.10567
R23499 VDD.n1436 VDD.t3633 8.10567
R23500 VDD.n1439 VDD.t3773 8.10567
R23501 VDD.n1438 VDD.t3773 8.10567
R23502 VDD.t3073 VDD.n1440 8.10567
R23503 VDD.t3967 VDD.n801 8.10567
R23504 VDD.n802 VDD.t3967 8.10567
R23505 VDD.t2914 VDD.n799 8.10567
R23506 VDD.n800 VDD.t2914 8.10567
R23507 VDD.t3225 VDD.n797 8.10567
R23508 VDD.n798 VDD.t3225 8.10567
R23509 VDD.t3115 VDD.n795 8.10567
R23510 VDD.n796 VDD.t3115 8.10567
R23511 VDD.t3231 VDD.n793 8.10567
R23512 VDD.n794 VDD.t3231 8.10567
R23513 VDD.n1325 VDD.t2071 8.10567
R23514 VDD.t2071 VDD.n745 8.10567
R23515 VDD.n1327 VDD.t2197 8.10567
R23516 VDD.t2197 VDD.n1326 8.10567
R23517 VDD.n1329 VDD.t1068 8.10567
R23518 VDD.t1068 VDD.n1328 8.10567
R23519 VDD.n1331 VDD.t3179 8.10567
R23520 VDD.t3179 VDD.n1330 8.10567
R23521 VDD.n1333 VDD.t2000 8.10567
R23522 VDD.t2000 VDD.n1332 8.10567
R23523 VDD.n1335 VDD.t4607 8.10567
R23524 VDD.t4607 VDD.n1334 8.10567
R23525 VDD.n801 VDD.t4715 8.10567
R23526 VDD.n802 VDD.t4715 8.10567
R23527 VDD.n799 VDD.t3617 8.10567
R23528 VDD.n800 VDD.t3617 8.10567
R23529 VDD.n797 VDD.t3951 8.10567
R23530 VDD.n798 VDD.t3951 8.10567
R23531 VDD.n795 VDD.t3821 8.10567
R23532 VDD.n796 VDD.t3821 8.10567
R23533 VDD.n793 VDD.t3959 8.10567
R23534 VDD.n794 VDD.t3959 8.10567
R23535 VDD.n1325 VDD.t2908 8.10567
R23536 VDD.t2908 VDD.n745 8.10567
R23537 VDD.n1327 VDD.t3031 8.10567
R23538 VDD.n1326 VDD.t3031 8.10567
R23539 VDD.n1329 VDD.t1811 8.10567
R23540 VDD.n1328 VDD.t1811 8.10567
R23541 VDD.n1331 VDD.t3893 8.10567
R23542 VDD.n1330 VDD.t3893 8.10567
R23543 VDD.n1333 VDD.t2856 8.10567
R23544 VDD.n1332 VDD.t2856 8.10567
R23545 VDD.n1335 VDD.t1220 8.10567
R23546 VDD.n1334 VDD.t1220 8.10567
R23547 VDD.n1665 VDD.t1519 8.10567
R23548 VDD.t1519 VDD.n1664 8.10567
R23549 VDD.t4551 VDD.n1662 8.10567
R23550 VDD.n1663 VDD.t4551 8.10567
R23551 VDD.t2472 VDD.n838 8.10567
R23552 VDD.n839 VDD.t2472 8.10567
R23553 VDD.t1246 VDD.n836 8.10567
R23554 VDD.n837 VDD.t1246 8.10567
R23555 VDD.t1582 VDD.n834 8.10567
R23556 VDD.n835 VDD.t1582 8.10567
R23557 VDD.t1452 VDD.n832 8.10567
R23558 VDD.n833 VDD.t1452 8.10567
R23559 VDD.t1586 VDD.n830 8.10567
R23560 VDD.n831 VDD.t1586 8.10567
R23561 VDD.n1372 VDD.t4631 8.10567
R23562 VDD.t4631 VDD.n1371 8.10567
R23563 VDD.n1374 VDD.t562 8.10567
R23564 VDD.t562 VDD.n1373 8.10567
R23565 VDD.n1376 VDD.t3635 8.10567
R23566 VDD.t3635 VDD.n1375 8.10567
R23567 VDD.n1378 VDD.t1523 8.10567
R23568 VDD.t1523 VDD.n1377 8.10567
R23569 VDD.n1380 VDD.t4563 8.10567
R23570 VDD.t4563 VDD.n1379 8.10567
R23571 VDD.n1382 VDD.t3119 8.10567
R23572 VDD.t3119 VDD.n1381 8.10567
R23573 VDD.n838 VDD.t1720 8.10567
R23574 VDD.n839 VDD.t1720 8.10567
R23575 VDD.n836 VDD.t605 8.10567
R23576 VDD.n837 VDD.t605 8.10567
R23577 VDD.n834 VDD.t987 8.10567
R23578 VDD.n835 VDD.t987 8.10567
R23579 VDD.n832 VDD.t870 8.10567
R23580 VDD.n833 VDD.t870 8.10567
R23581 VDD.n830 VDD.t996 8.10567
R23582 VDD.n831 VDD.t996 8.10567
R23583 VDD.n1372 VDD.t4021 8.10567
R23584 VDD.n1371 VDD.t4021 8.10567
R23585 VDD.n1374 VDD.t4145 8.10567
R23586 VDD.n1373 VDD.t4145 8.10567
R23587 VDD.n1376 VDD.t3085 8.10567
R23588 VDD.n1375 VDD.t3085 8.10567
R23589 VDD.n1378 VDD.t939 8.10567
R23590 VDD.n1377 VDD.t939 8.10567
R23591 VDD.n1380 VDD.t3971 8.10567
R23592 VDD.n1379 VDD.t3971 8.10567
R23593 VDD.n1382 VDD.t2511 8.10567
R23594 VDD.n1381 VDD.t2511 8.10567
R23595 VDD.n8070 VDD.t1358 6.64567
R23596 VDD.n2126 VDD.t2840 6.64567
R23597 VDD.n2125 VDD.t941 6.64567
R23598 VDD.n2127 VDD.t2083 6.64567
R23599 VDD.n2141 VDD.t1023 6.64567
R23600 VDD.n2139 VDD.t2409 6.64567
R23601 VDD.n2138 VDD.t3325 6.64567
R23602 VDD.n2138 VDD.t2296 6.64567
R23603 VDD.n2134 VDD.t771 6.64567
R23604 VDD.n2134 VDD.t3869 6.64567
R23605 VDD.n2133 VDD.t3801 6.64567
R23606 VDD.n2133 VDD.t2844 6.64567
R23607 VDD.n2131 VDD.t1989 6.64567
R23608 VDD.n2131 VDD.t961 6.64567
R23609 VDD.n8085 VDD.t1275 6.64567
R23610 VDD.n8080 VDD.t2769 6.64567
R23611 VDD.n2122 VDD.t859 6.64567
R23612 VDD.n8066 VDD.t567 6.64567
R23613 VDD.n2156 VDD.t1910 6.64567
R23614 VDD.n2158 VDD.t1828 6.64567
R23615 VDD.n2165 VDD.t3473 6.64567
R23616 VDD.n8016 VDD.t2426 6.64567
R23617 VDD.n8013 VDD.t4685 6.64567
R23618 VDD.n6021 VDD.t4878 6.58663
R23619 VDD.n6094 VDD.t4954 6.58663
R23620 VDD.n6846 VDD.t269 6.58663
R23621 VDD.n6796 VDD.t177 6.58663
R23622 VDD.n7009 VDD.n7005 6.50088
R23623 VDD.n6958 VDD.n6957 6.50088
R23624 VDD.n6548 VDD.n6547 6.50088
R23625 VDD.n6501 VDD.n6497 6.50088
R23626 VDD.n6116 VDD.n6109 6.45575
R23627 VDD.n6073 VDD.n6066 6.45575
R23628 VDD.n6801 VDD.n6800 6.45575
R23629 VDD.n6752 VDD.n6746 6.45575
R23630 VDD.n1719 VDD.n709 6.24156
R23631 VDD.n1415 VDD.n874 6.24156
R23632 VDD.n1429 VDD.n1428 6.24156
R23633 VDD.n1354 VDD.n1084 6.24156
R23634 VDD.n1346 VDD.n1345 6.24156
R23635 VDD.n6153 VDD.n6152 5.95439
R23636 VDD.n6096 VDD.n6095 5.95439
R23637 VDD.n6847 VDD.n6844 5.95439
R23638 VDD.n6797 VDD.n6794 5.95439
R23639 VDD.n8643 VDD.n8642 5.76894
R23640 VDD.n8702 VDD.n8701 5.76894
R23641 VDD.n1812 VDD.n1811 5.76894
R23642 VDD.n1868 VDD.n1867 5.76894
R23643 VDD.n5516 VDD.n5515 5.76894
R23644 VDD.n1960 VDD.n1959 5.76894
R23645 VDD.n2042 VDD.n2041 5.76894
R23646 VDD.n8752 VDD.n8751 5.76894
R23647 VDD.n8895 VDD.n8894 5.76894
R23648 VDD.n9068 VDD.n9067 5.76894
R23649 VDD.n8642 VDD.n8641 5.33948
R23650 VDD.n8701 VDD.n8700 5.33948
R23651 VDD.n1811 VDD.n1810 5.33948
R23652 VDD.n1867 VDD.n1866 5.33948
R23653 VDD.n5515 VDD.n5514 5.33948
R23654 VDD.n1959 VDD.n1958 5.33948
R23655 VDD.n2041 VDD.n2040 5.33948
R23656 VDD.n8751 VDD.n8750 5.33948
R23657 VDD.n8894 VDD.n8893 5.33948
R23658 VDD.n9067 VDD.n9066 5.33948
R23659 VDD.n6153 VDD.t4858 5.31528
R23660 VDD.n6096 VDD.t4936 5.31528
R23661 VDD.n6844 VDD.t90 5.31528
R23662 VDD.n6794 VDD.t225 5.31528
R23663 VDD.n2130 VDD.t414 5.19255
R23664 VDD.n983 VDD.t454 5.17005
R23665 VDD.n1034 VDD.t463 5.17005
R23666 VDD.n1044 VDD.t449 5.17005
R23667 VDD.n1105 VDD.t369 5.17005
R23668 VDD.n1620 VDD.t375 5.17005
R23669 VDD.n1086 VDD.t373 5.17005
R23670 VDD.n1419 VDD.t447 5.17005
R23671 VDD.n853 VDD.t460 5.17005
R23672 VDD.n1677 VDD.t347 5.17005
R23673 VDD.n1683 VDD.t342 5.17005
R23674 VDD.n1689 VDD.t340 5.17005
R23675 VDD.n1696 VDD.t440 5.17005
R23676 VDD.n979 VDD.t431 5.1669
R23677 VDD.n1039 VDD.t450 5.1669
R23678 VDD.n735 VDD.t466 5.1669
R23679 VDD.n784 VDD.t376 5.1669
R23680 VDD.n1625 VDD.t348 5.1669
R23681 VDD.n1091 VDD.t4976 5.1669
R23682 VDD.n1424 VDD.t448 5.1669
R23683 VDD.n858 VDD.t441 5.1669
R23684 VDD.n1673 VDD.t357 5.1669
R23685 VDD.n1679 VDD.t345 5.1669
R23686 VDD.n1685 VDD.t492 5.1669
R23687 VDD.n1692 VDD.t451 5.1669
R23688 VDD.n7952 VDD.t106 5.12594
R23689 VDD.n6370 VDD.n5376 5.12014
R23690 VDD.n7133 VDD.n2317 5.12014
R23691 VDD.n8057 VDD.t206 5.09041
R23692 VDD.n8069 VDD.t1359 5.0505
R23693 VDD.t942 VDD.n2145 5.0505
R23694 VDD.n2144 VDD.t2084 5.0505
R23695 VDD.t2084 VDD.n2143 5.0505
R23696 VDD.n2128 VDD.t860 5.0505
R23697 VDD.n8084 VDD.t1276 5.0505
R23698 VDD.n6743 VDD.n6742 4.96877
R23699 VDD.n6070 VDD.n6069 4.96877
R23700 VDD.n6113 VDD.n6112 4.96877
R23701 VDD.n6737 VDD.n6736 4.96877
R23702 VDD.n2379 VDD.n2377 4.92758
R23703 VDD.n6962 VDD.n6960 4.92758
R23704 VDD.n5292 VDD.n5290 4.92758
R23705 VDD.n6507 VDD.n6505 4.92758
R23706 VDD.n6887 VDD.n6886 4.78594
R23707 VDD.n6906 VDD.n6905 4.78594
R23708 VDD.n6420 VDD.n6419 4.78594
R23709 VDD.n6457 VDD.n6456 4.78594
R23710 VDD.n6744 VDD.n6743 4.61712
R23711 VDD.n6756 VDD.n6755 4.61712
R23712 VDD.n6071 VDD.n6070 4.61712
R23713 VDD.n6061 VDD.n6060 4.61712
R23714 VDD.n6114 VDD.n6113 4.61712
R23715 VDD.n6104 VDD.n6103 4.61712
R23716 VDD.n6738 VDD.n6737 4.61712
R23717 VDD.n6805 VDD.n6804 4.61712
R23718 VDD.n61 VDD.n60 4.61205
R23719 VDD.n70 VDD.n69 4.61205
R23720 VDD.n150 VDD.n149 4.61205
R23721 VDD.n159 VDD.n158 4.61205
R23722 VDD.n5769 VDD.n5768 4.61205
R23723 VDD.n5760 VDD.n5759 4.61205
R23724 VDD.n5836 VDD.n5835 4.61205
R23725 VDD.n5827 VDD.n5826 4.61205
R23726 VDD.n5653 VDD.n5652 4.61205
R23727 VDD.n5644 VDD.n5643 4.61205
R23728 VDD.n5571 VDD.n5570 4.61205
R23729 VDD.n5562 VDD.n5561 4.61205
R23730 VDD.n8157 VDD.n8156 4.61205
R23731 VDD.n8148 VDD.n8147 4.61205
R23732 VDD.n9105 VDD.n9104 4.61205
R23733 VDD.n9114 VDD.n9113 4.61205
R23734 VDD.n8818 VDD.n8817 4.61205
R23735 VDD.n8827 VDD.n8826 4.61205
R23736 VDD.n8958 VDD.n8957 4.61205
R23737 VDD.n8967 VDD.n8966 4.61205
R23738 VDD.n6754 VDD.n6753 4.61078
R23739 VDD.n6997 VDD.n6994 4.61078
R23740 VDD.n6992 VDD.n6989 4.61078
R23741 VDD.n6987 VDD.n6984 4.61078
R23742 VDD.n6982 VDD.n6979 4.61078
R23743 VDD.n6900 VDD.n6897 4.61078
R23744 VDD.n6895 VDD.n6892 4.61078
R23745 VDD.n6890 VDD.n6887 4.61078
R23746 VDD.n6949 VDD.n6946 4.61078
R23747 VDD.n6944 VDD.n6941 4.61078
R23748 VDD.n6939 VDD.n6936 4.61078
R23749 VDD.n6934 VDD.n6931 4.61078
R23750 VDD.n6919 VDD.n6916 4.61078
R23751 VDD.n6914 VDD.n6911 4.61078
R23752 VDD.n6909 VDD.n6906 4.61078
R23753 VDD.n6525 VDD.n6524 4.61078
R23754 VDD.n6528 VDD.n6527 4.61078
R23755 VDD.n6531 VDD.n6530 4.61078
R23756 VDD.n6534 VDD.n6533 4.61078
R23757 VDD.n6433 VDD.n6430 4.61078
R23758 VDD.n6428 VDD.n6425 4.61078
R23759 VDD.n6423 VDD.n6420 4.61078
R23760 VDD.n6485 VDD.n6484 4.61078
R23761 VDD.n6488 VDD.n6487 4.61078
R23762 VDD.n6491 VDD.n6490 4.61078
R23763 VDD.n6494 VDD.n6493 4.61078
R23764 VDD.n6470 VDD.n6467 4.61078
R23765 VDD.n6465 VDD.n6462 4.61078
R23766 VDD.n6460 VDD.n6457 4.61078
R23767 VDD.n6065 VDD.n6062 4.61078
R23768 VDD.n6108 VDD.n6105 4.61078
R23769 VDD.n7893 VDD.n7892 4.61078
R23770 VDD.n7896 VDD.n7895 4.61078
R23771 VDD.n7899 VDD.n7898 4.61078
R23772 VDD.n7902 VDD.n7901 4.61078
R23773 VDD.n7905 VDD.n7904 4.61078
R23774 VDD.n7908 VDD.n7907 4.61078
R23775 VDD.n8045 VDD.n8042 4.61078
R23776 VDD.n8040 VDD.n8037 4.61078
R23777 VDD.n8035 VDD.n8032 4.61078
R23778 VDD.n8030 VDD.n8028 4.61078
R23779 VDD.n8026 VDD.n8023 4.61078
R23780 VDD.n8021 VDD.n8018 4.61078
R23781 VDD.n6803 VDD.n6802 4.61078
R23782 VDD.n7940 VDD.n7937 4.60951
R23783 VDD.n7941 VDD.n7940 4.60951
R23784 VDD.n7935 VDD.n7932 4.60951
R23785 VDD.n7936 VDD.n7935 4.60951
R23786 VDD.n7930 VDD.n7927 4.60951
R23787 VDD.n7931 VDD.n7930 4.60951
R23788 VDD.n7925 VDD.n7923 4.60951
R23789 VDD.n7926 VDD.n7925 4.60951
R23790 VDD.n7921 VDD.n7918 4.60951
R23791 VDD.n7922 VDD.n7921 4.60951
R23792 VDD.n7916 VDD.n7913 4.60951
R23793 VDD.n7917 VDD.n7916 4.60951
R23794 VDD.n6753 VDD.n6752 4.60825
R23795 VDD.n6998 VDD.n6997 4.60825
R23796 VDD.n6993 VDD.n6992 4.60825
R23797 VDD.n6988 VDD.n6987 4.60825
R23798 VDD.n6983 VDD.n6982 4.60825
R23799 VDD.n6901 VDD.n6900 4.60825
R23800 VDD.n6896 VDD.n6895 4.60825
R23801 VDD.n6891 VDD.n6890 4.60825
R23802 VDD.n6950 VDD.n6949 4.60825
R23803 VDD.n6945 VDD.n6944 4.60825
R23804 VDD.n6940 VDD.n6939 4.60825
R23805 VDD.n6935 VDD.n6934 4.60825
R23806 VDD.n6920 VDD.n6919 4.60825
R23807 VDD.n6915 VDD.n6914 4.60825
R23808 VDD.n6910 VDD.n6909 4.60825
R23809 VDD.n6524 VDD.n6523 4.60825
R23810 VDD.n6527 VDD.n6526 4.60825
R23811 VDD.n6530 VDD.n6529 4.60825
R23812 VDD.n6533 VDD.n6532 4.60825
R23813 VDD.n6434 VDD.n6433 4.60825
R23814 VDD.n6429 VDD.n6428 4.60825
R23815 VDD.n6424 VDD.n6423 4.60825
R23816 VDD.n6484 VDD.n6447 4.60825
R23817 VDD.n6487 VDD.n6486 4.60825
R23818 VDD.n6490 VDD.n6489 4.60825
R23819 VDD.n6493 VDD.n6492 4.60825
R23820 VDD.n6471 VDD.n6470 4.60825
R23821 VDD.n6466 VDD.n6465 4.60825
R23822 VDD.n6461 VDD.n6460 4.60825
R23823 VDD.n6066 VDD.n6065 4.60825
R23824 VDD.n6109 VDD.n6108 4.60825
R23825 VDD.n7892 VDD.n7891 4.60825
R23826 VDD.n7895 VDD.n7894 4.60825
R23827 VDD.n7898 VDD.n7897 4.60825
R23828 VDD.n7901 VDD.n7900 4.60825
R23829 VDD.n7904 VDD.n7903 4.60825
R23830 VDD.n7907 VDD.n7906 4.60825
R23831 VDD.n8046 VDD.n8045 4.60825
R23832 VDD.n8041 VDD.n8040 4.60825
R23833 VDD.n8036 VDD.n8035 4.60825
R23834 VDD.n8031 VDD.n8030 4.60825
R23835 VDD.n8027 VDD.n8026 4.60825
R23836 VDD.n8022 VDD.n8021 4.60825
R23837 VDD.n6802 VDD.n6801 4.60825
R23838 VDD.n6745 VDD.n6744 4.60191
R23839 VDD.n6757 VDD.n6756 4.60191
R23840 VDD.n6072 VDD.n6071 4.60191
R23841 VDD.n6060 VDD.n6041 4.60191
R23842 VDD.n6115 VDD.n6114 4.60191
R23843 VDD.n6103 VDD.n6101 4.60191
R23844 VDD.n6739 VDD.n6738 4.60191
R23845 VDD.n6806 VDD.n6805 4.60191
R23846 VDD.n8644 VDD.n8643 4.57315
R23847 VDD.n8703 VDD.n8702 4.57315
R23848 VDD.n1813 VDD.n1812 4.57315
R23849 VDD.n1869 VDD.n1868 4.57315
R23850 VDD.n5517 VDD.n5516 4.57315
R23851 VDD.n1961 VDD.n1960 4.57315
R23852 VDD.n2043 VDD.n2042 4.57315
R23853 VDD.n8753 VDD.n8752 4.57315
R23854 VDD.n8896 VDD.n8895 4.57315
R23855 VDD.n9069 VDD.n9068 4.57315
R23856 VDD.n8643 VDD.n8639 4.56231
R23857 VDD.n8702 VDD.n8698 4.56231
R23858 VDD.n1812 VDD.n1780 4.56231
R23859 VDD.n1868 VDD.n1842 4.56231
R23860 VDD.n5516 VDD.n1907 4.56231
R23861 VDD.n1960 VDD.n1934 4.56231
R23862 VDD.n2042 VDD.n2007 4.56231
R23863 VDD.n8752 VDD.n8748 4.56231
R23864 VDD.n8895 VDD.n8891 4.56231
R23865 VDD.n9068 VDD.n9064 4.56231
R23866 VDD.n6156 VDD.n6155 4.50663
R23867 VDD.n6099 VDD.n6098 4.50663
R23868 VDD.n6843 VDD.n6841 4.50663
R23869 VDD.n6793 VDD.n6728 4.50663
R23870 VDD.n59 VDD.n58 4.5005
R23871 VDD.n68 VDD.n63 4.5005
R23872 VDD.n148 VDD.n147 4.5005
R23873 VDD.n157 VDD.n152 4.5005
R23874 VDD.n5763 VDD.n5762 4.5005
R23875 VDD.n5758 VDD.n5757 4.5005
R23876 VDD.n5830 VDD.n5829 4.5005
R23877 VDD.n5825 VDD.n5824 4.5005
R23878 VDD.n5647 VDD.n5646 4.5005
R23879 VDD.n5642 VDD.n5641 4.5005
R23880 VDD.n5565 VDD.n5564 4.5005
R23881 VDD.n5560 VDD.n5559 4.5005
R23882 VDD.n8151 VDD.n8150 4.5005
R23883 VDD.n8146 VDD.n8145 4.5005
R23884 VDD.n6889 VDD.n6885 4.5005
R23885 VDD.n6894 VDD.n6884 4.5005
R23886 VDD.n6899 VDD.n6883 4.5005
R23887 VDD.n6981 VDD.n6882 4.5005
R23888 VDD.n6986 VDD.n6881 4.5005
R23889 VDD.n6991 VDD.n6880 4.5005
R23890 VDD.n6996 VDD.n6879 4.5005
R23891 VDD.n6908 VDD.n6904 4.5005
R23892 VDD.n6913 VDD.n6903 4.5005
R23893 VDD.n6918 VDD.n6902 4.5005
R23894 VDD.n6933 VDD.n6930 4.5005
R23895 VDD.n6938 VDD.n6929 4.5005
R23896 VDD.n6943 VDD.n6928 4.5005
R23897 VDD.n6948 VDD.n6927 4.5005
R23898 VDD.n5983 VDD.n5914 4.5005
R23899 VDD.n6322 VDD.n5914 4.5005
R23900 VDD.n6323 VDD.n6322 4.5005
R23901 VDD.n6324 VDD.n5914 4.5005
R23902 VDD.n5981 VDD.n5914 4.5005
R23903 VDD.n6323 VDD.n5981 4.5005
R23904 VDD.n6324 VDD.n6323 4.5005
R23905 VDD.n6422 VDD.n6418 4.5005
R23906 VDD.n6427 VDD.n6417 4.5005
R23907 VDD.n6432 VDD.n6416 4.5005
R23908 VDD.n6437 VDD.n6435 4.5005
R23909 VDD.n6440 VDD.n6438 4.5005
R23910 VDD.n6443 VDD.n6441 4.5005
R23911 VDD.n6446 VDD.n6444 4.5005
R23912 VDD.n6459 VDD.n6455 4.5005
R23913 VDD.n6464 VDD.n6454 4.5005
R23914 VDD.n6469 VDD.n6453 4.5005
R23915 VDD.n6474 VDD.n6472 4.5005
R23916 VDD.n6477 VDD.n6475 4.5005
R23917 VDD.n6480 VDD.n6478 4.5005
R23918 VDD.n6483 VDD.n6481 4.5005
R23919 VDD.n6102 VDD.n6040 4.5005
R23920 VDD.n6107 VDD.n6039 4.5005
R23921 VDD.n6111 VDD.n6110 4.5005
R23922 VDD.n6059 VDD.n6058 4.5005
R23923 VDD.n6064 VDD.n6057 4.5005
R23924 VDD.n6068 VDD.n6067 4.5005
R23925 VDD.n6173 VDD.n6015 4.5005
R23926 VDD.n6179 VDD.n6015 4.5005
R23927 VDD.n6179 VDD.n6012 4.5005
R23928 VDD.n6179 VDD.n6011 4.5005
R23929 VDD.n6179 VDD.n6178 4.5005
R23930 VDD.n6178 VDD.n6177 4.5005
R23931 VDD.n6177 VDD.n6011 4.5005
R23932 VDD.n7915 VDD.n7860 4.5005
R23933 VDD.n7920 VDD.n7859 4.5005
R23934 VDD.n7924 VDD.n7858 4.5005
R23935 VDD.n7929 VDD.n7857 4.5005
R23936 VDD.n7934 VDD.n7856 4.5005
R23937 VDD.n7939 VDD.n7855 4.5005
R23938 VDD.n7867 VDD.n7865 4.5005
R23939 VDD.n7871 VDD.n7869 4.5005
R23940 VDD.n7874 VDD.n7873 4.5005
R23941 VDD.n7877 VDD.n7875 4.5005
R23942 VDD.n7881 VDD.n7879 4.5005
R23943 VDD.n7885 VDD.n7883 4.5005
R23944 VDD.n8020 VDD.n2155 4.5005
R23945 VDD.n8025 VDD.n2154 4.5005
R23946 VDD.n8029 VDD.n2153 4.5005
R23947 VDD.n8034 VDD.n2152 4.5005
R23948 VDD.n8039 VDD.n2151 4.5005
R23949 VDD.n8044 VDD.n2150 4.5005
R23950 VDD.n6730 VDD.n6729 4.5005
R23951 VDD.n6733 VDD.n6731 4.5005
R23952 VDD.n6735 VDD.n6734 4.5005
R23953 VDD.n6748 VDD.n6747 4.5005
R23954 VDD.n6751 VDD.n6749 4.5005
R23955 VDD.n6741 VDD.n6740 4.5005
R23956 VDD.n8161 VDD.n8160 4.5005
R23957 VDD.n8160 VDD.n8142 4.5005
R23958 VDD.n8143 VDD.n8140 4.5005
R23959 VDD.n8143 VDD.n2089 4.5005
R23960 VDD.n5575 VDD.n5574 4.5005
R23961 VDD.n5574 VDD.n5555 4.5005
R23962 VDD.n5557 VDD.n5553 4.5005
R23963 VDD.n5557 VDD.n5556 4.5005
R23964 VDD.n10817 VDD.n2002 4.5005
R23965 VDD.n8092 VDD.n8091 4.5005
R23966 VDD.n8092 VDD.n2109 4.5005
R23967 VDD.n8095 VDD.n2109 4.5005
R23968 VDD.n8095 VDD.n8094 4.5005
R23969 VDD.n8094 VDD.n2105 4.5005
R23970 VDD.n2110 VDD.n2105 4.5005
R23971 VDD.n8091 VDD.n2105 4.5005
R23972 VDD.n10819 VDD.n2004 4.5005
R23973 VDD.n2004 VDD.n1996 4.5005
R23974 VDD.n2004 VDD.n2001 4.5005
R23975 VDD.n10820 VDD.n2001 4.5005
R23976 VDD.n10820 VDD.n1997 4.5005
R23977 VDD.n10820 VDD.n2002 4.5005
R23978 VDD.n10820 VDD.n1996 4.5005
R23979 VDD.n10820 VDD.n10819 4.5005
R23980 VDD.n5657 VDD.n5656 4.5005
R23981 VDD.n5656 VDD.n5546 4.5005
R23982 VDD.n5639 VDD.n5638 4.5005
R23983 VDD.n5639 VDD.n5544 4.5005
R23984 VDD.n5907 VDD.n5540 4.5005
R23985 VDD.n5908 VDD.n5907 4.5005
R23986 VDD.n5534 VDD.n5533 4.5005
R23987 VDD.n5533 VDD.n5503 4.5005
R23988 VDD.n5883 VDD.n1919 4.5005
R23989 VDD.n5890 VDD.n5883 4.5005
R23990 VDD.n5531 VDD.n5503 4.5005
R23991 VDD.n5890 VDD.n5881 4.5005
R23992 VDD.n5904 VDD.n5902 4.5005
R23993 VDD.n5535 VDD.n5534 4.5005
R23994 VDD.n5529 VDD.n5489 4.5005
R23995 VDD.n5535 VDD.n5529 4.5005
R23996 VDD.n5902 VDD.n5540 4.5005
R23997 VDD.n5908 VDD.n5902 4.5005
R23998 VDD.n5890 VDD.n5885 4.5005
R23999 VDD.n5890 VDD.n5880 4.5005
R24000 VDD.n5885 VDD.n1919 4.5005
R24001 VDD.n5880 VDD.n1919 4.5005
R24002 VDD.n5503 VDD.n5489 4.5005
R24003 VDD.n5840 VDD.n5839 4.5005
R24004 VDD.n5839 VDD.n5821 4.5005
R24005 VDD.n5822 VDD.n5819 4.5005
R24006 VDD.n5822 VDD.n5680 4.5005
R24007 VDD.n5773 VDD.n5772 4.5005
R24008 VDD.n5772 VDD.n5754 4.5005
R24009 VDD.n5755 VDD.n5752 4.5005
R24010 VDD.n5755 VDD.n5704 4.5005
R24011 VDD.n11048 VDD.n11047 4.5005
R24012 VDD.n11047 VDD.n11046 4.5005
R24013 VDD.n11046 VDD.n675 4.5005
R24014 VDD.n11046 VDD.n1764 4.5005
R24015 VDD.n11046 VDD.n674 4.5005
R24016 VDD.n11046 VDD.n11045 4.5005
R24017 VDD.n11045 VDD.n11044 4.5005
R24018 VDD.n11044 VDD.n674 4.5005
R24019 VDD.n11044 VDD.n1764 4.5005
R24020 VDD.n11130 VDD.n636 4.5005
R24021 VDD.n640 VDD.n636 4.5005
R24022 VDD.n11129 VDD.n640 4.5005
R24023 VDD.n640 VDD.n635 4.5005
R24024 VDD.n11127 VDD.n634 4.5005
R24025 VDD.n11130 VDD.n635 4.5005
R24026 VDD.n11130 VDD.n637 4.5005
R24027 VDD.n11130 VDD.n634 4.5005
R24028 VDD.n11130 VDD.n11129 4.5005
R24029 VDD.n5220 VDD.n4593 4.5005
R24030 VDD.n5220 VDD.n4594 4.5005
R24031 VDD.n5220 VDD.n5219 4.5005
R24032 VDD.n5204 VDD.n2408 4.5005
R24033 VDD.n4599 VDD.n2408 4.5005
R24034 VDD.n4591 VDD.n2425 4.5005
R24035 VDD.n4592 VDD.n4591 4.5005
R24036 VDD.n5219 VDD.n5218 4.5005
R24037 VDD.n9103 VDD.n9102 4.5005
R24038 VDD.n9112 VDD.n9107 4.5005
R24039 VDD.n8816 VDD.n8815 4.5005
R24040 VDD.n8825 VDD.n8820 4.5005
R24041 VDD.n8956 VDD.n8955 4.5005
R24042 VDD.n8965 VDD.n8960 4.5005
R24043 VDD.n9003 VDD.n9002 4.5005
R24044 VDD.n9004 VDD.n9003 4.5005
R24045 VDD.n9001 VDD.n9000 4.5005
R24046 VDD.n9000 VDD.n8953 4.5005
R24047 VDD.n8832 VDD.n8831 4.5005
R24048 VDD.n8833 VDD.n8832 4.5005
R24049 VDD.n8813 VDD.n8525 4.5005
R24050 VDD.n8813 VDD.n8812 4.5005
R24051 VDD.n9100 VDD.n9090 4.5005
R24052 VDD.n9100 VDD.n9099 4.5005
R24053 VDD.n9120 VDD.n9119 4.5005
R24054 VDD.n9119 VDD.n9118 4.5005
R24055 VDD.n9200 VDD.n9184 4.5005
R24056 VDD.n9184 VDD.n8458 4.5005
R24057 VDD.n12448 VDD.n194 4.5005
R24058 VDD.n12448 VDD.n12447 4.5005
R24059 VDD.n164 VDD.n163 4.5005
R24060 VDD.n165 VDD.n164 4.5005
R24061 VDD.n145 VDD.n135 4.5005
R24062 VDD.n145 VDD.n144 4.5005
R24063 VDD.n75 VDD.n74 4.5005
R24064 VDD.n76 VDD.n75 4.5005
R24065 VDD.n56 VDD.n46 4.5005
R24066 VDD.n56 VDD.n55 4.5005
R24067 VDD.n12583 VDD.n12580 4.5005
R24068 VDD.n12584 VDD.n12583 4.5005
R24069 VDD.n12581 VDD.n12580 4.5005
R24070 VDD.n12581 VDD.n12561 4.5005
R24071 VDD.n12585 VDD.n12561 4.5005
R24072 VDD.n12585 VDD.n12559 4.5005
R24073 VDD.n12585 VDD.n12584 4.5005
R24074 VDD.n12626 VDD.n8 4.5005
R24075 VDD.n12628 VDD.n9 4.5005
R24076 VDD.n12630 VDD.n12628 4.5005
R24077 VDD.n12630 VDD.n12623 4.5005
R24078 VDD.n12630 VDD.n8 4.5005
R24079 VDD.n12631 VDD.n9 4.5005
R24080 VDD.n12629 VDD.n9 4.5005
R24081 VDD.n12631 VDD.n12630 4.5005
R24082 VDD.n12630 VDD.n12629 4.5005
R24083 VDD.n1757 VDD.n680 4.5005
R24084 VDD.n1759 VDD.n680 4.5005
R24085 VDD.n1755 VDD.n680 4.5005
R24086 VDD.n1757 VDD.n678 4.5005
R24087 VDD.n1759 VDD.n678 4.5005
R24088 VDD.n678 VDD.n677 4.5005
R24089 VDD.n1755 VDD.n678 4.5005
R24090 VDD.n1756 VDD.n677 4.5005
R24091 VDD.n1756 VDD.n1755 4.5005
R24092 VDD.n1002 VDD.n1001 4.5005
R24093 VDD.n1003 VDD.n1002 4.5005
R24094 VDD.n956 VDD.n954 4.5005
R24095 VDD.n956 VDD.n953 4.5005
R24096 VDD.n1001 VDD.n956 4.5005
R24097 VDD.n1003 VDD.n956 4.5005
R24098 VDD.n1004 VDD.n954 4.5005
R24099 VDD.n1004 VDD.n953 4.5005
R24100 VDD.n1004 VDD.n1003 4.5005
R24101 VDD.n12641 VDD.n1 4.5005
R24102 VDD.n12642 VDD.n5 4.5005
R24103 VDD.n12642 VDD.n3 4.5005
R24104 VDD.n12642 VDD.n12636 4.5005
R24105 VDD.n12642 VDD.n12641 4.5005
R24106 VDD.n12640 VDD.n5 4.5005
R24107 VDD.n12640 VDD.n3 4.5005
R24108 VDD.n12640 VDD.n12636 4.5005
R24109 VDD.n12641 VDD.n12640 4.5005
R24110 VDD.n6092 VDD.n6041 4.32507
R24111 VDD.n6758 VDD.n6757 4.32507
R24112 VDD.n823 VDD.t2745 4.07396
R24113 VDD.n6952 VDD.t197 4.06712
R24114 VDD.n6925 VDD.t247 4.06712
R24115 VDD.n7010 VDD.t286 4.06712
R24116 VDD.n7003 VDD.t112 4.06712
R24117 VDD.n6502 VDD.t4937 4.06712
R24118 VDD.n6451 VDD.t4921 4.06712
R24119 VDD.n6542 VDD.t4860 4.06712
R24120 VDD.n6540 VDD.t4838 4.06712
R24121 VDD.n1477 VDD.t3029 4.05637
R24122 VDD.n1611 VDD.t4123 4.05637
R24123 VDD.n1609 VDD.t2799 4.05637
R24124 VDD.n1478 VDD.t1529 4.05637
R24125 VDD.n1117 VDD.t1627 4.05408
R24126 VDD.n1116 VDD.t4565 4.05408
R24127 VDD.n1182 VDD.t1987 4.05408
R24128 VDD.n1115 VDD.t1759 4.05408
R24129 VDD.n1114 VDD.t4729 4.05408
R24130 VDD.n1138 VDD.t1215 4.05408
R24131 VDD.n1137 VDD.t1683 4.05408
R24132 VDD.n1169 VDD.t3002 4.05408
R24133 VDD.n1136 VDD.t4139 4.05408
R24134 VDD.n1135 VDD.t1476 4.05408
R24135 VDD.n1312 VDD.t2375 4.05408
R24136 VDD.n1313 VDD.t3847 4.05408
R24137 VDD.n757 VDD.t2743 4.05408
R24138 VDD.n756 VDD.t1088 4.05408
R24139 VDD.n755 VDD.t2708 4.05408
R24140 VDD.n754 VDD.t3117 4.05408
R24141 VDD.n1280 VDD.t880 4.05408
R24142 VDD.n1308 VDD.t588 4.05408
R24143 VDD.n1278 VDD.t863 4.05408
R24144 VDD.n1279 VDD.t3797 4.05408
R24145 VDD.n1311 VDD.t3572 4.05408
R24146 VDD.n1080 VDD.t3497 4.05408
R24147 VDD.n1081 VDD.t888 4.05408
R24148 VDD.n1359 VDD.t3477 4.05408
R24149 VDD.n1282 VDD.t3667 4.05408
R24150 VDD.n1281 VDD.t3811 4.05408
R24151 VDD.n878 VDD.t3285 4.05408
R24152 VDD.n1076 VDD.t578 4.05408
R24153 VDD.n876 VDD.t2025 4.05408
R24154 VDD.n877 VDD.t4591 4.05408
R24155 VDD.n1079 VDD.t1993 4.05408
R24156 VDD.n1244 VDD.t4597 4.05408
R24157 VDD.n1245 VDD.t3433 4.05408
R24158 VDD.n765 VDD.t3541 4.05408
R24159 VDD.n766 VDD.t3341 4.05408
R24160 VDD.n767 VDD.t2135 4.05408
R24161 VDD.n768 VDD.t2934 4.05408
R24162 VDD.n805 VDD.t2109 4.05408
R24163 VDD.n1497 VDD.t1307 4.05408
R24164 VDD.n1498 VDD.t3219 4.05408
R24165 VDD.n1499 VDD.t4695 4.05408
R24166 VDD.n1601 VDD.t3521 4.05408
R24167 VDD.n1502 VDD.t1940 4.05408
R24168 VDD.n1503 VDD.t3505 4.05408
R24169 VDD.n1504 VDD.t3923 4.05408
R24170 VDD.n805 VDD.t2405 4.05408
R24171 VDD.n1497 VDD.t1521 4.05408
R24172 VDD.n1498 VDD.t3394 4.05408
R24173 VDD.n1499 VDD.t782 4.05408
R24174 VDD.n1601 VDD.t3726 4.05408
R24175 VDD.n1502 VDD.t2184 4.05408
R24176 VDD.n1503 VDD.t3706 4.05408
R24177 VDD.n1504 VDD.t4149 4.05408
R24178 VDD.n1109 VDD.t3193 4.05408
R24179 VDD.n1240 VDD.t4673 4.05408
R24180 VDD.n1107 VDD.t1703 4.05408
R24181 VDD.n1108 VDD.t1843 4.05408
R24182 VDD.n1243 VDD.t3418 4.05408
R24183 VDD.n1113 VDD.t717 4.05408
R24184 VDD.n1112 VDD.t3657 4.05408
R24185 VDD.n1212 VDD.t3483 4.05408
R24186 VDD.n1111 VDD.t4669 4.05408
R24187 VDD.n1110 VDD.t2476 4.05408
R24188 VDD.n727 VDD.t3105 4.05408
R24189 VDD.n1396 VDD.t3661 4.05408
R24190 VDD.n1395 VDD.t4115 4.05408
R24191 VDD.n1394 VDD.t1446 4.05408
R24192 VDD.n1391 VDD.t2966 4.05408
R24193 VDD.n1393 VDD.t1294 4.05408
R24194 VDD.n1404 VDD.t2952 4.05408
R24195 VDD.n1405 VDD.t3311 4.05408
R24196 VDD.n822 VDD.t3931 4.05408
R24197 VDD.n1446 VDD.t4343 4.05408
R24198 VDD.n819 VDD.t1697 4.05408
R24199 VDD.n820 VDD.t4313 4.05408
R24200 VDD.n817 VDD.t4509 4.05408
R24201 VDD.n816 VDD.t4659 4.05408
R24202 VDD.n815 VDD.t2419 4.05408
R24203 VDD.n812 VDD.t1544 4.05408
R24204 VDD.n811 VDD.t1693 4.05408
R24205 VDD.n809 VDD.t1468 4.05408
R24206 VDD.n810 VDD.t1679 4.05408
R24207 VDD.n807 VDD.t4653 4.05408
R24208 VDD.n806 VDD.t4407 4.05408
R24209 VDD.n727 VDD.t3295 4.05408
R24210 VDD.n1396 VDD.t3889 4.05408
R24211 VDD.n1395 VDD.t4311 4.05408
R24212 VDD.n1394 VDD.t1673 4.05408
R24213 VDD.n1391 VDD.t3157 4.05408
R24214 VDD.n1393 VDD.t1507 4.05408
R24215 VDD.n1404 VDD.t3145 4.05408
R24216 VDD.n1405 VDD.t3509 4.05408
R24217 VDD.n822 VDD.t4155 4.05408
R24218 VDD.n1446 VDD.t4527 4.05408
R24219 VDD.n819 VDD.t1931 4.05408
R24220 VDD.n820 VDD.t4511 4.05408
R24221 VDD.n817 VDD.t4737 4.05408
R24222 VDD.n816 VDD.t739 4.05408
R24223 VDD.n815 VDD.t2657 4.05408
R24224 VDD.n812 VDD.t1769 4.05408
R24225 VDD.n811 VDD.t1927 4.05408
R24226 VDD.n809 VDD.t1681 4.05408
R24227 VDD.n810 VDD.t1906 4.05408
R24228 VDD.n807 VDD.t735 4.05408
R24229 VDD.n806 VDD.t4637 4.05408
R24230 VDD.n900 VDD.t3257 4.05408
R24231 VDD.n899 VDD.t1525 4.05408
R24232 VDD.n1065 VDD.t1744 4.05408
R24233 VDD.n898 VDD.t1983 4.05408
R24234 VDD.n897 VDD.t1722 4.05408
R24235 VDD.n904 VDD.t1646 4.05408
R24236 VDD.n903 VDD.t2824 4.05408
R24237 VDD.n910 VDD.t4377 4.05408
R24238 VDD.n902 VDD.t4581 4.05408
R24239 VDD.n901 VDD.t4461 4.05408
R24240 VDD.n943 VDD.t2619 4.05408
R24241 VDD.n944 VDD.t3598 4.05408
R24242 VDD.n693 VDD.t1103 4.05408
R24243 VDD.n695 VDD.t1285 4.05408
R24244 VDD.n697 VDD.t1150 4.05408
R24245 VDD.n943 VDD.t2828 4.05408
R24246 VDD.n944 VDD.t3815 4.05408
R24247 VDD.n693 VDD.t1287 4.05408
R24248 VDD.n695 VDD.t1502 4.05408
R24249 VDD.n697 VDD.t1367 4.05408
R24250 VDD.n698 VDD.t1572 4.05408
R24251 VDD.n718 VDD.t2248 4.05408
R24252 VDD.n717 VDD.t4067 4.05408
R24253 VDD.n716 VDD.t2505 4.05408
R24254 VDD.n713 VDD.t2718 4.05408
R24255 VDD.n715 VDD.t2938 4.05408
R24256 VDD.n726 VDD.t2698 4.05408
R24257 VDD.n698 VDD.t1782 4.05408
R24258 VDD.n718 VDD.t2533 4.05408
R24259 VDD.n717 VDD.t4285 4.05408
R24260 VDD.n716 VDD.t2720 4.05408
R24261 VDD.n713 VDD.t2942 4.05408
R24262 VDD.n715 VDD.t3135 4.05408
R24263 VDD.n726 VDD.t2910 4.05408
R24264 VDD.n683 VDD.t3049 4.05408
R24265 VDD.n684 VDD.t737 4.05408
R24266 VDD.n1745 VDD.t4639 4.05408
R24267 VDD.n1158 VDD.t1677 4.05408
R24268 VDD.n1157 VDD.t4197 4.05408
R24269 VDD.n57 VDD.t528 4.00905
R24270 VDD.n146 VDD.t4760 4.00905
R24271 VDD.n9101 VDD.t4981 4.00905
R24272 VDD.n8814 VDD.t10 4.00905
R24273 VDD.n8954 VDD.t4797 4.00905
R24274 VDD.n5756 VDD.t372 4.00848
R24275 VDD.n5823 VDD.t4789 4.00848
R24276 VDD.n5640 VDD.t4747 4.00848
R24277 VDD.n5558 VDD.t514 4.00848
R24278 VDD.n8144 VDD.t389 4.00848
R24279 VDD.n60 VDD.t534 4.00673
R24280 VDD.n149 VDD.t4758 4.00673
R24281 VDD.n9104 VDD.t4979 4.00673
R24282 VDD.n8817 VDD.t5 4.00673
R24283 VDD.n8957 VDD.t4793 4.00673
R24284 VDD.n5759 VDD.t323 4.00554
R24285 VDD.n5826 VDD.t4788 4.00554
R24286 VDD.n5643 VDD.t4752 4.00554
R24287 VDD.n5561 VDD.t517 4.00554
R24288 VDD.n8147 VDD.t388 4.00554
R24289 VDD.n7012 VDD.n7011 3.96014
R24290 VDD.n6953 VDD.n6951 3.96014
R24291 VDD.n6543 VDD.n5289 3.96014
R24292 VDD.n6504 VDD.n6503 3.96014
R24293 VDD.n6952 VDD.t59 3.86107
R24294 VDD.n6925 VDD.t124 3.86107
R24295 VDD.n7010 VDD.t234 3.86107
R24296 VDD.n7003 VDD.t279 3.86107
R24297 VDD.n6502 VDD.t4847 3.86107
R24298 VDD.n6451 VDD.t4830 3.86107
R24299 VDD.n6542 VDD.t4908 3.86107
R24300 VDD.n6540 VDD.t4893 3.86107
R24301 VDD.n8641 VDD.t539 3.8555
R24302 VDD.n8700 VDD.t4780 3.8555
R24303 VDD.n1810 VDD.t418 3.8555
R24304 VDD.n1866 VDD.t4763 3.8555
R24305 VDD.n5514 VDD.t4779 3.8555
R24306 VDD.n1958 VDD.t505 3.8555
R24307 VDD.n2040 VDD.t489 3.8555
R24308 VDD.n8750 VDD.t292 3.8555
R24309 VDD.n8893 VDD.t495 3.8555
R24310 VDD.n9066 VDD.t4769 3.8555
R24311 VDD.n8640 VDD.t540 3.85313
R24312 VDD.n8699 VDD.t4782 3.85313
R24313 VDD.n1809 VDD.t421 3.85313
R24314 VDD.n1865 VDD.t4764 3.85313
R24315 VDD.n5513 VDD.t4778 3.85313
R24316 VDD.n1957 VDD.t503 3.85313
R24317 VDD.n2039 VDD.t4761 3.85313
R24318 VDD.n8749 VDD.t291 3.85313
R24319 VDD.n8892 VDD.t518 3.85313
R24320 VDD.n9065 VDD.t4768 3.85313
R24321 VDD.n6741 VDD.t150 3.84568
R24322 VDD.n6748 VDD.t168 3.84568
R24323 VDD.n6068 VDD.t4817 3.84568
R24324 VDD.n6059 VDD.t4938 3.84568
R24325 VDD.n6111 VDD.t4869 3.84568
R24326 VDD.n6102 VDD.t4809 3.84568
R24327 VDD.n6735 VDD.t77 3.84568
R24328 VDD.n6730 VDD.t100 3.84568
R24329 VDD.n6021 VDD.n6020 3.84528
R24330 VDD.n6155 VDD.n6154 3.84528
R24331 VDD.n6094 VDD.n6093 3.84528
R24332 VDD.n6098 VDD.n6097 3.84528
R24333 VDD.n6846 VDD.n6845 3.84528
R24334 VDD.n6843 VDD.n6842 3.84528
R24335 VDD.n6796 VDD.n6795 3.84528
R24336 VDD.n6793 VDD.n6792 3.84528
R24337 VDD.n7901 VDD.t28 3.84449
R24338 VDD.n2381 VDD.n2379 3.79678
R24339 VDD.n7019 VDD.n7017 3.79678
R24340 VDD.n6964 VDD.n6962 3.79678
R24341 VDD.n6972 VDD.n6970 3.79678
R24342 VDD.n5294 VDD.n5292 3.79678
R24343 VDD.n6557 VDD.n6555 3.79678
R24344 VDD.n6509 VDD.n6507 3.79678
R24345 VDD.n6518 VDD.n6516 3.79678
R24346 VDD.n6129 VDD.n6125 3.79678
R24347 VDD.n6144 VDD.n6140 3.79678
R24348 VDD.n6087 VDD.n6083 3.79678
R24349 VDD.n6052 VDD.n6048 3.79678
R24350 VDD.n6835 VDD.n6831 3.79678
R24351 VDD.n6818 VDD.n6814 3.79678
R24352 VDD.n6770 VDD.n6766 3.79678
R24353 VDD.n6785 VDD.n6781 3.79678
R24354 VDD.n5756 VDD.t419 3.78097
R24355 VDD.n5823 VDD.t4787 3.78097
R24356 VDD.n5640 VDD.t4746 3.78097
R24357 VDD.n5558 VDD.t513 3.78097
R24358 VDD.n8144 VDD.t333 3.78097
R24359 VDD.n5764 VDD.t299 3.78097
R24360 VDD.n5831 VDD.t4786 3.78097
R24361 VDD.n5648 VDD.t4745 3.78097
R24362 VDD.n5566 VDD.t512 3.78097
R24363 VDD.n8152 VDD.t332 3.78097
R24364 VDD.n57 VDD.t525 3.7804
R24365 VDD.n64 VDD.t526 3.7804
R24366 VDD.n146 VDD.t4754 3.7804
R24367 VDD.n153 VDD.t4756 3.7804
R24368 VDD.n9101 VDD.t4983 3.7804
R24369 VDD.n9108 VDD.t4977 3.7804
R24370 VDD.n8814 VDD.t7 3.7804
R24371 VDD.n8821 VDD.t8 3.7804
R24372 VDD.n8954 VDD.t4794 3.7804
R24373 VDD.n8961 VDD.t4795 3.7804
R24374 VDD.n59 VDD.t530 3.77818
R24375 VDD.n68 VDD.t531 3.77818
R24376 VDD.n148 VDD.t4753 3.77818
R24377 VDD.n157 VDD.t4755 3.77818
R24378 VDD.n5763 VDD.t294 3.77818
R24379 VDD.n5758 VDD.t420 3.77818
R24380 VDD.n5830 VDD.t4784 3.77818
R24381 VDD.n5825 VDD.t4785 3.77818
R24382 VDD.n5647 VDD.t4750 3.77818
R24383 VDD.n5642 VDD.t4751 3.77818
R24384 VDD.n5565 VDD.t515 3.77818
R24385 VDD.n5560 VDD.t516 3.77818
R24386 VDD.n8151 VDD.t329 3.77818
R24387 VDD.n8146 VDD.t330 3.77818
R24388 VDD.n9103 VDD.t4982 3.77818
R24389 VDD.n9112 VDD.t4984 3.77818
R24390 VDD.n8816 VDD.t11 3.77818
R24391 VDD.n8825 VDD.t3 3.77818
R24392 VDD.n8956 VDD.t4798 3.77818
R24393 VDD.n8965 VDD.t4799 3.77818
R24394 VDD.n6101 VDD.n6100 3.74038
R24395 VDD.n6807 VDD.n6806 3.74038
R24396 VDD.n6149 VDD.n6133 3.73034
R24397 VDD.n6079 VDD.n6075 3.73034
R24398 VDD.n6827 VDD.n6823 3.73034
R24399 VDD.n6790 VDD.n6774 3.73034
R24400 VDD.n7995 VDD.t23 3.7109
R24401 VDD.n980 VDD.n978 3.70005
R24402 VDD.n1038 VDD.n1037 3.70005
R24403 VDD.n1041 VDD.n1040 3.70005
R24404 VDD.n1102 VDD.n1101 3.70005
R24405 VDD.n1624 VDD.n1623 3.70005
R24406 VDD.n1090 VDD.n1089 3.70005
R24407 VDD.n1423 VDD.n1422 3.70005
R24408 VDD.n857 VDD.n856 3.70005
R24409 VDD.n1674 VDD.n746 3.70005
R24410 VDD.n1680 VDD.n743 3.70005
R24411 VDD.n1686 VDD.n740 3.70005
R24412 VDD.n1693 VDD.n737 3.70005
R24413 VDD.n982 VDD.n981 3.6965
R24414 VDD.n1036 VDD.n1035 3.6965
R24415 VDD.n1043 VDD.n1042 3.6965
R24416 VDD.n1104 VDD.n1103 3.6965
R24417 VDD.n1622 VDD.n1621 3.6965
R24418 VDD.n1088 VDD.n1087 3.6965
R24419 VDD.n1421 VDD.n1420 3.6965
R24420 VDD.n855 VDD.n854 3.6965
R24421 VDD.n1676 VDD.n1675 3.6965
R24422 VDD.n1682 VDD.n1681 3.6965
R24423 VDD.n1688 VDD.n1687 3.6965
R24424 VDD.n1695 VDD.n1694 3.6965
R24425 VDD.n8640 VDD.t542 3.68497
R24426 VDD.n8699 VDD.t4781 3.68497
R24427 VDD.n1809 VDD.t300 3.68497
R24428 VDD.n1865 VDD.t4762 3.68497
R24429 VDD.n5513 VDD.t4776 3.68497
R24430 VDD.n1957 VDD.t506 3.68497
R24431 VDD.n2039 VDD.t490 3.68497
R24432 VDD.n8749 VDD.t295 3.68497
R24433 VDD.n8892 VDD.t494 3.68497
R24434 VDD.n9065 VDD.t4766 3.68497
R24435 VDD.n7874 VDD.t31 3.68344
R24436 VDD.n8641 VDD.t541 3.68261
R24437 VDD.n8700 VDD.t4783 3.68261
R24438 VDD.n1810 VDD.t422 3.68261
R24439 VDD.n1866 VDD.t4765 3.68261
R24440 VDD.n5514 VDD.t4777 3.68261
R24441 VDD.n1958 VDD.t504 3.68261
R24442 VDD.n2040 VDD.t488 3.68261
R24443 VDD.n8750 VDD.t296 3.68261
R24444 VDD.n8893 VDD.t493 3.68261
R24445 VDD.n9066 VDD.t4767 3.68261
R24446 VDD.n7954 VDD.n7953 3.65594
R24447 VDD.n7015 VDD.n7014 3.65581
R24448 VDD.n7017 VDD.n7016 3.65581
R24449 VDD.n7019 VDD.n7018 3.65581
R24450 VDD.n7021 VDD.n7020 3.65581
R24451 VDD.n2383 VDD.n2382 3.65581
R24452 VDD.n2381 VDD.n2380 3.65581
R24453 VDD.n2379 VDD.n2378 3.65581
R24454 VDD.n6968 VDD.n6967 3.65581
R24455 VDD.n6970 VDD.n6969 3.65581
R24456 VDD.n6972 VDD.n6971 3.65581
R24457 VDD.n6974 VDD.n6973 3.65581
R24458 VDD.n6966 VDD.n6965 3.65581
R24459 VDD.n6964 VDD.n6963 3.65581
R24460 VDD.n6962 VDD.n6961 3.65581
R24461 VDD.n6559 VDD.n6558 3.65581
R24462 VDD.n6557 VDD.n6556 3.65581
R24463 VDD.n6555 VDD.n6554 3.65581
R24464 VDD.n6553 VDD.n6552 3.65581
R24465 VDD.n5296 VDD.n5295 3.65581
R24466 VDD.n5294 VDD.n5293 3.65581
R24467 VDD.n5292 VDD.n5291 3.65581
R24468 VDD.n6520 VDD.n6519 3.65581
R24469 VDD.n6518 VDD.n6517 3.65581
R24470 VDD.n6516 VDD.n6515 3.65581
R24471 VDD.n6514 VDD.n6513 3.65581
R24472 VDD.n6511 VDD.n6510 3.65581
R24473 VDD.n6509 VDD.n6508 3.65581
R24474 VDD.n6507 VDD.n6506 3.65581
R24475 VDD.n7949 VDD.n7948 3.6512
R24476 VDD.n7958 VDD.n7957 3.6512
R24477 VDD.n7951 VDD.n7950 3.6512
R24478 VDD.n7956 VDD.n7955 3.6512
R24479 VDD.n7022 VDD.n7021 3.64443
R24480 VDD.n6975 VDD.n6974 3.64443
R24481 VDD.n6553 VDD.n6551 3.64443
R24482 VDD.n6514 VDD.n6512 3.64443
R24483 VDD.n8029 VDD.t166 3.6266
R24484 VDD.n8054 VDD.n8053 3.62041
R24485 VDD.n8056 VDD.n8055 3.62041
R24486 VDD.n8059 VDD.n8058 3.62041
R24487 VDD.n8061 VDD.n8060 3.62041
R24488 VDD.n8063 VDD.n8062 3.62041
R24489 VDD.n7924 VDD.t57 3.61594
R24490 VDD.n62 VDD.n61 3.54958
R24491 VDD.n151 VDD.n150 3.54958
R24492 VDD.n5761 VDD.n5760 3.54958
R24493 VDD.n5828 VDD.n5827 3.54958
R24494 VDD.n5645 VDD.n5644 3.54958
R24495 VDD.n5563 VDD.n5562 3.54958
R24496 VDD.n8149 VDD.n8148 3.54958
R24497 VDD.n9106 VDD.n9105 3.54958
R24498 VDD.n8819 VDD.n8818 3.54958
R24499 VDD.n8959 VDD.n8958 3.54958
R24500 VDD.n6892 VDD.n6891 3.524
R24501 VDD.n6989 VDD.n6988 3.524
R24502 VDD.n6911 VDD.n6910 3.524
R24503 VDD.n6941 VDD.n6940 3.524
R24504 VDD.n6425 VDD.n6424 3.524
R24505 VDD.n6529 VDD.n6528 3.524
R24506 VDD.n6462 VDD.n6461 3.524
R24507 VDD.n6489 VDD.n6488 3.524
R24508 VDD.n6979 VDD.n6978 3.506
R24509 VDD.n6931 VDD.n6921 3.506
R24510 VDD.n6535 VDD.n6534 3.506
R24511 VDD.n6495 VDD.n6494 3.506
R24512 VDD.n1441 VDD.t382 3.3982
R24513 VDD.n804 VDD.t381 3.3982
R24514 VDD.n803 VDD.t384 3.3982
R24515 VDD.n1479 VDD.t378 3.3982
R24516 VDD.n814 VDD.t308 3.3982
R24517 VDD.n751 VDD.t385 3.37007
R24518 VDD.n1506 VDD.t370 3.37007
R24519 VDD.n6326 VDD.n5912 3.31078
R24520 VDD.n968 VDD.t485 3.29673
R24521 VDD.n941 VDD.t486 3.29673
R24522 VDD.n1140 VDD.t484 3.29673
R24523 VDD.n1141 VDD.t477 3.29673
R24524 VDD.n927 VDD.t483 3.29673
R24525 VDD.n926 VDD.t481 3.29673
R24526 VDD.n730 VDD.t482 3.29673
R24527 VDD.n731 VDD.t475 3.29673
R24528 VDD.n1289 VDD.t380 3.29673
R24529 VDD.n1288 VDD.t379 3.29673
R24530 VDD.n1119 VDD.t480 3.29673
R24531 VDD.n1120 VDD.t479 3.29673
R24532 VDD.n1191 VDD.t478 3.29673
R24533 VDD.n1321 VDD.t383 3.29673
R24534 VDD.n1320 VDD.t377 3.29673
R24535 VDD.n826 VDD.t473 3.29673
R24536 VDD.n1366 VDD.t387 3.29673
R24537 VDD.n5766 VDD.n5761 3.27995
R24538 VDD.n5833 VDD.n5828 3.27995
R24539 VDD.n5650 VDD.n5645 3.27995
R24540 VDD.n5568 VDD.n5563 3.27995
R24541 VDD.n8154 VDD.n8149 3.27995
R24542 VDD.n66 VDD.n62 3.27994
R24543 VDD.n155 VDD.n151 3.27994
R24544 VDD.n9110 VDD.n9106 3.27994
R24545 VDD.n8823 VDD.n8819 3.27994
R24546 VDD.n8963 VDD.n8959 3.27994
R24547 VDD.n1661 VDD.t3118 3.22144
R24548 VDD.t2935 VDD.n1643 3.22144
R24549 VDD.t1005 VDD.n6714 3.21228
R24550 VDD.n8637 VDD.t1808 3.20383
R24551 VDD.t2640 VDD.n12 3.20383
R24552 VDD.n12616 VDD.t1465 3.20383
R24553 VDD.n12620 VDD.t2664 3.20383
R24554 VDD.n12598 VDD.t4188 3.20383
R24555 VDD.n12594 VDD.t753 3.20383
R24556 VDD.n12591 VDD.t3828 3.20383
R24557 VDD.n12587 VDD.t778 3.20383
R24558 VDD.n12544 VDD.t4266 3.20383
R24559 VDD.n12548 VDD.t846 3.20383
R24560 VDD.n12550 VDD.t3916 3.20383
R24561 VDD.n12554 VDD.t1291 3.20383
R24562 VDD.n8654 VDD.t1905 3.20383
R24563 VDD.n8650 VDD.t2734 3.20383
R24564 VDD.n8648 VDD.t1541 3.20383
R24565 VDD.n8623 VDD.t3190 3.20383
R24566 VDD.n8675 VDD.t3681 3.20383
R24567 VDD.n8671 VDD.t728 3.20383
R24568 VDD.n8669 VDD.t3346 3.20383
R24569 VDD.n8665 VDD.t764 3.20383
R24570 VDD.n65 VDD.t527 3.20383
R24571 VDD.n67 VDD.t533 3.20383
R24572 VDD.n79 VDD.t1853 3.20383
R24573 VDD.n53 VDD.t3128 3.20383
R24574 VDD.n51 VDD.t1492 3.20383
R24575 VDD.t3152 VDD.n26 3.20383
R24576 VDD.n12504 VDD.t796 3.20383
R24577 VDD.n12500 VDD.t2423 3.20383
R24578 VDD.n94 VDD.t2241 3.20383
R24579 VDD.n90 VDD.t1997 3.20383
R24580 VDD.n8687 VDD.t2683 3.20383
R24581 VDD.n8683 VDD.t4182 3.20383
R24582 VDD.n8681 VDD.t4048 3.20383
R24583 VDD.n8677 VDD.t3818 3.20383
R24584 VDD.n8713 VDD.t2788 3.20383
R24585 VDD.n8709 VDD.t4260 3.20383
R24586 VDD.n8707 VDD.t1632 3.20383
R24587 VDD.n8607 VDD.t1403 3.20383
R24588 VDD.n12488 VDD.t903 3.20383
R24589 VDD.n12492 VDD.t2522 3.20383
R24590 VDD.n12494 VDD.t3996 3.20383
R24591 VDD.n12498 VDD.t3772 3.20383
R24592 VDD.n154 VDD.t4759 3.20383
R24593 VDD.n156 VDD.t4757 3.20383
R24594 VDD.n168 VDD.t2730 3.20383
R24595 VDD.n142 VDD.t4228 3.20383
R24596 VDD.n140 VDD.t4078 3.20383
R24597 VDD.t3858 VDD.n106 3.20383
R24598 VDD.n8725 VDD.t4454 3.20383
R24599 VDD.n8721 VDD.t1851 3.20383
R24600 VDD.n8719 VDD.t1709 3.20383
R24601 VDD.n8715 VDD.t1487 3.20383
R24602 VDD.n8746 VDD.t2345 3.20383
R24603 VDD.n8742 VDD.t3850 3.20383
R24604 VDD.n8740 VDD.t2383 3.20383
R24605 VDD.n8736 VDD.t2097 3.20383
R24606 VDD.n5721 VDD.t4222 3.20383
R24607 VDD.t1754 VDD.n1770 3.20383
R24608 VDD.n11032 VDD.t1241 3.20383
R24609 VDD.n11036 VDD.t3591 3.20383
R24610 VDD.n11021 VDD.t3693 3.20383
R24611 VDD.n11025 VDD.t2614 3.20383
R24612 VDD.n1778 VDD.t581 3.20383
R24613 VDD.n1774 VDD.t3946 3.20383
R24614 VDD.n1823 VDD.t4452 3.20383
R24615 VDD.n1819 VDD.t3316 3.20383
R24616 VDD.n1817 VDD.t1357 3.20383
R24617 VDD.n1808 VDD.t1554 3.20383
R24618 VDD.n5733 VDD.t3648 3.20383
R24619 VDD.n5729 VDD.t1225 3.20383
R24620 VDD.n5727 VDD.t730 3.20383
R24621 VDD.n5723 VDD.t1616 3.20383
R24622 VDD.n5776 VDD.t1316 3.20383
R24623 VDD.n5750 VDD.t1661 3.20383
R24624 VDD.n5748 VDD.t2656 3.20383
R24625 VDD.n5744 VDD.t3490 3.20383
R24626 VDD.n5765 VDD.t325 3.20383
R24627 VDD.n5767 VDD.t324 3.20383
R24628 VDD.n10982 VDD.t1501 3.20383
R24629 VDD.n10978 VDD.t1385 3.20383
R24630 VDD.n1829 VDD.t2691 3.20383
R24631 VDD.n1825 VDD.t2887 3.20383
R24632 VDD.n10966 VDD.t1136 3.20383
R24633 VDD.n10970 VDD.t1329 3.20383
R24634 VDD.n10972 VDD.t3628 3.20383
R24635 VDD.n10976 VDD.t2518 3.20383
R24636 VDD.n5788 VDD.t1361 3.20383
R24637 VDD.n5784 VDD.t2364 3.20383
R24638 VDD.n5782 VDD.t2140 3.20383
R24639 VDD.n5778 VDD.t3524 3.20383
R24640 VDD.n5809 VDD.t869 3.20383
R24641 VDD.n5805 VDD.t1727 3.20383
R24642 VDD.n5803 VDD.t3984 3.20383
R24643 VDD.n5799 VDD.t1175 3.20383
R24644 VDD.n1879 VDD.t1900 3.20383
R24645 VDD.n1875 VDD.t2116 3.20383
R24646 VDD.n1873 VDD.t703 3.20383
R24647 VDD.n1864 VDD.t3654 3.20383
R24648 VDD.n10927 VDD.t3200 3.20383
R24649 VDD.n10923 VDD.t3355 3.20383
R24650 VDD.n1894 VDD.t1443 3.20383
R24651 VDD.n1890 VDD.t4402 3.20383
R24652 VDD.n5843 VDD.t2775 3.20383
R24653 VDD.n5817 VDD.t3593 3.20383
R24654 VDD.n5815 VDD.t3458 3.20383
R24655 VDD.n5811 VDD.t644 3.20383
R24656 VDD.n5832 VDD.t4791 3.20383
R24657 VDD.n5834 VDD.t4790 3.20383
R24658 VDD.n5864 VDD.t2925 3.20383
R24659 VDD.n5860 VDD.t3750 3.20383
R24660 VDD.n5858 VDD.t4626 3.20383
R24661 VDD.n5854 VDD.t1842 3.20383
R24662 VDD.n10911 VDD.t3369 3.20383
R24663 VDD.n10915 VDD.t3571 3.20383
R24664 VDD.n10917 VDD.t572 3.20383
R24665 VDD.n10921 VDD.t3568 3.20383
R24666 VDD.n5527 VDD.t4562 3.20383
R24667 VDD.n5523 VDD.t3399 3.20383
R24668 VDD.n5521 VDD.t2973 3.20383
R24669 VDD.n5512 VDD.t608 3.20383
R24670 VDD.n5876 VDD.t4676 3.20383
R24671 VDD.n5872 VDD.t1887 3.20383
R24672 VDD.n5870 VDD.t933 3.20383
R24673 VDD.n5866 VDD.t3697 3.20383
R24674 VDD.n5637 VDD.t2817 3.20383
R24675 VDD.n5660 VDD.t1339 3.20383
R24676 VDD.n5662 VDD.t867 3.20383
R24677 VDD.n5666 VDD.t3214 3.20383
R24678 VDD.n5649 VDD.t4749 3.20383
R24679 VDD.n5651 VDD.t4748 3.20383
R24680 VDD.n10872 VDD.t2262 3.20383
R24681 VDD.n10868 VDD.t4164 3.20383
R24682 VDD.n5505 VDD.t2259 3.20383
R24683 VDD.n5509 VDD.t1379 3.20383
R24684 VDD.n10856 VDD.t2543 3.20383
R24685 VDD.n10860 VDD.t665 3.20383
R24686 VDD.n10862 VDD.t3014 3.20383
R24687 VDD.n10866 VDD.t2095 3.20383
R24688 VDD.n5616 VDD.t2983 3.20383
R24689 VDD.n5620 VDD.t3906 3.20383
R24690 VDD.n5622 VDD.t3391 3.20383
R24691 VDD.n5626 VDD.t1513 3.20383
R24692 VDD.n5595 VDD.t4724 3.20383
R24693 VDD.n5599 VDD.t3365 3.20383
R24694 VDD.n5601 VDD.t2922 3.20383
R24695 VDD.n5605 VDD.t3748 3.20383
R24696 VDD.n1971 VDD.t3679 3.20383
R24697 VDD.n1967 VDD.t1406 3.20383
R24698 VDD.n1965 VDD.t3676 3.20383
R24699 VDD.n1956 VDD.t3888 3.20383
R24700 VDD.n10814 VDD.t4436 3.20383
R24701 VDD.n10810 VDD.t3290 3.20383
R24702 VDD.n1986 VDD.t4432 3.20383
R24703 VDD.n1982 VDD.t4634 3.20383
R24704 VDD.t4210 VDD.n2104 3.20383
R24705 VDD.n5578 VDD.t1391 3.20383
R24706 VDD.n5580 VDD.t2378 3.20383
R24707 VDD.n5584 VDD.t3266 3.20383
R24708 VDD.n5567 VDD.t509 3.20383
R24709 VDD.n5569 VDD.t511 3.20383
R24710 VDD.n8109 VDD.t4106 3.20383
R24711 VDD.n8105 VDD.t862 3.20383
R24712 VDD.n8103 VDD.t672 3.20383
R24713 VDD.n8099 VDD.t2082 3.20383
R24714 VDD.n10798 VDD.t2740 3.20383
R24715 VDD.n10802 VDD.t2937 3.20383
R24716 VDD.n10804 VDD.t1001 3.20383
R24717 VDD.n10808 VDD.t3938 3.20383
R24718 VDD.n2053 VDD.t3424 3.20383
R24719 VDD.n2049 VDD.t3614 3.20383
R24720 VDD.n2047 VDD.t1712 3.20383
R24721 VDD.n2038 VDD.t4682 3.20383
R24722 VDD.n8121 VDD.t3550 3.20383
R24723 VDD.n8117 VDD.t4450 3.20383
R24724 VDD.n8115 VDD.t4298 3.20383
R24725 VDD.n8111 VDD.t1495 3.20383
R24726 VDD.n8164 VDD.t1204 3.20383
R24727 VDD.n8138 VDD.t2147 3.20383
R24728 VDD.n8136 VDD.t1980 3.20383
R24729 VDD.n8132 VDD.t3367 3.20383
R24730 VDD.n8153 VDD.t304 3.20383
R24731 VDD.n8155 VDD.t327 3.20383
R24732 VDD.n10767 VDD.t4616 3.20383
R24733 VDD.n10771 VDD.t670 3.20383
R24734 VDD.n2059 VDD.t3040 3.20383
R24735 VDD.n2055 VDD.t1731 3.20383
R24736 VDD.t2330 VDD.n2241 3.20383
R24737 VDD.n7095 VDD.t2330 3.20383
R24738 VDD.n7096 VDD.t3108 3.20383
R24739 VDD.n7105 VDD.t3970 3.20383
R24740 VDD.t3046 VDD.n7106 3.20383
R24741 VDD.n7113 VDD.t1920 3.20383
R24742 VDD.n7114 VDD.t2425 3.20383
R24743 VDD.n7123 VDD.t2247 3.20383
R24744 VDD.t4336 VDD.n2241 3.20383
R24745 VDD.n7095 VDD.t4336 3.20383
R24746 VDD.n7096 VDD.t970 3.20383
R24747 VDD.n7105 VDD.t1839 3.20383
R24748 VDD.n7106 VDD.t901 3.20383
R24749 VDD.n7113 VDD.t4004 3.20383
R24750 VDD.n7114 VDD.t4392 3.20383
R24751 VDD.n7123 VDD.t4284 3.20383
R24752 VDD.t1814 VDD.n2265 3.20383
R24753 VDD.n7079 VDD.t2839 3.20383
R24754 VDD.t1735 VDD.n7080 3.20383
R24755 VDD.t732 VDD.n7064 3.20383
R24756 VDD.n7061 VDD.t1132 3.20383
R24757 VDD.n7051 VDD.t1022 3.20383
R24758 VDD.n7050 VDD.t1061 3.20383
R24759 VDD.t1061 VDD.n7049 3.20383
R24760 VDD.t695 VDD.n2342 3.20383
R24761 VDD.n6656 VDD.t695 3.20383
R24762 VDD.n6657 VDD.t1435 3.20383
R24763 VDD.n6666 VDD.t1314 3.20383
R24764 VDD.t831 VDD.n6667 3.20383
R24765 VDD.n6674 VDD.t4492 3.20383
R24766 VDD.n6675 VDD.t4012 3.20383
R24767 VDD.n6684 VDD.t3415 3.20383
R24768 VDD.t1833 VDD.n2265 3.20383
R24769 VDD.n7079 VDD.t2853 3.20383
R24770 VDD.n7080 VDD.t1750 3.20383
R24771 VDD.n7064 VDD.t758 3.20383
R24772 VDD.n7061 VDD.t1145 3.20383
R24773 VDD.t1034 VDD.n7051 3.20383
R24774 VDD.n7050 VDD.t1071 3.20383
R24775 VDD.n7049 VDD.t1071 3.20383
R24776 VDD.t716 VDD.n2342 3.20383
R24777 VDD.n6656 VDD.t716 3.20383
R24778 VDD.n6657 VDD.t1467 3.20383
R24779 VDD.n6666 VDD.t1327 3.20383
R24780 VDD.n6667 VDD.t858 3.20383
R24781 VDD.n6674 VDD.t4506 3.20383
R24782 VDD.n6675 VDD.t4026 3.20383
R24783 VDD.n6684 VDD.t3430 3.20383
R24784 VDD.n2396 VDD.t3270 3.20383
R24785 VDD.n7033 VDD.t3150 3.20383
R24786 VDD.t2650 VDD.n7034 3.20383
R24787 VDD.n6718 VDD.t2102 3.20383
R24788 VDD.t1552 VDD.n6719 3.20383
R24789 VDD.n6875 VDD.t3589 3.20383
R24790 VDD.n6866 VDD.t4478 3.20383
R24791 VDD.n6865 VDD.t3514 3.20383
R24792 VDD.t2555 VDD.n6858 3.20383
R24793 VDD.n6857 VDD.t2975 3.20383
R24794 VDD.n2403 VDD.t2843 3.20383
R24795 VDD.t2762 VDD.n2322 3.20383
R24796 VDD.n5244 VDD.t2636 3.20383
R24797 VDD.t2040 VDD.n5245 3.20383
R24798 VDD.n5252 VDD.t1532 3.20383
R24799 VDD.n5253 VDD.t1045 3.20383
R24800 VDD.n5262 VDD.t4572 3.20383
R24801 VDD.t4726 VDD.n2322 3.20383
R24802 VDD.n5244 VDD.t4578 3.20383
R24803 VDD.n5245 VDD.t4102 3.20383
R24804 VDD.n5252 VDD.t3622 3.20383
R24805 VDD.n5253 VDD.t3162 3.20383
R24806 VDD.n5262 VDD.t2592 3.20383
R24807 VDD.n6360 VDD.t4418 3.20383
R24808 VDD.n6350 VDD.t4300 3.20383
R24809 VDD.n6349 VDD.t3788 3.20383
R24810 VDD.t2334 VDD.n6342 3.20383
R24811 VDD.n6341 VDD.t3230 3.20383
R24812 VDD.n6331 VDD.t4096 3.20383
R24813 VDD.n6330 VDD.t4372 3.20383
R24814 VDD.t4372 VDD.n6329 3.20383
R24815 VDD.n6360 VDD.t3338 3.20383
R24816 VDD.t3264 VDD.n6350 3.20383
R24817 VDD.n6349 VDD.t2786 3.20383
R24818 VDD.n6342 VDD.t1167 3.20383
R24819 VDD.n6341 VDD.t2086 3.20383
R24820 VDD.t3056 VDD.n6331 3.20383
R24821 VDD.n6330 VDD.t3310 3.20383
R24822 VDD.n6329 VDD.t3310 3.20383
R24823 VDD.n5445 VDD.t628 3.20383
R24824 VDD.n5454 VDD.t4668 3.20383
R24825 VDD.t4176 VDD.n5455 3.20383
R24826 VDD.n5462 VDD.t3689 3.20383
R24827 VDD.n5463 VDD.t4542 3.20383
R24828 VDD.n5472 VDD.t3994 3.20383
R24829 VDD.n5445 VDD.t3701 3.20383
R24830 VDD.n5454 VDD.t3583 3.20383
R24831 VDD.n5455 VDD.t3122 3.20383
R24832 VDD.n5462 VDD.t2678 3.20383
R24833 VDD.n5463 VDD.t3500 3.20383
R24834 VDD.n5472 VDD.t2971 3.20383
R24835 VDD.n6593 VDD.t2458 3.20383
R24836 VDD.n6584 VDD.t2282 3.20383
R24837 VDD.n6583 VDD.t1700 3.20383
R24838 VDD.n5926 VDD.t1243 3.20383
R24839 VDD.n5927 VDD.t2171 3.20383
R24840 VDD.n5936 VDD.t1528 3.20383
R24841 VDD.t3900 VDD.n5265 3.20383
R24842 VDD.n6242 VDD.t3770 3.20383
R24843 VDD.t3292 VDD.n6243 3.20383
R24844 VDD.n6250 VDD.t2865 3.20383
R24845 VDD.n6251 VDD.t3664 3.20383
R24846 VDD.n6260 VDD.t3142 3.20383
R24847 VDD.t734 VDD.n6261 3.20383
R24848 VDD.n6262 VDD.t734 3.20383
R24849 VDD.t1690 VDD.n6267 3.20383
R24850 VDD.n6268 VDD.t1690 3.20383
R24851 VDD.n6269 VDD.t3534 3.20383
R24852 VDD.n6278 VDD.t3411 3.20383
R24853 VDD.t2963 VDD.n6279 3.20383
R24854 VDD.n6286 VDD.t1347 3.20383
R24855 VDD.n6287 VDD.t2309 3.20383
R24856 VDD.n6296 VDD.t3234 3.20383
R24857 VDD.t3492 VDD.n6297 3.20383
R24858 VDD.n6298 VDD.t3492 3.20383
R24859 VDD.t3918 VDD.n5265 3.20383
R24860 VDD.n6242 VDD.t3786 3.20383
R24861 VDD.n6243 VDD.t3300 3.20383
R24862 VDD.n6250 VDD.t2877 3.20383
R24863 VDD.n6251 VDD.t3683 3.20383
R24864 VDD.n6260 VDD.t3156 3.20383
R24865 VDD.n6261 VDD.t760 3.20383
R24866 VDD.n6262 VDD.t760 3.20383
R24867 VDD.n6267 VDD.t1706 3.20383
R24868 VDD.n6268 VDD.t1706 3.20383
R24869 VDD.n6269 VDD.t3544 3.20383
R24870 VDD.n6278 VDD.t3432 3.20383
R24871 VDD.n6279 VDD.t2979 3.20383
R24872 VDD.n6286 VDD.t1363 3.20383
R24873 VDD.n6287 VDD.t2332 3.20383
R24874 VDD.n6296 VDD.t3248 3.20383
R24875 VDD.n6297 VDD.t3502 3.20383
R24876 VDD.n6298 VDD.t3502 3.20383
R24877 VDD.n5951 VDD.t2009 3.20383
R24878 VDD.n5960 VDD.t1863 3.20383
R24879 VDD.t1336 VDD.n5961 3.20383
R24880 VDD.n5968 VDD.t4024 3.20383
R24881 VDD.n5969 VDD.t762 3.20383
R24882 VDD.n5978 VDD.t1645 3.20383
R24883 VDD.n6380 VDD.t4720 3.20383
R24884 VDD.n6389 VDD.t4570 3.20383
R24885 VDD.t4094 VDD.n6390 3.20383
R24886 VDD.n5997 VDD.t2660 3.20383
R24887 VDD.n5998 VDD.t3482 3.20383
R24888 VDD.n6007 VDD.t4368 3.20383
R24889 VDD.n6009 VDD.t4672 3.20383
R24890 VDD.t4672 VDD.n6008 3.20383
R24891 VDD.n6380 VDD.t2717 3.20383
R24892 VDD.n6389 VDD.t2590 3.20383
R24893 VDD.n6390 VDD.t1978 3.20383
R24894 VDD.n5997 VDD.t4614 3.20383
R24895 VDD.n5998 VDD.t1343 3.20383
R24896 VDD.n6007 VDD.t2338 3.20383
R24897 VDD.n6009 VDD.t2666 3.20383
R24898 VDD.n6008 VDD.t2666 3.20383
R24899 VDD.t960 VDD.n5263 3.20383
R24900 VDD.n5343 VDD.t821 3.20383
R24901 VDD.t4442 VDD.n5344 3.20383
R24902 VDD.n5351 VDD.t3998 3.20383
R24903 VDD.n5352 VDD.t714 3.20383
R24904 VDD.n5361 VDD.t4278 3.20383
R24905 VDD.t3078 VDD.n5263 3.20383
R24906 VDD.n5343 VDD.t2961 3.20383
R24907 VDD.n5344 VDD.t2431 3.20383
R24908 VDD.n5351 VDD.t1872 3.20383
R24909 VDD.n5352 VDD.t2861 3.20383
R24910 VDD.n5361 VDD.t2200 3.20383
R24911 VDD.n6412 VDD.t1108 3.20383
R24912 VDD.n6403 VDD.t1003 3.20383
R24913 VDD.n6402 VDD.t4596 3.20383
R24914 VDD.n6161 VDD.t3170 3.20383
R24915 VDD.n6162 VDD.t4014 3.20383
R24916 VDD.n6171 VDD.t776 3.20383
R24917 VDD.t1451 VDD.n2410 3.20383
R24918 VDD.n6570 VDD.t1318 3.20383
R24919 VDD.t850 VDD.n6571 3.20383
R24920 VDD.n6028 VDD.t4500 3.20383
R24921 VDD.t1231 VDD.n6029 3.20383
R24922 VDD.t646 VDD.n6024 3.20383
R24923 VDD.n2216 VDD.t1214 3.20383
R24924 VDD.n2227 VDD.t4386 3.20383
R24925 VDD.n2219 VDD.t3379 3.20383
R24926 VDD.n2218 VDD.t3792 3.20383
R24927 VDD.t3646 VDD.n7980 3.20383
R24928 VDD.n7976 VDD.t3687 3.20383
R24929 VDD.t3687 VDD.n7975 3.20383
R24930 VDD.n7969 VDD.t3350 3.20383
R24931 VDD.t3350 VDD.n7968 3.20383
R24932 VDD.n7965 VDD.t4132 3.20383
R24933 VDD.n7851 VDD.t2784 3.20383
R24934 VDD.t2784 VDD.n7850 3.20383
R24935 VDD.n2215 VDD.t4480 3.20383
R24936 VDD.t4360 VDD.n2193 3.20383
R24937 VDD.n7986 VDD.t1106 3.20383
R24938 VDD.t3401 VDD.n7983 3.20383
R24939 VDD.n7979 VDD.t1429 3.20383
R24940 VDD.n7966 VDD.t1882 3.20383
R24941 VDD.t2756 VDD.n2202 3.20383
R24942 VDD.n2203 VDD.t2756 3.20383
R24943 VDD.n6605 VDD.t3990 3.20383
R24944 VDD.t3480 VDD.n6606 3.20383
R24945 VDD.n6613 VDD.t3072 3.20383
R24946 VDD.n6614 VDD.t2564 3.20383
R24947 VDD.n6623 VDD.t1865 3.20383
R24948 VDD.t2460 VDD.n2310 3.20383
R24949 VDD.n5415 VDD.t2284 3.20383
R24950 VDD.t1702 VDD.n5416 3.20383
R24951 VDD.n5423 VDD.t1245 3.20383
R24952 VDD.n5424 VDD.t766 3.20383
R24953 VDD.n5433 VDD.t4302 3.20383
R24954 VDD.t1258 VDD.n2310 3.20383
R24955 VDD.n5415 VDD.t1134 3.20383
R24956 VDD.n5416 VDD.t601 3.20383
R24957 VDD.n5423 VDD.t4318 3.20383
R24958 VDD.n5424 VDD.t3808 3.20383
R24959 VDD.n5433 VDD.t3262 3.20383
R24960 VDD.n7174 VDD.t1976 3.20383
R24961 VDD.t1976 VDD.n7173 3.20383
R24962 VDD.n7172 VDD.t2833 3.20383
R24963 VDD.n7162 VDD.t3652 3.20383
R24964 VDD.n7161 VDD.t2760 3.20383
R24965 VDD.t1620 VDD.n7154 3.20383
R24966 VDD.n7153 VDD.t2074 3.20383
R24967 VDD.n7143 VDD.t1915 3.20383
R24968 VDD.n7174 VDD.t913 3.20383
R24969 VDD.n7173 VDD.t913 3.20383
R24970 VDD.n7172 VDD.t1634 3.20383
R24971 VDD.t2654 VDD.n7162 3.20383
R24972 VDD.n7161 VDD.t1547 3.20383
R24973 VDD.n7154 VDD.t4688 3.20383
R24974 VDD.n7153 VDD.t986 3.20383
R24975 VDD.t848 VDD.n7143 3.20383
R24976 VDD.n7843 VDD.t4466 3.20383
R24977 VDD.n2173 VDD.t2802 3.20383
R24978 VDD.n2182 VDD.t2670 3.20383
R24979 VDD.t3494 VDD.n2183 3.20383
R24980 VDD.n8000 VDD.t1585 3.20383
R24981 VDD.n8001 VDD.t3834 3.20383
R24982 VDD.n8010 VDD.t4276 3.20383
R24983 VDD.t3518 VDD.n8459 3.20383
R24984 VDD.t3322 VDD.n9130 3.20383
R24985 VDD.t2999 VDD.n8459 3.20383
R24986 VDD.n9130 VDD.t2794 3.20383
R24987 VDD.n9139 VDD.t2547 3.20383
R24988 VDD.n9143 VDD.t4042 3.20383
R24989 VDD.n9145 VDD.t3898 3.20383
R24990 VDD.n9149 VDD.t3672 3.20383
R24991 VDD.n9166 VDD.t3102 3.20383
R24992 VDD.n9162 VDD.t4568 3.20383
R24993 VDD.t4460 VDD.n8472 3.20383
R24994 VDD.n8488 VDD.t4256 3.20383
R24995 VDD.n9109 VDD.t4980 3.20383
R24996 VDD.n9111 VDD.t4978 3.20383
R24997 VDD.n8763 VDD.t4060 3.20383
R24998 VDD.n8759 VDD.t3840 3.20383
R24999 VDD.n8757 VDD.t4516 3.20383
R25000 VDD.n8582 VDD.t3860 3.20383
R25001 VDD.n8559 VDD.t2252 3.20383
R25002 VDD.n8555 VDD.t2022 3.20383
R25003 VDD.n8553 VDD.t2813 3.20383
R25004 VDD.t2059 VDD.n184 3.20383
R25005 VDD.n8822 VDD.t9 3.20383
R25006 VDD.n8824 VDD.t4 3.20383
R25007 VDD.n8836 VDD.t2869 3.20383
R25008 VDD.n8810 VDD.t2108 3.20383
R25009 VDD.t1032 VDD.n8526 3.20383
R25010 VDD.n8547 VDD.t2130 3.20383
R25011 VDD.n8799 VDD.t4584 3.20383
R25012 VDD.n8803 VDD.t3934 3.20383
R25013 VDD.n8769 VDD.t2941 3.20383
R25014 VDD.n8765 VDD.t3958 3.20383
R25015 VDD.n8889 VDD.t2520 3.20383
R25016 VDD.n8885 VDD.t3446 3.20383
R25017 VDD.t2437 VDD.n8518 3.20383
R25018 VDD.n8775 VDD.t3470 3.20383
R25019 VDD.n8872 VDD.t577 3.20383
R25020 VDD.n8876 VDD.t1591 3.20383
R25021 VDD.n8842 VDD.t4692 3.20383
R25022 VDD.n8838 VDD.t1618 3.20383
R25023 VDD.n8945 VDD.t2467 3.20383
R25024 VDD.n8941 VDD.t1676 3.20383
R25025 VDD.t596 VDD.n8507 3.20383
R25026 VDD.n8848 VDD.t2210 3.20383
R25027 VDD.n8930 VDD.t4226 3.20383
R25028 VDD.n8934 VDD.t3526 3.20383
R25029 VDD.n8900 VDD.t2528 3.20383
R25030 VDD.n8513 VDD.t4018 3.20383
R25031 VDD.n9020 VDD.t4290 3.20383
R25032 VDD.n9016 VDD.t4082 3.20383
R25033 VDD.t2624 VDD.n8499 3.20383
R25034 VDD.n8906 VDD.t4110 3.20383
R25035 VDD.n8962 VDD.t4796 3.20383
R25036 VDD.n8964 VDD.t4792 3.20383
R25037 VDD.n8999 VDD.t2560 3.20383
R25038 VDD.n9007 VDD.t2289 3.20383
R25039 VDD.n8951 VDD.t708 3.20383
R25040 VDD.n8947 VDD.t2326 3.20383
R25041 VDD.n9042 VDD.t3024 3.20383
R25042 VDD.n9038 VDD.t4486 3.20383
R25043 VDD.t4366 VDD.n8490 3.20383
R25044 VDD.n8975 VDD.t4178 3.20383
R25045 VDD.t561 VDD.n8476 3.20383
R25046 VDD.n9031 VDD.t2190 3.20383
R25047 VDD.n9026 VDD.t2062 3.20383
R25048 VDD.n9022 VDD.t1797 3.20383
R25049 VDD.n9151 VDD.t681 3.20383
R25050 VDD.n9155 VDD.t2303 3.20383
R25051 VDD.n9073 VDD.t2128 3.20383
R25052 VDD.n8475 VDD.t1894 3.20383
R25053 VDD.n190 VDD.t4604 3.20383
R25054 VDD.n186 VDD.t2044 3.20383
R25055 VDD.n174 VDD.t4630 3.20383
R25056 VDD.n170 VDD.t4406 3.20383
R25057 VDD.n9123 VDD.t623 3.20383
R25058 VDD.n9097 VDD.t2229 3.20383
R25059 VDD.n9095 VDD.t2089 3.20383
R25060 VDD.t1837 VDD.n8470 3.20383
R25061 VDD.n1162 VDD.t4198 3.20383
R25062 VDD.t4198 VDD.n1161 3.20383
R25063 VDD.n1160 VDD.t1678 3.20383
R25064 VDD.n1748 VDD.t738 3.20383
R25065 VDD.t3050 VDD.n1749 3.20383
R25066 VDD.n1750 VDD.t3050 3.20383
R25067 VDD.t2911 VDD.n1711 3.20383
R25068 VDD.n1712 VDD.t2911 3.20383
R25069 VDD.t3136 VDD.n1713 3.20383
R25070 VDD.n722 VDD.t2721 3.20383
R25071 VDD.n721 VDD.t4286 3.20383
R25072 VDD.t4286 VDD.n720 3.20383
R25073 VDD.n719 VDD.t2534 3.20383
R25074 VDD.t2534 VDD.n700 3.20383
R25075 VDD.t1783 VDD.n1733 3.20383
R25076 VDD.n1734 VDD.t1783 3.20383
R25077 VDD.n1711 VDD.t2699 3.20383
R25078 VDD.n1712 VDD.t2699 3.20383
R25079 VDD.n1713 VDD.t2939 3.20383
R25080 VDD.t2506 VDD.n722 3.20383
R25081 VDD.n721 VDD.t4068 3.20383
R25082 VDD.n720 VDD.t4068 3.20383
R25083 VDD.n719 VDD.t2249 3.20383
R25084 VDD.t2249 VDD.n700 3.20383
R25085 VDD.n1733 VDD.t1573 3.20383
R25086 VDD.n1734 VDD.t1573 3.20383
R25087 VDD.t1368 VDD.n1735 3.20383
R25088 VDD.n1736 VDD.t1368 3.20383
R25089 VDD.t1503 VDD.n1737 3.20383
R25090 VDD.n948 VDD.t3816 3.20383
R25091 VDD.t2829 VDD.n950 3.20383
R25092 VDD.n951 VDD.t2829 3.20383
R25093 VDD.n916 VDD.t4462 3.20383
R25094 VDD.t4462 VDD.n915 3.20383
R25095 VDD.n914 VDD.t4582 3.20383
R25096 VDD.t2825 VDD.n907 3.20383
R25097 VDD.n906 VDD.t1647 3.20383
R25098 VDD.t1647 VDD.n905 3.20383
R25099 VDD.n1071 VDD.t1723 3.20383
R25100 VDD.t1723 VDD.n1070 3.20383
R25101 VDD.n1069 VDD.t1984 3.20383
R25102 VDD.t1526 VDD.n1062 3.20383
R25103 VDD.n1061 VDD.t3258 3.20383
R25104 VDD.t3258 VDD.n1060 3.20383
R25105 VDD.n1494 VDD.t4638 3.20383
R25106 VDD.t4638 VDD.n1493 3.20383
R25107 VDD.n1492 VDD.t736 3.20383
R25108 VDD.t1682 VDD.n1485 3.20383
R25109 VDD.n1484 VDD.t1928 3.20383
R25110 VDD.t1928 VDD.n1483 3.20383
R25111 VDD.n1482 VDD.t1770 3.20383
R25112 VDD.t1770 VDD.n1481 3.20383
R25113 VDD.n1461 VDD.t2658 3.20383
R25114 VDD.t2658 VDD.n1460 3.20383
R25115 VDD.n1459 VDD.t740 3.20383
R25116 VDD.t740 VDD.n1458 3.20383
R25117 VDD.n1457 VDD.t4738 3.20383
R25118 VDD.t1932 VDD.n1450 3.20383
R25119 VDD.t4528 VDD.n821 3.20383
R25120 VDD.n1445 VDD.t4528 3.20383
R25121 VDD.n1444 VDD.t4156 3.20383
R25122 VDD.t4156 VDD.n1443 3.20383
R25123 VDD.t3510 VDD.n824 3.20383
R25124 VDD.n1406 VDD.t3510 3.20383
R25125 VDD.t3146 VDD.n1407 3.20383
R25126 VDD.n1408 VDD.t3146 3.20383
R25127 VDD.t1508 VDD.n1409 3.20383
R25128 VDD.n1400 VDD.t1674 3.20383
R25129 VDD.n1399 VDD.t4312 3.20383
R25130 VDD.t4312 VDD.n1398 3.20383
R25131 VDD.n1397 VDD.t3890 3.20383
R25132 VDD.t3890 VDD.n729 3.20383
R25133 VDD.t3296 VDD.n1709 3.20383
R25134 VDD.n1710 VDD.t3296 3.20383
R25135 VDD.n1494 VDD.t4408 3.20383
R25136 VDD.n1493 VDD.t4408 3.20383
R25137 VDD.n1492 VDD.t4654 3.20383
R25138 VDD.n1485 VDD.t1469 3.20383
R25139 VDD.n1484 VDD.t1694 3.20383
R25140 VDD.n1483 VDD.t1694 3.20383
R25141 VDD.n1482 VDD.t1545 3.20383
R25142 VDD.n1481 VDD.t1545 3.20383
R25143 VDD.n1461 VDD.t2420 3.20383
R25144 VDD.n1460 VDD.t2420 3.20383
R25145 VDD.n1459 VDD.t4660 3.20383
R25146 VDD.n1458 VDD.t4660 3.20383
R25147 VDD.n1457 VDD.t4510 3.20383
R25148 VDD.n1450 VDD.t1698 3.20383
R25149 VDD.t4344 VDD.n821 3.20383
R25150 VDD.n1445 VDD.t4344 3.20383
R25151 VDD.n1444 VDD.t3932 3.20383
R25152 VDD.n1443 VDD.t3932 3.20383
R25153 VDD.t3312 VDD.n824 3.20383
R25154 VDD.n1406 VDD.t3312 3.20383
R25155 VDD.n1407 VDD.t2953 3.20383
R25156 VDD.n1408 VDD.t2953 3.20383
R25157 VDD.n1409 VDD.t1295 3.20383
R25158 VDD.t1447 VDD.n1400 3.20383
R25159 VDD.n1399 VDD.t4116 3.20383
R25160 VDD.n1398 VDD.t4116 3.20383
R25161 VDD.n1397 VDD.t3662 3.20383
R25162 VDD.t3662 VDD.n729 3.20383
R25163 VDD.n1709 VDD.t3106 3.20383
R25164 VDD.n1710 VDD.t3106 3.20383
R25165 VDD.n1218 VDD.t2477 3.20383
R25166 VDD.t2477 VDD.n1217 3.20383
R25167 VDD.n1216 VDD.t4670 3.20383
R25168 VDD.t3658 VDD.n1209 3.20383
R25169 VDD.n1208 VDD.t718 3.20383
R25170 VDD.t718 VDD.n1207 3.20383
R25171 VDD.t3419 VDD.n1270 3.20383
R25172 VDD.n1271 VDD.t3419 3.20383
R25173 VDD.t1844 VDD.n1272 3.20383
R25174 VDD.n1239 VDD.t4674 3.20383
R25175 VDD.n1238 VDD.t3194 3.20383
R25176 VDD.t3194 VDD.n1237 3.20383
R25177 VDD.t4150 VDD.n1593 3.20383
R25178 VDD.n1594 VDD.t4150 3.20383
R25179 VDD.t3707 VDD.n1595 3.20383
R25180 VDD.n1596 VDD.t3707 3.20383
R25181 VDD.t2185 VDD.n1597 3.20383
R25182 VDD.n1604 VDD.t783 3.20383
R25183 VDD.t3395 VDD.n1605 3.20383
R25184 VDD.n1606 VDD.t3395 3.20383
R25185 VDD.t1522 VDD.n1607 3.20383
R25186 VDD.n1608 VDD.t1522 3.20383
R25187 VDD.n1496 VDD.t2406 3.20383
R25188 VDD.t2406 VDD.n1495 3.20383
R25189 VDD.n1593 VDD.t3924 3.20383
R25190 VDD.n1594 VDD.t3924 3.20383
R25191 VDD.n1595 VDD.t3506 3.20383
R25192 VDD.n1596 VDD.t3506 3.20383
R25193 VDD.n1597 VDD.t1941 3.20383
R25194 VDD.n1604 VDD.t4696 3.20383
R25195 VDD.n1605 VDD.t3220 3.20383
R25196 VDD.n1606 VDD.t3220 3.20383
R25197 VDD.n1607 VDD.t1308 3.20383
R25198 VDD.n1608 VDD.t1308 3.20383
R25199 VDD.n1496 VDD.t2110 3.20383
R25200 VDD.n1495 VDD.t2110 3.20383
R25201 VDD.n1528 VDD.t1624 3.20383
R25202 VDD.t1870 VDD.n1518 3.20383
R25203 VDD.n1517 VDD.t693 3.20383
R25204 VDD.t2429 VDD.n771 3.20383
R25205 VDD.n1555 VDD.t4773 3.20383
R25206 VDD.n1555 VDD.t4770 3.20383
R25207 VDD.n1556 VDD.t4775 3.20383
R25208 VDD.n1556 VDD.t4772 3.20383
R25209 VDD.n1557 VDD.t4774 3.20383
R25210 VDD.n1557 VDD.t4771 3.20383
R25211 VDD.n1541 VDD.t995 3.20383
R25212 VDD.n1537 VDD.t1189 3.20383
R25213 VDD.n1559 VDD.t4206 3.20383
R25214 VDD.n1563 VDD.t1666 3.20383
R25215 VDD.n1175 VDD.t1477 3.20383
R25216 VDD.t1477 VDD.n1174 3.20383
R25217 VDD.n1173 VDD.t4140 3.20383
R25218 VDD.t1684 VDD.n1166 3.20383
R25219 VDD.n1165 VDD.t1216 3.20383
R25220 VDD.t1216 VDD.n1164 3.20383
R25221 VDD.n1188 VDD.t4730 3.20383
R25222 VDD.t4730 VDD.n1187 3.20383
R25223 VDD.n1186 VDD.t1760 3.20383
R25224 VDD.t4566 VDD.n1179 3.20383
R25225 VDD.n1178 VDD.t1628 3.20383
R25226 VDD.t1628 VDD.n1177 3.20383
R25227 VDD.t3573 VDD.n1337 3.20383
R25228 VDD.n1338 VDD.t3573 3.20383
R25229 VDD.t3798 VDD.n1339 3.20383
R25230 VDD.n1307 VDD.t589 3.20383
R25231 VDD.n1306 VDD.t881 3.20383
R25232 VDD.t881 VDD.n1305 3.20383
R25233 VDD.t3118 VDD.n1660 3.20383
R25234 VDD.n1659 VDD.t2709 3.20383
R25235 VDD.t2709 VDD.n1658 3.20383
R25236 VDD.n1657 VDD.t1089 3.20383
R25237 VDD.n1316 VDD.t3848 3.20383
R25238 VDD.t2376 VDD.n1317 3.20383
R25239 VDD.n1318 VDD.t2376 3.20383
R25240 VDD.t1994 VDD.n1384 3.20383
R25241 VDD.n1385 VDD.t1994 3.20383
R25242 VDD.t4592 VDD.n1386 3.20383
R25243 VDD.n1075 VDD.t579 3.20383
R25244 VDD.n1074 VDD.t3286 3.20383
R25245 VDD.t3286 VDD.n1073 3.20383
R25246 VDD.n1286 VDD.t3812 3.20383
R25247 VDD.t3812 VDD.n1285 3.20383
R25248 VDD.n1284 VDD.t3668 3.20383
R25249 VDD.n1362 VDD.t889 3.20383
R25250 VDD.t3498 VDD.n1363 3.20383
R25251 VDD.n1364 VDD.t3498 3.20383
R25252 VDD.n1644 VDD.t2935 3.20383
R25253 VDD.t2136 VDD.n1645 3.20383
R25254 VDD.n1646 VDD.t2136 3.20383
R25255 VDD.t3342 VDD.n1647 3.20383
R25256 VDD.n1248 VDD.t3434 3.20383
R25257 VDD.t4598 VDD.n1249 3.20383
R25258 VDD.n1250 VDD.t4598 3.20383
R25259 VDD.n1735 VDD.t1151 3.20383
R25260 VDD.n1736 VDD.t1151 3.20383
R25261 VDD.n1737 VDD.t1286 3.20383
R25262 VDD.n948 VDD.t3599 3.20383
R25263 VDD.n950 VDD.t2620 3.20383
R25264 VDD.n951 VDD.t2620 3.20383
R25265 VDD.n71 VDD.n70 3.2012
R25266 VDD.n160 VDD.n159 3.2012
R25267 VDD.n5770 VDD.n5769 3.2012
R25268 VDD.n5837 VDD.n5836 3.2012
R25269 VDD.n5654 VDD.n5653 3.2012
R25270 VDD.n5572 VDD.n5571 3.2012
R25271 VDD.n8158 VDD.n8157 3.2012
R25272 VDD.n9115 VDD.n9114 3.2012
R25273 VDD.n8828 VDD.n8827 3.2012
R25274 VDD.n8968 VDD.n8967 3.2012
R25275 VDD.n5766 VDD.n5765 3.1154
R25276 VDD.n5833 VDD.n5832 3.1154
R25277 VDD.n5650 VDD.n5649 3.1154
R25278 VDD.n5568 VDD.n5567 3.1154
R25279 VDD.n8154 VDD.n8153 3.1154
R25280 VDD.n66 VDD.n65 3.11413
R25281 VDD.n155 VDD.n154 3.11413
R25282 VDD.n9110 VDD.n9109 3.11413
R25283 VDD.n8823 VDD.n8822 3.11413
R25284 VDD.n8963 VDD.n8962 3.11413
R25285 VDD.n6152 VDD.n6021 3.00663
R25286 VDD.n6095 VDD.n6094 3.00663
R25287 VDD.n6847 VDD.n6846 3.00663
R25288 VDD.n6797 VDD.n6796 3.00663
R25289 VDD.n1425 VDD.n1424 2.89741
R25290 VDD.n1418 VDD.n858 2.89677
R25291 VDD.n1679 VDD.n1678 2.89677
R25292 VDD.n1692 VDD.n1691 2.89677
R25293 VDD.n1626 VDD.n1625 2.89677
R25294 VDD.n1673 VDD.n1672 2.89677
R25295 VDD.n1619 VDD.n784 2.89677
R25296 VDD.n1106 VDD.n1091 2.89677
R25297 VDD.n1685 VDD.n1684 2.89677
R25298 VDD.n1697 VDD.n735 2.89677
R25299 VDD.n1045 VDD.n1039 2.89677
R25300 VDD.n979 VDD.n706 2.89677
R25301 VDD.n1086 VDD.n844 2.89406
R25302 VDD.n1419 VDD.n1418 2.89406
R25303 VDD.n1678 VDD.n1677 2.89406
R25304 VDD.n1690 VDD.n1689 2.89406
R25305 VDD.n1620 VDD.n1619 2.89406
R25306 VDD.n1106 VDD.n1105 2.89406
R25307 VDD.n1684 VDD.n1683 2.89406
R25308 VDD.n1697 VDD.n1696 2.89406
R25309 VDD.n1045 VDD.n1044 2.89406
R25310 VDD.n853 VDD.n706 2.89406
R25311 VDD.n984 VDD.n983 2.89406
R25312 VDD.n1034 VDD.n1033 2.89406
R25313 VDD.n6136 VDD.n6134 2.7866
R25314 VDD.n6139 VDD.n6137 2.7866
R25315 VDD.n6143 VDD.n6141 2.7866
R25316 VDD.n6147 VDD.n6145 2.7866
R25317 VDD.n6132 VDD.n6130 2.7866
R25318 VDD.n6128 VDD.n6126 2.7866
R25319 VDD.n6124 VDD.n6122 2.7866
R25320 VDD.n6120 VDD.n6118 2.7866
R25321 VDD.n6044 VDD.n6042 2.7866
R25322 VDD.n6047 VDD.n6045 2.7866
R25323 VDD.n6051 VDD.n6049 2.7866
R25324 VDD.n6055 VDD.n6053 2.7866
R25325 VDD.n6078 VDD.n6076 2.7866
R25326 VDD.n6082 VDD.n6080 2.7866
R25327 VDD.n6086 VDD.n6084 2.7866
R25328 VDD.n6090 VDD.n6088 2.7866
R25329 VDD.n6810 VDD.n6808 2.7866
R25330 VDD.n6813 VDD.n6811 2.7866
R25331 VDD.n6817 VDD.n6815 2.7866
R25332 VDD.n6821 VDD.n6819 2.7866
R25333 VDD.n6826 VDD.n6824 2.7866
R25334 VDD.n6830 VDD.n6828 2.7866
R25335 VDD.n6834 VDD.n6832 2.7866
R25336 VDD.n6838 VDD.n6836 2.7866
R25337 VDD.n6777 VDD.n6775 2.7866
R25338 VDD.n6780 VDD.n6778 2.7866
R25339 VDD.n6784 VDD.n6782 2.7866
R25340 VDD.n6788 VDD.n6786 2.7866
R25341 VDD.n6773 VDD.n6771 2.7866
R25342 VDD.n6769 VDD.n6767 2.7866
R25343 VDD.n6765 VDD.n6763 2.7866
R25344 VDD.n6761 VDD.n6759 2.7866
R25345 VDD.n7004 VDD.n7002 2.73714
R25346 VDD.n6926 VDD.n6924 2.73714
R25347 VDD.n6541 VDD.n6539 2.73714
R25348 VDD.n6452 VDD.n6450 2.73714
R25349 VDD.n6140 VDD.n6136 2.73672
R25350 VDD.n6048 VDD.n6044 2.73672
R25351 VDD.n6814 VDD.n6810 2.73672
R25352 VDD.n6781 VDD.n6777 2.73672
R25353 VDD.n58 VDD.n57 2.65954
R25354 VDD.n64 VDD.n63 2.65954
R25355 VDD.n147 VDD.n146 2.65954
R25356 VDD.n153 VDD.n152 2.65954
R25357 VDD.n9102 VDD.n9101 2.65954
R25358 VDD.n9108 VDD.n9107 2.65954
R25359 VDD.n8815 VDD.n8814 2.65954
R25360 VDD.n8821 VDD.n8820 2.65954
R25361 VDD.n8955 VDD.n8954 2.65954
R25362 VDD.n8961 VDD.n8960 2.65954
R25363 VDD.n5764 VDD.n5762 2.65924
R25364 VDD.n5757 VDD.n5756 2.65924
R25365 VDD.n5831 VDD.n5829 2.65924
R25366 VDD.n5824 VDD.n5823 2.65924
R25367 VDD.n5648 VDD.n5646 2.65924
R25368 VDD.n5641 VDD.n5640 2.65924
R25369 VDD.n5566 VDD.n5564 2.65924
R25370 VDD.n5559 VDD.n5558 2.65924
R25371 VDD.n8152 VDD.n8150 2.65924
R25372 VDD.n8145 VDD.n8144 2.65924
R25373 VDD.n5767 VDD.n5766 2.61766
R25374 VDD.n5834 VDD.n5833 2.61766
R25375 VDD.n5651 VDD.n5650 2.61766
R25376 VDD.n5569 VDD.n5568 2.61766
R25377 VDD.n8155 VDD.n8154 2.61766
R25378 VDD.n67 VDD.n66 2.61737
R25379 VDD.n156 VDD.n155 2.61737
R25380 VDD.n9111 VDD.n9110 2.61737
R25381 VDD.n8824 VDD.n8823 2.61737
R25382 VDD.n8964 VDD.n8963 2.61737
R25383 VDD.n8064 VDD.n8063 2.60496
R25384 VDD.n7959 VDD.n7958 2.60386
R25385 VDD.n8082 VDD.n8081 2.6005
R25386 VDD.n8083 VDD.n2120 2.6005
R25387 VDD.n8074 VDD.n8073 2.6005
R25388 VDD.n8072 VDD.n8071 2.6005
R25389 VDD.n8054 VDD.n8052 2.59852
R25390 VDD.n7949 VDD.n7947 2.59742
R25391 VDD.n6956 VDD.n6954 2.59712
R25392 VDD.n6924 VDD.n6922 2.59712
R25393 VDD.n7008 VDD.n7006 2.59712
R25394 VDD.n7002 VDD.n7000 2.59712
R25395 VDD.n6500 VDD.n6498 2.59712
R25396 VDD.n6450 VDD.n6448 2.59712
R25397 VDD.n6546 VDD.n6544 2.59712
R25398 VDD.n6539 VDD.n6537 2.59712
R25399 VDD.t3015 VDD.n1529 2.55028
R25400 VDD.t2298 VDD.n1542 2.55022
R25401 VDD.n772 VDD.t4521 2.54061
R25402 VDD.t4521 VDD.n770 2.54061
R25403 VDD.t4587 VDD.n1635 2.54061
R25404 VDD.n1636 VDD.t4587 2.54061
R25405 VDD.t1076 VDD.n1632 2.54061
R25406 VDD.n1633 VDD.t1076 2.54061
R25407 VDD.t919 VDD.n1629 2.54061
R25408 VDD.n1630 VDD.t919 2.54061
R25409 VDD.n1510 VDD.t3873 2.54061
R25410 VDD.t3873 VDD.n782 2.54061
R25411 VDD.n1530 VDD.t3015 2.54061
R25412 VDD.n1532 VDD.t3059 2.54061
R25413 VDD.t3059 VDD.n1531 2.54061
R25414 VDD.n1546 VDD.t3602 2.54061
R25415 VDD.t3602 VDD.n1533 2.54061
R25416 VDD.t3443 VDD.n1544 2.54061
R25417 VDD.n1545 VDD.t3443 2.54061
R25418 VDD.n1543 VDD.t2298 2.54061
R25419 VDD.n2142 VDD.t1024 2.5255
R25420 VDD.n2140 VDD.t2410 2.5255
R25421 VDD.n2137 VDD.t3326 2.5255
R25422 VDD.n2137 VDD.t2297 2.5255
R25423 VDD.n2135 VDD.t772 2.5255
R25424 VDD.n2135 VDD.t3870 2.5255
R25425 VDD.n2132 VDD.t3802 2.5255
R25426 VDD.n2132 VDD.t2845 2.5255
R25427 VDD.n2129 VDD.t1990 2.5255
R25428 VDD.n2129 VDD.t963 2.5255
R25429 VDD.n8067 VDD.t569 2.5255
R25430 VDD.n2147 VDD.t1911 2.5255
R25431 VDD.n2160 VDD.t1829 2.5255
R25432 VDD.n2164 VDD.t3474 2.5255
R25433 VDD.n8015 VDD.t2427 2.5255
R25434 VDD.n2121 VDD.t4686 2.5255
R25435 VDD.n7913 VDD.n7912 2.46986
R25436 VDD.n7909 VDD.n7908 2.46873
R25437 VDD.n8018 VDD.n8017 2.46873
R25438 VDD.n8047 VDD.n8046 2.46198
R25439 VDD.n7891 VDD.n7890 2.46198
R25440 VDD.n7942 VDD.n7941 2.46086
R25441 VDD.n7005 VDD.n7004 2.46014
R25442 VDD.n6958 VDD.n6926 2.46014
R25443 VDD.n6548 VDD.n6541 2.46014
R25444 VDD.n6497 VDD.n6452 2.46014
R25445 VDD.t2841 VDD.n8072 2.4505
R25446 VDD.n8072 VDD.t1359 2.4505
R25447 VDD.n8073 VDD.t942 2.4505
R25448 VDD.n8073 VDD.t2841 2.4505
R25449 VDD.n8083 VDD.t2770 2.4505
R25450 VDD.t1276 VDD.n8083 2.4505
R25451 VDD.n8082 VDD.t860 2.4505
R25452 VDD.t2770 VDD.n8082 2.4505
R25453 VDD.n6956 VDD.n6955 2.39107
R25454 VDD.n6924 VDD.n6923 2.39107
R25455 VDD.n7008 VDD.n7007 2.39107
R25456 VDD.n7002 VDD.n7001 2.39107
R25457 VDD.n6500 VDD.n6499 2.39107
R25458 VDD.n6450 VDD.n6449 2.39107
R25459 VDD.n6546 VDD.n6545 2.39107
R25460 VDD.n6539 VDD.n6538 2.39107
R25461 VDD.n6751 VDD.n6750 2.37568
R25462 VDD.n6064 VDD.n6063 2.37568
R25463 VDD.n6107 VDD.n6106 2.37568
R25464 VDD.n6733 VDD.n6732 2.37568
R25465 VDD.n7892 VDD.n7886 2.37449
R25466 VDD.n7895 VDD.n7882 2.37449
R25467 VDD.n7898 VDD.n7878 2.37449
R25468 VDD.n7904 VDD.n7872 2.37449
R25469 VDD.n7907 VDD.n7868 2.37449
R25470 VDD.n1448 VDD.n1447 2.30715
R25471 VDD.n7024 VDD.n2375 2.30165
R25472 VDD.n6877 VDD.n6876 2.30165
R25473 VDD.n6414 VDD.n6413 2.30165
R25474 VDD.n6561 VDD.n5288 2.30165
R25475 VDD.n5906 VDD.n5905 2.26828
R25476 VDD.n12582 VDD.n12560 2.26741
R25477 VDD.n6172 VDD.n6016 2.26689
R25478 VDD.n3630 VDD.n2745 2.2505
R25479 VDD.n3632 VDD.n3631 2.2505
R25480 VDD.n3633 VDD.n2744 2.2505
R25481 VDD.n3635 VDD.n3634 2.2505
R25482 VDD.n3636 VDD.n2743 2.2505
R25483 VDD.n3638 VDD.n3637 2.2505
R25484 VDD.n3639 VDD.n2742 2.2505
R25485 VDD.n3641 VDD.n3640 2.2505
R25486 VDD.n3642 VDD.n2741 2.2505
R25487 VDD.n3644 VDD.n3643 2.2505
R25488 VDD.n3645 VDD.n2740 2.2505
R25489 VDD.n3647 VDD.n3646 2.2505
R25490 VDD.n3648 VDD.n2739 2.2505
R25491 VDD.n3650 VDD.n3649 2.2505
R25492 VDD.n3651 VDD.n2738 2.2505
R25493 VDD.n3653 VDD.n3652 2.2505
R25494 VDD.n3654 VDD.n2737 2.2505
R25495 VDD.n3656 VDD.n3655 2.2505
R25496 VDD.n3657 VDD.n2736 2.2505
R25497 VDD.n3659 VDD.n3658 2.2505
R25498 VDD.n3660 VDD.n2735 2.2505
R25499 VDD.n3662 VDD.n3661 2.2505
R25500 VDD.n3663 VDD.n2734 2.2505
R25501 VDD.n3665 VDD.n3664 2.2505
R25502 VDD.n3666 VDD.n2733 2.2505
R25503 VDD.n3668 VDD.n3667 2.2505
R25504 VDD.n3669 VDD.n2732 2.2505
R25505 VDD.n3671 VDD.n3670 2.2505
R25506 VDD.n3672 VDD.n2731 2.2505
R25507 VDD.n3674 VDD.n3673 2.2505
R25508 VDD.n3675 VDD.n2730 2.2505
R25509 VDD.n3677 VDD.n3676 2.2505
R25510 VDD.n3678 VDD.n2729 2.2505
R25511 VDD.n3680 VDD.n3679 2.2505
R25512 VDD.n3681 VDD.n2728 2.2505
R25513 VDD.n3683 VDD.n3682 2.2505
R25514 VDD.n3684 VDD.n2727 2.2505
R25515 VDD.n3686 VDD.n3685 2.2505
R25516 VDD.n3687 VDD.n2726 2.2505
R25517 VDD.n3689 VDD.n3688 2.2505
R25518 VDD.n3690 VDD.n2725 2.2505
R25519 VDD.n3692 VDD.n3691 2.2505
R25520 VDD.n3693 VDD.n2724 2.2505
R25521 VDD.n3695 VDD.n3694 2.2505
R25522 VDD.n3696 VDD.n2723 2.2505
R25523 VDD.n3698 VDD.n3697 2.2505
R25524 VDD.n3699 VDD.n2722 2.2505
R25525 VDD.n3701 VDD.n3700 2.2505
R25526 VDD.n3702 VDD.n2721 2.2505
R25527 VDD.n3704 VDD.n3703 2.2505
R25528 VDD.n3705 VDD.n2720 2.2505
R25529 VDD.n3707 VDD.n3706 2.2505
R25530 VDD.n3708 VDD.n2719 2.2505
R25531 VDD.n3710 VDD.n3709 2.2505
R25532 VDD.n3711 VDD.n2718 2.2505
R25533 VDD.n3713 VDD.n3712 2.2505
R25534 VDD.n3714 VDD.n2717 2.2505
R25535 VDD.n3716 VDD.n3715 2.2505
R25536 VDD.n3717 VDD.n2716 2.2505
R25537 VDD.n3719 VDD.n3718 2.2505
R25538 VDD.n3720 VDD.n2715 2.2505
R25539 VDD.n3722 VDD.n3721 2.2505
R25540 VDD.n3723 VDD.n2714 2.2505
R25541 VDD.n3725 VDD.n3724 2.2505
R25542 VDD.n3726 VDD.n2713 2.2505
R25543 VDD.n3728 VDD.n3727 2.2505
R25544 VDD.n3729 VDD.n2712 2.2505
R25545 VDD.n3731 VDD.n3730 2.2505
R25546 VDD.n3732 VDD.n2711 2.2505
R25547 VDD.n3734 VDD.n3733 2.2505
R25548 VDD.n3735 VDD.n2710 2.2505
R25549 VDD.n3737 VDD.n3736 2.2505
R25550 VDD.n3738 VDD.n2709 2.2505
R25551 VDD.n3740 VDD.n3739 2.2505
R25552 VDD.n3741 VDD.n2708 2.2505
R25553 VDD.n3743 VDD.n3742 2.2505
R25554 VDD.n3744 VDD.n2707 2.2505
R25555 VDD.n3746 VDD.n3745 2.2505
R25556 VDD.n3747 VDD.n2706 2.2505
R25557 VDD.n3749 VDD.n3748 2.2505
R25558 VDD.n3750 VDD.n2705 2.2505
R25559 VDD.n3752 VDD.n3751 2.2505
R25560 VDD.n3753 VDD.n2704 2.2505
R25561 VDD.n3755 VDD.n3754 2.2505
R25562 VDD.n3756 VDD.n2703 2.2505
R25563 VDD.n3758 VDD.n3757 2.2505
R25564 VDD.n3759 VDD.n2702 2.2505
R25565 VDD.n3761 VDD.n3760 2.2505
R25566 VDD.n3762 VDD.n2701 2.2505
R25567 VDD.n3764 VDD.n3763 2.2505
R25568 VDD.n3765 VDD.n2700 2.2505
R25569 VDD.n3767 VDD.n3766 2.2505
R25570 VDD.n3768 VDD.n2699 2.2505
R25571 VDD.n3770 VDD.n3769 2.2505
R25572 VDD.n3771 VDD.n2698 2.2505
R25573 VDD.n3773 VDD.n3772 2.2505
R25574 VDD.n3774 VDD.n2697 2.2505
R25575 VDD.n3776 VDD.n3775 2.2505
R25576 VDD.n3777 VDD.n2696 2.2505
R25577 VDD.n3779 VDD.n3778 2.2505
R25578 VDD.n3780 VDD.n2695 2.2505
R25579 VDD.n3782 VDD.n3781 2.2505
R25580 VDD.n3783 VDD.n2694 2.2505
R25581 VDD.n3785 VDD.n3784 2.2505
R25582 VDD.n3786 VDD.n2693 2.2505
R25583 VDD.n3788 VDD.n3787 2.2505
R25584 VDD.n3789 VDD.n2692 2.2505
R25585 VDD.n3791 VDD.n3790 2.2505
R25586 VDD.n3792 VDD.n2691 2.2505
R25587 VDD.n3794 VDD.n3793 2.2505
R25588 VDD.n3795 VDD.n2690 2.2505
R25589 VDD.n3797 VDD.n3796 2.2505
R25590 VDD.n3798 VDD.n2689 2.2505
R25591 VDD.n3800 VDD.n3799 2.2505
R25592 VDD.n3801 VDD.n2688 2.2505
R25593 VDD.n3803 VDD.n3802 2.2505
R25594 VDD.n3804 VDD.n2687 2.2505
R25595 VDD.n3806 VDD.n3805 2.2505
R25596 VDD.n3807 VDD.n2686 2.2505
R25597 VDD.n3809 VDD.n3808 2.2505
R25598 VDD.n3810 VDD.n2685 2.2505
R25599 VDD.n3812 VDD.n3811 2.2505
R25600 VDD.n3813 VDD.n2684 2.2505
R25601 VDD.n3815 VDD.n3814 2.2505
R25602 VDD.n3816 VDD.n2683 2.2505
R25603 VDD.n3818 VDD.n3817 2.2505
R25604 VDD.n3819 VDD.n2682 2.2505
R25605 VDD.n3821 VDD.n3820 2.2505
R25606 VDD.n3822 VDD.n2681 2.2505
R25607 VDD.n3824 VDD.n3823 2.2505
R25608 VDD.n3825 VDD.n2680 2.2505
R25609 VDD.n3827 VDD.n3826 2.2505
R25610 VDD.n3828 VDD.n2679 2.2505
R25611 VDD.n3830 VDD.n3829 2.2505
R25612 VDD.n3831 VDD.n2678 2.2505
R25613 VDD.n3833 VDD.n3832 2.2505
R25614 VDD.n3834 VDD.n2677 2.2505
R25615 VDD.n3836 VDD.n3835 2.2505
R25616 VDD.n3837 VDD.n2676 2.2505
R25617 VDD.n3839 VDD.n3838 2.2505
R25618 VDD.n3840 VDD.n2675 2.2505
R25619 VDD.n3842 VDD.n3841 2.2505
R25620 VDD.n3843 VDD.n2674 2.2505
R25621 VDD.n3845 VDD.n3844 2.2505
R25622 VDD.n3846 VDD.n2673 2.2505
R25623 VDD.n3848 VDD.n3847 2.2505
R25624 VDD.n3849 VDD.n2672 2.2505
R25625 VDD.n3851 VDD.n3850 2.2505
R25626 VDD.n3852 VDD.n2671 2.2505
R25627 VDD.n3854 VDD.n3853 2.2505
R25628 VDD.n3855 VDD.n2670 2.2505
R25629 VDD.n3857 VDD.n3856 2.2505
R25630 VDD.n3858 VDD.n2669 2.2505
R25631 VDD.n3860 VDD.n3859 2.2505
R25632 VDD.n3861 VDD.n2668 2.2505
R25633 VDD.n3863 VDD.n3862 2.2505
R25634 VDD.n3864 VDD.n2667 2.2505
R25635 VDD.n3866 VDD.n3865 2.2505
R25636 VDD.n3867 VDD.n2666 2.2505
R25637 VDD.n3869 VDD.n3868 2.2505
R25638 VDD.n3870 VDD.n2665 2.2505
R25639 VDD.n3872 VDD.n3871 2.2505
R25640 VDD.n3873 VDD.n2664 2.2505
R25641 VDD.n3875 VDD.n3874 2.2505
R25642 VDD.n3876 VDD.n2663 2.2505
R25643 VDD.n3878 VDD.n3877 2.2505
R25644 VDD.n3879 VDD.n2662 2.2505
R25645 VDD.n3881 VDD.n3880 2.2505
R25646 VDD.n3882 VDD.n2661 2.2505
R25647 VDD.n3884 VDD.n3883 2.2505
R25648 VDD.n3885 VDD.n2660 2.2505
R25649 VDD.n3887 VDD.n3886 2.2505
R25650 VDD.n3888 VDD.n2659 2.2505
R25651 VDD.n3890 VDD.n3889 2.2505
R25652 VDD.n3891 VDD.n2658 2.2505
R25653 VDD.n3893 VDD.n3892 2.2505
R25654 VDD.n3894 VDD.n2657 2.2505
R25655 VDD.n3896 VDD.n3895 2.2505
R25656 VDD.n3897 VDD.n2656 2.2505
R25657 VDD.n3899 VDD.n3898 2.2505
R25658 VDD.n3900 VDD.n2655 2.2505
R25659 VDD.n3902 VDD.n3901 2.2505
R25660 VDD.n3903 VDD.n2654 2.2505
R25661 VDD.n3905 VDD.n3904 2.2505
R25662 VDD.n3906 VDD.n2653 2.2505
R25663 VDD.n3908 VDD.n3907 2.2505
R25664 VDD.n3909 VDD.n2652 2.2505
R25665 VDD.n3911 VDD.n3910 2.2505
R25666 VDD.n3912 VDD.n2651 2.2505
R25667 VDD.n3914 VDD.n3913 2.2505
R25668 VDD.n3915 VDD.n2650 2.2505
R25669 VDD.n3917 VDD.n3916 2.2505
R25670 VDD.n3918 VDD.n2649 2.2505
R25671 VDD.n3920 VDD.n3919 2.2505
R25672 VDD.n3921 VDD.n2648 2.2505
R25673 VDD.n3923 VDD.n3922 2.2505
R25674 VDD.n3924 VDD.n2647 2.2505
R25675 VDD.n3926 VDD.n3925 2.2505
R25676 VDD.n3927 VDD.n2646 2.2505
R25677 VDD.n3929 VDD.n3928 2.2505
R25678 VDD.n3930 VDD.n2645 2.2505
R25679 VDD.n3932 VDD.n3931 2.2505
R25680 VDD.n3933 VDD.n2644 2.2505
R25681 VDD.n3935 VDD.n3934 2.2505
R25682 VDD.n3936 VDD.n2643 2.2505
R25683 VDD.n3938 VDD.n3937 2.2505
R25684 VDD.n3939 VDD.n2642 2.2505
R25685 VDD.n3941 VDD.n3940 2.2505
R25686 VDD.n3942 VDD.n2641 2.2505
R25687 VDD.n3944 VDD.n3943 2.2505
R25688 VDD.n3945 VDD.n2640 2.2505
R25689 VDD.n3947 VDD.n3946 2.2505
R25690 VDD.n3948 VDD.n2639 2.2505
R25691 VDD.n3950 VDD.n3949 2.2505
R25692 VDD.n3951 VDD.n2638 2.2505
R25693 VDD.n3953 VDD.n3952 2.2505
R25694 VDD.n3954 VDD.n2637 2.2505
R25695 VDD.n3956 VDD.n3955 2.2505
R25696 VDD.n3957 VDD.n2636 2.2505
R25697 VDD.n3959 VDD.n3958 2.2505
R25698 VDD.n3960 VDD.n2635 2.2505
R25699 VDD.n3962 VDD.n3961 2.2505
R25700 VDD.n3963 VDD.n2634 2.2505
R25701 VDD.n3965 VDD.n3964 2.2505
R25702 VDD.n3966 VDD.n2633 2.2505
R25703 VDD.n3968 VDD.n3967 2.2505
R25704 VDD.n3969 VDD.n2632 2.2505
R25705 VDD.n3971 VDD.n3970 2.2505
R25706 VDD.n3972 VDD.n2631 2.2505
R25707 VDD.n3974 VDD.n3973 2.2505
R25708 VDD.n3975 VDD.n2630 2.2505
R25709 VDD.n3977 VDD.n3976 2.2505
R25710 VDD.n3978 VDD.n2629 2.2505
R25711 VDD.n3980 VDD.n3979 2.2505
R25712 VDD.n3981 VDD.n2628 2.2505
R25713 VDD.n3983 VDD.n3982 2.2505
R25714 VDD.n3984 VDD.n2627 2.2505
R25715 VDD.n3986 VDD.n3985 2.2505
R25716 VDD.n3987 VDD.n2626 2.2505
R25717 VDD.n3989 VDD.n3988 2.2505
R25718 VDD.n3990 VDD.n2625 2.2505
R25719 VDD.n3992 VDD.n3991 2.2505
R25720 VDD.n3993 VDD.n2624 2.2505
R25721 VDD.n3995 VDD.n3994 2.2505
R25722 VDD.n3996 VDD.n2623 2.2505
R25723 VDD.n3998 VDD.n3997 2.2505
R25724 VDD.n3999 VDD.n2622 2.2505
R25725 VDD.n4001 VDD.n4000 2.2505
R25726 VDD.n4002 VDD.n2621 2.2505
R25727 VDD.n4004 VDD.n4003 2.2505
R25728 VDD.n4005 VDD.n2620 2.2505
R25729 VDD.n4007 VDD.n4006 2.2505
R25730 VDD.n4008 VDD.n2619 2.2505
R25731 VDD.n4010 VDD.n4009 2.2505
R25732 VDD.n4011 VDD.n2618 2.2505
R25733 VDD.n4013 VDD.n4012 2.2505
R25734 VDD.n4014 VDD.n2617 2.2505
R25735 VDD.n4016 VDD.n4015 2.2505
R25736 VDD.n4017 VDD.n2616 2.2505
R25737 VDD.n4019 VDD.n4018 2.2505
R25738 VDD.n4020 VDD.n2615 2.2505
R25739 VDD.n4022 VDD.n4021 2.2505
R25740 VDD.n4023 VDD.n2614 2.2505
R25741 VDD.n4025 VDD.n4024 2.2505
R25742 VDD.n4026 VDD.n2613 2.2505
R25743 VDD.n4028 VDD.n4027 2.2505
R25744 VDD.n4029 VDD.n2612 2.2505
R25745 VDD.n4031 VDD.n4030 2.2505
R25746 VDD.n4032 VDD.n2611 2.2505
R25747 VDD.n4034 VDD.n4033 2.2505
R25748 VDD.n4035 VDD.n2610 2.2505
R25749 VDD.n4037 VDD.n4036 2.2505
R25750 VDD.n4038 VDD.n2609 2.2505
R25751 VDD.n4040 VDD.n4039 2.2505
R25752 VDD.n4041 VDD.n2608 2.2505
R25753 VDD.n4043 VDD.n4042 2.2505
R25754 VDD.n4044 VDD.n2607 2.2505
R25755 VDD.n4046 VDD.n4045 2.2505
R25756 VDD.n4047 VDD.n2606 2.2505
R25757 VDD.n4049 VDD.n4048 2.2505
R25758 VDD.n4050 VDD.n2605 2.2505
R25759 VDD.n4052 VDD.n4051 2.2505
R25760 VDD.n4053 VDD.n2604 2.2505
R25761 VDD.n4055 VDD.n4054 2.2505
R25762 VDD.n4056 VDD.n2603 2.2505
R25763 VDD.n4058 VDD.n4057 2.2505
R25764 VDD.n4059 VDD.n2602 2.2505
R25765 VDD.n4061 VDD.n4060 2.2505
R25766 VDD.n4062 VDD.n2601 2.2505
R25767 VDD.n4064 VDD.n4063 2.2505
R25768 VDD.n4065 VDD.n2600 2.2505
R25769 VDD.n4067 VDD.n4066 2.2505
R25770 VDD.n4068 VDD.n2599 2.2505
R25771 VDD.n4070 VDD.n4069 2.2505
R25772 VDD.n4071 VDD.n2598 2.2505
R25773 VDD.n4073 VDD.n4072 2.2505
R25774 VDD.n4074 VDD.n2597 2.2505
R25775 VDD.n4076 VDD.n4075 2.2505
R25776 VDD.n4077 VDD.n2596 2.2505
R25777 VDD.n4079 VDD.n4078 2.2505
R25778 VDD.n4080 VDD.n2595 2.2505
R25779 VDD.n4082 VDD.n4081 2.2505
R25780 VDD.n4083 VDD.n2594 2.2505
R25781 VDD.n4085 VDD.n4084 2.2505
R25782 VDD.n4086 VDD.n2593 2.2505
R25783 VDD.n4088 VDD.n4087 2.2505
R25784 VDD.n4089 VDD.n2592 2.2505
R25785 VDD.n4091 VDD.n4090 2.2505
R25786 VDD.n4092 VDD.n2591 2.2505
R25787 VDD.n4094 VDD.n4093 2.2505
R25788 VDD.n4095 VDD.n2590 2.2505
R25789 VDD.n4097 VDD.n4096 2.2505
R25790 VDD.n4098 VDD.n2589 2.2505
R25791 VDD.n4100 VDD.n4099 2.2505
R25792 VDD.n4101 VDD.n2588 2.2505
R25793 VDD.n4103 VDD.n4102 2.2505
R25794 VDD.n4104 VDD.n2587 2.2505
R25795 VDD.n4106 VDD.n4105 2.2505
R25796 VDD.n4107 VDD.n2586 2.2505
R25797 VDD.n4109 VDD.n4108 2.2505
R25798 VDD.n4110 VDD.n2585 2.2505
R25799 VDD.n4112 VDD.n4111 2.2505
R25800 VDD.n4113 VDD.n2584 2.2505
R25801 VDD.n4115 VDD.n4114 2.2505
R25802 VDD.n4116 VDD.n2583 2.2505
R25803 VDD.n4118 VDD.n4117 2.2505
R25804 VDD.n4119 VDD.n2582 2.2505
R25805 VDD.n4121 VDD.n4120 2.2505
R25806 VDD.n4122 VDD.n2581 2.2505
R25807 VDD.n4124 VDD.n4123 2.2505
R25808 VDD.n4125 VDD.n2580 2.2505
R25809 VDD.n4127 VDD.n4126 2.2505
R25810 VDD.n4128 VDD.n2579 2.2505
R25811 VDD.n4130 VDD.n4129 2.2505
R25812 VDD.n4131 VDD.n2578 2.2505
R25813 VDD.n4133 VDD.n4132 2.2505
R25814 VDD.n4134 VDD.n2577 2.2505
R25815 VDD.n4136 VDD.n4135 2.2505
R25816 VDD.n4137 VDD.n2576 2.2505
R25817 VDD.n4139 VDD.n4138 2.2505
R25818 VDD.n4140 VDD.n2575 2.2505
R25819 VDD.n4142 VDD.n4141 2.2505
R25820 VDD.n4143 VDD.n2574 2.2505
R25821 VDD.n4145 VDD.n4144 2.2505
R25822 VDD.n4146 VDD.n2573 2.2505
R25823 VDD.n4148 VDD.n4147 2.2505
R25824 VDD.n4149 VDD.n2572 2.2505
R25825 VDD.n4151 VDD.n4150 2.2505
R25826 VDD.n4152 VDD.n2571 2.2505
R25827 VDD.n4154 VDD.n4153 2.2505
R25828 VDD.n4155 VDD.n2570 2.2505
R25829 VDD.n4157 VDD.n4156 2.2505
R25830 VDD.n4158 VDD.n2569 2.2505
R25831 VDD.n4160 VDD.n4159 2.2505
R25832 VDD.n4161 VDD.n2568 2.2505
R25833 VDD.n4163 VDD.n4162 2.2505
R25834 VDD.n4164 VDD.n2567 2.2505
R25835 VDD.n4166 VDD.n4165 2.2505
R25836 VDD.n4167 VDD.n2566 2.2505
R25837 VDD.n4169 VDD.n4168 2.2505
R25838 VDD.n4170 VDD.n2565 2.2505
R25839 VDD.n4172 VDD.n4171 2.2505
R25840 VDD.n4173 VDD.n2564 2.2505
R25841 VDD.n4175 VDD.n4174 2.2505
R25842 VDD.n4176 VDD.n2563 2.2505
R25843 VDD.n4178 VDD.n4177 2.2505
R25844 VDD.n4179 VDD.n2562 2.2505
R25845 VDD.n4181 VDD.n4180 2.2505
R25846 VDD.n4182 VDD.n2561 2.2505
R25847 VDD.n4184 VDD.n4183 2.2505
R25848 VDD.n4185 VDD.n2560 2.2505
R25849 VDD.n4187 VDD.n4186 2.2505
R25850 VDD.n4188 VDD.n2559 2.2505
R25851 VDD.n4190 VDD.n4189 2.2505
R25852 VDD.n4191 VDD.n2558 2.2505
R25853 VDD.n4193 VDD.n4192 2.2505
R25854 VDD.n4194 VDD.n2557 2.2505
R25855 VDD.n4196 VDD.n4195 2.2505
R25856 VDD.n4197 VDD.n2556 2.2505
R25857 VDD.n4199 VDD.n4198 2.2505
R25858 VDD.n4200 VDD.n2555 2.2505
R25859 VDD.n4202 VDD.n4201 2.2505
R25860 VDD.n4203 VDD.n2554 2.2505
R25861 VDD.n4205 VDD.n4204 2.2505
R25862 VDD.n4206 VDD.n2553 2.2505
R25863 VDD.n4208 VDD.n4207 2.2505
R25864 VDD.n4209 VDD.n2552 2.2505
R25865 VDD.n4211 VDD.n4210 2.2505
R25866 VDD.n4212 VDD.n2551 2.2505
R25867 VDD.n4214 VDD.n4213 2.2505
R25868 VDD.n4215 VDD.n2550 2.2505
R25869 VDD.n4217 VDD.n4216 2.2505
R25870 VDD.n4218 VDD.n2549 2.2505
R25871 VDD.n4220 VDD.n4219 2.2505
R25872 VDD.n4221 VDD.n2548 2.2505
R25873 VDD.n4223 VDD.n4222 2.2505
R25874 VDD.n4224 VDD.n2547 2.2505
R25875 VDD.n4226 VDD.n4225 2.2505
R25876 VDD.n4227 VDD.n2546 2.2505
R25877 VDD.n4229 VDD.n4228 2.2505
R25878 VDD.n4230 VDD.n2545 2.2505
R25879 VDD.n4232 VDD.n4231 2.2505
R25880 VDD.n4233 VDD.n2544 2.2505
R25881 VDD.n4235 VDD.n4234 2.2505
R25882 VDD.n4236 VDD.n2543 2.2505
R25883 VDD.n4238 VDD.n4237 2.2505
R25884 VDD.n4239 VDD.n2542 2.2505
R25885 VDD.n4241 VDD.n4240 2.2505
R25886 VDD.n4242 VDD.n2541 2.2505
R25887 VDD.n4244 VDD.n4243 2.2505
R25888 VDD.n4245 VDD.n2540 2.2505
R25889 VDD.n4247 VDD.n4246 2.2505
R25890 VDD.n4248 VDD.n2539 2.2505
R25891 VDD.n4250 VDD.n4249 2.2505
R25892 VDD.n4251 VDD.n2538 2.2505
R25893 VDD.n4253 VDD.n4252 2.2505
R25894 VDD.n4254 VDD.n2537 2.2505
R25895 VDD.n4256 VDD.n4255 2.2505
R25896 VDD.n4257 VDD.n2536 2.2505
R25897 VDD.n4259 VDD.n4258 2.2505
R25898 VDD.n4260 VDD.n2535 2.2505
R25899 VDD.n4262 VDD.n4261 2.2505
R25900 VDD.n4263 VDD.n2534 2.2505
R25901 VDD.n4265 VDD.n4264 2.2505
R25902 VDD.n4266 VDD.n2533 2.2505
R25903 VDD.n4268 VDD.n4267 2.2505
R25904 VDD.n4269 VDD.n2532 2.2505
R25905 VDD.n4271 VDD.n4270 2.2505
R25906 VDD.n4272 VDD.n2531 2.2505
R25907 VDD.n4274 VDD.n4273 2.2505
R25908 VDD.n4275 VDD.n2530 2.2505
R25909 VDD.n4277 VDD.n4276 2.2505
R25910 VDD.n4278 VDD.n2529 2.2505
R25911 VDD.n4280 VDD.n4279 2.2505
R25912 VDD.n4281 VDD.n2528 2.2505
R25913 VDD.n4283 VDD.n4282 2.2505
R25914 VDD.n4284 VDD.n2527 2.2505
R25915 VDD.n4286 VDD.n4285 2.2505
R25916 VDD.n4287 VDD.n2526 2.2505
R25917 VDD.n4289 VDD.n4288 2.2505
R25918 VDD.n4290 VDD.n2525 2.2505
R25919 VDD.n4292 VDD.n4291 2.2505
R25920 VDD.n4293 VDD.n2524 2.2505
R25921 VDD.n4295 VDD.n4294 2.2505
R25922 VDD.n4296 VDD.n2523 2.2505
R25923 VDD.n4298 VDD.n4297 2.2505
R25924 VDD.n4299 VDD.n2522 2.2505
R25925 VDD.n4301 VDD.n4300 2.2505
R25926 VDD.n4302 VDD.n2521 2.2505
R25927 VDD.n4304 VDD.n4303 2.2505
R25928 VDD.n4305 VDD.n2520 2.2505
R25929 VDD.n4307 VDD.n4306 2.2505
R25930 VDD.n4308 VDD.n2519 2.2505
R25931 VDD.n4310 VDD.n4309 2.2505
R25932 VDD.n4311 VDD.n2518 2.2505
R25933 VDD.n4313 VDD.n4312 2.2505
R25934 VDD.n4314 VDD.n2517 2.2505
R25935 VDD.n4316 VDD.n4315 2.2505
R25936 VDD.n4317 VDD.n2516 2.2505
R25937 VDD.n4319 VDD.n4318 2.2505
R25938 VDD.n4320 VDD.n2515 2.2505
R25939 VDD.n4322 VDD.n4321 2.2505
R25940 VDD.n4323 VDD.n2514 2.2505
R25941 VDD.n4325 VDD.n4324 2.2505
R25942 VDD.n4326 VDD.n2513 2.2505
R25943 VDD.n4328 VDD.n4327 2.2505
R25944 VDD.n4329 VDD.n2512 2.2505
R25945 VDD.n4331 VDD.n4330 2.2505
R25946 VDD.n4332 VDD.n2511 2.2505
R25947 VDD.n4334 VDD.n4333 2.2505
R25948 VDD.n4335 VDD.n2510 2.2505
R25949 VDD.n4337 VDD.n4336 2.2505
R25950 VDD.n4338 VDD.n2509 2.2505
R25951 VDD.n4340 VDD.n4339 2.2505
R25952 VDD.n4341 VDD.n2508 2.2505
R25953 VDD.n4343 VDD.n4342 2.2505
R25954 VDD.n4344 VDD.n2507 2.2505
R25955 VDD.n4346 VDD.n4345 2.2505
R25956 VDD.n4347 VDD.n2506 2.2505
R25957 VDD.n4349 VDD.n4348 2.2505
R25958 VDD.n4350 VDD.n2505 2.2505
R25959 VDD.n4352 VDD.n4351 2.2505
R25960 VDD.n4353 VDD.n2504 2.2505
R25961 VDD.n4355 VDD.n4354 2.2505
R25962 VDD.n4356 VDD.n2503 2.2505
R25963 VDD.n4358 VDD.n4357 2.2505
R25964 VDD.n4359 VDD.n2502 2.2505
R25965 VDD.n4361 VDD.n4360 2.2505
R25966 VDD.n4362 VDD.n2501 2.2505
R25967 VDD.n4364 VDD.n4363 2.2505
R25968 VDD.n4365 VDD.n2500 2.2505
R25969 VDD.n4367 VDD.n4366 2.2505
R25970 VDD.n4368 VDD.n2499 2.2505
R25971 VDD.n4370 VDD.n4369 2.2505
R25972 VDD.n4371 VDD.n2498 2.2505
R25973 VDD.n4373 VDD.n4372 2.2505
R25974 VDD.n4374 VDD.n2497 2.2505
R25975 VDD.n4376 VDD.n4375 2.2505
R25976 VDD.n4377 VDD.n2496 2.2505
R25977 VDD.n4379 VDD.n4378 2.2505
R25978 VDD.n4380 VDD.n2495 2.2505
R25979 VDD.n4382 VDD.n4381 2.2505
R25980 VDD.n4383 VDD.n2494 2.2505
R25981 VDD.n4385 VDD.n4384 2.2505
R25982 VDD.n4386 VDD.n2493 2.2505
R25983 VDD.n4388 VDD.n4387 2.2505
R25984 VDD.n4389 VDD.n2492 2.2505
R25985 VDD.n4391 VDD.n4390 2.2505
R25986 VDD.n4392 VDD.n2491 2.2505
R25987 VDD.n4394 VDD.n4393 2.2505
R25988 VDD.n4395 VDD.n2490 2.2505
R25989 VDD.n4397 VDD.n4396 2.2505
R25990 VDD.n4398 VDD.n2489 2.2505
R25991 VDD.n4400 VDD.n4399 2.2505
R25992 VDD.n4401 VDD.n2488 2.2505
R25993 VDD.n4403 VDD.n4402 2.2505
R25994 VDD.n4404 VDD.n2487 2.2505
R25995 VDD.n4406 VDD.n4405 2.2505
R25996 VDD.n4407 VDD.n2486 2.2505
R25997 VDD.n4409 VDD.n4408 2.2505
R25998 VDD.n4410 VDD.n2485 2.2505
R25999 VDD.n4412 VDD.n4411 2.2505
R26000 VDD.n4413 VDD.n2484 2.2505
R26001 VDD.n4415 VDD.n4414 2.2505
R26002 VDD.n4416 VDD.n2483 2.2505
R26003 VDD.n4418 VDD.n4417 2.2505
R26004 VDD.n4419 VDD.n2482 2.2505
R26005 VDD.n4421 VDD.n4420 2.2505
R26006 VDD.n4422 VDD.n2481 2.2505
R26007 VDD.n4424 VDD.n4423 2.2505
R26008 VDD.n4425 VDD.n2480 2.2505
R26009 VDD.n4427 VDD.n4426 2.2505
R26010 VDD.n4428 VDD.n2479 2.2505
R26011 VDD.n4430 VDD.n4429 2.2505
R26012 VDD.n4431 VDD.n2478 2.2505
R26013 VDD.n4433 VDD.n4432 2.2505
R26014 VDD.n4434 VDD.n2477 2.2505
R26015 VDD.n4436 VDD.n4435 2.2505
R26016 VDD.n4437 VDD.n2476 2.2505
R26017 VDD.n4439 VDD.n4438 2.2505
R26018 VDD.n4440 VDD.n2475 2.2505
R26019 VDD.n4442 VDD.n4441 2.2505
R26020 VDD.n4443 VDD.n2474 2.2505
R26021 VDD.n4445 VDD.n4444 2.2505
R26022 VDD.n4446 VDD.n2473 2.2505
R26023 VDD.n4448 VDD.n4447 2.2505
R26024 VDD.n4449 VDD.n2472 2.2505
R26025 VDD.n4451 VDD.n4450 2.2505
R26026 VDD.n4452 VDD.n2471 2.2505
R26027 VDD.n4454 VDD.n4453 2.2505
R26028 VDD.n4455 VDD.n2470 2.2505
R26029 VDD.n4457 VDD.n4456 2.2505
R26030 VDD.n4458 VDD.n2469 2.2505
R26031 VDD.n4460 VDD.n4459 2.2505
R26032 VDD.n4461 VDD.n2468 2.2505
R26033 VDD.n4463 VDD.n4462 2.2505
R26034 VDD.n4464 VDD.n2467 2.2505
R26035 VDD.n4466 VDD.n4465 2.2505
R26036 VDD.n4467 VDD.n2466 2.2505
R26037 VDD.n4469 VDD.n4468 2.2505
R26038 VDD.n4470 VDD.n2465 2.2505
R26039 VDD.n4472 VDD.n4471 2.2505
R26040 VDD.n4473 VDD.n2464 2.2505
R26041 VDD.n4475 VDD.n4474 2.2505
R26042 VDD.n4476 VDD.n2463 2.2505
R26043 VDD.n4478 VDD.n4477 2.2505
R26044 VDD.n4479 VDD.n2462 2.2505
R26045 VDD.n4481 VDD.n4480 2.2505
R26046 VDD.n4482 VDD.n2461 2.2505
R26047 VDD.n4484 VDD.n4483 2.2505
R26048 VDD.n4485 VDD.n2460 2.2505
R26049 VDD.n4487 VDD.n4486 2.2505
R26050 VDD.n4488 VDD.n2459 2.2505
R26051 VDD.n4490 VDD.n4489 2.2505
R26052 VDD.n4491 VDD.n2458 2.2505
R26053 VDD.n4493 VDD.n4492 2.2505
R26054 VDD.n4494 VDD.n2457 2.2505
R26055 VDD.n4496 VDD.n4495 2.2505
R26056 VDD.n4497 VDD.n2456 2.2505
R26057 VDD.n4499 VDD.n4498 2.2505
R26058 VDD.n4500 VDD.n2455 2.2505
R26059 VDD.n4502 VDD.n4501 2.2505
R26060 VDD.n4503 VDD.n2454 2.2505
R26061 VDD.n4505 VDD.n4504 2.2505
R26062 VDD.n4506 VDD.n2453 2.2505
R26063 VDD.n4508 VDD.n4507 2.2505
R26064 VDD.n4509 VDD.n2452 2.2505
R26065 VDD.n4511 VDD.n4510 2.2505
R26066 VDD.n4512 VDD.n2451 2.2505
R26067 VDD.n4514 VDD.n4513 2.2505
R26068 VDD.n4515 VDD.n2450 2.2505
R26069 VDD.n4517 VDD.n4516 2.2505
R26070 VDD.n4518 VDD.n2449 2.2505
R26071 VDD.n4520 VDD.n4519 2.2505
R26072 VDD.n4521 VDD.n2448 2.2505
R26073 VDD.n4523 VDD.n4522 2.2505
R26074 VDD.n4524 VDD.n2447 2.2505
R26075 VDD.n4526 VDD.n4525 2.2505
R26076 VDD.n4527 VDD.n2446 2.2505
R26077 VDD.n4529 VDD.n4528 2.2505
R26078 VDD.n4530 VDD.n2445 2.2505
R26079 VDD.n4532 VDD.n4531 2.2505
R26080 VDD.n4533 VDD.n2444 2.2505
R26081 VDD.n4535 VDD.n4534 2.2505
R26082 VDD.n4536 VDD.n2443 2.2505
R26083 VDD.n4538 VDD.n4537 2.2505
R26084 VDD.n4539 VDD.n2442 2.2505
R26085 VDD.n4541 VDD.n4540 2.2505
R26086 VDD.n4542 VDD.n2441 2.2505
R26087 VDD.n4544 VDD.n4543 2.2505
R26088 VDD.n4545 VDD.n2440 2.2505
R26089 VDD.n4547 VDD.n4546 2.2505
R26090 VDD.n4548 VDD.n2439 2.2505
R26091 VDD.n4550 VDD.n4549 2.2505
R26092 VDD.n4551 VDD.n2438 2.2505
R26093 VDD.n4553 VDD.n4552 2.2505
R26094 VDD.n4554 VDD.n2437 2.2505
R26095 VDD.n4556 VDD.n4555 2.2505
R26096 VDD.n4557 VDD.n2436 2.2505
R26097 VDD.n4559 VDD.n4558 2.2505
R26098 VDD.n4560 VDD.n2435 2.2505
R26099 VDD.n4562 VDD.n4561 2.2505
R26100 VDD.n4563 VDD.n2434 2.2505
R26101 VDD.n4565 VDD.n4564 2.2505
R26102 VDD.n4566 VDD.n2433 2.2505
R26103 VDD.n4568 VDD.n4567 2.2505
R26104 VDD.n4569 VDD.n2432 2.2505
R26105 VDD.n4571 VDD.n4570 2.2505
R26106 VDD.n4572 VDD.n2431 2.2505
R26107 VDD.n4574 VDD.n4573 2.2505
R26108 VDD.n4575 VDD.n2430 2.2505
R26109 VDD.n4577 VDD.n4576 2.2505
R26110 VDD.n4578 VDD.n2429 2.2505
R26111 VDD.n4580 VDD.n4579 2.2505
R26112 VDD.n4581 VDD.n2428 2.2505
R26113 VDD.n4583 VDD.n4582 2.2505
R26114 VDD.n4584 VDD.n2427 2.2505
R26115 VDD.n4586 VDD.n4585 2.2505
R26116 VDD.n4587 VDD.n2426 2.2505
R26117 VDD.n4589 VDD.n4588 2.2505
R26118 VDD.n5200 VDD.n5199 2.2505
R26119 VDD.n5198 VDD.n4598 2.2505
R26120 VDD.n5197 VDD.n5196 2.2505
R26121 VDD.n5195 VDD.n4600 2.2505
R26122 VDD.n5194 VDD.n5193 2.2505
R26123 VDD.n5192 VDD.n4601 2.2505
R26124 VDD.n5191 VDD.n5190 2.2505
R26125 VDD.n5189 VDD.n4602 2.2505
R26126 VDD.n5188 VDD.n5187 2.2505
R26127 VDD.n5186 VDD.n4603 2.2505
R26128 VDD.n5185 VDD.n5184 2.2505
R26129 VDD.n5183 VDD.n4604 2.2505
R26130 VDD.n5182 VDD.n5181 2.2505
R26131 VDD.n5180 VDD.n4605 2.2505
R26132 VDD.n5179 VDD.n5178 2.2505
R26133 VDD.n5177 VDD.n4606 2.2505
R26134 VDD.n5176 VDD.n5175 2.2505
R26135 VDD.n5174 VDD.n4607 2.2505
R26136 VDD.n5173 VDD.n5172 2.2505
R26137 VDD.n5171 VDD.n4608 2.2505
R26138 VDD.n5170 VDD.n5169 2.2505
R26139 VDD.n5168 VDD.n4609 2.2505
R26140 VDD.n5167 VDD.n5166 2.2505
R26141 VDD.n5165 VDD.n4610 2.2505
R26142 VDD.n5164 VDD.n5163 2.2505
R26143 VDD.n5162 VDD.n4611 2.2505
R26144 VDD.n5161 VDD.n5160 2.2505
R26145 VDD.n5159 VDD.n4612 2.2505
R26146 VDD.n5158 VDD.n5157 2.2505
R26147 VDD.n5156 VDD.n4613 2.2505
R26148 VDD.n5155 VDD.n5154 2.2505
R26149 VDD.n5153 VDD.n4614 2.2505
R26150 VDD.n5152 VDD.n5151 2.2505
R26151 VDD.n5150 VDD.n4615 2.2505
R26152 VDD.n5149 VDD.n5148 2.2505
R26153 VDD.n5147 VDD.n4616 2.2505
R26154 VDD.n5146 VDD.n5145 2.2505
R26155 VDD.n5144 VDD.n4617 2.2505
R26156 VDD.n5143 VDD.n5142 2.2505
R26157 VDD.n5141 VDD.n4618 2.2505
R26158 VDD.n5140 VDD.n5139 2.2505
R26159 VDD.n5138 VDD.n4619 2.2505
R26160 VDD.n5137 VDD.n5136 2.2505
R26161 VDD.n5135 VDD.n4620 2.2505
R26162 VDD.n5134 VDD.n5133 2.2505
R26163 VDD.n5132 VDD.n4621 2.2505
R26164 VDD.n5131 VDD.n5130 2.2505
R26165 VDD.n5129 VDD.n4622 2.2505
R26166 VDD.n5128 VDD.n5127 2.2505
R26167 VDD.n5126 VDD.n4623 2.2505
R26168 VDD.n5125 VDD.n5124 2.2505
R26169 VDD.n5123 VDD.n4624 2.2505
R26170 VDD.n5122 VDD.n5121 2.2505
R26171 VDD.n5120 VDD.n4625 2.2505
R26172 VDD.n5119 VDD.n5118 2.2505
R26173 VDD.n5117 VDD.n4626 2.2505
R26174 VDD.n5116 VDD.n5115 2.2505
R26175 VDD.n5114 VDD.n4627 2.2505
R26176 VDD.n5113 VDD.n5112 2.2505
R26177 VDD.n5111 VDD.n4628 2.2505
R26178 VDD.n5110 VDD.n5109 2.2505
R26179 VDD.n5108 VDD.n4629 2.2505
R26180 VDD.n5107 VDD.n5106 2.2505
R26181 VDD.n5105 VDD.n4630 2.2505
R26182 VDD.n5104 VDD.n5103 2.2505
R26183 VDD.n5102 VDD.n4631 2.2505
R26184 VDD.n5101 VDD.n5100 2.2505
R26185 VDD.n5099 VDD.n4632 2.2505
R26186 VDD.n5098 VDD.n5097 2.2505
R26187 VDD.n5096 VDD.n4633 2.2505
R26188 VDD.n5095 VDD.n5094 2.2505
R26189 VDD.n5093 VDD.n4634 2.2505
R26190 VDD.n5092 VDD.n5091 2.2505
R26191 VDD.n5090 VDD.n4635 2.2505
R26192 VDD.n5089 VDD.n5088 2.2505
R26193 VDD.n5087 VDD.n4636 2.2505
R26194 VDD.n5086 VDD.n5085 2.2505
R26195 VDD.n5084 VDD.n4637 2.2505
R26196 VDD.n5083 VDD.n5082 2.2505
R26197 VDD.n5081 VDD.n4638 2.2505
R26198 VDD.n5080 VDD.n5079 2.2505
R26199 VDD.n5078 VDD.n4639 2.2505
R26200 VDD.n5077 VDD.n5076 2.2505
R26201 VDD.n5075 VDD.n4640 2.2505
R26202 VDD.n5074 VDD.n5073 2.2505
R26203 VDD.n5072 VDD.n4641 2.2505
R26204 VDD.n5071 VDD.n5070 2.2505
R26205 VDD.n5069 VDD.n4642 2.2505
R26206 VDD.n5068 VDD.n5067 2.2505
R26207 VDD.n5066 VDD.n4643 2.2505
R26208 VDD.n5065 VDD.n5064 2.2505
R26209 VDD.n5063 VDD.n4644 2.2505
R26210 VDD.n5062 VDD.n5061 2.2505
R26211 VDD.n5060 VDD.n4645 2.2505
R26212 VDD.n5059 VDD.n5058 2.2505
R26213 VDD.n5057 VDD.n4646 2.2505
R26214 VDD.n5056 VDD.n5055 2.2505
R26215 VDD.n5054 VDD.n4647 2.2505
R26216 VDD.n5053 VDD.n5052 2.2505
R26217 VDD.n5051 VDD.n4648 2.2505
R26218 VDD.n5050 VDD.n5049 2.2505
R26219 VDD.n5048 VDD.n4649 2.2505
R26220 VDD.n5047 VDD.n5046 2.2505
R26221 VDD.n5045 VDD.n4650 2.2505
R26222 VDD.n5044 VDD.n5043 2.2505
R26223 VDD.n5042 VDD.n4651 2.2505
R26224 VDD.n5041 VDD.n5040 2.2505
R26225 VDD.n5039 VDD.n4652 2.2505
R26226 VDD.n5038 VDD.n5037 2.2505
R26227 VDD.n5036 VDD.n4653 2.2505
R26228 VDD.n5035 VDD.n5034 2.2505
R26229 VDD.n5033 VDD.n4654 2.2505
R26230 VDD.n5032 VDD.n5031 2.2505
R26231 VDD.n5030 VDD.n4655 2.2505
R26232 VDD.n5029 VDD.n5028 2.2505
R26233 VDD.n5027 VDD.n4656 2.2505
R26234 VDD.n5026 VDD.n5025 2.2505
R26235 VDD.n5024 VDD.n4657 2.2505
R26236 VDD.n5023 VDD.n5022 2.2505
R26237 VDD.n5021 VDD.n4658 2.2505
R26238 VDD.n5020 VDD.n5019 2.2505
R26239 VDD.n5018 VDD.n4659 2.2505
R26240 VDD.n5017 VDD.n5016 2.2505
R26241 VDD.n5015 VDD.n4660 2.2505
R26242 VDD.n5014 VDD.n5013 2.2505
R26243 VDD.n5012 VDD.n4661 2.2505
R26244 VDD.n5011 VDD.n5010 2.2505
R26245 VDD.n5009 VDD.n4662 2.2505
R26246 VDD.n5008 VDD.n5007 2.2505
R26247 VDD.n5006 VDD.n4663 2.2505
R26248 VDD.n5005 VDD.n5004 2.2505
R26249 VDD.n5003 VDD.n4664 2.2505
R26250 VDD.n5002 VDD.n5001 2.2505
R26251 VDD.n5000 VDD.n4665 2.2505
R26252 VDD.n4999 VDD.n4998 2.2505
R26253 VDD.n4997 VDD.n4666 2.2505
R26254 VDD.n4996 VDD.n4995 2.2505
R26255 VDD.n4994 VDD.n4667 2.2505
R26256 VDD.n4993 VDD.n4992 2.2505
R26257 VDD.n4991 VDD.n4668 2.2505
R26258 VDD.n4990 VDD.n4989 2.2505
R26259 VDD.n4988 VDD.n4669 2.2505
R26260 VDD.n4987 VDD.n4986 2.2505
R26261 VDD.n4985 VDD.n4670 2.2505
R26262 VDD.n4984 VDD.n4983 2.2505
R26263 VDD.n4982 VDD.n4671 2.2505
R26264 VDD.n4981 VDD.n4980 2.2505
R26265 VDD.n4979 VDD.n4672 2.2505
R26266 VDD.n4978 VDD.n4977 2.2505
R26267 VDD.n4976 VDD.n4673 2.2505
R26268 VDD.n4975 VDD.n4974 2.2505
R26269 VDD.n4973 VDD.n4674 2.2505
R26270 VDD.n4972 VDD.n4971 2.2505
R26271 VDD.n4970 VDD.n4675 2.2505
R26272 VDD.n4969 VDD.n4968 2.2505
R26273 VDD.n4967 VDD.n4676 2.2505
R26274 VDD.n4966 VDD.n4965 2.2505
R26275 VDD.n4964 VDD.n4677 2.2505
R26276 VDD.n4963 VDD.n4962 2.2505
R26277 VDD.n4961 VDD.n4678 2.2505
R26278 VDD.n4960 VDD.n4959 2.2505
R26279 VDD.n4958 VDD.n4679 2.2505
R26280 VDD.n4957 VDD.n4956 2.2505
R26281 VDD.n4955 VDD.n4680 2.2505
R26282 VDD.n4954 VDD.n4953 2.2505
R26283 VDD.n4952 VDD.n4681 2.2505
R26284 VDD.n4951 VDD.n4950 2.2505
R26285 VDD.n4949 VDD.n4682 2.2505
R26286 VDD.n4948 VDD.n4947 2.2505
R26287 VDD.n4946 VDD.n4683 2.2505
R26288 VDD.n4945 VDD.n4944 2.2505
R26289 VDD.n4943 VDD.n4684 2.2505
R26290 VDD.n4942 VDD.n4941 2.2505
R26291 VDD.n4940 VDD.n4685 2.2505
R26292 VDD.n4939 VDD.n4938 2.2505
R26293 VDD.n4937 VDD.n4686 2.2505
R26294 VDD.n4936 VDD.n4935 2.2505
R26295 VDD.n4934 VDD.n4687 2.2505
R26296 VDD.n4933 VDD.n4932 2.2505
R26297 VDD.n4931 VDD.n4688 2.2505
R26298 VDD.n4930 VDD.n4929 2.2505
R26299 VDD.n4928 VDD.n4689 2.2505
R26300 VDD.n4927 VDD.n4926 2.2505
R26301 VDD.n4925 VDD.n4690 2.2505
R26302 VDD.n4924 VDD.n4923 2.2505
R26303 VDD.n4922 VDD.n4691 2.2505
R26304 VDD.n4921 VDD.n4920 2.2505
R26305 VDD.n4919 VDD.n4692 2.2505
R26306 VDD.n4918 VDD.n4917 2.2505
R26307 VDD.n4916 VDD.n4693 2.2505
R26308 VDD.n4915 VDD.n4914 2.2505
R26309 VDD.n4913 VDD.n4694 2.2505
R26310 VDD.n4912 VDD.n4911 2.2505
R26311 VDD.n4910 VDD.n4695 2.2505
R26312 VDD.n4909 VDD.n4908 2.2505
R26313 VDD.n4907 VDD.n4696 2.2505
R26314 VDD.n4906 VDD.n4905 2.2505
R26315 VDD.n1768 VDD.n1767 2.2505
R26316 VDD.n11039 VDD.n11038 2.2505
R26317 VDD.n11043 VDD.n11042 2.2505
R26318 VDD.n11041 VDD.n673 2.2505
R26319 VDD.n11040 VDD.n676 2.2505
R26320 VDD.n11049 VDD.n668 2.2505
R26321 VDD.n11051 VDD.n11050 2.2505
R26322 VDD.n11052 VDD.n667 2.2505
R26323 VDD.n11054 VDD.n11053 2.2505
R26324 VDD.n11055 VDD.n666 2.2505
R26325 VDD.n11059 VDD.n11058 2.2505
R26326 VDD.n11060 VDD.n665 2.2505
R26327 VDD.n11062 VDD.n11061 2.2505
R26328 VDD.n11064 VDD.n664 2.2505
R26329 VDD.n11066 VDD.n11065 2.2505
R26330 VDD.n11067 VDD.n663 2.2505
R26331 VDD.n11069 VDD.n11068 2.2505
R26332 VDD.n11070 VDD.n662 2.2505
R26333 VDD.n11072 VDD.n11071 2.2505
R26334 VDD.n11074 VDD.n11073 2.2505
R26335 VDD.n11075 VDD.n660 2.2505
R26336 VDD.n11079 VDD.n11078 2.2505
R26337 VDD.n11080 VDD.n659 2.2505
R26338 VDD.n11082 VDD.n11081 2.2505
R26339 VDD.n11083 VDD.n658 2.2505
R26340 VDD.n11085 VDD.n11084 2.2505
R26341 VDD.n11087 VDD.n11086 2.2505
R26342 VDD.n11088 VDD.n656 2.2505
R26343 VDD.n11092 VDD.n11091 2.2505
R26344 VDD.n11093 VDD.n655 2.2505
R26345 VDD.n11095 VDD.n11094 2.2505
R26346 VDD.n11096 VDD.n654 2.2505
R26347 VDD.n11099 VDD.n11098 2.2505
R26348 VDD.n11100 VDD.n653 2.2505
R26349 VDD.n11102 VDD.n11101 2.2505
R26350 VDD.n11103 VDD.n652 2.2505
R26351 VDD.n11105 VDD.n11104 2.2505
R26352 VDD.n11107 VDD.n11106 2.2505
R26353 VDD.n11108 VDD.n650 2.2505
R26354 VDD.n11110 VDD.n11109 2.2505
R26355 VDD.n11112 VDD.n11111 2.2505
R26356 VDD.n11113 VDD.n647 2.2505
R26357 VDD.n11115 VDD.n11114 2.2505
R26358 VDD.n11116 VDD.n646 2.2505
R26359 VDD.n11118 VDD.n11117 2.2505
R26360 VDD.n11120 VDD.n645 2.2505
R26361 VDD.n11122 VDD.n11121 2.2505
R26362 VDD.n11124 VDD.n11123 2.2505
R26363 VDD.n11126 VDD.n11125 2.2505
R26364 VDD.n633 VDD.n632 2.2505
R26365 VDD.n11132 VDD.n11131 2.2505
R26366 VDD.n11133 VDD.n631 2.2505
R26367 VDD.n3629 VDD.n3628 2.2505
R26368 VDD.n3627 VDD.n2746 2.2505
R26369 VDD.n3626 VDD.n3625 2.2505
R26370 VDD.n3624 VDD.n2747 2.2505
R26371 VDD.n3623 VDD.n3622 2.2505
R26372 VDD.n3621 VDD.n2748 2.2505
R26373 VDD.n3620 VDD.n3619 2.2505
R26374 VDD.n3618 VDD.n2749 2.2505
R26375 VDD.n3617 VDD.n3616 2.2505
R26376 VDD.n3615 VDD.n2750 2.2505
R26377 VDD.n3614 VDD.n3613 2.2505
R26378 VDD.n3612 VDD.n2751 2.2505
R26379 VDD.n3611 VDD.n3610 2.2505
R26380 VDD.n3609 VDD.n2752 2.2505
R26381 VDD.n3608 VDD.n3607 2.2505
R26382 VDD.n3606 VDD.n2753 2.2505
R26383 VDD.n3605 VDD.n3604 2.2505
R26384 VDD.n3603 VDD.n2754 2.2505
R26385 VDD.n3602 VDD.n3601 2.2505
R26386 VDD.n3600 VDD.n2755 2.2505
R26387 VDD.n3599 VDD.n3598 2.2505
R26388 VDD.n3597 VDD.n2756 2.2505
R26389 VDD.n3596 VDD.n3595 2.2505
R26390 VDD.n3594 VDD.n2757 2.2505
R26391 VDD.n3593 VDD.n3592 2.2505
R26392 VDD.n3591 VDD.n2758 2.2505
R26393 VDD.n3590 VDD.n3589 2.2505
R26394 VDD.n3588 VDD.n2759 2.2505
R26395 VDD.n3587 VDD.n3586 2.2505
R26396 VDD.n3585 VDD.n2760 2.2505
R26397 VDD.n3584 VDD.n3583 2.2505
R26398 VDD.n3582 VDD.n2761 2.2505
R26399 VDD.n3581 VDD.n3580 2.2505
R26400 VDD.n3579 VDD.n2762 2.2505
R26401 VDD.n3578 VDD.n3577 2.2505
R26402 VDD.n3576 VDD.n2763 2.2505
R26403 VDD.n3575 VDD.n3574 2.2505
R26404 VDD.n3573 VDD.n2764 2.2505
R26405 VDD.n3572 VDD.n3571 2.2505
R26406 VDD.n3570 VDD.n2765 2.2505
R26407 VDD.n3569 VDD.n3568 2.2505
R26408 VDD.n3567 VDD.n2766 2.2505
R26409 VDD.n3566 VDD.n3565 2.2505
R26410 VDD.n3564 VDD.n2767 2.2505
R26411 VDD.n3563 VDD.n3562 2.2505
R26412 VDD.n3561 VDD.n2768 2.2505
R26413 VDD.n3560 VDD.n3559 2.2505
R26414 VDD.n3558 VDD.n2769 2.2505
R26415 VDD.n3557 VDD.n3556 2.2505
R26416 VDD.n3555 VDD.n2770 2.2505
R26417 VDD.n3554 VDD.n3553 2.2505
R26418 VDD.n3552 VDD.n2771 2.2505
R26419 VDD.n3551 VDD.n3550 2.2505
R26420 VDD.n3549 VDD.n2772 2.2505
R26421 VDD.n3548 VDD.n3547 2.2505
R26422 VDD.n3546 VDD.n2773 2.2505
R26423 VDD.n3545 VDD.n3544 2.2505
R26424 VDD.n3543 VDD.n2774 2.2505
R26425 VDD.n3542 VDD.n3541 2.2505
R26426 VDD.n3540 VDD.n2775 2.2505
R26427 VDD.n3539 VDD.n3538 2.2505
R26428 VDD.n3537 VDD.n2776 2.2505
R26429 VDD.n3536 VDD.n3535 2.2505
R26430 VDD.n3534 VDD.n2777 2.2505
R26431 VDD.n3533 VDD.n3532 2.2505
R26432 VDD.n3531 VDD.n2778 2.2505
R26433 VDD.n3530 VDD.n3529 2.2505
R26434 VDD.n3528 VDD.n2779 2.2505
R26435 VDD.n3527 VDD.n3526 2.2505
R26436 VDD.n3525 VDD.n2780 2.2505
R26437 VDD.n3524 VDD.n3523 2.2505
R26438 VDD.n3522 VDD.n2781 2.2505
R26439 VDD.n3521 VDD.n3520 2.2505
R26440 VDD.n3519 VDD.n2782 2.2505
R26441 VDD.n3518 VDD.n3517 2.2505
R26442 VDD.n3516 VDD.n2783 2.2505
R26443 VDD.n3515 VDD.n3514 2.2505
R26444 VDD.n3513 VDD.n2784 2.2505
R26445 VDD.n3512 VDD.n3511 2.2505
R26446 VDD.n3510 VDD.n2785 2.2505
R26447 VDD.n3509 VDD.n3508 2.2505
R26448 VDD.n3507 VDD.n2786 2.2505
R26449 VDD.n3506 VDD.n3505 2.2505
R26450 VDD.n3504 VDD.n2787 2.2505
R26451 VDD.n3503 VDD.n3502 2.2505
R26452 VDD.n3501 VDD.n2788 2.2505
R26453 VDD.n3500 VDD.n3499 2.2505
R26454 VDD.n3498 VDD.n2789 2.2505
R26455 VDD.n3497 VDD.n3496 2.2505
R26456 VDD.n3495 VDD.n2790 2.2505
R26457 VDD.n3494 VDD.n3493 2.2505
R26458 VDD.n3492 VDD.n2791 2.2505
R26459 VDD.n3491 VDD.n3490 2.2505
R26460 VDD.n3489 VDD.n2792 2.2505
R26461 VDD.n3488 VDD.n3487 2.2505
R26462 VDD.n3486 VDD.n2793 2.2505
R26463 VDD.n3485 VDD.n3484 2.2505
R26464 VDD.n3483 VDD.n2794 2.2505
R26465 VDD.n3482 VDD.n3481 2.2505
R26466 VDD.n3480 VDD.n2795 2.2505
R26467 VDD.n3479 VDD.n3478 2.2505
R26468 VDD.n3477 VDD.n2796 2.2505
R26469 VDD.n3476 VDD.n3475 2.2505
R26470 VDD.n3474 VDD.n2797 2.2505
R26471 VDD.n3473 VDD.n3472 2.2505
R26472 VDD.n3471 VDD.n2798 2.2505
R26473 VDD.n3470 VDD.n3469 2.2505
R26474 VDD.n3468 VDD.n2799 2.2505
R26475 VDD.n3467 VDD.n3466 2.2505
R26476 VDD.n3465 VDD.n2800 2.2505
R26477 VDD.n3464 VDD.n3463 2.2505
R26478 VDD.n3462 VDD.n2801 2.2505
R26479 VDD.n3461 VDD.n3460 2.2505
R26480 VDD.n3459 VDD.n2802 2.2505
R26481 VDD.n3458 VDD.n3457 2.2505
R26482 VDD.n3456 VDD.n2803 2.2505
R26483 VDD.n3455 VDD.n3454 2.2505
R26484 VDD.n3453 VDD.n2804 2.2505
R26485 VDD.n3452 VDD.n3451 2.2505
R26486 VDD.n3450 VDD.n2805 2.2505
R26487 VDD.n3449 VDD.n3448 2.2505
R26488 VDD.n3447 VDD.n2806 2.2505
R26489 VDD.n3446 VDD.n3445 2.2505
R26490 VDD.n3444 VDD.n2807 2.2505
R26491 VDD.n3443 VDD.n3442 2.2505
R26492 VDD.n3441 VDD.n2808 2.2505
R26493 VDD.n3440 VDD.n3439 2.2505
R26494 VDD.n3438 VDD.n2809 2.2505
R26495 VDD.n3437 VDD.n3436 2.2505
R26496 VDD.n3435 VDD.n2810 2.2505
R26497 VDD.n3434 VDD.n3433 2.2505
R26498 VDD.n3432 VDD.n2811 2.2505
R26499 VDD.n3431 VDD.n3430 2.2505
R26500 VDD.n3429 VDD.n2812 2.2505
R26501 VDD.n3428 VDD.n3427 2.2505
R26502 VDD.n3426 VDD.n2813 2.2505
R26503 VDD.n3425 VDD.n3424 2.2505
R26504 VDD.n3423 VDD.n2814 2.2505
R26505 VDD.n3422 VDD.n3421 2.2505
R26506 VDD.n3420 VDD.n2815 2.2505
R26507 VDD.n3419 VDD.n3418 2.2505
R26508 VDD.n3417 VDD.n2816 2.2505
R26509 VDD.n3416 VDD.n3415 2.2505
R26510 VDD.n3414 VDD.n2817 2.2505
R26511 VDD.n3413 VDD.n3412 2.2505
R26512 VDD.n3411 VDD.n2818 2.2505
R26513 VDD.n3410 VDD.n3409 2.2505
R26514 VDD.n3408 VDD.n2819 2.2505
R26515 VDD.n3407 VDD.n3406 2.2505
R26516 VDD.n3405 VDD.n2820 2.2505
R26517 VDD.n3404 VDD.n3403 2.2505
R26518 VDD.n3402 VDD.n2821 2.2505
R26519 VDD.n3401 VDD.n3400 2.2505
R26520 VDD.n3399 VDD.n2822 2.2505
R26521 VDD.n3398 VDD.n3397 2.2505
R26522 VDD.n3396 VDD.n2823 2.2505
R26523 VDD.n3395 VDD.n3394 2.2505
R26524 VDD.n3393 VDD.n2824 2.2505
R26525 VDD.n3392 VDD.n3391 2.2505
R26526 VDD.n3390 VDD.n2825 2.2505
R26527 VDD.n3389 VDD.n3388 2.2505
R26528 VDD.n3387 VDD.n2826 2.2505
R26529 VDD.n3386 VDD.n3385 2.2505
R26530 VDD.n3384 VDD.n2827 2.2505
R26531 VDD.n3383 VDD.n3382 2.2505
R26532 VDD.n3381 VDD.n2828 2.2505
R26533 VDD.n3380 VDD.n3379 2.2505
R26534 VDD.n3378 VDD.n2829 2.2505
R26535 VDD.n3377 VDD.n3376 2.2505
R26536 VDD.n3375 VDD.n2830 2.2505
R26537 VDD.n3374 VDD.n3373 2.2505
R26538 VDD.n3372 VDD.n2831 2.2505
R26539 VDD.n3371 VDD.n3370 2.2505
R26540 VDD.n3369 VDD.n2832 2.2505
R26541 VDD.n3368 VDD.n3367 2.2505
R26542 VDD.n3366 VDD.n2833 2.2505
R26543 VDD.n3365 VDD.n3364 2.2505
R26544 VDD.n3363 VDD.n2834 2.2505
R26545 VDD.n3362 VDD.n3361 2.2505
R26546 VDD.n3360 VDD.n2835 2.2505
R26547 VDD.n3359 VDD.n3358 2.2505
R26548 VDD.n3357 VDD.n2836 2.2505
R26549 VDD.n3356 VDD.n3355 2.2505
R26550 VDD.n3354 VDD.n2837 2.2505
R26551 VDD.n3353 VDD.n3352 2.2505
R26552 VDD.n3351 VDD.n2838 2.2505
R26553 VDD.n3350 VDD.n3349 2.2505
R26554 VDD.n3348 VDD.n2839 2.2505
R26555 VDD.n3347 VDD.n3346 2.2505
R26556 VDD.n3345 VDD.n2840 2.2505
R26557 VDD.n3344 VDD.n3343 2.2505
R26558 VDD.n3342 VDD.n2841 2.2505
R26559 VDD.n3341 VDD.n3340 2.2505
R26560 VDD.n3339 VDD.n2842 2.2505
R26561 VDD.n3338 VDD.n3337 2.2505
R26562 VDD.n3336 VDD.n2843 2.2505
R26563 VDD.n3335 VDD.n3334 2.2505
R26564 VDD.n3333 VDD.n2844 2.2505
R26565 VDD.n3332 VDD.n3331 2.2505
R26566 VDD.n3330 VDD.n2845 2.2505
R26567 VDD.n3329 VDD.n3328 2.2505
R26568 VDD.n3327 VDD.n2846 2.2505
R26569 VDD.n3326 VDD.n3325 2.2505
R26570 VDD.n3324 VDD.n2847 2.2505
R26571 VDD.n3323 VDD.n3322 2.2505
R26572 VDD.n3321 VDD.n2848 2.2505
R26573 VDD.n3320 VDD.n3319 2.2505
R26574 VDD.n3318 VDD.n2849 2.2505
R26575 VDD.n3317 VDD.n3316 2.2505
R26576 VDD.n3315 VDD.n2850 2.2505
R26577 VDD.n3314 VDD.n3313 2.2505
R26578 VDD.n3312 VDD.n2851 2.2505
R26579 VDD.n3311 VDD.n3310 2.2505
R26580 VDD.n3309 VDD.n2852 2.2505
R26581 VDD.n3308 VDD.n3307 2.2505
R26582 VDD.n3306 VDD.n2853 2.2505
R26583 VDD.n3305 VDD.n3304 2.2505
R26584 VDD.n3303 VDD.n2854 2.2505
R26585 VDD.n3302 VDD.n3301 2.2505
R26586 VDD.n3300 VDD.n2855 2.2505
R26587 VDD.n3299 VDD.n3298 2.2505
R26588 VDD.n3297 VDD.n2856 2.2505
R26589 VDD.n3296 VDD.n3295 2.2505
R26590 VDD.n3294 VDD.n2857 2.2505
R26591 VDD.n3293 VDD.n3292 2.2505
R26592 VDD.n3291 VDD.n2858 2.2505
R26593 VDD.n3290 VDD.n3289 2.2505
R26594 VDD.n3288 VDD.n2859 2.2505
R26595 VDD.n3287 VDD.n3286 2.2505
R26596 VDD.n3285 VDD.n2860 2.2505
R26597 VDD.n3284 VDD.n3283 2.2505
R26598 VDD.n3282 VDD.n2861 2.2505
R26599 VDD.n3281 VDD.n3280 2.2505
R26600 VDD.n3279 VDD.n2862 2.2505
R26601 VDD.n3278 VDD.n3277 2.2505
R26602 VDD.n3276 VDD.n2863 2.2505
R26603 VDD.n3275 VDD.n3274 2.2505
R26604 VDD.n3273 VDD.n2864 2.2505
R26605 VDD.n3272 VDD.n3271 2.2505
R26606 VDD.n3270 VDD.n2865 2.2505
R26607 VDD.n3269 VDD.n3268 2.2505
R26608 VDD.n3267 VDD.n2866 2.2505
R26609 VDD.n3266 VDD.n3265 2.2505
R26610 VDD.n3264 VDD.n2867 2.2505
R26611 VDD.n3263 VDD.n3262 2.2505
R26612 VDD.n3261 VDD.n2868 2.2505
R26613 VDD.n3260 VDD.n3259 2.2505
R26614 VDD.n3258 VDD.n2869 2.2505
R26615 VDD.n3257 VDD.n3256 2.2505
R26616 VDD.n3255 VDD.n2870 2.2505
R26617 VDD.n3254 VDD.n3253 2.2505
R26618 VDD.n3252 VDD.n2871 2.2505
R26619 VDD.n3251 VDD.n3250 2.2505
R26620 VDD.n3249 VDD.n2872 2.2505
R26621 VDD.n3248 VDD.n3247 2.2505
R26622 VDD.n3246 VDD.n2873 2.2505
R26623 VDD.n3245 VDD.n3244 2.2505
R26624 VDD.n3243 VDD.n2874 2.2505
R26625 VDD.n3242 VDD.n3241 2.2505
R26626 VDD.n3240 VDD.n2875 2.2505
R26627 VDD.n3239 VDD.n3238 2.2505
R26628 VDD.n3237 VDD.n2876 2.2505
R26629 VDD.n3236 VDD.n3235 2.2505
R26630 VDD.n3234 VDD.n2877 2.2505
R26631 VDD.n3233 VDD.n3232 2.2505
R26632 VDD.n3231 VDD.n2878 2.2505
R26633 VDD.n3230 VDD.n3229 2.2505
R26634 VDD.n3228 VDD.n2879 2.2505
R26635 VDD.n3227 VDD.n3226 2.2505
R26636 VDD.n3225 VDD.n2880 2.2505
R26637 VDD.n3224 VDD.n3223 2.2505
R26638 VDD.n3222 VDD.n2881 2.2505
R26639 VDD.n3221 VDD.n3220 2.2505
R26640 VDD.n3219 VDD.n2882 2.2505
R26641 VDD.n3218 VDD.n3217 2.2505
R26642 VDD.n3216 VDD.n2883 2.2505
R26643 VDD.n3215 VDD.n3214 2.2505
R26644 VDD.n3213 VDD.n2884 2.2505
R26645 VDD.n3212 VDD.n3211 2.2505
R26646 VDD.n3210 VDD.n2885 2.2505
R26647 VDD.n3209 VDD.n3208 2.2505
R26648 VDD.n3207 VDD.n2886 2.2505
R26649 VDD.n3206 VDD.n3205 2.2505
R26650 VDD.n3204 VDD.n2887 2.2505
R26651 VDD.n3203 VDD.n3202 2.2505
R26652 VDD.n3201 VDD.n2888 2.2505
R26653 VDD.n3200 VDD.n3199 2.2505
R26654 VDD.n3198 VDD.n2889 2.2505
R26655 VDD.n3197 VDD.n3196 2.2505
R26656 VDD.n3195 VDD.n2890 2.2505
R26657 VDD.n3194 VDD.n3193 2.2505
R26658 VDD.n3192 VDD.n2891 2.2505
R26659 VDD.n3191 VDD.n3190 2.2505
R26660 VDD.n3189 VDD.n2892 2.2505
R26661 VDD.n3188 VDD.n3187 2.2505
R26662 VDD.n3186 VDD.n2893 2.2505
R26663 VDD.n3185 VDD.n3184 2.2505
R26664 VDD.n3183 VDD.n2894 2.2505
R26665 VDD.n3182 VDD.n3181 2.2505
R26666 VDD.n3180 VDD.n2895 2.2505
R26667 VDD.n3179 VDD.n3178 2.2505
R26668 VDD.n3177 VDD.n2896 2.2505
R26669 VDD.n3176 VDD.n3175 2.2505
R26670 VDD.n3174 VDD.n2897 2.2505
R26671 VDD.n3173 VDD.n3172 2.2505
R26672 VDD.n3171 VDD.n2898 2.2505
R26673 VDD.n3170 VDD.n3169 2.2505
R26674 VDD.n3168 VDD.n2899 2.2505
R26675 VDD.n3167 VDD.n3166 2.2505
R26676 VDD.n3165 VDD.n2900 2.2505
R26677 VDD.n3164 VDD.n3163 2.2505
R26678 VDD.n3162 VDD.n2901 2.2505
R26679 VDD.n3161 VDD.n3160 2.2505
R26680 VDD.n3159 VDD.n2902 2.2505
R26681 VDD.n3158 VDD.n3157 2.2505
R26682 VDD.n3156 VDD.n2903 2.2505
R26683 VDD.n3155 VDD.n3154 2.2505
R26684 VDD.n3153 VDD.n2904 2.2505
R26685 VDD.n3152 VDD.n3151 2.2505
R26686 VDD.n3150 VDD.n2905 2.2505
R26687 VDD.n3149 VDD.n3148 2.2505
R26688 VDD.n3147 VDD.n2906 2.2505
R26689 VDD.n3146 VDD.n3145 2.2505
R26690 VDD.n3144 VDD.n2907 2.2505
R26691 VDD.n3143 VDD.n3142 2.2505
R26692 VDD.n3141 VDD.n2908 2.2505
R26693 VDD.n3140 VDD.n3139 2.2505
R26694 VDD.n3138 VDD.n2909 2.2505
R26695 VDD.n3137 VDD.n3136 2.2505
R26696 VDD.n3135 VDD.n2910 2.2505
R26697 VDD.n3134 VDD.n3133 2.2505
R26698 VDD.n3132 VDD.n2911 2.2505
R26699 VDD.n3131 VDD.n3130 2.2505
R26700 VDD.n3129 VDD.n2912 2.2505
R26701 VDD.n3128 VDD.n3127 2.2505
R26702 VDD.n3126 VDD.n2913 2.2505
R26703 VDD.n3125 VDD.n3124 2.2505
R26704 VDD.n3123 VDD.n2914 2.2505
R26705 VDD.n3122 VDD.n3121 2.2505
R26706 VDD.n3120 VDD.n2915 2.2505
R26707 VDD.n3119 VDD.n3118 2.2505
R26708 VDD.n3117 VDD.n2916 2.2505
R26709 VDD.n3116 VDD.n3115 2.2505
R26710 VDD.n3114 VDD.n2917 2.2505
R26711 VDD.n3113 VDD.n3112 2.2505
R26712 VDD.n3111 VDD.n2918 2.2505
R26713 VDD.n3110 VDD.n3109 2.2505
R26714 VDD.n3108 VDD.n2919 2.2505
R26715 VDD.n3107 VDD.n3106 2.2505
R26716 VDD.n3105 VDD.n2920 2.2505
R26717 VDD.n3104 VDD.n3103 2.2505
R26718 VDD.n3102 VDD.n2921 2.2505
R26719 VDD.n3101 VDD.n3100 2.2505
R26720 VDD.n3099 VDD.n2922 2.2505
R26721 VDD.n3098 VDD.n3097 2.2505
R26722 VDD.n3096 VDD.n2923 2.2505
R26723 VDD.n3095 VDD.n3094 2.2505
R26724 VDD.n3093 VDD.n2924 2.2505
R26725 VDD.n3092 VDD.n3091 2.2505
R26726 VDD.n3090 VDD.n2925 2.2505
R26727 VDD.n3089 VDD.n3088 2.2505
R26728 VDD.n3087 VDD.n2926 2.2505
R26729 VDD.n3086 VDD.n3085 2.2505
R26730 VDD.n3084 VDD.n2927 2.2505
R26731 VDD.n3083 VDD.n3082 2.2505
R26732 VDD.n3081 VDD.n2928 2.2505
R26733 VDD.n3080 VDD.n3079 2.2505
R26734 VDD.n3078 VDD.n2929 2.2505
R26735 VDD.n3077 VDD.n3076 2.2505
R26736 VDD.n3075 VDD.n2930 2.2505
R26737 VDD.n3074 VDD.n3073 2.2505
R26738 VDD.n3072 VDD.n2931 2.2505
R26739 VDD.n3071 VDD.n3070 2.2505
R26740 VDD.n3069 VDD.n2932 2.2505
R26741 VDD.n3068 VDD.n3067 2.2505
R26742 VDD.n3066 VDD.n2933 2.2505
R26743 VDD.n3065 VDD.n3064 2.2505
R26744 VDD.n3063 VDD.n2934 2.2505
R26745 VDD.n3062 VDD.n3061 2.2505
R26746 VDD.n3060 VDD.n2935 2.2505
R26747 VDD.n3059 VDD.n3058 2.2505
R26748 VDD.n3057 VDD.n2936 2.2505
R26749 VDD.n3056 VDD.n3055 2.2505
R26750 VDD.n3054 VDD.n2937 2.2505
R26751 VDD.n3053 VDD.n3052 2.2505
R26752 VDD.n3051 VDD.n2938 2.2505
R26753 VDD.n3050 VDD.n3049 2.2505
R26754 VDD.n3048 VDD.n2939 2.2505
R26755 VDD.n3047 VDD.n3046 2.2505
R26756 VDD.n3045 VDD.n2940 2.2505
R26757 VDD.n3044 VDD.n3043 2.2505
R26758 VDD.n3042 VDD.n2941 2.2505
R26759 VDD.n3041 VDD.n3040 2.2505
R26760 VDD.n3039 VDD.n2942 2.2505
R26761 VDD.n3038 VDD.n3037 2.2505
R26762 VDD.n3036 VDD.n2943 2.2505
R26763 VDD.n3035 VDD.n3034 2.2505
R26764 VDD.n3033 VDD.n2944 2.2505
R26765 VDD.n3032 VDD.n3031 2.2505
R26766 VDD.n3030 VDD.n2945 2.2505
R26767 VDD.n3029 VDD.n3028 2.2505
R26768 VDD.n3027 VDD.n2946 2.2505
R26769 VDD.n3026 VDD.n3025 2.2505
R26770 VDD.n3024 VDD.n2947 2.2505
R26771 VDD.n3023 VDD.n3022 2.2505
R26772 VDD.n3021 VDD.n2948 2.2505
R26773 VDD.n3020 VDD.n3019 2.2505
R26774 VDD.n3018 VDD.n2949 2.2505
R26775 VDD.n3017 VDD.n3016 2.2505
R26776 VDD.n3015 VDD.n2950 2.2505
R26777 VDD.n3014 VDD.n3013 2.2505
R26778 VDD.n3012 VDD.n2951 2.2505
R26779 VDD.n3011 VDD.n3010 2.2505
R26780 VDD.n3009 VDD.n2952 2.2505
R26781 VDD.n3008 VDD.n3007 2.2505
R26782 VDD.n3006 VDD.n2953 2.2505
R26783 VDD.n3005 VDD.n3004 2.2505
R26784 VDD.n3003 VDD.n2954 2.2505
R26785 VDD.n3002 VDD.n3001 2.2505
R26786 VDD.n3000 VDD.n2955 2.2505
R26787 VDD.n2999 VDD.n2998 2.2505
R26788 VDD.n2997 VDD.n2956 2.2505
R26789 VDD.n2996 VDD.n2995 2.2505
R26790 VDD.n2994 VDD.n2957 2.2505
R26791 VDD.n2993 VDD.n2992 2.2505
R26792 VDD.n2991 VDD.n2958 2.2505
R26793 VDD.n2990 VDD.n2989 2.2505
R26794 VDD.n2988 VDD.n2959 2.2505
R26795 VDD.n2987 VDD.n2986 2.2505
R26796 VDD.n2985 VDD.n2960 2.2505
R26797 VDD.n2984 VDD.n2983 2.2505
R26798 VDD.n2982 VDD.n2961 2.2505
R26799 VDD.n2981 VDD.n2980 2.2505
R26800 VDD.n2979 VDD.n2962 2.2505
R26801 VDD.n2978 VDD.n2977 2.2505
R26802 VDD.n2976 VDD.n2963 2.2505
R26803 VDD.n2975 VDD.n2974 2.2505
R26804 VDD.n2973 VDD.n2964 2.2505
R26805 VDD.n2972 VDD.n2971 2.2505
R26806 VDD.n2970 VDD.n2965 2.2505
R26807 VDD.n2969 VDD.n2968 2.2505
R26808 VDD.n11135 VDD.n11134 2.2505
R26809 VDD.n11136 VDD.n630 2.2505
R26810 VDD.n11138 VDD.n11137 2.2505
R26811 VDD.n11139 VDD.n629 2.2505
R26812 VDD.n11141 VDD.n11140 2.2505
R26813 VDD.n11142 VDD.n628 2.2505
R26814 VDD.n11144 VDD.n11143 2.2505
R26815 VDD.n11145 VDD.n627 2.2505
R26816 VDD.n11147 VDD.n11146 2.2505
R26817 VDD.n11148 VDD.n626 2.2505
R26818 VDD.n11150 VDD.n11149 2.2505
R26819 VDD.n11151 VDD.n625 2.2505
R26820 VDD.n11153 VDD.n11152 2.2505
R26821 VDD.n11154 VDD.n624 2.2505
R26822 VDD.n11156 VDD.n11155 2.2505
R26823 VDD.n11157 VDD.n623 2.2505
R26824 VDD.n11159 VDD.n11158 2.2505
R26825 VDD.n11160 VDD.n622 2.2505
R26826 VDD.n11162 VDD.n11161 2.2505
R26827 VDD.n11163 VDD.n621 2.2505
R26828 VDD.n11165 VDD.n11164 2.2505
R26829 VDD.n11166 VDD.n620 2.2505
R26830 VDD.n11168 VDD.n11167 2.2505
R26831 VDD.n11169 VDD.n619 2.2505
R26832 VDD.n11171 VDD.n11170 2.2505
R26833 VDD.n11172 VDD.n618 2.2505
R26834 VDD.n11174 VDD.n11173 2.2505
R26835 VDD.n11175 VDD.n617 2.2505
R26836 VDD.n11177 VDD.n11176 2.2505
R26837 VDD.n11178 VDD.n616 2.2505
R26838 VDD.n11180 VDD.n11179 2.2505
R26839 VDD.n11181 VDD.n615 2.2505
R26840 VDD.n11183 VDD.n11182 2.2505
R26841 VDD.n11184 VDD.n614 2.2505
R26842 VDD.n11186 VDD.n11185 2.2505
R26843 VDD.n11187 VDD.n613 2.2505
R26844 VDD.n11189 VDD.n11188 2.2505
R26845 VDD.n11190 VDD.n612 2.2505
R26846 VDD.n11192 VDD.n11191 2.2505
R26847 VDD.n11193 VDD.n611 2.2505
R26848 VDD.n11195 VDD.n11194 2.2505
R26849 VDD.n11196 VDD.n610 2.2505
R26850 VDD.n11198 VDD.n11197 2.2505
R26851 VDD.n11199 VDD.n609 2.2505
R26852 VDD.n11201 VDD.n11200 2.2505
R26853 VDD.n11202 VDD.n608 2.2505
R26854 VDD.n11204 VDD.n11203 2.2505
R26855 VDD.n11205 VDD.n607 2.2505
R26856 VDD.n11207 VDD.n11206 2.2505
R26857 VDD.n11208 VDD.n606 2.2505
R26858 VDD.n11210 VDD.n11209 2.2505
R26859 VDD.n11211 VDD.n605 2.2505
R26860 VDD.n11213 VDD.n11212 2.2505
R26861 VDD.n11214 VDD.n604 2.2505
R26862 VDD.n11216 VDD.n11215 2.2505
R26863 VDD.n11217 VDD.n603 2.2505
R26864 VDD.n11219 VDD.n11218 2.2505
R26865 VDD.n11220 VDD.n602 2.2505
R26866 VDD.n11222 VDD.n11221 2.2505
R26867 VDD.n11223 VDD.n601 2.2505
R26868 VDD.n11225 VDD.n11224 2.2505
R26869 VDD.n11226 VDD.n600 2.2505
R26870 VDD.n11228 VDD.n11227 2.2505
R26871 VDD.n11229 VDD.n599 2.2505
R26872 VDD.n11231 VDD.n11230 2.2505
R26873 VDD.n11232 VDD.n598 2.2505
R26874 VDD.n11234 VDD.n11233 2.2505
R26875 VDD.n11235 VDD.n597 2.2505
R26876 VDD.n11237 VDD.n11236 2.2505
R26877 VDD.n11238 VDD.n596 2.2505
R26878 VDD.n11240 VDD.n11239 2.2505
R26879 VDD.n11241 VDD.n595 2.2505
R26880 VDD.n11243 VDD.n11242 2.2505
R26881 VDD.n11244 VDD.n594 2.2505
R26882 VDD.n11246 VDD.n11245 2.2505
R26883 VDD.n11247 VDD.n593 2.2505
R26884 VDD.n11249 VDD.n11248 2.2505
R26885 VDD.n11250 VDD.n592 2.2505
R26886 VDD.n11252 VDD.n11251 2.2505
R26887 VDD.n11253 VDD.n591 2.2505
R26888 VDD.n11255 VDD.n11254 2.2505
R26889 VDD.n11256 VDD.n590 2.2505
R26890 VDD.n11258 VDD.n11257 2.2505
R26891 VDD.n11259 VDD.n589 2.2505
R26892 VDD.n11261 VDD.n11260 2.2505
R26893 VDD.n11262 VDD.n588 2.2505
R26894 VDD.n11264 VDD.n11263 2.2505
R26895 VDD.n11265 VDD.n587 2.2505
R26896 VDD.n11267 VDD.n11266 2.2505
R26897 VDD.n11268 VDD.n586 2.2505
R26898 VDD.n11270 VDD.n11269 2.2505
R26899 VDD.n11271 VDD.n585 2.2505
R26900 VDD.n11273 VDD.n11272 2.2505
R26901 VDD.n11274 VDD.n584 2.2505
R26902 VDD.n11276 VDD.n11275 2.2505
R26903 VDD.n11277 VDD.n583 2.2505
R26904 VDD.n11279 VDD.n11278 2.2505
R26905 VDD.n11280 VDD.n582 2.2505
R26906 VDD.n11282 VDD.n11281 2.2505
R26907 VDD.n11283 VDD.n581 2.2505
R26908 VDD.n11285 VDD.n11284 2.2505
R26909 VDD.n11286 VDD.n580 2.2505
R26910 VDD.n11288 VDD.n11287 2.2505
R26911 VDD.n11289 VDD.n579 2.2505
R26912 VDD.n11291 VDD.n11290 2.2505
R26913 VDD.n11292 VDD.n578 2.2505
R26914 VDD.n11294 VDD.n11293 2.2505
R26915 VDD.n11295 VDD.n577 2.2505
R26916 VDD.n11297 VDD.n11296 2.2505
R26917 VDD.n11298 VDD.n576 2.2505
R26918 VDD.n11300 VDD.n11299 2.2505
R26919 VDD.n11301 VDD.n575 2.2505
R26920 VDD.n11303 VDD.n11302 2.2505
R26921 VDD.n11304 VDD.n574 2.2505
R26922 VDD.n11306 VDD.n11305 2.2505
R26923 VDD.n11307 VDD.n573 2.2505
R26924 VDD.n11309 VDD.n11308 2.2505
R26925 VDD.n11310 VDD.n572 2.2505
R26926 VDD.n11312 VDD.n11311 2.2505
R26927 VDD.n11313 VDD.n571 2.2505
R26928 VDD.n11315 VDD.n11314 2.2505
R26929 VDD.n11316 VDD.n570 2.2505
R26930 VDD.n11318 VDD.n11317 2.2505
R26931 VDD.n11319 VDD.n569 2.2505
R26932 VDD.n11321 VDD.n11320 2.2505
R26933 VDD.n11322 VDD.n568 2.2505
R26934 VDD.n11324 VDD.n11323 2.2505
R26935 VDD.n11325 VDD.n567 2.2505
R26936 VDD.n11327 VDD.n11326 2.2505
R26937 VDD.n11328 VDD.n566 2.2505
R26938 VDD.n11330 VDD.n11329 2.2505
R26939 VDD.n11331 VDD.n565 2.2505
R26940 VDD.n11333 VDD.n11332 2.2505
R26941 VDD.n11334 VDD.n564 2.2505
R26942 VDD.n11336 VDD.n11335 2.2505
R26943 VDD.n11337 VDD.n563 2.2505
R26944 VDD.n11339 VDD.n11338 2.2505
R26945 VDD.n11340 VDD.n562 2.2505
R26946 VDD.n11342 VDD.n11341 2.2505
R26947 VDD.n11343 VDD.n561 2.2505
R26948 VDD.n11345 VDD.n11344 2.2505
R26949 VDD.n11346 VDD.n560 2.2505
R26950 VDD.n11348 VDD.n11347 2.2505
R26951 VDD.n11349 VDD.n559 2.2505
R26952 VDD.n11351 VDD.n11350 2.2505
R26953 VDD.n11352 VDD.n558 2.2505
R26954 VDD.n11354 VDD.n11353 2.2505
R26955 VDD.n11355 VDD.n557 2.2505
R26956 VDD.n11357 VDD.n11356 2.2505
R26957 VDD.n11358 VDD.n556 2.2505
R26958 VDD.n11360 VDD.n11359 2.2505
R26959 VDD.n11361 VDD.n555 2.2505
R26960 VDD.n11363 VDD.n11362 2.2505
R26961 VDD.n11364 VDD.n554 2.2505
R26962 VDD.n11366 VDD.n11365 2.2505
R26963 VDD.n11367 VDD.n553 2.2505
R26964 VDD.n11369 VDD.n11368 2.2505
R26965 VDD.n11370 VDD.n552 2.2505
R26966 VDD.n11372 VDD.n11371 2.2505
R26967 VDD.n11373 VDD.n551 2.2505
R26968 VDD.n11375 VDD.n11374 2.2505
R26969 VDD.n11376 VDD.n550 2.2505
R26970 VDD.n11378 VDD.n11377 2.2505
R26971 VDD.n11379 VDD.n549 2.2505
R26972 VDD.n11381 VDD.n11380 2.2505
R26973 VDD.n11382 VDD.n548 2.2505
R26974 VDD.n11384 VDD.n11383 2.2505
R26975 VDD.n11385 VDD.n547 2.2505
R26976 VDD.n11387 VDD.n11386 2.2505
R26977 VDD.n11388 VDD.n546 2.2505
R26978 VDD.n11390 VDD.n11389 2.2505
R26979 VDD.n11391 VDD.n545 2.2505
R26980 VDD.n11393 VDD.n11392 2.2505
R26981 VDD.n11394 VDD.n544 2.2505
R26982 VDD.n11396 VDD.n11395 2.2505
R26983 VDD.n11397 VDD.n543 2.2505
R26984 VDD.n11399 VDD.n11398 2.2505
R26985 VDD.n11400 VDD.n542 2.2505
R26986 VDD.n11402 VDD.n11401 2.2505
R26987 VDD.n11403 VDD.n541 2.2505
R26988 VDD.n11405 VDD.n11404 2.2505
R26989 VDD.n11406 VDD.n540 2.2505
R26990 VDD.n11408 VDD.n11407 2.2505
R26991 VDD.n11409 VDD.n539 2.2505
R26992 VDD.n11411 VDD.n11410 2.2505
R26993 VDD.n11412 VDD.n538 2.2505
R26994 VDD.n11414 VDD.n11413 2.2505
R26995 VDD.n11415 VDD.n537 2.2505
R26996 VDD.n11417 VDD.n11416 2.2505
R26997 VDD.n11418 VDD.n536 2.2505
R26998 VDD.n11420 VDD.n11419 2.2505
R26999 VDD.n11421 VDD.n535 2.2505
R27000 VDD.n11423 VDD.n11422 2.2505
R27001 VDD.n11424 VDD.n534 2.2505
R27002 VDD.n11426 VDD.n11425 2.2505
R27003 VDD.n11427 VDD.n533 2.2505
R27004 VDD.n11429 VDD.n11428 2.2505
R27005 VDD.n11430 VDD.n532 2.2505
R27006 VDD.n11432 VDD.n11431 2.2505
R27007 VDD.n11433 VDD.n531 2.2505
R27008 VDD.n11435 VDD.n11434 2.2505
R27009 VDD.n11436 VDD.n530 2.2505
R27010 VDD.n11438 VDD.n11437 2.2505
R27011 VDD.n11439 VDD.n529 2.2505
R27012 VDD.n11441 VDD.n11440 2.2505
R27013 VDD.n11442 VDD.n528 2.2505
R27014 VDD.n11444 VDD.n11443 2.2505
R27015 VDD.n11445 VDD.n527 2.2505
R27016 VDD.n11447 VDD.n11446 2.2505
R27017 VDD.n11448 VDD.n526 2.2505
R27018 VDD.n11450 VDD.n11449 2.2505
R27019 VDD.n11451 VDD.n525 2.2505
R27020 VDD.n11453 VDD.n11452 2.2505
R27021 VDD.n11454 VDD.n524 2.2505
R27022 VDD.n11456 VDD.n11455 2.2505
R27023 VDD.n11457 VDD.n523 2.2505
R27024 VDD.n11459 VDD.n11458 2.2505
R27025 VDD.n11460 VDD.n522 2.2505
R27026 VDD.n11462 VDD.n11461 2.2505
R27027 VDD.n11463 VDD.n521 2.2505
R27028 VDD.n11465 VDD.n11464 2.2505
R27029 VDD.n11466 VDD.n520 2.2505
R27030 VDD.n11468 VDD.n11467 2.2505
R27031 VDD.n11469 VDD.n519 2.2505
R27032 VDD.n11471 VDD.n11470 2.2505
R27033 VDD.n11472 VDD.n518 2.2505
R27034 VDD.n11474 VDD.n11473 2.2505
R27035 VDD.n11475 VDD.n517 2.2505
R27036 VDD.n11477 VDD.n11476 2.2505
R27037 VDD.n11478 VDD.n516 2.2505
R27038 VDD.n11480 VDD.n11479 2.2505
R27039 VDD.n11481 VDD.n515 2.2505
R27040 VDD.n11483 VDD.n11482 2.2505
R27041 VDD.n11484 VDD.n514 2.2505
R27042 VDD.n11486 VDD.n11485 2.2505
R27043 VDD.n11487 VDD.n513 2.2505
R27044 VDD.n11489 VDD.n11488 2.2505
R27045 VDD.n11490 VDD.n512 2.2505
R27046 VDD.n11492 VDD.n11491 2.2505
R27047 VDD.n11493 VDD.n511 2.2505
R27048 VDD.n11495 VDD.n11494 2.2505
R27049 VDD.n11496 VDD.n510 2.2505
R27050 VDD.n11498 VDD.n11497 2.2505
R27051 VDD.n11499 VDD.n509 2.2505
R27052 VDD.n11501 VDD.n11500 2.2505
R27053 VDD.n11502 VDD.n508 2.2505
R27054 VDD.n11504 VDD.n11503 2.2505
R27055 VDD.n11505 VDD.n507 2.2505
R27056 VDD.n11507 VDD.n11506 2.2505
R27057 VDD.n11508 VDD.n506 2.2505
R27058 VDD.n11510 VDD.n11509 2.2505
R27059 VDD.n11511 VDD.n505 2.2505
R27060 VDD.n11513 VDD.n11512 2.2505
R27061 VDD.n11514 VDD.n504 2.2505
R27062 VDD.n11516 VDD.n11515 2.2505
R27063 VDD.n11517 VDD.n503 2.2505
R27064 VDD.n11519 VDD.n11518 2.2505
R27065 VDD.n11520 VDD.n502 2.2505
R27066 VDD.n11522 VDD.n11521 2.2505
R27067 VDD.n11523 VDD.n501 2.2505
R27068 VDD.n11525 VDD.n11524 2.2505
R27069 VDD.n11526 VDD.n500 2.2505
R27070 VDD.n11528 VDD.n11527 2.2505
R27071 VDD.n11529 VDD.n499 2.2505
R27072 VDD.n11531 VDD.n11530 2.2505
R27073 VDD.n11532 VDD.n498 2.2505
R27074 VDD.n11534 VDD.n11533 2.2505
R27075 VDD.n11535 VDD.n497 2.2505
R27076 VDD.n11537 VDD.n11536 2.2505
R27077 VDD.n11538 VDD.n496 2.2505
R27078 VDD.n11540 VDD.n11539 2.2505
R27079 VDD.n11541 VDD.n495 2.2505
R27080 VDD.n11543 VDD.n11542 2.2505
R27081 VDD.n11544 VDD.n494 2.2505
R27082 VDD.n11546 VDD.n11545 2.2505
R27083 VDD.n11547 VDD.n493 2.2505
R27084 VDD.n11549 VDD.n11548 2.2505
R27085 VDD.n11550 VDD.n492 2.2505
R27086 VDD.n11552 VDD.n11551 2.2505
R27087 VDD.n11553 VDD.n491 2.2505
R27088 VDD.n11555 VDD.n11554 2.2505
R27089 VDD.n11556 VDD.n490 2.2505
R27090 VDD.n11558 VDD.n11557 2.2505
R27091 VDD.n11559 VDD.n489 2.2505
R27092 VDD.n11561 VDD.n11560 2.2505
R27093 VDD.n11562 VDD.n488 2.2505
R27094 VDD.n11564 VDD.n11563 2.2505
R27095 VDD.n11565 VDD.n487 2.2505
R27096 VDD.n11567 VDD.n11566 2.2505
R27097 VDD.n11568 VDD.n486 2.2505
R27098 VDD.n11570 VDD.n11569 2.2505
R27099 VDD.n11571 VDD.n485 2.2505
R27100 VDD.n11573 VDD.n11572 2.2505
R27101 VDD.n11574 VDD.n484 2.2505
R27102 VDD.n11576 VDD.n11575 2.2505
R27103 VDD.n11577 VDD.n483 2.2505
R27104 VDD.n11579 VDD.n11578 2.2505
R27105 VDD.n11580 VDD.n482 2.2505
R27106 VDD.n11582 VDD.n11581 2.2505
R27107 VDD.n11583 VDD.n481 2.2505
R27108 VDD.n11585 VDD.n11584 2.2505
R27109 VDD.n11586 VDD.n480 2.2505
R27110 VDD.n11588 VDD.n11587 2.2505
R27111 VDD.n11589 VDD.n479 2.2505
R27112 VDD.n11591 VDD.n11590 2.2505
R27113 VDD.n11592 VDD.n478 2.2505
R27114 VDD.n11594 VDD.n11593 2.2505
R27115 VDD.n11595 VDD.n477 2.2505
R27116 VDD.n11597 VDD.n11596 2.2505
R27117 VDD.n11598 VDD.n476 2.2505
R27118 VDD.n11600 VDD.n11599 2.2505
R27119 VDD.n11601 VDD.n475 2.2505
R27120 VDD.n11603 VDD.n11602 2.2505
R27121 VDD.n11604 VDD.n474 2.2505
R27122 VDD.n11606 VDD.n11605 2.2505
R27123 VDD.n11607 VDD.n473 2.2505
R27124 VDD.n11609 VDD.n11608 2.2505
R27125 VDD.n11610 VDD.n472 2.2505
R27126 VDD.n11612 VDD.n11611 2.2505
R27127 VDD.n11613 VDD.n471 2.2505
R27128 VDD.n11615 VDD.n11614 2.2505
R27129 VDD.n11616 VDD.n470 2.2505
R27130 VDD.n11618 VDD.n11617 2.2505
R27131 VDD.n11619 VDD.n469 2.2505
R27132 VDD.n11621 VDD.n11620 2.2505
R27133 VDD.n11622 VDD.n468 2.2505
R27134 VDD.n11624 VDD.n11623 2.2505
R27135 VDD.n11625 VDD.n467 2.2505
R27136 VDD.n11627 VDD.n11626 2.2505
R27137 VDD.n11628 VDD.n466 2.2505
R27138 VDD.n11630 VDD.n11629 2.2505
R27139 VDD.n11631 VDD.n465 2.2505
R27140 VDD.n11633 VDD.n11632 2.2505
R27141 VDD.n11634 VDD.n464 2.2505
R27142 VDD.n11636 VDD.n11635 2.2505
R27143 VDD.n11637 VDD.n463 2.2505
R27144 VDD.n11639 VDD.n11638 2.2505
R27145 VDD.n11640 VDD.n462 2.2505
R27146 VDD.n11642 VDD.n11641 2.2505
R27147 VDD.n11643 VDD.n461 2.2505
R27148 VDD.n11645 VDD.n11644 2.2505
R27149 VDD.n11646 VDD.n460 2.2505
R27150 VDD.n11648 VDD.n11647 2.2505
R27151 VDD.n11649 VDD.n459 2.2505
R27152 VDD.n11651 VDD.n11650 2.2505
R27153 VDD.n11652 VDD.n458 2.2505
R27154 VDD.n11654 VDD.n11653 2.2505
R27155 VDD.n11655 VDD.n457 2.2505
R27156 VDD.n11657 VDD.n11656 2.2505
R27157 VDD.n11658 VDD.n456 2.2505
R27158 VDD.n11660 VDD.n11659 2.2505
R27159 VDD.n11661 VDD.n455 2.2505
R27160 VDD.n11663 VDD.n11662 2.2505
R27161 VDD.n11664 VDD.n454 2.2505
R27162 VDD.n11666 VDD.n11665 2.2505
R27163 VDD.n11667 VDD.n453 2.2505
R27164 VDD.n11669 VDD.n11668 2.2505
R27165 VDD.n11670 VDD.n452 2.2505
R27166 VDD.n11672 VDD.n11671 2.2505
R27167 VDD.n11673 VDD.n451 2.2505
R27168 VDD.n11675 VDD.n11674 2.2505
R27169 VDD.n11676 VDD.n450 2.2505
R27170 VDD.n11678 VDD.n11677 2.2505
R27171 VDD.n11679 VDD.n449 2.2505
R27172 VDD.n11681 VDD.n11680 2.2505
R27173 VDD.n11682 VDD.n448 2.2505
R27174 VDD.n11684 VDD.n11683 2.2505
R27175 VDD.n11685 VDD.n447 2.2505
R27176 VDD.n11687 VDD.n11686 2.2505
R27177 VDD.n11688 VDD.n446 2.2505
R27178 VDD.n11690 VDD.n11689 2.2505
R27179 VDD.n11691 VDD.n445 2.2505
R27180 VDD.n11693 VDD.n11692 2.2505
R27181 VDD.n11694 VDD.n444 2.2505
R27182 VDD.n11696 VDD.n11695 2.2505
R27183 VDD.n11697 VDD.n443 2.2505
R27184 VDD.n11699 VDD.n11698 2.2505
R27185 VDD.n11700 VDD.n442 2.2505
R27186 VDD.n11702 VDD.n11701 2.2505
R27187 VDD.n11703 VDD.n441 2.2505
R27188 VDD.n11705 VDD.n11704 2.2505
R27189 VDD.n11706 VDD.n440 2.2505
R27190 VDD.n11708 VDD.n11707 2.2505
R27191 VDD.n11709 VDD.n439 2.2505
R27192 VDD.n11711 VDD.n11710 2.2505
R27193 VDD.n11712 VDD.n438 2.2505
R27194 VDD.n11714 VDD.n11713 2.2505
R27195 VDD.n11715 VDD.n437 2.2505
R27196 VDD.n11717 VDD.n11716 2.2505
R27197 VDD.n11718 VDD.n436 2.2505
R27198 VDD.n11720 VDD.n11719 2.2505
R27199 VDD.n11721 VDD.n435 2.2505
R27200 VDD.n11723 VDD.n11722 2.2505
R27201 VDD.n11724 VDD.n434 2.2505
R27202 VDD.n11726 VDD.n11725 2.2505
R27203 VDD.n11727 VDD.n433 2.2505
R27204 VDD.n11729 VDD.n11728 2.2505
R27205 VDD.n11730 VDD.n432 2.2505
R27206 VDD.n11732 VDD.n11731 2.2505
R27207 VDD.n11733 VDD.n431 2.2505
R27208 VDD.n11735 VDD.n11734 2.2505
R27209 VDD.n11736 VDD.n430 2.2505
R27210 VDD.n11738 VDD.n11737 2.2505
R27211 VDD.n11739 VDD.n429 2.2505
R27212 VDD.n11741 VDD.n11740 2.2505
R27213 VDD.n11742 VDD.n428 2.2505
R27214 VDD.n11744 VDD.n11743 2.2505
R27215 VDD.n11745 VDD.n427 2.2505
R27216 VDD.n11747 VDD.n11746 2.2505
R27217 VDD.n11748 VDD.n426 2.2505
R27218 VDD.n11750 VDD.n11749 2.2505
R27219 VDD.n11751 VDD.n425 2.2505
R27220 VDD.n11753 VDD.n11752 2.2505
R27221 VDD.n11754 VDD.n424 2.2505
R27222 VDD.n11756 VDD.n11755 2.2505
R27223 VDD.n11757 VDD.n423 2.2505
R27224 VDD.n11759 VDD.n11758 2.2505
R27225 VDD.n11760 VDD.n422 2.2505
R27226 VDD.n11762 VDD.n11761 2.2505
R27227 VDD.n11763 VDD.n421 2.2505
R27228 VDD.n11765 VDD.n11764 2.2505
R27229 VDD.n11766 VDD.n420 2.2505
R27230 VDD.n11768 VDD.n11767 2.2505
R27231 VDD.n11769 VDD.n419 2.2505
R27232 VDD.n11771 VDD.n11770 2.2505
R27233 VDD.n11772 VDD.n418 2.2505
R27234 VDD.n11774 VDD.n11773 2.2505
R27235 VDD.n11775 VDD.n417 2.2505
R27236 VDD.n11777 VDD.n11776 2.2505
R27237 VDD.n11778 VDD.n416 2.2505
R27238 VDD.n11780 VDD.n11779 2.2505
R27239 VDD.n11781 VDD.n415 2.2505
R27240 VDD.n11783 VDD.n11782 2.2505
R27241 VDD.n11784 VDD.n414 2.2505
R27242 VDD.n11786 VDD.n11785 2.2505
R27243 VDD.n11787 VDD.n413 2.2505
R27244 VDD.n11789 VDD.n11788 2.2505
R27245 VDD.n11790 VDD.n412 2.2505
R27246 VDD.n11792 VDD.n11791 2.2505
R27247 VDD.n11793 VDD.n411 2.2505
R27248 VDD.n11795 VDD.n11794 2.2505
R27249 VDD.n11796 VDD.n410 2.2505
R27250 VDD.n11798 VDD.n11797 2.2505
R27251 VDD.n11799 VDD.n409 2.2505
R27252 VDD.n11801 VDD.n11800 2.2505
R27253 VDD.n11802 VDD.n408 2.2505
R27254 VDD.n11804 VDD.n11803 2.2505
R27255 VDD.n11805 VDD.n407 2.2505
R27256 VDD.n11807 VDD.n11806 2.2505
R27257 VDD.n11808 VDD.n406 2.2505
R27258 VDD.n11810 VDD.n11809 2.2505
R27259 VDD.n11811 VDD.n405 2.2505
R27260 VDD.n2967 VDD.n2966 2.2505
R27261 VDD.n10762 VDD.n10761 2.2505
R27262 VDD.n10763 VDD.n2062 2.2505
R27263 VDD.n10765 VDD.n10764 2.2505
R27264 VDD.n8253 VDD.n2061 2.2505
R27265 VDD.n8252 VDD.n8251 2.2505
R27266 VDD.n8248 VDD.n2063 2.2505
R27267 VDD.n8247 VDD.n8246 2.2505
R27268 VDD.n8245 VDD.n8244 2.2505
R27269 VDD.n8243 VDD.n2065 2.2505
R27270 VDD.n8242 VDD.n8241 2.2505
R27271 VDD.n8240 VDD.n2066 2.2505
R27272 VDD.n8239 VDD.n8238 2.2505
R27273 VDD.n8235 VDD.n2067 2.2505
R27274 VDD.n8234 VDD.n8233 2.2505
R27275 VDD.n8232 VDD.n2068 2.2505
R27276 VDD.n8231 VDD.n8230 2.2505
R27277 VDD.n8228 VDD.n2069 2.2505
R27278 VDD.n8227 VDD.n8226 2.2505
R27279 VDD.n8225 VDD.n2070 2.2505
R27280 VDD.n8224 VDD.n8223 2.2505
R27281 VDD.n8221 VDD.n2071 2.2505
R27282 VDD.n8220 VDD.n8219 2.2505
R27283 VDD.n8218 VDD.n2072 2.2505
R27284 VDD.n8217 VDD.n8216 2.2505
R27285 VDD.n8213 VDD.n2073 2.2505
R27286 VDD.n8212 VDD.n8211 2.2505
R27287 VDD.n8210 VDD.n8209 2.2505
R27288 VDD.n8208 VDD.n2075 2.2505
R27289 VDD.n8207 VDD.n8206 2.2505
R27290 VDD.n8205 VDD.n2076 2.2505
R27291 VDD.n8204 VDD.n8203 2.2505
R27292 VDD.n8200 VDD.n2077 2.2505
R27293 VDD.n8199 VDD.n8198 2.2505
R27294 VDD.n8197 VDD.n8196 2.2505
R27295 VDD.n8195 VDD.n2079 2.2505
R27296 VDD.n8194 VDD.n8193 2.2505
R27297 VDD.n8192 VDD.n2080 2.2505
R27298 VDD.n8191 VDD.n8190 2.2505
R27299 VDD.n8189 VDD.n2081 2.2505
R27300 VDD.n8187 VDD.n8186 2.2505
R27301 VDD.n8185 VDD.n2082 2.2505
R27302 VDD.n8184 VDD.n8183 2.2505
R27303 VDD.n8180 VDD.n2083 2.2505
R27304 VDD.n8179 VDD.n8178 2.2505
R27305 VDD.n8177 VDD.n2084 2.2505
R27306 VDD.n8176 VDD.n8175 2.2505
R27307 VDD.n8174 VDD.n2085 2.2505
R27308 VDD.n8172 VDD.n8171 2.2505
R27309 VDD.n8170 VDD.n2086 2.2505
R27310 VDD.n8169 VDD.n8168 2.2505
R27311 VDD.n2088 VDD.n2087 2.2505
R27312 VDD.n7304 VDD.n7303 2.2505
R27313 VDD.n7306 VDD.n7305 2.2505
R27314 VDD.n7307 VDD.n7302 2.2505
R27315 VDD.n7309 VDD.n7308 2.2505
R27316 VDD.n7310 VDD.n7301 2.2505
R27317 VDD.n7312 VDD.n7311 2.2505
R27318 VDD.n7313 VDD.n7300 2.2505
R27319 VDD.n7315 VDD.n7314 2.2505
R27320 VDD.n7316 VDD.n7299 2.2505
R27321 VDD.n7318 VDD.n7317 2.2505
R27322 VDD.n7319 VDD.n7298 2.2505
R27323 VDD.n7321 VDD.n7320 2.2505
R27324 VDD.n7322 VDD.n7297 2.2505
R27325 VDD.n7324 VDD.n7323 2.2505
R27326 VDD.n7325 VDD.n7296 2.2505
R27327 VDD.n7327 VDD.n7326 2.2505
R27328 VDD.n7328 VDD.n7295 2.2505
R27329 VDD.n7330 VDD.n7329 2.2505
R27330 VDD.n7331 VDD.n7294 2.2505
R27331 VDD.n7333 VDD.n7332 2.2505
R27332 VDD.n7334 VDD.n7293 2.2505
R27333 VDD.n7336 VDD.n7335 2.2505
R27334 VDD.n7337 VDD.n7292 2.2505
R27335 VDD.n7339 VDD.n7338 2.2505
R27336 VDD.n7340 VDD.n7291 2.2505
R27337 VDD.n7342 VDD.n7341 2.2505
R27338 VDD.n7343 VDD.n7290 2.2505
R27339 VDD.n7345 VDD.n7344 2.2505
R27340 VDD.n7346 VDD.n7289 2.2505
R27341 VDD.n7348 VDD.n7347 2.2505
R27342 VDD.n7349 VDD.n7288 2.2505
R27343 VDD.n7351 VDD.n7350 2.2505
R27344 VDD.n7352 VDD.n7287 2.2505
R27345 VDD.n7354 VDD.n7353 2.2505
R27346 VDD.n7355 VDD.n7286 2.2505
R27347 VDD.n7357 VDD.n7356 2.2505
R27348 VDD.n7358 VDD.n7285 2.2505
R27349 VDD.n7360 VDD.n7359 2.2505
R27350 VDD.n7361 VDD.n7284 2.2505
R27351 VDD.n7363 VDD.n7362 2.2505
R27352 VDD.n7364 VDD.n7283 2.2505
R27353 VDD.n7366 VDD.n7365 2.2505
R27354 VDD.n7367 VDD.n7282 2.2505
R27355 VDD.n7369 VDD.n7368 2.2505
R27356 VDD.n7370 VDD.n7281 2.2505
R27357 VDD.n7372 VDD.n7371 2.2505
R27358 VDD.n7373 VDD.n7280 2.2505
R27359 VDD.n7375 VDD.n7374 2.2505
R27360 VDD.n7376 VDD.n7279 2.2505
R27361 VDD.n7378 VDD.n7377 2.2505
R27362 VDD.n7379 VDD.n7278 2.2505
R27363 VDD.n7381 VDD.n7380 2.2505
R27364 VDD.n7382 VDD.n7277 2.2505
R27365 VDD.n7384 VDD.n7383 2.2505
R27366 VDD.n7385 VDD.n7276 2.2505
R27367 VDD.n7387 VDD.n7386 2.2505
R27368 VDD.n7388 VDD.n7275 2.2505
R27369 VDD.n7390 VDD.n7389 2.2505
R27370 VDD.n7391 VDD.n7274 2.2505
R27371 VDD.n7393 VDD.n7392 2.2505
R27372 VDD.n7394 VDD.n7273 2.2505
R27373 VDD.n7396 VDD.n7395 2.2505
R27374 VDD.n7397 VDD.n7272 2.2505
R27375 VDD.n7399 VDD.n7398 2.2505
R27376 VDD.n7400 VDD.n7271 2.2505
R27377 VDD.n7402 VDD.n7401 2.2505
R27378 VDD.n7403 VDD.n7270 2.2505
R27379 VDD.n7405 VDD.n7404 2.2505
R27380 VDD.n7406 VDD.n7269 2.2505
R27381 VDD.n7408 VDD.n7407 2.2505
R27382 VDD.n7409 VDD.n7268 2.2505
R27383 VDD.n7411 VDD.n7410 2.2505
R27384 VDD.n7412 VDD.n7267 2.2505
R27385 VDD.n7414 VDD.n7413 2.2505
R27386 VDD.n7415 VDD.n7266 2.2505
R27387 VDD.n7417 VDD.n7416 2.2505
R27388 VDD.n7418 VDD.n7265 2.2505
R27389 VDD.n7420 VDD.n7419 2.2505
R27390 VDD.n7421 VDD.n7264 2.2505
R27391 VDD.n7423 VDD.n7422 2.2505
R27392 VDD.n7424 VDD.n7263 2.2505
R27393 VDD.n7426 VDD.n7425 2.2505
R27394 VDD.n7427 VDD.n7262 2.2505
R27395 VDD.n7429 VDD.n7428 2.2505
R27396 VDD.n7430 VDD.n7261 2.2505
R27397 VDD.n7432 VDD.n7431 2.2505
R27398 VDD.n7433 VDD.n7260 2.2505
R27399 VDD.n7435 VDD.n7434 2.2505
R27400 VDD.n7436 VDD.n7259 2.2505
R27401 VDD.n7438 VDD.n7437 2.2505
R27402 VDD.n7439 VDD.n7258 2.2505
R27403 VDD.n7441 VDD.n7440 2.2505
R27404 VDD.n7442 VDD.n7257 2.2505
R27405 VDD.n7444 VDD.n7443 2.2505
R27406 VDD.n7445 VDD.n7256 2.2505
R27407 VDD.n7447 VDD.n7446 2.2505
R27408 VDD.n7448 VDD.n7255 2.2505
R27409 VDD.n7450 VDD.n7449 2.2505
R27410 VDD.n7451 VDD.n7254 2.2505
R27411 VDD.n7453 VDD.n7452 2.2505
R27412 VDD.n7454 VDD.n7253 2.2505
R27413 VDD.n7456 VDD.n7455 2.2505
R27414 VDD.n7457 VDD.n7252 2.2505
R27415 VDD.n7459 VDD.n7458 2.2505
R27416 VDD.n7460 VDD.n7251 2.2505
R27417 VDD.n7462 VDD.n7461 2.2505
R27418 VDD.n7463 VDD.n7250 2.2505
R27419 VDD.n7465 VDD.n7464 2.2505
R27420 VDD.n7466 VDD.n7249 2.2505
R27421 VDD.n7468 VDD.n7467 2.2505
R27422 VDD.n7469 VDD.n7248 2.2505
R27423 VDD.n7471 VDD.n7470 2.2505
R27424 VDD.n7472 VDD.n7247 2.2505
R27425 VDD.n7474 VDD.n7473 2.2505
R27426 VDD.n7475 VDD.n7246 2.2505
R27427 VDD.n7477 VDD.n7476 2.2505
R27428 VDD.n7478 VDD.n7245 2.2505
R27429 VDD.n7480 VDD.n7479 2.2505
R27430 VDD.n7481 VDD.n7244 2.2505
R27431 VDD.n7483 VDD.n7482 2.2505
R27432 VDD.n7484 VDD.n7243 2.2505
R27433 VDD.n7486 VDD.n7485 2.2505
R27434 VDD.n7487 VDD.n7242 2.2505
R27435 VDD.n7489 VDD.n7488 2.2505
R27436 VDD.n7490 VDD.n7241 2.2505
R27437 VDD.n7492 VDD.n7491 2.2505
R27438 VDD.n7493 VDD.n7240 2.2505
R27439 VDD.n7495 VDD.n7494 2.2505
R27440 VDD.n7496 VDD.n7239 2.2505
R27441 VDD.n7498 VDD.n7497 2.2505
R27442 VDD.n7499 VDD.n7238 2.2505
R27443 VDD.n7501 VDD.n7500 2.2505
R27444 VDD.n7502 VDD.n7237 2.2505
R27445 VDD.n7504 VDD.n7503 2.2505
R27446 VDD.n7505 VDD.n7236 2.2505
R27447 VDD.n7507 VDD.n7506 2.2505
R27448 VDD.n7508 VDD.n7235 2.2505
R27449 VDD.n7510 VDD.n7509 2.2505
R27450 VDD.n7511 VDD.n7234 2.2505
R27451 VDD.n7513 VDD.n7512 2.2505
R27452 VDD.n7514 VDD.n7233 2.2505
R27453 VDD.n7516 VDD.n7515 2.2505
R27454 VDD.n7517 VDD.n7232 2.2505
R27455 VDD.n7519 VDD.n7518 2.2505
R27456 VDD.n7520 VDD.n7231 2.2505
R27457 VDD.n7522 VDD.n7521 2.2505
R27458 VDD.n7523 VDD.n7230 2.2505
R27459 VDD.n7525 VDD.n7524 2.2505
R27460 VDD.n7526 VDD.n7229 2.2505
R27461 VDD.n7528 VDD.n7527 2.2505
R27462 VDD.n7529 VDD.n7228 2.2505
R27463 VDD.n7531 VDD.n7530 2.2505
R27464 VDD.n7532 VDD.n7227 2.2505
R27465 VDD.n7534 VDD.n7533 2.2505
R27466 VDD.n7535 VDD.n7226 2.2505
R27467 VDD.n7537 VDD.n7536 2.2505
R27468 VDD.n7538 VDD.n7225 2.2505
R27469 VDD.n7540 VDD.n7539 2.2505
R27470 VDD.n7541 VDD.n7224 2.2505
R27471 VDD.n7543 VDD.n7542 2.2505
R27472 VDD.n7544 VDD.n7223 2.2505
R27473 VDD.n7546 VDD.n7545 2.2505
R27474 VDD.n7547 VDD.n7222 2.2505
R27475 VDD.n7549 VDD.n7548 2.2505
R27476 VDD.n7550 VDD.n7221 2.2505
R27477 VDD.n7552 VDD.n7551 2.2505
R27478 VDD.n7553 VDD.n7220 2.2505
R27479 VDD.n7555 VDD.n7554 2.2505
R27480 VDD.n7556 VDD.n7219 2.2505
R27481 VDD.n7558 VDD.n7557 2.2505
R27482 VDD.n7559 VDD.n7218 2.2505
R27483 VDD.n7561 VDD.n7560 2.2505
R27484 VDD.n7562 VDD.n7217 2.2505
R27485 VDD.n7564 VDD.n7563 2.2505
R27486 VDD.n7565 VDD.n7216 2.2505
R27487 VDD.n7567 VDD.n7566 2.2505
R27488 VDD.n7568 VDD.n7215 2.2505
R27489 VDD.n7570 VDD.n7569 2.2505
R27490 VDD.n7571 VDD.n7214 2.2505
R27491 VDD.n7573 VDD.n7572 2.2505
R27492 VDD.n7574 VDD.n7213 2.2505
R27493 VDD.n7576 VDD.n7575 2.2505
R27494 VDD.n7577 VDD.n7212 2.2505
R27495 VDD.n7579 VDD.n7578 2.2505
R27496 VDD.n7580 VDD.n7211 2.2505
R27497 VDD.n7582 VDD.n7581 2.2505
R27498 VDD.n7583 VDD.n7210 2.2505
R27499 VDD.n7585 VDD.n7584 2.2505
R27500 VDD.n7586 VDD.n7209 2.2505
R27501 VDD.n7588 VDD.n7587 2.2505
R27502 VDD.n7589 VDD.n7208 2.2505
R27503 VDD.n7591 VDD.n7590 2.2505
R27504 VDD.n7592 VDD.n7207 2.2505
R27505 VDD.n7594 VDD.n7593 2.2505
R27506 VDD.n7595 VDD.n7206 2.2505
R27507 VDD.n7597 VDD.n7596 2.2505
R27508 VDD.n7598 VDD.n7205 2.2505
R27509 VDD.n7600 VDD.n7599 2.2505
R27510 VDD.n7601 VDD.n7204 2.2505
R27511 VDD.n7603 VDD.n7602 2.2505
R27512 VDD.n7604 VDD.n7203 2.2505
R27513 VDD.n7606 VDD.n7605 2.2505
R27514 VDD.n7607 VDD.n7202 2.2505
R27515 VDD.n7609 VDD.n7608 2.2505
R27516 VDD.n7610 VDD.n7201 2.2505
R27517 VDD.n7612 VDD.n7611 2.2505
R27518 VDD.n7613 VDD.n7200 2.2505
R27519 VDD.n7615 VDD.n7614 2.2505
R27520 VDD.n7616 VDD.n7199 2.2505
R27521 VDD.n7618 VDD.n7617 2.2505
R27522 VDD.n7619 VDD.n7198 2.2505
R27523 VDD.n7621 VDD.n7620 2.2505
R27524 VDD.n7622 VDD.n7197 2.2505
R27525 VDD.n7624 VDD.n7623 2.2505
R27526 VDD.n7625 VDD.n7196 2.2505
R27527 VDD.n7627 VDD.n7626 2.2505
R27528 VDD.n7628 VDD.n7195 2.2505
R27529 VDD.n7630 VDD.n7629 2.2505
R27530 VDD.n7631 VDD.n7194 2.2505
R27531 VDD.n7633 VDD.n7632 2.2505
R27532 VDD.n7634 VDD.n7193 2.2505
R27533 VDD.n7636 VDD.n7635 2.2505
R27534 VDD.n7637 VDD.n7192 2.2505
R27535 VDD.n7639 VDD.n7638 2.2505
R27536 VDD.n7640 VDD.n7191 2.2505
R27537 VDD.n7642 VDD.n7641 2.2505
R27538 VDD.n7643 VDD.n7190 2.2505
R27539 VDD.n7645 VDD.n7644 2.2505
R27540 VDD.n7646 VDD.n7189 2.2505
R27541 VDD.n7648 VDD.n7647 2.2505
R27542 VDD.n7649 VDD.n7188 2.2505
R27543 VDD.n7651 VDD.n7650 2.2505
R27544 VDD.n7652 VDD.n7187 2.2505
R27545 VDD.n7654 VDD.n7653 2.2505
R27546 VDD.n7655 VDD.n7186 2.2505
R27547 VDD.n7657 VDD.n7656 2.2505
R27548 VDD.n7658 VDD.n7185 2.2505
R27549 VDD.n7660 VDD.n7659 2.2505
R27550 VDD.n7661 VDD.n7184 2.2505
R27551 VDD.n7663 VDD.n7662 2.2505
R27552 VDD.n7664 VDD.n7183 2.2505
R27553 VDD.n7666 VDD.n7665 2.2505
R27554 VDD.n7667 VDD.n7182 2.2505
R27555 VDD.n7669 VDD.n7668 2.2505
R27556 VDD.n7670 VDD.n7181 2.2505
R27557 VDD.n7672 VDD.n7671 2.2505
R27558 VDD.n7673 VDD.n7180 2.2505
R27559 VDD.n7675 VDD.n7674 2.2505
R27560 VDD.n7676 VDD.n7179 2.2505
R27561 VDD.n7678 VDD.n7677 2.2505
R27562 VDD.n7679 VDD.n7178 2.2505
R27563 VDD.n7681 VDD.n7680 2.2505
R27564 VDD.n7682 VDD.n2293 2.2505
R27565 VDD.n7685 VDD.n7684 2.2505
R27566 VDD.n7750 VDD.n7749 2.2505
R27567 VDD.n7751 VDD.n2268 2.2505
R27568 VDD.n7753 VDD.n7752 2.2505
R27569 VDD.n7754 VDD.n2267 2.2505
R27570 VDD.n7756 VDD.n7755 2.2505
R27571 VDD.n7757 VDD.n2266 2.2505
R27572 VDD.n7759 VDD.n7758 2.2505
R27573 VDD.n7761 VDD.n2264 2.2505
R27574 VDD.n7763 VDD.n7762 2.2505
R27575 VDD.n7764 VDD.n2263 2.2505
R27576 VDD.n7766 VDD.n7765 2.2505
R27577 VDD.n7767 VDD.n2262 2.2505
R27578 VDD.n7769 VDD.n7768 2.2505
R27579 VDD.n7770 VDD.n2261 2.2505
R27580 VDD.n7772 VDD.n7771 2.2505
R27581 VDD.n7773 VDD.n2259 2.2505
R27582 VDD.n7775 VDD.n7774 2.2505
R27583 VDD.n7776 VDD.n2258 2.2505
R27584 VDD.n7778 VDD.n7777 2.2505
R27585 VDD.n7779 VDD.n2257 2.2505
R27586 VDD.n7782 VDD.n7781 2.2505
R27587 VDD.n7783 VDD.n2256 2.2505
R27588 VDD.n7785 VDD.n7784 2.2505
R27589 VDD.n7786 VDD.n2255 2.2505
R27590 VDD.n7788 VDD.n7787 2.2505
R27591 VDD.n7789 VDD.n2254 2.2505
R27592 VDD.n7791 VDD.n7790 2.2505
R27593 VDD.n7792 VDD.n2253 2.2505
R27594 VDD.n7794 VDD.n7793 2.2505
R27595 VDD.n7796 VDD.n7795 2.2505
R27596 VDD.n7797 VDD.n2251 2.2505
R27597 VDD.n7799 VDD.n7798 2.2505
R27598 VDD.n7801 VDD.n7800 2.2505
R27599 VDD.n7802 VDD.n2249 2.2505
R27600 VDD.n7804 VDD.n7803 2.2505
R27601 VDD.n7805 VDD.n2248 2.2505
R27602 VDD.n7807 VDD.n7806 2.2505
R27603 VDD.n7808 VDD.n2247 2.2505
R27604 VDD.n7811 VDD.n7810 2.2505
R27605 VDD.n7812 VDD.n2246 2.2505
R27606 VDD.n7814 VDD.n7813 2.2505
R27607 VDD.n7815 VDD.n2245 2.2505
R27608 VDD.n7817 VDD.n7816 2.2505
R27609 VDD.n7818 VDD.n2243 2.2505
R27610 VDD.n7820 VDD.n7819 2.2505
R27611 VDD.n2244 VDD.n2242 2.2505
R27612 VDD.n4750 VDD.n4749 2.2505
R27613 VDD.n4751 VDD.n4748 2.2505
R27614 VDD.n4753 VDD.n4752 2.2505
R27615 VDD.n4754 VDD.n4747 2.2505
R27616 VDD.n4756 VDD.n4755 2.2505
R27617 VDD.n4757 VDD.n4746 2.2505
R27618 VDD.n4759 VDD.n4758 2.2505
R27619 VDD.n4760 VDD.n4745 2.2505
R27620 VDD.n4762 VDD.n4761 2.2505
R27621 VDD.n4763 VDD.n4744 2.2505
R27622 VDD.n4765 VDD.n4764 2.2505
R27623 VDD.n4766 VDD.n4743 2.2505
R27624 VDD.n4768 VDD.n4767 2.2505
R27625 VDD.n4769 VDD.n4742 2.2505
R27626 VDD.n4771 VDD.n4770 2.2505
R27627 VDD.n4772 VDD.n4741 2.2505
R27628 VDD.n4774 VDD.n4773 2.2505
R27629 VDD.n4775 VDD.n4740 2.2505
R27630 VDD.n4777 VDD.n4776 2.2505
R27631 VDD.n4778 VDD.n4739 2.2505
R27632 VDD.n4780 VDD.n4779 2.2505
R27633 VDD.n4781 VDD.n4738 2.2505
R27634 VDD.n4783 VDD.n4782 2.2505
R27635 VDD.n4784 VDD.n4737 2.2505
R27636 VDD.n4786 VDD.n4785 2.2505
R27637 VDD.n4787 VDD.n4736 2.2505
R27638 VDD.n4789 VDD.n4788 2.2505
R27639 VDD.n4790 VDD.n4735 2.2505
R27640 VDD.n4792 VDD.n4791 2.2505
R27641 VDD.n4793 VDD.n4734 2.2505
R27642 VDD.n4795 VDD.n4794 2.2505
R27643 VDD.n4796 VDD.n4733 2.2505
R27644 VDD.n4798 VDD.n4797 2.2505
R27645 VDD.n4799 VDD.n4732 2.2505
R27646 VDD.n4801 VDD.n4800 2.2505
R27647 VDD.n4802 VDD.n4731 2.2505
R27648 VDD.n4804 VDD.n4803 2.2505
R27649 VDD.n4805 VDD.n4730 2.2505
R27650 VDD.n4807 VDD.n4806 2.2505
R27651 VDD.n4808 VDD.n4729 2.2505
R27652 VDD.n4810 VDD.n4809 2.2505
R27653 VDD.n4811 VDD.n4728 2.2505
R27654 VDD.n4813 VDD.n4812 2.2505
R27655 VDD.n4814 VDD.n4727 2.2505
R27656 VDD.n4816 VDD.n4815 2.2505
R27657 VDD.n4817 VDD.n4726 2.2505
R27658 VDD.n4819 VDD.n4818 2.2505
R27659 VDD.n4820 VDD.n4725 2.2505
R27660 VDD.n4822 VDD.n4821 2.2505
R27661 VDD.n4823 VDD.n4724 2.2505
R27662 VDD.n4825 VDD.n4824 2.2505
R27663 VDD.n4826 VDD.n4723 2.2505
R27664 VDD.n4828 VDD.n4827 2.2505
R27665 VDD.n4829 VDD.n4722 2.2505
R27666 VDD.n4831 VDD.n4830 2.2505
R27667 VDD.n4832 VDD.n4721 2.2505
R27668 VDD.n4834 VDD.n4833 2.2505
R27669 VDD.n4835 VDD.n4720 2.2505
R27670 VDD.n4837 VDD.n4836 2.2505
R27671 VDD.n4838 VDD.n4719 2.2505
R27672 VDD.n4840 VDD.n4839 2.2505
R27673 VDD.n4841 VDD.n4718 2.2505
R27674 VDD.n4843 VDD.n4842 2.2505
R27675 VDD.n4844 VDD.n4717 2.2505
R27676 VDD.n4846 VDD.n4845 2.2505
R27677 VDD.n4847 VDD.n4716 2.2505
R27678 VDD.n4849 VDD.n4848 2.2505
R27679 VDD.n4850 VDD.n4715 2.2505
R27680 VDD.n4852 VDD.n4851 2.2505
R27681 VDD.n4853 VDD.n4714 2.2505
R27682 VDD.n4855 VDD.n4854 2.2505
R27683 VDD.n4856 VDD.n4713 2.2505
R27684 VDD.n4858 VDD.n4857 2.2505
R27685 VDD.n4859 VDD.n4712 2.2505
R27686 VDD.n4861 VDD.n4860 2.2505
R27687 VDD.n4862 VDD.n4711 2.2505
R27688 VDD.n4864 VDD.n4863 2.2505
R27689 VDD.n4865 VDD.n4710 2.2505
R27690 VDD.n4867 VDD.n4866 2.2505
R27691 VDD.n4868 VDD.n4709 2.2505
R27692 VDD.n4870 VDD.n4869 2.2505
R27693 VDD.n4871 VDD.n4708 2.2505
R27694 VDD.n4873 VDD.n4872 2.2505
R27695 VDD.n4874 VDD.n4707 2.2505
R27696 VDD.n4876 VDD.n4875 2.2505
R27697 VDD.n4877 VDD.n4706 2.2505
R27698 VDD.n4879 VDD.n4878 2.2505
R27699 VDD.n4880 VDD.n4705 2.2505
R27700 VDD.n4882 VDD.n4881 2.2505
R27701 VDD.n4883 VDD.n4704 2.2505
R27702 VDD.n4885 VDD.n4884 2.2505
R27703 VDD.n4886 VDD.n4703 2.2505
R27704 VDD.n4888 VDD.n4887 2.2505
R27705 VDD.n4889 VDD.n4702 2.2505
R27706 VDD.n4891 VDD.n4890 2.2505
R27707 VDD.n4892 VDD.n4701 2.2505
R27708 VDD.n4894 VDD.n4893 2.2505
R27709 VDD.n4895 VDD.n4700 2.2505
R27710 VDD.n4897 VDD.n4896 2.2505
R27711 VDD.n4898 VDD.n4699 2.2505
R27712 VDD.n4900 VDD.n4899 2.2505
R27713 VDD.n4901 VDD.n4698 2.2505
R27714 VDD.n4903 VDD.n4902 2.2505
R27715 VDD.n4904 VDD.n4697 2.2505
R27716 VDD.n7748 VDD.n2269 2.2505
R27717 VDD.n7747 VDD.n7746 2.2505
R27718 VDD.n7745 VDD.n7744 2.2505
R27719 VDD.n7743 VDD.n2271 2.2505
R27720 VDD.n7742 VDD.n7741 2.2505
R27721 VDD.n7740 VDD.n7739 2.2505
R27722 VDD.n7738 VDD.n2273 2.2505
R27723 VDD.n7737 VDD.n7736 2.2505
R27724 VDD.n7735 VDD.n2274 2.2505
R27725 VDD.n7734 VDD.n7733 2.2505
R27726 VDD.n7732 VDD.n2275 2.2505
R27727 VDD.n7731 VDD.n7730 2.2505
R27728 VDD.n7729 VDD.n2276 2.2505
R27729 VDD.n7728 VDD.n7727 2.2505
R27730 VDD.n7726 VDD.n2277 2.2505
R27731 VDD.n7724 VDD.n7723 2.2505
R27732 VDD.n7722 VDD.n2278 2.2505
R27733 VDD.n7721 VDD.n7720 2.2505
R27734 VDD.n7718 VDD.n2279 2.2505
R27735 VDD.n7717 VDD.n7716 2.2505
R27736 VDD.n7715 VDD.n2280 2.2505
R27737 VDD.n7714 VDD.n7713 2.2505
R27738 VDD.n7712 VDD.n2281 2.2505
R27739 VDD.n7711 VDD.n7710 2.2505
R27740 VDD.n7709 VDD.n7708 2.2505
R27741 VDD.n7707 VDD.n2284 2.2505
R27742 VDD.n7706 VDD.n7705 2.2505
R27743 VDD.n7704 VDD.n2285 2.2505
R27744 VDD.n7703 VDD.n7702 2.2505
R27745 VDD.n7701 VDD.n2286 2.2505
R27746 VDD.n7699 VDD.n7698 2.2505
R27747 VDD.n7697 VDD.n2287 2.2505
R27748 VDD.n7696 VDD.n7695 2.2505
R27749 VDD.n7694 VDD.n2288 2.2505
R27750 VDD.n7693 VDD.n7692 2.2505
R27751 VDD.n7691 VDD.n2289 2.2505
R27752 VDD.n7690 VDD.n7689 2.2505
R27753 VDD.n7688 VDD.n2290 2.2505
R27754 VDD.n7687 VDD.n7686 2.2505
R27755 VDD.n10760 VDD.n8254 2.2505
R27756 VDD.n10759 VDD.n10758 2.2505
R27757 VDD.n10150 VDD.n10149 2.2505
R27758 VDD.n10151 VDD.n8457 2.2505
R27759 VDD.n10153 VDD.n10152 2.2505
R27760 VDD.n10154 VDD.n8456 2.2505
R27761 VDD.n10156 VDD.n10155 2.2505
R27762 VDD.n10157 VDD.n8455 2.2505
R27763 VDD.n10159 VDD.n10158 2.2505
R27764 VDD.n10160 VDD.n8454 2.2505
R27765 VDD.n10162 VDD.n10161 2.2505
R27766 VDD.n10163 VDD.n8453 2.2505
R27767 VDD.n10165 VDD.n10164 2.2505
R27768 VDD.n10166 VDD.n8452 2.2505
R27769 VDD.n10168 VDD.n10167 2.2505
R27770 VDD.n10169 VDD.n8451 2.2505
R27771 VDD.n10171 VDD.n10170 2.2505
R27772 VDD.n10172 VDD.n8450 2.2505
R27773 VDD.n10174 VDD.n10173 2.2505
R27774 VDD.n10175 VDD.n8449 2.2505
R27775 VDD.n10177 VDD.n10176 2.2505
R27776 VDD.n10178 VDD.n8448 2.2505
R27777 VDD.n10180 VDD.n10179 2.2505
R27778 VDD.n10181 VDD.n8447 2.2505
R27779 VDD.n10183 VDD.n10182 2.2505
R27780 VDD.n10184 VDD.n8446 2.2505
R27781 VDD.n10186 VDD.n10185 2.2505
R27782 VDD.n10187 VDD.n8445 2.2505
R27783 VDD.n10189 VDD.n10188 2.2505
R27784 VDD.n10190 VDD.n8444 2.2505
R27785 VDD.n10192 VDD.n10191 2.2505
R27786 VDD.n10193 VDD.n8443 2.2505
R27787 VDD.n10195 VDD.n10194 2.2505
R27788 VDD.n10196 VDD.n8442 2.2505
R27789 VDD.n10198 VDD.n10197 2.2505
R27790 VDD.n10199 VDD.n8441 2.2505
R27791 VDD.n10201 VDD.n10200 2.2505
R27792 VDD.n10202 VDD.n8440 2.2505
R27793 VDD.n10204 VDD.n10203 2.2505
R27794 VDD.n10205 VDD.n8439 2.2505
R27795 VDD.n10207 VDD.n10206 2.2505
R27796 VDD.n10208 VDD.n8438 2.2505
R27797 VDD.n10210 VDD.n10209 2.2505
R27798 VDD.n10211 VDD.n8437 2.2505
R27799 VDD.n10213 VDD.n10212 2.2505
R27800 VDD.n10214 VDD.n8436 2.2505
R27801 VDD.n10216 VDD.n10215 2.2505
R27802 VDD.n10217 VDD.n8435 2.2505
R27803 VDD.n10219 VDD.n10218 2.2505
R27804 VDD.n10220 VDD.n8434 2.2505
R27805 VDD.n10222 VDD.n10221 2.2505
R27806 VDD.n10223 VDD.n8433 2.2505
R27807 VDD.n10225 VDD.n10224 2.2505
R27808 VDD.n10226 VDD.n8432 2.2505
R27809 VDD.n10228 VDD.n10227 2.2505
R27810 VDD.n10229 VDD.n8431 2.2505
R27811 VDD.n10231 VDD.n10230 2.2505
R27812 VDD.n10232 VDD.n8430 2.2505
R27813 VDD.n10234 VDD.n10233 2.2505
R27814 VDD.n10235 VDD.n8429 2.2505
R27815 VDD.n10237 VDD.n10236 2.2505
R27816 VDD.n10238 VDD.n8428 2.2505
R27817 VDD.n10240 VDD.n10239 2.2505
R27818 VDD.n10241 VDD.n8427 2.2505
R27819 VDD.n10243 VDD.n10242 2.2505
R27820 VDD.n10244 VDD.n8426 2.2505
R27821 VDD.n10246 VDD.n10245 2.2505
R27822 VDD.n10247 VDD.n8425 2.2505
R27823 VDD.n10249 VDD.n10248 2.2505
R27824 VDD.n10250 VDD.n8424 2.2505
R27825 VDD.n10252 VDD.n10251 2.2505
R27826 VDD.n10253 VDD.n8423 2.2505
R27827 VDD.n10255 VDD.n10254 2.2505
R27828 VDD.n10256 VDD.n8422 2.2505
R27829 VDD.n10258 VDD.n10257 2.2505
R27830 VDD.n10259 VDD.n8421 2.2505
R27831 VDD.n10261 VDD.n10260 2.2505
R27832 VDD.n10262 VDD.n8420 2.2505
R27833 VDD.n10264 VDD.n10263 2.2505
R27834 VDD.n10265 VDD.n8419 2.2505
R27835 VDD.n10267 VDD.n10266 2.2505
R27836 VDD.n10268 VDD.n8418 2.2505
R27837 VDD.n10270 VDD.n10269 2.2505
R27838 VDD.n10271 VDD.n8417 2.2505
R27839 VDD.n10273 VDD.n10272 2.2505
R27840 VDD.n10274 VDD.n8416 2.2505
R27841 VDD.n10276 VDD.n10275 2.2505
R27842 VDD.n10277 VDD.n8415 2.2505
R27843 VDD.n10279 VDD.n10278 2.2505
R27844 VDD.n10280 VDD.n8414 2.2505
R27845 VDD.n10282 VDD.n10281 2.2505
R27846 VDD.n10283 VDD.n8413 2.2505
R27847 VDD.n10285 VDD.n10284 2.2505
R27848 VDD.n10286 VDD.n8412 2.2505
R27849 VDD.n10288 VDD.n10287 2.2505
R27850 VDD.n10289 VDD.n8411 2.2505
R27851 VDD.n10291 VDD.n10290 2.2505
R27852 VDD.n10292 VDD.n8410 2.2505
R27853 VDD.n10294 VDD.n10293 2.2505
R27854 VDD.n10295 VDD.n8409 2.2505
R27855 VDD.n10297 VDD.n10296 2.2505
R27856 VDD.n10298 VDD.n8408 2.2505
R27857 VDD.n10300 VDD.n10299 2.2505
R27858 VDD.n10301 VDD.n8407 2.2505
R27859 VDD.n10303 VDD.n10302 2.2505
R27860 VDD.n10304 VDD.n8406 2.2505
R27861 VDD.n10306 VDD.n10305 2.2505
R27862 VDD.n10307 VDD.n8405 2.2505
R27863 VDD.n10309 VDD.n10308 2.2505
R27864 VDD.n10310 VDD.n8404 2.2505
R27865 VDD.n10312 VDD.n10311 2.2505
R27866 VDD.n10313 VDD.n8403 2.2505
R27867 VDD.n10315 VDD.n10314 2.2505
R27868 VDD.n10316 VDD.n8402 2.2505
R27869 VDD.n10318 VDD.n10317 2.2505
R27870 VDD.n10319 VDD.n8401 2.2505
R27871 VDD.n10321 VDD.n10320 2.2505
R27872 VDD.n10322 VDD.n8400 2.2505
R27873 VDD.n10324 VDD.n10323 2.2505
R27874 VDD.n10325 VDD.n8399 2.2505
R27875 VDD.n10327 VDD.n10326 2.2505
R27876 VDD.n10328 VDD.n8398 2.2505
R27877 VDD.n10330 VDD.n10329 2.2505
R27878 VDD.n10331 VDD.n8397 2.2505
R27879 VDD.n10333 VDD.n10332 2.2505
R27880 VDD.n10334 VDD.n8396 2.2505
R27881 VDD.n10336 VDD.n10335 2.2505
R27882 VDD.n10337 VDD.n8395 2.2505
R27883 VDD.n10339 VDD.n10338 2.2505
R27884 VDD.n10340 VDD.n8394 2.2505
R27885 VDD.n10342 VDD.n10341 2.2505
R27886 VDD.n10343 VDD.n8393 2.2505
R27887 VDD.n10345 VDD.n10344 2.2505
R27888 VDD.n10346 VDD.n8392 2.2505
R27889 VDD.n10348 VDD.n10347 2.2505
R27890 VDD.n10349 VDD.n8391 2.2505
R27891 VDD.n10351 VDD.n10350 2.2505
R27892 VDD.n10352 VDD.n8390 2.2505
R27893 VDD.n10354 VDD.n10353 2.2505
R27894 VDD.n10355 VDD.n8389 2.2505
R27895 VDD.n10357 VDD.n10356 2.2505
R27896 VDD.n10358 VDD.n8388 2.2505
R27897 VDD.n10360 VDD.n10359 2.2505
R27898 VDD.n10361 VDD.n8387 2.2505
R27899 VDD.n10363 VDD.n10362 2.2505
R27900 VDD.n10364 VDD.n8386 2.2505
R27901 VDD.n10366 VDD.n10365 2.2505
R27902 VDD.n10367 VDD.n8385 2.2505
R27903 VDD.n10369 VDD.n10368 2.2505
R27904 VDD.n10370 VDD.n8384 2.2505
R27905 VDD.n10372 VDD.n10371 2.2505
R27906 VDD.n10373 VDD.n8383 2.2505
R27907 VDD.n10375 VDD.n10374 2.2505
R27908 VDD.n10376 VDD.n8382 2.2505
R27909 VDD.n10378 VDD.n10377 2.2505
R27910 VDD.n10379 VDD.n8381 2.2505
R27911 VDD.n10381 VDD.n10380 2.2505
R27912 VDD.n10382 VDD.n8380 2.2505
R27913 VDD.n10384 VDD.n10383 2.2505
R27914 VDD.n10385 VDD.n8379 2.2505
R27915 VDD.n10387 VDD.n10386 2.2505
R27916 VDD.n10388 VDD.n8378 2.2505
R27917 VDD.n10390 VDD.n10389 2.2505
R27918 VDD.n10391 VDD.n8377 2.2505
R27919 VDD.n10393 VDD.n10392 2.2505
R27920 VDD.n10394 VDD.n8376 2.2505
R27921 VDD.n10396 VDD.n10395 2.2505
R27922 VDD.n10397 VDD.n8375 2.2505
R27923 VDD.n10399 VDD.n10398 2.2505
R27924 VDD.n10400 VDD.n8374 2.2505
R27925 VDD.n10402 VDD.n10401 2.2505
R27926 VDD.n10403 VDD.n8373 2.2505
R27927 VDD.n10405 VDD.n10404 2.2505
R27928 VDD.n10406 VDD.n8372 2.2505
R27929 VDD.n10408 VDD.n10407 2.2505
R27930 VDD.n10409 VDD.n8371 2.2505
R27931 VDD.n10411 VDD.n10410 2.2505
R27932 VDD.n10412 VDD.n8370 2.2505
R27933 VDD.n10414 VDD.n10413 2.2505
R27934 VDD.n10415 VDD.n8369 2.2505
R27935 VDD.n10417 VDD.n10416 2.2505
R27936 VDD.n10418 VDD.n8368 2.2505
R27937 VDD.n10420 VDD.n10419 2.2505
R27938 VDD.n10421 VDD.n8367 2.2505
R27939 VDD.n10423 VDD.n10422 2.2505
R27940 VDD.n10424 VDD.n8366 2.2505
R27941 VDD.n10426 VDD.n10425 2.2505
R27942 VDD.n10427 VDD.n8365 2.2505
R27943 VDD.n10429 VDD.n10428 2.2505
R27944 VDD.n10430 VDD.n8364 2.2505
R27945 VDD.n10432 VDD.n10431 2.2505
R27946 VDD.n10433 VDD.n8363 2.2505
R27947 VDD.n10435 VDD.n10434 2.2505
R27948 VDD.n10436 VDD.n8362 2.2505
R27949 VDD.n10438 VDD.n10437 2.2505
R27950 VDD.n10439 VDD.n8361 2.2505
R27951 VDD.n10441 VDD.n10440 2.2505
R27952 VDD.n10442 VDD.n8360 2.2505
R27953 VDD.n10444 VDD.n10443 2.2505
R27954 VDD.n10445 VDD.n8359 2.2505
R27955 VDD.n10447 VDD.n10446 2.2505
R27956 VDD.n10448 VDD.n8358 2.2505
R27957 VDD.n10450 VDD.n10449 2.2505
R27958 VDD.n10451 VDD.n8357 2.2505
R27959 VDD.n10453 VDD.n10452 2.2505
R27960 VDD.n10454 VDD.n8356 2.2505
R27961 VDD.n10456 VDD.n10455 2.2505
R27962 VDD.n10457 VDD.n8355 2.2505
R27963 VDD.n10459 VDD.n10458 2.2505
R27964 VDD.n10460 VDD.n8354 2.2505
R27965 VDD.n10462 VDD.n10461 2.2505
R27966 VDD.n10463 VDD.n8353 2.2505
R27967 VDD.n10465 VDD.n10464 2.2505
R27968 VDD.n10466 VDD.n8352 2.2505
R27969 VDD.n10468 VDD.n10467 2.2505
R27970 VDD.n10469 VDD.n8351 2.2505
R27971 VDD.n10471 VDD.n10470 2.2505
R27972 VDD.n10472 VDD.n8350 2.2505
R27973 VDD.n10474 VDD.n10473 2.2505
R27974 VDD.n10475 VDD.n8349 2.2505
R27975 VDD.n10477 VDD.n10476 2.2505
R27976 VDD.n10478 VDD.n8348 2.2505
R27977 VDD.n10480 VDD.n10479 2.2505
R27978 VDD.n10481 VDD.n8347 2.2505
R27979 VDD.n10483 VDD.n10482 2.2505
R27980 VDD.n10484 VDD.n8346 2.2505
R27981 VDD.n10486 VDD.n10485 2.2505
R27982 VDD.n10487 VDD.n8345 2.2505
R27983 VDD.n10489 VDD.n10488 2.2505
R27984 VDD.n10490 VDD.n8344 2.2505
R27985 VDD.n10492 VDD.n10491 2.2505
R27986 VDD.n10493 VDD.n8343 2.2505
R27987 VDD.n10495 VDD.n10494 2.2505
R27988 VDD.n10496 VDD.n8342 2.2505
R27989 VDD.n10498 VDD.n10497 2.2505
R27990 VDD.n10499 VDD.n8341 2.2505
R27991 VDD.n10501 VDD.n10500 2.2505
R27992 VDD.n10502 VDD.n8340 2.2505
R27993 VDD.n10504 VDD.n10503 2.2505
R27994 VDD.n10505 VDD.n8339 2.2505
R27995 VDD.n10507 VDD.n10506 2.2505
R27996 VDD.n10508 VDD.n8338 2.2505
R27997 VDD.n10510 VDD.n10509 2.2505
R27998 VDD.n10511 VDD.n8337 2.2505
R27999 VDD.n10513 VDD.n10512 2.2505
R28000 VDD.n10514 VDD.n8336 2.2505
R28001 VDD.n10516 VDD.n10515 2.2505
R28002 VDD.n10517 VDD.n8335 2.2505
R28003 VDD.n10519 VDD.n10518 2.2505
R28004 VDD.n10520 VDD.n8334 2.2505
R28005 VDD.n10522 VDD.n10521 2.2505
R28006 VDD.n10523 VDD.n8333 2.2505
R28007 VDD.n10525 VDD.n10524 2.2505
R28008 VDD.n10526 VDD.n8332 2.2505
R28009 VDD.n10528 VDD.n10527 2.2505
R28010 VDD.n10529 VDD.n8331 2.2505
R28011 VDD.n10531 VDD.n10530 2.2505
R28012 VDD.n10532 VDD.n8330 2.2505
R28013 VDD.n10534 VDD.n10533 2.2505
R28014 VDD.n10535 VDD.n8329 2.2505
R28015 VDD.n10537 VDD.n10536 2.2505
R28016 VDD.n10538 VDD.n8328 2.2505
R28017 VDD.n10540 VDD.n10539 2.2505
R28018 VDD.n10541 VDD.n8327 2.2505
R28019 VDD.n10543 VDD.n10542 2.2505
R28020 VDD.n10544 VDD.n8326 2.2505
R28021 VDD.n10546 VDD.n10545 2.2505
R28022 VDD.n10547 VDD.n8325 2.2505
R28023 VDD.n10549 VDD.n10548 2.2505
R28024 VDD.n10550 VDD.n8324 2.2505
R28025 VDD.n10552 VDD.n10551 2.2505
R28026 VDD.n10553 VDD.n8323 2.2505
R28027 VDD.n10555 VDD.n10554 2.2505
R28028 VDD.n10556 VDD.n8322 2.2505
R28029 VDD.n10558 VDD.n10557 2.2505
R28030 VDD.n10559 VDD.n8321 2.2505
R28031 VDD.n10561 VDD.n10560 2.2505
R28032 VDD.n10562 VDD.n8320 2.2505
R28033 VDD.n10564 VDD.n10563 2.2505
R28034 VDD.n10565 VDD.n8319 2.2505
R28035 VDD.n10567 VDD.n10566 2.2505
R28036 VDD.n10568 VDD.n8318 2.2505
R28037 VDD.n10570 VDD.n10569 2.2505
R28038 VDD.n10571 VDD.n8317 2.2505
R28039 VDD.n10573 VDD.n10572 2.2505
R28040 VDD.n10574 VDD.n8316 2.2505
R28041 VDD.n10576 VDD.n10575 2.2505
R28042 VDD.n10577 VDD.n8315 2.2505
R28043 VDD.n10579 VDD.n10578 2.2505
R28044 VDD.n10580 VDD.n8314 2.2505
R28045 VDD.n10582 VDD.n10581 2.2505
R28046 VDD.n10583 VDD.n8313 2.2505
R28047 VDD.n10585 VDD.n10584 2.2505
R28048 VDD.n10586 VDD.n8312 2.2505
R28049 VDD.n10588 VDD.n10587 2.2505
R28050 VDD.n10589 VDD.n8311 2.2505
R28051 VDD.n10591 VDD.n10590 2.2505
R28052 VDD.n10592 VDD.n8310 2.2505
R28053 VDD.n10594 VDD.n10593 2.2505
R28054 VDD.n10595 VDD.n8309 2.2505
R28055 VDD.n10597 VDD.n10596 2.2505
R28056 VDD.n10598 VDD.n8308 2.2505
R28057 VDD.n10600 VDD.n10599 2.2505
R28058 VDD.n10601 VDD.n8307 2.2505
R28059 VDD.n10603 VDD.n10602 2.2505
R28060 VDD.n10604 VDD.n8306 2.2505
R28061 VDD.n10606 VDD.n10605 2.2505
R28062 VDD.n10607 VDD.n8305 2.2505
R28063 VDD.n10609 VDD.n10608 2.2505
R28064 VDD.n10610 VDD.n8304 2.2505
R28065 VDD.n10612 VDD.n10611 2.2505
R28066 VDD.n10613 VDD.n8303 2.2505
R28067 VDD.n10615 VDD.n10614 2.2505
R28068 VDD.n10616 VDD.n8302 2.2505
R28069 VDD.n10618 VDD.n10617 2.2505
R28070 VDD.n10619 VDD.n8301 2.2505
R28071 VDD.n10621 VDD.n10620 2.2505
R28072 VDD.n10622 VDD.n8300 2.2505
R28073 VDD.n10624 VDD.n10623 2.2505
R28074 VDD.n10625 VDD.n8299 2.2505
R28075 VDD.n10627 VDD.n10626 2.2505
R28076 VDD.n10628 VDD.n8298 2.2505
R28077 VDD.n10630 VDD.n10629 2.2505
R28078 VDD.n10631 VDD.n8297 2.2505
R28079 VDD.n10633 VDD.n10632 2.2505
R28080 VDD.n10634 VDD.n8296 2.2505
R28081 VDD.n10636 VDD.n10635 2.2505
R28082 VDD.n10637 VDD.n8295 2.2505
R28083 VDD.n10639 VDD.n10638 2.2505
R28084 VDD.n10640 VDD.n8294 2.2505
R28085 VDD.n10642 VDD.n10641 2.2505
R28086 VDD.n10643 VDD.n8293 2.2505
R28087 VDD.n10645 VDD.n10644 2.2505
R28088 VDD.n10646 VDD.n8292 2.2505
R28089 VDD.n10648 VDD.n10647 2.2505
R28090 VDD.n10649 VDD.n8291 2.2505
R28091 VDD.n10651 VDD.n10650 2.2505
R28092 VDD.n10652 VDD.n8290 2.2505
R28093 VDD.n10654 VDD.n10653 2.2505
R28094 VDD.n10655 VDD.n8289 2.2505
R28095 VDD.n10657 VDD.n10656 2.2505
R28096 VDD.n10658 VDD.n8288 2.2505
R28097 VDD.n10660 VDD.n10659 2.2505
R28098 VDD.n10661 VDD.n8287 2.2505
R28099 VDD.n10663 VDD.n10662 2.2505
R28100 VDD.n10664 VDD.n8286 2.2505
R28101 VDD.n10666 VDD.n10665 2.2505
R28102 VDD.n10667 VDD.n8285 2.2505
R28103 VDD.n10669 VDD.n10668 2.2505
R28104 VDD.n10670 VDD.n8284 2.2505
R28105 VDD.n10672 VDD.n10671 2.2505
R28106 VDD.n10673 VDD.n8283 2.2505
R28107 VDD.n10675 VDD.n10674 2.2505
R28108 VDD.n10676 VDD.n8282 2.2505
R28109 VDD.n10678 VDD.n10677 2.2505
R28110 VDD.n10679 VDD.n8281 2.2505
R28111 VDD.n10681 VDD.n10680 2.2505
R28112 VDD.n10682 VDD.n8280 2.2505
R28113 VDD.n10684 VDD.n10683 2.2505
R28114 VDD.n10685 VDD.n8279 2.2505
R28115 VDD.n10687 VDD.n10686 2.2505
R28116 VDD.n10688 VDD.n8278 2.2505
R28117 VDD.n10690 VDD.n10689 2.2505
R28118 VDD.n10691 VDD.n8277 2.2505
R28119 VDD.n10693 VDD.n10692 2.2505
R28120 VDD.n10694 VDD.n8276 2.2505
R28121 VDD.n10696 VDD.n10695 2.2505
R28122 VDD.n10697 VDD.n8275 2.2505
R28123 VDD.n10699 VDD.n10698 2.2505
R28124 VDD.n10700 VDD.n8274 2.2505
R28125 VDD.n10702 VDD.n10701 2.2505
R28126 VDD.n10703 VDD.n8273 2.2505
R28127 VDD.n10705 VDD.n10704 2.2505
R28128 VDD.n10706 VDD.n8272 2.2505
R28129 VDD.n10708 VDD.n10707 2.2505
R28130 VDD.n10709 VDD.n8271 2.2505
R28131 VDD.n10711 VDD.n10710 2.2505
R28132 VDD.n10712 VDD.n8270 2.2505
R28133 VDD.n10714 VDD.n10713 2.2505
R28134 VDD.n10715 VDD.n8269 2.2505
R28135 VDD.n10717 VDD.n10716 2.2505
R28136 VDD.n10718 VDD.n8268 2.2505
R28137 VDD.n10720 VDD.n10719 2.2505
R28138 VDD.n10721 VDD.n8267 2.2505
R28139 VDD.n10723 VDD.n10722 2.2505
R28140 VDD.n10724 VDD.n8266 2.2505
R28141 VDD.n10726 VDD.n10725 2.2505
R28142 VDD.n10727 VDD.n8265 2.2505
R28143 VDD.n10729 VDD.n10728 2.2505
R28144 VDD.n10730 VDD.n8264 2.2505
R28145 VDD.n10732 VDD.n10731 2.2505
R28146 VDD.n10733 VDD.n8263 2.2505
R28147 VDD.n10735 VDD.n10734 2.2505
R28148 VDD.n10736 VDD.n8262 2.2505
R28149 VDD.n10738 VDD.n10737 2.2505
R28150 VDD.n10739 VDD.n8261 2.2505
R28151 VDD.n10741 VDD.n10740 2.2505
R28152 VDD.n10742 VDD.n8260 2.2505
R28153 VDD.n10744 VDD.n10743 2.2505
R28154 VDD.n10745 VDD.n8259 2.2505
R28155 VDD.n10747 VDD.n10746 2.2505
R28156 VDD.n10748 VDD.n8258 2.2505
R28157 VDD.n10750 VDD.n10749 2.2505
R28158 VDD.n10751 VDD.n8257 2.2505
R28159 VDD.n10753 VDD.n10752 2.2505
R28160 VDD.n10754 VDD.n8256 2.2505
R28161 VDD.n10756 VDD.n10755 2.2505
R28162 VDD.n10757 VDD.n8255 2.2505
R28163 VDD.n10103 VDD.n9214 2.2505
R28164 VDD.n10105 VDD.n10104 2.2505
R28165 VDD.n10106 VDD.n9213 2.2505
R28166 VDD.n10108 VDD.n10107 2.2505
R28167 VDD.n10109 VDD.n9212 2.2505
R28168 VDD.n10111 VDD.n10110 2.2505
R28169 VDD.n10112 VDD.n9211 2.2505
R28170 VDD.n10114 VDD.n10113 2.2505
R28171 VDD.n10115 VDD.n9210 2.2505
R28172 VDD.n10117 VDD.n10116 2.2505
R28173 VDD.n10118 VDD.n9209 2.2505
R28174 VDD.n10120 VDD.n10119 2.2505
R28175 VDD.n10121 VDD.n9208 2.2505
R28176 VDD.n10123 VDD.n10122 2.2505
R28177 VDD.n10124 VDD.n9207 2.2505
R28178 VDD.n10126 VDD.n10125 2.2505
R28179 VDD.n10127 VDD.n9206 2.2505
R28180 VDD.n10129 VDD.n10128 2.2505
R28181 VDD.n10130 VDD.n9205 2.2505
R28182 VDD.n10132 VDD.n10131 2.2505
R28183 VDD.n10133 VDD.n9204 2.2505
R28184 VDD.n10135 VDD.n10134 2.2505
R28185 VDD.n10136 VDD.n9203 2.2505
R28186 VDD.n10138 VDD.n10137 2.2505
R28187 VDD.n10139 VDD.n9202 2.2505
R28188 VDD.n10141 VDD.n10140 2.2505
R28189 VDD.n10142 VDD.n9201 2.2505
R28190 VDD.n10144 VDD.n10143 2.2505
R28191 VDD.n10145 VDD.n9186 2.2505
R28192 VDD.n10147 VDD.n10146 2.2505
R28193 VDD.n10102 VDD.n10101 2.2505
R28194 VDD.n10100 VDD.n9215 2.2505
R28195 VDD.n10099 VDD.n10098 2.2505
R28196 VDD.n10097 VDD.n9216 2.2505
R28197 VDD.n10096 VDD.n10095 2.2505
R28198 VDD.n10094 VDD.n9217 2.2505
R28199 VDD.n10093 VDD.n10092 2.2505
R28200 VDD.n10091 VDD.n9218 2.2505
R28201 VDD.n10090 VDD.n10089 2.2505
R28202 VDD.n10088 VDD.n9219 2.2505
R28203 VDD.n10087 VDD.n10086 2.2505
R28204 VDD.n10085 VDD.n9220 2.2505
R28205 VDD.n10084 VDD.n10083 2.2505
R28206 VDD.n10082 VDD.n9221 2.2505
R28207 VDD.n10081 VDD.n10080 2.2505
R28208 VDD.n10079 VDD.n9222 2.2505
R28209 VDD.n10078 VDD.n10077 2.2505
R28210 VDD.n10076 VDD.n9223 2.2505
R28211 VDD.n10075 VDD.n10074 2.2505
R28212 VDD.n10073 VDD.n9224 2.2505
R28213 VDD.n10072 VDD.n10071 2.2505
R28214 VDD.n10070 VDD.n9225 2.2505
R28215 VDD.n10069 VDD.n10068 2.2505
R28216 VDD.n10067 VDD.n9226 2.2505
R28217 VDD.n10066 VDD.n10065 2.2505
R28218 VDD.n10064 VDD.n9227 2.2505
R28219 VDD.n10063 VDD.n10062 2.2505
R28220 VDD.n10061 VDD.n9228 2.2505
R28221 VDD.n10060 VDD.n10059 2.2505
R28222 VDD.n10058 VDD.n9229 2.2505
R28223 VDD.n10057 VDD.n10056 2.2505
R28224 VDD.n10055 VDD.n9230 2.2505
R28225 VDD.n10054 VDD.n10053 2.2505
R28226 VDD.n10052 VDD.n9231 2.2505
R28227 VDD.n10051 VDD.n10050 2.2505
R28228 VDD.n10049 VDD.n9232 2.2505
R28229 VDD.n10048 VDD.n10047 2.2505
R28230 VDD.n10046 VDD.n9233 2.2505
R28231 VDD.n10045 VDD.n10044 2.2505
R28232 VDD.n10043 VDD.n9234 2.2505
R28233 VDD.n10042 VDD.n10041 2.2505
R28234 VDD.n10040 VDD.n9235 2.2505
R28235 VDD.n10039 VDD.n10038 2.2505
R28236 VDD.n10037 VDD.n9236 2.2505
R28237 VDD.n10036 VDD.n10035 2.2505
R28238 VDD.n10034 VDD.n9237 2.2505
R28239 VDD.n10033 VDD.n10032 2.2505
R28240 VDD.n10031 VDD.n9238 2.2505
R28241 VDD.n10030 VDD.n10029 2.2505
R28242 VDD.n10028 VDD.n9239 2.2505
R28243 VDD.n10027 VDD.n10026 2.2505
R28244 VDD.n10025 VDD.n9240 2.2505
R28245 VDD.n10024 VDD.n10023 2.2505
R28246 VDD.n10022 VDD.n9241 2.2505
R28247 VDD.n10021 VDD.n10020 2.2505
R28248 VDD.n10019 VDD.n9242 2.2505
R28249 VDD.n10018 VDD.n10017 2.2505
R28250 VDD.n10016 VDD.n9243 2.2505
R28251 VDD.n10015 VDD.n10014 2.2505
R28252 VDD.n10013 VDD.n9244 2.2505
R28253 VDD.n10012 VDD.n10011 2.2505
R28254 VDD.n10010 VDD.n9245 2.2505
R28255 VDD.n10009 VDD.n10008 2.2505
R28256 VDD.n10007 VDD.n9246 2.2505
R28257 VDD.n10006 VDD.n10005 2.2505
R28258 VDD.n10004 VDD.n9247 2.2505
R28259 VDD.n10003 VDD.n10002 2.2505
R28260 VDD.n10001 VDD.n9248 2.2505
R28261 VDD.n10000 VDD.n9999 2.2505
R28262 VDD.n9998 VDD.n9249 2.2505
R28263 VDD.n9997 VDD.n9996 2.2505
R28264 VDD.n9995 VDD.n9250 2.2505
R28265 VDD.n9994 VDD.n9993 2.2505
R28266 VDD.n9992 VDD.n9251 2.2505
R28267 VDD.n9991 VDD.n9990 2.2505
R28268 VDD.n9989 VDD.n9252 2.2505
R28269 VDD.n9988 VDD.n9987 2.2505
R28270 VDD.n9986 VDD.n9253 2.2505
R28271 VDD.n9985 VDD.n9984 2.2505
R28272 VDD.n9983 VDD.n9254 2.2505
R28273 VDD.n9982 VDD.n9981 2.2505
R28274 VDD.n9980 VDD.n9255 2.2505
R28275 VDD.n9979 VDD.n9978 2.2505
R28276 VDD.n9977 VDD.n9256 2.2505
R28277 VDD.n9976 VDD.n9975 2.2505
R28278 VDD.n9974 VDD.n9257 2.2505
R28279 VDD.n9973 VDD.n9972 2.2505
R28280 VDD.n9971 VDD.n9258 2.2505
R28281 VDD.n9970 VDD.n9969 2.2505
R28282 VDD.n9968 VDD.n9259 2.2505
R28283 VDD.n9967 VDD.n9966 2.2505
R28284 VDD.n9965 VDD.n9260 2.2505
R28285 VDD.n9964 VDD.n9963 2.2505
R28286 VDD.n9962 VDD.n9261 2.2505
R28287 VDD.n9961 VDD.n9960 2.2505
R28288 VDD.n9959 VDD.n9262 2.2505
R28289 VDD.n9958 VDD.n9957 2.2505
R28290 VDD.n9956 VDD.n9263 2.2505
R28291 VDD.n9955 VDD.n9954 2.2505
R28292 VDD.n9953 VDD.n9264 2.2505
R28293 VDD.n9952 VDD.n9951 2.2505
R28294 VDD.n9950 VDD.n9265 2.2505
R28295 VDD.n9949 VDD.n9948 2.2505
R28296 VDD.n9947 VDD.n9266 2.2505
R28297 VDD.n9946 VDD.n9945 2.2505
R28298 VDD.n9944 VDD.n9267 2.2505
R28299 VDD.n9943 VDD.n9942 2.2505
R28300 VDD.n9941 VDD.n9268 2.2505
R28301 VDD.n9940 VDD.n9939 2.2505
R28302 VDD.n9938 VDD.n9269 2.2505
R28303 VDD.n9937 VDD.n9936 2.2505
R28304 VDD.n9935 VDD.n9270 2.2505
R28305 VDD.n9934 VDD.n9933 2.2505
R28306 VDD.n9932 VDD.n9271 2.2505
R28307 VDD.n9931 VDD.n9930 2.2505
R28308 VDD.n9929 VDD.n9272 2.2505
R28309 VDD.n9928 VDD.n9927 2.2505
R28310 VDD.n9926 VDD.n9273 2.2505
R28311 VDD.n9925 VDD.n9924 2.2505
R28312 VDD.n9923 VDD.n9274 2.2505
R28313 VDD.n9922 VDD.n9921 2.2505
R28314 VDD.n9920 VDD.n9275 2.2505
R28315 VDD.n9919 VDD.n9918 2.2505
R28316 VDD.n9917 VDD.n9276 2.2505
R28317 VDD.n9916 VDD.n9915 2.2505
R28318 VDD.n9914 VDD.n9277 2.2505
R28319 VDD.n9913 VDD.n9912 2.2505
R28320 VDD.n9911 VDD.n9278 2.2505
R28321 VDD.n9910 VDD.n9909 2.2505
R28322 VDD.n9908 VDD.n9279 2.2505
R28323 VDD.n9907 VDD.n9906 2.2505
R28324 VDD.n9905 VDD.n9280 2.2505
R28325 VDD.n9904 VDD.n9903 2.2505
R28326 VDD.n9902 VDD.n9281 2.2505
R28327 VDD.n9901 VDD.n9900 2.2505
R28328 VDD.n9899 VDD.n9282 2.2505
R28329 VDD.n9898 VDD.n9897 2.2505
R28330 VDD.n9896 VDD.n9283 2.2505
R28331 VDD.n9895 VDD.n9894 2.2505
R28332 VDD.n9893 VDD.n9284 2.2505
R28333 VDD.n9892 VDD.n9891 2.2505
R28334 VDD.n9890 VDD.n9285 2.2505
R28335 VDD.n9889 VDD.n9888 2.2505
R28336 VDD.n9887 VDD.n9286 2.2505
R28337 VDD.n9886 VDD.n9885 2.2505
R28338 VDD.n9884 VDD.n9287 2.2505
R28339 VDD.n9883 VDD.n9882 2.2505
R28340 VDD.n9881 VDD.n9288 2.2505
R28341 VDD.n9880 VDD.n9879 2.2505
R28342 VDD.n9878 VDD.n9289 2.2505
R28343 VDD.n9877 VDD.n9876 2.2505
R28344 VDD.n9875 VDD.n9290 2.2505
R28345 VDD.n9874 VDD.n9873 2.2505
R28346 VDD.n9872 VDD.n9291 2.2505
R28347 VDD.n9871 VDD.n9870 2.2505
R28348 VDD.n9869 VDD.n9292 2.2505
R28349 VDD.n9868 VDD.n9867 2.2505
R28350 VDD.n9866 VDD.n9293 2.2505
R28351 VDD.n9865 VDD.n9864 2.2505
R28352 VDD.n9863 VDD.n9294 2.2505
R28353 VDD.n9862 VDD.n9861 2.2505
R28354 VDD.n9860 VDD.n9295 2.2505
R28355 VDD.n9859 VDD.n9858 2.2505
R28356 VDD.n9857 VDD.n9296 2.2505
R28357 VDD.n9856 VDD.n9855 2.2505
R28358 VDD.n9854 VDD.n9297 2.2505
R28359 VDD.n9853 VDD.n9852 2.2505
R28360 VDD.n9851 VDD.n9298 2.2505
R28361 VDD.n9850 VDD.n9849 2.2505
R28362 VDD.n9848 VDD.n9299 2.2505
R28363 VDD.n9847 VDD.n9846 2.2505
R28364 VDD.n9845 VDD.n9300 2.2505
R28365 VDD.n9844 VDD.n9843 2.2505
R28366 VDD.n9842 VDD.n9301 2.2505
R28367 VDD.n9841 VDD.n9840 2.2505
R28368 VDD.n9839 VDD.n9302 2.2505
R28369 VDD.n9838 VDD.n9837 2.2505
R28370 VDD.n9836 VDD.n9303 2.2505
R28371 VDD.n9835 VDD.n9834 2.2505
R28372 VDD.n9833 VDD.n9304 2.2505
R28373 VDD.n9832 VDD.n9831 2.2505
R28374 VDD.n9830 VDD.n9305 2.2505
R28375 VDD.n9829 VDD.n9828 2.2505
R28376 VDD.n9827 VDD.n9306 2.2505
R28377 VDD.n9826 VDD.n9825 2.2505
R28378 VDD.n9824 VDD.n9307 2.2505
R28379 VDD.n9823 VDD.n9822 2.2505
R28380 VDD.n9821 VDD.n9308 2.2505
R28381 VDD.n9820 VDD.n9819 2.2505
R28382 VDD.n9818 VDD.n9309 2.2505
R28383 VDD.n9817 VDD.n9816 2.2505
R28384 VDD.n9815 VDD.n9310 2.2505
R28385 VDD.n9814 VDD.n9813 2.2505
R28386 VDD.n9812 VDD.n9311 2.2505
R28387 VDD.n9811 VDD.n9810 2.2505
R28388 VDD.n9809 VDD.n9312 2.2505
R28389 VDD.n9808 VDD.n9807 2.2505
R28390 VDD.n9806 VDD.n9313 2.2505
R28391 VDD.n9805 VDD.n9804 2.2505
R28392 VDD.n9803 VDD.n9314 2.2505
R28393 VDD.n9802 VDD.n9801 2.2505
R28394 VDD.n9800 VDD.n9315 2.2505
R28395 VDD.n9799 VDD.n9798 2.2505
R28396 VDD.n9797 VDD.n9316 2.2505
R28397 VDD.n9796 VDD.n9795 2.2505
R28398 VDD.n9794 VDD.n9317 2.2505
R28399 VDD.n9793 VDD.n9792 2.2505
R28400 VDD.n9791 VDD.n9318 2.2505
R28401 VDD.n9790 VDD.n9789 2.2505
R28402 VDD.n9788 VDD.n9319 2.2505
R28403 VDD.n9787 VDD.n9786 2.2505
R28404 VDD.n9785 VDD.n9320 2.2505
R28405 VDD.n9784 VDD.n9783 2.2505
R28406 VDD.n9782 VDD.n9321 2.2505
R28407 VDD.n9781 VDD.n9780 2.2505
R28408 VDD.n9779 VDD.n9322 2.2505
R28409 VDD.n9778 VDD.n9777 2.2505
R28410 VDD.n9776 VDD.n9323 2.2505
R28411 VDD.n9775 VDD.n9774 2.2505
R28412 VDD.n9773 VDD.n9324 2.2505
R28413 VDD.n9772 VDD.n9771 2.2505
R28414 VDD.n9770 VDD.n9325 2.2505
R28415 VDD.n9769 VDD.n9768 2.2505
R28416 VDD.n9767 VDD.n9326 2.2505
R28417 VDD.n9766 VDD.n9765 2.2505
R28418 VDD.n9764 VDD.n9327 2.2505
R28419 VDD.n9763 VDD.n9762 2.2505
R28420 VDD.n9761 VDD.n9328 2.2505
R28421 VDD.n9760 VDD.n9759 2.2505
R28422 VDD.n9758 VDD.n9329 2.2505
R28423 VDD.n9757 VDD.n9756 2.2505
R28424 VDD.n9755 VDD.n9330 2.2505
R28425 VDD.n9754 VDD.n9753 2.2505
R28426 VDD.n9752 VDD.n9331 2.2505
R28427 VDD.n9751 VDD.n9750 2.2505
R28428 VDD.n9749 VDD.n9332 2.2505
R28429 VDD.n9748 VDD.n9747 2.2505
R28430 VDD.n9746 VDD.n9333 2.2505
R28431 VDD.n9745 VDD.n9744 2.2505
R28432 VDD.n9743 VDD.n9334 2.2505
R28433 VDD.n9742 VDD.n9741 2.2505
R28434 VDD.n9740 VDD.n9335 2.2505
R28435 VDD.n9739 VDD.n9738 2.2505
R28436 VDD.n9737 VDD.n9336 2.2505
R28437 VDD.n9736 VDD.n9735 2.2505
R28438 VDD.n9734 VDD.n9337 2.2505
R28439 VDD.n9733 VDD.n9732 2.2505
R28440 VDD.n9731 VDD.n9338 2.2505
R28441 VDD.n9730 VDD.n9729 2.2505
R28442 VDD.n9728 VDD.n9339 2.2505
R28443 VDD.n9727 VDD.n9726 2.2505
R28444 VDD.n9725 VDD.n9340 2.2505
R28445 VDD.n9724 VDD.n9723 2.2505
R28446 VDD.n9722 VDD.n9341 2.2505
R28447 VDD.n9721 VDD.n9720 2.2505
R28448 VDD.n9719 VDD.n9342 2.2505
R28449 VDD.n9718 VDD.n9717 2.2505
R28450 VDD.n9716 VDD.n9343 2.2505
R28451 VDD.n9715 VDD.n9714 2.2505
R28452 VDD.n9713 VDD.n9344 2.2505
R28453 VDD.n9712 VDD.n9711 2.2505
R28454 VDD.n9710 VDD.n9345 2.2505
R28455 VDD.n9709 VDD.n9708 2.2505
R28456 VDD.n9707 VDD.n9346 2.2505
R28457 VDD.n9706 VDD.n9705 2.2505
R28458 VDD.n9704 VDD.n9347 2.2505
R28459 VDD.n9703 VDD.n9702 2.2505
R28460 VDD.n9701 VDD.n9348 2.2505
R28461 VDD.n9700 VDD.n9699 2.2505
R28462 VDD.n9698 VDD.n9349 2.2505
R28463 VDD.n9697 VDD.n9696 2.2505
R28464 VDD.n9695 VDD.n9350 2.2505
R28465 VDD.n9694 VDD.n9693 2.2505
R28466 VDD.n9692 VDD.n9351 2.2505
R28467 VDD.n9691 VDD.n9690 2.2505
R28468 VDD.n9689 VDD.n9352 2.2505
R28469 VDD.n9688 VDD.n9687 2.2505
R28470 VDD.n9686 VDD.n9353 2.2505
R28471 VDD.n9685 VDD.n9684 2.2505
R28472 VDD.n9683 VDD.n9354 2.2505
R28473 VDD.n9682 VDD.n9681 2.2505
R28474 VDD.n9680 VDD.n9355 2.2505
R28475 VDD.n9679 VDD.n9678 2.2505
R28476 VDD.n9677 VDD.n9356 2.2505
R28477 VDD.n9676 VDD.n9675 2.2505
R28478 VDD.n9674 VDD.n9357 2.2505
R28479 VDD.n9673 VDD.n9672 2.2505
R28480 VDD.n9671 VDD.n9358 2.2505
R28481 VDD.n9670 VDD.n9669 2.2505
R28482 VDD.n9668 VDD.n9359 2.2505
R28483 VDD.n9667 VDD.n9666 2.2505
R28484 VDD.n9665 VDD.n9360 2.2505
R28485 VDD.n9664 VDD.n9663 2.2505
R28486 VDD.n9662 VDD.n9361 2.2505
R28487 VDD.n9661 VDD.n9660 2.2505
R28488 VDD.n9659 VDD.n9362 2.2505
R28489 VDD.n9658 VDD.n9657 2.2505
R28490 VDD.n9656 VDD.n9363 2.2505
R28491 VDD.n9655 VDD.n9654 2.2505
R28492 VDD.n9653 VDD.n9364 2.2505
R28493 VDD.n9652 VDD.n9651 2.2505
R28494 VDD.n9650 VDD.n9365 2.2505
R28495 VDD.n9649 VDD.n9648 2.2505
R28496 VDD.n9647 VDD.n9366 2.2505
R28497 VDD.n9646 VDD.n9645 2.2505
R28498 VDD.n9644 VDD.n9367 2.2505
R28499 VDD.n9643 VDD.n9642 2.2505
R28500 VDD.n9641 VDD.n9368 2.2505
R28501 VDD.n9640 VDD.n9639 2.2505
R28502 VDD.n9638 VDD.n9369 2.2505
R28503 VDD.n9637 VDD.n9636 2.2505
R28504 VDD.n9635 VDD.n9370 2.2505
R28505 VDD.n9634 VDD.n9633 2.2505
R28506 VDD.n9632 VDD.n9371 2.2505
R28507 VDD.n9631 VDD.n9630 2.2505
R28508 VDD.n9629 VDD.n9372 2.2505
R28509 VDD.n9628 VDD.n9627 2.2505
R28510 VDD.n9626 VDD.n9373 2.2505
R28511 VDD.n9625 VDD.n9624 2.2505
R28512 VDD.n9623 VDD.n9374 2.2505
R28513 VDD.n9622 VDD.n9621 2.2505
R28514 VDD.n9620 VDD.n9375 2.2505
R28515 VDD.n9619 VDD.n9618 2.2505
R28516 VDD.n9617 VDD.n9376 2.2505
R28517 VDD.n9616 VDD.n9615 2.2505
R28518 VDD.n9614 VDD.n9377 2.2505
R28519 VDD.n9613 VDD.n9612 2.2505
R28520 VDD.n9611 VDD.n9378 2.2505
R28521 VDD.n9610 VDD.n9609 2.2505
R28522 VDD.n9608 VDD.n9379 2.2505
R28523 VDD.n9607 VDD.n9606 2.2505
R28524 VDD.n9605 VDD.n9380 2.2505
R28525 VDD.n9604 VDD.n9603 2.2505
R28526 VDD.n9602 VDD.n9381 2.2505
R28527 VDD.n9601 VDD.n9600 2.2505
R28528 VDD.n9599 VDD.n9382 2.2505
R28529 VDD.n9598 VDD.n9597 2.2505
R28530 VDD.n9596 VDD.n9383 2.2505
R28531 VDD.n9595 VDD.n9594 2.2505
R28532 VDD.n9593 VDD.n9384 2.2505
R28533 VDD.n9592 VDD.n9591 2.2505
R28534 VDD.n9590 VDD.n9385 2.2505
R28535 VDD.n9589 VDD.n9588 2.2505
R28536 VDD.n9587 VDD.n9386 2.2505
R28537 VDD.n9586 VDD.n9585 2.2505
R28538 VDD.n9584 VDD.n9387 2.2505
R28539 VDD.n9583 VDD.n9582 2.2505
R28540 VDD.n9581 VDD.n9388 2.2505
R28541 VDD.n9580 VDD.n9579 2.2505
R28542 VDD.n9578 VDD.n9389 2.2505
R28543 VDD.n9577 VDD.n9576 2.2505
R28544 VDD.n9575 VDD.n9390 2.2505
R28545 VDD.n9574 VDD.n9573 2.2505
R28546 VDD.n9572 VDD.n9391 2.2505
R28547 VDD.n9571 VDD.n9570 2.2505
R28548 VDD.n9569 VDD.n9392 2.2505
R28549 VDD.n9568 VDD.n9567 2.2505
R28550 VDD.n9566 VDD.n9393 2.2505
R28551 VDD.n9565 VDD.n9564 2.2505
R28552 VDD.n9563 VDD.n9394 2.2505
R28553 VDD.n9562 VDD.n9561 2.2505
R28554 VDD.n9560 VDD.n9395 2.2505
R28555 VDD.n9559 VDD.n9558 2.2505
R28556 VDD.n9557 VDD.n9396 2.2505
R28557 VDD.n9556 VDD.n9555 2.2505
R28558 VDD.n9554 VDD.n9397 2.2505
R28559 VDD.n9553 VDD.n9552 2.2505
R28560 VDD.n9551 VDD.n9398 2.2505
R28561 VDD.n9550 VDD.n9549 2.2505
R28562 VDD.n9548 VDD.n9399 2.2505
R28563 VDD.n9547 VDD.n9546 2.2505
R28564 VDD.n9545 VDD.n9400 2.2505
R28565 VDD.n9544 VDD.n9543 2.2505
R28566 VDD.n9542 VDD.n9401 2.2505
R28567 VDD.n9541 VDD.n9540 2.2505
R28568 VDD.n9539 VDD.n9402 2.2505
R28569 VDD.n9538 VDD.n9537 2.2505
R28570 VDD.n9536 VDD.n9403 2.2505
R28571 VDD.n9535 VDD.n9534 2.2505
R28572 VDD.n9533 VDD.n9404 2.2505
R28573 VDD.n9532 VDD.n9531 2.2505
R28574 VDD.n9530 VDD.n9405 2.2505
R28575 VDD.n9529 VDD.n9528 2.2505
R28576 VDD.n9527 VDD.n9406 2.2505
R28577 VDD.n9526 VDD.n9525 2.2505
R28578 VDD.n9524 VDD.n9407 2.2505
R28579 VDD.n9523 VDD.n9522 2.2505
R28580 VDD.n9521 VDD.n9408 2.2505
R28581 VDD.n9520 VDD.n9519 2.2505
R28582 VDD.n9518 VDD.n9409 2.2505
R28583 VDD.n9517 VDD.n9516 2.2505
R28584 VDD.n9515 VDD.n9410 2.2505
R28585 VDD.n9514 VDD.n9513 2.2505
R28586 VDD.n9512 VDD.n9411 2.2505
R28587 VDD.n9511 VDD.n9510 2.2505
R28588 VDD.n9509 VDD.n9412 2.2505
R28589 VDD.n9508 VDD.n9507 2.2505
R28590 VDD.n9506 VDD.n9413 2.2505
R28591 VDD.n9505 VDD.n9504 2.2505
R28592 VDD.n9503 VDD.n9414 2.2505
R28593 VDD.n9502 VDD.n9501 2.2505
R28594 VDD.n9500 VDD.n9415 2.2505
R28595 VDD.n9499 VDD.n9498 2.2505
R28596 VDD.n9497 VDD.n9416 2.2505
R28597 VDD.n9496 VDD.n9495 2.2505
R28598 VDD.n9494 VDD.n9417 2.2505
R28599 VDD.n9493 VDD.n9492 2.2505
R28600 VDD.n9491 VDD.n9418 2.2505
R28601 VDD.n9490 VDD.n9489 2.2505
R28602 VDD.n9488 VDD.n9419 2.2505
R28603 VDD.n9487 VDD.n9486 2.2505
R28604 VDD.n9485 VDD.n9420 2.2505
R28605 VDD.n9484 VDD.n9483 2.2505
R28606 VDD.n9482 VDD.n9421 2.2505
R28607 VDD.n9481 VDD.n9480 2.2505
R28608 VDD.n9479 VDD.n9422 2.2505
R28609 VDD.n9478 VDD.n9477 2.2505
R28610 VDD.n9476 VDD.n9423 2.2505
R28611 VDD.n9475 VDD.n9474 2.2505
R28612 VDD.n9473 VDD.n9424 2.2505
R28613 VDD.n9472 VDD.n9471 2.2505
R28614 VDD.n9470 VDD.n9425 2.2505
R28615 VDD.n9469 VDD.n9468 2.2505
R28616 VDD.n9467 VDD.n9426 2.2505
R28617 VDD.n9466 VDD.n9465 2.2505
R28618 VDD.n9464 VDD.n9427 2.2505
R28619 VDD.n9463 VDD.n9462 2.2505
R28620 VDD.n9461 VDD.n9428 2.2505
R28621 VDD.n9460 VDD.n9459 2.2505
R28622 VDD.n9458 VDD.n9429 2.2505
R28623 VDD.n9457 VDD.n9456 2.2505
R28624 VDD.n9455 VDD.n9430 2.2505
R28625 VDD.n9454 VDD.n9453 2.2505
R28626 VDD.n9452 VDD.n9431 2.2505
R28627 VDD.n9451 VDD.n9450 2.2505
R28628 VDD.n9449 VDD.n9432 2.2505
R28629 VDD.n9448 VDD.n9447 2.2505
R28630 VDD.n9446 VDD.n9433 2.2505
R28631 VDD.n9445 VDD.n9444 2.2505
R28632 VDD.n9443 VDD.n9434 2.2505
R28633 VDD.n9442 VDD.n9441 2.2505
R28634 VDD.n9440 VDD.n9435 2.2505
R28635 VDD.n9439 VDD.n9438 2.2505
R28636 VDD.n9437 VDD.n9436 2.2505
R28637 VDD.n12441 VDD.n12440 2.2505
R28638 VDD.n12439 VDD.n196 2.2505
R28639 VDD.n12438 VDD.n12437 2.2505
R28640 VDD.n12436 VDD.n197 2.2505
R28641 VDD.n12435 VDD.n12434 2.2505
R28642 VDD.n12433 VDD.n198 2.2505
R28643 VDD.n12432 VDD.n12431 2.2505
R28644 VDD.n12430 VDD.n199 2.2505
R28645 VDD.n12429 VDD.n12428 2.2505
R28646 VDD.n12427 VDD.n200 2.2505
R28647 VDD.n12426 VDD.n12425 2.2505
R28648 VDD.n12424 VDD.n201 2.2505
R28649 VDD.n12423 VDD.n12422 2.2505
R28650 VDD.n12421 VDD.n202 2.2505
R28651 VDD.n12420 VDD.n12419 2.2505
R28652 VDD.n12418 VDD.n203 2.2505
R28653 VDD.n12417 VDD.n12416 2.2505
R28654 VDD.n12415 VDD.n204 2.2505
R28655 VDD.n12414 VDD.n12413 2.2505
R28656 VDD.n12412 VDD.n205 2.2505
R28657 VDD.n12411 VDD.n12410 2.2505
R28658 VDD.n12409 VDD.n206 2.2505
R28659 VDD.n12408 VDD.n12407 2.2505
R28660 VDD.n12406 VDD.n207 2.2505
R28661 VDD.n12405 VDD.n12404 2.2505
R28662 VDD.n12403 VDD.n208 2.2505
R28663 VDD.n12402 VDD.n12401 2.2505
R28664 VDD.n12400 VDD.n209 2.2505
R28665 VDD.n12399 VDD.n12398 2.2505
R28666 VDD.n12397 VDD.n210 2.2505
R28667 VDD.n12396 VDD.n12395 2.2505
R28668 VDD.n12394 VDD.n211 2.2505
R28669 VDD.n12393 VDD.n12392 2.2505
R28670 VDD.n12391 VDD.n212 2.2505
R28671 VDD.n12390 VDD.n12389 2.2505
R28672 VDD.n12388 VDD.n213 2.2505
R28673 VDD.n12387 VDD.n12386 2.2505
R28674 VDD.n12385 VDD.n214 2.2505
R28675 VDD.n12384 VDD.n12383 2.2505
R28676 VDD.n12382 VDD.n215 2.2505
R28677 VDD.n12381 VDD.n12380 2.2505
R28678 VDD.n12379 VDD.n216 2.2505
R28679 VDD.n12378 VDD.n12377 2.2505
R28680 VDD.n12376 VDD.n217 2.2505
R28681 VDD.n12375 VDD.n12374 2.2505
R28682 VDD.n12373 VDD.n218 2.2505
R28683 VDD.n12372 VDD.n12371 2.2505
R28684 VDD.n12370 VDD.n219 2.2505
R28685 VDD.n12369 VDD.n12368 2.2505
R28686 VDD.n12367 VDD.n220 2.2505
R28687 VDD.n12366 VDD.n12365 2.2505
R28688 VDD.n12364 VDD.n221 2.2505
R28689 VDD.n12363 VDD.n12362 2.2505
R28690 VDD.n12361 VDD.n222 2.2505
R28691 VDD.n12360 VDD.n12359 2.2505
R28692 VDD.n12358 VDD.n223 2.2505
R28693 VDD.n12357 VDD.n12356 2.2505
R28694 VDD.n12355 VDD.n224 2.2505
R28695 VDD.n12354 VDD.n12353 2.2505
R28696 VDD.n12352 VDD.n225 2.2505
R28697 VDD.n12351 VDD.n12350 2.2505
R28698 VDD.n12349 VDD.n226 2.2505
R28699 VDD.n12348 VDD.n12347 2.2505
R28700 VDD.n12346 VDD.n227 2.2505
R28701 VDD.n12345 VDD.n12344 2.2505
R28702 VDD.n12343 VDD.n228 2.2505
R28703 VDD.n12342 VDD.n12341 2.2505
R28704 VDD.n12340 VDD.n229 2.2505
R28705 VDD.n12339 VDD.n12338 2.2505
R28706 VDD.n12337 VDD.n230 2.2505
R28707 VDD.n12336 VDD.n12335 2.2505
R28708 VDD.n12334 VDD.n231 2.2505
R28709 VDD.n12333 VDD.n12332 2.2505
R28710 VDD.n12331 VDD.n232 2.2505
R28711 VDD.n12330 VDD.n12329 2.2505
R28712 VDD.n12328 VDD.n233 2.2505
R28713 VDD.n12327 VDD.n12326 2.2505
R28714 VDD.n12325 VDD.n234 2.2505
R28715 VDD.n12324 VDD.n12323 2.2505
R28716 VDD.n12322 VDD.n235 2.2505
R28717 VDD.n12321 VDD.n12320 2.2505
R28718 VDD.n12319 VDD.n236 2.2505
R28719 VDD.n12318 VDD.n12317 2.2505
R28720 VDD.n12316 VDD.n237 2.2505
R28721 VDD.n12315 VDD.n12314 2.2505
R28722 VDD.n12313 VDD.n238 2.2505
R28723 VDD.n12312 VDD.n12311 2.2505
R28724 VDD.n12310 VDD.n239 2.2505
R28725 VDD.n12309 VDD.n12308 2.2505
R28726 VDD.n12307 VDD.n240 2.2505
R28727 VDD.n12306 VDD.n12305 2.2505
R28728 VDD.n12304 VDD.n241 2.2505
R28729 VDD.n12303 VDD.n12302 2.2505
R28730 VDD.n12301 VDD.n242 2.2505
R28731 VDD.n12300 VDD.n12299 2.2505
R28732 VDD.n12298 VDD.n243 2.2505
R28733 VDD.n12297 VDD.n12296 2.2505
R28734 VDD.n12295 VDD.n244 2.2505
R28735 VDD.n12294 VDD.n12293 2.2505
R28736 VDD.n12292 VDD.n245 2.2505
R28737 VDD.n12291 VDD.n12290 2.2505
R28738 VDD.n12289 VDD.n246 2.2505
R28739 VDD.n12288 VDD.n12287 2.2505
R28740 VDD.n12286 VDD.n247 2.2505
R28741 VDD.n12285 VDD.n12284 2.2505
R28742 VDD.n12283 VDD.n248 2.2505
R28743 VDD.n12282 VDD.n12281 2.2505
R28744 VDD.n12280 VDD.n249 2.2505
R28745 VDD.n12279 VDD.n12278 2.2505
R28746 VDD.n12277 VDD.n250 2.2505
R28747 VDD.n12276 VDD.n12275 2.2505
R28748 VDD.n12274 VDD.n251 2.2505
R28749 VDD.n12273 VDD.n12272 2.2505
R28750 VDD.n12271 VDD.n252 2.2505
R28751 VDD.n12270 VDD.n12269 2.2505
R28752 VDD.n12268 VDD.n253 2.2505
R28753 VDD.n12267 VDD.n12266 2.2505
R28754 VDD.n12265 VDD.n254 2.2505
R28755 VDD.n12264 VDD.n12263 2.2505
R28756 VDD.n12262 VDD.n255 2.2505
R28757 VDD.n12261 VDD.n12260 2.2505
R28758 VDD.n12259 VDD.n256 2.2505
R28759 VDD.n12258 VDD.n12257 2.2505
R28760 VDD.n12256 VDD.n257 2.2505
R28761 VDD.n12255 VDD.n12254 2.2505
R28762 VDD.n12253 VDD.n258 2.2505
R28763 VDD.n12252 VDD.n12251 2.2505
R28764 VDD.n12250 VDD.n259 2.2505
R28765 VDD.n12249 VDD.n12248 2.2505
R28766 VDD.n12247 VDD.n260 2.2505
R28767 VDD.n12246 VDD.n12245 2.2505
R28768 VDD.n12244 VDD.n261 2.2505
R28769 VDD.n12243 VDD.n12242 2.2505
R28770 VDD.n12241 VDD.n262 2.2505
R28771 VDD.n12240 VDD.n12239 2.2505
R28772 VDD.n12238 VDD.n263 2.2505
R28773 VDD.n12237 VDD.n12236 2.2505
R28774 VDD.n12235 VDD.n264 2.2505
R28775 VDD.n12234 VDD.n12233 2.2505
R28776 VDD.n12232 VDD.n265 2.2505
R28777 VDD.n12231 VDD.n12230 2.2505
R28778 VDD.n12229 VDD.n266 2.2505
R28779 VDD.n12228 VDD.n12227 2.2505
R28780 VDD.n12226 VDD.n267 2.2505
R28781 VDD.n12225 VDD.n12224 2.2505
R28782 VDD.n12223 VDD.n268 2.2505
R28783 VDD.n12222 VDD.n12221 2.2505
R28784 VDD.n12220 VDD.n269 2.2505
R28785 VDD.n12219 VDD.n12218 2.2505
R28786 VDD.n12217 VDD.n270 2.2505
R28787 VDD.n12216 VDD.n12215 2.2505
R28788 VDD.n12214 VDD.n271 2.2505
R28789 VDD.n12213 VDD.n12212 2.2505
R28790 VDD.n12211 VDD.n272 2.2505
R28791 VDD.n12210 VDD.n12209 2.2505
R28792 VDD.n12208 VDD.n273 2.2505
R28793 VDD.n12207 VDD.n12206 2.2505
R28794 VDD.n12205 VDD.n274 2.2505
R28795 VDD.n12204 VDD.n12203 2.2505
R28796 VDD.n12202 VDD.n275 2.2505
R28797 VDD.n12201 VDD.n12200 2.2505
R28798 VDD.n12199 VDD.n276 2.2505
R28799 VDD.n12198 VDD.n12197 2.2505
R28800 VDD.n12196 VDD.n277 2.2505
R28801 VDD.n12195 VDD.n12194 2.2505
R28802 VDD.n12193 VDD.n278 2.2505
R28803 VDD.n12192 VDD.n12191 2.2505
R28804 VDD.n12190 VDD.n279 2.2505
R28805 VDD.n12189 VDD.n12188 2.2505
R28806 VDD.n12187 VDD.n280 2.2505
R28807 VDD.n12186 VDD.n12185 2.2505
R28808 VDD.n12184 VDD.n281 2.2505
R28809 VDD.n12183 VDD.n12182 2.2505
R28810 VDD.n12181 VDD.n282 2.2505
R28811 VDD.n12180 VDD.n12179 2.2505
R28812 VDD.n12178 VDD.n283 2.2505
R28813 VDD.n12177 VDD.n12176 2.2505
R28814 VDD.n12175 VDD.n284 2.2505
R28815 VDD.n12174 VDD.n12173 2.2505
R28816 VDD.n12172 VDD.n285 2.2505
R28817 VDD.n12171 VDD.n12170 2.2505
R28818 VDD.n12169 VDD.n286 2.2505
R28819 VDD.n12168 VDD.n12167 2.2505
R28820 VDD.n12166 VDD.n287 2.2505
R28821 VDD.n12165 VDD.n12164 2.2505
R28822 VDD.n12163 VDD.n288 2.2505
R28823 VDD.n12162 VDD.n12161 2.2505
R28824 VDD.n12160 VDD.n289 2.2505
R28825 VDD.n12159 VDD.n12158 2.2505
R28826 VDD.n12157 VDD.n290 2.2505
R28827 VDD.n12156 VDD.n12155 2.2505
R28828 VDD.n12154 VDD.n291 2.2505
R28829 VDD.n12153 VDD.n12152 2.2505
R28830 VDD.n12151 VDD.n292 2.2505
R28831 VDD.n12150 VDD.n12149 2.2505
R28832 VDD.n12148 VDD.n293 2.2505
R28833 VDD.n12147 VDD.n12146 2.2505
R28834 VDD.n12145 VDD.n294 2.2505
R28835 VDD.n12144 VDD.n12143 2.2505
R28836 VDD.n12142 VDD.n295 2.2505
R28837 VDD.n12141 VDD.n12140 2.2505
R28838 VDD.n12139 VDD.n296 2.2505
R28839 VDD.n12138 VDD.n12137 2.2505
R28840 VDD.n12136 VDD.n297 2.2505
R28841 VDD.n12135 VDD.n12134 2.2505
R28842 VDD.n12133 VDD.n298 2.2505
R28843 VDD.n12132 VDD.n12131 2.2505
R28844 VDD.n12130 VDD.n299 2.2505
R28845 VDD.n12129 VDD.n12128 2.2505
R28846 VDD.n12127 VDD.n300 2.2505
R28847 VDD.n12126 VDD.n12125 2.2505
R28848 VDD.n12124 VDD.n301 2.2505
R28849 VDD.n12123 VDD.n12122 2.2505
R28850 VDD.n12121 VDD.n302 2.2505
R28851 VDD.n12120 VDD.n12119 2.2505
R28852 VDD.n12118 VDD.n303 2.2505
R28853 VDD.n12117 VDD.n12116 2.2505
R28854 VDD.n12115 VDD.n304 2.2505
R28855 VDD.n12114 VDD.n12113 2.2505
R28856 VDD.n12112 VDD.n305 2.2505
R28857 VDD.n12111 VDD.n12110 2.2505
R28858 VDD.n12109 VDD.n306 2.2505
R28859 VDD.n12108 VDD.n12107 2.2505
R28860 VDD.n12106 VDD.n307 2.2505
R28861 VDD.n12105 VDD.n12104 2.2505
R28862 VDD.n12103 VDD.n308 2.2505
R28863 VDD.n12102 VDD.n12101 2.2505
R28864 VDD.n12100 VDD.n309 2.2505
R28865 VDD.n12099 VDD.n12098 2.2505
R28866 VDD.n12097 VDD.n310 2.2505
R28867 VDD.n12096 VDD.n12095 2.2505
R28868 VDD.n12094 VDD.n311 2.2505
R28869 VDD.n12093 VDD.n12092 2.2505
R28870 VDD.n12091 VDD.n312 2.2505
R28871 VDD.n12090 VDD.n12089 2.2505
R28872 VDD.n12088 VDD.n313 2.2505
R28873 VDD.n12087 VDD.n12086 2.2505
R28874 VDD.n12085 VDD.n314 2.2505
R28875 VDD.n12084 VDD.n12083 2.2505
R28876 VDD.n12082 VDD.n315 2.2505
R28877 VDD.n12081 VDD.n12080 2.2505
R28878 VDD.n12079 VDD.n316 2.2505
R28879 VDD.n12078 VDD.n12077 2.2505
R28880 VDD.n12076 VDD.n317 2.2505
R28881 VDD.n12075 VDD.n12074 2.2505
R28882 VDD.n12073 VDD.n318 2.2505
R28883 VDD.n12072 VDD.n12071 2.2505
R28884 VDD.n12070 VDD.n319 2.2505
R28885 VDD.n12069 VDD.n12068 2.2505
R28886 VDD.n12067 VDD.n320 2.2505
R28887 VDD.n12066 VDD.n12065 2.2505
R28888 VDD.n12064 VDD.n321 2.2505
R28889 VDD.n12063 VDD.n12062 2.2505
R28890 VDD.n12061 VDD.n322 2.2505
R28891 VDD.n12060 VDD.n12059 2.2505
R28892 VDD.n12058 VDD.n323 2.2505
R28893 VDD.n12057 VDD.n12056 2.2505
R28894 VDD.n12055 VDD.n324 2.2505
R28895 VDD.n12054 VDD.n12053 2.2505
R28896 VDD.n12052 VDD.n325 2.2505
R28897 VDD.n12051 VDD.n12050 2.2505
R28898 VDD.n12049 VDD.n326 2.2505
R28899 VDD.n12048 VDD.n12047 2.2505
R28900 VDD.n12046 VDD.n327 2.2505
R28901 VDD.n12045 VDD.n12044 2.2505
R28902 VDD.n12043 VDD.n328 2.2505
R28903 VDD.n12042 VDD.n12041 2.2505
R28904 VDD.n12040 VDD.n329 2.2505
R28905 VDD.n12039 VDD.n12038 2.2505
R28906 VDD.n12037 VDD.n330 2.2505
R28907 VDD.n12036 VDD.n12035 2.2505
R28908 VDD.n12034 VDD.n331 2.2505
R28909 VDD.n12033 VDD.n12032 2.2505
R28910 VDD.n12031 VDD.n332 2.2505
R28911 VDD.n12030 VDD.n12029 2.2505
R28912 VDD.n12028 VDD.n333 2.2505
R28913 VDD.n12027 VDD.n12026 2.2505
R28914 VDD.n12025 VDD.n334 2.2505
R28915 VDD.n12024 VDD.n12023 2.2505
R28916 VDD.n12022 VDD.n335 2.2505
R28917 VDD.n12021 VDD.n12020 2.2505
R28918 VDD.n12019 VDD.n336 2.2505
R28919 VDD.n12018 VDD.n12017 2.2505
R28920 VDD.n12016 VDD.n337 2.2505
R28921 VDD.n12015 VDD.n12014 2.2505
R28922 VDD.n12013 VDD.n338 2.2505
R28923 VDD.n12012 VDD.n12011 2.2505
R28924 VDD.n12010 VDD.n339 2.2505
R28925 VDD.n12009 VDD.n12008 2.2505
R28926 VDD.n12007 VDD.n340 2.2505
R28927 VDD.n12006 VDD.n12005 2.2505
R28928 VDD.n12004 VDD.n341 2.2505
R28929 VDD.n12003 VDD.n12002 2.2505
R28930 VDD.n12001 VDD.n342 2.2505
R28931 VDD.n12000 VDD.n11999 2.2505
R28932 VDD.n11998 VDD.n343 2.2505
R28933 VDD.n11997 VDD.n11996 2.2505
R28934 VDD.n11995 VDD.n344 2.2505
R28935 VDD.n11994 VDD.n11993 2.2505
R28936 VDD.n11992 VDD.n345 2.2505
R28937 VDD.n11991 VDD.n11990 2.2505
R28938 VDD.n11989 VDD.n346 2.2505
R28939 VDD.n11988 VDD.n11987 2.2505
R28940 VDD.n11986 VDD.n347 2.2505
R28941 VDD.n11985 VDD.n11984 2.2505
R28942 VDD.n11983 VDD.n348 2.2505
R28943 VDD.n11982 VDD.n11981 2.2505
R28944 VDD.n11980 VDD.n349 2.2505
R28945 VDD.n11979 VDD.n11978 2.2505
R28946 VDD.n11977 VDD.n350 2.2505
R28947 VDD.n11976 VDD.n11975 2.2505
R28948 VDD.n11974 VDD.n351 2.2505
R28949 VDD.n11973 VDD.n11972 2.2505
R28950 VDD.n11971 VDD.n352 2.2505
R28951 VDD.n11970 VDD.n11969 2.2505
R28952 VDD.n11968 VDD.n353 2.2505
R28953 VDD.n11967 VDD.n11966 2.2505
R28954 VDD.n11965 VDD.n354 2.2505
R28955 VDD.n11964 VDD.n11963 2.2505
R28956 VDD.n11962 VDD.n355 2.2505
R28957 VDD.n11961 VDD.n11960 2.2505
R28958 VDD.n11959 VDD.n356 2.2505
R28959 VDD.n11958 VDD.n11957 2.2505
R28960 VDD.n11956 VDD.n357 2.2505
R28961 VDD.n11955 VDD.n11954 2.2505
R28962 VDD.n11953 VDD.n358 2.2505
R28963 VDD.n11952 VDD.n11951 2.2505
R28964 VDD.n11950 VDD.n359 2.2505
R28965 VDD.n11949 VDD.n11948 2.2505
R28966 VDD.n11947 VDD.n360 2.2505
R28967 VDD.n11946 VDD.n11945 2.2505
R28968 VDD.n11944 VDD.n361 2.2505
R28969 VDD.n11943 VDD.n11942 2.2505
R28970 VDD.n11941 VDD.n362 2.2505
R28971 VDD.n11940 VDD.n11939 2.2505
R28972 VDD.n11938 VDD.n363 2.2505
R28973 VDD.n11937 VDD.n11936 2.2505
R28974 VDD.n11935 VDD.n364 2.2505
R28975 VDD.n11934 VDD.n11933 2.2505
R28976 VDD.n11932 VDD.n365 2.2505
R28977 VDD.n11931 VDD.n11930 2.2505
R28978 VDD.n11929 VDD.n366 2.2505
R28979 VDD.n11928 VDD.n11927 2.2505
R28980 VDD.n11926 VDD.n367 2.2505
R28981 VDD.n11925 VDD.n11924 2.2505
R28982 VDD.n11923 VDD.n368 2.2505
R28983 VDD.n11922 VDD.n11921 2.2505
R28984 VDD.n11920 VDD.n369 2.2505
R28985 VDD.n11919 VDD.n11918 2.2505
R28986 VDD.n11917 VDD.n370 2.2505
R28987 VDD.n11916 VDD.n11915 2.2505
R28988 VDD.n11914 VDD.n371 2.2505
R28989 VDD.n11913 VDD.n11912 2.2505
R28990 VDD.n11911 VDD.n372 2.2505
R28991 VDD.n11910 VDD.n11909 2.2505
R28992 VDD.n11908 VDD.n373 2.2505
R28993 VDD.n11907 VDD.n11906 2.2505
R28994 VDD.n11905 VDD.n374 2.2505
R28995 VDD.n11904 VDD.n11903 2.2505
R28996 VDD.n11902 VDD.n375 2.2505
R28997 VDD.n11901 VDD.n11900 2.2505
R28998 VDD.n11899 VDD.n376 2.2505
R28999 VDD.n11898 VDD.n11897 2.2505
R29000 VDD.n11896 VDD.n377 2.2505
R29001 VDD.n11895 VDD.n11894 2.2505
R29002 VDD.n11893 VDD.n378 2.2505
R29003 VDD.n11892 VDD.n11891 2.2505
R29004 VDD.n11890 VDD.n379 2.2505
R29005 VDD.n11889 VDD.n11888 2.2505
R29006 VDD.n11887 VDD.n380 2.2505
R29007 VDD.n11886 VDD.n11885 2.2505
R29008 VDD.n11884 VDD.n381 2.2505
R29009 VDD.n11883 VDD.n11882 2.2505
R29010 VDD.n11881 VDD.n382 2.2505
R29011 VDD.n11880 VDD.n11879 2.2505
R29012 VDD.n11878 VDD.n383 2.2505
R29013 VDD.n11877 VDD.n11876 2.2505
R29014 VDD.n11875 VDD.n384 2.2505
R29015 VDD.n11874 VDD.n11873 2.2505
R29016 VDD.n11871 VDD.n385 2.2505
R29017 VDD.n11870 VDD.n11869 2.2505
R29018 VDD.n11868 VDD.n386 2.2505
R29019 VDD.n11867 VDD.n11866 2.2505
R29020 VDD.n11865 VDD.n387 2.2505
R29021 VDD.n11864 VDD.n11863 2.2505
R29022 VDD.n11862 VDD.n388 2.2505
R29023 VDD.n11861 VDD.n11860 2.2505
R29024 VDD.n11859 VDD.n389 2.2505
R29025 VDD.n11858 VDD.n11857 2.2505
R29026 VDD.n11856 VDD.n390 2.2505
R29027 VDD.n11855 VDD.n11854 2.2505
R29028 VDD.n11853 VDD.n391 2.2505
R29029 VDD.n11852 VDD.n11851 2.2505
R29030 VDD.n11850 VDD.n392 2.2505
R29031 VDD.n11849 VDD.n11848 2.2505
R29032 VDD.n11847 VDD.n393 2.2505
R29033 VDD.n11846 VDD.n11845 2.2505
R29034 VDD.n11844 VDD.n394 2.2505
R29035 VDD.n11843 VDD.n11842 2.2505
R29036 VDD.n11841 VDD.n395 2.2505
R29037 VDD.n11840 VDD.n11839 2.2505
R29038 VDD.n11838 VDD.n396 2.2505
R29039 VDD.n11837 VDD.n11836 2.2505
R29040 VDD.n11835 VDD.n397 2.2505
R29041 VDD.n11834 VDD.n11833 2.2505
R29042 VDD.n11832 VDD.n398 2.2505
R29043 VDD.n11831 VDD.n11830 2.2505
R29044 VDD.n11829 VDD.n399 2.2505
R29045 VDD.n11828 VDD.n11827 2.2505
R29046 VDD.n11826 VDD.n400 2.2505
R29047 VDD.n11825 VDD.n11824 2.2505
R29048 VDD.n11823 VDD.n401 2.2505
R29049 VDD.n11822 VDD.n11821 2.2505
R29050 VDD.n11820 VDD.n402 2.2505
R29051 VDD.n11819 VDD.n11818 2.2505
R29052 VDD.n11817 VDD.n403 2.2505
R29053 VDD.n11816 VDD.n11815 2.2505
R29054 VDD.n11814 VDD.n404 2.2505
R29055 VDD.n11813 VDD.n11812 2.2505
R29056 VDD.n1449 VDD.n1448 2.2505
R29057 VDD.n1754 VDD.n681 2.25019
R29058 VDD.n998 VDD.n957 2.25019
R29059 VDD.n12638 VDD.n2 2.25019
R29060 VDD.n4595 VDD.n2411 2.25018
R29061 VDD.n2118 VDD.n2108 2.25015
R29062 VDD.n5537 VDD.n5490 2.25014
R29063 VDD.n5910 VDD.n5541 2.25014
R29064 VDD.n5889 VDD.n5888 2.25014
R29065 VDD.n6319 VDD.n5913 2.24874
R29066 VDD.n6321 VDD.n6320 2.24218
R29067 VDD.n6323 VDD.n5982 2.24218
R29068 VDD.n6320 VDD.n5915 2.24218
R29069 VDD.n6173 VDD.n6172 2.24218
R29070 VDD.n6177 VDD.n6176 2.24218
R29071 VDD.n6173 VDD.n6017 2.24218
R29072 VDD.n10817 VDD.n10816 2.24218
R29073 VDD.n10818 VDD.n10817 2.24218
R29074 VDD.n8093 VDD.n8092 2.24218
R29075 VDD.n8095 VDD.n2107 2.24218
R29076 VDD.n2117 VDD.n2105 2.24218
R29077 VDD.n2004 VDD.n2003 2.24218
R29078 VDD.n5907 VDD.n5906 2.24218
R29079 VDD.n5534 VDD.n5530 2.24218
R29080 VDD.n5532 VDD.n5529 2.24218
R29081 VDD.n5887 VDD.n1919 2.24218
R29082 VDD.n5882 VDD.n1918 2.24218
R29083 VDD.n5909 VDD.n5901 2.24218
R29084 VDD.n5903 VDD.n5901 2.24218
R29085 VDD.n5884 VDD.n1918 2.24218
R29086 VDD.n5536 VDD.n5503 2.24218
R29087 VDD.n11048 VDD.n671 2.24218
R29088 VDD.n11048 VDD.n670 2.24218
R29089 VDD.n11044 VDD.n672 2.24218
R29090 VDD.n11128 VDD.n11127 2.24218
R29091 VDD.n640 VDD.n639 2.24218
R29092 VDD.n11127 VDD.n643 2.24218
R29093 VDD.n12583 VDD.n12578 2.24218
R29094 VDD.n12585 VDD.n12560 2.24218
R29095 VDD.n12581 VDD.n12562 2.24218
R29096 VDD.n12626 VDD.n10 2.24218
R29097 VDD.n12627 VDD.n12626 2.24218
R29098 VDD.n12622 VDD.n9 2.24218
R29099 VDD.n1753 VDD.n680 2.24218
R29100 VDD.n1758 VDD.n1756 2.24218
R29101 VDD.n1002 VDD.n999 2.24218
R29102 VDD.n1004 VDD.n955 2.24218
R29103 VDD.n4 VDD.n1 2.24218
R29104 VDD.n12637 VDD.n1 2.24218
R29105 VDD.n2424 VDD.n2409 2.24111
R29106 VDD.n5220 VDD.n2423 2.24111
R29107 VDD.n5220 VDD.n2422 2.24111
R29108 VDD.n5220 VDD.n2421 2.24111
R29109 VDD.n5220 VDD.n2420 2.24111
R29110 VDD.n5220 VDD.n2419 2.24111
R29111 VDD.n5220 VDD.n2418 2.24111
R29112 VDD.n5220 VDD.n2417 2.24111
R29113 VDD.n5220 VDD.n2416 2.24111
R29114 VDD.n5220 VDD.n2415 2.24111
R29115 VDD.n5220 VDD.n2414 2.24111
R29116 VDD.n5220 VDD.n2413 2.24111
R29117 VDD.n5220 VDD.n2412 2.24111
R29118 VDD.n4596 VDD.n2408 2.24111
R29119 VDD.n5218 VDD.n5217 2.24111
R29120 VDD.n5218 VDD.n5216 2.24111
R29121 VDD.n5218 VDD.n5215 2.24111
R29122 VDD.n5218 VDD.n5214 2.24111
R29123 VDD.n5218 VDD.n5213 2.24111
R29124 VDD.n5218 VDD.n5212 2.24111
R29125 VDD.n5218 VDD.n5211 2.24111
R29126 VDD.n5218 VDD.n5210 2.24111
R29127 VDD.n5218 VDD.n5209 2.24111
R29128 VDD.n5218 VDD.n5208 2.24111
R29129 VDD.n5218 VDD.n5207 2.24111
R29130 VDD.n5218 VDD.n5206 2.24111
R29131 VDD.n5218 VDD.n5205 2.24111
R29132 VDD.n5203 VDD.n5202 2.24111
R29133 VDD.n5202 VDD.n4597 2.24111
R29134 VDD.n9199 VDD.n9185 2.24111
R29135 VDD.n9198 VDD.n9184 2.24111
R29136 VDD.n9187 VDD.n9185 2.24111
R29137 VDD.n9188 VDD.n9184 2.24111
R29138 VDD.n9189 VDD.n9185 2.24111
R29139 VDD.n9190 VDD.n9184 2.24111
R29140 VDD.n9191 VDD.n9185 2.24111
R29141 VDD.n9192 VDD.n9184 2.24111
R29142 VDD.n9193 VDD.n9185 2.24111
R29143 VDD.n9194 VDD.n9184 2.24111
R29144 VDD.n9195 VDD.n9185 2.24111
R29145 VDD.n9196 VDD.n9184 2.24111
R29146 VDD.n9197 VDD.n9185 2.24111
R29147 VDD.n12448 VDD.n193 2.24111
R29148 VDD.n12448 VDD.n192 2.24111
R29149 VDD.n12448 VDD.n191 2.24111
R29150 VDD.n12445 VDD.n12444 2.24111
R29151 VDD.n12445 VDD.n12443 2.24111
R29152 VDD.n12445 VDD.n12442 2.24111
R29153 VDD.n12446 VDD.n12445 2.24111
R29154 VDD.n6116 VDD.n6115 2.24038
R29155 VDD.n6073 VDD.n6072 2.24038
R29156 VDD.n6800 VDD.n6739 2.24038
R29157 VDD.n6746 VDD.n6745 2.24038
R29158 VDD.n7885 VDD.n7884 2.21344
R29159 VDD.n7881 VDD.n7880 2.21344
R29160 VDD.n7877 VDD.n7876 2.21344
R29161 VDD.n7871 VDD.n7870 2.21344
R29162 VDD.n7867 VDD.n7866 2.21344
R29163 VDD.n6136 VDD.n6135 2.2016
R29164 VDD.n6139 VDD.n6138 2.2016
R29165 VDD.n6143 VDD.n6142 2.2016
R29166 VDD.n6147 VDD.n6146 2.2016
R29167 VDD.n6132 VDD.n6131 2.2016
R29168 VDD.n6128 VDD.n6127 2.2016
R29169 VDD.n6124 VDD.n6123 2.2016
R29170 VDD.n6120 VDD.n6119 2.2016
R29171 VDD.n6044 VDD.n6043 2.2016
R29172 VDD.n6047 VDD.n6046 2.2016
R29173 VDD.n6051 VDD.n6050 2.2016
R29174 VDD.n6055 VDD.n6054 2.2016
R29175 VDD.n6078 VDD.n6077 2.2016
R29176 VDD.n6082 VDD.n6081 2.2016
R29177 VDD.n6086 VDD.n6085 2.2016
R29178 VDD.n6090 VDD.n6089 2.2016
R29179 VDD.n6810 VDD.n6809 2.2016
R29180 VDD.n6813 VDD.n6812 2.2016
R29181 VDD.n6817 VDD.n6816 2.2016
R29182 VDD.n6821 VDD.n6820 2.2016
R29183 VDD.n6826 VDD.n6825 2.2016
R29184 VDD.n6830 VDD.n6829 2.2016
R29185 VDD.n6834 VDD.n6833 2.2016
R29186 VDD.n6838 VDD.n6837 2.2016
R29187 VDD.n6777 VDD.n6776 2.2016
R29188 VDD.n6780 VDD.n6779 2.2016
R29189 VDD.n6784 VDD.n6783 2.2016
R29190 VDD.n6788 VDD.n6787 2.2016
R29191 VDD.n6773 VDD.n6772 2.2016
R29192 VDD.n6769 VDD.n6768 2.2016
R29193 VDD.n6765 VDD.n6764 2.2016
R29194 VDD.n6761 VDD.n6760 2.2016
R29195 VDD.n6951 VDD.n6950 2.18645
R29196 VDD.n6504 VDD.n6447 2.18645
R29197 VDD.n6996 VDD.n6995 2.18502
R29198 VDD.n6991 VDD.n6990 2.18502
R29199 VDD.n6986 VDD.n6985 2.18502
R29200 VDD.n6981 VDD.n6980 2.18502
R29201 VDD.n6899 VDD.n6898 2.18502
R29202 VDD.n6894 VDD.n6893 2.18502
R29203 VDD.n6889 VDD.n6888 2.18502
R29204 VDD.n6948 VDD.n6947 2.18502
R29205 VDD.n6943 VDD.n6942 2.18502
R29206 VDD.n6938 VDD.n6937 2.18502
R29207 VDD.n6933 VDD.n6932 2.18502
R29208 VDD.n6918 VDD.n6917 2.18502
R29209 VDD.n6913 VDD.n6912 2.18502
R29210 VDD.n6908 VDD.n6907 2.18502
R29211 VDD.n6446 VDD.n6445 2.18502
R29212 VDD.n6443 VDD.n6442 2.18502
R29213 VDD.n6440 VDD.n6439 2.18502
R29214 VDD.n6437 VDD.n6436 2.18502
R29215 VDD.n6432 VDD.n6431 2.18502
R29216 VDD.n6427 VDD.n6426 2.18502
R29217 VDD.n6422 VDD.n6421 2.18502
R29218 VDD.n6483 VDD.n6482 2.18502
R29219 VDD.n6480 VDD.n6479 2.18502
R29220 VDD.n6477 VDD.n6476 2.18502
R29221 VDD.n6474 VDD.n6473 2.18502
R29222 VDD.n6469 VDD.n6468 2.18502
R29223 VDD.n6464 VDD.n6463 2.18502
R29224 VDD.n6459 VDD.n6458 2.18502
R29225 VDD.n8044 VDD.n8043 2.1566
R29226 VDD.n8039 VDD.n8038 2.1566
R29227 VDD.n8034 VDD.n8033 2.1566
R29228 VDD.n8025 VDD.n8024 2.1566
R29229 VDD.n8020 VDD.n8019 2.1566
R29230 VDD.n7939 VDD.n7938 2.14594
R29231 VDD.n7934 VDD.n7933 2.14594
R29232 VDD.n7929 VDD.n7928 2.14594
R29233 VDD.n7920 VDD.n7919 2.14594
R29234 VDD.n7915 VDD.n7914 2.14594
R29235 VDD.n6959 VDD.n6921 2.0852
R29236 VDD.n6496 VDD.n6495 2.0852
R29237 VDD.n6074 VDD.n6073 2.0852
R29238 VDD.n6791 VDD.n6746 2.0852
R29239 VDD.n1761 VDD.n6 1.9774
R29240 VDD.n12634 VDD.n6 1.9617
R29241 VDD.n12634 VDD.n12633 1.84997
R29242 VDD.n1762 VDD.n1761 1.83884
R29243 VDD.n8089 VDD.n8087 1.78866
R29244 VDD.n7015 VDD.n7013 1.73609
R29245 VDD.n6968 VDD.n6878 1.73609
R29246 VDD.n6560 VDD.n6559 1.73609
R29247 VDD.n6521 VDD.n6520 1.73609
R29248 VDD.n2058 VDD.n2057 1.73383
R29249 VDD.n10770 VDD.n10769 1.73383
R29250 VDD.n5260 VDD.n5223 1.73383
R29251 VDD.n5258 VDD.n5224 1.73383
R29252 VDD.n5255 VDD.n5226 1.73383
R29253 VDD.n5250 VDD.n5228 1.73383
R29254 VDD.n5247 VDD.n5229 1.73383
R29255 VDD.n5242 VDD.n5232 1.73383
R29256 VDD.n5240 VDD.n5233 1.73383
R29257 VDD.n5237 VDD.n5235 1.73383
R29258 VDD.n5261 VDD.n5260 1.73383
R29259 VDD.n5258 VDD.n5257 1.73383
R29260 VDD.n5256 VDD.n5255 1.73383
R29261 VDD.n5251 VDD.n5250 1.73383
R29262 VDD.n5247 VDD.n5246 1.73383
R29263 VDD.n5243 VDD.n5242 1.73383
R29264 VDD.n5240 VDD.n5239 1.73383
R29265 VDD.n5238 VDD.n5237 1.73383
R29266 VDD.n5470 VDD.n5380 1.73383
R29267 VDD.n5468 VDD.n5381 1.73383
R29268 VDD.n5465 VDD.n5383 1.73383
R29269 VDD.n5460 VDD.n5385 1.73383
R29270 VDD.n5457 VDD.n5386 1.73383
R29271 VDD.n5452 VDD.n5389 1.73383
R29272 VDD.n5450 VDD.n5390 1.73383
R29273 VDD.n5447 VDD.n5392 1.73383
R29274 VDD.n5471 VDD.n5470 1.73383
R29275 VDD.n5468 VDD.n5467 1.73383
R29276 VDD.n5466 VDD.n5465 1.73383
R29277 VDD.n5461 VDD.n5460 1.73383
R29278 VDD.n5457 VDD.n5456 1.73383
R29279 VDD.n5453 VDD.n5452 1.73383
R29280 VDD.n5450 VDD.n5449 1.73383
R29281 VDD.n5448 VDD.n5447 1.73383
R29282 VDD.n5935 VDD.n5934 1.73383
R29283 VDD.n5932 VDD.n5931 1.73383
R29284 VDD.n5930 VDD.n5929 1.73383
R29285 VDD.n5925 VDD.n5274 1.73383
R29286 VDD.n6582 VDD.n6581 1.73383
R29287 VDD.n6587 VDD.n6586 1.73383
R29288 VDD.n6589 VDD.n6588 1.73383
R29289 VDD.n6592 VDD.n6591 1.73383
R29290 VDD.n5977 VDD.n5976 1.73383
R29291 VDD.n5974 VDD.n5973 1.73383
R29292 VDD.n5972 VDD.n5971 1.73383
R29293 VDD.n5967 VDD.n5966 1.73383
R29294 VDD.n5963 VDD.n5962 1.73383
R29295 VDD.n5959 VDD.n5958 1.73383
R29296 VDD.n5956 VDD.n5955 1.73383
R29297 VDD.n5954 VDD.n5953 1.73383
R29298 VDD.n5359 VDD.n5322 1.73383
R29299 VDD.n5357 VDD.n5323 1.73383
R29300 VDD.n5354 VDD.n5325 1.73383
R29301 VDD.n5349 VDD.n5327 1.73383
R29302 VDD.n5346 VDD.n5328 1.73383
R29303 VDD.n5341 VDD.n5331 1.73383
R29304 VDD.n5339 VDD.n5332 1.73383
R29305 VDD.n5336 VDD.n5334 1.73383
R29306 VDD.n5360 VDD.n5359 1.73383
R29307 VDD.n5357 VDD.n5356 1.73383
R29308 VDD.n5355 VDD.n5354 1.73383
R29309 VDD.n5350 VDD.n5349 1.73383
R29310 VDD.n5346 VDD.n5345 1.73383
R29311 VDD.n5342 VDD.n5341 1.73383
R29312 VDD.n5339 VDD.n5338 1.73383
R29313 VDD.n5337 VDD.n5336 1.73383
R29314 VDD.n6036 VDD.n6035 1.73383
R29315 VDD.n6034 VDD.n6033 1.73383
R29316 VDD.n6031 VDD.n6030 1.73383
R29317 VDD.n6027 VDD.n5283 1.73383
R29318 VDD.n6573 VDD.n6572 1.73383
R29319 VDD.n6569 VDD.n6568 1.73383
R29320 VDD.n6566 VDD.n6565 1.73383
R29321 VDD.n6564 VDD.n6563 1.73383
R29322 VDD.n6170 VDD.n6169 1.73383
R29323 VDD.n6167 VDD.n6166 1.73383
R29324 VDD.n6165 VDD.n6164 1.73383
R29325 VDD.n6160 VDD.n5302 1.73383
R29326 VDD.n6401 VDD.n6400 1.73383
R29327 VDD.n6406 VDD.n6405 1.73383
R29328 VDD.n6408 VDD.n6407 1.73383
R29329 VDD.n6411 VDD.n6410 1.73383
R29330 VDD.n6005 VDD.n5990 1.73383
R29331 VDD.n6003 VDD.n5991 1.73383
R29332 VDD.n6000 VDD.n5993 1.73383
R29333 VDD.n5994 VDD.n5313 1.73383
R29334 VDD.n6392 VDD.n5314 1.73383
R29335 VDD.n6387 VDD.n5317 1.73383
R29336 VDD.n6385 VDD.n5318 1.73383
R29337 VDD.n6382 VDD.n5320 1.73383
R29338 VDD.n6006 VDD.n6005 1.73383
R29339 VDD.n6003 VDD.n6002 1.73383
R29340 VDD.n6001 VDD.n6000 1.73383
R29341 VDD.n5996 VDD.n5313 1.73383
R29342 VDD.n6392 VDD.n6391 1.73383
R29343 VDD.n6388 VDD.n6387 1.73383
R29344 VDD.n6385 VDD.n6384 1.73383
R29345 VDD.n6383 VDD.n6382 1.73383
R29346 VDD.n6294 VDD.n6202 1.73383
R29347 VDD.n6292 VDD.n6203 1.73383
R29348 VDD.n6289 VDD.n6205 1.73383
R29349 VDD.n6284 VDD.n6207 1.73383
R29350 VDD.n6281 VDD.n6208 1.73383
R29351 VDD.n6276 VDD.n6211 1.73383
R29352 VDD.n6274 VDD.n6212 1.73383
R29353 VDD.n6271 VDD.n6214 1.73383
R29354 VDD.n6258 VDD.n6221 1.73383
R29355 VDD.n6256 VDD.n6222 1.73383
R29356 VDD.n6253 VDD.n6224 1.73383
R29357 VDD.n6248 VDD.n6226 1.73383
R29358 VDD.n6245 VDD.n6227 1.73383
R29359 VDD.n6240 VDD.n6230 1.73383
R29360 VDD.n6238 VDD.n6231 1.73383
R29361 VDD.n6235 VDD.n6233 1.73383
R29362 VDD.n6295 VDD.n6294 1.73383
R29363 VDD.n6292 VDD.n6291 1.73383
R29364 VDD.n6290 VDD.n6289 1.73383
R29365 VDD.n6285 VDD.n6284 1.73383
R29366 VDD.n6281 VDD.n6280 1.73383
R29367 VDD.n6277 VDD.n6276 1.73383
R29368 VDD.n6274 VDD.n6273 1.73383
R29369 VDD.n6272 VDD.n6271 1.73383
R29370 VDD.n6259 VDD.n6258 1.73383
R29371 VDD.n6256 VDD.n6255 1.73383
R29372 VDD.n6254 VDD.n6253 1.73383
R29373 VDD.n6249 VDD.n6248 1.73383
R29374 VDD.n6245 VDD.n6244 1.73383
R29375 VDD.n6241 VDD.n6240 1.73383
R29376 VDD.n6238 VDD.n6237 1.73383
R29377 VDD.n6236 VDD.n6235 1.73383
R29378 VDD.n6333 VDD.n6332 1.73383
R29379 VDD.n6337 VDD.n6336 1.73383
R29380 VDD.n6339 VDD.n6338 1.73383
R29381 VDD.n6345 VDD.n6344 1.73383
R29382 VDD.n6347 VDD.n6346 1.73383
R29383 VDD.n6352 VDD.n6351 1.73383
R29384 VDD.n6356 VDD.n6355 1.73383
R29385 VDD.n6358 VDD.n6357 1.73383
R29386 VDD.n6334 VDD.n6333 1.73383
R29387 VDD.n6336 VDD.n6335 1.73383
R29388 VDD.n6340 VDD.n6339 1.73383
R29389 VDD.n6344 VDD.n6343 1.73383
R29390 VDD.n6348 VDD.n6347 1.73383
R29391 VDD.n6353 VDD.n6352 1.73383
R29392 VDD.n6355 VDD.n6354 1.73383
R29393 VDD.n6359 VDD.n6358 1.73383
R29394 VDD.n6622 VDD.n6621 1.73383
R29395 VDD.n6619 VDD.n6618 1.73383
R29396 VDD.n6617 VDD.n6616 1.73383
R29397 VDD.n6612 VDD.n6611 1.73383
R29398 VDD.n6608 VDD.n6607 1.73383
R29399 VDD.n6604 VDD.n6603 1.73383
R29400 VDD.n6601 VDD.n6600 1.73383
R29401 VDD.n7846 VDD.n7845 1.73383
R29402 VDD.n7145 VDD.n7144 1.73383
R29403 VDD.n7149 VDD.n7148 1.73383
R29404 VDD.n7151 VDD.n7150 1.73383
R29405 VDD.n7157 VDD.n7156 1.73383
R29406 VDD.n7159 VDD.n7158 1.73383
R29407 VDD.n7164 VDD.n7163 1.73383
R29408 VDD.n7168 VDD.n7167 1.73383
R29409 VDD.n7170 VDD.n7169 1.73383
R29410 VDD.n7146 VDD.n7145 1.73383
R29411 VDD.n7148 VDD.n7147 1.73383
R29412 VDD.n7152 VDD.n7151 1.73383
R29413 VDD.n7156 VDD.n7155 1.73383
R29414 VDD.n7160 VDD.n7159 1.73383
R29415 VDD.n7165 VDD.n7164 1.73383
R29416 VDD.n7167 VDD.n7166 1.73383
R29417 VDD.n7171 VDD.n7170 1.73383
R29418 VDD.n5431 VDD.n5394 1.73383
R29419 VDD.n5429 VDD.n5395 1.73383
R29420 VDD.n5426 VDD.n5397 1.73383
R29421 VDD.n5421 VDD.n5399 1.73383
R29422 VDD.n5418 VDD.n5400 1.73383
R29423 VDD.n5413 VDD.n5403 1.73383
R29424 VDD.n5411 VDD.n5404 1.73383
R29425 VDD.n5408 VDD.n5406 1.73383
R29426 VDD.n5432 VDD.n5431 1.73383
R29427 VDD.n5429 VDD.n5428 1.73383
R29428 VDD.n5427 VDD.n5426 1.73383
R29429 VDD.n5422 VDD.n5421 1.73383
R29430 VDD.n5418 VDD.n5417 1.73383
R29431 VDD.n5414 VDD.n5413 1.73383
R29432 VDD.n5411 VDD.n5410 1.73383
R29433 VDD.n5409 VDD.n5408 1.73383
R29434 VDD.n8009 VDD.n8008 1.73383
R29435 VDD.n8006 VDD.n8005 1.73383
R29436 VDD.n8004 VDD.n8003 1.73383
R29437 VDD.n7999 VDD.n7998 1.73383
R29438 VDD.n2185 VDD.n2184 1.73383
R29439 VDD.n2181 VDD.n2180 1.73383
R29440 VDD.n2178 VDD.n2177 1.73383
R29441 VDD.n2176 VDD.n2175 1.73383
R29442 VDD.n7971 VDD.n7970 1.73383
R29443 VDD.n7973 VDD.n7972 1.73383
R29444 VDD.n7978 VDD.n7977 1.73383
R29445 VDD.n7984 VDD.n2189 1.73383
R29446 VDD.n7985 VDD.n2192 1.73383
R29447 VDD.n2223 VDD.n2222 1.73383
R29448 VDD.n2231 VDD.n2230 1.73383
R29449 VDD.n2229 VDD.n2228 1.73383
R29450 VDD.n7964 VDD.n7963 1.73383
R29451 VDD.n7982 VDD.n7981 1.73383
R29452 VDD.n7992 VDD.n7991 1.73383
R29453 VDD.n7990 VDD.n7989 1.73383
R29454 VDD.n2225 VDD.n2224 1.73383
R29455 VDD.n2226 VDD.n2212 1.73383
R29456 VDD.n7849 VDD.n7848 1.73383
R29457 VDD.n7847 VDD.n2206 1.73383
R29458 VDD.n6851 VDD.n6850 1.73383
R29459 VDD.n6853 VDD.n6852 1.73383
R29460 VDD.n6856 VDD.n6855 1.73383
R29461 VDD.n6860 VDD.n6859 1.73383
R29462 VDD.n6864 VDD.n6863 1.73383
R29463 VDD.n6869 VDD.n6868 1.73383
R29464 VDD.n6871 VDD.n6870 1.73383
R29465 VDD.n6874 VDD.n6873 1.73383
R29466 VDD.n6726 VDD.n6725 1.73383
R29467 VDD.n6724 VDD.n6723 1.73383
R29468 VDD.n6721 VDD.n6720 1.73383
R29469 VDD.n6717 VDD.n2370 1.73383
R29470 VDD.n7036 VDD.n7035 1.73383
R29471 VDD.n7032 VDD.n7031 1.73383
R29472 VDD.n7029 VDD.n7028 1.73383
R29473 VDD.n7027 VDD.n7026 1.73383
R29474 VDD.n6682 VDD.n6643 1.73383
R29475 VDD.n6680 VDD.n6644 1.73383
R29476 VDD.n6677 VDD.n6646 1.73383
R29477 VDD.n6672 VDD.n6671 1.73383
R29478 VDD.n6670 VDD.n6669 1.73383
R29479 VDD.n6664 VDD.n6651 1.73383
R29480 VDD.n6662 VDD.n6652 1.73383
R29481 VDD.n6659 VDD.n6654 1.73383
R29482 VDD.n7053 VDD.n7052 1.73383
R29483 VDD.n7057 VDD.n7056 1.73383
R29484 VDD.n7059 VDD.n7058 1.73383
R29485 VDD.n7062 VDD.n2333 1.73383
R29486 VDD.n7082 VDD.n2334 1.73383
R29487 VDD.n7077 VDD.n7067 1.73383
R29488 VDD.n7075 VDD.n7068 1.73383
R29489 VDD.n7072 VDD.n7070 1.73383
R29490 VDD.n6683 VDD.n6682 1.73383
R29491 VDD.n6680 VDD.n6679 1.73383
R29492 VDD.n6678 VDD.n6677 1.73383
R29493 VDD.n6673 VDD.n6672 1.73383
R29494 VDD.n6669 VDD.n6668 1.73383
R29495 VDD.n6665 VDD.n6664 1.73383
R29496 VDD.n6662 VDD.n6661 1.73383
R29497 VDD.n6660 VDD.n6659 1.73383
R29498 VDD.n7054 VDD.n7053 1.73383
R29499 VDD.n7056 VDD.n7055 1.73383
R29500 VDD.n7060 VDD.n7059 1.73383
R29501 VDD.n7065 VDD.n2333 1.73383
R29502 VDD.n7082 VDD.n7081 1.73383
R29503 VDD.n7078 VDD.n7077 1.73383
R29504 VDD.n7075 VDD.n7074 1.73383
R29505 VDD.n7073 VDD.n7072 1.73383
R29506 VDD.n7121 VDD.n2325 1.73383
R29507 VDD.n7119 VDD.n2326 1.73383
R29508 VDD.n7116 VDD.n2328 1.73383
R29509 VDD.n7111 VDD.n2330 1.73383
R29510 VDD.n7108 VDD.n7088 1.73383
R29511 VDD.n7103 VDD.n7091 1.73383
R29512 VDD.n7101 VDD.n7092 1.73383
R29513 VDD.n7098 VDD.n7094 1.73383
R29514 VDD.n7122 VDD.n7121 1.73383
R29515 VDD.n7119 VDD.n7118 1.73383
R29516 VDD.n7117 VDD.n7116 1.73383
R29517 VDD.n7112 VDD.n7111 1.73383
R29518 VDD.n7108 VDD.n7107 1.73383
R29519 VDD.n7104 VDD.n7103 1.73383
R29520 VDD.n7101 VDD.n7100 1.73383
R29521 VDD.n7099 VDD.n7098 1.73383
R29522 VDD.n8135 VDD.n8134 1.73383
R29523 VDD.n8163 VDD.n8162 1.73383
R29524 VDD.n8114 VDD.n8113 1.73383
R29525 VDD.n8120 VDD.n8119 1.73383
R29526 VDD.n2046 VDD.n2045 1.73383
R29527 VDD.n2052 VDD.n2051 1.73383
R29528 VDD.n10807 VDD.n10806 1.73383
R29529 VDD.n10801 VDD.n10800 1.73383
R29530 VDD.n8102 VDD.n8101 1.73383
R29531 VDD.n8108 VDD.n8107 1.73383
R29532 VDD.n5583 VDD.n5582 1.73383
R29533 VDD.n5577 VDD.n5576 1.73383
R29534 VDD.n1985 VDD.n1984 1.73383
R29535 VDD.n10813 VDD.n10812 1.73383
R29536 VDD.n1964 VDD.n1963 1.73383
R29537 VDD.n1970 VDD.n1969 1.73383
R29538 VDD.n5604 VDD.n5603 1.73383
R29539 VDD.n5598 VDD.n5597 1.73383
R29540 VDD.n5625 VDD.n5624 1.73383
R29541 VDD.n5619 VDD.n5618 1.73383
R29542 VDD.n10865 VDD.n10864 1.73383
R29543 VDD.n10859 VDD.n10858 1.73383
R29544 VDD.n5508 VDD.n5507 1.73383
R29545 VDD.n10871 VDD.n10870 1.73383
R29546 VDD.n5665 VDD.n5664 1.73383
R29547 VDD.n5659 VDD.n5658 1.73383
R29548 VDD.n5869 VDD.n5868 1.73383
R29549 VDD.n5875 VDD.n5874 1.73383
R29550 VDD.n5520 VDD.n5519 1.73383
R29551 VDD.n5526 VDD.n5525 1.73383
R29552 VDD.n10920 VDD.n10919 1.73383
R29553 VDD.n10914 VDD.n10913 1.73383
R29554 VDD.n5857 VDD.n5856 1.73383
R29555 VDD.n5863 VDD.n5862 1.73383
R29556 VDD.n5814 VDD.n5813 1.73383
R29557 VDD.n5842 VDD.n5841 1.73383
R29558 VDD.n1893 VDD.n1892 1.73383
R29559 VDD.n10926 VDD.n10925 1.73383
R29560 VDD.n1872 VDD.n1871 1.73383
R29561 VDD.n1878 VDD.n1877 1.73383
R29562 VDD.n5802 VDD.n5801 1.73383
R29563 VDD.n5808 VDD.n5807 1.73383
R29564 VDD.n5781 VDD.n5780 1.73383
R29565 VDD.n5787 VDD.n5786 1.73383
R29566 VDD.n10975 VDD.n10974 1.73383
R29567 VDD.n10969 VDD.n10968 1.73383
R29568 VDD.n1828 VDD.n1827 1.73383
R29569 VDD.n10981 VDD.n10980 1.73383
R29570 VDD.n5747 VDD.n5746 1.73383
R29571 VDD.n5775 VDD.n5774 1.73383
R29572 VDD.n5726 VDD.n5725 1.73383
R29573 VDD.n5732 VDD.n5731 1.73383
R29574 VDD.n1816 VDD.n1815 1.73383
R29575 VDD.n1822 VDD.n1821 1.73383
R29576 VDD.n1777 VDD.n1776 1.73383
R29577 VDD.n11024 VDD.n11023 1.73383
R29578 VDD.n11035 VDD.n11034 1.73383
R29579 VDD.n5720 VDD.n5719 1.73383
R29580 VDD.n9072 VDD.n9071 1.73383
R29581 VDD.n9154 VDD.n9153 1.73383
R29582 VDD.n9025 VDD.n9024 1.73383
R29583 VDD.n9030 VDD.n9029 1.73383
R29584 VDD.n8974 VDD.n8973 1.73383
R29585 VDD.n9041 VDD.n9040 1.73383
R29586 VDD.n8950 VDD.n8949 1.73383
R29587 VDD.n9006 VDD.n9005 1.73383
R29588 VDD.n8905 VDD.n8904 1.73383
R29589 VDD.n9019 VDD.n9018 1.73383
R29590 VDD.n8899 VDD.n8898 1.73383
R29591 VDD.n8933 VDD.n8932 1.73383
R29592 VDD.n8847 VDD.n8846 1.73383
R29593 VDD.n8944 VDD.n8943 1.73383
R29594 VDD.n8841 VDD.n8840 1.73383
R29595 VDD.n8875 VDD.n8874 1.73383
R29596 VDD.n8774 VDD.n8773 1.73383
R29597 VDD.n8888 VDD.n8887 1.73383
R29598 VDD.n8768 VDD.n8767 1.73383
R29599 VDD.n8802 VDD.n8801 1.73383
R29600 VDD.n8546 VDD.n8545 1.73383
R29601 VDD.n8835 VDD.n8834 1.73383
R29602 VDD.n8552 VDD.n8551 1.73383
R29603 VDD.n8558 VDD.n8557 1.73383
R29604 VDD.n8756 VDD.n8755 1.73383
R29605 VDD.n8762 VDD.n8761 1.73383
R29606 VDD.n173 VDD.n172 1.73383
R29607 VDD.n189 VDD.n188 1.73383
R29608 VDD.n9094 VDD.n9093 1.73383
R29609 VDD.n9122 VDD.n9121 1.73383
R29610 VDD.n8487 VDD.n8486 1.73383
R29611 VDD.n9165 VDD.n9164 1.73383
R29612 VDD.n9148 VDD.n9147 1.73383
R29613 VDD.n9142 VDD.n9141 1.73383
R29614 VDD.n9132 VDD.n9129 1.73383
R29615 VDD.n9132 VDD.n9131 1.73383
R29616 VDD.n8739 VDD.n8738 1.73383
R29617 VDD.n8745 VDD.n8744 1.73383
R29618 VDD.n8718 VDD.n8717 1.73383
R29619 VDD.n8724 VDD.n8723 1.73383
R29620 VDD.n139 VDD.n138 1.73383
R29621 VDD.n167 VDD.n166 1.73383
R29622 VDD.n12497 VDD.n12496 1.73383
R29623 VDD.n12491 VDD.n12490 1.73383
R29624 VDD.n8706 VDD.n8705 1.73383
R29625 VDD.n8712 VDD.n8711 1.73383
R29626 VDD.n8680 VDD.n8679 1.73383
R29627 VDD.n8686 VDD.n8685 1.73383
R29628 VDD.n93 VDD.n92 1.73383
R29629 VDD.n12503 VDD.n12502 1.73383
R29630 VDD.n50 VDD.n49 1.73383
R29631 VDD.n78 VDD.n77 1.73383
R29632 VDD.n8668 VDD.n8667 1.73383
R29633 VDD.n8674 VDD.n8673 1.73383
R29634 VDD.n8647 VDD.n8646 1.73383
R29635 VDD.n8653 VDD.n8652 1.73383
R29636 VDD.n12553 VDD.n12552 1.73383
R29637 VDD.n12547 VDD.n12546 1.73383
R29638 VDD.n12590 VDD.n12589 1.73383
R29639 VDD.n12597 VDD.n12596 1.73383
R29640 VDD.n12619 VDD.n12618 1.73383
R29641 VDD.n8636 VDD.n8635 1.73383
R29642 VDD.n1562 VDD.n1561 1.73383
R29643 VDD.n1540 VDD.n1539 1.73383
R29644 VDD.n1516 VDD.n1515 1.73383
R29645 VDD.n1527 VDD.n1526 1.73383
R29646 VDD.n1181 VDD.n1180 1.73383
R29647 VDD.n1185 VDD.n1184 1.73383
R29648 VDD.n1168 VDD.n1167 1.73383
R29649 VDD.n1172 VDD.n1171 1.73383
R29650 VDD.n1315 VDD.n1314 1.73383
R29651 VDD.n1656 VDD.n1655 1.73383
R29652 VDD.n1310 VDD.n1309 1.73383
R29653 VDD.n1341 VDD.n1340 1.73383
R29654 VDD.n1361 VDD.n1360 1.73383
R29655 VDD.n1283 VDD.n1082 1.73383
R29656 VDD.n1078 VDD.n1077 1.73383
R29657 VDD.n1388 VDD.n1387 1.73383
R29658 VDD.n1247 VDD.n1246 1.73383
R29659 VDD.n1649 VDD.n1648 1.73383
R29660 VDD.n1602 VDD.n1500 1.73383
R29661 VDD.n1599 VDD.n1501 1.73383
R29662 VDD.n1603 VDD.n1602 1.73383
R29663 VDD.n1599 VDD.n1598 1.73383
R29664 VDD.n1242 VDD.n1241 1.73383
R29665 VDD.n1274 VDD.n1273 1.73383
R29666 VDD.n1211 VDD.n1210 1.73383
R29667 VDD.n1215 VDD.n1214 1.73383
R29668 VDD.n1402 VDD.n1401 1.73383
R29669 VDD.n1411 VDD.n1392 1.73383
R29670 VDD.n1453 VDD.n1452 1.73383
R29671 VDD.n1455 VDD.n1454 1.73383
R29672 VDD.n1488 VDD.n1487 1.73383
R29673 VDD.n1490 VDD.n1489 1.73383
R29674 VDD.n1403 VDD.n1402 1.73383
R29675 VDD.n1411 VDD.n1410 1.73383
R29676 VDD.n1452 VDD.n1451 1.73383
R29677 VDD.n1456 VDD.n1455 1.73383
R29678 VDD.n1487 VDD.n1486 1.73383
R29679 VDD.n1491 VDD.n1490 1.73383
R29680 VDD.n1064 VDD.n1063 1.73383
R29681 VDD.n1068 VDD.n1067 1.73383
R29682 VDD.n909 VDD.n908 1.73383
R29683 VDD.n913 VDD.n912 1.73383
R29684 VDD.n946 VDD.n945 1.73383
R29685 VDD.n1739 VDD.n694 1.73383
R29686 VDD.n947 VDD.n946 1.73383
R29687 VDD.n1739 VDD.n1738 1.73383
R29688 VDD.n724 VDD.n723 1.73383
R29689 VDD.n1715 VDD.n714 1.73383
R29690 VDD.n725 VDD.n724 1.73383
R29691 VDD.n1715 VDD.n1714 1.73383
R29692 VDD.n1747 VDD.n1746 1.73383
R29693 VDD.n1159 VDD.n685 1.73383
R29694 VDD.n1442 VDD.t2746 1.7314
R29695 VDD.n1610 VDD.t2800 1.7314
R29696 VDD.n1610 VDD.t1067 1.7314
R29697 VDD.n1480 VDD.t1530 1.7314
R29698 VDD.n1480 VDD.t4070 1.7314
R29699 VDD.n6157 VDD.n6156 1.69136
R29700 VDD.n6151 VDD.n6037 1.69136
R29701 VDD.n6849 VDD.n6848 1.69136
R29702 VDD.n6841 VDD.n6727 1.69136
R29703 VDD.n6121 VDD.n6019 1.65018
R29704 VDD.n6092 VDD.n6091 1.65018
R29705 VDD.n6840 VDD.n6839 1.65018
R29706 VDD.n6762 VDD.n6758 1.65018
R29707 VDD.n679 VDD.t1169 1.60217
R29708 VDD.n968 VDD.t3581 1.60217
R29709 VDD.n967 VDD.t2545 1.60217
R29710 VDD.n966 VDD.t2668 1.60217
R29711 VDD.n965 VDD.t1431 1.60217
R29712 VDD.n964 VDD.t1560 1.60217
R29713 VDD.n963 VDD.t4610 1.60217
R29714 VDD.n962 VDD.t806 1.60217
R29715 VDD.n961 VDD.t3846 1.60217
R29716 VDD.n960 VDD.t3978 1.60217
R29717 VDD.n959 VDD.t2931 1.60217
R29718 VDD.n958 VDD.t938 1.60217
R29719 VDD.n942 VDD.t684 1.60217
R29720 VDD.n941 VDD.t3330 1.60217
R29721 VDD.n940 VDD.t2224 1.60217
R29722 VDD.n939 VDD.t2622 1.60217
R29723 VDD.n938 VDD.t2498 1.60217
R29724 VDD.n937 VDD.t2628 1.60217
R29725 VDD.n1017 VDD.t1397 1.60217
R29726 VDD.n1018 VDD.t1510 1.60217
R29727 VDD.n1019 VDD.t4544 1.60217
R29728 VDD.n1020 VDD.t2566 1.60217
R29729 VDD.n1021 VDD.t1341 1.60217
R29730 VDD.n12639 VDD.t4000 1.60217
R29731 VDD.n7809 VDD.t3954 1.60217
R29732 VDD.n2252 VDD.t3587 1.60217
R29733 VDD.n2260 VDD.t1079 1.60217
R29734 VDD.n2270 VDD.t1091 1.60217
R29735 VDD.n7725 VDD.t2827 1.60217
R29736 VDD.n2283 VDD.t2452 1.60217
R29737 VDD.n2291 VDD.t2711 1.60217
R29738 VDD.n7826 VDD.t2052 1.60217
R29739 VDD.n7823 VDD.t1663 1.60217
R29740 VDD.n2401 VDD.t2873 1.60217
R29741 VDD.n2399 VDD.t4426 1.60217
R29742 VDD.n2320 VDD.t4092 1.60217
R29743 VDD.n7130 VDD.t992 1.60217
R29744 VDD.n7127 VDD.t4742 1.60217
R29745 VDD.n7125 VDD.t2293 1.60217
R29746 VDD.n2401 VDD.t2526 1.60217
R29747 VDD.n2399 VDD.t4114 1.60217
R29748 VDD.n2320 VDD.t3733 1.60217
R29749 VDD.n7130 VDD.t584 1.60217
R29750 VDD.n7127 VDD.t4396 1.60217
R29751 VDD.n7125 VDD.t1889 1.60217
R29752 VDD.n2323 VDD.t4310 1.60217
R29753 VDD.n2344 VDD.t2017 1.60217
R29754 VDD.n2347 VDD.t1640 1.60217
R29755 VDD.n7044 VDD.t3930 1.60217
R29756 VDD.n7047 VDD.t3562 1.60217
R29757 VDD.n2323 VDD.t3980 1.60217
R29758 VDD.n2344 VDD.t1656 1.60217
R29759 VDD.n2347 VDD.t1284 1.60217
R29760 VDD.n7044 VDD.t3577 1.60217
R29761 VDD.n7047 VDD.t3268 1.60217
R29762 VDD.n6712 VDD.t2871 1.60217
R29763 VDD.n6710 VDD.t4424 1.60217
R29764 VDD.n6707 VDD.t4090 1.60217
R29765 VDD.n6705 VDD.t990 1.60217
R29766 VDD.n6702 VDD.t4740 1.60217
R29767 VDD.n6700 VDD.t2291 1.60217
R29768 VDD.n6712 VDD.t705 1.60217
R29769 VDD.n6710 VDD.t2445 1.60217
R29770 VDD.n6707 VDD.t1999 1.60217
R29771 VDD.n6705 VDD.t3110 1.60217
R29772 VDD.n6702 VDD.t2780 1.60217
R29773 VDD.n6700 VDD.t4330 1.60217
R29774 VDD.n6698 VDD.t4308 1.60217
R29775 VDD.n6696 VDD.t2015 1.60217
R29776 VDD.n6693 VDD.t1638 1.60217
R29777 VDD.n6691 VDD.t3928 1.60217
R29778 VDD.n6688 VDD.t3560 1.60217
R29779 VDD.n6686 VDD.t1059 1.60217
R29780 VDD.n6698 VDD.t2257 1.60217
R29781 VDD.n6696 VDD.t4112 1.60217
R29782 VDD.n6693 VDD.t3731 1.60217
R29783 VDD.n6691 VDD.t1816 1.60217
R29784 VDD.n6688 VDD.t1449 1.60217
R29785 VDD.n6686 VDD.t3188 1.60217
R29786 VDD.n6641 VDD.t1073 1.60217
R29787 VDD.n6639 VDD.t2806 1.60217
R29788 VDD.n6636 VDD.t2435 1.60217
R29789 VDD.n5267 VDD.t2689 1.60217
R29790 VDD.n5436 VDD.t2274 1.60217
R29791 VDD.n5438 VDD.t1953 1.60217
R29792 VDD.n6641 VDD.t3206 1.60217
R29793 VDD.n6639 VDD.t614 1.60217
R29794 VDD.n6636 VDD.t4410 1.60217
R29795 VDD.n5267 VDD.t4678 1.60217
R29796 VDD.n5436 VDD.t4316 1.60217
R29797 VDD.n5438 VDD.t4050 1.60217
R29798 VDD.n5443 VDD.t887 1.60217
R29799 VDD.n5441 VDD.t2604 1.60217
R29800 VDD.n5269 VDD.t2165 1.60217
R29801 VDD.n6630 VDD.t2216 1.60217
R29802 VDD.n6627 VDD.t1806 1.60217
R29803 VDD.n6625 VDD.t3685 1.60217
R29804 VDD.n5443 VDD.t3022 1.60217
R29805 VDD.n5441 VDD.t4558 1.60217
R29806 VDD.n5269 VDD.t4242 1.60217
R29807 VDD.n6630 VDD.t4274 1.60217
R29808 VDD.n6627 VDD.t3920 1.60217
R29809 VDD.n6625 VDD.t1593 1.60217
R29810 VDD.n6265 VDD.t2479 1.60217
R29811 VDD.n5377 VDD.t2048 1.60217
R29812 VDD.n6367 VDD.t2342 1.60217
R29813 VDD.n6364 VDD.t1909 1.60217
R29814 VDD.n6362 VDD.t1622 1.60217
R29815 VDD.n6265 VDD.t3389 1.60217
R29816 VDD.n5377 VDD.t3090 1.60217
R29817 VDD.n6367 VDD.t3304 1.60217
R29818 VDD.n6364 VDD.t3001 1.60217
R29819 VDD.n6362 VDD.t2707 1.60217
R29820 VDD.n5473 VDD.t4690 1.60217
R29821 VDD.n5938 VDD.t2212 1.60217
R29822 VDD.n5941 VDD.t1802 1.60217
R29823 VDD.n5944 VDD.t1855 1.60217
R29824 VDD.n5947 VDD.t1484 1.60217
R29825 VDD.n5949 VDD.t3381 1.60217
R29826 VDD.n5473 VDD.t1499 1.60217
R29827 VDD.n5938 VDD.t3238 1.60217
R29828 VDD.n5941 VDD.t2897 1.60217
R29829 VDD.n5944 VDD.t2951 1.60217
R29830 VDD.n5947 VDD.t2584 1.60217
R29831 VDD.n5949 VDD.t4352 1.60217
R29832 VDD.n6301 VDD.t1007 1.60217
R29833 VDD.n6304 VDD.t587 1.60217
R29834 VDD.n6308 VDD.t896 1.60217
R29835 VDD.n6305 VDD.t4652 1.60217
R29836 VDD.n5984 VDD.t787 1.60217
R29837 VDD.n5987 VDD.t4536 1.60217
R29838 VDD.n6314 VDD.t4594 1.60217
R29839 VDD.n6317 VDD.t4262 1.60217
R29840 VDD.n5979 VDD.t1949 1.60217
R29841 VDD.n6175 VDD.t1065 1.60217
R29842 VDD.n6181 VDD.t2796 1.60217
R29843 VDD.n6184 VDD.t2418 1.60217
R29844 VDD.n6186 VDD.t3405 1.60217
R29845 VDD.n6189 VDD.t3092 1.60217
R29846 VDD.n6191 VDD.t4420 1.60217
R29847 VDD.n6194 VDD.t4086 1.60217
R29848 VDD.n6196 VDD.t2206 1.60217
R29849 VDD.n6199 VDD.t1792 1.60217
R29850 VDD.n5362 VDD.t2557 1.60217
R29851 VDD.n5364 VDD.t4138 1.60217
R29852 VDD.n5367 VDD.t3764 1.60217
R29853 VDD.n5369 VDD.t617 1.60217
R29854 VDD.n5372 VDD.t4422 1.60217
R29855 VDD.n5374 VDD.t1922 1.60217
R29856 VDD.n5362 VDD.t3472 1.60217
R29857 VDD.n5364 VDD.t974 1.60217
R29858 VDD.n5367 VDD.t4734 1.60217
R29859 VDD.n5369 VDD.t1609 1.60217
R29860 VDD.n5372 VDD.t1249 1.60217
R29861 VDD.n5374 VDD.t3009 1.60217
R29862 VDD.n6378 VDD.t4006 1.60217
R29863 VDD.n6376 VDD.t1672 1.60217
R29864 VDD.n6373 VDD.t1306 1.60217
R29865 VDD.n5375 VDD.t3597 1.60217
R29866 VDD.n6218 VDD.t3288 1.60217
R29867 VDD.n6378 VDD.t840 1.60217
R29868 VDD.n6376 VDD.t2772 1.60217
R29869 VDD.n6373 VDD.t2395 1.60217
R29870 VDD.n5375 VDD.t4546 1.60217
R29871 VDD.n6218 VDD.t4238 1.60217
R29872 VDD.n2146 VDD.t1097 1.60217
R29873 VDD.n2157 VDD.t3752 1.60217
R29874 VDD.n2163 VDD.t2169 1.60217
R29875 VDD.n8012 VDD.t911 1.60217
R29876 VDD.n2204 VDD.t1381 1.60217
R29877 VDD.n7863 VDD.t3966 1.60217
R29878 VDD.n7910 VDD.t2305 1.60217
R29879 VDD.n2341 VDD.t2804 1.60217
R29880 VDD.n2360 VDD.t2433 1.60217
R29881 VDD.n2365 VDD.t2687 1.60217
R29882 VDD.n2362 VDD.t2272 1.60217
R29883 VDD.n2311 VDD.t1951 1.60217
R29884 VDD.n2341 VDD.t2450 1.60217
R29885 VDD.n2360 VDD.t2005 1.60217
R29886 VDD.n2365 VDD.t2307 1.60217
R29887 VDD.n2362 VDD.t1880 1.60217
R29888 VDD.n2311 VDD.t1595 1.60217
R29889 VDD.n7141 VDD.t884 1.60217
R29890 VDD.n7139 VDD.t2602 1.60217
R29891 VDD.n7136 VDD.t2163 1.60217
R29892 VDD.n2316 VDD.t2214 1.60217
R29893 VDD.n2313 VDD.t1804 1.60217
R29894 VDD.n7141 VDD.t4664 1.60217
R29895 VDD.n7139 VDD.t2177 1.60217
R29896 VDD.n7136 VDD.t1774 1.60217
R29897 VDD.n2316 VDD.t1827 1.60217
R29898 VDD.n2313 VDD.t1463 1.60217
R29899 VDD.n2296 VDD.t2626 1.60217
R29900 VDD.n2209 VDD.t2192 1.60217
R29901 VDD.n7837 VDD.t2243 1.60217
R29902 VDD.n7840 VDD.t1835 1.60217
R29903 VDD.n7842 VDD.t3711 1.60217
R29904 VDD.n7176 VDD.t2313 1.60217
R29905 VDD.n7946 VDD.t1395 1.60217
R29906 VDD.n7943 VDD.t3986 1.60217
R29907 VDD.n7887 VDD.t2336 1.60217
R29908 VDD.n7888 VDD.t1117 1.60217
R29909 VDD.n8051 VDD.t3780 1.60217
R29910 VDD.n8048 VDD.t2196 1.60217
R29911 VDD.n2172 VDD.t926 1.60217
R29912 VDD.n2390 VDD.t2895 1.60217
R29913 VDD.n2388 VDD.t4458 1.60217
R29914 VDD.n2239 VDD.t4120 1.60217
R29915 VDD.n7831 VDD.t1009 1.60217
R29916 VDD.n7828 VDD.t594 1.60217
R29917 VDD.n1156 VDD.t3607 1.60217
R29918 VDD.n1140 VDD.t4264 1.60217
R29919 VDD.n1141 VDD.t3196 1.60217
R29920 VDD.n1142 VDD.t3302 1.60217
R29921 VDD.n1143 VDD.t2158 1.60217
R29922 VDD.n1144 VDD.t2321 1.60217
R29923 VDD.n705 VDD.t1140 1.60217
R29924 VDD.n704 VDD.t1457 1.60217
R29925 VDD.n703 VDD.t4502 1.60217
R29926 VDD.n702 VDD.t4636 1.60217
R29927 VDD.n701 VDD.t3536 1.60217
R29928 VDD.n1156 VDD.t751 1.60217
R29929 VDD.n1140 VDD.t3914 1.60217
R29930 VDD.n1141 VDD.t2875 1.60217
R29931 VDD.n1142 VDD.t3005 1.60217
R29932 VDD.n1143 VDD.t1772 1.60217
R29933 VDD.n1144 VDD.t1913 1.60217
R29934 VDD.n705 VDD.t816 1.60217
R29935 VDD.n704 VDD.t1130 1.60217
R29936 VDD.n703 VDD.t4192 1.60217
R29937 VDD.n702 VDD.t4294 1.60217
R29938 VDD.n701 VDD.t3244 1.60217
R29939 VDD.n927 VDD.t690 1.60217
R29940 VDD.n926 VDD.t3739 1.60217
R29941 VDD.n925 VDD.t4072 1.60217
R29942 VDD.n924 VDD.t3962 1.60217
R29943 VDD.n923 VDD.t4080 1.60217
R29944 VDD.n922 VDD.t3034 1.60217
R29945 VDD.n921 VDD.t3144 1.60217
R29946 VDD.n920 VDD.t1962 1.60217
R29947 VDD.n919 VDD.t4036 1.60217
R29948 VDD.n918 VDD.t2993 1.60217
R29949 VDD.n917 VDD.t1345 1.60217
R29950 VDD.n927 VDD.t4232 1.60217
R29951 VDD.n926 VDD.t3160 1.60217
R29952 VDD.n925 VDD.t3452 1.60217
R29953 VDD.n924 VDD.t3328 1.60217
R29954 VDD.n923 VDD.t3456 1.60217
R29955 VDD.n922 VDD.t2397 1.60217
R29956 VDD.n921 VDD.t2524 1.60217
R29957 VDD.n920 VDD.t1297 1.60217
R29958 VDD.n919 VDD.t3397 1.60217
R29959 VDD.n918 VDD.t2315 1.60217
R29960 VDD.n917 VDD.t743 1.60217
R29961 VDD.n730 VDD.t2145 1.60217
R29962 VDD.n731 VDD.t1026 1.60217
R29963 VDD.n732 VDD.t1320 1.60217
R29964 VDD.n733 VDD.t1212 1.60217
R29965 VDD.n734 VDD.t1325 1.60217
R29966 VDD.n884 VDD.t4380 1.60217
R29967 VDD.n883 VDD.t4498 1.60217
R29968 VDD.n882 VDD.t3421 1.60217
R29969 VDD.n881 VDD.t1280 1.60217
R29970 VDD.n880 VDD.t4346 1.60217
R29971 VDD.n879 VDD.t2889 1.60217
R29972 VDD.n730 VDD.t1473 1.60217
R29973 VDD.n731 VDD.t4514 1.60217
R29974 VDD.n732 VDD.t710 1.60217
R29975 VDD.n733 VDD.t4736 1.60217
R29976 VDD.n734 VDD.t712 1.60217
R29977 VDD.n884 VDD.t3766 1.60217
R29978 VDD.n883 VDD.t3886 1.60217
R29979 VDD.n882 VDD.t2851 1.60217
R29980 VDD.n881 VDD.t657 1.60217
R29981 VDD.n880 VDD.t3705 1.60217
R29982 VDD.n879 VDD.t2194 1.60217
R29983 VDD.n1462 VDD.t4214 1.60217
R29984 VDD.n1463 VDD.t3148 1.60217
R29985 VDD.n1464 VDD.t3428 1.60217
R29986 VDD.n1465 VDD.t3324 1.60217
R29987 VDD.n1466 VDD.t3436 1.60217
R29988 VDD.n1292 VDD.t2368 1.60217
R29989 VDD.n1291 VDD.t2508 1.60217
R29990 VDD.n1290 VDD.t1278 1.60217
R29991 VDD.n1289 VDD.t3363 1.60217
R29992 VDD.n1288 VDD.t2276 1.60217
R29993 VDD.n1287 VDD.t701 1.60217
R29994 VDD.n1462 VDD.t819 1.60217
R29995 VDD.n1463 VDD.t3856 1.60217
R29996 VDD.n1464 VDD.t4200 1.60217
R29997 VDD.n1465 VDD.t4066 1.60217
R29998 VDD.n1466 VDD.t4208 1.60217
R29999 VDD.n1292 VDD.t3138 1.60217
R30000 VDD.n1291 VDD.t3252 1.60217
R30001 VDD.n1290 VDD.t2091 1.60217
R30002 VDD.n1289 VDD.t4154 1.60217
R30003 VDD.n1288 VDD.t3088 1.60217
R30004 VDD.n1287 VDD.t1455 1.60217
R30005 VDD.n1235 VDD.t1785 1.60217
R30006 VDD.n1220 VDD.t3670 1.60217
R30007 VDD.n1221 VDD.t2648 1.60217
R30008 VDD.n1222 VDD.t2782 1.60217
R30009 VDD.n1223 VDD.t1534 1.60217
R30010 VDD.n1224 VDD.t1668 1.60217
R30011 VDD.n1092 VDD.t4718 1.60217
R30012 VDD.n1093 VDD.t923 1.60217
R30013 VDD.n1094 VDD.t3956 1.60217
R30014 VDD.n1235 VDD.t4204 1.60217
R30015 VDD.n1220 VDD.t2358 1.60217
R30016 VDD.n1221 VDD.t1149 1.60217
R30017 VDD.n1222 VDD.t1268 1.60217
R30018 VDD.n1223 VDD.t4334 1.60217
R30019 VDD.n1224 VDD.t4446 1.60217
R30020 VDD.n1092 VDD.t3344 1.60217
R30021 VDD.n1093 VDD.t3656 1.60217
R30022 VDD.n1094 VDD.t2638 1.60217
R30023 VDD.n1268 VDD.t2905 1.60217
R30024 VDD.n1252 VDD.t662 1.60217
R30025 VDD.n1253 VDD.t3715 1.60217
R30026 VDD.n1254 VDD.t3838 1.60217
R30027 VDD.n1255 VDD.t2810 1.60217
R30028 VDD.n1256 VDD.t2917 1.60217
R30029 VDD.n785 VDD.t1696 1.60217
R30030 VDD.n786 VDD.t2070 1.60217
R30031 VDD.n787 VDD.t958 1.60217
R30032 VDD.n1268 VDD.t1040 1.60217
R30033 VDD.n1252 VDD.t3466 1.60217
R30034 VDD.n1253 VDD.t2404 1.60217
R30035 VDD.n1254 VDD.t2530 1.60217
R30036 VDD.n1255 VDD.t1302 1.60217
R30037 VDD.n1256 VDD.t1427 1.60217
R30038 VDD.n785 VDD.t4476 1.60217
R30039 VDD.n786 VDD.t654 1.60217
R30040 VDD.n787 VDD.t3699 1.60217
R30041 VDD.n1577 VDD.t2462 1.60217
R30042 VDD.n1578 VDD.t1237 1.60217
R30043 VDD.n1579 VDD.t1568 1.60217
R30044 VDD.n1580 VDD.t1445 1.60217
R30045 VDD.n1581 VDD.t1579 1.60217
R30046 VDD.n748 VDD.t4620 1.60217
R30047 VDD.n749 VDD.t4744 1.60217
R30048 VDD.n750 VDD.t3632 1.60217
R30049 VDD.n1505 VDD.t2754 1.60217
R30050 VDD.n1509 VDD.t575 1.60217
R30051 VDD.n1508 VDD.t3642 1.60217
R30052 VDD.n1639 VDD.t4522 1.60217
R30053 VDD.n775 VDD.t4588 1.60217
R30054 VDD.n1519 VDD.t1077 1.60217
R30055 VDD.n780 VDD.t921 1.60217
R30056 VDD.n1566 VDD.t3874 1.60217
R30057 VDD.n769 VDD.t3409 1.60217
R30058 VDD.n773 VDD.t2323 1.60217
R30059 VDD.n776 VDD.t2481 1.60217
R30060 VDD.n778 VDD.t1256 1.60217
R30061 VDD.n781 VDD.t1387 1.60217
R30062 VDD.n1565 VDD.t4428 1.60217
R30063 VDD.n1523 VDD.t3016 1.60217
R30064 VDD.n1522 VDD.t3060 1.60217
R30065 VDD.n1547 VDD.t3603 1.60217
R30066 VDD.n1534 VDD.t3444 1.60217
R30067 VDD.n1535 VDD.t2300 1.60217
R30068 VDD.n1134 VDD.t951 1.60217
R30069 VDD.n1119 VDD.t3626 1.60217
R30070 VDD.n1120 VDD.t2606 1.60217
R30071 VDD.n1121 VDD.t2725 1.60217
R30072 VDD.n1122 VDD.t1497 1.60217
R30073 VDD.n1123 VDD.t1630 1.60217
R30074 VDD.n860 VDD.t4680 1.60217
R30075 VDD.n861 VDD.t879 1.60217
R30076 VDD.n862 VDD.t3904 1.60217
R30077 VDD.n863 VDD.t4038 1.60217
R30078 VDD.n864 VDD.t2997 1.60217
R30079 VDD.n1134 VDD.t2245 1.60217
R30080 VDD.n1119 VDD.t3318 1.60217
R30081 VDD.n1120 VDD.t2187 1.60217
R30082 VDD.n1121 VDD.t2366 1.60217
R30083 VDD.n1122 VDD.t1160 1.60217
R30084 VDD.n1123 VDD.t1274 1.60217
R30085 VDD.n860 VDD.t4338 1.60217
R30086 VDD.n861 VDD.t4658 1.60217
R30087 VDD.n862 VDD.t3554 1.60217
R30088 VDD.n863 VDD.t3666 1.60217
R30089 VDD.n864 VDD.t2646 1.60217
R30090 VDD.n1205 VDD.t4180 1.60217
R30091 VDD.n1190 VDD.t3723 1.60217
R30092 VDD.n1191 VDD.t2697 1.60217
R30093 VDD.n1192 VDD.t2819 1.60217
R30094 VDD.n1193 VDD.t1599 1.60217
R30095 VDD.n1194 VDD.t1717 1.60217
R30096 VDD.n843 VDD.t591 1.60217
R30097 VDD.n842 VDD.t982 1.60217
R30098 VDD.n841 VDD.t4010 1.60217
R30099 VDD.n840 VDD.t4136 1.60217
R30100 VDD.n1205 VDD.t1270 1.60217
R30101 VDD.n1190 VDD.t3387 1.60217
R30102 VDD.n1191 VDD.t2311 1.60217
R30103 VDD.n1192 VDD.t2475 1.60217
R30104 VDD.n1193 VDD.t1254 1.60217
R30105 VDD.n1194 VDD.t1376 1.60217
R30106 VDD.n843 VDD.t4414 1.60217
R30107 VDD.n842 VDD.t558 1.60217
R30108 VDD.n841 VDD.t3634 1.60217
R30109 VDD.n840 VDD.t3774 1.60217
R30110 VDD.n788 VDD.t3968 1.60217
R30111 VDD.n789 VDD.t2915 1.60217
R30112 VDD.n790 VDD.t3226 1.60217
R30113 VDD.n791 VDD.t3116 1.60217
R30114 VDD.n792 VDD.t3232 1.60217
R30115 VDD.n1324 VDD.t2072 1.60217
R30116 VDD.n1323 VDD.t2198 1.60217
R30117 VDD.n1322 VDD.t1069 1.60217
R30118 VDD.n1321 VDD.t3180 1.60217
R30119 VDD.n1320 VDD.t2001 1.60217
R30120 VDD.n1319 VDD.t4608 1.60217
R30121 VDD.n788 VDD.t4716 1.60217
R30122 VDD.n789 VDD.t3618 1.60217
R30123 VDD.n790 VDD.t3952 1.60217
R30124 VDD.n791 VDD.t3822 1.60217
R30125 VDD.n792 VDD.t3960 1.60217
R30126 VDD.n1324 VDD.t2909 1.60217
R30127 VDD.n1323 VDD.t3032 1.60217
R30128 VDD.n1322 VDD.t1812 1.60217
R30129 VDD.n1321 VDD.t3894 1.60217
R30130 VDD.n1320 VDD.t2857 1.60217
R30131 VDD.n1319 VDD.t1221 1.60217
R30132 VDD.n753 VDD.t4552 1.60217
R30133 VDD.n825 VDD.t2473 1.60217
R30134 VDD.n826 VDD.t1247 1.60217
R30135 VDD.n827 VDD.t1583 1.60217
R30136 VDD.n828 VDD.t1453 1.60217
R30137 VDD.n829 VDD.t1587 1.60217
R30138 VDD.n1370 VDD.t4632 1.60217
R30139 VDD.n1369 VDD.t564 1.60217
R30140 VDD.n1368 VDD.t3636 1.60217
R30141 VDD.n1367 VDD.t1524 1.60217
R30142 VDD.n1366 VDD.t4564 1.60217
R30143 VDD.n1365 VDD.t3120 1.60217
R30144 VDD.n825 VDD.t1721 1.60217
R30145 VDD.n826 VDD.t606 1.60217
R30146 VDD.n827 VDD.t988 1.60217
R30147 VDD.n828 VDD.t871 1.60217
R30148 VDD.n829 VDD.t997 1.60217
R30149 VDD.n1370 VDD.t4022 1.60217
R30150 VDD.n1369 VDD.t4146 1.60217
R30151 VDD.n1368 VDD.t3086 1.60217
R30152 VDD.n1367 VDD.t940 1.60217
R30153 VDD.n1366 VDD.t3972 1.60217
R30154 VDD.n1365 VDD.t2512 1.60217
R30155 VDD.n6999 VDD.n6998 1.60175
R30156 VDD.n6523 VDD.n6522 1.60175
R30157 VDD.n72 VDD.n71 1.59478
R30158 VDD.n161 VDD.n160 1.59478
R30159 VDD.n5771 VDD.n5770 1.59478
R30160 VDD.n5838 VDD.n5837 1.59478
R30161 VDD.n5655 VDD.n5654 1.59478
R30162 VDD.n5573 VDD.n5572 1.59478
R30163 VDD.n8159 VDD.n8158 1.59478
R30164 VDD.n9116 VDD.n9115 1.59478
R30165 VDD.n8829 VDD.n8828 1.59478
R30166 VDD.n8969 VDD.n8968 1.59478
R30167 VDD.n751 VDD.t1520 1.58642
R30168 VDD.n1506 VDD.t3784 1.58642
R30169 VDD.n7956 VDD.n7954 1.57603
R30170 VDD.n8061 VDD.n8059 1.57603
R30171 VDD.n2356 VDD.n2317 1.56483
R30172 VDD.n1441 VDD.t3074 1.55829
R30173 VDD.n804 VDD.t4124 1.55829
R30174 VDD.n803 VDD.t3836 1.55829
R30175 VDD.n1479 VDD.t3030 1.55829
R30176 VDD.n814 VDD.t2764 1.55829
R30177 VDD.n6014 VDD.n6013 1.52779
R30178 VDD.n7005 VDD.n2376 1.5005
R30179 VDD.n6976 VDD.n6975 1.5005
R30180 VDD.n6978 VDD.n6977 1.5005
R30181 VDD.n7023 VDD.n7022 1.5005
R30182 VDD.n6959 VDD.n6958 1.5005
R30183 VDD.n6549 VDD.n6548 1.5005
R30184 VDD.n6512 VDD.n6415 1.5005
R30185 VDD.n6536 VDD.n6535 1.5005
R30186 VDD.n6551 VDD.n6550 1.5005
R30187 VDD.n6497 VDD.n6496 1.5005
R30188 VDD.n6095 VDD.n6038 1.5005
R30189 VDD.n6117 VDD.n6116 1.5005
R30190 VDD.n6152 VDD.n6151 1.5005
R30191 VDD.n6075 VDD.n6074 1.5005
R30192 VDD.n6150 VDD.n6149 1.5005
R30193 VDD.n6798 VDD.n6797 1.5005
R30194 VDD.n6800 VDD.n6799 1.5005
R30195 VDD.n6848 VDD.n6847 1.5005
R30196 VDD.n6791 VDD.n6790 1.5005
R30197 VDD.n6823 VDD.n2405 1.5005
R30198 VDD.n8642 VDD.n8640 1.49396
R30199 VDD.n8701 VDD.n8699 1.49396
R30200 VDD.n1811 VDD.n1809 1.49396
R30201 VDD.n1867 VDD.n1865 1.49396
R30202 VDD.n5515 VDD.n5513 1.49396
R30203 VDD.n1959 VDD.n1957 1.49396
R30204 VDD.n2041 VDD.n2039 1.49396
R30205 VDD.n8751 VDD.n8749 1.49396
R30206 VDD.n8894 VDD.n8892 1.49396
R30207 VDD.n9067 VDD.n9065 1.49396
R30208 VDD.n8636 VDD.t2640 1.4705
R30209 VDD.t1808 VDD.n8636 1.4705
R30210 VDD.t2664 VDD.n12619 1.4705
R30211 VDD.n12619 VDD.t1465 1.4705
R30212 VDD.n12597 VDD.t753 1.4705
R30213 VDD.t4188 VDD.n12597 1.4705
R30214 VDD.n12590 VDD.t778 1.4705
R30215 VDD.t3828 VDD.n12590 1.4705
R30216 VDD.t846 VDD.n12547 1.4705
R30217 VDD.n12547 VDD.t4266 1.4705
R30218 VDD.t1291 VDD.n12553 1.4705
R30219 VDD.n12553 VDD.t3916 1.4705
R30220 VDD.n8653 VDD.t2734 1.4705
R30221 VDD.t1905 VDD.n8653 1.4705
R30222 VDD.n8647 VDD.t3190 1.4705
R30223 VDD.t1541 VDD.n8647 1.4705
R30224 VDD.n8674 VDD.t728 1.4705
R30225 VDD.t3681 VDD.n8674 1.4705
R30226 VDD.n8668 VDD.t764 1.4705
R30227 VDD.t3346 VDD.n8668 1.4705
R30228 VDD.n78 VDD.t3128 1.4705
R30229 VDD.t1853 VDD.n78 1.4705
R30230 VDD.n50 VDD.t3152 1.4705
R30231 VDD.t1492 VDD.n50 1.4705
R30232 VDD.n12503 VDD.t2423 1.4705
R30233 VDD.t796 VDD.n12503 1.4705
R30234 VDD.n93 VDD.t1997 1.4705
R30235 VDD.t2241 VDD.n93 1.4705
R30236 VDD.n8686 VDD.t4182 1.4705
R30237 VDD.t2683 VDD.n8686 1.4705
R30238 VDD.n8680 VDD.t3818 1.4705
R30239 VDD.t4048 VDD.n8680 1.4705
R30240 VDD.n8712 VDD.t4260 1.4705
R30241 VDD.t2788 VDD.n8712 1.4705
R30242 VDD.n8706 VDD.t1403 1.4705
R30243 VDD.t1632 VDD.n8706 1.4705
R30244 VDD.t2522 VDD.n12491 1.4705
R30245 VDD.n12491 VDD.t903 1.4705
R30246 VDD.t3772 VDD.n12497 1.4705
R30247 VDD.n12497 VDD.t3996 1.4705
R30248 VDD.n167 VDD.t4228 1.4705
R30249 VDD.t2730 VDD.n167 1.4705
R30250 VDD.n139 VDD.t3858 1.4705
R30251 VDD.t4078 VDD.n139 1.4705
R30252 VDD.n8724 VDD.t1851 1.4705
R30253 VDD.t4454 VDD.n8724 1.4705
R30254 VDD.n8718 VDD.t1487 1.4705
R30255 VDD.t1709 VDD.n8718 1.4705
R30256 VDD.n8745 VDD.t3850 1.4705
R30257 VDD.t2345 VDD.n8745 1.4705
R30258 VDD.n8739 VDD.t2097 1.4705
R30259 VDD.t2383 VDD.n8739 1.4705
R30260 VDD.n5720 VDD.t1754 1.4705
R30261 VDD.t4222 VDD.n5720 1.4705
R30262 VDD.t3591 VDD.n11035 1.4705
R30263 VDD.n11035 VDD.t1241 1.4705
R30264 VDD.t2614 VDD.n11024 1.4705
R30265 VDD.n11024 VDD.t3693 1.4705
R30266 VDD.n1777 VDD.t3946 1.4705
R30267 VDD.t581 VDD.n1777 1.4705
R30268 VDD.n1822 VDD.t3316 1.4705
R30269 VDD.t4452 VDD.n1822 1.4705
R30270 VDD.n1816 VDD.t1554 1.4705
R30271 VDD.t1357 VDD.n1816 1.4705
R30272 VDD.n5732 VDD.t1225 1.4705
R30273 VDD.t3648 VDD.n5732 1.4705
R30274 VDD.n5726 VDD.t1616 1.4705
R30275 VDD.t730 VDD.n5726 1.4705
R30276 VDD.n5775 VDD.t1661 1.4705
R30277 VDD.t1316 VDD.n5775 1.4705
R30278 VDD.n5747 VDD.t3490 1.4705
R30279 VDD.t2656 VDD.n5747 1.4705
R30280 VDD.n10981 VDD.t1385 1.4705
R30281 VDD.t1501 VDD.n10981 1.4705
R30282 VDD.n1828 VDD.t2887 1.4705
R30283 VDD.t2691 VDD.n1828 1.4705
R30284 VDD.t1329 VDD.n10969 1.4705
R30285 VDD.n10969 VDD.t1136 1.4705
R30286 VDD.t2518 VDD.n10975 1.4705
R30287 VDD.n10975 VDD.t3628 1.4705
R30288 VDD.n5787 VDD.t2364 1.4705
R30289 VDD.t1361 VDD.n5787 1.4705
R30290 VDD.n5781 VDD.t3524 1.4705
R30291 VDD.t2140 VDD.n5781 1.4705
R30292 VDD.n5808 VDD.t1727 1.4705
R30293 VDD.t869 VDD.n5808 1.4705
R30294 VDD.n5802 VDD.t1175 1.4705
R30295 VDD.t3984 VDD.n5802 1.4705
R30296 VDD.n1878 VDD.t2116 1.4705
R30297 VDD.t1900 VDD.n1878 1.4705
R30298 VDD.n1872 VDD.t3654 1.4705
R30299 VDD.t703 VDD.n1872 1.4705
R30300 VDD.n10926 VDD.t3355 1.4705
R30301 VDD.t3200 VDD.n10926 1.4705
R30302 VDD.n1893 VDD.t4402 1.4705
R30303 VDD.t1443 VDD.n1893 1.4705
R30304 VDD.n5842 VDD.t3593 1.4705
R30305 VDD.t2775 VDD.n5842 1.4705
R30306 VDD.n5814 VDD.t644 1.4705
R30307 VDD.t3458 VDD.n5814 1.4705
R30308 VDD.n5863 VDD.t3750 1.4705
R30309 VDD.t2925 VDD.n5863 1.4705
R30310 VDD.n5857 VDD.t1842 1.4705
R30311 VDD.t4626 VDD.n5857 1.4705
R30312 VDD.t3571 VDD.n10914 1.4705
R30313 VDD.n10914 VDD.t3369 1.4705
R30314 VDD.t3568 VDD.n10920 1.4705
R30315 VDD.n10920 VDD.t572 1.4705
R30316 VDD.n5526 VDD.t3399 1.4705
R30317 VDD.t4562 VDD.n5526 1.4705
R30318 VDD.n5520 VDD.t608 1.4705
R30319 VDD.t2973 VDD.n5520 1.4705
R30320 VDD.n5875 VDD.t1887 1.4705
R30321 VDD.t4676 VDD.n5875 1.4705
R30322 VDD.n5869 VDD.t3697 1.4705
R30323 VDD.t933 VDD.n5869 1.4705
R30324 VDD.t1339 VDD.n5659 1.4705
R30325 VDD.n5659 VDD.t2817 1.4705
R30326 VDD.t3214 VDD.n5665 1.4705
R30327 VDD.n5665 VDD.t867 1.4705
R30328 VDD.n10871 VDD.t4164 1.4705
R30329 VDD.t2262 VDD.n10871 1.4705
R30330 VDD.t1379 VDD.n5508 1.4705
R30331 VDD.n5508 VDD.t2259 1.4705
R30332 VDD.t665 VDD.n10859 1.4705
R30333 VDD.n10859 VDD.t2543 1.4705
R30334 VDD.t2095 VDD.n10865 1.4705
R30335 VDD.n10865 VDD.t3014 1.4705
R30336 VDD.t3906 VDD.n5619 1.4705
R30337 VDD.n5619 VDD.t2983 1.4705
R30338 VDD.t1513 VDD.n5625 1.4705
R30339 VDD.n5625 VDD.t3391 1.4705
R30340 VDD.t3365 VDD.n5598 1.4705
R30341 VDD.n5598 VDD.t4724 1.4705
R30342 VDD.t3748 VDD.n5604 1.4705
R30343 VDD.n5604 VDD.t2922 1.4705
R30344 VDD.n1970 VDD.t1406 1.4705
R30345 VDD.t3679 VDD.n1970 1.4705
R30346 VDD.n1964 VDD.t3888 1.4705
R30347 VDD.t3676 VDD.n1964 1.4705
R30348 VDD.n10813 VDD.t3290 1.4705
R30349 VDD.t4436 VDD.n10813 1.4705
R30350 VDD.n1985 VDD.t4634 1.4705
R30351 VDD.t4432 VDD.n1985 1.4705
R30352 VDD.t1391 VDD.n5577 1.4705
R30353 VDD.n5577 VDD.t4210 1.4705
R30354 VDD.t3266 VDD.n5583 1.4705
R30355 VDD.n5583 VDD.t2378 1.4705
R30356 VDD.n8108 VDD.t862 1.4705
R30357 VDD.t4106 VDD.n8108 1.4705
R30358 VDD.n8102 VDD.t2082 1.4705
R30359 VDD.t672 VDD.n8102 1.4705
R30360 VDD.t2937 VDD.n10801 1.4705
R30361 VDD.n10801 VDD.t2740 1.4705
R30362 VDD.t3938 VDD.n10807 1.4705
R30363 VDD.n10807 VDD.t1001 1.4705
R30364 VDD.n2052 VDD.t3614 1.4705
R30365 VDD.t3424 VDD.n2052 1.4705
R30366 VDD.n2046 VDD.t4682 1.4705
R30367 VDD.t1712 VDD.n2046 1.4705
R30368 VDD.n8120 VDD.t4450 1.4705
R30369 VDD.t3550 VDD.n8120 1.4705
R30370 VDD.n8114 VDD.t1495 1.4705
R30371 VDD.t4298 VDD.n8114 1.4705
R30372 VDD.n8163 VDD.t2147 1.4705
R30373 VDD.t1204 VDD.n8163 1.4705
R30374 VDD.n8135 VDD.t3367 1.4705
R30375 VDD.t1980 VDD.n8135 1.4705
R30376 VDD.t670 VDD.n10770 1.4705
R30377 VDD.n10770 VDD.t4616 1.4705
R30378 VDD.n2058 VDD.t1731 1.4705
R30379 VDD.t3040 VDD.n2058 1.4705
R30380 VDD.t3964 VDD.n7099 1.4705
R30381 VDD.n7099 VDD.t3108 1.4705
R30382 VDD.n7100 VDD.t1147 1.4705
R30383 VDD.n7100 VDD.t3964 1.4705
R30384 VDD.t3970 VDD.n7104 1.4705
R30385 VDD.n7104 VDD.t1147 1.4705
R30386 VDD.n7107 VDD.t4700 1.4705
R30387 VDD.n7107 VDD.t3046 1.4705
R30388 VDD.t1920 VDD.n7112 1.4705
R30389 VDD.n7112 VDD.t4700 1.4705
R30390 VDD.t3725 VDD.n7117 1.4705
R30391 VDD.n7117 VDD.t2425 1.4705
R30392 VDD.n7118 VDD.t972 1.4705
R30393 VDD.n7118 VDD.t3725 1.4705
R30394 VDD.t2247 VDD.n7122 1.4705
R30395 VDD.n7122 VDD.t972 1.4705
R30396 VDD.n7094 VDD.t1831 1.4705
R30397 VDD.t970 VDD.n7094 1.4705
R30398 VDD.n7092 VDD.t3282 1.4705
R30399 VDD.t1831 VDD.n7092 1.4705
R30400 VDD.n7091 VDD.t1839 1.4705
R30401 VDD.t3282 VDD.n7091 1.4705
R30402 VDD.n7088 VDD.t2701 1.4705
R30403 VDD.t901 VDD.n7088 1.4705
R30404 VDD.n2330 VDD.t4004 1.4705
R30405 VDD.t2701 VDD.n2330 1.4705
R30406 VDD.n2328 VDD.t1614 1.4705
R30407 VDD.t4392 VDD.n2328 1.4705
R30408 VDD.n2326 VDD.t3082 1.4705
R30409 VDD.t1614 VDD.n2326 1.4705
R30410 VDD.n2325 VDD.t4284 1.4705
R30411 VDD.t3082 VDD.n2325 1.4705
R30412 VDD.t2831 VDD.n7073 1.4705
R30413 VDD.n7073 VDD.t1814 1.4705
R30414 VDD.n7074 VDD.t4142 1.4705
R30415 VDD.n7074 VDD.t2831 1.4705
R30416 VDD.t2839 VDD.n7078 1.4705
R30417 VDD.n7078 VDD.t4142 1.4705
R30418 VDD.n7081 VDD.t3520 1.4705
R30419 VDD.n7081 VDD.t1735 1.4705
R30420 VDD.n7065 VDD.t732 1.4705
R30421 VDD.t3520 VDD.n7065 1.4705
R30422 VDD.n7060 VDD.t2616 1.4705
R30423 VDD.t1132 VDD.n7060 1.4705
R30424 VDD.n7055 VDD.t3908 1.4705
R30425 VDD.n7055 VDD.t2616 1.4705
R30426 VDD.n7054 VDD.t1022 1.4705
R30427 VDD.t3908 VDD.n7054 1.4705
R30428 VDD.t2929 VDD.n6660 1.4705
R30429 VDD.n6660 VDD.t1435 1.4705
R30430 VDD.n6661 VDD.t3756 1.4705
R30431 VDD.n6661 VDD.t2929 1.4705
R30432 VDD.t1314 VDD.n6665 1.4705
R30433 VDD.n6665 VDD.t3756 1.4705
R30434 VDD.n6668 VDD.t3192 1.4705
R30435 VDD.n6668 VDD.t831 1.4705
R30436 VDD.t4492 VDD.n6673 1.4705
R30437 VDD.n6673 VDD.t3192 1.4705
R30438 VDD.t1110 VDD.n6678 1.4705
R30439 VDD.n6678 VDD.t4012 1.4705
R30440 VDD.n6679 VDD.t2576 1.4705
R30441 VDD.n6679 VDD.t1110 1.4705
R30442 VDD.t3415 VDD.n6683 1.4705
R30443 VDD.n6683 VDD.t2576 1.4705
R30444 VDD.n7070 VDD.t2847 1.4705
R30445 VDD.n7070 VDD.t1833 1.4705
R30446 VDD.n7068 VDD.t4158 1.4705
R30447 VDD.t2847 VDD.n7068 1.4705
R30448 VDD.n7067 VDD.t2853 1.4705
R30449 VDD.t4158 VDD.n7067 1.4705
R30450 VDD.t3532 VDD.n2334 1.4705
R30451 VDD.t1750 VDD.n2334 1.4705
R30452 VDD.t758 VDD.n7062 1.4705
R30453 VDD.n7062 VDD.t3532 1.4705
R30454 VDD.n7058 VDD.t2632 1.4705
R30455 VDD.n7058 VDD.t1145 1.4705
R30456 VDD.n7057 VDD.t3926 1.4705
R30457 VDD.t2632 VDD.n7057 1.4705
R30458 VDD.n7052 VDD.t1034 1.4705
R30459 VDD.n7052 VDD.t3926 1.4705
R30460 VDD.n6654 VDD.t2957 1.4705
R30461 VDD.t1467 VDD.n6654 1.4705
R30462 VDD.n6652 VDD.t3776 1.4705
R30463 VDD.t2957 VDD.n6652 1.4705
R30464 VDD.n6651 VDD.t1327 1.4705
R30465 VDD.t3776 VDD.n6651 1.4705
R30466 VDD.t3212 VDD.n6670 1.4705
R30467 VDD.n6670 VDD.t858 1.4705
R30468 VDD.n6671 VDD.t4506 1.4705
R30469 VDD.n6671 VDD.t3212 1.4705
R30470 VDD.n6646 VDD.t1121 1.4705
R30471 VDD.t4026 VDD.n6646 1.4705
R30472 VDD.n6644 VDD.t2594 1.4705
R30473 VDD.t1121 VDD.n6644 1.4705
R30474 VDD.n6643 VDD.t3430 1.4705
R30475 VDD.t2594 VDD.n6643 1.4705
R30476 VDD.t4554 VDD.n7027 1.4705
R30477 VDD.n7027 VDD.t3270 1.4705
R30478 VDD.n7028 VDD.t1312 1.4705
R30479 VDD.n7028 VDD.t4554 1.4705
R30480 VDD.t3150 VDD.n7032 1.4705
R30481 VDD.n7032 VDD.t1312 1.4705
R30482 VDD.n7035 VDD.t723 1.4705
R30483 VDD.n7035 VDD.t2650 1.4705
R30484 VDD.t2102 VDD.n6717 1.4705
R30485 VDD.n6717 VDD.t723 1.4705
R30486 VDD.n6720 VDD.t2945 1.4705
R30487 VDD.n6720 VDD.t1552 1.4705
R30488 VDD.t4244 VDD.n6724 1.4705
R30489 VDD.n6724 VDD.t2945 1.4705
R30490 VDD.n6725 VDD.t1005 1.4705
R30491 VDD.n6725 VDD.t4244 1.4705
R30492 VDD.n6742 VDD.t223 1.4705
R30493 VDD.n6742 VDD.t89 1.4705
R30494 VDD.n6750 VDD.t243 1.4705
R30495 VDD.n6750 VDD.t146 1.4705
R30496 VDD.n6874 VDD.t4474 1.4705
R30497 VDD.t3589 VDD.n6874 1.4705
R30498 VDD.n6870 VDD.t1688 1.4705
R30499 VDD.n6870 VDD.t4474 1.4705
R30500 VDD.n6869 VDD.t4478 1.4705
R30501 VDD.t1688 VDD.n6869 1.4705
R30502 VDD.n6864 VDD.t1093 1.4705
R30503 VDD.t3514 VDD.n6864 1.4705
R30504 VDD.n6859 VDD.t2555 1.4705
R30505 VDD.n6859 VDD.t1093 1.4705
R30506 VDD.n6856 VDD.t4268 1.4705
R30507 VDD.t2975 VDD.n6856 1.4705
R30508 VDD.n6852 VDD.t1461 1.4705
R30509 VDD.n6852 VDD.t4268 1.4705
R30510 VDD.n6851 VDD.t2843 1.4705
R30511 VDD.t1461 VDD.n6851 1.4705
R30512 VDD.n6954 VDD.t253 1.4705
R30513 VDD.n6954 VDD.t95 1.4705
R30514 VDD.n6955 VDD.t130 1.4705
R30515 VDD.n6955 VDD.t205 1.4705
R30516 VDD.n6922 VDD.t270 1.4705
R30517 VDD.n6922 VDD.t119 1.4705
R30518 VDD.n6923 VDD.t152 1.4705
R30519 VDD.n6923 VDD.t224 1.4705
R30520 VDD.n7014 VDD.t220 1.4705
R30521 VDD.n7014 VDD.t264 1.4705
R30522 VDD.n7016 VDD.t218 1.4705
R30523 VDD.n7016 VDD.t143 1.4705
R30524 VDD.n7018 VDD.t226 1.4705
R30525 VDD.n7018 VDD.t63 1.4705
R30526 VDD.n7020 VDD.t80 1.4705
R30527 VDD.n7020 VDD.t154 1.4705
R30528 VDD.n2382 VDD.t211 1.4705
R30529 VDD.n2382 VDD.t282 1.4705
R30530 VDD.n2380 VDD.t48 1.4705
R30531 VDD.n2380 VDD.t162 1.4705
R30532 VDD.n2378 VDD.t69 1.4705
R30533 VDD.n2378 VDD.t151 1.4705
R30534 VDD.n2377 VDD.t182 1.4705
R30535 VDD.n2377 VDD.t230 1.4705
R30536 VDD.n6995 VDD.t201 1.4705
R30537 VDD.n6995 VDD.t250 1.4705
R30538 VDD.n6990 VDD.t199 1.4705
R30539 VDD.n6990 VDD.t125 1.4705
R30540 VDD.n6985 VDD.t212 1.4705
R30541 VDD.n6985 VDD.t283 1.4705
R30542 VDD.n6980 VDD.t50 1.4705
R30543 VDD.n6980 VDD.t136 1.4705
R30544 VDD.n6898 VDD.t193 1.4705
R30545 VDD.n6898 VDD.t268 1.4705
R30546 VDD.n6893 VDD.t273 1.4705
R30547 VDD.n6893 VDD.t148 1.4705
R30548 VDD.n6888 VDD.t284 1.4705
R30549 VDD.n6888 VDD.t132 1.4705
R30550 VDD.n6886 VDD.t164 1.4705
R30551 VDD.n6886 VDD.t216 1.4705
R30552 VDD.n6967 VDD.t123 1.4705
R30553 VDD.n6967 VDD.t170 1.4705
R30554 VDD.n6969 VDD.t121 1.4705
R30555 VDD.n6969 VDD.t272 1.4705
R30556 VDD.n6971 VDD.t135 1.4705
R30557 VDD.n6971 VDD.t208 1.4705
R30558 VDD.n6973 VDD.t219 1.4705
R30559 VDD.n6973 VDD.t281 1.4705
R30560 VDD.n6965 VDD.t116 1.4705
R30561 VDD.n6965 VDD.t191 1.4705
R30562 VDD.n6963 VDD.t200 1.4705
R30563 VDD.n6963 VDD.t54 1.4705
R30564 VDD.n6961 VDD.t213 1.4705
R30565 VDD.n6961 VDD.t276 1.4705
R30566 VDD.n6960 VDD.t83 1.4705
R30567 VDD.n6960 VDD.t138 1.4705
R30568 VDD.n6947 VDD.t263 1.4705
R30569 VDD.n6947 VDD.t85 1.4705
R30570 VDD.n6942 VDD.t262 1.4705
R30571 VDD.n6942 VDD.t187 1.4705
R30572 VDD.n6937 VDD.t274 1.4705
R30573 VDD.n6937 VDD.t127 1.4705
R30574 VDD.n6932 VDD.t133 1.4705
R30575 VDD.n6932 VDD.t204 1.4705
R30576 VDD.n6917 VDD.t261 1.4705
R30577 VDD.n6917 VDD.t108 1.4705
R30578 VDD.n6912 VDD.t113 1.4705
R30579 VDD.n6912 VDD.t210 1.4705
R30580 VDD.n6907 VDD.t129 1.4705
R30581 VDD.n6907 VDD.t198 1.4705
R30582 VDD.n6905 VDD.t229 1.4705
R30583 VDD.n6905 VDD.t275 1.4705
R30584 VDD.n7006 VDD.t117 1.4705
R30585 VDD.n7006 VDD.t195 1.4705
R30586 VDD.n7007 VDD.t285 1.4705
R30587 VDD.n7007 VDD.t141 1.4705
R30588 VDD.n7000 VDD.t142 1.4705
R30589 VDD.n7000 VDD.t217 1.4705
R30590 VDD.n7001 VDD.t79 1.4705
R30591 VDD.n7001 VDD.t159 1.4705
R30592 VDD.t4058 VDD.n5238 1.4705
R30593 VDD.n5238 VDD.t2762 1.4705
R30594 VDD.n5239 VDD.t808 1.4705
R30595 VDD.n5239 VDD.t4058 1.4705
R30596 VDD.t2636 VDD.n5243 1.4705
R30597 VDD.n5243 VDD.t808 1.4705
R30598 VDD.n5246 VDD.t4340 1.4705
R30599 VDD.n5246 VDD.t2040 1.4705
R30600 VDD.t1532 VDD.n5251 1.4705
R30601 VDD.n5251 VDD.t4340 1.4705
R30602 VDD.t2389 VDD.n5256 1.4705
R30603 VDD.n5256 VDD.t1045 1.4705
R30604 VDD.n5257 VDD.t3691 1.4705
R30605 VDD.n5257 VDD.t2389 1.4705
R30606 VDD.t4572 VDD.n5261 1.4705
R30607 VDD.n5261 VDD.t3691 1.4705
R30608 VDD.n5235 VDD.t1947 1.4705
R30609 VDD.n5235 VDD.t4726 1.4705
R30610 VDD.n5233 VDD.t2955 1.4705
R30611 VDD.t1947 VDD.n5233 1.4705
R30612 VDD.n5232 VDD.t4578 1.4705
R30613 VDD.t2955 VDD.n5232 1.4705
R30614 VDD.n5229 VDD.t2278 1.4705
R30615 VDD.t4102 VDD.n5229 1.4705
R30616 VDD.n5228 VDD.t3622 1.4705
R30617 VDD.t2278 VDD.n5228 1.4705
R30618 VDD.n5226 VDD.t4364 1.4705
R30619 VDD.t3162 VDD.n5226 1.4705
R30620 VDD.n5224 VDD.t1575 1.4705
R30621 VDD.t4364 VDD.n5224 1.4705
R30622 VDD.n5223 VDD.t2592 1.4705
R30623 VDD.t1575 VDD.n5223 1.4705
R30624 VDD.n6359 VDD.t566 1.4705
R30625 VDD.t4418 VDD.n6359 1.4705
R30626 VDD.n6354 VDD.t1986 1.4705
R30627 VDD.n6354 VDD.t566 1.4705
R30628 VDD.n6353 VDD.t4300 1.4705
R30629 VDD.t1986 VDD.n6353 1.4705
R30630 VDD.n6348 VDD.t1934 1.4705
R30631 VDD.t3788 VDD.n6348 1.4705
R30632 VDD.n6343 VDD.t2334 1.4705
R30633 VDD.n6343 VDD.t1934 1.4705
R30634 VDD.n6340 VDD.t4088 1.4705
R30635 VDD.t3230 VDD.n6340 1.4705
R30636 VDD.n6335 VDD.t1272 1.4705
R30637 VDD.n6335 VDD.t4088 1.4705
R30638 VDD.n6334 VDD.t4096 1.4705
R30639 VDD.t1272 VDD.n6334 1.4705
R30640 VDD.n6357 VDD.t3660 1.4705
R30641 VDD.n6357 VDD.t3338 1.4705
R30642 VDD.n6356 VDD.t915 1.4705
R30643 VDD.t3660 VDD.n6356 1.4705
R30644 VDD.n6351 VDD.t3264 1.4705
R30645 VDD.n6351 VDD.t915 1.4705
R30646 VDD.n6346 VDD.t873 1.4705
R30647 VDD.n6346 VDD.t2786 1.4705
R30648 VDD.n6345 VDD.t1167 1.4705
R30649 VDD.t873 VDD.n6345 1.4705
R30650 VDD.n6338 VDD.t3052 1.4705
R30651 VDD.n6338 VDD.t2086 1.4705
R30652 VDD.n6337 VDD.t4350 1.4705
R30653 VDD.t3052 VDD.n6337 1.4705
R30654 VDD.n6332 VDD.t3056 1.4705
R30655 VDD.n6332 VDD.t4350 1.4705
R30656 VDD.t2038 VDD.n5448 1.4705
R30657 VDD.n5448 VDD.t628 1.4705
R30658 VDD.n5449 VDD.t3018 1.4705
R30659 VDD.n5449 VDD.t2038 1.4705
R30660 VDD.t4668 VDD.n5453 1.4705
R30661 VDD.n5453 VDD.t3018 1.4705
R30662 VDD.n5456 VDD.t2387 1.4705
R30663 VDD.n5456 VDD.t4176 1.4705
R30664 VDD.t3689 VDD.n5461 1.4705
R30665 VDD.n5461 VDD.t2387 1.4705
R30666 VDD.t4438 VDD.n5466 1.4705
R30667 VDD.n5466 VDD.t4542 1.4705
R30668 VDD.n5467 VDD.t1651 1.4705
R30669 VDD.n5467 VDD.t4438 1.4705
R30670 VDD.t3994 VDD.n5471 1.4705
R30671 VDD.n5471 VDD.t1651 1.4705
R30672 VDD.n5392 VDD.t949 1.4705
R30673 VDD.t3701 VDD.n5392 1.4705
R30674 VDD.n5390 VDD.t1810 1.4705
R30675 VDD.t949 VDD.n5390 1.4705
R30676 VDD.n5389 VDD.t3583 1.4705
R30677 VDD.t1810 VDD.n5389 1.4705
R30678 VDD.n5386 VDD.t1193 1.4705
R30679 VDD.t3122 VDD.n5386 1.4705
R30680 VDD.n5385 VDD.t2678 1.4705
R30681 VDD.t1193 VDD.n5385 1.4705
R30682 VDD.n5383 VDD.t3359 1.4705
R30683 VDD.t3500 VDD.n5383 1.4705
R30684 VDD.n5381 VDD.t4714 1.4705
R30685 VDD.t3359 VDD.n5381 1.4705
R30686 VDD.n5380 VDD.t2971 1.4705
R30687 VDD.t4714 VDD.n5380 1.4705
R30688 VDD.n6592 VDD.t3758 1.4705
R30689 VDD.t2458 VDD.n6592 1.4705
R30690 VDD.n6588 VDD.t4648 1.4705
R30691 VDD.n6588 VDD.t3758 1.4705
R30692 VDD.n6587 VDD.t2282 1.4705
R30693 VDD.t4648 VDD.n6587 1.4705
R30694 VDD.n6582 VDD.t4052 1.4705
R30695 VDD.t1700 VDD.n6582 1.4705
R30696 VDD.t1243 VDD.n5925 1.4705
R30697 VDD.n5925 VDD.t4052 1.4705
R30698 VDD.t2028 VDD.n5930 1.4705
R30699 VDD.n5930 VDD.t2171 1.4705
R30700 VDD.n5931 VDD.t3413 1.4705
R30701 VDD.n5931 VDD.t2028 1.4705
R30702 VDD.t1528 VDD.n5935 1.4705
R30703 VDD.n5935 VDD.t3413 1.4705
R30704 VDD.t1115 VDD.n6236 1.4705
R30705 VDD.n6236 VDD.t3900 1.4705
R30706 VDD.n6237 VDD.t2036 1.4705
R30707 VDD.n6237 VDD.t1115 1.4705
R30708 VDD.t3770 VDD.n6241 1.4705
R30709 VDD.n6241 VDD.t2036 1.4705
R30710 VDD.n6244 VDD.t1389 1.4705
R30711 VDD.n6244 VDD.t3292 1.4705
R30712 VDD.t2865 VDD.n6249 1.4705
R30713 VDD.n6249 VDD.t1389 1.4705
R30714 VDD.t3540 VDD.n6254 1.4705
R30715 VDD.n6254 VDD.t3664 1.4705
R30716 VDD.n6255 VDD.t774 1.4705
R30717 VDD.n6255 VDD.t3540 1.4705
R30718 VDD.t3142 VDD.n6259 1.4705
R30719 VDD.n6259 VDD.t774 1.4705
R30720 VDD.t3862 VDD.n6272 1.4705
R30721 VDD.n6272 VDD.t3534 1.4705
R30722 VDD.n6273 VDD.t1084 1.4705
R30723 VDD.n6273 VDD.t3862 1.4705
R30724 VDD.t3411 VDD.n6277 1.4705
R30725 VDD.n6277 VDD.t1084 1.4705
R30726 VDD.n6280 VDD.t1038 1.4705
R30727 VDD.n6280 VDD.t2963 1.4705
R30728 VDD.t1347 VDD.n6285 1.4705
R30729 VDD.n6285 VDD.t1038 1.4705
R30730 VDD.t3228 VDD.n6290 1.4705
R30731 VDD.n6290 VDD.t2309 1.4705
R30732 VDD.n6291 VDD.t4520 1.4705
R30733 VDD.n6291 VDD.t3228 1.4705
R30734 VDD.t3234 VDD.n6295 1.4705
R30735 VDD.n6295 VDD.t4520 1.4705
R30736 VDD.n6233 VDD.t1125 1.4705
R30737 VDD.n6233 VDD.t3918 1.4705
R30738 VDD.n6231 VDD.t2056 1.4705
R30739 VDD.t1125 VDD.n6231 1.4705
R30740 VDD.n6230 VDD.t3786 1.4705
R30741 VDD.t2056 VDD.n6230 1.4705
R30742 VDD.n6227 VDD.t1401 1.4705
R30743 VDD.t3300 VDD.n6227 1.4705
R30744 VDD.n6226 VDD.t2877 1.4705
R30745 VDD.t1401 VDD.n6226 1.4705
R30746 VDD.n6224 VDD.t3552 1.4705
R30747 VDD.t3683 VDD.n6224 1.4705
R30748 VDD.n6222 VDD.t785 1.4705
R30749 VDD.t3552 VDD.n6222 1.4705
R30750 VDD.n6221 VDD.t3156 1.4705
R30751 VDD.t785 VDD.n6221 1.4705
R30752 VDD.n6214 VDD.t3876 1.4705
R30753 VDD.t3544 VDD.n6214 1.4705
R30754 VDD.n6212 VDD.t1102 1.4705
R30755 VDD.t3876 VDD.n6212 1.4705
R30756 VDD.n6211 VDD.t3432 1.4705
R30757 VDD.t1102 VDD.n6211 1.4705
R30758 VDD.n6208 VDD.t1063 1.4705
R30759 VDD.t2979 VDD.n6208 1.4705
R30760 VDD.n6207 VDD.t1363 1.4705
R30761 VDD.t1063 VDD.n6207 1.4705
R30762 VDD.n6205 VDD.t3242 1.4705
R30763 VDD.t2332 VDD.n6205 1.4705
R30764 VDD.n6203 VDD.t4526 1.4705
R30765 VDD.t3242 VDD.n6203 1.4705
R30766 VDD.n6202 VDD.t3248 1.4705
R30767 VDD.t4526 VDD.n6202 1.4705
R30768 VDD.t2416 VDD.n5954 1.4705
R30769 VDD.n5954 VDD.t2009 1.4705
R30770 VDD.n5955 VDD.t3721 1.4705
R30771 VDD.n5955 VDD.t2416 1.4705
R30772 VDD.t1863 VDD.n5959 1.4705
R30773 VDD.n5959 VDD.t3721 1.4705
R30774 VDD.n5962 VDD.t3674 1.4705
R30775 VDD.n5962 VDD.t1336 1.4705
R30776 VDD.t4024 VDD.n5967 1.4705
R30777 VDD.n5967 VDD.t3674 1.4705
R30778 VDD.t1636 VDD.n5972 1.4705
R30779 VDD.n5972 VDD.t762 1.4705
R30780 VDD.n5973 VDD.t3098 1.4705
R30781 VDD.n5973 VDD.t1636 1.4705
R30782 VDD.t1645 VDD.n5977 1.4705
R30783 VDD.n5977 VDD.t3098 1.4705
R30784 VDD.t928 VDD.n6383 1.4705
R30785 VDD.n6383 VDD.t4720 1.4705
R30786 VDD.n6384 VDD.t2340 1.4705
R30787 VDD.n6384 VDD.t928 1.4705
R30788 VDD.t4570 VDD.n6388 1.4705
R30789 VDD.n6388 VDD.t2340 1.4705
R30790 VDD.n6391 VDD.t2270 1.4705
R30791 VDD.n6391 VDD.t4094 1.4705
R30792 VDD.t2660 VDD.n5996 1.4705
R30793 VDD.n5996 VDD.t2270 1.4705
R30794 VDD.t4362 VDD.n6001 1.4705
R30795 VDD.n6001 VDD.t3482 1.4705
R30796 VDD.n6002 VDD.t1566 1.4705
R30797 VDD.n6002 VDD.t4362 1.4705
R30798 VDD.t4368 VDD.n6006 1.4705
R30799 VDD.n6006 VDD.t1566 1.4705
R30800 VDD.n5320 VDD.t3044 1.4705
R30801 VDD.t2717 VDD.n5320 1.4705
R30802 VDD.n5318 VDD.t4342 1.4705
R30803 VDD.t3044 VDD.n5318 1.4705
R30804 VDD.n5317 VDD.t2590 1.4705
R30805 VDD.t4342 VDD.n5317 1.4705
R30806 VDD.t4296 VDD.n5314 1.4705
R30807 VDD.t1978 VDD.n5314 1.4705
R30808 VDD.t4614 VDD.n5994 1.4705
R30809 VDD.n5994 VDD.t4296 1.4705
R30810 VDD.n5993 VDD.t2328 1.4705
R30811 VDD.t1343 VDD.n5993 1.4705
R30812 VDD.n5991 VDD.t3640 1.4705
R30813 VDD.t2328 VDD.n5991 1.4705
R30814 VDD.n5990 VDD.t2338 1.4705
R30815 VDD.t3640 VDD.n5990 1.4705
R30816 VDD.t2393 VDD.n5337 1.4705
R30817 VDD.n5337 VDD.t960 1.4705
R30818 VDD.n5338 VDD.t3278 1.4705
R30819 VDD.n5338 VDD.t2393 1.4705
R30820 VDD.t821 VDD.n5342 1.4705
R30821 VDD.n5342 VDD.t3278 1.4705
R30822 VDD.n5345 VDD.t2695 1.4705
R30823 VDD.n5345 VDD.t4442 1.4705
R30824 VDD.t3998 VDD.n5350 1.4705
R30825 VDD.n5350 VDD.t2695 1.4705
R30826 VDD.t4732 VDD.n5355 1.4705
R30827 VDD.n5355 VDD.t714 1.4705
R30828 VDD.n5356 VDD.t1960 1.4705
R30829 VDD.n5356 VDD.t4732 1.4705
R30830 VDD.t4278 VDD.n5360 1.4705
R30831 VDD.n5360 VDD.t1960 1.4705
R30832 VDD.n5334 VDD.t4370 1.4705
R30833 VDD.n5334 VDD.t3078 1.4705
R30834 VDD.n5332 VDD.t1123 1.4705
R30835 VDD.t4370 VDD.n5332 1.4705
R30836 VDD.n5331 VDD.t2961 1.4705
R30837 VDD.t1123 VDD.n5331 1.4705
R30838 VDD.n5328 VDD.t4662 1.4705
R30839 VDD.t2431 VDD.n5328 1.4705
R30840 VDD.n5327 VDD.t1872 1.4705
R30841 VDD.t4662 VDD.n5327 1.4705
R30842 VDD.n5325 VDD.t2736 1.4705
R30843 VDD.t2861 VDD.n5325 1.4705
R30844 VDD.n5323 VDD.t4040 1.4705
R30845 VDD.t2736 VDD.n5323 1.4705
R30846 VDD.n5322 VDD.t2200 1.4705
R30847 VDD.t4040 VDD.n5322 1.4705
R30848 VDD.n6411 VDD.t1417 1.4705
R30849 VDD.t1108 VDD.n6411 1.4705
R30850 VDD.n6407 VDD.t2899 1.4705
R30851 VDD.n6407 VDD.t1417 1.4705
R30852 VDD.n6406 VDD.t1003 1.4705
R30853 VDD.t2899 VDD.n6406 1.4705
R30854 VDD.n6401 VDD.t2859 1.4705
R30855 VDD.t4596 VDD.n6401 1.4705
R30856 VDD.t3170 VDD.n6160 1.4705
R30857 VDD.n6160 VDD.t2859 1.4705
R30858 VDD.t768 VDD.n6165 1.4705
R30859 VDD.n6165 VDD.t4014 1.4705
R30860 VDD.n6166 VDD.t2132 1.4705
R30861 VDD.n6166 VDD.t768 1.4705
R30862 VDD.t776 VDD.n6170 1.4705
R30863 VDD.n6170 VDD.t2132 1.4705
R30864 VDD.t2947 VDD.n6564 1.4705
R30865 VDD.n6564 VDD.t1451 1.4705
R30866 VDD.n6565 VDD.t3768 1.4705
R30867 VDD.n6565 VDD.t2947 1.4705
R30868 VDD.t1318 VDD.n6569 1.4705
R30869 VDD.n6569 VDD.t3768 1.4705
R30870 VDD.n6572 VDD.t3210 1.4705
R30871 VDD.n6572 VDD.t850 1.4705
R30872 VDD.t4500 VDD.n6027 1.4705
R30873 VDD.n6027 VDD.t3210 1.4705
R30874 VDD.n6030 VDD.t1119 1.4705
R30875 VDD.n6030 VDD.t1231 1.4705
R30876 VDD.t2582 VDD.n6034 1.4705
R30877 VDD.n6034 VDD.t1119 1.4705
R30878 VDD.n6035 VDD.t646 1.4705
R30879 VDD.n6035 VDD.t2582 1.4705
R30880 VDD.n6498 VDD.t4915 1.4705
R30881 VDD.n6498 VDD.t4850 1.4705
R30882 VDD.n6499 VDD.t4826 1.4705
R30883 VDD.n6499 VDD.t4956 1.4705
R30884 VDD.n6448 VDD.t4848 1.4705
R30885 VDD.n6448 VDD.t4832 1.4705
R30886 VDD.n6449 VDD.t4955 1.4705
R30887 VDD.n6449 VDD.t4939 1.4705
R30888 VDD.n6558 VDD.t4970 1.4705
R30889 VDD.n6558 VDD.t4907 1.4705
R30890 VDD.n6556 VDD.t4901 1.4705
R30891 VDD.n6556 VDD.t4819 1.4705
R30892 VDD.n6554 VDD.t4892 1.4705
R30893 VDD.n6554 VDD.t4897 1.4705
R30894 VDD.n6552 VDD.t4867 1.4705
R30895 VDD.n6552 VDD.t4953 1.4705
R30896 VDD.n5295 VDD.t4906 1.4705
R30897 VDD.n5295 VDD.t4890 1.4705
R30898 VDD.n5293 VDD.t4884 1.4705
R30899 VDD.n5293 VDD.t4966 1.4705
R30900 VDD.n5291 VDD.t4873 1.4705
R30901 VDD.n5291 VDD.t4825 1.4705
R30902 VDD.n5290 VDD.t4874 1.4705
R30903 VDD.n5290 VDD.t4933 1.4705
R30904 VDD.n6445 VDD.t4804 1.4705
R30905 VDD.n6445 VDD.t4919 1.4705
R30906 VDD.n6442 VDD.t4914 1.4705
R30907 VDD.n6442 VDD.t4829 1.4705
R30908 VDD.n6439 VDD.t4905 1.4705
R30909 VDD.n6439 VDD.t4910 1.4705
R30910 VDD.n6436 VDD.t4883 1.4705
R30911 VDD.n6436 VDD.t4965 1.4705
R30912 VDD.n6431 VDD.t4916 1.4705
R30913 VDD.n6431 VDD.t4902 1.4705
R30914 VDD.n6426 VDD.t4898 1.4705
R30915 VDD.n6426 VDD.t4801 1.4705
R30916 VDD.n6421 VDD.t4887 1.4705
R30917 VDD.n6421 VDD.t4840 1.4705
R30918 VDD.n6419 VDD.t4888 1.4705
R30919 VDD.n6419 VDD.t4946 1.4705
R30920 VDD.n6519 VDD.t4856 1.4705
R30921 VDD.n6519 VDD.t4806 1.4705
R30922 VDD.n6517 VDD.t4973 1.4705
R30923 VDD.n6517 VDD.t4899 1.4705
R30924 VDD.n6515 VDD.t4969 1.4705
R30925 VDD.n6515 VDD.t4972 1.4705
R30926 VDD.n6513 VDD.t4944 1.4705
R30927 VDD.n6513 VDD.t4836 1.4705
R30928 VDD.n6510 VDD.t4803 1.4705
R30929 VDD.n6510 VDD.t4967 1.4705
R30930 VDD.n6508 VDD.t4958 1.4705
R30931 VDD.n6508 VDD.t4854 1.4705
R30932 VDD.n6506 VDD.t4949 1.4705
R30933 VDD.n6506 VDD.t4909 1.4705
R30934 VDD.n6505 VDD.t4950 1.4705
R30935 VDD.n6505 VDD.t4822 1.4705
R30936 VDD.n6482 VDD.t4925 1.4705
R30937 VDD.n6482 VDD.t4864 1.4705
R30938 VDD.n6479 VDD.t4859 1.4705
R30939 VDD.n6479 VDD.t4971 1.4705
R30940 VDD.n6476 VDD.t4844 1.4705
R30941 VDD.n6476 VDD.t4852 1.4705
R30942 VDD.n6473 VDD.t4824 1.4705
R30943 VDD.n6473 VDD.t4912 1.4705
R30944 VDD.n6468 VDD.t4862 1.4705
R30945 VDD.n6468 VDD.t4841 1.4705
R30946 VDD.n6463 VDD.t4837 1.4705
R30947 VDD.n6463 VDD.t4923 1.4705
R30948 VDD.n6458 VDD.t4827 1.4705
R30949 VDD.n6458 VDD.t4800 1.4705
R30950 VDD.n6456 VDD.t4828 1.4705
R30951 VDD.n6456 VDD.t4896 1.4705
R30952 VDD.n6544 VDD.t4833 1.4705
R30953 VDD.n6544 VDD.t4962 1.4705
R30954 VDD.n6545 VDD.t4886 1.4705
R30955 VDD.n6545 VDD.t4821 1.4705
R30956 VDD.n6537 VDD.t4960 1.4705
R30957 VDD.n6537 VDD.t4945 1.4705
R30958 VDD.n6538 VDD.t4820 1.4705
R30959 VDD.n6538 VDD.t4810 1.4705
R30960 VDD.n6069 VDD.t4940 1.4705
R30961 VDD.n6069 VDD.t4831 1.4705
R30962 VDD.n6063 VDD.t4922 1.4705
R30963 VDD.n6063 VDD.t4818 1.4705
R30964 VDD.n6134 VDD.t4952 1.4705
R30965 VDD.n6134 VDD.t4891 1.4705
R30966 VDD.n6135 VDD.t4815 1.4705
R30967 VDD.n6135 VDD.t4935 1.4705
R30968 VDD.n6137 VDD.t4885 1.4705
R30969 VDD.n6137 VDD.t4808 1.4705
R30970 VDD.n6138 VDD.t4928 1.4705
R30971 VDD.n6138 VDD.t4845 1.4705
R30972 VDD.n6141 VDD.t4875 1.4705
R30973 VDD.n6141 VDD.t4879 1.4705
R30974 VDD.n6142 VDD.t4920 1.4705
R30975 VDD.n6142 VDD.t4924 1.4705
R30976 VDD.n6145 VDD.t4846 1.4705
R30977 VDD.n6145 VDD.t4934 1.4705
R30978 VDD.n6146 VDD.t4900 1.4705
R30979 VDD.n6146 VDD.t4805 1.4705
R30980 VDD.n6130 VDD.t4889 1.4705
R30981 VDD.n6130 VDD.t4872 1.4705
R30982 VDD.n6131 VDD.t4931 1.4705
R30983 VDD.n6131 VDD.t4918 1.4705
R30984 VDD.n6126 VDD.t4866 1.4705
R30985 VDD.n6126 VDD.t4947 1.4705
R30986 VDD.n6127 VDD.t4913 1.4705
R30987 VDD.n6127 VDD.t4814 1.4705
R30988 VDD.n6122 VDD.t4853 1.4705
R30989 VDD.n6122 VDD.t4816 1.4705
R30990 VDD.n6123 VDD.t4903 1.4705
R30991 VDD.n6123 VDD.t4861 1.4705
R30992 VDD.n6118 VDD.t4855 1.4705
R30993 VDD.n6118 VDD.t4917 1.4705
R30994 VDD.n6119 VDD.t4904 1.4705
R30995 VDD.n6119 VDD.t4963 1.4705
R30996 VDD.n6042 VDD.t4835 1.4705
R30997 VDD.n6042 VDD.t4968 1.4705
R30998 VDD.n6043 VDD.t4942 1.4705
R30999 VDD.n6043 VDD.t4881 1.4705
R31000 VDD.n6045 VDD.t4959 1.4705
R31001 VDD.n6045 VDD.t4882 1.4705
R31002 VDD.n6046 VDD.t4877 1.4705
R31003 VDD.n6046 VDD.t4807 1.4705
R31004 VDD.n6049 VDD.t4951 1.4705
R31005 VDD.n6049 VDD.t4957 1.4705
R31006 VDD.n6050 VDD.t4865 1.4705
R31007 VDD.n6050 VDD.t4871 1.4705
R31008 VDD.n6053 VDD.t4927 1.4705
R31009 VDD.n6053 VDD.t4823 1.4705
R31010 VDD.n6054 VDD.t4839 1.4705
R31011 VDD.n6054 VDD.t4926 1.4705
R31012 VDD.n6076 VDD.t4964 1.4705
R31013 VDD.n6076 VDD.t4948 1.4705
R31014 VDD.n6077 VDD.t4880 1.4705
R31015 VDD.n6077 VDD.t4863 1.4705
R31016 VDD.n6080 VDD.t4943 1.4705
R31017 VDD.n6080 VDD.t4834 1.4705
R31018 VDD.n6081 VDD.t4857 1.4705
R31019 VDD.n6081 VDD.t4941 1.4705
R31020 VDD.n6084 VDD.t4930 1.4705
R31021 VDD.n6084 VDD.t4895 1.4705
R31022 VDD.n6085 VDD.t4842 1.4705
R31023 VDD.n6085 VDD.t4812 1.4705
R31024 VDD.n6088 VDD.t4932 1.4705
R31025 VDD.n6088 VDD.t4813 1.4705
R31026 VDD.n6089 VDD.t4843 1.4705
R31027 VDD.n6089 VDD.t4911 1.4705
R31028 VDD.n6020 VDD.t4851 1.4705
R31029 VDD.n6020 VDD.t4802 1.4705
R31030 VDD.n6154 VDD.t4975 1.4705
R31031 VDD.n6154 VDD.t4961 1.4705
R31032 VDD.n6112 VDD.t4811 1.4705
R31033 VDD.n6112 VDD.t4894 1.4705
R31034 VDD.n6106 VDD.t4974 1.4705
R31035 VDD.n6106 VDD.t4876 1.4705
R31036 VDD.n6093 VDD.t4929 1.4705
R31037 VDD.n6093 VDD.t4870 1.4705
R31038 VDD.n6097 VDD.t4868 1.4705
R31039 VDD.n6097 VDD.t4849 1.4705
R31040 VDD.t2693 VDD.n7847 1.4705
R31041 VDD.n7847 VDD.t1202 1.4705
R31042 VDD.n7848 VDD.t1214 1.4705
R31043 VDD.n7848 VDD.t2693 1.4705
R31044 VDD.n2226 VDD.t1992 1.4705
R31045 VDD.t4386 VDD.n2226 1.4705
R31046 VDD.n2225 VDD.t3379 1.4705
R31047 VDD.t1992 VDD.n2225 1.4705
R31048 VDD.t1018 VDD.n7990 1.4705
R31049 VDD.n7990 VDD.t3792 1.4705
R31050 VDD.n7991 VDD.t2471 1.4705
R31051 VDD.n7991 VDD.t1018 1.4705
R31052 VDD.n7981 VDD.t3646 1.4705
R31053 VDD.n7981 VDD.t2471 1.4705
R31054 VDD.n7964 VDD.t1304 1.4705
R31055 VDD.t4132 VDD.n7964 1.4705
R31056 VDD.t1692 VDD.n2229 1.4705
R31057 VDD.n2229 VDD.t4480 1.4705
R31058 VDD.n2230 VDD.t3062 1.4705
R31059 VDD.n2230 VDD.t1692 1.4705
R31060 VDD.n2222 VDD.t4360 1.4705
R31061 VDD.n2222 VDD.t3062 1.4705
R31062 VDD.n7985 VDD.t2007 1.4705
R31063 VDD.t1106 VDD.n7985 1.4705
R31064 VDD.n7984 VDD.t3401 1.4705
R31065 VDD.t2007 VDD.n7984 1.4705
R31066 VDD.n7978 VDD.t2439 1.4705
R31067 VDD.t1429 VDD.n7978 1.4705
R31068 VDD.n7972 VDD.t1011 1.4705
R31069 VDD.n7972 VDD.t2439 1.4705
R31070 VDD.n7971 VDD.t1882 1.4705
R31071 VDD.t1011 VDD.n7971 1.4705
R31072 VDD.n6600 VDD.t2266 1.4705
R31073 VDD.n6600 VDD.t1304 1.4705
R31074 VDD.t3990 VDD.n6604 1.4705
R31075 VDD.n6604 VDD.t2266 1.4705
R31076 VDD.n6607 VDD.t1603 1.4705
R31077 VDD.n6607 VDD.t3480 1.4705
R31078 VDD.t3072 VDD.n6612 1.4705
R31079 VDD.n6612 VDD.t1603 1.4705
R31080 VDD.t3754 VDD.n6617 1.4705
R31081 VDD.n6617 VDD.t2564 1.4705
R31082 VDD.n6618 VDD.t999 1.4705
R31083 VDD.n6618 VDD.t3754 1.4705
R31084 VDD.t1865 VDD.n6622 1.4705
R31085 VDD.n6622 VDD.t999 1.4705
R31086 VDD.t3762 VDD.n5409 1.4705
R31087 VDD.n5409 VDD.t2460 1.4705
R31088 VDD.n5410 VDD.t4650 1.4705
R31089 VDD.n5410 VDD.t3762 1.4705
R31090 VDD.t2284 VDD.n5414 1.4705
R31091 VDD.n5414 VDD.t4650 1.4705
R31092 VDD.n5417 VDD.t4054 1.4705
R31093 VDD.n5417 VDD.t1702 1.4705
R31094 VDD.t1245 VDD.n5422 1.4705
R31095 VDD.n5422 VDD.t4054 1.4705
R31096 VDD.t2030 VDD.n5427 1.4705
R31097 VDD.n5427 VDD.t766 1.4705
R31098 VDD.n5428 VDD.t3417 1.4705
R31099 VDD.n5428 VDD.t2030 1.4705
R31100 VDD.t4302 VDD.n5432 1.4705
R31101 VDD.n5432 VDD.t3417 1.4705
R31102 VDD.n5406 VDD.t2750 1.4705
R31103 VDD.n5406 VDD.t1258 1.4705
R31104 VDD.n5404 VDD.t3575 1.4705
R31105 VDD.t2750 VDD.n5404 1.4705
R31106 VDD.n5403 VDD.t1134 1.4705
R31107 VDD.t3575 VDD.n5403 1.4705
R31108 VDD.n5400 VDD.t3026 1.4705
R31109 VDD.t601 VDD.n5400 1.4705
R31110 VDD.n5399 VDD.t4318 1.4705
R31111 VDD.t3026 VDD.n5399 1.4705
R31112 VDD.n5397 VDD.t947 1.4705
R31113 VDD.t3808 VDD.n5397 1.4705
R31114 VDD.n5395 VDD.t2370 1.4705
R31115 VDD.t947 VDD.n5395 1.4705
R31116 VDD.n5394 VDD.t3262 1.4705
R31117 VDD.t2370 VDD.n5394 1.4705
R31118 VDD.n7171 VDD.t3644 1.4705
R31119 VDD.t2833 VDD.n7171 1.4705
R31120 VDD.n7166 VDD.t908 1.4705
R31121 VDD.n7166 VDD.t3644 1.4705
R31122 VDD.n7165 VDD.t3652 1.4705
R31123 VDD.t908 VDD.n7165 1.4705
R31124 VDD.n7160 VDD.t4398 1.4705
R31125 VDD.t2760 VDD.n7160 1.4705
R31126 VDD.n7155 VDD.t1620 1.4705
R31127 VDD.n7155 VDD.t4398 1.4705
R31128 VDD.n7152 VDD.t3454 1.4705
R31129 VDD.t2074 VDD.n7152 1.4705
R31130 VDD.n7147 VDD.t641 1.4705
R31131 VDD.n7147 VDD.t3454 1.4705
R31132 VDD.n7146 VDD.t1915 1.4705
R31133 VDD.t641 VDD.n7146 1.4705
R31134 VDD.n7169 VDD.t2642 1.4705
R31135 VDD.n7169 VDD.t1634 1.4705
R31136 VDD.n7168 VDD.t3950 1.4705
R31137 VDD.t2642 VDD.n7168 1.4705
R31138 VDD.n7163 VDD.t2654 1.4705
R31139 VDD.n7163 VDD.t3950 1.4705
R31140 VDD.n7158 VDD.t3332 1.4705
R31141 VDD.n7158 VDD.t1547 1.4705
R31142 VDD.n7157 VDD.t4688 1.4705
R31143 VDD.t3332 VDD.n7157 1.4705
R31144 VDD.n7150 VDD.t2412 1.4705
R31145 VDD.n7150 VDD.t986 1.4705
R31146 VDD.n7149 VDD.t3713 1.4705
R31147 VDD.t2412 VDD.n7149 1.4705
R31148 VDD.n7144 VDD.t848 1.4705
R31149 VDD.n7144 VDD.t3713 1.4705
R31150 VDD.t1202 VDD.n7846 1.4705
R31151 VDD.n7846 VDD.t4466 1.4705
R31152 VDD.n7948 VDD.t43 1.4705
R31153 VDD.n7948 VDD.t35 1.4705
R31154 VDD.n7950 VDD.t33 1.4705
R31155 VDD.n7950 VDD.t26 1.4705
R31156 VDD.n7953 VDD.t207 1.4705
R31157 VDD.n7953 VDD.t278 1.4705
R31158 VDD.n7955 VDD.t19 1.4705
R31159 VDD.n7955 VDD.t41 1.4705
R31160 VDD.n7957 VDD.t13 1.4705
R31161 VDD.n7957 VDD.t39 1.4705
R31162 VDD.n7938 VDD.t160 1.4705
R31163 VDD.n7938 VDD.t235 1.4705
R31164 VDD.n7933 VDD.t240 1.4705
R31165 VDD.n7933 VDD.t88 1.4705
R31166 VDD.n7928 VDD.t149 1.4705
R31167 VDD.n7928 VDD.t194 1.4705
R31168 VDD.n7919 VDD.t128 1.4705
R31169 VDD.n7919 VDD.t175 1.4705
R31170 VDD.n7914 VDD.t153 1.4705
R31171 VDD.n7914 VDD.t202 1.4705
R31172 VDD.n7884 VDD.t256 1.4705
R31173 VDD.n7884 VDD.t98 1.4705
R31174 VDD.n7886 VDD.t87 1.4705
R31175 VDD.n7886 VDD.t165 1.4705
R31176 VDD.n7880 VDD.t109 1.4705
R31177 VDD.n7880 VDD.t185 1.4705
R31178 VDD.n7882 VDD.t172 1.4705
R31179 VDD.n7882 VDD.t248 1.4705
R31180 VDD.n7876 VDD.t24 1.4705
R31181 VDD.n7876 VDD.t15 1.4705
R31182 VDD.n7878 VDD.t42 1.4705
R31183 VDD.n7878 VDD.t36 1.4705
R31184 VDD.n7870 VDD.t221 1.4705
R31185 VDD.n7870 VDD.t266 1.4705
R31186 VDD.n7872 VDD.t277 1.4705
R31187 VDD.n7872 VDD.t102 1.4705
R31188 VDD.n7866 VDD.t242 1.4705
R31189 VDD.n7866 VDD.t46 1.4705
R31190 VDD.n7868 VDD.t72 1.4705
R31191 VDD.n7868 VDD.t131 1.4705
R31192 VDD.n8053 VDD.t171 1.4705
R31193 VDD.n8053 VDD.t246 1.4705
R31194 VDD.n8055 VDD.t257 1.4705
R31195 VDD.n8055 VDD.t99 1.4705
R31196 VDD.n8058 VDD.t75 1.4705
R31197 VDD.n8058 VDD.t156 1.4705
R31198 VDD.n8060 VDD.t140 1.4705
R31199 VDD.n8060 VDD.t186 1.4705
R31200 VDD.n8062 VDD.t163 1.4705
R31201 VDD.n8062 VDD.t214 1.4705
R31202 VDD.n8043 VDD.t21 1.4705
R31203 VDD.n8043 VDD.t40 1.4705
R31204 VDD.n8038 VDD.t37 1.4705
R31205 VDD.n8038 VDD.t30 1.4705
R31206 VDD.n8033 VDD.t241 1.4705
R31207 VDD.n8033 VDD.t45 1.4705
R31208 VDD.n8024 VDD.t29 1.4705
R31209 VDD.n8024 VDD.t17 1.4705
R31210 VDD.n8019 VDD.t22 1.4705
R31211 VDD.n8019 VDD.t44 1.4705
R31212 VDD.t4108 VDD.n2176 1.4705
R31213 VDD.n2176 VDD.t2802 1.4705
R31214 VDD.n2177 VDD.t1186 1.4705
R31215 VDD.n2177 VDD.t4108 1.4705
R31216 VDD.t2670 VDD.n2181 1.4705
R31217 VDD.n2181 VDD.t1186 1.4705
R31218 VDD.n2184 VDD.t4374 1.4705
R31219 VDD.n2184 VDD.t3494 1.4705
R31220 VDD.t1585 VDD.n7999 1.4705
R31221 VDD.n7999 VDD.t4374 1.4705
R31222 VDD.t4728 VDD.n8004 1.4705
R31223 VDD.n8004 VDD.t3834 1.4705
R31224 VDD.n8005 VDD.t3377 1.4705
R31225 VDD.n8005 VDD.t4728 1.4705
R31226 VDD.t4276 VDD.n8009 1.4705
R31227 VDD.n8009 VDD.t3377 1.4705
R31228 VDD.n6808 VDD.t238 1.4705
R31229 VDD.n6808 VDD.t280 1.4705
R31230 VDD.n6809 VDD.t181 1.4705
R31231 VDD.n6809 VDD.t227 1.4705
R31232 VDD.n6811 VDD.t236 1.4705
R31233 VDD.n6811 VDD.t161 1.4705
R31234 VDD.n6812 VDD.t180 1.4705
R31235 VDD.n6812 VDD.t103 1.4705
R31236 VDD.n6815 VDD.t249 1.4705
R31237 VDD.n6815 VDD.t92 1.4705
R31238 VDD.n6816 VDD.t190 1.4705
R31239 VDD.n6816 VDD.t265 1.4705
R31240 VDD.n6819 VDD.t101 1.4705
R31241 VDD.n6819 VDD.t173 1.4705
R31242 VDD.n6820 VDD.t271 1.4705
R31243 VDD.n6820 VDD.t114 1.4705
R31244 VDD.n6824 VDD.t231 1.4705
R31245 VDD.n6824 VDD.t71 1.4705
R31246 VDD.n6825 VDD.t174 1.4705
R31247 VDD.n6825 VDD.t251 1.4705
R31248 VDD.n6828 VDD.t81 1.4705
R31249 VDD.n6828 VDD.t183 1.4705
R31250 VDD.n6829 VDD.t258 1.4705
R31251 VDD.n6829 VDD.t126 1.4705
R31252 VDD.n6832 VDD.t93 1.4705
R31253 VDD.n6832 VDD.t167 1.4705
R31254 VDD.n6833 VDD.t267 1.4705
R31255 VDD.n6833 VDD.t110 1.4705
R31256 VDD.n6836 VDD.t203 1.4705
R31257 VDD.n6836 VDD.t252 1.4705
R31258 VDD.n6837 VDD.t147 1.4705
R31259 VDD.n6837 VDD.t192 1.4705
R31260 VDD.n6775 VDD.t145 1.4705
R31261 VDD.n6775 VDD.t189 1.4705
R31262 VDD.n6776 VDD.t245 1.4705
R31263 VDD.n6776 VDD.t56 1.4705
R31264 VDD.n6778 VDD.t144 1.4705
R31265 VDD.n6778 VDD.t52 1.4705
R31266 VDD.n6779 VDD.t244 1.4705
R31267 VDD.n6779 VDD.t169 1.4705
R31268 VDD.n6782 VDD.t155 1.4705
R31269 VDD.n6782 VDD.t228 1.4705
R31270 VDD.n6783 VDD.t259 1.4705
R31271 VDD.n6783 VDD.t104 1.4705
R31272 VDD.n6786 VDD.t237 1.4705
R31273 VDD.n6786 VDD.t67 1.4705
R31274 VDD.n6787 VDD.t111 1.4705
R31275 VDD.n6787 VDD.t184 1.4705
R31276 VDD.n6771 VDD.t139 1.4705
R31277 VDD.n6771 VDD.t215 1.4705
R31278 VDD.n6772 VDD.t239 1.4705
R31279 VDD.n6772 VDD.t86 1.4705
R31280 VDD.n6767 VDD.t222 1.4705
R31281 VDD.n6767 VDD.t84 1.4705
R31282 VDD.n6768 VDD.t91 1.4705
R31283 VDD.n6768 VDD.t188 1.4705
R31284 VDD.n6763 VDD.t232 1.4705
R31285 VDD.n6763 VDD.t61 1.4705
R31286 VDD.n6764 VDD.t107 1.4705
R31287 VDD.n6764 VDD.t178 1.4705
R31288 VDD.n6759 VDD.t105 1.4705
R31289 VDD.n6759 VDD.t157 1.4705
R31290 VDD.n6760 VDD.t209 1.4705
R31291 VDD.n6760 VDD.t260 1.4705
R31292 VDD.n6845 VDD.t94 1.4705
R31293 VDD.n6845 VDD.t176 1.4705
R31294 VDD.n6842 VDD.t118 1.4705
R31295 VDD.n6842 VDD.t196 1.4705
R31296 VDD.n6736 VDD.t158 1.4705
R31297 VDD.n6736 VDD.t255 1.4705
R31298 VDD.n6732 VDD.t179 1.4705
R31299 VDD.n6732 VDD.t65 1.4705
R31300 VDD.n6795 VDD.t233 1.4705
R31301 VDD.n6795 VDD.t74 1.4705
R31302 VDD.n6792 VDD.t254 1.4705
R31303 VDD.n6792 VDD.t97 1.4705
R31304 VDD.n9131 VDD.t3322 1.4705
R31305 VDD.n9131 VDD.t3518 1.4705
R31306 VDD.t2794 VDD.n9129 1.4705
R31307 VDD.n9129 VDD.t2999 1.4705
R31308 VDD.t4042 VDD.n9142 1.4705
R31309 VDD.n9142 VDD.t2547 1.4705
R31310 VDD.t3672 VDD.n9148 1.4705
R31311 VDD.n9148 VDD.t3898 1.4705
R31312 VDD.n9165 VDD.t4568 1.4705
R31313 VDD.t3102 VDD.n9165 1.4705
R31314 VDD.t4256 VDD.n8487 1.4705
R31315 VDD.n8487 VDD.t4460 1.4705
R31316 VDD.n8762 VDD.t3840 1.4705
R31317 VDD.t4060 VDD.n8762 1.4705
R31318 VDD.n8756 VDD.t3860 1.4705
R31319 VDD.t4516 VDD.n8756 1.4705
R31320 VDD.n8558 VDD.t2022 1.4705
R31321 VDD.t2252 VDD.n8558 1.4705
R31322 VDD.n8552 VDD.t2059 1.4705
R31323 VDD.t2813 VDD.n8552 1.4705
R31324 VDD.n8835 VDD.t2108 1.4705
R31325 VDD.t2869 VDD.n8835 1.4705
R31326 VDD.t2130 VDD.n8546 1.4705
R31327 VDD.n8546 VDD.t1032 1.4705
R31328 VDD.t3934 VDD.n8802 1.4705
R31329 VDD.n8802 VDD.t4584 1.4705
R31330 VDD.n8768 VDD.t3958 1.4705
R31331 VDD.t2941 VDD.n8768 1.4705
R31332 VDD.n8888 VDD.t3446 1.4705
R31333 VDD.t2520 VDD.n8888 1.4705
R31334 VDD.t3470 VDD.n8774 1.4705
R31335 VDD.n8774 VDD.t2437 1.4705
R31336 VDD.t1591 VDD.n8875 1.4705
R31337 VDD.n8875 VDD.t577 1.4705
R31338 VDD.n8841 VDD.t1618 1.4705
R31339 VDD.t4692 VDD.n8841 1.4705
R31340 VDD.n8944 VDD.t1676 1.4705
R31341 VDD.t2467 VDD.n8944 1.4705
R31342 VDD.t2210 VDD.n8847 1.4705
R31343 VDD.n8847 VDD.t596 1.4705
R31344 VDD.t3526 VDD.n8933 1.4705
R31345 VDD.n8933 VDD.t4226 1.4705
R31346 VDD.n8899 VDD.t4018 1.4705
R31347 VDD.t2528 VDD.n8899 1.4705
R31348 VDD.n9019 VDD.t4082 1.4705
R31349 VDD.t4290 VDD.n9019 1.4705
R31350 VDD.t4110 VDD.n8905 1.4705
R31351 VDD.n8905 VDD.t2624 1.4705
R31352 VDD.t2289 VDD.n9006 1.4705
R31353 VDD.n9006 VDD.t2560 1.4705
R31354 VDD.n8950 VDD.t2326 1.4705
R31355 VDD.t708 VDD.n8950 1.4705
R31356 VDD.n9041 VDD.t4486 1.4705
R31357 VDD.t3024 VDD.n9041 1.4705
R31358 VDD.t4178 VDD.n8974 1.4705
R31359 VDD.n8974 VDD.t4366 1.4705
R31360 VDD.t2190 VDD.n9030 1.4705
R31361 VDD.n9030 VDD.t561 1.4705
R31362 VDD.n9025 VDD.t1797 1.4705
R31363 VDD.t2062 VDD.n9025 1.4705
R31364 VDD.t2303 VDD.n9154 1.4705
R31365 VDD.n9154 VDD.t681 1.4705
R31366 VDD.n9072 VDD.t1894 1.4705
R31367 VDD.t2128 VDD.n9072 1.4705
R31368 VDD.n189 VDD.t2044 1.4705
R31369 VDD.t4604 VDD.n189 1.4705
R31370 VDD.n173 VDD.t4406 1.4705
R31371 VDD.t4630 VDD.n173 1.4705
R31372 VDD.n9122 VDD.t2229 1.4705
R31373 VDD.t623 VDD.n9122 1.4705
R31374 VDD.n9094 VDD.t1837 1.4705
R31375 VDD.t2089 VDD.n9094 1.4705
R31376 VDD.n1159 VDD.t4640 1.4705
R31377 VDD.t1678 VDD.n1159 1.4705
R31378 VDD.t738 VDD.n1747 1.4705
R31379 VDD.n1747 VDD.t4640 1.4705
R31380 VDD.n981 VDD.t464 1.4705
R31381 VDD.n981 VDD.t452 1.4705
R31382 VDD.n978 VDD.t438 1.4705
R31383 VDD.n978 VDD.t424 1.4705
R31384 VDD.n1714 VDD.t2943 1.4705
R31385 VDD.n1714 VDD.t3136 1.4705
R31386 VDD.n725 VDD.t2721 1.4705
R31387 VDD.t2943 VDD.n725 1.4705
R31388 VDD.t2719 VDD.n714 1.4705
R31389 VDD.t2939 VDD.n714 1.4705
R31390 VDD.n723 VDD.t2506 1.4705
R31391 VDD.n723 VDD.t2719 1.4705
R31392 VDD.n1738 VDD.t1288 1.4705
R31393 VDD.n1738 VDD.t1503 1.4705
R31394 VDD.t3816 VDD.n947 1.4705
R31395 VDD.n947 VDD.t1288 1.4705
R31396 VDD.n1035 VDD.t428 1.4705
R31397 VDD.n1035 VDD.t446 1.4705
R31398 VDD.n1037 VDD.t433 1.4705
R31399 VDD.n1037 VDD.t436 1.4705
R31400 VDD.n913 VDD.t4378 1.4705
R31401 VDD.t4582 VDD.n913 1.4705
R31402 VDD.n908 VDD.t2825 1.4705
R31403 VDD.n908 VDD.t4378 1.4705
R31404 VDD.n1068 VDD.t1745 1.4705
R31405 VDD.t1984 VDD.n1068 1.4705
R31406 VDD.n1063 VDD.t1526 1.4705
R31407 VDD.n1063 VDD.t1745 1.4705
R31408 VDD.n1042 VDD.t462 1.4705
R31409 VDD.n1042 VDD.t465 1.4705
R31410 VDD.n1040 VDD.t455 1.4705
R31411 VDD.n1040 VDD.t456 1.4705
R31412 VDD.n1491 VDD.t1907 1.4705
R31413 VDD.t736 VDD.n1491 1.4705
R31414 VDD.n1486 VDD.t1682 1.4705
R31415 VDD.n1486 VDD.t1907 1.4705
R31416 VDD.n1456 VDD.t4512 1.4705
R31417 VDD.t4738 VDD.n1456 1.4705
R31418 VDD.n1451 VDD.t1932 1.4705
R31419 VDD.n1451 VDD.t4512 1.4705
R31420 VDD.n1410 VDD.t3158 1.4705
R31421 VDD.n1410 VDD.t1508 1.4705
R31422 VDD.n1403 VDD.t1674 1.4705
R31423 VDD.t3158 VDD.n1403 1.4705
R31424 VDD.n1489 VDD.t1680 1.4705
R31425 VDD.n1489 VDD.t4654 1.4705
R31426 VDD.n1488 VDD.t1469 1.4705
R31427 VDD.t1680 VDD.n1488 1.4705
R31428 VDD.n1454 VDD.t4314 1.4705
R31429 VDD.n1454 VDD.t4510 1.4705
R31430 VDD.n1453 VDD.t1698 1.4705
R31431 VDD.t4314 VDD.n1453 1.4705
R31432 VDD.t2967 VDD.n1392 1.4705
R31433 VDD.t1295 VDD.n1392 1.4705
R31434 VDD.n1401 VDD.t1447 1.4705
R31435 VDD.n1401 VDD.t2967 1.4705
R31436 VDD.n1215 VDD.t3484 1.4705
R31437 VDD.t4670 VDD.n1215 1.4705
R31438 VDD.n1210 VDD.t3658 1.4705
R31439 VDD.n1210 VDD.t3484 1.4705
R31440 VDD.n1273 VDD.t1704 1.4705
R31441 VDD.n1273 VDD.t1844 1.4705
R31442 VDD.n1242 VDD.t4674 1.4705
R31443 VDD.t1704 VDD.n1242 1.4705
R31444 VDD.n1101 VDD.t364 1.4705
R31445 VDD.n1101 VDD.t331 1.4705
R31446 VDD.n1103 VDD.t362 1.4705
R31447 VDD.n1103 VDD.t343 1.4705
R31448 VDD.n1598 VDD.t3727 1.4705
R31449 VDD.n1598 VDD.t2185 1.4705
R31450 VDD.t783 VDD.n1603 1.4705
R31451 VDD.n1603 VDD.t3727 1.4705
R31452 VDD.n1501 VDD.t3522 1.4705
R31453 VDD.t1941 VDD.n1501 1.4705
R31454 VDD.n1500 VDD.t4696 1.4705
R31455 VDD.t3522 VDD.n1500 1.4705
R31456 VDD.n1623 VDD.t361 1.4705
R31457 VDD.n1623 VDD.t339 1.4705
R31458 VDD.n1621 VDD.t354 1.4705
R31459 VDD.n1621 VDD.t355 1.4705
R31460 VDD.n1527 VDD.t1870 1.4705
R31461 VDD.t1624 VDD.n1527 1.4705
R31462 VDD.n1516 VDD.t2429 1.4705
R31463 VDD.t693 VDD.n1516 1.4705
R31464 VDD.n1540 VDD.t1189 1.4705
R31465 VDD.t995 VDD.n1540 1.4705
R31466 VDD.t1666 VDD.n1562 1.4705
R31467 VDD.n1562 VDD.t4206 1.4705
R31468 VDD.n1172 VDD.t3003 1.4705
R31469 VDD.t4140 VDD.n1172 1.4705
R31470 VDD.n1167 VDD.t1684 1.4705
R31471 VDD.n1167 VDD.t3003 1.4705
R31472 VDD.n1185 VDD.t1988 1.4705
R31473 VDD.t1760 VDD.n1185 1.4705
R31474 VDD.n1180 VDD.t4566 1.4705
R31475 VDD.n1180 VDD.t1988 1.4705
R31476 VDD.n1089 VDD.t334 1.4705
R31477 VDD.n1089 VDD.t328 1.4705
R31478 VDD.n1087 VDD.t356 1.4705
R31479 VDD.n1087 VDD.t350 1.4705
R31480 VDD.n1420 VDD.t461 1.4705
R31481 VDD.n1420 VDD.t459 1.4705
R31482 VDD.n1422 VDD.t445 1.4705
R31483 VDD.n1422 VDD.t435 1.4705
R31484 VDD.n854 VDD.t426 1.4705
R31485 VDD.n854 VDD.t458 1.4705
R31486 VDD.n856 VDD.t443 1.4705
R31487 VDD.n856 VDD.t430 1.4705
R31488 VDD.n746 VDD.t365 1.4705
R31489 VDD.n746 VDD.t374 1.4705
R31490 VDD.n1675 VDD.t358 1.4705
R31491 VDD.n1675 VDD.t366 1.4705
R31492 VDD.n743 VDD.t368 1.4705
R31493 VDD.n743 VDD.t360 1.4705
R31494 VDD.n1681 VDD.t359 1.4705
R31495 VDD.n1681 VDD.t349 1.4705
R31496 VDD.n1340 VDD.t864 1.4705
R31497 VDD.n1340 VDD.t3798 1.4705
R31498 VDD.n1310 VDD.t589 1.4705
R31499 VDD.t864 VDD.n1310 1.4705
R31500 VDD.n1656 VDD.t2744 1.4705
R31501 VDD.t1089 VDD.n1656 1.4705
R31502 VDD.t3848 VDD.n1315 1.4705
R31503 VDD.n1315 VDD.t2744 1.4705
R31504 VDD.n740 VDD.t371 1.4705
R31505 VDD.n740 VDD.t346 1.4705
R31506 VDD.n1687 VDD.t344 1.4705
R31507 VDD.n1687 VDD.t491 1.4705
R31508 VDD.n1694 VDD.t453 1.4705
R31509 VDD.n1694 VDD.t467 1.4705
R31510 VDD.n737 VDD.t457 1.4705
R31511 VDD.n737 VDD.t437 1.4705
R31512 VDD.n1387 VDD.t2026 1.4705
R31513 VDD.n1387 VDD.t4592 1.4705
R31514 VDD.n1078 VDD.t579 1.4705
R31515 VDD.t2026 VDD.n1078 1.4705
R31516 VDD.n1283 VDD.t3478 1.4705
R31517 VDD.t3668 VDD.n1283 1.4705
R31518 VDD.t889 VDD.n1361 1.4705
R31519 VDD.n1361 VDD.t3478 1.4705
R31520 VDD.n1648 VDD.t3542 1.4705
R31521 VDD.n1648 VDD.t3342 1.4705
R31522 VDD.t3434 VDD.n1247 1.4705
R31523 VDD.n1247 VDD.t3542 1.4705
R31524 VDD.t1104 VDD.n694 1.4705
R31525 VDD.t1286 VDD.n694 1.4705
R31526 VDD.n945 VDD.t3599 1.4705
R31527 VDD.n945 VDD.t1104 1.4705
R31528 VDD.n6953 VDD.n6952 1.46537
R31529 VDD.n6957 VDD.n6956 1.46537
R31530 VDD.n6926 VDD.n6925 1.46537
R31531 VDD.n7011 VDD.n7010 1.46537
R31532 VDD.n7009 VDD.n7008 1.46537
R31533 VDD.n7004 VDD.n7003 1.46537
R31534 VDD.n6503 VDD.n6502 1.46537
R31535 VDD.n6501 VDD.n6500 1.46537
R31536 VDD.n6452 VDD.n6451 1.46537
R31537 VDD.n6543 VDD.n6542 1.46537
R31538 VDD.n6547 VDD.n6546 1.46537
R31539 VDD.n6541 VDD.n6540 1.46537
R31540 VDD.n6140 VDD.n6139 1.46537
R31541 VDD.n6144 VDD.n6143 1.46537
R31542 VDD.n6148 VDD.n6147 1.46537
R31543 VDD.n6133 VDD.n6132 1.46537
R31544 VDD.n6129 VDD.n6128 1.46537
R31545 VDD.n6125 VDD.n6124 1.46537
R31546 VDD.n6121 VDD.n6120 1.46537
R31547 VDD.n6048 VDD.n6047 1.46537
R31548 VDD.n6052 VDD.n6051 1.46537
R31549 VDD.n6056 VDD.n6055 1.46537
R31550 VDD.n6079 VDD.n6078 1.46537
R31551 VDD.n6083 VDD.n6082 1.46537
R31552 VDD.n6087 VDD.n6086 1.46537
R31553 VDD.n6091 VDD.n6090 1.46537
R31554 VDD.n6814 VDD.n6813 1.46537
R31555 VDD.n6818 VDD.n6817 1.46537
R31556 VDD.n6822 VDD.n6821 1.46537
R31557 VDD.n6827 VDD.n6826 1.46537
R31558 VDD.n6831 VDD.n6830 1.46537
R31559 VDD.n6835 VDD.n6834 1.46537
R31560 VDD.n6839 VDD.n6838 1.46537
R31561 VDD.n6781 VDD.n6780 1.46537
R31562 VDD.n6785 VDD.n6784 1.46537
R31563 VDD.n6789 VDD.n6788 1.46537
R31564 VDD.n6774 VDD.n6773 1.46537
R31565 VDD.n6770 VDD.n6769 1.46537
R31566 VDD.n6766 VDD.n6765 1.46537
R31567 VDD.n6762 VDD.n6761 1.46537
R31568 VDD.n6327 VDD.n5488 1.3379
R31569 VDD.n6013 VDD.n5488 1.3306
R31570 VDD.n7932 VDD.n7931 1.30325
R31571 VDD.n7897 VDD.n7896 1.30325
R31572 VDD.n8037 VDD.n8036 1.30325
R31573 VDD.n7951 VDD.n7949 1.27338
R31574 VDD.n7958 VDD.n7956 1.27338
R31575 VDD.n7954 VDD.n7952 1.27228
R31576 VDD.n8063 VDD.n8061 1.27228
R31577 VDD.n8059 VDD.n8057 1.27228
R31578 VDD.n8056 VDD.n8054 1.27228
R31579 VDD.n2383 VDD.n2381 1.27228
R31580 VDD.n7021 VDD.n7019 1.27228
R31581 VDD.n7017 VDD.n7015 1.27228
R31582 VDD.n6966 VDD.n6964 1.27228
R31583 VDD.n6974 VDD.n6972 1.27228
R31584 VDD.n6970 VDD.n6968 1.27228
R31585 VDD.n7011 VDD.n7009 1.27228
R31586 VDD.n6957 VDD.n6953 1.27228
R31587 VDD.n5296 VDD.n5294 1.27228
R31588 VDD.n6555 VDD.n6553 1.27228
R31589 VDD.n6559 VDD.n6557 1.27228
R31590 VDD.n6511 VDD.n6509 1.27228
R31591 VDD.n6516 VDD.n6514 1.27228
R31592 VDD.n6520 VDD.n6518 1.27228
R31593 VDD.n6547 VDD.n6543 1.27228
R31594 VDD.n6503 VDD.n6501 1.27228
R31595 VDD.n6125 VDD.n6121 1.27228
R31596 VDD.n6133 VDD.n6129 1.27228
R31597 VDD.n6148 VDD.n6144 1.27228
R31598 VDD.n6091 VDD.n6087 1.27228
R31599 VDD.n6083 VDD.n6079 1.27228
R31600 VDD.n6056 VDD.n6052 1.27228
R31601 VDD.n6155 VDD.n6153 1.27228
R31602 VDD.n6098 VDD.n6096 1.27228
R31603 VDD.n6839 VDD.n6835 1.27228
R31604 VDD.n6831 VDD.n6827 1.27228
R31605 VDD.n6822 VDD.n6818 1.27228
R31606 VDD.n6766 VDD.n6762 1.27228
R31607 VDD.n6774 VDD.n6770 1.27228
R31608 VDD.n6789 VDD.n6785 1.27228
R31609 VDD.n6844 VDD.n6843 1.27228
R31610 VDD.n6794 VDD.n6793 1.27228
R31611 VDD.n1511 VDD.t1664 1.27155
R31612 VDD.n1560 VDD.t4205 1.27155
R31613 VDD.n1538 VDD.t1187 1.27155
R31614 VDD.n1536 VDD.t993 1.27155
R31615 VDD.n1514 VDD.t2428 1.27155
R31616 VDD.n1513 VDD.t691 1.27155
R31617 VDD.n1525 VDD.t1869 1.27155
R31618 VDD.n1524 VDD.t1623 1.27155
R31619 VDD.n8089 VDD.n8088 1.26911
R31620 VDD.n1763 VDD.n1762 1.23698
R31621 VDD.n6327 VDD.n6326 1.14768
R31622 VDD.n6396 VDD.t413 1.1382
R31623 VDD.n6577 VDD.t409 1.1382
R31624 VDD.n7040 VDD.t96 1.1382
R31625 VDD.n7086 VDD.t73 1.1382
R31626 VDD.n7025 VDD.n7024 1.13692
R31627 VDD.n6414 VDD.n5297 1.13692
R31628 VDD.n6562 VDD.n6561 1.13692
R31629 VDD.n6877 VDD.n2384 1.13692
R31630 VDD.n12624 VDD.t834 1.00929
R31631 VDD.n12564 VDD.t1162 1.00929
R31632 VDD.n12568 VDD.t1766 1.00929
R31633 VDD.n12571 VDD.t1173 1.00929
R31634 VDD.n12575 VDD.t1536 1.00929
R31635 VDD.n12557 VDD.t3218 1.00929
R31636 VDD.n8624 VDD.t3124 1.00929
R31637 VDD.n8625 VDD.t3438 1.00929
R31638 VDD.n18 VDD.t4044 1.00929
R31639 VDD.n21 VDD.t3448 1.00929
R31640 VDD.n22 VDD.t3806 1.00929
R31641 VDD.n23 VDD.t1219 1.00929
R31642 VDD.n8631 VDD.t2995 1.00929
R31643 VDD.n8628 VDD.t3298 1.00929
R31644 VDD.n19 VDD.t3872 1.00929
R31645 VDD.n12607 VDD.t3308 1.00929
R31646 VDD.n12603 VDD.t3638 1.00929
R31647 VDD.n12600 VDD.t1087 1.00929
R31648 VDD.n8655 VDD.t3208 1.00929
R31649 VDD.n8656 VDD.t3508 1.00929
R31650 VDD.n27 VDD.t4134 1.00929
R31651 VDD.n12531 VDD.t3528 1.00929
R31652 VDD.n12536 VDD.t3892 1.00929
R31653 VDD.n12540 VDD.t1300 1.00929
R31654 VDD.n8662 VDD.t3064 1.00929
R31655 VDD.n8659 VDD.t3357 1.00929
R31656 VDD.n28 VDD.t3974 1.00929
R31657 VDD.n12532 VDD.t3373 1.00929
R31658 VDD.n12537 VDD.t3741 1.00929
R31659 VDD.n12541 VDD.t1156 1.00929
R31660 VDD.n8610 VDD.t3842 1.00929
R31661 VDD.n8611 VDD.t4212 1.00929
R31662 VDD.n37 VDD.t636 1.00929
R31663 VDD.n40 VDD.t4230 1.00929
R31664 VDD.n82 VDD.t4550 1.00929
R31665 VDD.n86 VDD.t2032 1.00929
R31666 VDD.n8617 VDD.t3468 1.00929
R31667 VDD.n8614 VDD.t3800 1.00929
R31668 VDD.n38 VDD.t4400 1.00929
R31669 VDD.n41 VDD.t3820 1.00929
R31670 VDD.n83 VDD.t4220 1.00929
R31671 VDD.n87 VDD.t1612 1.00929
R31672 VDD.n8688 VDD.t1425 1.00929
R31673 VDD.n8689 VDD.t1776 1.00929
R31674 VDD.n98 VDD.t2510 1.00929
R31675 VDD.n101 VDD.t1790 1.00929
R31676 VDD.n102 VDD.t2220 1.00929
R31677 VDD.n103 VDD.t3794 1.00929
R31678 VDD.n8695 VDD.t4166 1.00929
R31679 VDD.n8692 VDD.t4482 1.00929
R31680 VDD.n99 VDD.t984 1.00929
R31681 VDD.n12513 VDD.t4490 1.00929
R31682 VDD.n12509 VDD.t749 1.00929
R31683 VDD.n12506 VDD.t2408 1.00929
R31684 VDD.n8596 VDD.t1506 1.00929
R31685 VDD.n8597 VDD.t1874 1.00929
R31686 VDD.n107 VDD.t2598 1.00929
R31687 VDD.n12475 VDD.t1891 1.00929
R31688 VDD.n12480 VDD.t2347 1.00929
R31689 VDD.n12484 VDD.t3878 1.00929
R31690 VDD.n8603 VDD.t4246 1.00929
R31691 VDD.n8600 VDD.t4548 1.00929
R31692 VDD.n108 VDD.t1047 1.00929
R31693 VDD.n12476 VDD.t4574 1.00929
R31694 VDD.n12481 VDD.t829 1.00929
R31695 VDD.n12485 VDD.t2496 1.00929
R31696 VDD.n8726 VDD.t1053 1.00929
R31697 VDD.n8727 VDD.t1383 1.00929
R31698 VDD.n117 VDD.t2013 1.00929
R31699 VDD.n120 VDD.t1393 1.00929
R31700 VDD.n128 VDD.t1764 1.00929
R31701 VDD.n132 VDD.t3393 1.00929
R31702 VDD.n8733 VDD.t1822 1.00929
R31703 VDD.n8730 VDD.t2218 1.00929
R31704 VDD.n118 VDD.t2891 1.00929
R31705 VDD.n121 VDD.t2236 1.00929
R31706 VDD.n129 VDD.t2672 1.00929
R31707 VDD.n133 VDD.t4196 1.00929
R31708 VDD.n8583 VDD.t1128 1.00929
R31709 VDD.n8584 VDD.t1459 1.00929
R31710 VDD.n178 VDD.t2106 1.00929
R31711 VDD.n181 VDD.t1475 1.00929
R31712 VDD.n182 VDD.t1859 1.00929
R31713 VDD.n183 VDD.t3486 1.00929
R31714 VDD.n8590 VDD.t3826 1.00929
R31715 VDD.n8587 VDD.t4194 1.00929
R31716 VDD.n179 VDD.t611 1.00929
R31717 VDD.n12457 VDD.t4216 1.00929
R31718 VDD.n12453 VDD.t4534 1.00929
R31719 VDD.n12450 VDD.t2003 1.00929
R31720 VDD.n1765 VDD.t1670 1.00929
R31721 VDD.n11056 VDD.t1310 1.00929
R31722 VDD.n11076 VDD.t3882 1.00929
R31723 VDD.n11089 VDD.t1293 1.00929
R31724 VDD.n648 VDD.t966 1.00929
R31725 VDD.n641 VDD.t3942 1.00929
R31726 VDD.n5708 VDD.t2125 1.00929
R31727 VDD.n5709 VDD.t1739 1.00929
R31728 VDD.n1781 VDD.t4306 1.00929
R31729 VDD.n11008 VDD.t1729 1.00929
R31730 VDD.n11013 VDD.t1355 1.00929
R31731 VDD.n11017 VDD.t2068 1.00929
R31732 VDD.n5715 VDD.t4706 1.00929
R31733 VDD.n5712 VDD.t4358 1.00929
R31734 VDD.n1782 VDD.t2835 1.00929
R31735 VDD.n11009 VDD.t4348 1.00929
R31736 VDD.n11014 VDD.t3982 1.00929
R31737 VDD.n11018 VDD.t1420 1.00929
R31738 VDD.n5734 VDD.t1558 1.00929
R31739 VDD.n5735 VDD.t1200 1.00929
R31740 VDD.n1788 VDD.t3778 1.00929
R31741 VDD.n1791 VDD.t1191 1.00929
R31742 VDD.n1799 VDD.t853 1.00929
R31743 VDD.n1803 VDD.t2885 1.00929
R31744 VDD.n5741 VDD.t4190 1.00929
R31745 VDD.n5738 VDD.t3824 1.00929
R31746 VDD.n1789 VDD.t2234 1.00929
R31747 VDD.n1792 VDD.t3810 1.00929
R31748 VDD.n1800 VDD.t3450 1.00929
R31749 VDD.n1804 VDD.t2232 1.00929
R31750 VDD.n5695 VDD.t1138 1.00929
R31751 VDD.n5696 VDD.t804 1.00929
R31752 VDD.n1834 VDD.t3352 1.00929
R31753 VDD.n1837 VDD.t790 1.00929
R31754 VDD.n1838 VDD.t4530 1.00929
R31755 VDD.n1839 VDD.t3844 1.00929
R31756 VDD.n5702 VDD.t945 1.00929
R31757 VDD.n5699 VDD.t4712 1.00929
R31758 VDD.n1835 VDD.t3168 1.00929
R31759 VDD.n10991 VDD.t4698 1.00929
R31760 VDD.n10987 VDD.t4326 1.00929
R31761 VDD.n10984 VDD.t3140 1.00929
R31762 VDD.n5789 VDD.t3068 1.00929
R31763 VDD.n5790 VDD.t2727 1.00929
R31764 VDD.n1843 VDD.t1030 1.00929
R31765 VDD.n10953 VDD.t2705 1.00929
R31766 VDD.n10958 VDD.t2280 1.00929
R31767 VDD.n10962 VDD.t936 1.00929
R31768 VDD.n5796 VDD.t4642 1.00929
R31769 VDD.n5793 VDD.t4292 1.00929
R31770 VDD.n1844 VDD.t2778 1.00929
R31771 VDD.n10954 VDD.t4280 1.00929
R31772 VDD.n10959 VDD.t3910 1.00929
R31773 VDD.n10963 VDD.t4126 1.00929
R31774 VDD.n5682 VDD.t2540 1.00929
R31775 VDD.n5683 VDD.t2104 1.00929
R31776 VDD.n1853 VDD.t4628 1.00929
R31777 VDD.n1856 VDD.t2093 1.00929
R31778 VDD.n1882 VDD.t1686 1.00929
R31779 VDD.n1886 VDD.t1659 1.00929
R31780 VDD.n5689 VDD.t4130 1.00929
R31781 VDD.n5686 VDD.t3760 1.00929
R31782 VDD.n1854 VDD.t2153 1.00929
R31783 VDD.n1857 VDD.t3743 1.00929
R31784 VDD.n1883 VDD.t3375 1.00929
R31785 VDD.n1887 VDD.t698 1.00929
R31786 VDD.n5844 VDD.t856 1.00929
R31787 VDD.n5845 VDD.t4622 1.00929
R31788 VDD.n1899 VDD.t3094 1.00929
R31789 VDD.n1902 VDD.t4602 1.00929
R31790 VDD.n1903 VDD.t4254 1.00929
R31791 VDD.n1904 VDD.t2441 1.00929
R31792 VDD.n5851 VDD.t1768 1.00929
R31793 VDD.n5848 VDD.t1411 1.00929
R31794 VDD.n1900 VDD.t3992 1.00929
R31795 VDD.n10936 VDD.t1399 1.00929
R31796 VDD.n10932 VDD.t1050 1.00929
R31797 VDD.n10929 VDD.t1924 1.00929
R31798 VDD.n5669 VDD.t4444 1.00929
R31799 VDD.n5670 VDD.t4118 1.00929
R31800 VDD.n1908 VDD.t2571 1.00929
R31801 VDD.n10898 VDD.t4098 1.00929
R31802 VDD.n10903 VDD.t3703 1.00929
R31803 VDD.n10907 VDD.t3182 1.00929
R31804 VDD.n5676 VDD.t1945 1.00929
R31805 VDD.n5673 VDD.t1581 1.00929
R31806 VDD.n1909 VDD.t4160 1.00929
R31807 VDD.n10899 VDD.t1556 1.00929
R31808 VDD.n10904 VDD.t1184 1.00929
R31809 VDD.n10908 VDD.t2173 1.00929
R31810 VDD.n5877 VDD.t3922 1.00929
R31811 VDD.n5878 VDD.t3564 1.00929
R31812 VDD.n5879 VDD.t1937 1.00929
R31813 VDD.n5491 VDD.t3546 1.00929
R31814 VDD.n5496 VDD.t3224 1.00929
R31815 VDD.n5500 VDD.t3884 1.00929
R31816 VDD.n5898 VDD.t3796 1.00929
R31817 VDD.n5895 VDD.t3462 1.00929
R31818 VDD.n5891 VDD.t1800 1.00929
R31819 VDD.n5492 VDD.t3442 1.00929
R31820 VDD.n5497 VDD.t3112 1.00929
R31821 VDD.n5501 VDD.t3403 1.00929
R31822 VDD.n5627 VDD.t2849 1.00929
R31823 VDD.n5628 VDD.t2492 1.00929
R31824 VDD.n1926 VDD.t799 1.00929
R31825 VDD.n1929 VDD.t2483 1.00929
R31826 VDD.n1930 VDD.t2024 1.00929
R31827 VDD.n1931 VDD.t3216 1.00929
R31828 VDD.n5634 VDD.t3294 1.00929
R31829 VDD.n5631 VDD.t2987 1.00929
R31830 VDD.n1927 VDD.t1263 1.00929
R31831 VDD.n10881 VDD.t2965 1.00929
R31832 VDD.n10877 VDD.t2596 1.00929
R31833 VDD.n10874 VDD.t4168 1.00929
R31834 VDD.n5606 VDD.t826 1.00929
R31835 VDD.n5607 VDD.t4600 1.00929
R31836 VDD.n1935 VDD.t3080 1.00929
R31837 VDD.n10843 VDD.t4576 1.00929
R31838 VDD.n10848 VDD.t4240 1.00929
R31839 VDD.n10852 VDD.t814 1.00929
R31840 VDD.n5613 VDD.t4448 1.00929
R31841 VDD.n5610 VDD.t4122 1.00929
R31842 VDD.n1936 VDD.t2574 1.00929
R31843 VDD.n10844 VDD.t4100 1.00929
R31844 VDD.n10849 VDD.t3709 1.00929
R31845 VDD.n10853 VDD.t3320 1.00929
R31846 VDD.n5585 VDD.t2748 1.00929
R31847 VDD.n5586 VDD.t2374 1.00929
R31848 VDD.n1945 VDD.t675 1.00929
R31849 VDD.n1948 VDD.t2354 1.00929
R31850 VDD.n1974 VDD.t1896 1.00929
R31851 VDD.n1978 VDD.t2050 1.00929
R31852 VDD.n5592 VDD.t2149 1.00929
R31853 VDD.n5589 VDD.t1756 1.00929
R31854 VDD.n1946 VDD.t4322 1.00929
R31855 VDD.n1949 VDD.t1741 1.00929
R31856 VDD.n1975 VDD.t1371 1.00929
R31857 VDD.n1979 VDD.t4494 1.00929
R31858 VDD.n2106 VDD.t3864 1.00929
R31859 VDD.n2111 VDD.t3516 1.00929
R31860 VDD.n1991 VDD.t1876 1.00929
R31861 VDD.n1994 VDD.t3504 1.00929
R31862 VDD.n1995 VDD.t3174 1.00929
R31863 VDD.n1998 VDD.t1165 1.00929
R31864 VDD.n8096 VDD.t649 1.00929
R31865 VDD.n2114 VDD.t4456 1.00929
R31866 VDD.n1992 VDD.t2933 1.00929
R31867 VDD.n10826 VDD.t4430 1.00929
R31868 VDD.n10822 VDD.t4074 1.00929
R31869 VDD.n1999 VDD.t770 1.00929
R31870 VDD.n2093 VDD.t3334 1.00929
R31871 VDD.n2094 VDD.t3042 1.00929
R31872 VDD.n2008 VDD.t1323 1.00929
R31873 VDD.n10785 VDD.t3028 1.00929
R31874 VDD.n10790 VDD.t2662 1.00929
R31875 VDD.n10794 VDD.t1926 1.00929
R31876 VDD.n2100 VDD.t3256 1.00929
R31877 VDD.n2097 VDD.t2927 1.00929
R31878 VDD.n2009 VDD.t1207 1.00929
R31879 VDD.n10786 VDD.t2907 1.00929
R31880 VDD.n10791 VDD.t2538 1.00929
R31881 VDD.n10795 VDD.t1413 1.00929
R31882 VDD.n8122 VDD.t1013 1.00929
R31883 VDD.n8123 VDD.t633 1.00929
R31884 VDD.n2018 VDD.t3250 1.00929
R31885 VDD.n2021 VDD.t599 1.00929
R31886 VDD.n2029 VDD.t4394 1.00929
R31887 VDD.n2033 VDD.t3222 1.00929
R31888 VDD.n8129 VDD.t2752 1.00929
R31889 VDD.n8126 VDD.t2380 1.00929
R31890 VDD.n2019 VDD.t678 1.00929
R31891 VDD.n2022 VDD.t2360 1.00929
R31892 VDD.n2030 VDD.t1898 1.00929
R31893 VDD.n2034 VDD.t2226 1.00929
R31894 VDD.n8166 VDD.t2121 1.00929
R31895 VDD.n8181 VDD.t1733 1.00929
R31896 VDD.n8201 VDD.t4304 1.00929
R31897 VDD.n8214 VDD.t1719 1.00929
R31898 VDD.n8236 VDD.t1350 1.00929
R31899 VDD.n8249 VDD.t3036 1.00929
R31900 VDD.n9088 VDD.t3134 1.00929
R31901 VDD.n9089 VDD.t4646 1.00929
R31902 VDD.n9086 VDD.t2400 1.00929
R31903 VDD.n9087 VDD.t2766 1.00929
R31904 VDD.n9075 VDD.t3695 1.00929
R31905 VDD.n9076 VDD.t4062 1.00929
R31906 VDD.n8463 VDD.t4656 1.00929
R31907 VDD.n8467 VDD.t4076 1.00929
R31908 VDD.n8468 VDD.t4434 1.00929
R31909 VDD.n8469 VDD.t1868 1.00929
R31910 VDD.n9082 VDD.t2255 1.00929
R31911 VDD.n9079 VDD.t2674 1.00929
R31912 VDD.n8464 VDD.t3260 1.00929
R31913 VDD.n9175 VDD.t2685 1.00929
R31914 VDD.n9171 VDD.t3054 1.00929
R31915 VDD.n9168 VDD.t4540 1.00929
R31916 VDD.n8532 VDD.t1196 1.00929
R31917 VDD.n8533 VDD.t1538 1.00929
R31918 VDD.n8534 VDD.t2208 1.00929
R31919 VDD.n8540 VDD.t1562 1.00929
R31920 VDD.n8541 VDD.t1964 1.00929
R31921 VDD.n8542 VDD.t3558 1.00929
R31922 VDD.n8578 VDD.t1409 1.00929
R31923 VDD.n8575 VDD.t1762 1.00929
R31924 VDD.n8571 VDD.t2490 1.00929
R31925 VDD.n8568 VDD.t1778 1.00929
R31926 VDD.n8564 VDD.t2202 1.00929
R31927 VDD.n8561 VDD.t3782 1.00929
R31928 VDD.n8776 VDD.t3164 1.00929
R31929 VDD.n8777 VDD.t3476 1.00929
R31930 VDD.n8778 VDD.t4084 1.00929
R31931 VDD.n8779 VDD.t3496 1.00929
R31932 VDD.n8780 VDD.t3854 1.00929
R31933 VDD.n8522 VDD.t1266 1.00929
R31934 VDD.n8796 VDD.t1490 1.00929
R31935 VDD.n8793 VDD.t1857 1.00929
R31936 VDD.n8789 VDD.t2578 1.00929
R31937 VDD.n8786 VDD.t1878 1.00929
R31938 VDD.n8782 VDD.t2317 1.00929
R31939 VDD.n8523 VDD.t3866 1.00929
R31940 VDD.n8514 VDD.t3650 1.00929
R31941 VDD.n8850 VDD.t4032 1.00929
R31942 VDD.n8855 VDD.t4612 1.00929
R31943 VDD.n8859 VDD.t4046 1.00929
R31944 VDD.n8864 VDD.t4388 1.00929
R31945 VDD.n8868 VDD.t1819 1.00929
R31946 VDD.n8515 VDD.t2100 1.00929
R31947 VDD.n8851 VDD.t2532 1.00929
R31948 VDD.n8856 VDD.t3130 1.00929
R31949 VDD.n8860 VDD.t2551 1.00929
R31950 VDD.n8865 VDD.t2919 1.00929
R31951 VDD.n8869 VDD.t4416 1.00929
R31952 VDD.n8907 VDD.t1252 1.00929
R31953 VDD.n8908 VDD.t1607 1.00929
R31954 VDD.n8909 VDD.t2268 1.00929
R31955 VDD.n8910 VDD.t1626 1.00929
R31956 VDD.n8911 VDD.t2019 1.00929
R31957 VDD.n8503 VDD.t3611 1.00929
R31958 VDD.n8927 VDD.t3868 1.00929
R31959 VDD.n8924 VDD.t4236 1.00929
R31960 VDD.n8920 VDD.t668 1.00929
R31961 VDD.n8917 VDD.t4248 1.00929
R31962 VDD.n8913 VDD.t4590 1.00929
R31963 VDD.n8504 VDD.t2064 1.00929
R31964 VDD.n8495 VDD.t1825 1.00929
R31965 VDD.n8977 VDD.t2222 1.00929
R31966 VDD.n8982 VDD.t2893 1.00929
R31967 VDD.n8986 VDD.t2238 1.00929
R31968 VDD.n8991 VDD.t2676 1.00929
R31969 VDD.n8995 VDD.t4202 1.00929
R31970 VDD.n8496 VDD.t2732 1.00929
R31971 VDD.n8978 VDD.t3070 1.00929
R31972 VDD.n8983 VDD.t3616 1.00929
R31973 VDD.n8987 VDD.t3084 1.00929
R31974 VDD.n8992 VDD.t3407 1.00929
R31975 VDD.n8996 VDD.t837 1.00929
R31976 VDD.n8477 VDD.t1918 1.00929
R31977 VDD.n8478 VDD.t2352 1.00929
R31978 VDD.n8479 VDD.t2989 1.00929
R31979 VDD.n8481 VDD.t2372 1.00929
R31980 VDD.n8482 VDD.t2768 1.00929
R31981 VDD.n8483 VDD.t4270 1.00929
R31982 VDD.n9061 VDD.t2161 1.00929
R31983 VDD.n9058 VDD.t2588 1.00929
R31984 VDD.n9054 VDD.t3178 1.00929
R31985 VDD.n9051 VDD.t2610 1.00929
R31986 VDD.n9047 VDD.t2985 1.00929
R31987 VDD.n9044 VDD.t4472 1.00929
R31988 VDD.n12624 VDD.t1482 1.00871
R31989 VDD.n12564 VDD.t1848 1.00871
R31990 VDD.n12568 VDD.t2562 1.00871
R31991 VDD.n12571 VDD.t1861 1.00871
R31992 VDD.n12575 VDD.t2295 1.00871
R31993 VDD.n12557 VDD.t3852 1.00871
R31994 VDD.n8624 VDD.t1571 1.00871
R31995 VDD.n8625 VDD.t1939 1.00871
R31996 VDD.n18 VDD.t2652 1.00871
R31997 VDD.n21 VDD.t1966 1.00871
R31998 VDD.n22 VDD.t2414 1.00871
R31999 VDD.n23 VDD.t3944 1.00871
R32000 VDD.n8631 VDD.t1781 1.00871
R32001 VDD.n8628 VDD.t2181 1.00871
R32002 VDD.n19 VDD.t2863 1.00871
R32003 VDD.n12607 VDD.t2204 1.00871
R32004 VDD.n12603 VDD.t2644 1.00871
R32005 VDD.n12600 VDD.t4172 1.00871
R32006 VDD.n8655 VDD.t3371 1.00871
R32007 VDD.n8656 VDD.t3719 1.00871
R32008 VDD.n27 VDD.t4328 1.00871
R32009 VDD.n12531 VDD.t3735 1.00871
R32010 VDD.n12536 VDD.t4128 1.00871
R32011 VDD.n12540 VDD.t1516 1.00871
R32012 VDD.n8662 VDD.t1885 1.00871
R32013 VDD.n8659 VDD.t2286 1.00871
R32014 VDD.n28 VDD.t2959 1.00871
R32015 VDD.n12532 VDD.t2319 1.00871
R32016 VDD.n12537 VDD.t2738 1.00871
R32017 VDD.n12541 VDD.t4252 1.00871
R32018 VDD.n8610 VDD.t4064 1.00871
R32019 VDD.n8611 VDD.t4390 1.00871
R32020 VDD.n37 VDD.t891 1.00871
R32021 VDD.n40 VDD.t4404 1.00871
R32022 VDD.n82 VDD.t626 1.00871
R32023 VDD.n86 VDD.t2264 1.00871
R32024 VDD.n8617 VDD.t687 1.00871
R32025 VDD.n8614 VDD.t1057 1.00871
R32026 VDD.n38 VDD.t1649 1.00871
R32027 VDD.n41 VDD.t1075 1.00871
R32028 VDD.n83 VDD.t1415 1.00871
R32029 VDD.n87 VDD.t3104 1.00871
R32030 VDD.n8688 VDD.t1654 1.00871
R32031 VDD.n8689 VDD.t2034 1.00871
R32032 VDD.n98 VDD.t2723 1.00871
R32033 VDD.n101 VDD.t2054 1.00871
R32034 VDD.n102 VDD.t2500 1.00871
R32035 VDD.n103 VDD.t4016 1.00871
R32036 VDD.n8695 VDD.t4354 1.00871
R32037 VDD.n8692 VDD.t4704 1.00871
R32038 VDD.n99 VDD.t1153 1.00871
R32039 VDD.n12513 VDD.t4722 1.00871
R32040 VDD.n12509 VDD.t977 1.00871
R32041 VDD.n12506 VDD.t2634 1.00871
R32042 VDD.n8596 VDD.t4148 1.00871
R32043 VDD.n8597 VDD.t4470 1.00871
R32044 VDD.n107 VDD.t968 1.00871
R32045 VDD.n12475 VDD.t4484 1.00871
R32046 VDD.n12480 VDD.t726 1.00871
R32047 VDD.n12484 VDD.t2385 1.00871
R32048 VDD.n8603 VDD.t4440 1.00871
R32049 VDD.n8600 VDD.t620 1.00871
R32050 VDD.n108 VDD.t1233 1.00871
R32051 VDD.n12476 VDD.t651 1.00871
R32052 VDD.n12481 VDD.t1036 1.00871
R32053 VDD.n12485 VDD.t2713 1.00871
R32054 VDD.n8726 VDD.t3630 1.00871
R32055 VDD.n8727 VDD.t4008 1.00871
R32056 VDD.n117 VDD.t4586 1.00871
R32057 VDD.n120 VDD.t4030 1.00871
R32058 VDD.n128 VDD.t4376 1.00871
R32059 VDD.n132 VDD.t1788 1.00871
R32060 VDD.n8733 VDD.t2077 1.00871
R32061 VDD.n8730 VDD.t2494 1.00871
R32062 VDD.n118 VDD.t3096 1.00871
R32063 VDD.n121 VDD.t2514 1.00871
R32064 VDD.n129 VDD.t2879 1.00871
R32065 VDD.n133 VDD.t4382 1.00871
R32066 VDD.n8583 VDD.t4218 1.00871
R32067 VDD.n8584 VDD.t4524 1.00871
R32068 VDD.n178 VDD.t1020 1.00871
R32069 VDD.n181 VDD.t4532 1.00871
R32070 VDD.n182 VDD.t793 1.00871
R32071 VDD.n183 VDD.t2454 1.00871
R32072 VDD.n8590 VDD.t2715 1.00871
R32073 VDD.n8587 VDD.t3058 1.00871
R32074 VDD.n179 VDD.t3601 1.00871
R32075 VDD.n12457 VDD.t3076 1.00871
R32076 VDD.n12453 VDD.t3385 1.00871
R32077 VDD.n12450 VDD.t824 1.00871
R32078 VDD.n1765 VDD.t3126 1.00871
R32079 VDD.n11056 VDD.t2798 1.00871
R32080 VDD.n11076 VDD.t1100 1.00871
R32081 VDD.n11089 VDD.t2790 1.00871
R32082 VDD.n648 VDD.t2391 1.00871
R32083 VDD.n641 VDD.t2042 1.00871
R32084 VDD.n5708 VDD.t2612 1.00871
R32085 VDD.n5709 VDD.t2183 1.00871
R32086 VDD.n1781 VDD.t4702 1.00871
R32087 VDD.n11008 VDD.t2167 1.00871
R32088 VDD.n11013 VDD.t1748 1.00871
R32089 VDD.n11017 VDD.t2867 1.00871
R32090 VDD.n5715 VDD.t2488 1.00871
R32091 VDD.n5712 VDD.t2066 1.00871
R32092 VDD.n1782 VDD.t4560 1.00871
R32093 VDD.n11009 VDD.t2046 1.00871
R32094 VDD.n11014 VDD.t1643 1.00871
R32095 VDD.n11018 VDD.t2362 1.00871
R32096 VDD.n5734 VDD.t4356 1.00871
R32097 VDD.n5735 VDD.t4020 1.00871
R32098 VDD.n1788 VDD.t2486 1.00871
R32099 VDD.n1791 VDD.t4002 1.00871
R32100 VDD.n1799 VDD.t3620 1.00871
R32101 VDD.n1803 VDD.t4034 1.00871
R32102 VDD.n5741 VDD.t1846 1.00871
R32103 VDD.n5738 VDD.t1479 1.00871
R32104 VDD.n1789 VDD.t4056 1.00871
R32105 VDD.n1792 VDD.t1471 1.00871
R32106 VDD.n1800 VDD.t1113 1.00871
R32107 VDD.n1804 VDD.t3114 1.00871
R32108 VDD.n5695 VDD.t3948 1.00871
R32109 VDD.n5696 VDD.t3585 1.00871
R32110 VDD.n1834 VDD.t1968 1.00871
R32111 VDD.n1837 VDD.t3566 1.00871
R32112 VDD.n1838 VDD.t3246 1.00871
R32113 VDD.n1839 VDD.t918 1.00871
R32114 VDD.n5702 VDD.t746 1.00871
R32115 VDD.n5699 VDD.t4508 1.00871
R32116 VDD.n1835 VDD.t3011 1.00871
R32117 VDD.n10991 VDD.t4496 1.00871
R32118 VDD.n10987 VDD.t4162 1.00871
R32119 VDD.n10984 VDD.t4606 1.00871
R32120 VDD.n5789 VDD.t1597 1.00871
R32121 VDD.n5790 VDD.t1235 1.00871
R32122 VDD.n1843 VDD.t3804 1.00871
R32123 VDD.n10953 VDD.t1227 1.00871
R32124 VDD.n10958 VDD.t894 1.00871
R32125 VDD.n10962 VDD.t2123 1.00871
R32126 VDD.n5796 VDD.t3306 1.00871
R32127 VDD.n5793 VDD.t3007 1.00871
R32128 VDD.n1844 VDD.t1282 1.00871
R32129 VDD.n10954 VDD.t2991 1.00871
R32130 VDD.n10959 VDD.t2618 1.00871
R32131 VDD.n10963 VDD.t1143 1.00871
R32132 VDD.n5682 VDD.t1518 1.00871
R32133 VDD.n5683 VDD.t1171 1.00871
R32134 VDD.n1853 VDD.t3737 1.00871
R32135 VDD.n1856 VDD.t1158 1.00871
R32136 VDD.n1882 VDD.t802 1.00871
R32137 VDD.n1886 VDD.t1437 1.00871
R32138 VDD.n5689 VDD.t2815 1.00871
R32139 VDD.n5686 VDD.t2456 1.00871
R32140 VDD.n1854 VDD.t781 1.00871
R32141 VDD.n1857 VDD.t2443 1.00871
R32142 VDD.n1883 VDD.t1982 1.00871
R32143 VDD.n1887 VDD.t1902 1.00871
R32144 VDD.n5844 VDD.t4104 1.00871
R32145 VDD.n5845 VDD.t3729 1.00871
R32146 VDD.n1899 VDD.t2119 1.00871
R32147 VDD.n1902 VDD.t3717 1.00871
R32148 VDD.n1903 VDD.t3340 1.00871
R32149 VDD.n1904 VDD.t2175 1.00871
R32150 VDD.n5851 VDD.t4538 1.00871
R32151 VDD.n5848 VDD.t4234 1.00871
R32152 VDD.n1900 VDD.t2681 1.00871
R32153 VDD.n10936 VDD.t4224 1.00871
R32154 VDD.n10932 VDD.t3830 1.00871
R32155 VDD.n10929 VDD.t3202 1.00871
R32156 VDD.n5669 VDD.t2138 1.00871
R32157 VDD.n5670 VDD.t1752 1.00871
R32158 VDD.n1908 VDD.t4320 1.00871
R32159 VDD.n10898 VDD.t1737 1.00871
R32160 VDD.n10903 VDD.t1366 1.00871
R32161 VDD.n10907 VDD.t3976 1.00871
R32162 VDD.n5676 VDD.t1601 1.00871
R32163 VDD.n5673 VDD.t1239 1.00871
R32164 VDD.n1909 VDD.t3814 1.00871
R32165 VDD.n10899 VDD.t1229 1.00871
R32166 VDD.n10904 VDD.t906 1.00871
R32167 VDD.n10908 VDD.t2356 1.00871
R32168 VDD.n5877 VDD.t1577 1.00871
R32169 VDD.n5878 VDD.t1223 1.00871
R32170 VDD.n5879 VDD.t3790 1.00871
R32171 VDD.n5491 VDD.t1198 1.00871
R32172 VDD.n5496 VDD.t876 1.00871
R32173 VDD.n5500 VDD.t4710 1.00871
R32174 VDD.n5898 VDD.t3940 1.00871
R32175 VDD.n5895 VDD.t3579 1.00871
R32176 VDD.n5891 VDD.t1958 1.00871
R32177 VDD.n5492 VDD.t3556 1.00871
R32178 VDD.n5497 VDD.t3240 1.00871
R32179 VDD.n5501 VDD.t2112 1.00871
R32180 VDD.n5627 VDD.t1028 1.00871
R32181 VDD.n5628 VDD.t659 1.00871
R32182 VDD.n1926 VDD.t3274 1.00871
R32183 VDD.n1929 VDD.t639 1.00871
R32184 VDD.n1930 VDD.t4412 1.00871
R32185 VDD.n1931 VDD.t4332 1.00871
R32186 VDD.n5634 VDD.t1974 1.00871
R32187 VDD.n5631 VDD.t1605 1.00871
R32188 VDD.n1927 VDD.t4186 1.00871
R32189 VDD.n10881 VDD.t1589 1.00871
R32190 VDD.n10877 VDD.t1210 1.00871
R32191 VDD.n10874 VDD.t3912 1.00871
R32192 VDD.n5606 VDD.t4624 1.00871
R32193 VDD.n5607 VDD.t4288 1.00871
R32194 VDD.n1935 VDD.t2758 1.00871
R32195 VDD.n10843 VDD.t4272 1.00871
R32196 VDD.n10848 VDD.t3896 1.00871
R32197 VDD.n10852 VDD.t956 1.00871
R32198 VDD.n5613 VDD.t2151 1.00871
R32199 VDD.n5610 VDD.t1758 1.00871
R32200 VDD.n1936 VDD.t4324 1.00871
R32201 VDD.n10844 VDD.t1743 1.00871
R32202 VDD.n10849 VDD.t1374 1.00871
R32203 VDD.n10853 VDD.t4144 1.00871
R32204 VDD.n5585 VDD.t2402 1.00871
R32205 VDD.n5586 VDD.t1970 1.00871
R32206 VDD.n1945 VDD.t4488 1.00871
R32207 VDD.n1948 VDD.t1943 1.00871
R32208 VDD.n1974 VDD.t1550 1.00871
R32209 VDD.n1978 VDD.t2179 1.00871
R32210 VDD.n5592 VDD.t3988 1.00871
R32211 VDD.n5589 VDD.t3624 1.00871
R32212 VDD.n1946 VDD.t2011 1.00871
R32213 VDD.n1949 VDD.t3609 1.00871
R32214 VDD.n1975 VDD.t3284 1.00871
R32215 VDD.n1979 VDD.t1181 1.00871
R32216 VDD.n2106 VDD.t2568 1.00871
R32217 VDD.n2111 VDD.t2134 1.00871
R32218 VDD.n1991 VDD.t4666 1.00871
R32219 VDD.n1994 VDD.t2114 1.00871
R32220 VDD.n1995 VDD.t1715 1.00871
R32221 VDD.n1998 VDD.t2469 1.00871
R32222 VDD.n8096 VDD.t3464 1.00871
R32223 VDD.n2114 VDD.t3154 1.00871
R32224 VDD.n1992 VDD.t1440 1.00871
R32225 VDD.n10826 VDD.t3132 1.00871
R32226 VDD.n10822 VDD.t2792 1.00871
R32227 VDD.n1999 VDD.t1955 1.00871
R32228 VDD.n2093 VDD.t1930 1.00871
R32229 VDD.n2094 VDD.t1564 1.00871
R32230 VDD.n2008 VDD.t4152 1.00871
R32231 VDD.n10785 VDD.t1543 1.00871
R32232 VDD.n10790 VDD.t1178 1.00871
R32233 VDD.n10794 VDD.t3204 1.00871
R32234 VDD.n2100 VDD.t1794 1.00871
R32235 VDD.n2097 VDD.t1433 1.00871
R32236 VDD.n2009 VDD.t4028 1.00871
R32237 VDD.n10786 VDD.t1422 1.00871
R32238 VDD.n10791 VDD.t1082 1.00871
R32239 VDD.n10795 VDD.t2742 1.00871
R32240 VDD.n8122 VDD.t4258 1.00871
R32241 VDD.n8123 VDD.t3902 1.00871
R32242 VDD.n2018 VDD.t2350 1.00871
R32243 VDD.n2021 VDD.t3880 1.00871
R32244 VDD.n2029 VDD.t3512 1.00871
R32245 VDD.n2033 VDD.t3038 1.00871
R32246 VDD.n8129 VDD.t1260 1.00871
R32247 VDD.n8126 VDD.t953 1.00871
R32248 VDD.n2019 VDD.t3488 1.00871
R32249 VDD.n2022 VDD.t931 1.00871
R32250 VDD.n2030 VDD.t4684 1.00871
R32251 VDD.n2034 VDD.t3426 1.00871
R32252 VDD.n8166 VDD.t756 1.00871
R32253 VDD.n8181 VDD.t4518 1.00871
R32254 VDD.n8201 VDD.t3020 1.00871
R32255 VDD.n8214 VDD.t4504 1.00871
R32256 VDD.n8236 VDD.t4174 1.00871
R32257 VDD.n8249 VDD.t4184 1.00871
R32258 VDD.n9088 VDD.t3314 1.00871
R32259 VDD.n9089 VDD.t721 1.00871
R32260 VDD.n9086 VDD.t2630 1.00871
R32261 VDD.n9087 VDD.t2977 1.00871
R32262 VDD.n9075 VDD.t2143 1.00871
R32263 VDD.n9076 VDD.t2580 1.00871
R32264 VDD.n8463 VDD.t3166 1.00871
R32265 VDD.n8467 VDD.t2600 1.00871
R32266 VDD.n8468 VDD.t2969 1.00871
R32267 VDD.n8469 VDD.t4464 1.00871
R32268 VDD.n9082 VDD.t2536 1.00871
R32269 VDD.n9079 VDD.t2881 1.00871
R32270 VDD.n8464 VDD.t3440 1.00871
R32271 VDD.n9175 VDD.t2903 1.00871
R32272 VDD.n9171 VDD.t3254 1.00871
R32273 VDD.n9168 VDD.t604 1.00871
R32274 VDD.n8532 VDD.t4282 1.00871
R32275 VDD.n8533 VDD.t4618 1.00871
R32276 VDD.n8534 VDD.t1095 1.00871
R32277 VDD.n8540 VDD.t4644 1.00871
R32278 VDD.n8541 VDD.t899 1.00871
R32279 VDD.n8542 VDD.t2549 1.00871
R32280 VDD.n8578 VDD.t2703 1.00871
R32281 VDD.n8575 VDD.t3048 1.00871
R32282 VDD.n8571 VDD.t3595 1.00871
R32283 VDD.n8568 VDD.t3066 1.00871
R32284 VDD.n8564 VDD.t3383 1.00871
R32285 VDD.n8561 VDD.t811 1.00871
R32286 VDD.n8776 VDD.t2465 1.00871
R32287 VDD.n8777 VDD.t2821 1.00871
R32288 VDD.n8778 VDD.t3361 1.00871
R32289 VDD.n8779 VDD.t2837 1.00871
R32290 VDD.n8780 VDD.t3186 1.00871
R32291 VDD.n8522 VDD.t4708 1.00871
R32292 VDD.n8796 VDD.t3236 1.00871
R32293 VDD.n8793 VDD.t3538 1.00871
R32294 VDD.n8789 VDD.t4170 1.00871
R32295 VDD.n8786 VDD.t3548 1.00871
R32296 VDD.n8782 VDD.t3936 1.00871
R32297 VDD.n8523 VDD.t1334 1.00871
R32298 VDD.n8514 VDD.t2553 1.00871
R32299 VDD.n8850 VDD.t2901 1.00871
R32300 VDD.n8855 VDD.t3460 1.00871
R32301 VDD.n8859 VDD.t2913 1.00871
R32302 VDD.n8864 VDD.t3276 1.00871
R32303 VDD.n8868 VDD.t631 1.00871
R32304 VDD.n8515 VDD.t1016 1.00871
R32305 VDD.n8851 VDD.t1331 1.00871
R32306 VDD.n8856 VDD.t1972 1.00871
R32307 VDD.n8860 VDD.t1352 1.00871
R32308 VDD.n8865 VDD.t1725 1.00871
R32309 VDD.n8869 VDD.t3348 1.00871
R32310 VDD.n8907 VDD.t4250 1.00871
R32311 VDD.n8908 VDD.t4556 1.00871
R32312 VDD.n8909 VDD.t1055 1.00871
R32313 VDD.n8910 VDD.t4580 1.00871
R32314 VDD.n8911 VDD.t843 1.00871
R32315 VDD.n8503 VDD.t2504 1.00871
R32316 VDD.n8927 VDD.t2855 1.00871
R32317 VDD.n8924 VDD.t3184 1.00871
R32318 VDD.n8920 VDD.t3745 1.00871
R32319 VDD.n8917 VDD.t3198 1.00871
R32320 VDD.n8913 VDD.t3530 1.00871
R32321 VDD.n8504 VDD.t980 1.00871
R32322 VDD.n8495 VDD.t2080 1.00871
R32323 VDD.n8977 VDD.t2502 1.00871
R32324 VDD.n8982 VDD.t3100 1.00871
R32325 VDD.n8986 VDD.t2516 1.00871
R32326 VDD.n8991 VDD.t2883 1.00871
R32327 VDD.n8995 VDD.t4384 1.00871
R32328 VDD.n8496 VDD.t2949 1.00871
R32329 VDD.n8978 VDD.t3272 1.00871
R32330 VDD.n8983 VDD.t3832 1.00871
R32331 VDD.n8987 VDD.t3280 1.00871
R32332 VDD.n8992 VDD.t3605 1.00871
R32333 VDD.n8996 VDD.t1043 1.00871
R32334 VDD.n8477 VDD.t2156 1.00871
R32335 VDD.n8478 VDD.t2586 1.00871
R32336 VDD.n8479 VDD.t3176 1.00871
R32337 VDD.n8481 VDD.t2608 1.00871
R32338 VDD.n8482 VDD.t2981 1.00871
R32339 VDD.n8483 VDD.t4468 1.00871
R32340 VDD.n9061 VDD.t2448 1.00871
R32341 VDD.n9058 VDD.t2808 1.00871
R32342 VDD.n9054 VDD.t3336 1.00871
R32343 VDD.n9051 VDD.t2823 1.00871
R32344 VDD.n9047 VDD.t3172 1.00871
R32345 VDD.n9044 VDD.t4694 1.00871
R32346 VDD.n6897 VDD.n6896 0.9995
R32347 VDD.n6984 VDD.n6983 0.9995
R32348 VDD.n6994 VDD.n6993 0.9995
R32349 VDD.n6916 VDD.n6915 0.9995
R32350 VDD.n6936 VDD.n6935 0.9995
R32351 VDD.n6946 VDD.n6945 0.9995
R32352 VDD.n6430 VDD.n6429 0.9995
R32353 VDD.n6532 VDD.n6531 0.9995
R32354 VDD.n6526 VDD.n6525 0.9995
R32355 VDD.n6467 VDD.n6466 0.9995
R32356 VDD.n6492 VDD.n6491 0.9995
R32357 VDD.n6486 VDD.n6485 0.9995
R32358 VDD.n7918 VDD.n7917 0.9995
R32359 VDD.n7927 VDD.n7926 0.9995
R32360 VDD.n7937 VDD.n7936 0.9995
R32361 VDD.n7906 VDD.n7905 0.9995
R32362 VDD.n7900 VDD.n7899 0.9995
R32363 VDD.n7894 VDD.n7893 0.9995
R32364 VDD.n8023 VDD.n8022 0.9995
R32365 VDD.n8032 VDD.n8031 0.9995
R32366 VDD.n8042 VDD.n8041 0.9995
R32367 VDD.n6105 VDD.n6104 0.991625
R32368 VDD.n6062 VDD.n6061 0.991625
R32369 VDD.n6804 VDD.n6803 0.991625
R32370 VDD.n6755 VDD.n6754 0.991625
R32371 VDD.n7024 VDD.n7023 0.983405
R32372 VDD.n7013 VDD.n6877 0.983405
R32373 VDD.n6550 VDD.n6414 0.983405
R32374 VDD.n6561 VDD.n6560 0.983405
R32375 VDD.n7952 VDD.n7951 0.937025
R32376 VDD.n8057 VDD.n8056 0.937025
R32377 VDD.n12633 VDD.n7 0.897031
R32378 VDD.n11872 VDD.n7 0.884663
R32379 VDD.n5539 VDD.n5538 0.851788
R32380 VDD.n6977 VDD.n6976 0.822966
R32381 VDD.n6999 VDD.n6878 0.822966
R32382 VDD.n6536 VDD.n6415 0.822966
R32383 VDD.n6522 VDD.n6521 0.822966
R32384 VDD.n65 VDD.n64 0.805721
R32385 VDD.n154 VDD.n153 0.805721
R32386 VDD.n9109 VDD.n9108 0.805721
R32387 VDD.n8822 VDD.n8821 0.805721
R32388 VDD.n8962 VDD.n8961 0.805721
R32389 VDD.n5765 VDD.n5764 0.805146
R32390 VDD.n5832 VDD.n5831 0.805146
R32391 VDD.n5649 VDD.n5648 0.805146
R32392 VDD.n5567 VDD.n5566 0.805146
R32393 VDD.n8153 VDD.n8152 0.805146
R32394 VDD.n69 VDD.n67 0.803395
R32395 VDD.n158 VDD.n156 0.803395
R32396 VDD.n9113 VDD.n9111 0.803395
R32397 VDD.n8826 VDD.n8824 0.803395
R32398 VDD.n8966 VDD.n8964 0.803395
R32399 VDD.n5768 VDD.n5767 0.80221
R32400 VDD.n5835 VDD.n5834 0.80221
R32401 VDD.n5652 VDD.n5651 0.80221
R32402 VDD.n5570 VDD.n5569 0.80221
R32403 VDD.n8156 VDD.n8155 0.80221
R32404 VDD.n8087 VDD.n8086 0.789456
R32405 VDD.n6156 VDD.n6019 0.737223
R32406 VDD.n6099 VDD.n6092 0.737223
R32407 VDD.n6151 VDD.n6150 0.737223
R32408 VDD.n6074 VDD.n6038 0.737223
R32409 VDD.n6848 VDD.n2405 0.737223
R32410 VDD.n6798 VDD.n6791 0.737223
R32411 VDD.n6841 VDD.n6840 0.737223
R32412 VDD.n6758 VDD.n6728 0.737223
R32413 VDD.n6100 VDD.n6099 0.725061
R32414 VDD.n6117 VDD.n6038 0.725061
R32415 VDD.n6799 VDD.n6798 0.725061
R32416 VDD.n6807 VDD.n6728 0.725061
R32417 VDD.n6328 VDD.n6327 0.699146
R32418 VDD.n6013 VDD.n5988 0.697565
R32419 VDD.n6299 VDD.n5488 0.694506
R32420 VDD.n7923 VDD.n7922 0.66425
R32421 VDD.n7903 VDD.n7902 0.66425
R32422 VDD.n8028 VDD.n8027 0.66425
R32423 VDD.n7023 VDD.n2376 0.639318
R32424 VDD.n6976 VDD.n6959 0.639318
R32425 VDD.n7013 VDD.n7012 0.639318
R32426 VDD.n6951 VDD.n6878 0.639318
R32427 VDD.n6550 VDD.n6549 0.639318
R32428 VDD.n6496 VDD.n6415 0.639318
R32429 VDD.n6560 VDD.n5289 0.639318
R32430 VDD.n6521 VDD.n6504 0.639318
R32431 VDD.n980 VDD.n979 0.636255
R32432 VDD.n1039 VDD.n1038 0.636255
R32433 VDD.n1041 VDD.n735 0.636255
R32434 VDD.n1102 VDD.n784 0.636255
R32435 VDD.n1625 VDD.n1624 0.636255
R32436 VDD.n1091 VDD.n1090 0.636255
R32437 VDD.n1424 VDD.n1423 0.636255
R32438 VDD.n858 VDD.n857 0.636255
R32439 VDD.n1674 VDD.n1673 0.636255
R32440 VDD.n1680 VDD.n1679 0.636255
R32441 VDD.n1686 VDD.n1685 0.636255
R32442 VDD.n1693 VDD.n1692 0.636255
R32443 VDD.n983 VDD.n982 0.63334
R32444 VDD.n1036 VDD.n1034 0.63334
R32445 VDD.n1044 VDD.n1043 0.63334
R32446 VDD.n1105 VDD.n1104 0.63334
R32447 VDD.n1622 VDD.n1620 0.63334
R32448 VDD.n1088 VDD.n1086 0.63334
R32449 VDD.n1421 VDD.n1419 0.63334
R32450 VDD.n855 VDD.n853 0.63334
R32451 VDD.n1677 VDD.n1676 0.63334
R32452 VDD.n1683 VDD.n1682 0.63334
R32453 VDD.n1689 VDD.n1688 0.63334
R32454 VDD.n1696 VDD.n1695 0.63334
R32455 VDD.n982 VDD.n980 0.631515
R32456 VDD.n1038 VDD.n1036 0.631515
R32457 VDD.n1043 VDD.n1041 0.631515
R32458 VDD.n1104 VDD.n1102 0.631515
R32459 VDD.n1624 VDD.n1622 0.631515
R32460 VDD.n1090 VDD.n1088 0.631515
R32461 VDD.n1423 VDD.n1421 0.631515
R32462 VDD.n857 VDD.n855 0.631515
R32463 VDD.n1676 VDD.n1674 0.631515
R32464 VDD.n1682 VDD.n1680 0.631515
R32465 VDD.n1688 VDD.n1686 0.631515
R32466 VDD.n1695 VDD.n1693 0.631515
R32467 VDD.n1742 VDD.t432 0.60727
R32468 VDD.t442 VDD.n1718 0.60727
R32469 VDD.t444 VDD.n1414 0.60727
R32470 VDD.n1356 VDD.t318 0.60727
R32471 VDD.n1349 VDD.t319 0.60727
R32472 VDD.n1652 VDD.t313 0.60727
R32473 VDD.n6977 VDD.n2376 0.585196
R32474 VDD.n7012 VDD.n6999 0.585196
R32475 VDD.n6549 VDD.n6536 0.585196
R32476 VDD.n6522 VDD.n5289 0.585196
R32477 VDD.n6100 VDD.n6019 0.585196
R32478 VDD.n6150 VDD.n6117 0.585196
R32479 VDD.n6799 VDD.n2405 0.585196
R32480 VDD.n6840 VDD.n6807 0.585196
R32481 VDD.n8087 VDD.n2119 0.51351
R32482 VDD.n5912 VDD.n5539 0.48482
R32483 VDD.n8250 VDD.n8249 0.468749
R32484 VDD.n8237 VDD.n8236 0.468749
R32485 VDD.n8215 VDD.n8214 0.468749
R32486 VDD.n8202 VDD.n8201 0.468749
R32487 VDD.n8182 VDD.n8181 0.468749
R32488 VDD.n8167 VDD.n8166 0.468749
R32489 VDD.n2035 VDD.n2034 0.468749
R32490 VDD.n2031 VDD.n2030 0.468749
R32491 VDD.n2023 VDD.n2022 0.468749
R32492 VDD.n2020 VDD.n2019 0.468749
R32493 VDD.n8127 VDD.n8126 0.468749
R32494 VDD.n8130 VDD.n8129 0.468749
R32495 VDD.n2035 VDD.n2033 0.468749
R32496 VDD.n2031 VDD.n2029 0.468749
R32497 VDD.n2023 VDD.n2021 0.468749
R32498 VDD.n2020 VDD.n2018 0.468749
R32499 VDD.n8127 VDD.n8123 0.468749
R32500 VDD.n8130 VDD.n8122 0.468749
R32501 VDD.n10796 VDD.n10795 0.468749
R32502 VDD.n10792 VDD.n10791 0.468749
R32503 VDD.n10787 VDD.n10786 0.468749
R32504 VDD.n2010 VDD.n2009 0.468749
R32505 VDD.n2098 VDD.n2097 0.468749
R32506 VDD.n2101 VDD.n2100 0.468749
R32507 VDD.n10796 VDD.n10794 0.468749
R32508 VDD.n10792 VDD.n10790 0.468749
R32509 VDD.n10787 VDD.n10785 0.468749
R32510 VDD.n2010 VDD.n2008 0.468749
R32511 VDD.n2098 VDD.n2094 0.468749
R32512 VDD.n2101 VDD.n2093 0.468749
R32513 VDD.n2000 VDD.n1999 0.468749
R32514 VDD.n10823 VDD.n10822 0.468749
R32515 VDD.n10827 VDD.n10826 0.468749
R32516 VDD.n1993 VDD.n1992 0.468749
R32517 VDD.n2115 VDD.n2114 0.468749
R32518 VDD.n8097 VDD.n8096 0.468749
R32519 VDD.n2000 VDD.n1998 0.468749
R32520 VDD.n10823 VDD.n1995 0.468749
R32521 VDD.n10827 VDD.n1994 0.468749
R32522 VDD.n1993 VDD.n1991 0.468749
R32523 VDD.n2115 VDD.n2111 0.468749
R32524 VDD.n8097 VDD.n2106 0.468749
R32525 VDD.n1980 VDD.n1979 0.468749
R32526 VDD.n1976 VDD.n1975 0.468749
R32527 VDD.n1950 VDD.n1949 0.468749
R32528 VDD.n1947 VDD.n1946 0.468749
R32529 VDD.n5590 VDD.n5589 0.468749
R32530 VDD.n5593 VDD.n5592 0.468749
R32531 VDD.n1980 VDD.n1978 0.468749
R32532 VDD.n1976 VDD.n1974 0.468749
R32533 VDD.n1950 VDD.n1948 0.468749
R32534 VDD.n1947 VDD.n1945 0.468749
R32535 VDD.n5590 VDD.n5586 0.468749
R32536 VDD.n5593 VDD.n5585 0.468749
R32537 VDD.n10854 VDD.n10853 0.468749
R32538 VDD.n10850 VDD.n10849 0.468749
R32539 VDD.n10845 VDD.n10844 0.468749
R32540 VDD.n1937 VDD.n1936 0.468749
R32541 VDD.n5611 VDD.n5610 0.468749
R32542 VDD.n5614 VDD.n5613 0.468749
R32543 VDD.n10854 VDD.n10852 0.468749
R32544 VDD.n10850 VDD.n10848 0.468749
R32545 VDD.n10845 VDD.n10843 0.468749
R32546 VDD.n1937 VDD.n1935 0.468749
R32547 VDD.n5611 VDD.n5607 0.468749
R32548 VDD.n5614 VDD.n5606 0.468749
R32549 VDD.n10875 VDD.n10874 0.468749
R32550 VDD.n10878 VDD.n10877 0.468749
R32551 VDD.n10882 VDD.n10881 0.468749
R32552 VDD.n1928 VDD.n1927 0.468749
R32553 VDD.n5632 VDD.n5631 0.468749
R32554 VDD.n5635 VDD.n5634 0.468749
R32555 VDD.n10875 VDD.n1931 0.468749
R32556 VDD.n10878 VDD.n1930 0.468749
R32557 VDD.n10882 VDD.n1929 0.468749
R32558 VDD.n1928 VDD.n1926 0.468749
R32559 VDD.n5632 VDD.n5628 0.468749
R32560 VDD.n5635 VDD.n5627 0.468749
R32561 VDD.n5502 VDD.n5501 0.468749
R32562 VDD.n5498 VDD.n5497 0.468749
R32563 VDD.n5493 VDD.n5492 0.468749
R32564 VDD.n5892 VDD.n5891 0.468749
R32565 VDD.n5896 VDD.n5895 0.468749
R32566 VDD.n5899 VDD.n5898 0.468749
R32567 VDD.n5502 VDD.n5500 0.468749
R32568 VDD.n5498 VDD.n5496 0.468749
R32569 VDD.n5493 VDD.n5491 0.468749
R32570 VDD.n5892 VDD.n5879 0.468749
R32571 VDD.n5896 VDD.n5878 0.468749
R32572 VDD.n5899 VDD.n5877 0.468749
R32573 VDD.n10909 VDD.n10908 0.468749
R32574 VDD.n10905 VDD.n10904 0.468749
R32575 VDD.n10900 VDD.n10899 0.468749
R32576 VDD.n1910 VDD.n1909 0.468749
R32577 VDD.n5674 VDD.n5673 0.468749
R32578 VDD.n5677 VDD.n5676 0.468749
R32579 VDD.n10909 VDD.n10907 0.468749
R32580 VDD.n10905 VDD.n10903 0.468749
R32581 VDD.n10900 VDD.n10898 0.468749
R32582 VDD.n1910 VDD.n1908 0.468749
R32583 VDD.n5674 VDD.n5670 0.468749
R32584 VDD.n5677 VDD.n5669 0.468749
R32585 VDD.n10930 VDD.n10929 0.468749
R32586 VDD.n10933 VDD.n10932 0.468749
R32587 VDD.n10937 VDD.n10936 0.468749
R32588 VDD.n1901 VDD.n1900 0.468749
R32589 VDD.n5849 VDD.n5848 0.468749
R32590 VDD.n5852 VDD.n5851 0.468749
R32591 VDD.n10930 VDD.n1904 0.468749
R32592 VDD.n10933 VDD.n1903 0.468749
R32593 VDD.n10937 VDD.n1902 0.468749
R32594 VDD.n1901 VDD.n1899 0.468749
R32595 VDD.n5849 VDD.n5845 0.468749
R32596 VDD.n5852 VDD.n5844 0.468749
R32597 VDD.n1888 VDD.n1887 0.468749
R32598 VDD.n1884 VDD.n1883 0.468749
R32599 VDD.n1858 VDD.n1857 0.468749
R32600 VDD.n1855 VDD.n1854 0.468749
R32601 VDD.n5687 VDD.n5686 0.468749
R32602 VDD.n5690 VDD.n5689 0.468749
R32603 VDD.n1888 VDD.n1886 0.468749
R32604 VDD.n1884 VDD.n1882 0.468749
R32605 VDD.n1858 VDD.n1856 0.468749
R32606 VDD.n1855 VDD.n1853 0.468749
R32607 VDD.n5687 VDD.n5683 0.468749
R32608 VDD.n5690 VDD.n5682 0.468749
R32609 VDD.n10964 VDD.n10963 0.468749
R32610 VDD.n10960 VDD.n10959 0.468749
R32611 VDD.n10955 VDD.n10954 0.468749
R32612 VDD.n1845 VDD.n1844 0.468749
R32613 VDD.n5794 VDD.n5793 0.468749
R32614 VDD.n5797 VDD.n5796 0.468749
R32615 VDD.n10964 VDD.n10962 0.468749
R32616 VDD.n10960 VDD.n10958 0.468749
R32617 VDD.n10955 VDD.n10953 0.468749
R32618 VDD.n1845 VDD.n1843 0.468749
R32619 VDD.n5794 VDD.n5790 0.468749
R32620 VDD.n5797 VDD.n5789 0.468749
R32621 VDD.n10985 VDD.n10984 0.468749
R32622 VDD.n10988 VDD.n10987 0.468749
R32623 VDD.n10992 VDD.n10991 0.468749
R32624 VDD.n1836 VDD.n1835 0.468749
R32625 VDD.n5700 VDD.n5699 0.468749
R32626 VDD.n5703 VDD.n5702 0.468749
R32627 VDD.n10985 VDD.n1839 0.468749
R32628 VDD.n10988 VDD.n1838 0.468749
R32629 VDD.n10992 VDD.n1837 0.468749
R32630 VDD.n1836 VDD.n1834 0.468749
R32631 VDD.n5700 VDD.n5696 0.468749
R32632 VDD.n5703 VDD.n5695 0.468749
R32633 VDD.n1805 VDD.n1804 0.468749
R32634 VDD.n1801 VDD.n1800 0.468749
R32635 VDD.n1793 VDD.n1792 0.468749
R32636 VDD.n1790 VDD.n1789 0.468749
R32637 VDD.n5739 VDD.n5738 0.468749
R32638 VDD.n5742 VDD.n5741 0.468749
R32639 VDD.n1805 VDD.n1803 0.468749
R32640 VDD.n1801 VDD.n1799 0.468749
R32641 VDD.n1793 VDD.n1791 0.468749
R32642 VDD.n1790 VDD.n1788 0.468749
R32643 VDD.n5739 VDD.n5735 0.468749
R32644 VDD.n5742 VDD.n5734 0.468749
R32645 VDD.n11019 VDD.n11018 0.468749
R32646 VDD.n11015 VDD.n11014 0.468749
R32647 VDD.n11010 VDD.n11009 0.468749
R32648 VDD.n1783 VDD.n1782 0.468749
R32649 VDD.n5713 VDD.n5712 0.468749
R32650 VDD.n5716 VDD.n5715 0.468749
R32651 VDD.n11019 VDD.n11017 0.468749
R32652 VDD.n11015 VDD.n11013 0.468749
R32653 VDD.n11010 VDD.n11008 0.468749
R32654 VDD.n1783 VDD.n1781 0.468749
R32655 VDD.n5713 VDD.n5709 0.468749
R32656 VDD.n5716 VDD.n5708 0.468749
R32657 VDD.n642 VDD.n641 0.468749
R32658 VDD.n649 VDD.n648 0.468749
R32659 VDD.n11090 VDD.n11089 0.468749
R32660 VDD.n11077 VDD.n11076 0.468749
R32661 VDD.n11057 VDD.n11056 0.468749
R32662 VDD.n1766 VDD.n1765 0.468749
R32663 VDD.n9045 VDD.n9044 0.468749
R32664 VDD.n9048 VDD.n9047 0.468749
R32665 VDD.n9052 VDD.n9051 0.468749
R32666 VDD.n9055 VDD.n9054 0.468749
R32667 VDD.n9059 VDD.n9058 0.468749
R32668 VDD.n9062 VDD.n9061 0.468749
R32669 VDD.n9045 VDD.n8483 0.468749
R32670 VDD.n9048 VDD.n8482 0.468749
R32671 VDD.n9052 VDD.n8481 0.468749
R32672 VDD.n9055 VDD.n8479 0.468749
R32673 VDD.n9059 VDD.n8478 0.468749
R32674 VDD.n9062 VDD.n8477 0.468749
R32675 VDD.n8997 VDD.n8996 0.468749
R32676 VDD.n8993 VDD.n8992 0.468749
R32677 VDD.n8988 VDD.n8987 0.468749
R32678 VDD.n8984 VDD.n8983 0.468749
R32679 VDD.n8979 VDD.n8978 0.468749
R32680 VDD.n8497 VDD.n8496 0.468749
R32681 VDD.n8997 VDD.n8995 0.468749
R32682 VDD.n8993 VDD.n8991 0.468749
R32683 VDD.n8988 VDD.n8986 0.468749
R32684 VDD.n8984 VDD.n8982 0.468749
R32685 VDD.n8979 VDD.n8977 0.468749
R32686 VDD.n8497 VDD.n8495 0.468749
R32687 VDD.n8505 VDD.n8504 0.468749
R32688 VDD.n8914 VDD.n8913 0.468749
R32689 VDD.n8918 VDD.n8917 0.468749
R32690 VDD.n8921 VDD.n8920 0.468749
R32691 VDD.n8925 VDD.n8924 0.468749
R32692 VDD.n8928 VDD.n8927 0.468749
R32693 VDD.n8505 VDD.n8503 0.468749
R32694 VDD.n8914 VDD.n8911 0.468749
R32695 VDD.n8918 VDD.n8910 0.468749
R32696 VDD.n8921 VDD.n8909 0.468749
R32697 VDD.n8925 VDD.n8908 0.468749
R32698 VDD.n8928 VDD.n8907 0.468749
R32699 VDD.n8870 VDD.n8869 0.468749
R32700 VDD.n8866 VDD.n8865 0.468749
R32701 VDD.n8861 VDD.n8860 0.468749
R32702 VDD.n8857 VDD.n8856 0.468749
R32703 VDD.n8852 VDD.n8851 0.468749
R32704 VDD.n8516 VDD.n8515 0.468749
R32705 VDD.n8870 VDD.n8868 0.468749
R32706 VDD.n8866 VDD.n8864 0.468749
R32707 VDD.n8861 VDD.n8859 0.468749
R32708 VDD.n8857 VDD.n8855 0.468749
R32709 VDD.n8852 VDD.n8850 0.468749
R32710 VDD.n8516 VDD.n8514 0.468749
R32711 VDD.n8524 VDD.n8523 0.468749
R32712 VDD.n8783 VDD.n8782 0.468749
R32713 VDD.n8787 VDD.n8786 0.468749
R32714 VDD.n8790 VDD.n8789 0.468749
R32715 VDD.n8794 VDD.n8793 0.468749
R32716 VDD.n8797 VDD.n8796 0.468749
R32717 VDD.n8524 VDD.n8522 0.468749
R32718 VDD.n8783 VDD.n8780 0.468749
R32719 VDD.n8787 VDD.n8779 0.468749
R32720 VDD.n8790 VDD.n8778 0.468749
R32721 VDD.n8794 VDD.n8777 0.468749
R32722 VDD.n8797 VDD.n8776 0.468749
R32723 VDD.n8562 VDD.n8561 0.468749
R32724 VDD.n8565 VDD.n8564 0.468749
R32725 VDD.n8569 VDD.n8568 0.468749
R32726 VDD.n8572 VDD.n8571 0.468749
R32727 VDD.n8576 VDD.n8575 0.468749
R32728 VDD.n8579 VDD.n8578 0.468749
R32729 VDD.n8562 VDD.n8542 0.468749
R32730 VDD.n8565 VDD.n8541 0.468749
R32731 VDD.n8569 VDD.n8540 0.468749
R32732 VDD.n8572 VDD.n8534 0.468749
R32733 VDD.n8576 VDD.n8533 0.468749
R32734 VDD.n8579 VDD.n8532 0.468749
R32735 VDD.n9169 VDD.n9168 0.468749
R32736 VDD.n9172 VDD.n9171 0.468749
R32737 VDD.n9176 VDD.n9175 0.468749
R32738 VDD.n8465 VDD.n8464 0.468749
R32739 VDD.n9080 VDD.n9079 0.468749
R32740 VDD.n9083 VDD.n9082 0.468749
R32741 VDD.n9169 VDD.n8469 0.468749
R32742 VDD.n9172 VDD.n8468 0.468749
R32743 VDD.n9176 VDD.n8467 0.468749
R32744 VDD.n8465 VDD.n8463 0.468749
R32745 VDD.n9080 VDD.n9076 0.468749
R32746 VDD.n9083 VDD.n9075 0.468749
R32747 VDD.n9136 VDD.n9087 0.468749
R32748 VDD.n9138 VDD.n9086 0.468749
R32749 VDD.n9124 VDD.n9089 0.468749
R32750 VDD.n9126 VDD.n9088 0.468749
R32751 VDD.n12451 VDD.n12450 0.468749
R32752 VDD.n12454 VDD.n12453 0.468749
R32753 VDD.n12458 VDD.n12457 0.468749
R32754 VDD.n180 VDD.n179 0.468749
R32755 VDD.n8588 VDD.n8587 0.468749
R32756 VDD.n8591 VDD.n8590 0.468749
R32757 VDD.n12451 VDD.n183 0.468749
R32758 VDD.n12454 VDD.n182 0.468749
R32759 VDD.n12458 VDD.n181 0.468749
R32760 VDD.n180 VDD.n178 0.468749
R32761 VDD.n8588 VDD.n8584 0.468749
R32762 VDD.n8591 VDD.n8583 0.468749
R32763 VDD.n134 VDD.n133 0.468749
R32764 VDD.n130 VDD.n129 0.468749
R32765 VDD.n122 VDD.n121 0.468749
R32766 VDD.n119 VDD.n118 0.468749
R32767 VDD.n8731 VDD.n8730 0.468749
R32768 VDD.n8734 VDD.n8733 0.468749
R32769 VDD.n134 VDD.n132 0.468749
R32770 VDD.n130 VDD.n128 0.468749
R32771 VDD.n122 VDD.n120 0.468749
R32772 VDD.n119 VDD.n117 0.468749
R32773 VDD.n8731 VDD.n8727 0.468749
R32774 VDD.n8734 VDD.n8726 0.468749
R32775 VDD.n12486 VDD.n12485 0.468749
R32776 VDD.n12482 VDD.n12481 0.468749
R32777 VDD.n12477 VDD.n12476 0.468749
R32778 VDD.n109 VDD.n108 0.468749
R32779 VDD.n8601 VDD.n8600 0.468749
R32780 VDD.n8604 VDD.n8603 0.468749
R32781 VDD.n12486 VDD.n12484 0.468749
R32782 VDD.n12482 VDD.n12480 0.468749
R32783 VDD.n12477 VDD.n12475 0.468749
R32784 VDD.n109 VDD.n107 0.468749
R32785 VDD.n8601 VDD.n8597 0.468749
R32786 VDD.n8604 VDD.n8596 0.468749
R32787 VDD.n12507 VDD.n12506 0.468749
R32788 VDD.n12510 VDD.n12509 0.468749
R32789 VDD.n12514 VDD.n12513 0.468749
R32790 VDD.n100 VDD.n99 0.468749
R32791 VDD.n8693 VDD.n8692 0.468749
R32792 VDD.n8696 VDD.n8695 0.468749
R32793 VDD.n12507 VDD.n103 0.468749
R32794 VDD.n12510 VDD.n102 0.468749
R32795 VDD.n12514 VDD.n101 0.468749
R32796 VDD.n100 VDD.n98 0.468749
R32797 VDD.n8693 VDD.n8689 0.468749
R32798 VDD.n8696 VDD.n8688 0.468749
R32799 VDD.n88 VDD.n87 0.468749
R32800 VDD.n84 VDD.n83 0.468749
R32801 VDD.n42 VDD.n41 0.468749
R32802 VDD.n39 VDD.n38 0.468749
R32803 VDD.n8615 VDD.n8614 0.468749
R32804 VDD.n8618 VDD.n8617 0.468749
R32805 VDD.n88 VDD.n86 0.468749
R32806 VDD.n84 VDD.n82 0.468749
R32807 VDD.n42 VDD.n40 0.468749
R32808 VDD.n39 VDD.n37 0.468749
R32809 VDD.n8615 VDD.n8611 0.468749
R32810 VDD.n8618 VDD.n8610 0.468749
R32811 VDD.n12542 VDD.n12541 0.468749
R32812 VDD.n12538 VDD.n12537 0.468749
R32813 VDD.n12533 VDD.n12532 0.468749
R32814 VDD.n29 VDD.n28 0.468749
R32815 VDD.n8660 VDD.n8659 0.468749
R32816 VDD.n8663 VDD.n8662 0.468749
R32817 VDD.n12542 VDD.n12540 0.468749
R32818 VDD.n12538 VDD.n12536 0.468749
R32819 VDD.n12533 VDD.n12531 0.468749
R32820 VDD.n29 VDD.n27 0.468749
R32821 VDD.n8660 VDD.n8656 0.468749
R32822 VDD.n8663 VDD.n8655 0.468749
R32823 VDD.n12601 VDD.n12600 0.468749
R32824 VDD.n12604 VDD.n12603 0.468749
R32825 VDD.n12608 VDD.n12607 0.468749
R32826 VDD.n20 VDD.n19 0.468749
R32827 VDD.n8629 VDD.n8628 0.468749
R32828 VDD.n8632 VDD.n8631 0.468749
R32829 VDD.n12601 VDD.n23 0.468749
R32830 VDD.n12604 VDD.n22 0.468749
R32831 VDD.n12608 VDD.n21 0.468749
R32832 VDD.n20 VDD.n18 0.468749
R32833 VDD.n8629 VDD.n8625 0.468749
R32834 VDD.n8632 VDD.n8624 0.468749
R32835 VDD.n12558 VDD.n12557 0.468749
R32836 VDD.n12576 VDD.n12575 0.468749
R32837 VDD.n12572 VDD.n12571 0.468749
R32838 VDD.n12569 VDD.n12568 0.468749
R32839 VDD.n12565 VDD.n12564 0.468749
R32840 VDD.n12625 VDD.n12624 0.468749
R32841 VDD.n71 VDD.n62 0.3755
R32842 VDD.n160 VDD.n151 0.3755
R32843 VDD.n5770 VDD.n5761 0.3755
R32844 VDD.n5837 VDD.n5828 0.3755
R32845 VDD.n5654 VDD.n5645 0.3755
R32846 VDD.n5572 VDD.n5563 0.3755
R32847 VDD.n8158 VDD.n8149 0.3755
R32848 VDD.n5912 VDD.n5911 0.3755
R32849 VDD.n5886 VDD.n5539 0.3755
R32850 VDD.n6326 VDD.n6325 0.3755
R32851 VDD.n8090 VDD.n8089 0.3755
R32852 VDD.n9115 VDD.n9106 0.3755
R32853 VDD.n8828 VDD.n8819 0.3755
R32854 VDD.n8968 VDD.n8959 0.3755
R32855 VDD.n1000 VDD.n6 0.3755
R32856 VDD.n12635 VDD.n12634 0.3755
R32857 VDD.n12633 VDD.n12632 0.3755
R32858 VDD.n12579 VDD.n7 0.3755
R32859 VDD.n1762 VDD.n638 0.3755
R32860 VDD.n1761 VDD.n1760 0.3755
R32861 VDD.n6713 VDD.n2409 0.355763
R32862 VDD.n6713 VDD.n2410 0.281286
R32863 VDD.n1556 VDD.n1555 0.249951
R32864 VDD.n1557 VDD.n1556 0.249951
R32865 VDD.n7022 VDD.n2383 0.236091
R32866 VDD.n6975 VDD.n6966 0.236091
R32867 VDD.n6551 VDD.n5296 0.236091
R32868 VDD.n6512 VDD.n6511 0.236091
R32869 VDD.n1555 VDD.n1554 0.192465
R32870 VDD.n1558 VDD.n1557 0.192465
R32871 VDD.n6713 VDD.n2408 0.177356
R32872 VDD.n1442 VDD.n1441 0.174614
R32873 VDD.n1610 VDD.n804 0.174614
R32874 VDD.n1610 VDD.n803 0.174614
R32875 VDD.n1480 VDD.n814 0.174614
R32876 VDD.n1480 VDD.n1479 0.174614
R32877 VDD.n2136 VDD.n2123 0.166289
R32878 VDD.n2162 VDD.n2124 0.166289
R32879 VDD.n2354 VDD.n2124 0.166289
R32880 VDD.n61 VDD.n58 0.157683
R32881 VDD.n70 VDD.n63 0.157683
R32882 VDD.n150 VDD.n147 0.157683
R32883 VDD.n159 VDD.n152 0.157683
R32884 VDD.n5769 VDD.n5762 0.157683
R32885 VDD.n5760 VDD.n5757 0.157683
R32886 VDD.n5836 VDD.n5829 0.157683
R32887 VDD.n5827 VDD.n5824 0.157683
R32888 VDD.n5653 VDD.n5646 0.157683
R32889 VDD.n5644 VDD.n5641 0.157683
R32890 VDD.n5571 VDD.n5564 0.157683
R32891 VDD.n5562 VDD.n5559 0.157683
R32892 VDD.n8157 VDD.n8150 0.157683
R32893 VDD.n8148 VDD.n8145 0.157683
R32894 VDD.n9105 VDD.n9102 0.157683
R32895 VDD.n9114 VDD.n9107 0.157683
R32896 VDD.n8818 VDD.n8815 0.157683
R32897 VDD.n8827 VDD.n8820 0.157683
R32898 VDD.n8958 VDD.n8955 0.157683
R32899 VDD.n8967 VDD.n8960 0.157683
R32900 VDD.n6149 VDD.n6148 0.150184
R32901 VDD.n6075 VDD.n6056 0.150184
R32902 VDD.n6823 VDD.n6822 0.150184
R32903 VDD.n6790 VDD.n6789 0.150184
R32904 VDD.n12449 VDD.n12448 0.143306
R32905 VDD.n6887 VDD.n6885 0.14
R32906 VDD.n6891 VDD.n6885 0.14
R32907 VDD.n6892 VDD.n6884 0.14
R32908 VDD.n6896 VDD.n6884 0.14
R32909 VDD.n6897 VDD.n6883 0.14
R32910 VDD.n6901 VDD.n6883 0.14
R32911 VDD.n6979 VDD.n6882 0.14
R32912 VDD.n6983 VDD.n6882 0.14
R32913 VDD.n6984 VDD.n6881 0.14
R32914 VDD.n6988 VDD.n6881 0.14
R32915 VDD.n6989 VDD.n6880 0.14
R32916 VDD.n6993 VDD.n6880 0.14
R32917 VDD.n6994 VDD.n6879 0.14
R32918 VDD.n6998 VDD.n6879 0.14
R32919 VDD.n6906 VDD.n6904 0.14
R32920 VDD.n6910 VDD.n6904 0.14
R32921 VDD.n6911 VDD.n6903 0.14
R32922 VDD.n6915 VDD.n6903 0.14
R32923 VDD.n6916 VDD.n6902 0.14
R32924 VDD.n6920 VDD.n6902 0.14
R32925 VDD.n6931 VDD.n6930 0.14
R32926 VDD.n6935 VDD.n6930 0.14
R32927 VDD.n6936 VDD.n6929 0.14
R32928 VDD.n6940 VDD.n6929 0.14
R32929 VDD.n6941 VDD.n6928 0.14
R32930 VDD.n6945 VDD.n6928 0.14
R32931 VDD.n6946 VDD.n6927 0.14
R32932 VDD.n6950 VDD.n6927 0.14
R32933 VDD.n6420 VDD.n6418 0.14
R32934 VDD.n6424 VDD.n6418 0.14
R32935 VDD.n6425 VDD.n6417 0.14
R32936 VDD.n6429 VDD.n6417 0.14
R32937 VDD.n6430 VDD.n6416 0.14
R32938 VDD.n6434 VDD.n6416 0.14
R32939 VDD.n6534 VDD.n6435 0.14
R32940 VDD.n6532 VDD.n6435 0.14
R32941 VDD.n6531 VDD.n6438 0.14
R32942 VDD.n6529 VDD.n6438 0.14
R32943 VDD.n6528 VDD.n6441 0.14
R32944 VDD.n6526 VDD.n6441 0.14
R32945 VDD.n6525 VDD.n6444 0.14
R32946 VDD.n6523 VDD.n6444 0.14
R32947 VDD.n6457 VDD.n6455 0.14
R32948 VDD.n6461 VDD.n6455 0.14
R32949 VDD.n6462 VDD.n6454 0.14
R32950 VDD.n6466 VDD.n6454 0.14
R32951 VDD.n6467 VDD.n6453 0.14
R32952 VDD.n6471 VDD.n6453 0.14
R32953 VDD.n6494 VDD.n6472 0.14
R32954 VDD.n6492 VDD.n6472 0.14
R32955 VDD.n6491 VDD.n6475 0.14
R32956 VDD.n6489 VDD.n6475 0.14
R32957 VDD.n6488 VDD.n6478 0.14
R32958 VDD.n6486 VDD.n6478 0.14
R32959 VDD.n6485 VDD.n6481 0.14
R32960 VDD.n6481 VDD.n6447 0.14
R32961 VDD.n6101 VDD.n6040 0.14
R32962 VDD.n6104 VDD.n6040 0.14
R32963 VDD.n6105 VDD.n6039 0.14
R32964 VDD.n6109 VDD.n6039 0.14
R32965 VDD.n6115 VDD.n6110 0.14
R32966 VDD.n6113 VDD.n6110 0.14
R32967 VDD.n6058 VDD.n6041 0.14
R32968 VDD.n6061 VDD.n6058 0.14
R32969 VDD.n6062 VDD.n6057 0.14
R32970 VDD.n6066 VDD.n6057 0.14
R32971 VDD.n6072 VDD.n6067 0.14
R32972 VDD.n6070 VDD.n6067 0.14
R32973 VDD.n7913 VDD.n7860 0.14
R32974 VDD.n7917 VDD.n7860 0.14
R32975 VDD.n7918 VDD.n7859 0.14
R32976 VDD.n7922 VDD.n7859 0.14
R32977 VDD.n7923 VDD.n7858 0.14
R32978 VDD.n7926 VDD.n7858 0.14
R32979 VDD.n7927 VDD.n7857 0.14
R32980 VDD.n7931 VDD.n7857 0.14
R32981 VDD.n7932 VDD.n7856 0.14
R32982 VDD.n7936 VDD.n7856 0.14
R32983 VDD.n7937 VDD.n7855 0.14
R32984 VDD.n7941 VDD.n7855 0.14
R32985 VDD.n7908 VDD.n7865 0.14
R32986 VDD.n7906 VDD.n7865 0.14
R32987 VDD.n7905 VDD.n7869 0.14
R32988 VDD.n7903 VDD.n7869 0.14
R32989 VDD.n7902 VDD.n7873 0.14
R32990 VDD.n7900 VDD.n7873 0.14
R32991 VDD.n7899 VDD.n7875 0.14
R32992 VDD.n7897 VDD.n7875 0.14
R32993 VDD.n7896 VDD.n7879 0.14
R32994 VDD.n7894 VDD.n7879 0.14
R32995 VDD.n7893 VDD.n7883 0.14
R32996 VDD.n7891 VDD.n7883 0.14
R32997 VDD.n8018 VDD.n2155 0.14
R32998 VDD.n8022 VDD.n2155 0.14
R32999 VDD.n8023 VDD.n2154 0.14
R33000 VDD.n8027 VDD.n2154 0.14
R33001 VDD.n8028 VDD.n2153 0.14
R33002 VDD.n8031 VDD.n2153 0.14
R33003 VDD.n8032 VDD.n2152 0.14
R33004 VDD.n8036 VDD.n2152 0.14
R33005 VDD.n8037 VDD.n2151 0.14
R33006 VDD.n8041 VDD.n2151 0.14
R33007 VDD.n8042 VDD.n2150 0.14
R33008 VDD.n8046 VDD.n2150 0.14
R33009 VDD.n6806 VDD.n6729 0.14
R33010 VDD.n6804 VDD.n6729 0.14
R33011 VDD.n6803 VDD.n6731 0.14
R33012 VDD.n6801 VDD.n6731 0.14
R33013 VDD.n6739 VDD.n6734 0.14
R33014 VDD.n6737 VDD.n6734 0.14
R33015 VDD.n6757 VDD.n6747 0.14
R33016 VDD.n6755 VDD.n6747 0.14
R33017 VDD.n6754 VDD.n6749 0.14
R33018 VDD.n6752 VDD.n6749 0.14
R33019 VDD.n6745 VDD.n6740 0.14
R33020 VDD.n6743 VDD.n6740 0.14
R33021 VDD.n6714 VDD.n6713 0.136679
R33022 VDD.n8076 VDD.n8075 0.13175
R33023 VDD.n8077 VDD.n8076 0.13175
R33024 VDD.n8079 VDD.n8078 0.13175
R33025 VDD.n8078 VDD.n8077 0.13175
R33026 VDD.n1549 VDD.n1548 0.119368
R33027 VDD.n1521 VDD.n1520 0.119368
R33028 VDD.n4906 VDD.n4697 0.110375
R33029 VDD.n4905 VDD.n4904 0.110375
R33030 VDD.n3630 VDD.n3629 0.11
R33031 VDD.n3628 VDD.n2745 0.11
R33032 VDD.n10103 VDD.n10102 0.11
R33033 VDD.n10101 VDD.n9214 0.11
R33034 VDD.n11813 VDD.n405 0.109625
R33035 VDD.n11812 VDD.n11811 0.109625
R33036 VDD.n1390 VDD.n1389 0.109121
R33037 VDD.n1414 VDD.n1390 0.109121
R33038 VDD.n1358 VDD.n1357 0.109121
R33039 VDD.n1357 VDD.n1356 0.109121
R33040 VDD.n1343 VDD.n1342 0.109121
R33041 VDD.n1349 VDD.n1343 0.109121
R33042 VDD.n1654 VDD.n1653 0.109121
R33043 VDD.n1653 VDD.n1652 0.109121
R33044 VDD.n1170 VDD.n707 0.109121
R33045 VDD.n1718 VDD.n707 0.109121
R33046 VDD.n1183 VDD.n845 0.109121
R33047 VDD.n1414 VDD.n845 0.109121
R33048 VDD.n1651 VDD.n1650 0.109121
R33049 VDD.n1652 VDD.n1651 0.109121
R33050 VDD.n1600 VDD.n761 0.109121
R33051 VDD.n1652 VDD.n761 0.109121
R33052 VDD.n1600 VDD.n760 0.109121
R33053 VDD.n1652 VDD.n760 0.109121
R33054 VDD.n1276 VDD.n1275 0.109121
R33055 VDD.n1349 VDD.n1276 0.109121
R33056 VDD.n1213 VDD.n849 0.109121
R33057 VDD.n1356 VDD.n849 0.109121
R33058 VDD.n1413 VDD.n1412 0.109121
R33059 VDD.n1414 VDD.n1413 0.109121
R33060 VDD.n1355 VDD.n818 0.109121
R33061 VDD.n1356 VDD.n1355 0.109121
R33062 VDD.n1348 VDD.n808 0.109121
R33063 VDD.n1349 VDD.n1348 0.109121
R33064 VDD.n1412 VDD.n846 0.109121
R33065 VDD.n1414 VDD.n846 0.109121
R33066 VDD.n850 VDD.n818 0.109121
R33067 VDD.n1356 VDD.n850 0.109121
R33068 VDD.n1350 VDD.n808 0.109121
R33069 VDD.n1350 VDD.n1349 0.109121
R33070 VDD.n1066 VDD.n711 0.109121
R33071 VDD.n1718 VDD.n711 0.109121
R33072 VDD.n911 VDD.n689 0.109121
R33073 VDD.n1742 VDD.n689 0.109121
R33074 VDD.n1741 VDD.n1740 0.109121
R33075 VDD.n1742 VDD.n1741 0.109121
R33076 VDD.n1740 VDD.n688 0.109121
R33077 VDD.n1742 VDD.n688 0.109121
R33078 VDD.n1717 VDD.n1716 0.109121
R33079 VDD.n1718 VDD.n1717 0.109121
R33080 VDD.n1716 VDD.n708 0.109121
R33081 VDD.n1718 VDD.n708 0.109121
R33082 VDD.n1744 VDD.n1743 0.109121
R33083 VDD.n1743 VDD.n1742 0.109121
R33084 VDD.n2074 VDD.n2025 0.10728
R33085 VDD.n8137 VDD.n2024 0.10728
R33086 VDD.n10773 VDD.n2024 0.10728
R33087 VDD.n8116 VDD.n2012 0.10728
R33088 VDD.n10781 VDD.n2012 0.10728
R33089 VDD.n10778 VDD.n10777 0.10728
R33090 VDD.n10779 VDD.n10778 0.10728
R33091 VDD.n10777 VDD.n10776 0.10728
R33092 VDD.n10776 VDD.n2017 0.10728
R33093 VDD.n10784 VDD.n2011 0.10728
R33094 VDD.n2016 VDD.n2011 0.10728
R33095 VDD.n10784 VDD.n10783 0.10728
R33096 VDD.n10783 VDD.n10782 0.10728
R33097 VDD.n8104 VDD.n1989 0.10728
R33098 VDD.n2014 VDD.n1989 0.10728
R33099 VDD.n5579 VDD.n1951 0.10728
R33100 VDD.n1988 VDD.n1951 0.10728
R33101 VDD.n10828 VDD.n1952 0.10728
R33102 VDD.n10831 VDD.n1952 0.10728
R33103 VDD.n10829 VDD.n10828 0.10728
R33104 VDD.n10830 VDD.n10829 0.10728
R33105 VDD.n10836 VDD.n10835 0.10728
R33106 VDD.n10837 VDD.n10836 0.10728
R33107 VDD.n10835 VDD.n10834 0.10728
R33108 VDD.n10834 VDD.n1944 0.10728
R33109 VDD.n5600 VDD.n1939 0.10728
R33110 VDD.n10839 VDD.n1939 0.10728
R33111 VDD.n5621 VDD.n1924 0.10728
R33112 VDD.n1941 VDD.n1924 0.10728
R33113 VDD.n10842 VDD.n1938 0.10728
R33114 VDD.n1943 VDD.n1938 0.10728
R33115 VDD.n10842 VDD.n10841 0.10728
R33116 VDD.n10841 VDD.n10840 0.10728
R33117 VDD.n10883 VDD.n1921 0.10728
R33118 VDD.n10886 VDD.n1921 0.10728
R33119 VDD.n10884 VDD.n10883 0.10728
R33120 VDD.n10885 VDD.n10884 0.10728
R33121 VDD.n5661 VDD.n1920 0.10728
R33122 VDD.n1923 VDD.n1920 0.10728
R33123 VDD.n5871 VDD.n1912 0.10728
R33124 VDD.n10894 VDD.n1912 0.10728
R33125 VDD.n10891 VDD.n10890 0.10728
R33126 VDD.n10892 VDD.n10891 0.10728
R33127 VDD.n10890 VDD.n10889 0.10728
R33128 VDD.n10889 VDD.n1917 0.10728
R33129 VDD.n10897 VDD.n1911 0.10728
R33130 VDD.n1916 VDD.n1911 0.10728
R33131 VDD.n10897 VDD.n10896 0.10728
R33132 VDD.n10896 VDD.n10895 0.10728
R33133 VDD.n5859 VDD.n1897 0.10728
R33134 VDD.n1914 VDD.n1897 0.10728
R33135 VDD.n5816 VDD.n1859 0.10728
R33136 VDD.n1896 VDD.n1859 0.10728
R33137 VDD.n10938 VDD.n1860 0.10728
R33138 VDD.n10941 VDD.n1860 0.10728
R33139 VDD.n10939 VDD.n10938 0.10728
R33140 VDD.n10940 VDD.n10939 0.10728
R33141 VDD.n10946 VDD.n10945 0.10728
R33142 VDD.n10947 VDD.n10946 0.10728
R33143 VDD.n10945 VDD.n10944 0.10728
R33144 VDD.n10944 VDD.n1852 0.10728
R33145 VDD.n5804 VDD.n1847 0.10728
R33146 VDD.n10949 VDD.n1847 0.10728
R33147 VDD.n5783 VDD.n1832 0.10728
R33148 VDD.n1849 VDD.n1832 0.10728
R33149 VDD.n10952 VDD.n1846 0.10728
R33150 VDD.n1851 VDD.n1846 0.10728
R33151 VDD.n10952 VDD.n10951 0.10728
R33152 VDD.n10951 VDD.n10950 0.10728
R33153 VDD.n10993 VDD.n1795 0.10728
R33154 VDD.n10996 VDD.n1795 0.10728
R33155 VDD.n10994 VDD.n10993 0.10728
R33156 VDD.n10995 VDD.n10994 0.10728
R33157 VDD.n5749 VDD.n1794 0.10728
R33158 VDD.n1831 VDD.n1794 0.10728
R33159 VDD.n5728 VDD.n1784 0.10728
R33160 VDD.n11004 VDD.n1784 0.10728
R33161 VDD.n11001 VDD.n11000 0.10728
R33162 VDD.n11002 VDD.n11001 0.10728
R33163 VDD.n11000 VDD.n10999 0.10728
R33164 VDD.n10999 VDD.n1787 0.10728
R33165 VDD.n11007 VDD.n1772 0.10728
R33166 VDD.n1786 VDD.n1772 0.10728
R33167 VDD.n11007 VDD.n11006 0.10728
R33168 VDD.n11006 VDD.n11005 0.10728
R33169 VDD.n11031 VDD.n11030 0.10728
R33170 VDD.n11030 VDD.n11029 0.10728
R33171 VDD.n1771 VDD.n657 0.10728
R33172 VDD.n12465 VDD.n175 0.10728
R33173 VDD.n12465 VDD.n12464 0.10728
R33174 VDD.n8570 VDD.n8539 0.10728
R33175 VDD.n8539 VDD.n8538 0.10728
R33176 VDD.n8554 VDD.n177 0.10728
R33177 VDD.n8535 VDD.n177 0.10728
R33178 VDD.n8570 VDD.n8527 0.10728
R33179 VDD.n8537 VDD.n8527 0.10728
R33180 VDD.n8788 VDD.n8528 0.10728
R33181 VDD.n8530 VDD.n8528 0.10728
R33182 VDD.n8809 VDD.n8808 0.10728
R33183 VDD.n8808 VDD.n8807 0.10728
R33184 VDD.n8788 VDD.n8519 0.10728
R33185 VDD.n8529 VDD.n8519 0.10728
R33186 VDD.n8858 VDD.n8520 0.10728
R33187 VDD.n8881 VDD.n8520 0.10728
R33188 VDD.n8878 VDD.n8877 0.10728
R33189 VDD.n8879 VDD.n8878 0.10728
R33190 VDD.n8858 VDD.n8508 0.10728
R33191 VDD.n8880 VDD.n8508 0.10728
R33192 VDD.n8919 VDD.n8509 0.10728
R33193 VDD.n8511 VDD.n8509 0.10728
R33194 VDD.n8940 VDD.n8939 0.10728
R33195 VDD.n8939 VDD.n8938 0.10728
R33196 VDD.n8919 VDD.n8500 0.10728
R33197 VDD.n8510 VDD.n8500 0.10728
R33198 VDD.n8985 VDD.n8501 0.10728
R33199 VDD.n9012 VDD.n8501 0.10728
R33200 VDD.n9009 VDD.n9008 0.10728
R33201 VDD.n9010 VDD.n9009 0.10728
R33202 VDD.n8985 VDD.n8491 0.10728
R33203 VDD.n9011 VDD.n8491 0.10728
R33204 VDD.n9053 VDD.n8480 0.10728
R33205 VDD.n8493 VDD.n8480 0.10728
R33206 VDD.n9037 VDD.n9036 0.10728
R33207 VDD.n9036 VDD.n9035 0.10728
R33208 VDD.n9053 VDD.n8473 0.10728
R33209 VDD.n8492 VDD.n8473 0.10728
R33210 VDD.n9096 VDD.n8461 0.10728
R33211 VDD.n9180 VDD.n8461 0.10728
R33212 VDD.n9161 VDD.n9160 0.10728
R33213 VDD.n9160 VDD.n9159 0.10728
R33214 VDD.n9177 VDD.n8466 0.10728
R33215 VDD.n8466 VDD.n8462 0.10728
R33216 VDD.n9178 VDD.n9177 0.10728
R33217 VDD.n9179 VDD.n9178 0.10728
R33218 VDD.n9183 VDD.n9182 0.10728
R33219 VDD.n12459 VDD.n124 0.10728
R33220 VDD.n12462 VDD.n124 0.10728
R33221 VDD.n12460 VDD.n12459 0.10728
R33222 VDD.n12461 VDD.n12460 0.10728
R33223 VDD.n12468 VDD.n12467 0.10728
R33224 VDD.n12469 VDD.n12468 0.10728
R33225 VDD.n12467 VDD.n12466 0.10728
R33226 VDD.n12466 VDD.n116 0.10728
R33227 VDD.n141 VDD.n112 0.10728
R33228 VDD.n12471 VDD.n112 0.10728
R33229 VDD.n12493 VDD.n97 0.10728
R33230 VDD.n113 VDD.n97 0.10728
R33231 VDD.n12474 VDD.n110 0.10728
R33232 VDD.n115 VDD.n110 0.10728
R33233 VDD.n12474 VDD.n12473 0.10728
R33234 VDD.n12473 VDD.n12472 0.10728
R33235 VDD.n12515 VDD.n44 0.10728
R33236 VDD.n12518 VDD.n44 0.10728
R33237 VDD.n12516 VDD.n12515 0.10728
R33238 VDD.n12517 VDD.n12516 0.10728
R33239 VDD.n12521 VDD.n95 0.10728
R33240 VDD.n12521 VDD.n12520 0.10728
R33241 VDD.n52 VDD.n32 0.10728
R33242 VDD.n12527 VDD.n32 0.10728
R33243 VDD.n12524 VDD.n12523 0.10728
R33244 VDD.n12525 VDD.n12524 0.10728
R33245 VDD.n12523 VDD.n12522 0.10728
R33246 VDD.n12522 VDD.n36 0.10728
R33247 VDD.n12530 VDD.n30 0.10728
R33248 VDD.n35 VDD.n30 0.10728
R33249 VDD.n12530 VDD.n12529 0.10728
R33250 VDD.n12529 VDD.n12528 0.10728
R33251 VDD.n12549 VDD.n17 0.10728
R33252 VDD.n33 VDD.n17 0.10728
R33253 VDD.n12593 VDD.n12592 0.10728
R33254 VDD.n12592 VDD.n15 0.10728
R33255 VDD.n12609 VDD.n14 0.10728
R33256 VDD.n12612 VDD.n14 0.10728
R33257 VDD.n12610 VDD.n12609 0.10728
R33258 VDD.n12611 VDD.n12610 0.10728
R33259 VDD.n12570 VDD.n13 0.10728
R33260 VDD.n7841 VDD.n7840 0.105779
R33261 VDD.n2389 VDD.n2388 0.105779
R33262 VDD.n10775 VDD.n10772 0.1055
R33263 VDD.n10775 VDD.n10774 0.1055
R33264 VDD.n2048 VDD.n2013 0.1055
R33265 VDD.n10780 VDD.n2013 0.1055
R33266 VDD.n10803 VDD.n1990 0.1055
R33267 VDD.n2015 VDD.n1990 0.1055
R33268 VDD.n10833 VDD.n1987 0.1055
R33269 VDD.n10833 VDD.n10832 0.1055
R33270 VDD.n1966 VDD.n1940 0.1055
R33271 VDD.n10838 VDD.n1940 0.1055
R33272 VDD.n10861 VDD.n1925 0.1055
R33273 VDD.n1942 VDD.n1925 0.1055
R33274 VDD.n10888 VDD.n1922 0.1055
R33275 VDD.n10888 VDD.n10887 0.1055
R33276 VDD.n5522 VDD.n1913 0.1055
R33277 VDD.n10893 VDD.n1913 0.1055
R33278 VDD.n10916 VDD.n1898 0.1055
R33279 VDD.n1915 VDD.n1898 0.1055
R33280 VDD.n10943 VDD.n1895 0.1055
R33281 VDD.n10943 VDD.n10942 0.1055
R33282 VDD.n1874 VDD.n1848 0.1055
R33283 VDD.n10948 VDD.n1848 0.1055
R33284 VDD.n10971 VDD.n1833 0.1055
R33285 VDD.n1850 VDD.n1833 0.1055
R33286 VDD.n10998 VDD.n1830 0.1055
R33287 VDD.n10998 VDD.n10997 0.1055
R33288 VDD.n1818 VDD.n1785 0.1055
R33289 VDD.n11003 VDD.n1785 0.1055
R33290 VDD.n11027 VDD.n11026 0.1055
R33291 VDD.n11028 VDD.n11027 0.1055
R33292 VDD.n8758 VDD.n176 0.1055
R33293 VDD.n8536 VDD.n176 0.1055
R33294 VDD.n8805 VDD.n8804 0.1055
R33295 VDD.n8806 VDD.n8805 0.1055
R33296 VDD.n8884 VDD.n8883 0.1055
R33297 VDD.n8883 VDD.n8882 0.1055
R33298 VDD.n8936 VDD.n8935 0.1055
R33299 VDD.n8937 VDD.n8936 0.1055
R33300 VDD.n9015 VDD.n9014 0.1055
R33301 VDD.n9014 VDD.n9013 0.1055
R33302 VDD.n9033 VDD.n9032 0.1055
R33303 VDD.n9034 VDD.n9033 0.1055
R33304 VDD.n9157 VDD.n9156 0.1055
R33305 VDD.n9158 VDD.n9157 0.1055
R33306 VDD.n9144 VDD.n8460 0.1055
R33307 VDD.n9181 VDD.n8460 0.1055
R33308 VDD.n8741 VDD.n123 0.1055
R33309 VDD.n12463 VDD.n123 0.1055
R33310 VDD.n8720 VDD.n111 0.1055
R33311 VDD.n12470 VDD.n111 0.1055
R33312 VDD.n8708 VDD.n96 0.1055
R33313 VDD.n114 VDD.n96 0.1055
R33314 VDD.n8682 VDD.n43 0.1055
R33315 VDD.n12519 VDD.n43 0.1055
R33316 VDD.n8670 VDD.n31 0.1055
R33317 VDD.n12526 VDD.n31 0.1055
R33318 VDD.n8649 VDD.n16 0.1055
R33319 VDD.n34 VDD.n16 0.1055
R33320 VDD.n12615 VDD.n12614 0.1055
R33321 VDD.n12614 VDD.n12613 0.1055
R33322 VDD.n7176 VDD.n7175 0.101802
R33323 VDD.n7175 VDD.n2296 0.101802
R33324 VDD.n7828 VDD.n7827 0.101802
R33325 VDD.n7827 VDD.n7826 0.101802
R33326 VDD.n6978 VDD.n6901 0.10175
R33327 VDD.n6921 VDD.n6920 0.10175
R33328 VDD.n6535 VDD.n6434 0.10175
R33329 VDD.n6495 VDD.n6471 0.10175
R33330 VDD.n6313 VDD.n6312 0.0931471
R33331 VDD.n6312 VDD.n6311 0.0931471
R33332 VDD.n5943 VDD.n5942 0.0931471
R33333 VDD.n5942 VDD.n5376 0.0931471
R33334 VDD.n5943 VDD.n5275 0.0931471
R33335 VDD.n6370 VDD.n5275 0.0931471
R33336 VDD.n7135 VDD.n2312 0.0931471
R33337 VDD.n2317 VDD.n2312 0.0931471
R33338 VDD.n7135 VDD.n7134 0.0931471
R33339 VDD.n7134 VDD.n7133 0.0931471
R33340 VDD.n7836 VDD.n7835 0.0931471
R33341 VDD.n7835 VDD.n7834 0.0931471
R33342 VDD.n6310 VDD.n6309 0.0931471
R33343 VDD.n6311 VDD.n6310 0.0931471
R33344 VDD.n6368 VDD.n5378 0.0931471
R33345 VDD.n5378 VDD.n5376 0.0931471
R33346 VDD.n6369 VDD.n6368 0.0931471
R33347 VDD.n6370 VDD.n6369 0.0931471
R33348 VDD.n2367 VDD.n2366 0.0931471
R33349 VDD.n2367 VDD.n2317 0.0931471
R33350 VDD.n2366 VDD.n2319 0.0931471
R33351 VDD.n7133 VDD.n2319 0.0931471
R33352 VDD.n6195 VDD.n5311 0.0931471
R33353 VDD.n6311 VDD.n5311 0.0931471
R33354 VDD.n6372 VDD.n5312 0.0931471
R33355 VDD.n5376 VDD.n5312 0.0931471
R33356 VDD.n6372 VDD.n6371 0.0931471
R33357 VDD.n6371 VDD.n6370 0.0931471
R33358 VDD.n6185 VDD.n5303 0.0931471
R33359 VDD.n6311 VDD.n5303 0.0931471
R33360 VDD.n5368 VDD.n5304 0.0931471
R33361 VDD.n5376 VDD.n5304 0.0931471
R33362 VDD.n5368 VDD.n5282 0.0931471
R33363 VDD.n6370 VDD.n5282 0.0931471
R33364 VDD.n7833 VDD.n7832 0.0931471
R33365 VDD.n7834 VDD.n7833 0.0931471
R33366 VDD.n6631 VDD.n5270 0.0931471
R33367 VDD.n5270 VDD.n5268 0.0931471
R33368 VDD.n6632 VDD.n6631 0.0931471
R33369 VDD.n6633 VDD.n6632 0.0931471
R33370 VDD.n6635 VDD.n5266 0.0931471
R33371 VDD.n5268 VDD.n5266 0.0931471
R33372 VDD.n6635 VDD.n6634 0.0931471
R33373 VDD.n6634 VDD.n6633 0.0931471
R33374 VDD.n6692 VDD.n5264 0.0931471
R33375 VDD.n5268 VDD.n5264 0.0931471
R33376 VDD.n6692 VDD.n2349 0.0931471
R33377 VDD.n6633 VDD.n2349 0.0931471
R33378 VDD.n6706 VDD.n5221 0.0931471
R33379 VDD.n5268 VDD.n5221 0.0931471
R33380 VDD.n6706 VDD.n2369 0.0931471
R33381 VDD.n6633 VDD.n2369 0.0931471
R33382 VDD.n7043 VDD.n7042 0.0931471
R33383 VDD.n7042 VDD.n2317 0.0931471
R33384 VDD.n7043 VDD.n2318 0.0931471
R33385 VDD.n7133 VDD.n2318 0.0931471
R33386 VDD.n7131 VDD.n2321 0.0931471
R33387 VDD.n2321 VDD.n2317 0.0931471
R33388 VDD.n7132 VDD.n7131 0.0931471
R33389 VDD.n7133 VDD.n7132 0.0931471
R33390 VDD.n7700 VDD.n2236 0.0931471
R33391 VDD.n7834 VDD.n2236 0.0931471
R33392 VDD.n7821 VDD.n2235 0.0931471
R33393 VDD.n7834 VDD.n2235 0.0931471
R33394 VDD.n6318 VDD.n6317 0.0831095
R33395 VDD.n6181 VDD.n6180 0.0831095
R33396 VDD.n6301 VDD.n6300 0.0799891
R33397 VDD.n6305 VDD.n5487 0.0799891
R33398 VDD.n5984 VDD.n5487 0.0799891
R33399 VDD.n6191 VDD.n6190 0.0799891
R33400 VDD.n6300 VDD.n6199 0.0799891
R33401 VDD.n6190 VDD.n6189 0.0799891
R33402 VDD.n7864 VDD.n2187 0.0737558
R33403 VDD.n2355 VDD.n2187 0.0737558
R33404 VDD.n7889 VDD.n2188 0.0737558
R33405 VDD.n7837 VDD.n7836 0.0723953
R33406 VDD.n7832 VDD.n7831 0.0723953
R33407 VDD.n2130 VDD.n2128 0.0720299
R33408 VDD.n8047 VDD.n2149 0.0692176
R33409 VDD.n7994 VDD.n7993 0.0682419
R33410 VDD.n7995 VDD.n7994 0.0682419
R33411 VDD.n7997 VDD.n7996 0.0682419
R33412 VDD.n7996 VDD.n7995 0.0682419
R33413 VDD.n5481 VDD.n5309 0.0682419
R33414 VDD.n6396 VDD.n5309 0.0682419
R33415 VDD.n5459 VDD.n5279 0.0682419
R33416 VDD.n6577 VDD.n5279 0.0682419
R33417 VDD.n5420 VDD.n2357 0.0682419
R33418 VDD.n7040 VDD.n2357 0.0682419
R33419 VDD.n2305 VDD.n2210 0.0682419
R33420 VDD.n7086 VDD.n2210 0.0682419
R33421 VDD.n6283 VDD.n5310 0.0682419
R33422 VDD.n6396 VDD.n5310 0.0682419
R33423 VDD.n6247 VDD.n5280 0.0682419
R33424 VDD.n6577 VDD.n5280 0.0682419
R33425 VDD.n6395 VDD.n6394 0.0682419
R33426 VDD.n6396 VDD.n6395 0.0682419
R33427 VDD.n5348 VDD.n5281 0.0682419
R33428 VDD.n6577 VDD.n5281 0.0682419
R33429 VDD.n5249 VDD.n2348 0.0682419
R33430 VDD.n7040 VDD.n2348 0.0682419
R33431 VDD.n6398 VDD.n6397 0.0682419
R33432 VDD.n6397 VDD.n6396 0.0682419
R33433 VDD.n6576 VDD.n6575 0.0682419
R33434 VDD.n6577 VDD.n6576 0.0682419
R33435 VDD.n6861 VDD.n2237 0.0682419
R33436 VDD.n7086 VDD.n2237 0.0682419
R33437 VDD.n7039 VDD.n7038 0.0682419
R33438 VDD.n7040 VDD.n7039 0.0682419
R33439 VDD.n2368 VDD.n2350 0.0682419
R33440 VDD.n7040 VDD.n2368 0.0682419
R33441 VDD.n7085 VDD.n7084 0.0682419
R33442 VDD.n7086 VDD.n7085 0.0682419
R33443 VDD.n7110 VDD.n7087 0.0682419
R33444 VDD.n7087 VDD.n7086 0.0682419
R33445 VDD.n1563 VDD.n1511 0.0677787
R33446 VDD.n1561 VDD.n1511 0.0677787
R33447 VDD.n1561 VDD.n1560 0.0677787
R33448 VDD.n1560 VDD.n1559 0.0677787
R33449 VDD.n1538 VDD.n1537 0.0677787
R33450 VDD.n1539 VDD.n1538 0.0677787
R33451 VDD.n1539 VDD.n1536 0.0677787
R33452 VDD.n1541 VDD.n1536 0.0677787
R33453 VDD.n1514 VDD.n771 0.0677787
R33454 VDD.n1515 VDD.n1514 0.0677787
R33455 VDD.n1515 VDD.n1513 0.0677787
R33456 VDD.n1517 VDD.n1513 0.0677787
R33457 VDD.n1525 VDD.n1518 0.0677787
R33458 VDD.n1526 VDD.n1525 0.0677787
R33459 VDD.n1526 VDD.n1524 0.0677787
R33460 VDD.n1528 VDD.n1524 0.0677787
R33461 VDD.n5965 VDD.n5308 0.0668158
R33462 VDD.n6396 VDD.n5308 0.0668158
R33463 VDD.n6579 VDD.n6578 0.0668158
R33464 VDD.n6578 VDD.n6577 0.0668158
R33465 VDD.n6610 VDD.n2353 0.0668158
R33466 VDD.n7040 VDD.n2353 0.0668158
R33467 VDD.n2234 VDD.n2233 0.0668158
R33468 VDD.n7086 VDD.n2234 0.0668158
R33469 VDD.n5481 VDD.n5307 0.0668158
R33470 VDD.n6396 VDD.n5307 0.0668158
R33471 VDD.n5459 VDD.n5278 0.0668158
R33472 VDD.n6577 VDD.n5278 0.0668158
R33473 VDD.n5420 VDD.n2352 0.0668158
R33474 VDD.n7040 VDD.n2352 0.0668158
R33475 VDD.n2332 VDD.n2305 0.0668158
R33476 VDD.n7086 VDD.n2332 0.0668158
R33477 VDD.n6283 VDD.n5306 0.0668158
R33478 VDD.n6396 VDD.n5306 0.0668158
R33479 VDD.n6247 VDD.n5277 0.0668158
R33480 VDD.n6577 VDD.n5277 0.0668158
R33481 VDD.n6394 VDD.n5305 0.0668158
R33482 VDD.n6396 VDD.n5305 0.0668158
R33483 VDD.n5348 VDD.n5276 0.0668158
R33484 VDD.n6577 VDD.n5276 0.0668158
R33485 VDD.n5249 VDD.n2351 0.0668158
R33486 VDD.n7040 VDD.n2351 0.0668158
R33487 VDD.n7041 VDD.n2350 0.0668158
R33488 VDD.n7041 VDD.n7040 0.0668158
R33489 VDD.n7084 VDD.n2331 0.0668158
R33490 VDD.n7086 VDD.n2331 0.0668158
R33491 VDD.n7110 VDD.n2238 0.0668158
R33492 VDD.n7086 VDD.n2238 0.0668158
R33493 VDD.n7836 VDD.n2209 0.0629767
R33494 VDD.n7832 VDD.n2239 0.0629767
R33495 VDD.n1553 VDD.n1552 0.0628762
R33496 VDD.n1552 VDD.n1551 0.0628762
R33497 VDD.n752 VDD.n751 0.0627244
R33498 VDD.n1507 VDD.n1506 0.0627244
R33499 VDD.n7947 VDD.n7853 0.0619118
R33500 VDD.n1550 VDD.n1512 0.061665
R33501 VDD.n1551 VDD.n1550 0.061665
R33502 VDD.n7960 VDD.n7959 0.0616241
R33503 VDD.n7823 VDD.n7822 0.0585814
R33504 VDD.n6309 VDD.n6308 0.0569142
R33505 VDD.n6314 VDD.n6313 0.0569142
R33506 VDD.n6196 VDD.n6195 0.0569142
R33507 VDD.n6186 VDD.n6185 0.0569142
R33508 VDD.n847 VDD.n739 0.0543462
R33509 VDD.n1429 VDD.n847 0.0543462
R33510 VDD.n848 VDD.n738 0.0543462
R33511 VDD.n1428 VDD.n848 0.0543462
R33512 VDD.n1347 VDD.n744 0.0543462
R33513 VDD.n1347 VDD.n1346 0.0543462
R33514 VDD.n758 VDD.n744 0.0543462
R33515 VDD.n1345 VDD.n758 0.0543462
R33516 VDD.n1417 VDD.n859 0.0543462
R33517 VDD.n874 VDD.n859 0.0543462
R33518 VDD.n1417 VDD.n1416 0.0543462
R33519 VDD.n1416 VDD.n1415 0.0543462
R33520 VDD.n1431 VDD.n1430 0.0543462
R33521 VDD.n1430 VDD.n1429 0.0543462
R33522 VDD.n1427 VDD.n1426 0.0543462
R33523 VDD.n1428 VDD.n1427 0.0543462
R33524 VDD.n1627 VDD.n764 0.0543462
R33525 VDD.n764 VDD.n763 0.0543462
R33526 VDD.n759 VDD.n747 0.0543462
R33527 VDD.n763 VDD.n759 0.0543462
R33528 VDD.n1277 VDD.n783 0.0543462
R33529 VDD.n1346 VDD.n1277 0.0543462
R33530 VDD.n783 VDD.n762 0.0543462
R33531 VDD.n1345 VDD.n762 0.0543462
R33532 VDD.n1353 VDD.n1352 0.0543462
R33533 VDD.n1354 VDD.n1353 0.0543462
R33534 VDD.n1352 VDD.n1351 0.0543462
R33535 VDD.n1351 VDD.n1084 0.0543462
R33536 VDD.n1083 VDD.n741 0.0543462
R33537 VDD.n1354 VDD.n1083 0.0543462
R33538 VDD.n1344 VDD.n741 0.0543462
R33539 VDD.n1344 VDD.n1084 0.0543462
R33540 VDD.n736 VDD.n712 0.0543462
R33541 VDD.n874 VDD.n712 0.0543462
R33542 VDD.n875 VDD.n736 0.0543462
R33543 VDD.n1415 VDD.n875 0.0543462
R33544 VDD.n1046 VDD.n710 0.0543462
R33545 VDD.n1719 VDD.n710 0.0543462
R33546 VDD.n1046 VDD.n692 0.0543462
R33547 VDD.n709 VDD.n692 0.0543462
R33548 VDD.n1721 VDD.n687 0.0543462
R33549 VDD.n709 VDD.n687 0.0543462
R33550 VDD.n1721 VDD.n1720 0.0543462
R33551 VDD.n1720 VDD.n1719 0.0543462
R33552 VDD.n1032 VDD.n691 0.0543462
R33553 VDD.n691 VDD.n690 0.0543462
R33554 VDD.n985 VDD.n686 0.0543462
R33555 VDD.n690 VDD.n686 0.0543462
R33556 VDD.n5364 VDD.n5363 0.0525345
R33557 VDD.n5373 VDD.n5372 0.0525345
R33558 VDD.n6377 VDD.n6376 0.0525345
R33559 VDD.n6364 VDD.n6363 0.0525345
R33560 VDD.n5938 VDD.n5937 0.0525345
R33561 VDD.n5948 VDD.n5947 0.0525345
R33562 VDD.n2362 VDD.n2361 0.0525345
R33563 VDD.n7140 VDD.n7139 0.0525345
R33564 VDD.n2400 VDD.n2399 0.0525345
R33565 VDD.n7127 VDD.n7126 0.0525345
R33566 VDD.n2344 VDD.n2343 0.0525345
R33567 VDD.n2128 VDD.n2122 0.0513315
R33568 VDD.n7889 VDD.n7888 0.0507941
R33569 VDD.n6266 VDD.n6218 0.050569
R33570 VDD.n6266 VDD.n6265 0.050569
R33571 VDD.n7048 VDD.n2341 0.050569
R33572 VDD.n2313 VDD.n2199 0.050569
R33573 VDD.n7048 VDD.n7047 0.050569
R33574 VDD.n6309 VDD.n6304 0.0495237
R33575 VDD.n6313 VDD.n5987 0.0495237
R33576 VDD.n6195 VDD.n6194 0.0495237
R33577 VDD.n6185 VDD.n6184 0.0495237
R33578 VDD.n8084 VDD.n2121 0.0465048
R33579 VDD.n2141 VDD.n2140 0.0445515
R33580 VDD.n8069 VDD.n8068 0.0440678
R33581 VDD.n8081 VDD.n8080 0.0436757
R33582 VDD.n8085 VDD.n8084 0.0436757
R33583 VDD.n2143 VDD.n2127 0.0433141
R33584 VDD.n2144 VDD.n2127 0.0433141
R33585 VDD.n2145 VDD.n2125 0.0433141
R33586 VDD.n8074 VDD.n2126 0.0433141
R33587 VDD.n8071 VDD.n2126 0.0433141
R33588 VDD.n8071 VDD.n8070 0.0433141
R33589 VDD.n8070 VDD.n8069 0.0433141
R33590 VDD.n2143 VDD.n2142 0.0430669
R33591 VDD.n7890 VDD.n7887 0.0430647
R33592 VDD.n7910 VDD.n7909 0.0428653
R33593 VDD.n7945 VDD.n7944 0.0417941
R33594 VDD.n8050 VDD.n8049 0.0417941
R33595 VDD.n1662 VDD.n1661 0.0416398
R33596 VDD.n1643 VDD.n1642 0.0416398
R33597 VDD.n1592 VDD.n1576 0.0416398
R33598 VDD.n1592 VDD.n1591 0.0416398
R33599 VDD.n7862 VDD.n7861 0.0416007
R33600 VDD.n7947 VDD.n7946 0.0415824
R33601 VDD.n7959 VDD.n2204 0.0413899
R33602 VDD.n2295 VDD.n2294 0.041314
R33603 VDD.n7839 VDD.n7838 0.041314
R33604 VDD.n2387 VDD.n2386 0.041314
R33605 VDD.n7830 VDD.n7829 0.041314
R33606 VDD.n7825 VDD.n7824 0.041314
R33607 VDD.n5216 VDD.n2423 0.0410752
R33608 VDD.n5215 VDD.n2422 0.0410752
R33609 VDD.n5214 VDD.n2421 0.0410752
R33610 VDD.n5213 VDD.n2420 0.0410752
R33611 VDD.n5212 VDD.n2419 0.0410752
R33612 VDD.n5211 VDD.n2418 0.0410752
R33613 VDD.n5210 VDD.n2417 0.0410752
R33614 VDD.n5209 VDD.n2416 0.0410752
R33615 VDD.n5208 VDD.n2415 0.0410752
R33616 VDD.n5207 VDD.n2414 0.0410752
R33617 VDD.n5206 VDD.n2413 0.0410752
R33618 VDD.n5205 VDD.n2412 0.0410752
R33619 VDD.n4597 VDD.n4596 0.0410752
R33620 VDD.n5217 VDD.n2423 0.0410752
R33621 VDD.n5216 VDD.n2422 0.0410752
R33622 VDD.n5215 VDD.n2421 0.0410752
R33623 VDD.n5214 VDD.n2420 0.0410752
R33624 VDD.n5213 VDD.n2419 0.0410752
R33625 VDD.n5212 VDD.n2418 0.0410752
R33626 VDD.n5211 VDD.n2417 0.0410752
R33627 VDD.n5210 VDD.n2416 0.0410752
R33628 VDD.n5209 VDD.n2415 0.0410752
R33629 VDD.n5208 VDD.n2414 0.0410752
R33630 VDD.n5207 VDD.n2413 0.0410752
R33631 VDD.n5206 VDD.n2412 0.0410752
R33632 VDD.n5203 VDD.n4596 0.0410752
R33633 VDD.n12446 VDD.n191 0.0410752
R33634 VDD.n12442 VDD.n192 0.0410752
R33635 VDD.n12443 VDD.n193 0.0410752
R33636 VDD.n9188 VDD.n9187 0.0410752
R33637 VDD.n9190 VDD.n9189 0.0410752
R33638 VDD.n9192 VDD.n9191 0.0410752
R33639 VDD.n9194 VDD.n9193 0.0410752
R33640 VDD.n9196 VDD.n9195 0.0410752
R33641 VDD.n9198 VDD.n9197 0.0410752
R33642 VDD.n9199 VDD.n9198 0.0410752
R33643 VDD.n9189 VDD.n9188 0.0410752
R33644 VDD.n9191 VDD.n9190 0.0410752
R33645 VDD.n9193 VDD.n9192 0.0410752
R33646 VDD.n9195 VDD.n9194 0.0410752
R33647 VDD.n9197 VDD.n9196 0.0410752
R33648 VDD.n12444 VDD.n193 0.0410752
R33649 VDD.n12443 VDD.n192 0.0410752
R33650 VDD.n12442 VDD.n191 0.0410752
R33651 VDD.n2145 VDD.n2144 0.040902
R33652 VDD.n1480 VDD.n1477 0.0404831
R33653 VDD.n1611 VDD.n1610 0.0404831
R33654 VDD.n1610 VDD.n1609 0.0404831
R33655 VDD.n1480 VDD.n1478 0.0404831
R33656 VDD.n5200 VDD.n4598 0.04025
R33657 VDD.n5196 VDD.n4598 0.04025
R33658 VDD.n5196 VDD.n5195 0.04025
R33659 VDD.n5195 VDD.n5194 0.04025
R33660 VDD.n5194 VDD.n4601 0.04025
R33661 VDD.n5190 VDD.n4601 0.04025
R33662 VDD.n5190 VDD.n5189 0.04025
R33663 VDD.n5189 VDD.n5188 0.04025
R33664 VDD.n5188 VDD.n4603 0.04025
R33665 VDD.n5184 VDD.n4603 0.04025
R33666 VDD.n5184 VDD.n5183 0.04025
R33667 VDD.n5183 VDD.n5182 0.04025
R33668 VDD.n5182 VDD.n4605 0.04025
R33669 VDD.n5178 VDD.n4605 0.04025
R33670 VDD.n5178 VDD.n5177 0.04025
R33671 VDD.n5177 VDD.n5176 0.04025
R33672 VDD.n5176 VDD.n4607 0.04025
R33673 VDD.n5172 VDD.n4607 0.04025
R33674 VDD.n5172 VDD.n5171 0.04025
R33675 VDD.n5171 VDD.n5170 0.04025
R33676 VDD.n5170 VDD.n4609 0.04025
R33677 VDD.n5166 VDD.n4609 0.04025
R33678 VDD.n5166 VDD.n5165 0.04025
R33679 VDD.n5165 VDD.n5164 0.04025
R33680 VDD.n5164 VDD.n4611 0.04025
R33681 VDD.n5160 VDD.n4611 0.04025
R33682 VDD.n5160 VDD.n5159 0.04025
R33683 VDD.n5159 VDD.n5158 0.04025
R33684 VDD.n5158 VDD.n4613 0.04025
R33685 VDD.n5154 VDD.n4613 0.04025
R33686 VDD.n5154 VDD.n5153 0.04025
R33687 VDD.n5153 VDD.n5152 0.04025
R33688 VDD.n5152 VDD.n4615 0.04025
R33689 VDD.n5148 VDD.n4615 0.04025
R33690 VDD.n5148 VDD.n5147 0.04025
R33691 VDD.n5147 VDD.n5146 0.04025
R33692 VDD.n5146 VDD.n4617 0.04025
R33693 VDD.n5142 VDD.n4617 0.04025
R33694 VDD.n5142 VDD.n5141 0.04025
R33695 VDD.n5141 VDD.n5140 0.04025
R33696 VDD.n5140 VDD.n4619 0.04025
R33697 VDD.n5136 VDD.n4619 0.04025
R33698 VDD.n5136 VDD.n5135 0.04025
R33699 VDD.n5135 VDD.n5134 0.04025
R33700 VDD.n5134 VDD.n4621 0.04025
R33701 VDD.n5130 VDD.n4621 0.04025
R33702 VDD.n5130 VDD.n5129 0.04025
R33703 VDD.n5129 VDD.n5128 0.04025
R33704 VDD.n5128 VDD.n4623 0.04025
R33705 VDD.n5124 VDD.n4623 0.04025
R33706 VDD.n5124 VDD.n5123 0.04025
R33707 VDD.n5123 VDD.n5122 0.04025
R33708 VDD.n5122 VDD.n4625 0.04025
R33709 VDD.n5118 VDD.n4625 0.04025
R33710 VDD.n5118 VDD.n5117 0.04025
R33711 VDD.n5117 VDD.n5116 0.04025
R33712 VDD.n5116 VDD.n4627 0.04025
R33713 VDD.n5112 VDD.n4627 0.04025
R33714 VDD.n5112 VDD.n5111 0.04025
R33715 VDD.n5111 VDD.n5110 0.04025
R33716 VDD.n5110 VDD.n4629 0.04025
R33717 VDD.n5106 VDD.n4629 0.04025
R33718 VDD.n5106 VDD.n5105 0.04025
R33719 VDD.n5105 VDD.n5104 0.04025
R33720 VDD.n5104 VDD.n4631 0.04025
R33721 VDD.n5100 VDD.n4631 0.04025
R33722 VDD.n5100 VDD.n5099 0.04025
R33723 VDD.n5099 VDD.n5098 0.04025
R33724 VDD.n5098 VDD.n4633 0.04025
R33725 VDD.n5094 VDD.n4633 0.04025
R33726 VDD.n5094 VDD.n5093 0.04025
R33727 VDD.n5093 VDD.n5092 0.04025
R33728 VDD.n5092 VDD.n4635 0.04025
R33729 VDD.n5088 VDD.n4635 0.04025
R33730 VDD.n5088 VDD.n5087 0.04025
R33731 VDD.n5087 VDD.n5086 0.04025
R33732 VDD.n5086 VDD.n4637 0.04025
R33733 VDD.n5082 VDD.n4637 0.04025
R33734 VDD.n5082 VDD.n5081 0.04025
R33735 VDD.n5081 VDD.n5080 0.04025
R33736 VDD.n5080 VDD.n4639 0.04025
R33737 VDD.n5076 VDD.n4639 0.04025
R33738 VDD.n5076 VDD.n5075 0.04025
R33739 VDD.n5075 VDD.n5074 0.04025
R33740 VDD.n5074 VDD.n4641 0.04025
R33741 VDD.n5070 VDD.n4641 0.04025
R33742 VDD.n5070 VDD.n5069 0.04025
R33743 VDD.n5069 VDD.n5068 0.04025
R33744 VDD.n5068 VDD.n4643 0.04025
R33745 VDD.n5064 VDD.n4643 0.04025
R33746 VDD.n5064 VDD.n5063 0.04025
R33747 VDD.n5063 VDD.n5062 0.04025
R33748 VDD.n5062 VDD.n4645 0.04025
R33749 VDD.n5058 VDD.n4645 0.04025
R33750 VDD.n5058 VDD.n5057 0.04025
R33751 VDD.n5057 VDD.n5056 0.04025
R33752 VDD.n5056 VDD.n4647 0.04025
R33753 VDD.n5052 VDD.n4647 0.04025
R33754 VDD.n5052 VDD.n5051 0.04025
R33755 VDD.n5051 VDD.n5050 0.04025
R33756 VDD.n5050 VDD.n4649 0.04025
R33757 VDD.n5046 VDD.n4649 0.04025
R33758 VDD.n5046 VDD.n5045 0.04025
R33759 VDD.n5045 VDD.n5044 0.04025
R33760 VDD.n5044 VDD.n4651 0.04025
R33761 VDD.n5040 VDD.n4651 0.04025
R33762 VDD.n5040 VDD.n5039 0.04025
R33763 VDD.n5039 VDD.n5038 0.04025
R33764 VDD.n5038 VDD.n4653 0.04025
R33765 VDD.n5034 VDD.n4653 0.04025
R33766 VDD.n5034 VDD.n5033 0.04025
R33767 VDD.n5033 VDD.n5032 0.04025
R33768 VDD.n5032 VDD.n4655 0.04025
R33769 VDD.n5028 VDD.n4655 0.04025
R33770 VDD.n5028 VDD.n5027 0.04025
R33771 VDD.n5027 VDD.n5026 0.04025
R33772 VDD.n5026 VDD.n4657 0.04025
R33773 VDD.n5022 VDD.n4657 0.04025
R33774 VDD.n5022 VDD.n5021 0.04025
R33775 VDD.n5021 VDD.n5020 0.04025
R33776 VDD.n5020 VDD.n4659 0.04025
R33777 VDD.n5016 VDD.n4659 0.04025
R33778 VDD.n5016 VDD.n5015 0.04025
R33779 VDD.n5015 VDD.n5014 0.04025
R33780 VDD.n5014 VDD.n4661 0.04025
R33781 VDD.n5010 VDD.n4661 0.04025
R33782 VDD.n5010 VDD.n5009 0.04025
R33783 VDD.n5009 VDD.n5008 0.04025
R33784 VDD.n5008 VDD.n4663 0.04025
R33785 VDD.n5004 VDD.n4663 0.04025
R33786 VDD.n5004 VDD.n5003 0.04025
R33787 VDD.n5003 VDD.n5002 0.04025
R33788 VDD.n5002 VDD.n4665 0.04025
R33789 VDD.n4998 VDD.n4665 0.04025
R33790 VDD.n4998 VDD.n4997 0.04025
R33791 VDD.n4997 VDD.n4996 0.04025
R33792 VDD.n4996 VDD.n4667 0.04025
R33793 VDD.n4992 VDD.n4667 0.04025
R33794 VDD.n4992 VDD.n4991 0.04025
R33795 VDD.n4991 VDD.n4990 0.04025
R33796 VDD.n4990 VDD.n4669 0.04025
R33797 VDD.n4986 VDD.n4669 0.04025
R33798 VDD.n4986 VDD.n4985 0.04025
R33799 VDD.n4985 VDD.n4984 0.04025
R33800 VDD.n4984 VDD.n4671 0.04025
R33801 VDD.n4980 VDD.n4671 0.04025
R33802 VDD.n4980 VDD.n4979 0.04025
R33803 VDD.n4979 VDD.n4978 0.04025
R33804 VDD.n4978 VDD.n4673 0.04025
R33805 VDD.n4974 VDD.n4673 0.04025
R33806 VDD.n4974 VDD.n4973 0.04025
R33807 VDD.n4973 VDD.n4972 0.04025
R33808 VDD.n4972 VDD.n4675 0.04025
R33809 VDD.n4968 VDD.n4675 0.04025
R33810 VDD.n4968 VDD.n4967 0.04025
R33811 VDD.n4967 VDD.n4966 0.04025
R33812 VDD.n4966 VDD.n4677 0.04025
R33813 VDD.n4962 VDD.n4677 0.04025
R33814 VDD.n4962 VDD.n4961 0.04025
R33815 VDD.n4961 VDD.n4960 0.04025
R33816 VDD.n4960 VDD.n4679 0.04025
R33817 VDD.n4956 VDD.n4679 0.04025
R33818 VDD.n4956 VDD.n4955 0.04025
R33819 VDD.n4955 VDD.n4954 0.04025
R33820 VDD.n4954 VDD.n4681 0.04025
R33821 VDD.n4950 VDD.n4681 0.04025
R33822 VDD.n4950 VDD.n4949 0.04025
R33823 VDD.n4949 VDD.n4948 0.04025
R33824 VDD.n4948 VDD.n4683 0.04025
R33825 VDD.n4944 VDD.n4683 0.04025
R33826 VDD.n4944 VDD.n4943 0.04025
R33827 VDD.n4943 VDD.n4942 0.04025
R33828 VDD.n4942 VDD.n4685 0.04025
R33829 VDD.n4938 VDD.n4685 0.04025
R33830 VDD.n4938 VDD.n4937 0.04025
R33831 VDD.n4937 VDD.n4936 0.04025
R33832 VDD.n4936 VDD.n4687 0.04025
R33833 VDD.n4932 VDD.n4687 0.04025
R33834 VDD.n4932 VDD.n4931 0.04025
R33835 VDD.n4931 VDD.n4930 0.04025
R33836 VDD.n4930 VDD.n4689 0.04025
R33837 VDD.n4926 VDD.n4689 0.04025
R33838 VDD.n4926 VDD.n4925 0.04025
R33839 VDD.n4925 VDD.n4924 0.04025
R33840 VDD.n4924 VDD.n4691 0.04025
R33841 VDD.n4920 VDD.n4691 0.04025
R33842 VDD.n4920 VDD.n4919 0.04025
R33843 VDD.n4919 VDD.n4918 0.04025
R33844 VDD.n4918 VDD.n4693 0.04025
R33845 VDD.n4914 VDD.n4693 0.04025
R33846 VDD.n4914 VDD.n4913 0.04025
R33847 VDD.n4913 VDD.n4912 0.04025
R33848 VDD.n4912 VDD.n4695 0.04025
R33849 VDD.n4908 VDD.n4695 0.04025
R33850 VDD.n4908 VDD.n4907 0.04025
R33851 VDD.n4907 VDD.n4906 0.04025
R33852 VDD.n4902 VDD.n4697 0.04025
R33853 VDD.n4902 VDD.n4901 0.04025
R33854 VDD.n4901 VDD.n4900 0.04025
R33855 VDD.n4900 VDD.n4699 0.04025
R33856 VDD.n4896 VDD.n4699 0.04025
R33857 VDD.n4896 VDD.n4895 0.04025
R33858 VDD.n4895 VDD.n4894 0.04025
R33859 VDD.n4894 VDD.n4701 0.04025
R33860 VDD.n4890 VDD.n4701 0.04025
R33861 VDD.n4890 VDD.n4889 0.04025
R33862 VDD.n4889 VDD.n4888 0.04025
R33863 VDD.n4888 VDD.n4703 0.04025
R33864 VDD.n4884 VDD.n4703 0.04025
R33865 VDD.n4884 VDD.n4883 0.04025
R33866 VDD.n4883 VDD.n4882 0.04025
R33867 VDD.n4882 VDD.n4705 0.04025
R33868 VDD.n4878 VDD.n4705 0.04025
R33869 VDD.n4878 VDD.n4877 0.04025
R33870 VDD.n4877 VDD.n4876 0.04025
R33871 VDD.n4876 VDD.n4707 0.04025
R33872 VDD.n4872 VDD.n4707 0.04025
R33873 VDD.n4872 VDD.n4871 0.04025
R33874 VDD.n4871 VDD.n4870 0.04025
R33875 VDD.n4870 VDD.n4709 0.04025
R33876 VDD.n4866 VDD.n4709 0.04025
R33877 VDD.n4866 VDD.n4865 0.04025
R33878 VDD.n4865 VDD.n4864 0.04025
R33879 VDD.n4864 VDD.n4711 0.04025
R33880 VDD.n4860 VDD.n4711 0.04025
R33881 VDD.n4860 VDD.n4859 0.04025
R33882 VDD.n4859 VDD.n4858 0.04025
R33883 VDD.n4858 VDD.n4713 0.04025
R33884 VDD.n4854 VDD.n4713 0.04025
R33885 VDD.n4854 VDD.n4853 0.04025
R33886 VDD.n4853 VDD.n4852 0.04025
R33887 VDD.n4852 VDD.n4715 0.04025
R33888 VDD.n4848 VDD.n4715 0.04025
R33889 VDD.n4848 VDD.n4847 0.04025
R33890 VDD.n4847 VDD.n4846 0.04025
R33891 VDD.n4846 VDD.n4717 0.04025
R33892 VDD.n4842 VDD.n4717 0.04025
R33893 VDD.n4842 VDD.n4841 0.04025
R33894 VDD.n4841 VDD.n4840 0.04025
R33895 VDD.n4840 VDD.n4719 0.04025
R33896 VDD.n4836 VDD.n4719 0.04025
R33897 VDD.n4836 VDD.n4835 0.04025
R33898 VDD.n4835 VDD.n4834 0.04025
R33899 VDD.n4834 VDD.n4721 0.04025
R33900 VDD.n4830 VDD.n4721 0.04025
R33901 VDD.n4830 VDD.n4829 0.04025
R33902 VDD.n4829 VDD.n4828 0.04025
R33903 VDD.n4828 VDD.n4723 0.04025
R33904 VDD.n4824 VDD.n4723 0.04025
R33905 VDD.n4824 VDD.n4823 0.04025
R33906 VDD.n4823 VDD.n4822 0.04025
R33907 VDD.n4822 VDD.n4725 0.04025
R33908 VDD.n4818 VDD.n4725 0.04025
R33909 VDD.n4818 VDD.n4817 0.04025
R33910 VDD.n4817 VDD.n4816 0.04025
R33911 VDD.n4816 VDD.n4727 0.04025
R33912 VDD.n4812 VDD.n4727 0.04025
R33913 VDD.n4812 VDD.n4811 0.04025
R33914 VDD.n4811 VDD.n4810 0.04025
R33915 VDD.n4810 VDD.n4729 0.04025
R33916 VDD.n4806 VDD.n4729 0.04025
R33917 VDD.n4806 VDD.n4805 0.04025
R33918 VDD.n4805 VDD.n4804 0.04025
R33919 VDD.n4804 VDD.n4731 0.04025
R33920 VDD.n4800 VDD.n4731 0.04025
R33921 VDD.n4800 VDD.n4799 0.04025
R33922 VDD.n4799 VDD.n4798 0.04025
R33923 VDD.n4798 VDD.n4733 0.04025
R33924 VDD.n4794 VDD.n4733 0.04025
R33925 VDD.n4794 VDD.n4793 0.04025
R33926 VDD.n4793 VDD.n4792 0.04025
R33927 VDD.n4792 VDD.n4735 0.04025
R33928 VDD.n4788 VDD.n4735 0.04025
R33929 VDD.n4788 VDD.n4787 0.04025
R33930 VDD.n4787 VDD.n4786 0.04025
R33931 VDD.n4786 VDD.n4737 0.04025
R33932 VDD.n4782 VDD.n4737 0.04025
R33933 VDD.n4782 VDD.n4781 0.04025
R33934 VDD.n4781 VDD.n4780 0.04025
R33935 VDD.n4780 VDD.n4739 0.04025
R33936 VDD.n4776 VDD.n4739 0.04025
R33937 VDD.n4776 VDD.n4775 0.04025
R33938 VDD.n4775 VDD.n4774 0.04025
R33939 VDD.n4774 VDD.n4741 0.04025
R33940 VDD.n4770 VDD.n4741 0.04025
R33941 VDD.n4770 VDD.n4769 0.04025
R33942 VDD.n4769 VDD.n4768 0.04025
R33943 VDD.n4768 VDD.n4743 0.04025
R33944 VDD.n4764 VDD.n4743 0.04025
R33945 VDD.n4764 VDD.n4763 0.04025
R33946 VDD.n4763 VDD.n4762 0.04025
R33947 VDD.n4762 VDD.n4745 0.04025
R33948 VDD.n4758 VDD.n4745 0.04025
R33949 VDD.n4758 VDD.n4757 0.04025
R33950 VDD.n4757 VDD.n4756 0.04025
R33951 VDD.n4756 VDD.n4747 0.04025
R33952 VDD.n4752 VDD.n4747 0.04025
R33953 VDD.n4752 VDD.n4751 0.04025
R33954 VDD.n4751 VDD.n4750 0.04025
R33955 VDD.n4750 VDD.n2242 0.04025
R33956 VDD.n7682 VDD.n7681 0.04025
R33957 VDD.n7681 VDD.n7178 0.04025
R33958 VDD.n7677 VDD.n7178 0.04025
R33959 VDD.n7677 VDD.n7676 0.04025
R33960 VDD.n7676 VDD.n7675 0.04025
R33961 VDD.n7675 VDD.n7180 0.04025
R33962 VDD.n7671 VDD.n7180 0.04025
R33963 VDD.n7671 VDD.n7670 0.04025
R33964 VDD.n7670 VDD.n7669 0.04025
R33965 VDD.n7669 VDD.n7182 0.04025
R33966 VDD.n7665 VDD.n7182 0.04025
R33967 VDD.n7665 VDD.n7664 0.04025
R33968 VDD.n7664 VDD.n7663 0.04025
R33969 VDD.n7663 VDD.n7184 0.04025
R33970 VDD.n7659 VDD.n7184 0.04025
R33971 VDD.n7659 VDD.n7658 0.04025
R33972 VDD.n7658 VDD.n7657 0.04025
R33973 VDD.n7657 VDD.n7186 0.04025
R33974 VDD.n7653 VDD.n7186 0.04025
R33975 VDD.n7653 VDD.n7652 0.04025
R33976 VDD.n7652 VDD.n7651 0.04025
R33977 VDD.n7651 VDD.n7188 0.04025
R33978 VDD.n7647 VDD.n7188 0.04025
R33979 VDD.n7647 VDD.n7646 0.04025
R33980 VDD.n7646 VDD.n7645 0.04025
R33981 VDD.n7645 VDD.n7190 0.04025
R33982 VDD.n7641 VDD.n7190 0.04025
R33983 VDD.n7641 VDD.n7640 0.04025
R33984 VDD.n7640 VDD.n7639 0.04025
R33985 VDD.n7639 VDD.n7192 0.04025
R33986 VDD.n7635 VDD.n7192 0.04025
R33987 VDD.n7635 VDD.n7634 0.04025
R33988 VDD.n7634 VDD.n7633 0.04025
R33989 VDD.n7633 VDD.n7194 0.04025
R33990 VDD.n7629 VDD.n7194 0.04025
R33991 VDD.n7629 VDD.n7628 0.04025
R33992 VDD.n7628 VDD.n7627 0.04025
R33993 VDD.n7627 VDD.n7196 0.04025
R33994 VDD.n7623 VDD.n7196 0.04025
R33995 VDD.n7623 VDD.n7622 0.04025
R33996 VDD.n7622 VDD.n7621 0.04025
R33997 VDD.n7621 VDD.n7198 0.04025
R33998 VDD.n7617 VDD.n7198 0.04025
R33999 VDD.n7617 VDD.n7616 0.04025
R34000 VDD.n7616 VDD.n7615 0.04025
R34001 VDD.n7615 VDD.n7200 0.04025
R34002 VDD.n7611 VDD.n7200 0.04025
R34003 VDD.n7611 VDD.n7610 0.04025
R34004 VDD.n7610 VDD.n7609 0.04025
R34005 VDD.n7609 VDD.n7202 0.04025
R34006 VDD.n7605 VDD.n7202 0.04025
R34007 VDD.n7605 VDD.n7604 0.04025
R34008 VDD.n7604 VDD.n7603 0.04025
R34009 VDD.n7603 VDD.n7204 0.04025
R34010 VDD.n7599 VDD.n7204 0.04025
R34011 VDD.n7599 VDD.n7598 0.04025
R34012 VDD.n7598 VDD.n7597 0.04025
R34013 VDD.n7597 VDD.n7206 0.04025
R34014 VDD.n7593 VDD.n7206 0.04025
R34015 VDD.n7593 VDD.n7592 0.04025
R34016 VDD.n7592 VDD.n7591 0.04025
R34017 VDD.n7591 VDD.n7208 0.04025
R34018 VDD.n7587 VDD.n7208 0.04025
R34019 VDD.n7587 VDD.n7586 0.04025
R34020 VDD.n7586 VDD.n7585 0.04025
R34021 VDD.n7585 VDD.n7210 0.04025
R34022 VDD.n7581 VDD.n7210 0.04025
R34023 VDD.n7581 VDD.n7580 0.04025
R34024 VDD.n7580 VDD.n7579 0.04025
R34025 VDD.n7579 VDD.n7212 0.04025
R34026 VDD.n7575 VDD.n7212 0.04025
R34027 VDD.n7575 VDD.n7574 0.04025
R34028 VDD.n7574 VDD.n7573 0.04025
R34029 VDD.n7573 VDD.n7214 0.04025
R34030 VDD.n7569 VDD.n7214 0.04025
R34031 VDD.n7569 VDD.n7568 0.04025
R34032 VDD.n7568 VDD.n7567 0.04025
R34033 VDD.n7567 VDD.n7216 0.04025
R34034 VDD.n7563 VDD.n7216 0.04025
R34035 VDD.n7563 VDD.n7562 0.04025
R34036 VDD.n7562 VDD.n7561 0.04025
R34037 VDD.n7561 VDD.n7218 0.04025
R34038 VDD.n7557 VDD.n7218 0.04025
R34039 VDD.n7557 VDD.n7556 0.04025
R34040 VDD.n7556 VDD.n7555 0.04025
R34041 VDD.n7555 VDD.n7220 0.04025
R34042 VDD.n7551 VDD.n7220 0.04025
R34043 VDD.n7551 VDD.n7550 0.04025
R34044 VDD.n7550 VDD.n7549 0.04025
R34045 VDD.n7549 VDD.n7222 0.04025
R34046 VDD.n7545 VDD.n7222 0.04025
R34047 VDD.n7545 VDD.n7544 0.04025
R34048 VDD.n7544 VDD.n7543 0.04025
R34049 VDD.n7543 VDD.n7224 0.04025
R34050 VDD.n7539 VDD.n7224 0.04025
R34051 VDD.n7539 VDD.n7538 0.04025
R34052 VDD.n7538 VDD.n7537 0.04025
R34053 VDD.n7537 VDD.n7226 0.04025
R34054 VDD.n7533 VDD.n7226 0.04025
R34055 VDD.n7533 VDD.n7532 0.04025
R34056 VDD.n7532 VDD.n7531 0.04025
R34057 VDD.n7531 VDD.n7228 0.04025
R34058 VDD.n7527 VDD.n7228 0.04025
R34059 VDD.n7527 VDD.n7526 0.04025
R34060 VDD.n7526 VDD.n7525 0.04025
R34061 VDD.n7525 VDD.n7230 0.04025
R34062 VDD.n7521 VDD.n7230 0.04025
R34063 VDD.n7521 VDD.n7520 0.04025
R34064 VDD.n7520 VDD.n7519 0.04025
R34065 VDD.n7519 VDD.n7232 0.04025
R34066 VDD.n7515 VDD.n7232 0.04025
R34067 VDD.n7515 VDD.n7514 0.04025
R34068 VDD.n7514 VDD.n7513 0.04025
R34069 VDD.n7513 VDD.n7234 0.04025
R34070 VDD.n7509 VDD.n7234 0.04025
R34071 VDD.n7509 VDD.n7508 0.04025
R34072 VDD.n7508 VDD.n7507 0.04025
R34073 VDD.n7507 VDD.n7236 0.04025
R34074 VDD.n7503 VDD.n7236 0.04025
R34075 VDD.n7503 VDD.n7502 0.04025
R34076 VDD.n7502 VDD.n7501 0.04025
R34077 VDD.n7501 VDD.n7238 0.04025
R34078 VDD.n7497 VDD.n7238 0.04025
R34079 VDD.n7497 VDD.n7496 0.04025
R34080 VDD.n7496 VDD.n7495 0.04025
R34081 VDD.n7495 VDD.n7240 0.04025
R34082 VDD.n7491 VDD.n7240 0.04025
R34083 VDD.n7491 VDD.n7490 0.04025
R34084 VDD.n7490 VDD.n7489 0.04025
R34085 VDD.n7489 VDD.n7242 0.04025
R34086 VDD.n7485 VDD.n7242 0.04025
R34087 VDD.n7485 VDD.n7484 0.04025
R34088 VDD.n7484 VDD.n7483 0.04025
R34089 VDD.n7483 VDD.n7244 0.04025
R34090 VDD.n7479 VDD.n7244 0.04025
R34091 VDD.n7479 VDD.n7478 0.04025
R34092 VDD.n7478 VDD.n7477 0.04025
R34093 VDD.n7477 VDD.n7246 0.04025
R34094 VDD.n7473 VDD.n7246 0.04025
R34095 VDD.n7473 VDD.n7472 0.04025
R34096 VDD.n7472 VDD.n7471 0.04025
R34097 VDD.n7471 VDD.n7248 0.04025
R34098 VDD.n7467 VDD.n7248 0.04025
R34099 VDD.n7467 VDD.n7466 0.04025
R34100 VDD.n7466 VDD.n7465 0.04025
R34101 VDD.n7465 VDD.n7250 0.04025
R34102 VDD.n7461 VDD.n7250 0.04025
R34103 VDD.n7461 VDD.n7460 0.04025
R34104 VDD.n7460 VDD.n7459 0.04025
R34105 VDD.n7459 VDD.n7252 0.04025
R34106 VDD.n7455 VDD.n7252 0.04025
R34107 VDD.n7455 VDD.n7454 0.04025
R34108 VDD.n7454 VDD.n7453 0.04025
R34109 VDD.n7453 VDD.n7254 0.04025
R34110 VDD.n7449 VDD.n7254 0.04025
R34111 VDD.n7449 VDD.n7448 0.04025
R34112 VDD.n7448 VDD.n7447 0.04025
R34113 VDD.n7447 VDD.n7256 0.04025
R34114 VDD.n7443 VDD.n7256 0.04025
R34115 VDD.n7443 VDD.n7442 0.04025
R34116 VDD.n7442 VDD.n7441 0.04025
R34117 VDD.n7441 VDD.n7258 0.04025
R34118 VDD.n7437 VDD.n7258 0.04025
R34119 VDD.n7437 VDD.n7436 0.04025
R34120 VDD.n7436 VDD.n7435 0.04025
R34121 VDD.n7435 VDD.n7260 0.04025
R34122 VDD.n7431 VDD.n7260 0.04025
R34123 VDD.n7431 VDD.n7430 0.04025
R34124 VDD.n7430 VDD.n7429 0.04025
R34125 VDD.n7429 VDD.n7262 0.04025
R34126 VDD.n7425 VDD.n7262 0.04025
R34127 VDD.n7425 VDD.n7424 0.04025
R34128 VDD.n7424 VDD.n7423 0.04025
R34129 VDD.n7423 VDD.n7264 0.04025
R34130 VDD.n7419 VDD.n7264 0.04025
R34131 VDD.n7419 VDD.n7418 0.04025
R34132 VDD.n7418 VDD.n7417 0.04025
R34133 VDD.n7417 VDD.n7266 0.04025
R34134 VDD.n7413 VDD.n7266 0.04025
R34135 VDD.n7413 VDD.n7412 0.04025
R34136 VDD.n7412 VDD.n7411 0.04025
R34137 VDD.n7411 VDD.n7268 0.04025
R34138 VDD.n7407 VDD.n7268 0.04025
R34139 VDD.n7407 VDD.n7406 0.04025
R34140 VDD.n7406 VDD.n7405 0.04025
R34141 VDD.n7405 VDD.n7270 0.04025
R34142 VDD.n7401 VDD.n7270 0.04025
R34143 VDD.n7401 VDD.n7400 0.04025
R34144 VDD.n7400 VDD.n7399 0.04025
R34145 VDD.n7399 VDD.n7272 0.04025
R34146 VDD.n7395 VDD.n7272 0.04025
R34147 VDD.n7395 VDD.n7394 0.04025
R34148 VDD.n7394 VDD.n7393 0.04025
R34149 VDD.n7393 VDD.n7274 0.04025
R34150 VDD.n7389 VDD.n7274 0.04025
R34151 VDD.n7389 VDD.n7388 0.04025
R34152 VDD.n7388 VDD.n7387 0.04025
R34153 VDD.n7387 VDD.n7276 0.04025
R34154 VDD.n7383 VDD.n7276 0.04025
R34155 VDD.n7383 VDD.n7382 0.04025
R34156 VDD.n7382 VDD.n7381 0.04025
R34157 VDD.n7381 VDD.n7278 0.04025
R34158 VDD.n7377 VDD.n7278 0.04025
R34159 VDD.n7377 VDD.n7376 0.04025
R34160 VDD.n7376 VDD.n7375 0.04025
R34161 VDD.n7375 VDD.n7280 0.04025
R34162 VDD.n7371 VDD.n7280 0.04025
R34163 VDD.n7371 VDD.n7370 0.04025
R34164 VDD.n7370 VDD.n7369 0.04025
R34165 VDD.n7369 VDD.n7282 0.04025
R34166 VDD.n7365 VDD.n7282 0.04025
R34167 VDD.n7365 VDD.n7364 0.04025
R34168 VDD.n7364 VDD.n7363 0.04025
R34169 VDD.n7363 VDD.n7284 0.04025
R34170 VDD.n7359 VDD.n7284 0.04025
R34171 VDD.n7359 VDD.n7358 0.04025
R34172 VDD.n7358 VDD.n7357 0.04025
R34173 VDD.n7357 VDD.n7286 0.04025
R34174 VDD.n7353 VDD.n7286 0.04025
R34175 VDD.n7353 VDD.n7352 0.04025
R34176 VDD.n7352 VDD.n7351 0.04025
R34177 VDD.n7351 VDD.n7288 0.04025
R34178 VDD.n7347 VDD.n7288 0.04025
R34179 VDD.n7347 VDD.n7346 0.04025
R34180 VDD.n7346 VDD.n7345 0.04025
R34181 VDD.n7345 VDD.n7290 0.04025
R34182 VDD.n7341 VDD.n7290 0.04025
R34183 VDD.n7341 VDD.n7340 0.04025
R34184 VDD.n7340 VDD.n7339 0.04025
R34185 VDD.n7339 VDD.n7292 0.04025
R34186 VDD.n7335 VDD.n7292 0.04025
R34187 VDD.n7335 VDD.n7334 0.04025
R34188 VDD.n7334 VDD.n7333 0.04025
R34189 VDD.n7333 VDD.n7294 0.04025
R34190 VDD.n7329 VDD.n7294 0.04025
R34191 VDD.n7329 VDD.n7328 0.04025
R34192 VDD.n7328 VDD.n7327 0.04025
R34193 VDD.n7327 VDD.n7296 0.04025
R34194 VDD.n7323 VDD.n7296 0.04025
R34195 VDD.n7323 VDD.n7322 0.04025
R34196 VDD.n7322 VDD.n7321 0.04025
R34197 VDD.n7321 VDD.n7298 0.04025
R34198 VDD.n7317 VDD.n7298 0.04025
R34199 VDD.n7317 VDD.n7316 0.04025
R34200 VDD.n7316 VDD.n7315 0.04025
R34201 VDD.n7315 VDD.n7300 0.04025
R34202 VDD.n7311 VDD.n7300 0.04025
R34203 VDD.n7311 VDD.n7310 0.04025
R34204 VDD.n7310 VDD.n7309 0.04025
R34205 VDD.n10759 VDD.n8255 0.04025
R34206 VDD.n10755 VDD.n8255 0.04025
R34207 VDD.n10755 VDD.n10754 0.04025
R34208 VDD.n10754 VDD.n10753 0.04025
R34209 VDD.n10753 VDD.n8257 0.04025
R34210 VDD.n10749 VDD.n8257 0.04025
R34211 VDD.n10749 VDD.n10748 0.04025
R34212 VDD.n10748 VDD.n10747 0.04025
R34213 VDD.n10747 VDD.n8259 0.04025
R34214 VDD.n10743 VDD.n8259 0.04025
R34215 VDD.n10743 VDD.n10742 0.04025
R34216 VDD.n10742 VDD.n10741 0.04025
R34217 VDD.n10741 VDD.n8261 0.04025
R34218 VDD.n10737 VDD.n8261 0.04025
R34219 VDD.n10737 VDD.n10736 0.04025
R34220 VDD.n10736 VDD.n10735 0.04025
R34221 VDD.n10735 VDD.n8263 0.04025
R34222 VDD.n10731 VDD.n8263 0.04025
R34223 VDD.n10731 VDD.n10730 0.04025
R34224 VDD.n10730 VDD.n10729 0.04025
R34225 VDD.n10729 VDD.n8265 0.04025
R34226 VDD.n10725 VDD.n8265 0.04025
R34227 VDD.n10725 VDD.n10724 0.04025
R34228 VDD.n10724 VDD.n10723 0.04025
R34229 VDD.n10723 VDD.n8267 0.04025
R34230 VDD.n10719 VDD.n8267 0.04025
R34231 VDD.n10719 VDD.n10718 0.04025
R34232 VDD.n10718 VDD.n10717 0.04025
R34233 VDD.n10717 VDD.n8269 0.04025
R34234 VDD.n10713 VDD.n8269 0.04025
R34235 VDD.n10713 VDD.n10712 0.04025
R34236 VDD.n10712 VDD.n10711 0.04025
R34237 VDD.n10711 VDD.n8271 0.04025
R34238 VDD.n10707 VDD.n8271 0.04025
R34239 VDD.n10707 VDD.n10706 0.04025
R34240 VDD.n10706 VDD.n10705 0.04025
R34241 VDD.n10705 VDD.n8273 0.04025
R34242 VDD.n10701 VDD.n8273 0.04025
R34243 VDD.n10701 VDD.n10700 0.04025
R34244 VDD.n10700 VDD.n10699 0.04025
R34245 VDD.n10699 VDD.n8275 0.04025
R34246 VDD.n10695 VDD.n8275 0.04025
R34247 VDD.n10695 VDD.n10694 0.04025
R34248 VDD.n10694 VDD.n10693 0.04025
R34249 VDD.n10693 VDD.n8277 0.04025
R34250 VDD.n10689 VDD.n8277 0.04025
R34251 VDD.n10689 VDD.n10688 0.04025
R34252 VDD.n10688 VDD.n10687 0.04025
R34253 VDD.n10687 VDD.n8279 0.04025
R34254 VDD.n10683 VDD.n8279 0.04025
R34255 VDD.n10683 VDD.n10682 0.04025
R34256 VDD.n10682 VDD.n10681 0.04025
R34257 VDD.n10681 VDD.n8281 0.04025
R34258 VDD.n10677 VDD.n8281 0.04025
R34259 VDD.n10677 VDD.n10676 0.04025
R34260 VDD.n10676 VDD.n10675 0.04025
R34261 VDD.n10675 VDD.n8283 0.04025
R34262 VDD.n10671 VDD.n8283 0.04025
R34263 VDD.n10671 VDD.n10670 0.04025
R34264 VDD.n10670 VDD.n10669 0.04025
R34265 VDD.n10669 VDD.n8285 0.04025
R34266 VDD.n10665 VDD.n8285 0.04025
R34267 VDD.n10665 VDD.n10664 0.04025
R34268 VDD.n10664 VDD.n10663 0.04025
R34269 VDD.n10663 VDD.n8287 0.04025
R34270 VDD.n10659 VDD.n8287 0.04025
R34271 VDD.n10659 VDD.n10658 0.04025
R34272 VDD.n10658 VDD.n10657 0.04025
R34273 VDD.n10657 VDD.n8289 0.04025
R34274 VDD.n10653 VDD.n8289 0.04025
R34275 VDD.n10653 VDD.n10652 0.04025
R34276 VDD.n10652 VDD.n10651 0.04025
R34277 VDD.n10651 VDD.n8291 0.04025
R34278 VDD.n10647 VDD.n8291 0.04025
R34279 VDD.n10647 VDD.n10646 0.04025
R34280 VDD.n10646 VDD.n10645 0.04025
R34281 VDD.n10645 VDD.n8293 0.04025
R34282 VDD.n10641 VDD.n8293 0.04025
R34283 VDD.n10641 VDD.n10640 0.04025
R34284 VDD.n10640 VDD.n10639 0.04025
R34285 VDD.n10639 VDD.n8295 0.04025
R34286 VDD.n10635 VDD.n8295 0.04025
R34287 VDD.n10635 VDD.n10634 0.04025
R34288 VDD.n10634 VDD.n10633 0.04025
R34289 VDD.n10633 VDD.n8297 0.04025
R34290 VDD.n10629 VDD.n8297 0.04025
R34291 VDD.n10629 VDD.n10628 0.04025
R34292 VDD.n10628 VDD.n10627 0.04025
R34293 VDD.n10627 VDD.n8299 0.04025
R34294 VDD.n10623 VDD.n8299 0.04025
R34295 VDD.n10623 VDD.n10622 0.04025
R34296 VDD.n10622 VDD.n10621 0.04025
R34297 VDD.n10621 VDD.n8301 0.04025
R34298 VDD.n10617 VDD.n8301 0.04025
R34299 VDD.n10617 VDD.n10616 0.04025
R34300 VDD.n10616 VDD.n10615 0.04025
R34301 VDD.n10615 VDD.n8303 0.04025
R34302 VDD.n10611 VDD.n8303 0.04025
R34303 VDD.n10611 VDD.n10610 0.04025
R34304 VDD.n10610 VDD.n10609 0.04025
R34305 VDD.n10609 VDD.n8305 0.04025
R34306 VDD.n10605 VDD.n8305 0.04025
R34307 VDD.n10605 VDD.n10604 0.04025
R34308 VDD.n10604 VDD.n10603 0.04025
R34309 VDD.n10603 VDD.n8307 0.04025
R34310 VDD.n10599 VDD.n8307 0.04025
R34311 VDD.n10599 VDD.n10598 0.04025
R34312 VDD.n10598 VDD.n10597 0.04025
R34313 VDD.n10597 VDD.n8309 0.04025
R34314 VDD.n10593 VDD.n8309 0.04025
R34315 VDD.n10593 VDD.n10592 0.04025
R34316 VDD.n10592 VDD.n10591 0.04025
R34317 VDD.n10591 VDD.n8311 0.04025
R34318 VDD.n10587 VDD.n8311 0.04025
R34319 VDD.n10587 VDD.n10586 0.04025
R34320 VDD.n10586 VDD.n10585 0.04025
R34321 VDD.n10585 VDD.n8313 0.04025
R34322 VDD.n10581 VDD.n8313 0.04025
R34323 VDD.n10581 VDD.n10580 0.04025
R34324 VDD.n10580 VDD.n10579 0.04025
R34325 VDD.n10579 VDD.n8315 0.04025
R34326 VDD.n10575 VDD.n8315 0.04025
R34327 VDD.n10575 VDD.n10574 0.04025
R34328 VDD.n10574 VDD.n10573 0.04025
R34329 VDD.n10573 VDD.n8317 0.04025
R34330 VDD.n10569 VDD.n8317 0.04025
R34331 VDD.n10569 VDD.n10568 0.04025
R34332 VDD.n10568 VDD.n10567 0.04025
R34333 VDD.n10567 VDD.n8319 0.04025
R34334 VDD.n10563 VDD.n8319 0.04025
R34335 VDD.n10563 VDD.n10562 0.04025
R34336 VDD.n10562 VDD.n10561 0.04025
R34337 VDD.n10561 VDD.n8321 0.04025
R34338 VDD.n10557 VDD.n8321 0.04025
R34339 VDD.n10557 VDD.n10556 0.04025
R34340 VDD.n10556 VDD.n10555 0.04025
R34341 VDD.n10555 VDD.n8323 0.04025
R34342 VDD.n10551 VDD.n8323 0.04025
R34343 VDD.n10551 VDD.n10550 0.04025
R34344 VDD.n10550 VDD.n10549 0.04025
R34345 VDD.n10549 VDD.n8325 0.04025
R34346 VDD.n10545 VDD.n8325 0.04025
R34347 VDD.n10545 VDD.n10544 0.04025
R34348 VDD.n10544 VDD.n10543 0.04025
R34349 VDD.n10543 VDD.n8327 0.04025
R34350 VDD.n10539 VDD.n8327 0.04025
R34351 VDD.n10539 VDD.n10538 0.04025
R34352 VDD.n10538 VDD.n10537 0.04025
R34353 VDD.n10537 VDD.n8329 0.04025
R34354 VDD.n10533 VDD.n8329 0.04025
R34355 VDD.n10533 VDD.n10532 0.04025
R34356 VDD.n10532 VDD.n10531 0.04025
R34357 VDD.n10531 VDD.n8331 0.04025
R34358 VDD.n10527 VDD.n8331 0.04025
R34359 VDD.n10527 VDD.n10526 0.04025
R34360 VDD.n10526 VDD.n10525 0.04025
R34361 VDD.n10525 VDD.n8333 0.04025
R34362 VDD.n10521 VDD.n8333 0.04025
R34363 VDD.n10521 VDD.n10520 0.04025
R34364 VDD.n10520 VDD.n10519 0.04025
R34365 VDD.n10519 VDD.n8335 0.04025
R34366 VDD.n10515 VDD.n8335 0.04025
R34367 VDD.n10515 VDD.n10514 0.04025
R34368 VDD.n10514 VDD.n10513 0.04025
R34369 VDD.n10513 VDD.n8337 0.04025
R34370 VDD.n10509 VDD.n8337 0.04025
R34371 VDD.n10509 VDD.n10508 0.04025
R34372 VDD.n10508 VDD.n10507 0.04025
R34373 VDD.n10507 VDD.n8339 0.04025
R34374 VDD.n10503 VDD.n8339 0.04025
R34375 VDD.n10503 VDD.n10502 0.04025
R34376 VDD.n10502 VDD.n10501 0.04025
R34377 VDD.n10501 VDD.n8341 0.04025
R34378 VDD.n10497 VDD.n8341 0.04025
R34379 VDD.n10497 VDD.n10496 0.04025
R34380 VDD.n10496 VDD.n10495 0.04025
R34381 VDD.n10495 VDD.n8343 0.04025
R34382 VDD.n10491 VDD.n8343 0.04025
R34383 VDD.n10491 VDD.n10490 0.04025
R34384 VDD.n10490 VDD.n10489 0.04025
R34385 VDD.n10489 VDD.n8345 0.04025
R34386 VDD.n10485 VDD.n8345 0.04025
R34387 VDD.n10485 VDD.n10484 0.04025
R34388 VDD.n10484 VDD.n10483 0.04025
R34389 VDD.n10483 VDD.n8347 0.04025
R34390 VDD.n10479 VDD.n8347 0.04025
R34391 VDD.n10479 VDD.n10478 0.04025
R34392 VDD.n10478 VDD.n10477 0.04025
R34393 VDD.n10477 VDD.n8349 0.04025
R34394 VDD.n10473 VDD.n8349 0.04025
R34395 VDD.n10473 VDD.n10472 0.04025
R34396 VDD.n10472 VDD.n10471 0.04025
R34397 VDD.n10471 VDD.n8351 0.04025
R34398 VDD.n10467 VDD.n8351 0.04025
R34399 VDD.n10467 VDD.n10466 0.04025
R34400 VDD.n10466 VDD.n10465 0.04025
R34401 VDD.n10465 VDD.n8353 0.04025
R34402 VDD.n10461 VDD.n8353 0.04025
R34403 VDD.n10461 VDD.n10460 0.04025
R34404 VDD.n10460 VDD.n10459 0.04025
R34405 VDD.n10459 VDD.n8355 0.04025
R34406 VDD.n10455 VDD.n8355 0.04025
R34407 VDD.n10455 VDD.n10454 0.04025
R34408 VDD.n10454 VDD.n10453 0.04025
R34409 VDD.n10453 VDD.n8357 0.04025
R34410 VDD.n10449 VDD.n8357 0.04025
R34411 VDD.n10449 VDD.n10448 0.04025
R34412 VDD.n10448 VDD.n10447 0.04025
R34413 VDD.n10447 VDD.n8359 0.04025
R34414 VDD.n10443 VDD.n8359 0.04025
R34415 VDD.n10443 VDD.n10442 0.04025
R34416 VDD.n10442 VDD.n10441 0.04025
R34417 VDD.n10441 VDD.n8361 0.04025
R34418 VDD.n10437 VDD.n8361 0.04025
R34419 VDD.n10437 VDD.n10436 0.04025
R34420 VDD.n10436 VDD.n10435 0.04025
R34421 VDD.n10435 VDD.n8363 0.04025
R34422 VDD.n10431 VDD.n8363 0.04025
R34423 VDD.n10431 VDD.n10430 0.04025
R34424 VDD.n10430 VDD.n10429 0.04025
R34425 VDD.n10429 VDD.n8365 0.04025
R34426 VDD.n10425 VDD.n8365 0.04025
R34427 VDD.n10425 VDD.n10424 0.04025
R34428 VDD.n10424 VDD.n10423 0.04025
R34429 VDD.n10423 VDD.n8367 0.04025
R34430 VDD.n10419 VDD.n8367 0.04025
R34431 VDD.n10419 VDD.n10418 0.04025
R34432 VDD.n10418 VDD.n10417 0.04025
R34433 VDD.n10417 VDD.n8369 0.04025
R34434 VDD.n10413 VDD.n8369 0.04025
R34435 VDD.n10413 VDD.n10412 0.04025
R34436 VDD.n10412 VDD.n10411 0.04025
R34437 VDD.n10411 VDD.n8371 0.04025
R34438 VDD.n10407 VDD.n8371 0.04025
R34439 VDD.n10407 VDD.n10406 0.04025
R34440 VDD.n10406 VDD.n10405 0.04025
R34441 VDD.n10405 VDD.n8373 0.04025
R34442 VDD.n10401 VDD.n8373 0.04025
R34443 VDD.n10401 VDD.n10400 0.04025
R34444 VDD.n10400 VDD.n10399 0.04025
R34445 VDD.n10399 VDD.n8375 0.04025
R34446 VDD.n10395 VDD.n8375 0.04025
R34447 VDD.n10395 VDD.n10394 0.04025
R34448 VDD.n10394 VDD.n10393 0.04025
R34449 VDD.n10393 VDD.n8377 0.04025
R34450 VDD.n10389 VDD.n8377 0.04025
R34451 VDD.n10389 VDD.n10388 0.04025
R34452 VDD.n10388 VDD.n10387 0.04025
R34453 VDD.n10387 VDD.n8379 0.04025
R34454 VDD.n10383 VDD.n8379 0.04025
R34455 VDD.n10383 VDD.n10382 0.04025
R34456 VDD.n10382 VDD.n10381 0.04025
R34457 VDD.n10381 VDD.n8381 0.04025
R34458 VDD.n10377 VDD.n8381 0.04025
R34459 VDD.n10377 VDD.n10376 0.04025
R34460 VDD.n10376 VDD.n10375 0.04025
R34461 VDD.n10375 VDD.n8383 0.04025
R34462 VDD.n10371 VDD.n8383 0.04025
R34463 VDD.n10371 VDD.n10370 0.04025
R34464 VDD.n10370 VDD.n10369 0.04025
R34465 VDD.n10369 VDD.n8385 0.04025
R34466 VDD.n10365 VDD.n8385 0.04025
R34467 VDD.n10365 VDD.n10364 0.04025
R34468 VDD.n10364 VDD.n10363 0.04025
R34469 VDD.n10363 VDD.n8387 0.04025
R34470 VDD.n10359 VDD.n8387 0.04025
R34471 VDD.n10359 VDD.n10358 0.04025
R34472 VDD.n10358 VDD.n10357 0.04025
R34473 VDD.n10357 VDD.n8389 0.04025
R34474 VDD.n10353 VDD.n8389 0.04025
R34475 VDD.n10353 VDD.n10352 0.04025
R34476 VDD.n10352 VDD.n10351 0.04025
R34477 VDD.n10351 VDD.n8391 0.04025
R34478 VDD.n10347 VDD.n8391 0.04025
R34479 VDD.n10347 VDD.n10346 0.04025
R34480 VDD.n10346 VDD.n10345 0.04025
R34481 VDD.n10345 VDD.n8393 0.04025
R34482 VDD.n10341 VDD.n8393 0.04025
R34483 VDD.n10341 VDD.n10340 0.04025
R34484 VDD.n10340 VDD.n10339 0.04025
R34485 VDD.n10339 VDD.n8395 0.04025
R34486 VDD.n10335 VDD.n8395 0.04025
R34487 VDD.n10335 VDD.n10334 0.04025
R34488 VDD.n10334 VDD.n10333 0.04025
R34489 VDD.n10333 VDD.n8397 0.04025
R34490 VDD.n10329 VDD.n8397 0.04025
R34491 VDD.n10329 VDD.n10328 0.04025
R34492 VDD.n10328 VDD.n10327 0.04025
R34493 VDD.n10327 VDD.n8399 0.04025
R34494 VDD.n10323 VDD.n8399 0.04025
R34495 VDD.n10323 VDD.n10322 0.04025
R34496 VDD.n10322 VDD.n10321 0.04025
R34497 VDD.n10321 VDD.n8401 0.04025
R34498 VDD.n10317 VDD.n8401 0.04025
R34499 VDD.n10317 VDD.n10316 0.04025
R34500 VDD.n10316 VDD.n10315 0.04025
R34501 VDD.n10315 VDD.n8403 0.04025
R34502 VDD.n10311 VDD.n8403 0.04025
R34503 VDD.n10311 VDD.n10310 0.04025
R34504 VDD.n10310 VDD.n10309 0.04025
R34505 VDD.n10309 VDD.n8405 0.04025
R34506 VDD.n10305 VDD.n8405 0.04025
R34507 VDD.n10305 VDD.n10304 0.04025
R34508 VDD.n10304 VDD.n10303 0.04025
R34509 VDD.n10303 VDD.n8407 0.04025
R34510 VDD.n10299 VDD.n8407 0.04025
R34511 VDD.n10299 VDD.n10298 0.04025
R34512 VDD.n10298 VDD.n10297 0.04025
R34513 VDD.n10297 VDD.n8409 0.04025
R34514 VDD.n10293 VDD.n8409 0.04025
R34515 VDD.n10293 VDD.n10292 0.04025
R34516 VDD.n10292 VDD.n10291 0.04025
R34517 VDD.n10291 VDD.n8411 0.04025
R34518 VDD.n10287 VDD.n8411 0.04025
R34519 VDD.n10287 VDD.n10286 0.04025
R34520 VDD.n10286 VDD.n10285 0.04025
R34521 VDD.n10285 VDD.n8413 0.04025
R34522 VDD.n10281 VDD.n8413 0.04025
R34523 VDD.n10281 VDD.n10280 0.04025
R34524 VDD.n10280 VDD.n10279 0.04025
R34525 VDD.n10279 VDD.n8415 0.04025
R34526 VDD.n10275 VDD.n8415 0.04025
R34527 VDD.n10275 VDD.n10274 0.04025
R34528 VDD.n10274 VDD.n10273 0.04025
R34529 VDD.n10273 VDD.n8417 0.04025
R34530 VDD.n10269 VDD.n8417 0.04025
R34531 VDD.n10269 VDD.n10268 0.04025
R34532 VDD.n10268 VDD.n10267 0.04025
R34533 VDD.n10267 VDD.n8419 0.04025
R34534 VDD.n10263 VDD.n8419 0.04025
R34535 VDD.n10263 VDD.n10262 0.04025
R34536 VDD.n10262 VDD.n10261 0.04025
R34537 VDD.n10261 VDD.n8421 0.04025
R34538 VDD.n10257 VDD.n8421 0.04025
R34539 VDD.n10257 VDD.n10256 0.04025
R34540 VDD.n10256 VDD.n10255 0.04025
R34541 VDD.n10255 VDD.n8423 0.04025
R34542 VDD.n10251 VDD.n8423 0.04025
R34543 VDD.n10251 VDD.n10250 0.04025
R34544 VDD.n10250 VDD.n10249 0.04025
R34545 VDD.n10249 VDD.n8425 0.04025
R34546 VDD.n10245 VDD.n8425 0.04025
R34547 VDD.n10245 VDD.n10244 0.04025
R34548 VDD.n10244 VDD.n10243 0.04025
R34549 VDD.n10243 VDD.n8427 0.04025
R34550 VDD.n10239 VDD.n8427 0.04025
R34551 VDD.n10239 VDD.n10238 0.04025
R34552 VDD.n10238 VDD.n10237 0.04025
R34553 VDD.n10237 VDD.n8429 0.04025
R34554 VDD.n10233 VDD.n8429 0.04025
R34555 VDD.n10233 VDD.n10232 0.04025
R34556 VDD.n10232 VDD.n10231 0.04025
R34557 VDD.n10231 VDD.n8431 0.04025
R34558 VDD.n10227 VDD.n8431 0.04025
R34559 VDD.n10227 VDD.n10226 0.04025
R34560 VDD.n10226 VDD.n10225 0.04025
R34561 VDD.n10225 VDD.n8433 0.04025
R34562 VDD.n10221 VDD.n8433 0.04025
R34563 VDD.n10221 VDD.n10220 0.04025
R34564 VDD.n10220 VDD.n10219 0.04025
R34565 VDD.n10219 VDD.n8435 0.04025
R34566 VDD.n10215 VDD.n8435 0.04025
R34567 VDD.n10215 VDD.n10214 0.04025
R34568 VDD.n10214 VDD.n10213 0.04025
R34569 VDD.n10213 VDD.n8437 0.04025
R34570 VDD.n10209 VDD.n8437 0.04025
R34571 VDD.n10209 VDD.n10208 0.04025
R34572 VDD.n10208 VDD.n10207 0.04025
R34573 VDD.n10207 VDD.n8439 0.04025
R34574 VDD.n10203 VDD.n8439 0.04025
R34575 VDD.n10203 VDD.n10202 0.04025
R34576 VDD.n10202 VDD.n10201 0.04025
R34577 VDD.n10201 VDD.n8441 0.04025
R34578 VDD.n10197 VDD.n8441 0.04025
R34579 VDD.n10197 VDD.n10196 0.04025
R34580 VDD.n10196 VDD.n10195 0.04025
R34581 VDD.n10195 VDD.n8443 0.04025
R34582 VDD.n10191 VDD.n8443 0.04025
R34583 VDD.n10191 VDD.n10190 0.04025
R34584 VDD.n10190 VDD.n10189 0.04025
R34585 VDD.n10189 VDD.n8445 0.04025
R34586 VDD.n10185 VDD.n8445 0.04025
R34587 VDD.n10185 VDD.n10184 0.04025
R34588 VDD.n10184 VDD.n10183 0.04025
R34589 VDD.n10183 VDD.n8447 0.04025
R34590 VDD.n10179 VDD.n8447 0.04025
R34591 VDD.n10179 VDD.n10178 0.04025
R34592 VDD.n10178 VDD.n10177 0.04025
R34593 VDD.n10177 VDD.n8449 0.04025
R34594 VDD.n10173 VDD.n8449 0.04025
R34595 VDD.n10173 VDD.n10172 0.04025
R34596 VDD.n10172 VDD.n10171 0.04025
R34597 VDD.n10171 VDD.n8451 0.04025
R34598 VDD.n10167 VDD.n8451 0.04025
R34599 VDD.n10167 VDD.n10166 0.04025
R34600 VDD.n10166 VDD.n10165 0.04025
R34601 VDD.n10165 VDD.n8453 0.04025
R34602 VDD.n10161 VDD.n8453 0.04025
R34603 VDD.n10161 VDD.n10160 0.04025
R34604 VDD.n10160 VDD.n10159 0.04025
R34605 VDD.n10159 VDD.n8455 0.04025
R34606 VDD.n10155 VDD.n8455 0.04025
R34607 VDD.n10155 VDD.n10154 0.04025
R34608 VDD.n10154 VDD.n10153 0.04025
R34609 VDD.n10153 VDD.n8457 0.04025
R34610 VDD.n10149 VDD.n8457 0.04025
R34611 VDD.n11137 VDD.n11136 0.04025
R34612 VDD.n11137 VDD.n629 0.04025
R34613 VDD.n11141 VDD.n629 0.04025
R34614 VDD.n11142 VDD.n11141 0.04025
R34615 VDD.n11143 VDD.n11142 0.04025
R34616 VDD.n11143 VDD.n627 0.04025
R34617 VDD.n11147 VDD.n627 0.04025
R34618 VDD.n11148 VDD.n11147 0.04025
R34619 VDD.n11149 VDD.n11148 0.04025
R34620 VDD.n11149 VDD.n625 0.04025
R34621 VDD.n11153 VDD.n625 0.04025
R34622 VDD.n11154 VDD.n11153 0.04025
R34623 VDD.n11155 VDD.n11154 0.04025
R34624 VDD.n11155 VDD.n623 0.04025
R34625 VDD.n11159 VDD.n623 0.04025
R34626 VDD.n11160 VDD.n11159 0.04025
R34627 VDD.n11161 VDD.n11160 0.04025
R34628 VDD.n11161 VDD.n621 0.04025
R34629 VDD.n11165 VDD.n621 0.04025
R34630 VDD.n11166 VDD.n11165 0.04025
R34631 VDD.n11167 VDD.n11166 0.04025
R34632 VDD.n11167 VDD.n619 0.04025
R34633 VDD.n11171 VDD.n619 0.04025
R34634 VDD.n11172 VDD.n11171 0.04025
R34635 VDD.n11173 VDD.n11172 0.04025
R34636 VDD.n11173 VDD.n617 0.04025
R34637 VDD.n11177 VDD.n617 0.04025
R34638 VDD.n11178 VDD.n11177 0.04025
R34639 VDD.n11179 VDD.n11178 0.04025
R34640 VDD.n11179 VDD.n615 0.04025
R34641 VDD.n11183 VDD.n615 0.04025
R34642 VDD.n11184 VDD.n11183 0.04025
R34643 VDD.n11185 VDD.n11184 0.04025
R34644 VDD.n11185 VDD.n613 0.04025
R34645 VDD.n11189 VDD.n613 0.04025
R34646 VDD.n11190 VDD.n11189 0.04025
R34647 VDD.n11191 VDD.n11190 0.04025
R34648 VDD.n11191 VDD.n611 0.04025
R34649 VDD.n11195 VDD.n611 0.04025
R34650 VDD.n11196 VDD.n11195 0.04025
R34651 VDD.n11197 VDD.n11196 0.04025
R34652 VDD.n11197 VDD.n609 0.04025
R34653 VDD.n11201 VDD.n609 0.04025
R34654 VDD.n11202 VDD.n11201 0.04025
R34655 VDD.n11203 VDD.n11202 0.04025
R34656 VDD.n11203 VDD.n607 0.04025
R34657 VDD.n11207 VDD.n607 0.04025
R34658 VDD.n11208 VDD.n11207 0.04025
R34659 VDD.n11209 VDD.n11208 0.04025
R34660 VDD.n11209 VDD.n605 0.04025
R34661 VDD.n11213 VDD.n605 0.04025
R34662 VDD.n11214 VDD.n11213 0.04025
R34663 VDD.n11215 VDD.n11214 0.04025
R34664 VDD.n11215 VDD.n603 0.04025
R34665 VDD.n11219 VDD.n603 0.04025
R34666 VDD.n11220 VDD.n11219 0.04025
R34667 VDD.n11221 VDD.n11220 0.04025
R34668 VDD.n11221 VDD.n601 0.04025
R34669 VDD.n11225 VDD.n601 0.04025
R34670 VDD.n11226 VDD.n11225 0.04025
R34671 VDD.n11227 VDD.n11226 0.04025
R34672 VDD.n11227 VDD.n599 0.04025
R34673 VDD.n11231 VDD.n599 0.04025
R34674 VDD.n11232 VDD.n11231 0.04025
R34675 VDD.n11233 VDD.n11232 0.04025
R34676 VDD.n11233 VDD.n597 0.04025
R34677 VDD.n11237 VDD.n597 0.04025
R34678 VDD.n11238 VDD.n11237 0.04025
R34679 VDD.n11239 VDD.n11238 0.04025
R34680 VDD.n11239 VDD.n595 0.04025
R34681 VDD.n11243 VDD.n595 0.04025
R34682 VDD.n11244 VDD.n11243 0.04025
R34683 VDD.n11245 VDD.n11244 0.04025
R34684 VDD.n11245 VDD.n593 0.04025
R34685 VDD.n11249 VDD.n593 0.04025
R34686 VDD.n11250 VDD.n11249 0.04025
R34687 VDD.n11251 VDD.n11250 0.04025
R34688 VDD.n11251 VDD.n591 0.04025
R34689 VDD.n11255 VDD.n591 0.04025
R34690 VDD.n11256 VDD.n11255 0.04025
R34691 VDD.n11257 VDD.n11256 0.04025
R34692 VDD.n11257 VDD.n589 0.04025
R34693 VDD.n11261 VDD.n589 0.04025
R34694 VDD.n11262 VDD.n11261 0.04025
R34695 VDD.n11263 VDD.n11262 0.04025
R34696 VDD.n11263 VDD.n587 0.04025
R34697 VDD.n11267 VDD.n587 0.04025
R34698 VDD.n11268 VDD.n11267 0.04025
R34699 VDD.n11269 VDD.n11268 0.04025
R34700 VDD.n11269 VDD.n585 0.04025
R34701 VDD.n11273 VDD.n585 0.04025
R34702 VDD.n11274 VDD.n11273 0.04025
R34703 VDD.n11275 VDD.n11274 0.04025
R34704 VDD.n11275 VDD.n583 0.04025
R34705 VDD.n11279 VDD.n583 0.04025
R34706 VDD.n11280 VDD.n11279 0.04025
R34707 VDD.n11281 VDD.n11280 0.04025
R34708 VDD.n11281 VDD.n581 0.04025
R34709 VDD.n11285 VDD.n581 0.04025
R34710 VDD.n11286 VDD.n11285 0.04025
R34711 VDD.n11287 VDD.n11286 0.04025
R34712 VDD.n11287 VDD.n579 0.04025
R34713 VDD.n11291 VDD.n579 0.04025
R34714 VDD.n11292 VDD.n11291 0.04025
R34715 VDD.n11293 VDD.n11292 0.04025
R34716 VDD.n11293 VDD.n577 0.04025
R34717 VDD.n11297 VDD.n577 0.04025
R34718 VDD.n11298 VDD.n11297 0.04025
R34719 VDD.n11299 VDD.n11298 0.04025
R34720 VDD.n11299 VDD.n575 0.04025
R34721 VDD.n11303 VDD.n575 0.04025
R34722 VDD.n11304 VDD.n11303 0.04025
R34723 VDD.n11305 VDD.n11304 0.04025
R34724 VDD.n11305 VDD.n573 0.04025
R34725 VDD.n11309 VDD.n573 0.04025
R34726 VDD.n11310 VDD.n11309 0.04025
R34727 VDD.n11311 VDD.n11310 0.04025
R34728 VDD.n11311 VDD.n571 0.04025
R34729 VDD.n11315 VDD.n571 0.04025
R34730 VDD.n11316 VDD.n11315 0.04025
R34731 VDD.n11317 VDD.n11316 0.04025
R34732 VDD.n11317 VDD.n569 0.04025
R34733 VDD.n11321 VDD.n569 0.04025
R34734 VDD.n11322 VDD.n11321 0.04025
R34735 VDD.n11323 VDD.n11322 0.04025
R34736 VDD.n11323 VDD.n567 0.04025
R34737 VDD.n11327 VDD.n567 0.04025
R34738 VDD.n11328 VDD.n11327 0.04025
R34739 VDD.n11329 VDD.n11328 0.04025
R34740 VDD.n11329 VDD.n565 0.04025
R34741 VDD.n11333 VDD.n565 0.04025
R34742 VDD.n11334 VDD.n11333 0.04025
R34743 VDD.n11335 VDD.n11334 0.04025
R34744 VDD.n11335 VDD.n563 0.04025
R34745 VDD.n11339 VDD.n563 0.04025
R34746 VDD.n11340 VDD.n11339 0.04025
R34747 VDD.n11341 VDD.n11340 0.04025
R34748 VDD.n11341 VDD.n561 0.04025
R34749 VDD.n11345 VDD.n561 0.04025
R34750 VDD.n11346 VDD.n11345 0.04025
R34751 VDD.n11347 VDD.n11346 0.04025
R34752 VDD.n11347 VDD.n559 0.04025
R34753 VDD.n11351 VDD.n559 0.04025
R34754 VDD.n11352 VDD.n11351 0.04025
R34755 VDD.n11353 VDD.n11352 0.04025
R34756 VDD.n11353 VDD.n557 0.04025
R34757 VDD.n11357 VDD.n557 0.04025
R34758 VDD.n11358 VDD.n11357 0.04025
R34759 VDD.n11359 VDD.n11358 0.04025
R34760 VDD.n11359 VDD.n555 0.04025
R34761 VDD.n11363 VDD.n555 0.04025
R34762 VDD.n11364 VDD.n11363 0.04025
R34763 VDD.n11365 VDD.n11364 0.04025
R34764 VDD.n11365 VDD.n553 0.04025
R34765 VDD.n11369 VDD.n553 0.04025
R34766 VDD.n11370 VDD.n11369 0.04025
R34767 VDD.n11371 VDD.n11370 0.04025
R34768 VDD.n11371 VDD.n551 0.04025
R34769 VDD.n11375 VDD.n551 0.04025
R34770 VDD.n11376 VDD.n11375 0.04025
R34771 VDD.n11377 VDD.n11376 0.04025
R34772 VDD.n11377 VDD.n549 0.04025
R34773 VDD.n11381 VDD.n549 0.04025
R34774 VDD.n11382 VDD.n11381 0.04025
R34775 VDD.n11383 VDD.n11382 0.04025
R34776 VDD.n11383 VDD.n547 0.04025
R34777 VDD.n11387 VDD.n547 0.04025
R34778 VDD.n11388 VDD.n11387 0.04025
R34779 VDD.n11389 VDD.n11388 0.04025
R34780 VDD.n11389 VDD.n545 0.04025
R34781 VDD.n11393 VDD.n545 0.04025
R34782 VDD.n11394 VDD.n11393 0.04025
R34783 VDD.n11395 VDD.n11394 0.04025
R34784 VDD.n11395 VDD.n543 0.04025
R34785 VDD.n11399 VDD.n543 0.04025
R34786 VDD.n11400 VDD.n11399 0.04025
R34787 VDD.n11401 VDD.n11400 0.04025
R34788 VDD.n11401 VDD.n541 0.04025
R34789 VDD.n11405 VDD.n541 0.04025
R34790 VDD.n11406 VDD.n11405 0.04025
R34791 VDD.n11407 VDD.n11406 0.04025
R34792 VDD.n11407 VDD.n539 0.04025
R34793 VDD.n11411 VDD.n539 0.04025
R34794 VDD.n11412 VDD.n11411 0.04025
R34795 VDD.n11413 VDD.n11412 0.04025
R34796 VDD.n11413 VDD.n537 0.04025
R34797 VDD.n11417 VDD.n537 0.04025
R34798 VDD.n11418 VDD.n11417 0.04025
R34799 VDD.n11419 VDD.n11418 0.04025
R34800 VDD.n11419 VDD.n535 0.04025
R34801 VDD.n11423 VDD.n535 0.04025
R34802 VDD.n11424 VDD.n11423 0.04025
R34803 VDD.n11425 VDD.n11424 0.04025
R34804 VDD.n11425 VDD.n533 0.04025
R34805 VDD.n11429 VDD.n533 0.04025
R34806 VDD.n11430 VDD.n11429 0.04025
R34807 VDD.n11431 VDD.n11430 0.04025
R34808 VDD.n11431 VDD.n531 0.04025
R34809 VDD.n11435 VDD.n531 0.04025
R34810 VDD.n11436 VDD.n11435 0.04025
R34811 VDD.n11437 VDD.n11436 0.04025
R34812 VDD.n11437 VDD.n529 0.04025
R34813 VDD.n11441 VDD.n529 0.04025
R34814 VDD.n11442 VDD.n11441 0.04025
R34815 VDD.n11443 VDD.n11442 0.04025
R34816 VDD.n11443 VDD.n527 0.04025
R34817 VDD.n11447 VDD.n527 0.04025
R34818 VDD.n11448 VDD.n11447 0.04025
R34819 VDD.n11449 VDD.n11448 0.04025
R34820 VDD.n11449 VDD.n525 0.04025
R34821 VDD.n11453 VDD.n525 0.04025
R34822 VDD.n11454 VDD.n11453 0.04025
R34823 VDD.n11455 VDD.n11454 0.04025
R34824 VDD.n11455 VDD.n523 0.04025
R34825 VDD.n11459 VDD.n523 0.04025
R34826 VDD.n11460 VDD.n11459 0.04025
R34827 VDD.n11461 VDD.n11460 0.04025
R34828 VDD.n11461 VDD.n521 0.04025
R34829 VDD.n11465 VDD.n521 0.04025
R34830 VDD.n11466 VDD.n11465 0.04025
R34831 VDD.n11467 VDD.n11466 0.04025
R34832 VDD.n11467 VDD.n519 0.04025
R34833 VDD.n11471 VDD.n519 0.04025
R34834 VDD.n11472 VDD.n11471 0.04025
R34835 VDD.n11473 VDD.n11472 0.04025
R34836 VDD.n11473 VDD.n517 0.04025
R34837 VDD.n11477 VDD.n517 0.04025
R34838 VDD.n11478 VDD.n11477 0.04025
R34839 VDD.n11479 VDD.n11478 0.04025
R34840 VDD.n11479 VDD.n515 0.04025
R34841 VDD.n11483 VDD.n515 0.04025
R34842 VDD.n11484 VDD.n11483 0.04025
R34843 VDD.n11485 VDD.n11484 0.04025
R34844 VDD.n11485 VDD.n513 0.04025
R34845 VDD.n11489 VDD.n513 0.04025
R34846 VDD.n11490 VDD.n11489 0.04025
R34847 VDD.n11491 VDD.n11490 0.04025
R34848 VDD.n11491 VDD.n511 0.04025
R34849 VDD.n11495 VDD.n511 0.04025
R34850 VDD.n11496 VDD.n11495 0.04025
R34851 VDD.n11497 VDD.n11496 0.04025
R34852 VDD.n11497 VDD.n509 0.04025
R34853 VDD.n11501 VDD.n509 0.04025
R34854 VDD.n11502 VDD.n11501 0.04025
R34855 VDD.n11503 VDD.n11502 0.04025
R34856 VDD.n11503 VDD.n507 0.04025
R34857 VDD.n11507 VDD.n507 0.04025
R34858 VDD.n11508 VDD.n11507 0.04025
R34859 VDD.n11509 VDD.n11508 0.04025
R34860 VDD.n11509 VDD.n505 0.04025
R34861 VDD.n11513 VDD.n505 0.04025
R34862 VDD.n11514 VDD.n11513 0.04025
R34863 VDD.n11515 VDD.n11514 0.04025
R34864 VDD.n11515 VDD.n503 0.04025
R34865 VDD.n11519 VDD.n503 0.04025
R34866 VDD.n11520 VDD.n11519 0.04025
R34867 VDD.n11521 VDD.n11520 0.04025
R34868 VDD.n11521 VDD.n501 0.04025
R34869 VDD.n11525 VDD.n501 0.04025
R34870 VDD.n11526 VDD.n11525 0.04025
R34871 VDD.n11527 VDD.n11526 0.04025
R34872 VDD.n11527 VDD.n499 0.04025
R34873 VDD.n11531 VDD.n499 0.04025
R34874 VDD.n11532 VDD.n11531 0.04025
R34875 VDD.n11533 VDD.n11532 0.04025
R34876 VDD.n11533 VDD.n497 0.04025
R34877 VDD.n11537 VDD.n497 0.04025
R34878 VDD.n11538 VDD.n11537 0.04025
R34879 VDD.n11539 VDD.n11538 0.04025
R34880 VDD.n11539 VDD.n495 0.04025
R34881 VDD.n11543 VDD.n495 0.04025
R34882 VDD.n11544 VDD.n11543 0.04025
R34883 VDD.n11545 VDD.n11544 0.04025
R34884 VDD.n11545 VDD.n493 0.04025
R34885 VDD.n11549 VDD.n493 0.04025
R34886 VDD.n11550 VDD.n11549 0.04025
R34887 VDD.n11551 VDD.n11550 0.04025
R34888 VDD.n11551 VDD.n491 0.04025
R34889 VDD.n11555 VDD.n491 0.04025
R34890 VDD.n11556 VDD.n11555 0.04025
R34891 VDD.n11557 VDD.n11556 0.04025
R34892 VDD.n11557 VDD.n489 0.04025
R34893 VDD.n11561 VDD.n489 0.04025
R34894 VDD.n11562 VDD.n11561 0.04025
R34895 VDD.n11563 VDD.n11562 0.04025
R34896 VDD.n11563 VDD.n487 0.04025
R34897 VDD.n11567 VDD.n487 0.04025
R34898 VDD.n11568 VDD.n11567 0.04025
R34899 VDD.n11569 VDD.n11568 0.04025
R34900 VDD.n11569 VDD.n485 0.04025
R34901 VDD.n11573 VDD.n485 0.04025
R34902 VDD.n11574 VDD.n11573 0.04025
R34903 VDD.n11575 VDD.n11574 0.04025
R34904 VDD.n11575 VDD.n483 0.04025
R34905 VDD.n11579 VDD.n483 0.04025
R34906 VDD.n11580 VDD.n11579 0.04025
R34907 VDD.n11581 VDD.n11580 0.04025
R34908 VDD.n11581 VDD.n481 0.04025
R34909 VDD.n11585 VDD.n481 0.04025
R34910 VDD.n11586 VDD.n11585 0.04025
R34911 VDD.n11587 VDD.n11586 0.04025
R34912 VDD.n11587 VDD.n479 0.04025
R34913 VDD.n11591 VDD.n479 0.04025
R34914 VDD.n11592 VDD.n11591 0.04025
R34915 VDD.n11593 VDD.n11592 0.04025
R34916 VDD.n11593 VDD.n477 0.04025
R34917 VDD.n11597 VDD.n477 0.04025
R34918 VDD.n11598 VDD.n11597 0.04025
R34919 VDD.n11599 VDD.n11598 0.04025
R34920 VDD.n11599 VDD.n475 0.04025
R34921 VDD.n11603 VDD.n475 0.04025
R34922 VDD.n11604 VDD.n11603 0.04025
R34923 VDD.n11605 VDD.n11604 0.04025
R34924 VDD.n11605 VDD.n473 0.04025
R34925 VDD.n11609 VDD.n473 0.04025
R34926 VDD.n11610 VDD.n11609 0.04025
R34927 VDD.n11611 VDD.n11610 0.04025
R34928 VDD.n11611 VDD.n471 0.04025
R34929 VDD.n11615 VDD.n471 0.04025
R34930 VDD.n11616 VDD.n11615 0.04025
R34931 VDD.n11617 VDD.n11616 0.04025
R34932 VDD.n11617 VDD.n469 0.04025
R34933 VDD.n11621 VDD.n469 0.04025
R34934 VDD.n11622 VDD.n11621 0.04025
R34935 VDD.n11623 VDD.n11622 0.04025
R34936 VDD.n11623 VDD.n467 0.04025
R34937 VDD.n11627 VDD.n467 0.04025
R34938 VDD.n11628 VDD.n11627 0.04025
R34939 VDD.n11629 VDD.n11628 0.04025
R34940 VDD.n11629 VDD.n465 0.04025
R34941 VDD.n11633 VDD.n465 0.04025
R34942 VDD.n11634 VDD.n11633 0.04025
R34943 VDD.n11635 VDD.n11634 0.04025
R34944 VDD.n11635 VDD.n463 0.04025
R34945 VDD.n11639 VDD.n463 0.04025
R34946 VDD.n11640 VDD.n11639 0.04025
R34947 VDD.n11641 VDD.n11640 0.04025
R34948 VDD.n11641 VDD.n461 0.04025
R34949 VDD.n11645 VDD.n461 0.04025
R34950 VDD.n11646 VDD.n11645 0.04025
R34951 VDD.n11647 VDD.n11646 0.04025
R34952 VDD.n11647 VDD.n459 0.04025
R34953 VDD.n11651 VDD.n459 0.04025
R34954 VDD.n11652 VDD.n11651 0.04025
R34955 VDD.n11653 VDD.n11652 0.04025
R34956 VDD.n11653 VDD.n457 0.04025
R34957 VDD.n11657 VDD.n457 0.04025
R34958 VDD.n11658 VDD.n11657 0.04025
R34959 VDD.n11659 VDD.n11658 0.04025
R34960 VDD.n11659 VDD.n455 0.04025
R34961 VDD.n11663 VDD.n455 0.04025
R34962 VDD.n11664 VDD.n11663 0.04025
R34963 VDD.n11665 VDD.n11664 0.04025
R34964 VDD.n11665 VDD.n453 0.04025
R34965 VDD.n11669 VDD.n453 0.04025
R34966 VDD.n11670 VDD.n11669 0.04025
R34967 VDD.n11671 VDD.n11670 0.04025
R34968 VDD.n11671 VDD.n451 0.04025
R34969 VDD.n11675 VDD.n451 0.04025
R34970 VDD.n11676 VDD.n11675 0.04025
R34971 VDD.n11677 VDD.n11676 0.04025
R34972 VDD.n11677 VDD.n449 0.04025
R34973 VDD.n11681 VDD.n449 0.04025
R34974 VDD.n11682 VDD.n11681 0.04025
R34975 VDD.n11683 VDD.n11682 0.04025
R34976 VDD.n11683 VDD.n447 0.04025
R34977 VDD.n11687 VDD.n447 0.04025
R34978 VDD.n11688 VDD.n11687 0.04025
R34979 VDD.n11689 VDD.n11688 0.04025
R34980 VDD.n11689 VDD.n445 0.04025
R34981 VDD.n11693 VDD.n445 0.04025
R34982 VDD.n11694 VDD.n11693 0.04025
R34983 VDD.n11695 VDD.n11694 0.04025
R34984 VDD.n11695 VDD.n443 0.04025
R34985 VDD.n11699 VDD.n443 0.04025
R34986 VDD.n11700 VDD.n11699 0.04025
R34987 VDD.n11701 VDD.n11700 0.04025
R34988 VDD.n11701 VDD.n441 0.04025
R34989 VDD.n11705 VDD.n441 0.04025
R34990 VDD.n11706 VDD.n11705 0.04025
R34991 VDD.n11707 VDD.n11706 0.04025
R34992 VDD.n11707 VDD.n439 0.04025
R34993 VDD.n11711 VDD.n439 0.04025
R34994 VDD.n11712 VDD.n11711 0.04025
R34995 VDD.n11713 VDD.n11712 0.04025
R34996 VDD.n11713 VDD.n437 0.04025
R34997 VDD.n11717 VDD.n437 0.04025
R34998 VDD.n11718 VDD.n11717 0.04025
R34999 VDD.n11719 VDD.n11718 0.04025
R35000 VDD.n11719 VDD.n435 0.04025
R35001 VDD.n11723 VDD.n435 0.04025
R35002 VDD.n11724 VDD.n11723 0.04025
R35003 VDD.n11725 VDD.n11724 0.04025
R35004 VDD.n11725 VDD.n433 0.04025
R35005 VDD.n11729 VDD.n433 0.04025
R35006 VDD.n11730 VDD.n11729 0.04025
R35007 VDD.n11731 VDD.n11730 0.04025
R35008 VDD.n11731 VDD.n431 0.04025
R35009 VDD.n11735 VDD.n431 0.04025
R35010 VDD.n11736 VDD.n11735 0.04025
R35011 VDD.n11737 VDD.n11736 0.04025
R35012 VDD.n11737 VDD.n429 0.04025
R35013 VDD.n11741 VDD.n429 0.04025
R35014 VDD.n11742 VDD.n11741 0.04025
R35015 VDD.n11743 VDD.n11742 0.04025
R35016 VDD.n11743 VDD.n427 0.04025
R35017 VDD.n11747 VDD.n427 0.04025
R35018 VDD.n11748 VDD.n11747 0.04025
R35019 VDD.n11749 VDD.n11748 0.04025
R35020 VDD.n11749 VDD.n425 0.04025
R35021 VDD.n11753 VDD.n425 0.04025
R35022 VDD.n11754 VDD.n11753 0.04025
R35023 VDD.n11755 VDD.n11754 0.04025
R35024 VDD.n11755 VDD.n423 0.04025
R35025 VDD.n11759 VDD.n423 0.04025
R35026 VDD.n11760 VDD.n11759 0.04025
R35027 VDD.n11761 VDD.n11760 0.04025
R35028 VDD.n11761 VDD.n421 0.04025
R35029 VDD.n11765 VDD.n421 0.04025
R35030 VDD.n11766 VDD.n11765 0.04025
R35031 VDD.n11767 VDD.n11766 0.04025
R35032 VDD.n11767 VDD.n419 0.04025
R35033 VDD.n11771 VDD.n419 0.04025
R35034 VDD.n11772 VDD.n11771 0.04025
R35035 VDD.n11773 VDD.n11772 0.04025
R35036 VDD.n11773 VDD.n417 0.04025
R35037 VDD.n11777 VDD.n417 0.04025
R35038 VDD.n11778 VDD.n11777 0.04025
R35039 VDD.n11779 VDD.n11778 0.04025
R35040 VDD.n11779 VDD.n415 0.04025
R35041 VDD.n11783 VDD.n415 0.04025
R35042 VDD.n11784 VDD.n11783 0.04025
R35043 VDD.n11785 VDD.n11784 0.04025
R35044 VDD.n11785 VDD.n413 0.04025
R35045 VDD.n11789 VDD.n413 0.04025
R35046 VDD.n11790 VDD.n11789 0.04025
R35047 VDD.n11791 VDD.n11790 0.04025
R35048 VDD.n11791 VDD.n411 0.04025
R35049 VDD.n11795 VDD.n411 0.04025
R35050 VDD.n11796 VDD.n11795 0.04025
R35051 VDD.n11797 VDD.n11796 0.04025
R35052 VDD.n11797 VDD.n409 0.04025
R35053 VDD.n11801 VDD.n409 0.04025
R35054 VDD.n11802 VDD.n11801 0.04025
R35055 VDD.n11803 VDD.n11802 0.04025
R35056 VDD.n11803 VDD.n407 0.04025
R35057 VDD.n11807 VDD.n407 0.04025
R35058 VDD.n11808 VDD.n11807 0.04025
R35059 VDD.n11809 VDD.n11808 0.04025
R35060 VDD.n11809 VDD.n405 0.04025
R35061 VDD.n3629 VDD.n2746 0.04025
R35062 VDD.n3625 VDD.n2746 0.04025
R35063 VDD.n3625 VDD.n3624 0.04025
R35064 VDD.n3624 VDD.n3623 0.04025
R35065 VDD.n3623 VDD.n2748 0.04025
R35066 VDD.n3619 VDD.n2748 0.04025
R35067 VDD.n3619 VDD.n3618 0.04025
R35068 VDD.n3618 VDD.n3617 0.04025
R35069 VDD.n3617 VDD.n2750 0.04025
R35070 VDD.n3613 VDD.n2750 0.04025
R35071 VDD.n3613 VDD.n3612 0.04025
R35072 VDD.n3612 VDD.n3611 0.04025
R35073 VDD.n3611 VDD.n2752 0.04025
R35074 VDD.n3607 VDD.n2752 0.04025
R35075 VDD.n3607 VDD.n3606 0.04025
R35076 VDD.n3606 VDD.n3605 0.04025
R35077 VDD.n3605 VDD.n2754 0.04025
R35078 VDD.n3601 VDD.n2754 0.04025
R35079 VDD.n3601 VDD.n3600 0.04025
R35080 VDD.n3600 VDD.n3599 0.04025
R35081 VDD.n3599 VDD.n2756 0.04025
R35082 VDD.n3595 VDD.n2756 0.04025
R35083 VDD.n3595 VDD.n3594 0.04025
R35084 VDD.n3594 VDD.n3593 0.04025
R35085 VDD.n3593 VDD.n2758 0.04025
R35086 VDD.n3589 VDD.n2758 0.04025
R35087 VDD.n3589 VDD.n3588 0.04025
R35088 VDD.n3588 VDD.n3587 0.04025
R35089 VDD.n3587 VDD.n2760 0.04025
R35090 VDD.n3583 VDD.n2760 0.04025
R35091 VDD.n3583 VDD.n3582 0.04025
R35092 VDD.n3582 VDD.n3581 0.04025
R35093 VDD.n3581 VDD.n2762 0.04025
R35094 VDD.n3577 VDD.n2762 0.04025
R35095 VDD.n3577 VDD.n3576 0.04025
R35096 VDD.n3576 VDD.n3575 0.04025
R35097 VDD.n3575 VDD.n2764 0.04025
R35098 VDD.n3571 VDD.n2764 0.04025
R35099 VDD.n3571 VDD.n3570 0.04025
R35100 VDD.n3570 VDD.n3569 0.04025
R35101 VDD.n3569 VDD.n2766 0.04025
R35102 VDD.n3565 VDD.n2766 0.04025
R35103 VDD.n3565 VDD.n3564 0.04025
R35104 VDD.n3564 VDD.n3563 0.04025
R35105 VDD.n3563 VDD.n2768 0.04025
R35106 VDD.n3559 VDD.n2768 0.04025
R35107 VDD.n3559 VDD.n3558 0.04025
R35108 VDD.n3558 VDD.n3557 0.04025
R35109 VDD.n3557 VDD.n2770 0.04025
R35110 VDD.n3553 VDD.n2770 0.04025
R35111 VDD.n3553 VDD.n3552 0.04025
R35112 VDD.n3552 VDD.n3551 0.04025
R35113 VDD.n3551 VDD.n2772 0.04025
R35114 VDD.n3547 VDD.n2772 0.04025
R35115 VDD.n3547 VDD.n3546 0.04025
R35116 VDD.n3546 VDD.n3545 0.04025
R35117 VDD.n3545 VDD.n2774 0.04025
R35118 VDD.n3541 VDD.n2774 0.04025
R35119 VDD.n3541 VDD.n3540 0.04025
R35120 VDD.n3540 VDD.n3539 0.04025
R35121 VDD.n3539 VDD.n2776 0.04025
R35122 VDD.n3535 VDD.n2776 0.04025
R35123 VDD.n3535 VDD.n3534 0.04025
R35124 VDD.n3534 VDD.n3533 0.04025
R35125 VDD.n3533 VDD.n2778 0.04025
R35126 VDD.n3529 VDD.n2778 0.04025
R35127 VDD.n3529 VDD.n3528 0.04025
R35128 VDD.n3528 VDD.n3527 0.04025
R35129 VDD.n3527 VDD.n2780 0.04025
R35130 VDD.n3523 VDD.n2780 0.04025
R35131 VDD.n3523 VDD.n3522 0.04025
R35132 VDD.n3522 VDD.n3521 0.04025
R35133 VDD.n3521 VDD.n2782 0.04025
R35134 VDD.n3517 VDD.n2782 0.04025
R35135 VDD.n3517 VDD.n3516 0.04025
R35136 VDD.n3516 VDD.n3515 0.04025
R35137 VDD.n3515 VDD.n2784 0.04025
R35138 VDD.n3511 VDD.n2784 0.04025
R35139 VDD.n3511 VDD.n3510 0.04025
R35140 VDD.n3510 VDD.n3509 0.04025
R35141 VDD.n3509 VDD.n2786 0.04025
R35142 VDD.n3505 VDD.n2786 0.04025
R35143 VDD.n3505 VDD.n3504 0.04025
R35144 VDD.n3504 VDD.n3503 0.04025
R35145 VDD.n3503 VDD.n2788 0.04025
R35146 VDD.n3499 VDD.n2788 0.04025
R35147 VDD.n3499 VDD.n3498 0.04025
R35148 VDD.n3498 VDD.n3497 0.04025
R35149 VDD.n3497 VDD.n2790 0.04025
R35150 VDD.n3493 VDD.n2790 0.04025
R35151 VDD.n3493 VDD.n3492 0.04025
R35152 VDD.n3492 VDD.n3491 0.04025
R35153 VDD.n3491 VDD.n2792 0.04025
R35154 VDD.n3487 VDD.n2792 0.04025
R35155 VDD.n3487 VDD.n3486 0.04025
R35156 VDD.n3486 VDD.n3485 0.04025
R35157 VDD.n3485 VDD.n2794 0.04025
R35158 VDD.n3481 VDD.n2794 0.04025
R35159 VDD.n3481 VDD.n3480 0.04025
R35160 VDD.n3480 VDD.n3479 0.04025
R35161 VDD.n3479 VDD.n2796 0.04025
R35162 VDD.n3475 VDD.n2796 0.04025
R35163 VDD.n3475 VDD.n3474 0.04025
R35164 VDD.n3474 VDD.n3473 0.04025
R35165 VDD.n3473 VDD.n2798 0.04025
R35166 VDD.n3469 VDD.n2798 0.04025
R35167 VDD.n3469 VDD.n3468 0.04025
R35168 VDD.n3468 VDD.n3467 0.04025
R35169 VDD.n3467 VDD.n2800 0.04025
R35170 VDD.n3463 VDD.n2800 0.04025
R35171 VDD.n3463 VDD.n3462 0.04025
R35172 VDD.n3462 VDD.n3461 0.04025
R35173 VDD.n3461 VDD.n2802 0.04025
R35174 VDD.n3457 VDD.n2802 0.04025
R35175 VDD.n3457 VDD.n3456 0.04025
R35176 VDD.n3456 VDD.n3455 0.04025
R35177 VDD.n3455 VDD.n2804 0.04025
R35178 VDD.n3451 VDD.n2804 0.04025
R35179 VDD.n3451 VDD.n3450 0.04025
R35180 VDD.n3450 VDD.n3449 0.04025
R35181 VDD.n3449 VDD.n2806 0.04025
R35182 VDD.n3445 VDD.n2806 0.04025
R35183 VDD.n3445 VDD.n3444 0.04025
R35184 VDD.n3444 VDD.n3443 0.04025
R35185 VDD.n3443 VDD.n2808 0.04025
R35186 VDD.n3439 VDD.n2808 0.04025
R35187 VDD.n3439 VDD.n3438 0.04025
R35188 VDD.n3438 VDD.n3437 0.04025
R35189 VDD.n3437 VDD.n2810 0.04025
R35190 VDD.n3433 VDD.n2810 0.04025
R35191 VDD.n3433 VDD.n3432 0.04025
R35192 VDD.n3432 VDD.n3431 0.04025
R35193 VDD.n3431 VDD.n2812 0.04025
R35194 VDD.n3427 VDD.n2812 0.04025
R35195 VDD.n3427 VDD.n3426 0.04025
R35196 VDD.n3426 VDD.n3425 0.04025
R35197 VDD.n3425 VDD.n2814 0.04025
R35198 VDD.n3421 VDD.n2814 0.04025
R35199 VDD.n3421 VDD.n3420 0.04025
R35200 VDD.n3420 VDD.n3419 0.04025
R35201 VDD.n3419 VDD.n2816 0.04025
R35202 VDD.n3415 VDD.n2816 0.04025
R35203 VDD.n3415 VDD.n3414 0.04025
R35204 VDD.n3414 VDD.n3413 0.04025
R35205 VDD.n3413 VDD.n2818 0.04025
R35206 VDD.n3409 VDD.n2818 0.04025
R35207 VDD.n3409 VDD.n3408 0.04025
R35208 VDD.n3408 VDD.n3407 0.04025
R35209 VDD.n3407 VDD.n2820 0.04025
R35210 VDD.n3403 VDD.n2820 0.04025
R35211 VDD.n3403 VDD.n3402 0.04025
R35212 VDD.n3402 VDD.n3401 0.04025
R35213 VDD.n3401 VDD.n2822 0.04025
R35214 VDD.n3397 VDD.n2822 0.04025
R35215 VDD.n3397 VDD.n3396 0.04025
R35216 VDD.n3396 VDD.n3395 0.04025
R35217 VDD.n3395 VDD.n2824 0.04025
R35218 VDD.n3391 VDD.n2824 0.04025
R35219 VDD.n3391 VDD.n3390 0.04025
R35220 VDD.n3390 VDD.n3389 0.04025
R35221 VDD.n3389 VDD.n2826 0.04025
R35222 VDD.n3385 VDD.n2826 0.04025
R35223 VDD.n3385 VDD.n3384 0.04025
R35224 VDD.n3384 VDD.n3383 0.04025
R35225 VDD.n3383 VDD.n2828 0.04025
R35226 VDD.n3379 VDD.n2828 0.04025
R35227 VDD.n3379 VDD.n3378 0.04025
R35228 VDD.n3378 VDD.n3377 0.04025
R35229 VDD.n3377 VDD.n2830 0.04025
R35230 VDD.n3373 VDD.n2830 0.04025
R35231 VDD.n3373 VDD.n3372 0.04025
R35232 VDD.n3372 VDD.n3371 0.04025
R35233 VDD.n3371 VDD.n2832 0.04025
R35234 VDD.n3367 VDD.n2832 0.04025
R35235 VDD.n3367 VDD.n3366 0.04025
R35236 VDD.n3366 VDD.n3365 0.04025
R35237 VDD.n3365 VDD.n2834 0.04025
R35238 VDD.n3361 VDD.n2834 0.04025
R35239 VDD.n3361 VDD.n3360 0.04025
R35240 VDD.n3360 VDD.n3359 0.04025
R35241 VDD.n3359 VDD.n2836 0.04025
R35242 VDD.n3355 VDD.n2836 0.04025
R35243 VDD.n3355 VDD.n3354 0.04025
R35244 VDD.n3354 VDD.n3353 0.04025
R35245 VDD.n3353 VDD.n2838 0.04025
R35246 VDD.n3349 VDD.n2838 0.04025
R35247 VDD.n3349 VDD.n3348 0.04025
R35248 VDD.n3348 VDD.n3347 0.04025
R35249 VDD.n3347 VDD.n2840 0.04025
R35250 VDD.n3343 VDD.n2840 0.04025
R35251 VDD.n3343 VDD.n3342 0.04025
R35252 VDD.n3342 VDD.n3341 0.04025
R35253 VDD.n3341 VDD.n2842 0.04025
R35254 VDD.n3337 VDD.n2842 0.04025
R35255 VDD.n3337 VDD.n3336 0.04025
R35256 VDD.n3336 VDD.n3335 0.04025
R35257 VDD.n3335 VDD.n2844 0.04025
R35258 VDD.n3331 VDD.n2844 0.04025
R35259 VDD.n3331 VDD.n3330 0.04025
R35260 VDD.n3330 VDD.n3329 0.04025
R35261 VDD.n3329 VDD.n2846 0.04025
R35262 VDD.n3325 VDD.n2846 0.04025
R35263 VDD.n3325 VDD.n3324 0.04025
R35264 VDD.n3324 VDD.n3323 0.04025
R35265 VDD.n3323 VDD.n2848 0.04025
R35266 VDD.n3319 VDD.n2848 0.04025
R35267 VDD.n3319 VDD.n3318 0.04025
R35268 VDD.n3318 VDD.n3317 0.04025
R35269 VDD.n3317 VDD.n2850 0.04025
R35270 VDD.n3313 VDD.n2850 0.04025
R35271 VDD.n3313 VDD.n3312 0.04025
R35272 VDD.n3312 VDD.n3311 0.04025
R35273 VDD.n3311 VDD.n2852 0.04025
R35274 VDD.n3307 VDD.n2852 0.04025
R35275 VDD.n3307 VDD.n3306 0.04025
R35276 VDD.n3306 VDD.n3305 0.04025
R35277 VDD.n3305 VDD.n2854 0.04025
R35278 VDD.n3301 VDD.n2854 0.04025
R35279 VDD.n3301 VDD.n3300 0.04025
R35280 VDD.n3300 VDD.n3299 0.04025
R35281 VDD.n3299 VDD.n2856 0.04025
R35282 VDD.n3295 VDD.n2856 0.04025
R35283 VDD.n3295 VDD.n3294 0.04025
R35284 VDD.n3294 VDD.n3293 0.04025
R35285 VDD.n3293 VDD.n2858 0.04025
R35286 VDD.n3289 VDD.n2858 0.04025
R35287 VDD.n3289 VDD.n3288 0.04025
R35288 VDD.n3288 VDD.n3287 0.04025
R35289 VDD.n3287 VDD.n2860 0.04025
R35290 VDD.n3283 VDD.n2860 0.04025
R35291 VDD.n3283 VDD.n3282 0.04025
R35292 VDD.n3282 VDD.n3281 0.04025
R35293 VDD.n3281 VDD.n2862 0.04025
R35294 VDD.n3277 VDD.n2862 0.04025
R35295 VDD.n3277 VDD.n3276 0.04025
R35296 VDD.n3276 VDD.n3275 0.04025
R35297 VDD.n3275 VDD.n2864 0.04025
R35298 VDD.n3271 VDD.n2864 0.04025
R35299 VDD.n3271 VDD.n3270 0.04025
R35300 VDD.n3270 VDD.n3269 0.04025
R35301 VDD.n3269 VDD.n2866 0.04025
R35302 VDD.n3265 VDD.n2866 0.04025
R35303 VDD.n3265 VDD.n3264 0.04025
R35304 VDD.n3264 VDD.n3263 0.04025
R35305 VDD.n3263 VDD.n2868 0.04025
R35306 VDD.n3259 VDD.n2868 0.04025
R35307 VDD.n3259 VDD.n3258 0.04025
R35308 VDD.n3258 VDD.n3257 0.04025
R35309 VDD.n3257 VDD.n2870 0.04025
R35310 VDD.n3253 VDD.n2870 0.04025
R35311 VDD.n3253 VDD.n3252 0.04025
R35312 VDD.n3252 VDD.n3251 0.04025
R35313 VDD.n3251 VDD.n2872 0.04025
R35314 VDD.n3247 VDD.n2872 0.04025
R35315 VDD.n3247 VDD.n3246 0.04025
R35316 VDD.n3246 VDD.n3245 0.04025
R35317 VDD.n3245 VDD.n2874 0.04025
R35318 VDD.n3241 VDD.n2874 0.04025
R35319 VDD.n3241 VDD.n3240 0.04025
R35320 VDD.n3240 VDD.n3239 0.04025
R35321 VDD.n3239 VDD.n2876 0.04025
R35322 VDD.n3235 VDD.n2876 0.04025
R35323 VDD.n3235 VDD.n3234 0.04025
R35324 VDD.n3234 VDD.n3233 0.04025
R35325 VDD.n3233 VDD.n2878 0.04025
R35326 VDD.n3229 VDD.n2878 0.04025
R35327 VDD.n3229 VDD.n3228 0.04025
R35328 VDD.n3228 VDD.n3227 0.04025
R35329 VDD.n3227 VDD.n2880 0.04025
R35330 VDD.n3223 VDD.n2880 0.04025
R35331 VDD.n3223 VDD.n3222 0.04025
R35332 VDD.n3222 VDD.n3221 0.04025
R35333 VDD.n3221 VDD.n2882 0.04025
R35334 VDD.n3217 VDD.n2882 0.04025
R35335 VDD.n3217 VDD.n3216 0.04025
R35336 VDD.n3216 VDD.n3215 0.04025
R35337 VDD.n3215 VDD.n2884 0.04025
R35338 VDD.n3211 VDD.n2884 0.04025
R35339 VDD.n3211 VDD.n3210 0.04025
R35340 VDD.n3210 VDD.n3209 0.04025
R35341 VDD.n3209 VDD.n2886 0.04025
R35342 VDD.n3205 VDD.n2886 0.04025
R35343 VDD.n3205 VDD.n3204 0.04025
R35344 VDD.n3204 VDD.n3203 0.04025
R35345 VDD.n3203 VDD.n2888 0.04025
R35346 VDD.n3199 VDD.n2888 0.04025
R35347 VDD.n3199 VDD.n3198 0.04025
R35348 VDD.n3198 VDD.n3197 0.04025
R35349 VDD.n3197 VDD.n2890 0.04025
R35350 VDD.n3193 VDD.n2890 0.04025
R35351 VDD.n3193 VDD.n3192 0.04025
R35352 VDD.n3192 VDD.n3191 0.04025
R35353 VDD.n3191 VDD.n2892 0.04025
R35354 VDD.n3187 VDD.n2892 0.04025
R35355 VDD.n3187 VDD.n3186 0.04025
R35356 VDD.n3186 VDD.n3185 0.04025
R35357 VDD.n3185 VDD.n2894 0.04025
R35358 VDD.n3181 VDD.n2894 0.04025
R35359 VDD.n3181 VDD.n3180 0.04025
R35360 VDD.n3180 VDD.n3179 0.04025
R35361 VDD.n3179 VDD.n2896 0.04025
R35362 VDD.n3175 VDD.n2896 0.04025
R35363 VDD.n3175 VDD.n3174 0.04025
R35364 VDD.n3174 VDD.n3173 0.04025
R35365 VDD.n3173 VDD.n2898 0.04025
R35366 VDD.n3169 VDD.n2898 0.04025
R35367 VDD.n3169 VDD.n3168 0.04025
R35368 VDD.n3168 VDD.n3167 0.04025
R35369 VDD.n3167 VDD.n2900 0.04025
R35370 VDD.n3163 VDD.n2900 0.04025
R35371 VDD.n3163 VDD.n3162 0.04025
R35372 VDD.n3162 VDD.n3161 0.04025
R35373 VDD.n3161 VDD.n2902 0.04025
R35374 VDD.n3157 VDD.n2902 0.04025
R35375 VDD.n3157 VDD.n3156 0.04025
R35376 VDD.n3156 VDD.n3155 0.04025
R35377 VDD.n3155 VDD.n2904 0.04025
R35378 VDD.n3151 VDD.n2904 0.04025
R35379 VDD.n3151 VDD.n3150 0.04025
R35380 VDD.n3150 VDD.n3149 0.04025
R35381 VDD.n3149 VDD.n2906 0.04025
R35382 VDD.n3145 VDD.n2906 0.04025
R35383 VDD.n3145 VDD.n3144 0.04025
R35384 VDD.n3144 VDD.n3143 0.04025
R35385 VDD.n3143 VDD.n2908 0.04025
R35386 VDD.n3139 VDD.n2908 0.04025
R35387 VDD.n3139 VDD.n3138 0.04025
R35388 VDD.n3138 VDD.n3137 0.04025
R35389 VDD.n3137 VDD.n2910 0.04025
R35390 VDD.n3133 VDD.n2910 0.04025
R35391 VDD.n3133 VDD.n3132 0.04025
R35392 VDD.n3132 VDD.n3131 0.04025
R35393 VDD.n3131 VDD.n2912 0.04025
R35394 VDD.n3127 VDD.n2912 0.04025
R35395 VDD.n3127 VDD.n3126 0.04025
R35396 VDD.n3126 VDD.n3125 0.04025
R35397 VDD.n3125 VDD.n2914 0.04025
R35398 VDD.n3121 VDD.n2914 0.04025
R35399 VDD.n3121 VDD.n3120 0.04025
R35400 VDD.n3120 VDD.n3119 0.04025
R35401 VDD.n3119 VDD.n2916 0.04025
R35402 VDD.n3115 VDD.n2916 0.04025
R35403 VDD.n3115 VDD.n3114 0.04025
R35404 VDD.n3114 VDD.n3113 0.04025
R35405 VDD.n3113 VDD.n2918 0.04025
R35406 VDD.n3109 VDD.n2918 0.04025
R35407 VDD.n3109 VDD.n3108 0.04025
R35408 VDD.n3108 VDD.n3107 0.04025
R35409 VDD.n3107 VDD.n2920 0.04025
R35410 VDD.n3103 VDD.n2920 0.04025
R35411 VDD.n3103 VDD.n3102 0.04025
R35412 VDD.n3102 VDD.n3101 0.04025
R35413 VDD.n3101 VDD.n2922 0.04025
R35414 VDD.n3097 VDD.n2922 0.04025
R35415 VDD.n3097 VDD.n3096 0.04025
R35416 VDD.n3096 VDD.n3095 0.04025
R35417 VDD.n3095 VDD.n2924 0.04025
R35418 VDD.n3091 VDD.n2924 0.04025
R35419 VDD.n3091 VDD.n3090 0.04025
R35420 VDD.n3090 VDD.n3089 0.04025
R35421 VDD.n3089 VDD.n2926 0.04025
R35422 VDD.n3085 VDD.n2926 0.04025
R35423 VDD.n3085 VDD.n3084 0.04025
R35424 VDD.n3084 VDD.n3083 0.04025
R35425 VDD.n3083 VDD.n2928 0.04025
R35426 VDD.n3079 VDD.n2928 0.04025
R35427 VDD.n3079 VDD.n3078 0.04025
R35428 VDD.n3078 VDD.n3077 0.04025
R35429 VDD.n3077 VDD.n2930 0.04025
R35430 VDD.n3073 VDD.n2930 0.04025
R35431 VDD.n3073 VDD.n3072 0.04025
R35432 VDD.n3072 VDD.n3071 0.04025
R35433 VDD.n3071 VDD.n2932 0.04025
R35434 VDD.n3067 VDD.n2932 0.04025
R35435 VDD.n3067 VDD.n3066 0.04025
R35436 VDD.n3066 VDD.n3065 0.04025
R35437 VDD.n3065 VDD.n2934 0.04025
R35438 VDD.n3061 VDD.n2934 0.04025
R35439 VDD.n3061 VDD.n3060 0.04025
R35440 VDD.n3060 VDD.n3059 0.04025
R35441 VDD.n3059 VDD.n2936 0.04025
R35442 VDD.n3055 VDD.n2936 0.04025
R35443 VDD.n3055 VDD.n3054 0.04025
R35444 VDD.n3054 VDD.n3053 0.04025
R35445 VDD.n3053 VDD.n2938 0.04025
R35446 VDD.n3049 VDD.n2938 0.04025
R35447 VDD.n3049 VDD.n3048 0.04025
R35448 VDD.n3048 VDD.n3047 0.04025
R35449 VDD.n3047 VDD.n2940 0.04025
R35450 VDD.n3043 VDD.n2940 0.04025
R35451 VDD.n3043 VDD.n3042 0.04025
R35452 VDD.n3042 VDD.n3041 0.04025
R35453 VDD.n3041 VDD.n2942 0.04025
R35454 VDD.n3037 VDD.n2942 0.04025
R35455 VDD.n3037 VDD.n3036 0.04025
R35456 VDD.n3036 VDD.n3035 0.04025
R35457 VDD.n3035 VDD.n2944 0.04025
R35458 VDD.n3031 VDD.n2944 0.04025
R35459 VDD.n3031 VDD.n3030 0.04025
R35460 VDD.n3030 VDD.n3029 0.04025
R35461 VDD.n3029 VDD.n2946 0.04025
R35462 VDD.n3025 VDD.n2946 0.04025
R35463 VDD.n3025 VDD.n3024 0.04025
R35464 VDD.n3024 VDD.n3023 0.04025
R35465 VDD.n3023 VDD.n2948 0.04025
R35466 VDD.n3019 VDD.n2948 0.04025
R35467 VDD.n3019 VDD.n3018 0.04025
R35468 VDD.n3018 VDD.n3017 0.04025
R35469 VDD.n3017 VDD.n2950 0.04025
R35470 VDD.n3013 VDD.n2950 0.04025
R35471 VDD.n3013 VDD.n3012 0.04025
R35472 VDD.n3012 VDD.n3011 0.04025
R35473 VDD.n3011 VDD.n2952 0.04025
R35474 VDD.n3007 VDD.n2952 0.04025
R35475 VDD.n3007 VDD.n3006 0.04025
R35476 VDD.n3006 VDD.n3005 0.04025
R35477 VDD.n3005 VDD.n2954 0.04025
R35478 VDD.n3001 VDD.n2954 0.04025
R35479 VDD.n3001 VDD.n3000 0.04025
R35480 VDD.n3000 VDD.n2999 0.04025
R35481 VDD.n2999 VDD.n2956 0.04025
R35482 VDD.n2995 VDD.n2956 0.04025
R35483 VDD.n2995 VDD.n2994 0.04025
R35484 VDD.n2994 VDD.n2993 0.04025
R35485 VDD.n2993 VDD.n2958 0.04025
R35486 VDD.n2989 VDD.n2958 0.04025
R35487 VDD.n2989 VDD.n2988 0.04025
R35488 VDD.n2988 VDD.n2987 0.04025
R35489 VDD.n2987 VDD.n2960 0.04025
R35490 VDD.n2983 VDD.n2960 0.04025
R35491 VDD.n2983 VDD.n2982 0.04025
R35492 VDD.n2982 VDD.n2981 0.04025
R35493 VDD.n2981 VDD.n2962 0.04025
R35494 VDD.n2977 VDD.n2962 0.04025
R35495 VDD.n2977 VDD.n2976 0.04025
R35496 VDD.n2976 VDD.n2975 0.04025
R35497 VDD.n2975 VDD.n2964 0.04025
R35498 VDD.n2971 VDD.n2964 0.04025
R35499 VDD.n2971 VDD.n2970 0.04025
R35500 VDD.n3631 VDD.n3630 0.04025
R35501 VDD.n3631 VDD.n2744 0.04025
R35502 VDD.n3635 VDD.n2744 0.04025
R35503 VDD.n3636 VDD.n3635 0.04025
R35504 VDD.n3637 VDD.n3636 0.04025
R35505 VDD.n3637 VDD.n2742 0.04025
R35506 VDD.n3641 VDD.n2742 0.04025
R35507 VDD.n3642 VDD.n3641 0.04025
R35508 VDD.n3643 VDD.n3642 0.04025
R35509 VDD.n3643 VDD.n2740 0.04025
R35510 VDD.n3647 VDD.n2740 0.04025
R35511 VDD.n3648 VDD.n3647 0.04025
R35512 VDD.n3649 VDD.n3648 0.04025
R35513 VDD.n3649 VDD.n2738 0.04025
R35514 VDD.n3653 VDD.n2738 0.04025
R35515 VDD.n3654 VDD.n3653 0.04025
R35516 VDD.n3655 VDD.n3654 0.04025
R35517 VDD.n3655 VDD.n2736 0.04025
R35518 VDD.n3659 VDD.n2736 0.04025
R35519 VDD.n3660 VDD.n3659 0.04025
R35520 VDD.n3661 VDD.n3660 0.04025
R35521 VDD.n3661 VDD.n2734 0.04025
R35522 VDD.n3665 VDD.n2734 0.04025
R35523 VDD.n3666 VDD.n3665 0.04025
R35524 VDD.n3667 VDD.n3666 0.04025
R35525 VDD.n3667 VDD.n2732 0.04025
R35526 VDD.n3671 VDD.n2732 0.04025
R35527 VDD.n3672 VDD.n3671 0.04025
R35528 VDD.n3673 VDD.n3672 0.04025
R35529 VDD.n3673 VDD.n2730 0.04025
R35530 VDD.n3677 VDD.n2730 0.04025
R35531 VDD.n3678 VDD.n3677 0.04025
R35532 VDD.n3679 VDD.n3678 0.04025
R35533 VDD.n3679 VDD.n2728 0.04025
R35534 VDD.n3683 VDD.n2728 0.04025
R35535 VDD.n3684 VDD.n3683 0.04025
R35536 VDD.n3685 VDD.n3684 0.04025
R35537 VDD.n3685 VDD.n2726 0.04025
R35538 VDD.n3689 VDD.n2726 0.04025
R35539 VDD.n3690 VDD.n3689 0.04025
R35540 VDD.n3691 VDD.n3690 0.04025
R35541 VDD.n3691 VDD.n2724 0.04025
R35542 VDD.n3695 VDD.n2724 0.04025
R35543 VDD.n3696 VDD.n3695 0.04025
R35544 VDD.n3697 VDD.n3696 0.04025
R35545 VDD.n3697 VDD.n2722 0.04025
R35546 VDD.n3701 VDD.n2722 0.04025
R35547 VDD.n3702 VDD.n3701 0.04025
R35548 VDD.n3703 VDD.n3702 0.04025
R35549 VDD.n3703 VDD.n2720 0.04025
R35550 VDD.n3707 VDD.n2720 0.04025
R35551 VDD.n3708 VDD.n3707 0.04025
R35552 VDD.n3709 VDD.n3708 0.04025
R35553 VDD.n3709 VDD.n2718 0.04025
R35554 VDD.n3713 VDD.n2718 0.04025
R35555 VDD.n3714 VDD.n3713 0.04025
R35556 VDD.n3715 VDD.n3714 0.04025
R35557 VDD.n3715 VDD.n2716 0.04025
R35558 VDD.n3719 VDD.n2716 0.04025
R35559 VDD.n3720 VDD.n3719 0.04025
R35560 VDD.n3721 VDD.n3720 0.04025
R35561 VDD.n3721 VDD.n2714 0.04025
R35562 VDD.n3725 VDD.n2714 0.04025
R35563 VDD.n3726 VDD.n3725 0.04025
R35564 VDD.n3727 VDD.n3726 0.04025
R35565 VDD.n3727 VDD.n2712 0.04025
R35566 VDD.n3731 VDD.n2712 0.04025
R35567 VDD.n3732 VDD.n3731 0.04025
R35568 VDD.n3733 VDD.n3732 0.04025
R35569 VDD.n3733 VDD.n2710 0.04025
R35570 VDD.n3737 VDD.n2710 0.04025
R35571 VDD.n3738 VDD.n3737 0.04025
R35572 VDD.n3739 VDD.n3738 0.04025
R35573 VDD.n3739 VDD.n2708 0.04025
R35574 VDD.n3743 VDD.n2708 0.04025
R35575 VDD.n3744 VDD.n3743 0.04025
R35576 VDD.n3745 VDD.n3744 0.04025
R35577 VDD.n3745 VDD.n2706 0.04025
R35578 VDD.n3749 VDD.n2706 0.04025
R35579 VDD.n3750 VDD.n3749 0.04025
R35580 VDD.n3751 VDD.n3750 0.04025
R35581 VDD.n3751 VDD.n2704 0.04025
R35582 VDD.n3755 VDD.n2704 0.04025
R35583 VDD.n3756 VDD.n3755 0.04025
R35584 VDD.n3757 VDD.n3756 0.04025
R35585 VDD.n3757 VDD.n2702 0.04025
R35586 VDD.n3761 VDD.n2702 0.04025
R35587 VDD.n3762 VDD.n3761 0.04025
R35588 VDD.n3763 VDD.n3762 0.04025
R35589 VDD.n3763 VDD.n2700 0.04025
R35590 VDD.n3767 VDD.n2700 0.04025
R35591 VDD.n3768 VDD.n3767 0.04025
R35592 VDD.n3769 VDD.n3768 0.04025
R35593 VDD.n3769 VDD.n2698 0.04025
R35594 VDD.n3773 VDD.n2698 0.04025
R35595 VDD.n3774 VDD.n3773 0.04025
R35596 VDD.n3775 VDD.n3774 0.04025
R35597 VDD.n3775 VDD.n2696 0.04025
R35598 VDD.n3779 VDD.n2696 0.04025
R35599 VDD.n3780 VDD.n3779 0.04025
R35600 VDD.n3781 VDD.n3780 0.04025
R35601 VDD.n3781 VDD.n2694 0.04025
R35602 VDD.n3785 VDD.n2694 0.04025
R35603 VDD.n3786 VDD.n3785 0.04025
R35604 VDD.n3787 VDD.n3786 0.04025
R35605 VDD.n3787 VDD.n2692 0.04025
R35606 VDD.n3791 VDD.n2692 0.04025
R35607 VDD.n3792 VDD.n3791 0.04025
R35608 VDD.n3793 VDD.n3792 0.04025
R35609 VDD.n3793 VDD.n2690 0.04025
R35610 VDD.n3797 VDD.n2690 0.04025
R35611 VDD.n3798 VDD.n3797 0.04025
R35612 VDD.n3799 VDD.n3798 0.04025
R35613 VDD.n3799 VDD.n2688 0.04025
R35614 VDD.n3803 VDD.n2688 0.04025
R35615 VDD.n3804 VDD.n3803 0.04025
R35616 VDD.n3805 VDD.n3804 0.04025
R35617 VDD.n3805 VDD.n2686 0.04025
R35618 VDD.n3809 VDD.n2686 0.04025
R35619 VDD.n3810 VDD.n3809 0.04025
R35620 VDD.n3811 VDD.n3810 0.04025
R35621 VDD.n3811 VDD.n2684 0.04025
R35622 VDD.n3815 VDD.n2684 0.04025
R35623 VDD.n3816 VDD.n3815 0.04025
R35624 VDD.n3817 VDD.n3816 0.04025
R35625 VDD.n3817 VDD.n2682 0.04025
R35626 VDD.n3821 VDD.n2682 0.04025
R35627 VDD.n3822 VDD.n3821 0.04025
R35628 VDD.n3823 VDD.n3822 0.04025
R35629 VDD.n3823 VDD.n2680 0.04025
R35630 VDD.n3827 VDD.n2680 0.04025
R35631 VDD.n3828 VDD.n3827 0.04025
R35632 VDD.n3829 VDD.n3828 0.04025
R35633 VDD.n3829 VDD.n2678 0.04025
R35634 VDD.n3833 VDD.n2678 0.04025
R35635 VDD.n3834 VDD.n3833 0.04025
R35636 VDD.n3835 VDD.n3834 0.04025
R35637 VDD.n3835 VDD.n2676 0.04025
R35638 VDD.n3839 VDD.n2676 0.04025
R35639 VDD.n3840 VDD.n3839 0.04025
R35640 VDD.n3841 VDD.n3840 0.04025
R35641 VDD.n3841 VDD.n2674 0.04025
R35642 VDD.n3845 VDD.n2674 0.04025
R35643 VDD.n3846 VDD.n3845 0.04025
R35644 VDD.n3847 VDD.n3846 0.04025
R35645 VDD.n3847 VDD.n2672 0.04025
R35646 VDD.n3851 VDD.n2672 0.04025
R35647 VDD.n3852 VDD.n3851 0.04025
R35648 VDD.n3853 VDD.n3852 0.04025
R35649 VDD.n3853 VDD.n2670 0.04025
R35650 VDD.n3857 VDD.n2670 0.04025
R35651 VDD.n3858 VDD.n3857 0.04025
R35652 VDD.n3859 VDD.n3858 0.04025
R35653 VDD.n3859 VDD.n2668 0.04025
R35654 VDD.n3863 VDD.n2668 0.04025
R35655 VDD.n3864 VDD.n3863 0.04025
R35656 VDD.n3865 VDD.n3864 0.04025
R35657 VDD.n3865 VDD.n2666 0.04025
R35658 VDD.n3869 VDD.n2666 0.04025
R35659 VDD.n3870 VDD.n3869 0.04025
R35660 VDD.n3871 VDD.n3870 0.04025
R35661 VDD.n3871 VDD.n2664 0.04025
R35662 VDD.n3875 VDD.n2664 0.04025
R35663 VDD.n3876 VDD.n3875 0.04025
R35664 VDD.n3877 VDD.n3876 0.04025
R35665 VDD.n3877 VDD.n2662 0.04025
R35666 VDD.n3881 VDD.n2662 0.04025
R35667 VDD.n3882 VDD.n3881 0.04025
R35668 VDD.n3883 VDD.n3882 0.04025
R35669 VDD.n3883 VDD.n2660 0.04025
R35670 VDD.n3887 VDD.n2660 0.04025
R35671 VDD.n3888 VDD.n3887 0.04025
R35672 VDD.n3889 VDD.n3888 0.04025
R35673 VDD.n3889 VDD.n2658 0.04025
R35674 VDD.n3893 VDD.n2658 0.04025
R35675 VDD.n3894 VDD.n3893 0.04025
R35676 VDD.n3895 VDD.n3894 0.04025
R35677 VDD.n3895 VDD.n2656 0.04025
R35678 VDD.n3899 VDD.n2656 0.04025
R35679 VDD.n3900 VDD.n3899 0.04025
R35680 VDD.n3901 VDD.n3900 0.04025
R35681 VDD.n3901 VDD.n2654 0.04025
R35682 VDD.n3905 VDD.n2654 0.04025
R35683 VDD.n3906 VDD.n3905 0.04025
R35684 VDD.n3907 VDD.n3906 0.04025
R35685 VDD.n3907 VDD.n2652 0.04025
R35686 VDD.n3911 VDD.n2652 0.04025
R35687 VDD.n3912 VDD.n3911 0.04025
R35688 VDD.n3913 VDD.n3912 0.04025
R35689 VDD.n3913 VDD.n2650 0.04025
R35690 VDD.n3917 VDD.n2650 0.04025
R35691 VDD.n3918 VDD.n3917 0.04025
R35692 VDD.n3919 VDD.n3918 0.04025
R35693 VDD.n3919 VDD.n2648 0.04025
R35694 VDD.n3923 VDD.n2648 0.04025
R35695 VDD.n3924 VDD.n3923 0.04025
R35696 VDD.n3925 VDD.n3924 0.04025
R35697 VDD.n3925 VDD.n2646 0.04025
R35698 VDD.n3929 VDD.n2646 0.04025
R35699 VDD.n3930 VDD.n3929 0.04025
R35700 VDD.n3931 VDD.n3930 0.04025
R35701 VDD.n3931 VDD.n2644 0.04025
R35702 VDD.n3935 VDD.n2644 0.04025
R35703 VDD.n3936 VDD.n3935 0.04025
R35704 VDD.n3937 VDD.n3936 0.04025
R35705 VDD.n3937 VDD.n2642 0.04025
R35706 VDD.n3941 VDD.n2642 0.04025
R35707 VDD.n3942 VDD.n3941 0.04025
R35708 VDD.n3943 VDD.n3942 0.04025
R35709 VDD.n3943 VDD.n2640 0.04025
R35710 VDD.n3947 VDD.n2640 0.04025
R35711 VDD.n3948 VDD.n3947 0.04025
R35712 VDD.n3949 VDD.n3948 0.04025
R35713 VDD.n3949 VDD.n2638 0.04025
R35714 VDD.n3953 VDD.n2638 0.04025
R35715 VDD.n3954 VDD.n3953 0.04025
R35716 VDD.n3955 VDD.n3954 0.04025
R35717 VDD.n3955 VDD.n2636 0.04025
R35718 VDD.n3959 VDD.n2636 0.04025
R35719 VDD.n3960 VDD.n3959 0.04025
R35720 VDD.n3961 VDD.n3960 0.04025
R35721 VDD.n3961 VDD.n2634 0.04025
R35722 VDD.n3965 VDD.n2634 0.04025
R35723 VDD.n3966 VDD.n3965 0.04025
R35724 VDD.n3967 VDD.n3966 0.04025
R35725 VDD.n3967 VDD.n2632 0.04025
R35726 VDD.n3971 VDD.n2632 0.04025
R35727 VDD.n3972 VDD.n3971 0.04025
R35728 VDD.n3973 VDD.n3972 0.04025
R35729 VDD.n3973 VDD.n2630 0.04025
R35730 VDD.n3977 VDD.n2630 0.04025
R35731 VDD.n3978 VDD.n3977 0.04025
R35732 VDD.n3979 VDD.n3978 0.04025
R35733 VDD.n3979 VDD.n2628 0.04025
R35734 VDD.n3983 VDD.n2628 0.04025
R35735 VDD.n3984 VDD.n3983 0.04025
R35736 VDD.n3985 VDD.n3984 0.04025
R35737 VDD.n3985 VDD.n2626 0.04025
R35738 VDD.n3989 VDD.n2626 0.04025
R35739 VDD.n3990 VDD.n3989 0.04025
R35740 VDD.n3991 VDD.n3990 0.04025
R35741 VDD.n3991 VDD.n2624 0.04025
R35742 VDD.n3995 VDD.n2624 0.04025
R35743 VDD.n3996 VDD.n3995 0.04025
R35744 VDD.n3997 VDD.n3996 0.04025
R35745 VDD.n3997 VDD.n2622 0.04025
R35746 VDD.n4001 VDD.n2622 0.04025
R35747 VDD.n4002 VDD.n4001 0.04025
R35748 VDD.n4003 VDD.n4002 0.04025
R35749 VDD.n4003 VDD.n2620 0.04025
R35750 VDD.n4007 VDD.n2620 0.04025
R35751 VDD.n4008 VDD.n4007 0.04025
R35752 VDD.n4009 VDD.n4008 0.04025
R35753 VDD.n4009 VDD.n2618 0.04025
R35754 VDD.n4013 VDD.n2618 0.04025
R35755 VDD.n4014 VDD.n4013 0.04025
R35756 VDD.n4015 VDD.n4014 0.04025
R35757 VDD.n4015 VDD.n2616 0.04025
R35758 VDD.n4019 VDD.n2616 0.04025
R35759 VDD.n4020 VDD.n4019 0.04025
R35760 VDD.n4021 VDD.n4020 0.04025
R35761 VDD.n4021 VDD.n2614 0.04025
R35762 VDD.n4025 VDD.n2614 0.04025
R35763 VDD.n4026 VDD.n4025 0.04025
R35764 VDD.n4027 VDD.n4026 0.04025
R35765 VDD.n4027 VDD.n2612 0.04025
R35766 VDD.n4031 VDD.n2612 0.04025
R35767 VDD.n4032 VDD.n4031 0.04025
R35768 VDD.n4033 VDD.n4032 0.04025
R35769 VDD.n4033 VDD.n2610 0.04025
R35770 VDD.n4037 VDD.n2610 0.04025
R35771 VDD.n4038 VDD.n4037 0.04025
R35772 VDD.n4039 VDD.n4038 0.04025
R35773 VDD.n4039 VDD.n2608 0.04025
R35774 VDD.n4043 VDD.n2608 0.04025
R35775 VDD.n4044 VDD.n4043 0.04025
R35776 VDD.n4045 VDD.n4044 0.04025
R35777 VDD.n4045 VDD.n2606 0.04025
R35778 VDD.n4049 VDD.n2606 0.04025
R35779 VDD.n4050 VDD.n4049 0.04025
R35780 VDD.n4051 VDD.n4050 0.04025
R35781 VDD.n4051 VDD.n2604 0.04025
R35782 VDD.n4055 VDD.n2604 0.04025
R35783 VDD.n4056 VDD.n4055 0.04025
R35784 VDD.n4057 VDD.n4056 0.04025
R35785 VDD.n4057 VDD.n2602 0.04025
R35786 VDD.n4061 VDD.n2602 0.04025
R35787 VDD.n4062 VDD.n4061 0.04025
R35788 VDD.n4063 VDD.n4062 0.04025
R35789 VDD.n4063 VDD.n2600 0.04025
R35790 VDD.n4067 VDD.n2600 0.04025
R35791 VDD.n4068 VDD.n4067 0.04025
R35792 VDD.n4069 VDD.n4068 0.04025
R35793 VDD.n4069 VDD.n2598 0.04025
R35794 VDD.n4073 VDD.n2598 0.04025
R35795 VDD.n4074 VDD.n4073 0.04025
R35796 VDD.n4075 VDD.n4074 0.04025
R35797 VDD.n4075 VDD.n2596 0.04025
R35798 VDD.n4079 VDD.n2596 0.04025
R35799 VDD.n4080 VDD.n4079 0.04025
R35800 VDD.n4081 VDD.n4080 0.04025
R35801 VDD.n4081 VDD.n2594 0.04025
R35802 VDD.n4085 VDD.n2594 0.04025
R35803 VDD.n4086 VDD.n4085 0.04025
R35804 VDD.n4087 VDD.n4086 0.04025
R35805 VDD.n4087 VDD.n2592 0.04025
R35806 VDD.n4091 VDD.n2592 0.04025
R35807 VDD.n4092 VDD.n4091 0.04025
R35808 VDD.n4093 VDD.n4092 0.04025
R35809 VDD.n4093 VDD.n2590 0.04025
R35810 VDD.n4097 VDD.n2590 0.04025
R35811 VDD.n4098 VDD.n4097 0.04025
R35812 VDD.n4099 VDD.n4098 0.04025
R35813 VDD.n4099 VDD.n2588 0.04025
R35814 VDD.n4103 VDD.n2588 0.04025
R35815 VDD.n4104 VDD.n4103 0.04025
R35816 VDD.n4105 VDD.n4104 0.04025
R35817 VDD.n4105 VDD.n2586 0.04025
R35818 VDD.n4109 VDD.n2586 0.04025
R35819 VDD.n4110 VDD.n4109 0.04025
R35820 VDD.n4111 VDD.n4110 0.04025
R35821 VDD.n4111 VDD.n2584 0.04025
R35822 VDD.n4115 VDD.n2584 0.04025
R35823 VDD.n4116 VDD.n4115 0.04025
R35824 VDD.n4117 VDD.n4116 0.04025
R35825 VDD.n4117 VDD.n2582 0.04025
R35826 VDD.n4121 VDD.n2582 0.04025
R35827 VDD.n4122 VDD.n4121 0.04025
R35828 VDD.n4123 VDD.n4122 0.04025
R35829 VDD.n4123 VDD.n2580 0.04025
R35830 VDD.n4127 VDD.n2580 0.04025
R35831 VDD.n4128 VDD.n4127 0.04025
R35832 VDD.n4129 VDD.n4128 0.04025
R35833 VDD.n4129 VDD.n2578 0.04025
R35834 VDD.n4133 VDD.n2578 0.04025
R35835 VDD.n4134 VDD.n4133 0.04025
R35836 VDD.n4135 VDD.n4134 0.04025
R35837 VDD.n4135 VDD.n2576 0.04025
R35838 VDD.n4139 VDD.n2576 0.04025
R35839 VDD.n4140 VDD.n4139 0.04025
R35840 VDD.n4141 VDD.n4140 0.04025
R35841 VDD.n4141 VDD.n2574 0.04025
R35842 VDD.n4145 VDD.n2574 0.04025
R35843 VDD.n4146 VDD.n4145 0.04025
R35844 VDD.n4147 VDD.n4146 0.04025
R35845 VDD.n4147 VDD.n2572 0.04025
R35846 VDD.n4151 VDD.n2572 0.04025
R35847 VDD.n4152 VDD.n4151 0.04025
R35848 VDD.n4153 VDD.n4152 0.04025
R35849 VDD.n4153 VDD.n2570 0.04025
R35850 VDD.n4157 VDD.n2570 0.04025
R35851 VDD.n4158 VDD.n4157 0.04025
R35852 VDD.n4159 VDD.n4158 0.04025
R35853 VDD.n4159 VDD.n2568 0.04025
R35854 VDD.n4163 VDD.n2568 0.04025
R35855 VDD.n4164 VDD.n4163 0.04025
R35856 VDD.n4165 VDD.n4164 0.04025
R35857 VDD.n4165 VDD.n2566 0.04025
R35858 VDD.n4169 VDD.n2566 0.04025
R35859 VDD.n4170 VDD.n4169 0.04025
R35860 VDD.n4171 VDD.n4170 0.04025
R35861 VDD.n4171 VDD.n2564 0.04025
R35862 VDD.n4175 VDD.n2564 0.04025
R35863 VDD.n4176 VDD.n4175 0.04025
R35864 VDD.n4177 VDD.n4176 0.04025
R35865 VDD.n4177 VDD.n2562 0.04025
R35866 VDD.n4181 VDD.n2562 0.04025
R35867 VDD.n4182 VDD.n4181 0.04025
R35868 VDD.n4183 VDD.n4182 0.04025
R35869 VDD.n4183 VDD.n2560 0.04025
R35870 VDD.n4187 VDD.n2560 0.04025
R35871 VDD.n4188 VDD.n4187 0.04025
R35872 VDD.n4189 VDD.n4188 0.04025
R35873 VDD.n4189 VDD.n2558 0.04025
R35874 VDD.n4193 VDD.n2558 0.04025
R35875 VDD.n4194 VDD.n4193 0.04025
R35876 VDD.n4195 VDD.n4194 0.04025
R35877 VDD.n4195 VDD.n2556 0.04025
R35878 VDD.n4199 VDD.n2556 0.04025
R35879 VDD.n4200 VDD.n4199 0.04025
R35880 VDD.n4201 VDD.n4200 0.04025
R35881 VDD.n4201 VDD.n2554 0.04025
R35882 VDD.n4205 VDD.n2554 0.04025
R35883 VDD.n4206 VDD.n4205 0.04025
R35884 VDD.n4207 VDD.n4206 0.04025
R35885 VDD.n4207 VDD.n2552 0.04025
R35886 VDD.n4211 VDD.n2552 0.04025
R35887 VDD.n4212 VDD.n4211 0.04025
R35888 VDD.n4213 VDD.n4212 0.04025
R35889 VDD.n4213 VDD.n2550 0.04025
R35890 VDD.n4217 VDD.n2550 0.04025
R35891 VDD.n4218 VDD.n4217 0.04025
R35892 VDD.n4219 VDD.n4218 0.04025
R35893 VDD.n4219 VDD.n2548 0.04025
R35894 VDD.n4223 VDD.n2548 0.04025
R35895 VDD.n4224 VDD.n4223 0.04025
R35896 VDD.n4225 VDD.n4224 0.04025
R35897 VDD.n4225 VDD.n2546 0.04025
R35898 VDD.n4229 VDD.n2546 0.04025
R35899 VDD.n4230 VDD.n4229 0.04025
R35900 VDD.n4231 VDD.n4230 0.04025
R35901 VDD.n4231 VDD.n2544 0.04025
R35902 VDD.n4235 VDD.n2544 0.04025
R35903 VDD.n4236 VDD.n4235 0.04025
R35904 VDD.n4237 VDD.n4236 0.04025
R35905 VDD.n4237 VDD.n2542 0.04025
R35906 VDD.n4241 VDD.n2542 0.04025
R35907 VDD.n4242 VDD.n4241 0.04025
R35908 VDD.n4243 VDD.n4242 0.04025
R35909 VDD.n4243 VDD.n2540 0.04025
R35910 VDD.n4247 VDD.n2540 0.04025
R35911 VDD.n4248 VDD.n4247 0.04025
R35912 VDD.n4249 VDD.n4248 0.04025
R35913 VDD.n4249 VDD.n2538 0.04025
R35914 VDD.n4253 VDD.n2538 0.04025
R35915 VDD.n4254 VDD.n4253 0.04025
R35916 VDD.n4255 VDD.n4254 0.04025
R35917 VDD.n4255 VDD.n2536 0.04025
R35918 VDD.n4259 VDD.n2536 0.04025
R35919 VDD.n4260 VDD.n4259 0.04025
R35920 VDD.n4261 VDD.n4260 0.04025
R35921 VDD.n4261 VDD.n2534 0.04025
R35922 VDD.n4265 VDD.n2534 0.04025
R35923 VDD.n4266 VDD.n4265 0.04025
R35924 VDD.n4267 VDD.n4266 0.04025
R35925 VDD.n4267 VDD.n2532 0.04025
R35926 VDD.n4271 VDD.n2532 0.04025
R35927 VDD.n4272 VDD.n4271 0.04025
R35928 VDD.n4273 VDD.n4272 0.04025
R35929 VDD.n4273 VDD.n2530 0.04025
R35930 VDD.n4277 VDD.n2530 0.04025
R35931 VDD.n4278 VDD.n4277 0.04025
R35932 VDD.n4279 VDD.n4278 0.04025
R35933 VDD.n4279 VDD.n2528 0.04025
R35934 VDD.n4283 VDD.n2528 0.04025
R35935 VDD.n4284 VDD.n4283 0.04025
R35936 VDD.n4285 VDD.n4284 0.04025
R35937 VDD.n4285 VDD.n2526 0.04025
R35938 VDD.n4289 VDD.n2526 0.04025
R35939 VDD.n4290 VDD.n4289 0.04025
R35940 VDD.n4291 VDD.n4290 0.04025
R35941 VDD.n4291 VDD.n2524 0.04025
R35942 VDD.n4295 VDD.n2524 0.04025
R35943 VDD.n4296 VDD.n4295 0.04025
R35944 VDD.n4297 VDD.n4296 0.04025
R35945 VDD.n4297 VDD.n2522 0.04025
R35946 VDD.n4301 VDD.n2522 0.04025
R35947 VDD.n4302 VDD.n4301 0.04025
R35948 VDD.n4303 VDD.n4302 0.04025
R35949 VDD.n4303 VDD.n2520 0.04025
R35950 VDD.n4307 VDD.n2520 0.04025
R35951 VDD.n4308 VDD.n4307 0.04025
R35952 VDD.n4309 VDD.n4308 0.04025
R35953 VDD.n4309 VDD.n2518 0.04025
R35954 VDD.n4313 VDD.n2518 0.04025
R35955 VDD.n4314 VDD.n4313 0.04025
R35956 VDD.n4315 VDD.n4314 0.04025
R35957 VDD.n4315 VDD.n2516 0.04025
R35958 VDD.n4319 VDD.n2516 0.04025
R35959 VDD.n4320 VDD.n4319 0.04025
R35960 VDD.n4321 VDD.n4320 0.04025
R35961 VDD.n4321 VDD.n2514 0.04025
R35962 VDD.n4325 VDD.n2514 0.04025
R35963 VDD.n4326 VDD.n4325 0.04025
R35964 VDD.n4327 VDD.n4326 0.04025
R35965 VDD.n4327 VDD.n2512 0.04025
R35966 VDD.n4331 VDD.n2512 0.04025
R35967 VDD.n4332 VDD.n4331 0.04025
R35968 VDD.n4333 VDD.n4332 0.04025
R35969 VDD.n4333 VDD.n2510 0.04025
R35970 VDD.n4337 VDD.n2510 0.04025
R35971 VDD.n4338 VDD.n4337 0.04025
R35972 VDD.n4339 VDD.n4338 0.04025
R35973 VDD.n4339 VDD.n2508 0.04025
R35974 VDD.n4343 VDD.n2508 0.04025
R35975 VDD.n4344 VDD.n4343 0.04025
R35976 VDD.n4345 VDD.n4344 0.04025
R35977 VDD.n4345 VDD.n2506 0.04025
R35978 VDD.n4349 VDD.n2506 0.04025
R35979 VDD.n4350 VDD.n4349 0.04025
R35980 VDD.n4351 VDD.n4350 0.04025
R35981 VDD.n4351 VDD.n2504 0.04025
R35982 VDD.n4355 VDD.n2504 0.04025
R35983 VDD.n4356 VDD.n4355 0.04025
R35984 VDD.n4357 VDD.n4356 0.04025
R35985 VDD.n4357 VDD.n2502 0.04025
R35986 VDD.n4361 VDD.n2502 0.04025
R35987 VDD.n4362 VDD.n4361 0.04025
R35988 VDD.n4363 VDD.n4362 0.04025
R35989 VDD.n4363 VDD.n2500 0.04025
R35990 VDD.n4367 VDD.n2500 0.04025
R35991 VDD.n4368 VDD.n4367 0.04025
R35992 VDD.n4369 VDD.n4368 0.04025
R35993 VDD.n4369 VDD.n2498 0.04025
R35994 VDD.n4373 VDD.n2498 0.04025
R35995 VDD.n4374 VDD.n4373 0.04025
R35996 VDD.n4375 VDD.n4374 0.04025
R35997 VDD.n4375 VDD.n2496 0.04025
R35998 VDD.n4379 VDD.n2496 0.04025
R35999 VDD.n4380 VDD.n4379 0.04025
R36000 VDD.n4381 VDD.n4380 0.04025
R36001 VDD.n4381 VDD.n2494 0.04025
R36002 VDD.n4385 VDD.n2494 0.04025
R36003 VDD.n4386 VDD.n4385 0.04025
R36004 VDD.n4387 VDD.n4386 0.04025
R36005 VDD.n4387 VDD.n2492 0.04025
R36006 VDD.n4391 VDD.n2492 0.04025
R36007 VDD.n4392 VDD.n4391 0.04025
R36008 VDD.n4393 VDD.n4392 0.04025
R36009 VDD.n4393 VDD.n2490 0.04025
R36010 VDD.n4397 VDD.n2490 0.04025
R36011 VDD.n4398 VDD.n4397 0.04025
R36012 VDD.n4399 VDD.n4398 0.04025
R36013 VDD.n4399 VDD.n2488 0.04025
R36014 VDD.n4403 VDD.n2488 0.04025
R36015 VDD.n4404 VDD.n4403 0.04025
R36016 VDD.n4405 VDD.n4404 0.04025
R36017 VDD.n4405 VDD.n2486 0.04025
R36018 VDD.n4409 VDD.n2486 0.04025
R36019 VDD.n4410 VDD.n4409 0.04025
R36020 VDD.n4411 VDD.n4410 0.04025
R36021 VDD.n4411 VDD.n2484 0.04025
R36022 VDD.n4415 VDD.n2484 0.04025
R36023 VDD.n4416 VDD.n4415 0.04025
R36024 VDD.n4417 VDD.n4416 0.04025
R36025 VDD.n4417 VDD.n2482 0.04025
R36026 VDD.n4421 VDD.n2482 0.04025
R36027 VDD.n4422 VDD.n4421 0.04025
R36028 VDD.n4423 VDD.n4422 0.04025
R36029 VDD.n4423 VDD.n2480 0.04025
R36030 VDD.n4427 VDD.n2480 0.04025
R36031 VDD.n4428 VDD.n4427 0.04025
R36032 VDD.n4429 VDD.n4428 0.04025
R36033 VDD.n4429 VDD.n2478 0.04025
R36034 VDD.n4433 VDD.n2478 0.04025
R36035 VDD.n4434 VDD.n4433 0.04025
R36036 VDD.n4435 VDD.n4434 0.04025
R36037 VDD.n4435 VDD.n2476 0.04025
R36038 VDD.n4439 VDD.n2476 0.04025
R36039 VDD.n4440 VDD.n4439 0.04025
R36040 VDD.n4441 VDD.n4440 0.04025
R36041 VDD.n4441 VDD.n2474 0.04025
R36042 VDD.n4445 VDD.n2474 0.04025
R36043 VDD.n4446 VDD.n4445 0.04025
R36044 VDD.n4447 VDD.n4446 0.04025
R36045 VDD.n4447 VDD.n2472 0.04025
R36046 VDD.n4451 VDD.n2472 0.04025
R36047 VDD.n4452 VDD.n4451 0.04025
R36048 VDD.n4453 VDD.n4452 0.04025
R36049 VDD.n4453 VDD.n2470 0.04025
R36050 VDD.n4457 VDD.n2470 0.04025
R36051 VDD.n4458 VDD.n4457 0.04025
R36052 VDD.n4459 VDD.n4458 0.04025
R36053 VDD.n4459 VDD.n2468 0.04025
R36054 VDD.n4463 VDD.n2468 0.04025
R36055 VDD.n4464 VDD.n4463 0.04025
R36056 VDD.n4465 VDD.n4464 0.04025
R36057 VDD.n4465 VDD.n2466 0.04025
R36058 VDD.n4469 VDD.n2466 0.04025
R36059 VDD.n4470 VDD.n4469 0.04025
R36060 VDD.n4471 VDD.n4470 0.04025
R36061 VDD.n4471 VDD.n2464 0.04025
R36062 VDD.n4475 VDD.n2464 0.04025
R36063 VDD.n4476 VDD.n4475 0.04025
R36064 VDD.n4477 VDD.n4476 0.04025
R36065 VDD.n4477 VDD.n2462 0.04025
R36066 VDD.n4481 VDD.n2462 0.04025
R36067 VDD.n4482 VDD.n4481 0.04025
R36068 VDD.n4483 VDD.n4482 0.04025
R36069 VDD.n4483 VDD.n2460 0.04025
R36070 VDD.n4487 VDD.n2460 0.04025
R36071 VDD.n4488 VDD.n4487 0.04025
R36072 VDD.n4489 VDD.n4488 0.04025
R36073 VDD.n4489 VDD.n2458 0.04025
R36074 VDD.n4493 VDD.n2458 0.04025
R36075 VDD.n4494 VDD.n4493 0.04025
R36076 VDD.n4495 VDD.n4494 0.04025
R36077 VDD.n4495 VDD.n2456 0.04025
R36078 VDD.n4499 VDD.n2456 0.04025
R36079 VDD.n4500 VDD.n4499 0.04025
R36080 VDD.n4501 VDD.n4500 0.04025
R36081 VDD.n4501 VDD.n2454 0.04025
R36082 VDD.n4505 VDD.n2454 0.04025
R36083 VDD.n4506 VDD.n4505 0.04025
R36084 VDD.n4507 VDD.n4506 0.04025
R36085 VDD.n4507 VDD.n2452 0.04025
R36086 VDD.n4511 VDD.n2452 0.04025
R36087 VDD.n4512 VDD.n4511 0.04025
R36088 VDD.n4513 VDD.n4512 0.04025
R36089 VDD.n4513 VDD.n2450 0.04025
R36090 VDD.n4517 VDD.n2450 0.04025
R36091 VDD.n4518 VDD.n4517 0.04025
R36092 VDD.n4519 VDD.n4518 0.04025
R36093 VDD.n4519 VDD.n2448 0.04025
R36094 VDD.n4523 VDD.n2448 0.04025
R36095 VDD.n4524 VDD.n4523 0.04025
R36096 VDD.n4525 VDD.n4524 0.04025
R36097 VDD.n4525 VDD.n2446 0.04025
R36098 VDD.n4529 VDD.n2446 0.04025
R36099 VDD.n4530 VDD.n4529 0.04025
R36100 VDD.n4531 VDD.n4530 0.04025
R36101 VDD.n4531 VDD.n2444 0.04025
R36102 VDD.n4535 VDD.n2444 0.04025
R36103 VDD.n4536 VDD.n4535 0.04025
R36104 VDD.n4537 VDD.n4536 0.04025
R36105 VDD.n4537 VDD.n2442 0.04025
R36106 VDD.n4541 VDD.n2442 0.04025
R36107 VDD.n4542 VDD.n4541 0.04025
R36108 VDD.n4543 VDD.n4542 0.04025
R36109 VDD.n4543 VDD.n2440 0.04025
R36110 VDD.n4547 VDD.n2440 0.04025
R36111 VDD.n4548 VDD.n4547 0.04025
R36112 VDD.n4549 VDD.n4548 0.04025
R36113 VDD.n4549 VDD.n2438 0.04025
R36114 VDD.n4553 VDD.n2438 0.04025
R36115 VDD.n4554 VDD.n4553 0.04025
R36116 VDD.n4555 VDD.n4554 0.04025
R36117 VDD.n4555 VDD.n2436 0.04025
R36118 VDD.n4559 VDD.n2436 0.04025
R36119 VDD.n4560 VDD.n4559 0.04025
R36120 VDD.n4561 VDD.n4560 0.04025
R36121 VDD.n4561 VDD.n2434 0.04025
R36122 VDD.n4565 VDD.n2434 0.04025
R36123 VDD.n4566 VDD.n4565 0.04025
R36124 VDD.n4567 VDD.n4566 0.04025
R36125 VDD.n4567 VDD.n2432 0.04025
R36126 VDD.n4571 VDD.n2432 0.04025
R36127 VDD.n4572 VDD.n4571 0.04025
R36128 VDD.n4573 VDD.n4572 0.04025
R36129 VDD.n4573 VDD.n2430 0.04025
R36130 VDD.n4577 VDD.n2430 0.04025
R36131 VDD.n4578 VDD.n4577 0.04025
R36132 VDD.n4579 VDD.n4578 0.04025
R36133 VDD.n4579 VDD.n2428 0.04025
R36134 VDD.n4583 VDD.n2428 0.04025
R36135 VDD.n4584 VDD.n4583 0.04025
R36136 VDD.n4585 VDD.n4584 0.04025
R36137 VDD.n4585 VDD.n2426 0.04025
R36138 VDD.n4589 VDD.n2426 0.04025
R36139 VDD.n3632 VDD.n2745 0.04025
R36140 VDD.n3633 VDD.n3632 0.04025
R36141 VDD.n3634 VDD.n3633 0.04025
R36142 VDD.n3634 VDD.n2743 0.04025
R36143 VDD.n3638 VDD.n2743 0.04025
R36144 VDD.n3639 VDD.n3638 0.04025
R36145 VDD.n3640 VDD.n3639 0.04025
R36146 VDD.n3640 VDD.n2741 0.04025
R36147 VDD.n3644 VDD.n2741 0.04025
R36148 VDD.n3645 VDD.n3644 0.04025
R36149 VDD.n3646 VDD.n3645 0.04025
R36150 VDD.n3646 VDD.n2739 0.04025
R36151 VDD.n3650 VDD.n2739 0.04025
R36152 VDD.n3651 VDD.n3650 0.04025
R36153 VDD.n3652 VDD.n3651 0.04025
R36154 VDD.n3652 VDD.n2737 0.04025
R36155 VDD.n3656 VDD.n2737 0.04025
R36156 VDD.n3657 VDD.n3656 0.04025
R36157 VDD.n3658 VDD.n3657 0.04025
R36158 VDD.n3658 VDD.n2735 0.04025
R36159 VDD.n3662 VDD.n2735 0.04025
R36160 VDD.n3663 VDD.n3662 0.04025
R36161 VDD.n3664 VDD.n3663 0.04025
R36162 VDD.n3664 VDD.n2733 0.04025
R36163 VDD.n3668 VDD.n2733 0.04025
R36164 VDD.n3669 VDD.n3668 0.04025
R36165 VDD.n3670 VDD.n3669 0.04025
R36166 VDD.n3670 VDD.n2731 0.04025
R36167 VDD.n3674 VDD.n2731 0.04025
R36168 VDD.n3675 VDD.n3674 0.04025
R36169 VDD.n3676 VDD.n3675 0.04025
R36170 VDD.n3676 VDD.n2729 0.04025
R36171 VDD.n3680 VDD.n2729 0.04025
R36172 VDD.n3681 VDD.n3680 0.04025
R36173 VDD.n3682 VDD.n3681 0.04025
R36174 VDD.n3682 VDD.n2727 0.04025
R36175 VDD.n3686 VDD.n2727 0.04025
R36176 VDD.n3687 VDD.n3686 0.04025
R36177 VDD.n3688 VDD.n3687 0.04025
R36178 VDD.n3688 VDD.n2725 0.04025
R36179 VDD.n3692 VDD.n2725 0.04025
R36180 VDD.n3693 VDD.n3692 0.04025
R36181 VDD.n3694 VDD.n3693 0.04025
R36182 VDD.n3694 VDD.n2723 0.04025
R36183 VDD.n3698 VDD.n2723 0.04025
R36184 VDD.n3699 VDD.n3698 0.04025
R36185 VDD.n3700 VDD.n3699 0.04025
R36186 VDD.n3700 VDD.n2721 0.04025
R36187 VDD.n3704 VDD.n2721 0.04025
R36188 VDD.n3705 VDD.n3704 0.04025
R36189 VDD.n3706 VDD.n3705 0.04025
R36190 VDD.n3706 VDD.n2719 0.04025
R36191 VDD.n3710 VDD.n2719 0.04025
R36192 VDD.n3711 VDD.n3710 0.04025
R36193 VDD.n3712 VDD.n3711 0.04025
R36194 VDD.n3712 VDD.n2717 0.04025
R36195 VDD.n3716 VDD.n2717 0.04025
R36196 VDD.n3717 VDD.n3716 0.04025
R36197 VDD.n3718 VDD.n3717 0.04025
R36198 VDD.n3718 VDD.n2715 0.04025
R36199 VDD.n3722 VDD.n2715 0.04025
R36200 VDD.n3723 VDD.n3722 0.04025
R36201 VDD.n3724 VDD.n3723 0.04025
R36202 VDD.n3724 VDD.n2713 0.04025
R36203 VDD.n3728 VDD.n2713 0.04025
R36204 VDD.n3729 VDD.n3728 0.04025
R36205 VDD.n3730 VDD.n3729 0.04025
R36206 VDD.n3730 VDD.n2711 0.04025
R36207 VDD.n3734 VDD.n2711 0.04025
R36208 VDD.n3735 VDD.n3734 0.04025
R36209 VDD.n3736 VDD.n3735 0.04025
R36210 VDD.n3736 VDD.n2709 0.04025
R36211 VDD.n3740 VDD.n2709 0.04025
R36212 VDD.n3741 VDD.n3740 0.04025
R36213 VDD.n3742 VDD.n3741 0.04025
R36214 VDD.n3742 VDD.n2707 0.04025
R36215 VDD.n3746 VDD.n2707 0.04025
R36216 VDD.n3747 VDD.n3746 0.04025
R36217 VDD.n3748 VDD.n3747 0.04025
R36218 VDD.n3748 VDD.n2705 0.04025
R36219 VDD.n3752 VDD.n2705 0.04025
R36220 VDD.n3753 VDD.n3752 0.04025
R36221 VDD.n3754 VDD.n3753 0.04025
R36222 VDD.n3754 VDD.n2703 0.04025
R36223 VDD.n3758 VDD.n2703 0.04025
R36224 VDD.n3759 VDD.n3758 0.04025
R36225 VDD.n3760 VDD.n3759 0.04025
R36226 VDD.n3760 VDD.n2701 0.04025
R36227 VDD.n3764 VDD.n2701 0.04025
R36228 VDD.n3765 VDD.n3764 0.04025
R36229 VDD.n3766 VDD.n3765 0.04025
R36230 VDD.n3766 VDD.n2699 0.04025
R36231 VDD.n3770 VDD.n2699 0.04025
R36232 VDD.n3771 VDD.n3770 0.04025
R36233 VDD.n3772 VDD.n3771 0.04025
R36234 VDD.n3772 VDD.n2697 0.04025
R36235 VDD.n3776 VDD.n2697 0.04025
R36236 VDD.n3777 VDD.n3776 0.04025
R36237 VDD.n3778 VDD.n3777 0.04025
R36238 VDD.n3778 VDD.n2695 0.04025
R36239 VDD.n3782 VDD.n2695 0.04025
R36240 VDD.n3783 VDD.n3782 0.04025
R36241 VDD.n3784 VDD.n3783 0.04025
R36242 VDD.n3784 VDD.n2693 0.04025
R36243 VDD.n3788 VDD.n2693 0.04025
R36244 VDD.n3789 VDD.n3788 0.04025
R36245 VDD.n3790 VDD.n3789 0.04025
R36246 VDD.n3790 VDD.n2691 0.04025
R36247 VDD.n3794 VDD.n2691 0.04025
R36248 VDD.n3795 VDD.n3794 0.04025
R36249 VDD.n3796 VDD.n3795 0.04025
R36250 VDD.n3796 VDD.n2689 0.04025
R36251 VDD.n3800 VDD.n2689 0.04025
R36252 VDD.n3801 VDD.n3800 0.04025
R36253 VDD.n3802 VDD.n3801 0.04025
R36254 VDD.n3802 VDD.n2687 0.04025
R36255 VDD.n3806 VDD.n2687 0.04025
R36256 VDD.n3807 VDD.n3806 0.04025
R36257 VDD.n3808 VDD.n3807 0.04025
R36258 VDD.n3808 VDD.n2685 0.04025
R36259 VDD.n3812 VDD.n2685 0.04025
R36260 VDD.n3813 VDD.n3812 0.04025
R36261 VDD.n3814 VDD.n3813 0.04025
R36262 VDD.n3814 VDD.n2683 0.04025
R36263 VDD.n3818 VDD.n2683 0.04025
R36264 VDD.n3819 VDD.n3818 0.04025
R36265 VDD.n3820 VDD.n3819 0.04025
R36266 VDD.n3820 VDD.n2681 0.04025
R36267 VDD.n3824 VDD.n2681 0.04025
R36268 VDD.n3825 VDD.n3824 0.04025
R36269 VDD.n3826 VDD.n3825 0.04025
R36270 VDD.n3826 VDD.n2679 0.04025
R36271 VDD.n3830 VDD.n2679 0.04025
R36272 VDD.n3831 VDD.n3830 0.04025
R36273 VDD.n3832 VDD.n3831 0.04025
R36274 VDD.n3832 VDD.n2677 0.04025
R36275 VDD.n3836 VDD.n2677 0.04025
R36276 VDD.n3837 VDD.n3836 0.04025
R36277 VDD.n3838 VDD.n3837 0.04025
R36278 VDD.n3838 VDD.n2675 0.04025
R36279 VDD.n3842 VDD.n2675 0.04025
R36280 VDD.n3843 VDD.n3842 0.04025
R36281 VDD.n3844 VDD.n3843 0.04025
R36282 VDD.n3844 VDD.n2673 0.04025
R36283 VDD.n3848 VDD.n2673 0.04025
R36284 VDD.n3849 VDD.n3848 0.04025
R36285 VDD.n3850 VDD.n3849 0.04025
R36286 VDD.n3850 VDD.n2671 0.04025
R36287 VDD.n3854 VDD.n2671 0.04025
R36288 VDD.n3855 VDD.n3854 0.04025
R36289 VDD.n3856 VDD.n3855 0.04025
R36290 VDD.n3856 VDD.n2669 0.04025
R36291 VDD.n3860 VDD.n2669 0.04025
R36292 VDD.n3861 VDD.n3860 0.04025
R36293 VDD.n3862 VDD.n3861 0.04025
R36294 VDD.n3862 VDD.n2667 0.04025
R36295 VDD.n3866 VDD.n2667 0.04025
R36296 VDD.n3867 VDD.n3866 0.04025
R36297 VDD.n3868 VDD.n3867 0.04025
R36298 VDD.n3868 VDD.n2665 0.04025
R36299 VDD.n3872 VDD.n2665 0.04025
R36300 VDD.n3873 VDD.n3872 0.04025
R36301 VDD.n3874 VDD.n3873 0.04025
R36302 VDD.n3874 VDD.n2663 0.04025
R36303 VDD.n3878 VDD.n2663 0.04025
R36304 VDD.n3879 VDD.n3878 0.04025
R36305 VDD.n3880 VDD.n3879 0.04025
R36306 VDD.n3880 VDD.n2661 0.04025
R36307 VDD.n3884 VDD.n2661 0.04025
R36308 VDD.n3885 VDD.n3884 0.04025
R36309 VDD.n3886 VDD.n3885 0.04025
R36310 VDD.n3886 VDD.n2659 0.04025
R36311 VDD.n3890 VDD.n2659 0.04025
R36312 VDD.n3891 VDD.n3890 0.04025
R36313 VDD.n3892 VDD.n3891 0.04025
R36314 VDD.n3892 VDD.n2657 0.04025
R36315 VDD.n3896 VDD.n2657 0.04025
R36316 VDD.n3897 VDD.n3896 0.04025
R36317 VDD.n3898 VDD.n3897 0.04025
R36318 VDD.n3898 VDD.n2655 0.04025
R36319 VDD.n3902 VDD.n2655 0.04025
R36320 VDD.n3903 VDD.n3902 0.04025
R36321 VDD.n3904 VDD.n3903 0.04025
R36322 VDD.n3904 VDD.n2653 0.04025
R36323 VDD.n3908 VDD.n2653 0.04025
R36324 VDD.n3909 VDD.n3908 0.04025
R36325 VDD.n3910 VDD.n3909 0.04025
R36326 VDD.n3910 VDD.n2651 0.04025
R36327 VDD.n3914 VDD.n2651 0.04025
R36328 VDD.n3915 VDD.n3914 0.04025
R36329 VDD.n3916 VDD.n3915 0.04025
R36330 VDD.n3916 VDD.n2649 0.04025
R36331 VDD.n3920 VDD.n2649 0.04025
R36332 VDD.n3921 VDD.n3920 0.04025
R36333 VDD.n3922 VDD.n3921 0.04025
R36334 VDD.n3922 VDD.n2647 0.04025
R36335 VDD.n3926 VDD.n2647 0.04025
R36336 VDD.n3927 VDD.n3926 0.04025
R36337 VDD.n3928 VDD.n3927 0.04025
R36338 VDD.n3928 VDD.n2645 0.04025
R36339 VDD.n3932 VDD.n2645 0.04025
R36340 VDD.n3933 VDD.n3932 0.04025
R36341 VDD.n3934 VDD.n3933 0.04025
R36342 VDD.n3934 VDD.n2643 0.04025
R36343 VDD.n3938 VDD.n2643 0.04025
R36344 VDD.n3939 VDD.n3938 0.04025
R36345 VDD.n3940 VDD.n3939 0.04025
R36346 VDD.n3940 VDD.n2641 0.04025
R36347 VDD.n3944 VDD.n2641 0.04025
R36348 VDD.n3945 VDD.n3944 0.04025
R36349 VDD.n3946 VDD.n3945 0.04025
R36350 VDD.n3946 VDD.n2639 0.04025
R36351 VDD.n3950 VDD.n2639 0.04025
R36352 VDD.n3951 VDD.n3950 0.04025
R36353 VDD.n3952 VDD.n3951 0.04025
R36354 VDD.n3952 VDD.n2637 0.04025
R36355 VDD.n3956 VDD.n2637 0.04025
R36356 VDD.n3957 VDD.n3956 0.04025
R36357 VDD.n3958 VDD.n3957 0.04025
R36358 VDD.n3958 VDD.n2635 0.04025
R36359 VDD.n3962 VDD.n2635 0.04025
R36360 VDD.n3963 VDD.n3962 0.04025
R36361 VDD.n3964 VDD.n3963 0.04025
R36362 VDD.n3964 VDD.n2633 0.04025
R36363 VDD.n3968 VDD.n2633 0.04025
R36364 VDD.n3969 VDD.n3968 0.04025
R36365 VDD.n3970 VDD.n3969 0.04025
R36366 VDD.n3970 VDD.n2631 0.04025
R36367 VDD.n3974 VDD.n2631 0.04025
R36368 VDD.n3975 VDD.n3974 0.04025
R36369 VDD.n3976 VDD.n3975 0.04025
R36370 VDD.n3976 VDD.n2629 0.04025
R36371 VDD.n3980 VDD.n2629 0.04025
R36372 VDD.n3981 VDD.n3980 0.04025
R36373 VDD.n3982 VDD.n3981 0.04025
R36374 VDD.n3982 VDD.n2627 0.04025
R36375 VDD.n3986 VDD.n2627 0.04025
R36376 VDD.n3987 VDD.n3986 0.04025
R36377 VDD.n3988 VDD.n3987 0.04025
R36378 VDD.n3988 VDD.n2625 0.04025
R36379 VDD.n3992 VDD.n2625 0.04025
R36380 VDD.n3993 VDD.n3992 0.04025
R36381 VDD.n3994 VDD.n3993 0.04025
R36382 VDD.n3994 VDD.n2623 0.04025
R36383 VDD.n3998 VDD.n2623 0.04025
R36384 VDD.n3999 VDD.n3998 0.04025
R36385 VDD.n4000 VDD.n3999 0.04025
R36386 VDD.n4000 VDD.n2621 0.04025
R36387 VDD.n4004 VDD.n2621 0.04025
R36388 VDD.n4005 VDD.n4004 0.04025
R36389 VDD.n4006 VDD.n4005 0.04025
R36390 VDD.n4006 VDD.n2619 0.04025
R36391 VDD.n4010 VDD.n2619 0.04025
R36392 VDD.n4011 VDD.n4010 0.04025
R36393 VDD.n4012 VDD.n4011 0.04025
R36394 VDD.n4012 VDD.n2617 0.04025
R36395 VDD.n4016 VDD.n2617 0.04025
R36396 VDD.n4017 VDD.n4016 0.04025
R36397 VDD.n4018 VDD.n4017 0.04025
R36398 VDD.n4018 VDD.n2615 0.04025
R36399 VDD.n4022 VDD.n2615 0.04025
R36400 VDD.n4023 VDD.n4022 0.04025
R36401 VDD.n4024 VDD.n4023 0.04025
R36402 VDD.n4024 VDD.n2613 0.04025
R36403 VDD.n4028 VDD.n2613 0.04025
R36404 VDD.n4029 VDD.n4028 0.04025
R36405 VDD.n4030 VDD.n4029 0.04025
R36406 VDD.n4030 VDD.n2611 0.04025
R36407 VDD.n4034 VDD.n2611 0.04025
R36408 VDD.n4035 VDD.n4034 0.04025
R36409 VDD.n4036 VDD.n4035 0.04025
R36410 VDD.n4036 VDD.n2609 0.04025
R36411 VDD.n4040 VDD.n2609 0.04025
R36412 VDD.n4041 VDD.n4040 0.04025
R36413 VDD.n4042 VDD.n4041 0.04025
R36414 VDD.n4042 VDD.n2607 0.04025
R36415 VDD.n4046 VDD.n2607 0.04025
R36416 VDD.n4047 VDD.n4046 0.04025
R36417 VDD.n4048 VDD.n4047 0.04025
R36418 VDD.n4048 VDD.n2605 0.04025
R36419 VDD.n4052 VDD.n2605 0.04025
R36420 VDD.n4053 VDD.n4052 0.04025
R36421 VDD.n4054 VDD.n4053 0.04025
R36422 VDD.n4054 VDD.n2603 0.04025
R36423 VDD.n4058 VDD.n2603 0.04025
R36424 VDD.n4059 VDD.n4058 0.04025
R36425 VDD.n4060 VDD.n4059 0.04025
R36426 VDD.n4060 VDD.n2601 0.04025
R36427 VDD.n4064 VDD.n2601 0.04025
R36428 VDD.n4065 VDD.n4064 0.04025
R36429 VDD.n4066 VDD.n4065 0.04025
R36430 VDD.n4066 VDD.n2599 0.04025
R36431 VDD.n4070 VDD.n2599 0.04025
R36432 VDD.n4071 VDD.n4070 0.04025
R36433 VDD.n4072 VDD.n4071 0.04025
R36434 VDD.n4072 VDD.n2597 0.04025
R36435 VDD.n4076 VDD.n2597 0.04025
R36436 VDD.n4077 VDD.n4076 0.04025
R36437 VDD.n4078 VDD.n4077 0.04025
R36438 VDD.n4078 VDD.n2595 0.04025
R36439 VDD.n4082 VDD.n2595 0.04025
R36440 VDD.n4083 VDD.n4082 0.04025
R36441 VDD.n4084 VDD.n4083 0.04025
R36442 VDD.n4084 VDD.n2593 0.04025
R36443 VDD.n4088 VDD.n2593 0.04025
R36444 VDD.n4089 VDD.n4088 0.04025
R36445 VDD.n4090 VDD.n4089 0.04025
R36446 VDD.n4090 VDD.n2591 0.04025
R36447 VDD.n4094 VDD.n2591 0.04025
R36448 VDD.n4095 VDD.n4094 0.04025
R36449 VDD.n4096 VDD.n4095 0.04025
R36450 VDD.n4096 VDD.n2589 0.04025
R36451 VDD.n4100 VDD.n2589 0.04025
R36452 VDD.n4101 VDD.n4100 0.04025
R36453 VDD.n4102 VDD.n4101 0.04025
R36454 VDD.n4102 VDD.n2587 0.04025
R36455 VDD.n4106 VDD.n2587 0.04025
R36456 VDD.n4107 VDD.n4106 0.04025
R36457 VDD.n4108 VDD.n4107 0.04025
R36458 VDD.n4108 VDD.n2585 0.04025
R36459 VDD.n4112 VDD.n2585 0.04025
R36460 VDD.n4113 VDD.n4112 0.04025
R36461 VDD.n4114 VDD.n4113 0.04025
R36462 VDD.n4114 VDD.n2583 0.04025
R36463 VDD.n4118 VDD.n2583 0.04025
R36464 VDD.n4119 VDD.n4118 0.04025
R36465 VDD.n4120 VDD.n4119 0.04025
R36466 VDD.n4120 VDD.n2581 0.04025
R36467 VDD.n4124 VDD.n2581 0.04025
R36468 VDD.n4125 VDD.n4124 0.04025
R36469 VDD.n4126 VDD.n4125 0.04025
R36470 VDD.n4126 VDD.n2579 0.04025
R36471 VDD.n4130 VDD.n2579 0.04025
R36472 VDD.n4131 VDD.n4130 0.04025
R36473 VDD.n4132 VDD.n4131 0.04025
R36474 VDD.n4132 VDD.n2577 0.04025
R36475 VDD.n4136 VDD.n2577 0.04025
R36476 VDD.n4137 VDD.n4136 0.04025
R36477 VDD.n4138 VDD.n4137 0.04025
R36478 VDD.n4138 VDD.n2575 0.04025
R36479 VDD.n4142 VDD.n2575 0.04025
R36480 VDD.n4143 VDD.n4142 0.04025
R36481 VDD.n4144 VDD.n4143 0.04025
R36482 VDD.n4144 VDD.n2573 0.04025
R36483 VDD.n4148 VDD.n2573 0.04025
R36484 VDD.n4149 VDD.n4148 0.04025
R36485 VDD.n4150 VDD.n4149 0.04025
R36486 VDD.n4150 VDD.n2571 0.04025
R36487 VDD.n4154 VDD.n2571 0.04025
R36488 VDD.n4155 VDD.n4154 0.04025
R36489 VDD.n4156 VDD.n4155 0.04025
R36490 VDD.n4156 VDD.n2569 0.04025
R36491 VDD.n4160 VDD.n2569 0.04025
R36492 VDD.n4161 VDD.n4160 0.04025
R36493 VDD.n4162 VDD.n4161 0.04025
R36494 VDD.n4162 VDD.n2567 0.04025
R36495 VDD.n4166 VDD.n2567 0.04025
R36496 VDD.n4167 VDD.n4166 0.04025
R36497 VDD.n4168 VDD.n4167 0.04025
R36498 VDD.n4168 VDD.n2565 0.04025
R36499 VDD.n4172 VDD.n2565 0.04025
R36500 VDD.n4173 VDD.n4172 0.04025
R36501 VDD.n4174 VDD.n4173 0.04025
R36502 VDD.n4174 VDD.n2563 0.04025
R36503 VDD.n4178 VDD.n2563 0.04025
R36504 VDD.n4179 VDD.n4178 0.04025
R36505 VDD.n4180 VDD.n4179 0.04025
R36506 VDD.n4180 VDD.n2561 0.04025
R36507 VDD.n4184 VDD.n2561 0.04025
R36508 VDD.n4185 VDD.n4184 0.04025
R36509 VDD.n4186 VDD.n4185 0.04025
R36510 VDD.n4186 VDD.n2559 0.04025
R36511 VDD.n4190 VDD.n2559 0.04025
R36512 VDD.n4191 VDD.n4190 0.04025
R36513 VDD.n4192 VDD.n4191 0.04025
R36514 VDD.n4192 VDD.n2557 0.04025
R36515 VDD.n4196 VDD.n2557 0.04025
R36516 VDD.n4197 VDD.n4196 0.04025
R36517 VDD.n4198 VDD.n4197 0.04025
R36518 VDD.n4198 VDD.n2555 0.04025
R36519 VDD.n4202 VDD.n2555 0.04025
R36520 VDD.n4203 VDD.n4202 0.04025
R36521 VDD.n4204 VDD.n4203 0.04025
R36522 VDD.n4204 VDD.n2553 0.04025
R36523 VDD.n4208 VDD.n2553 0.04025
R36524 VDD.n4209 VDD.n4208 0.04025
R36525 VDD.n4210 VDD.n4209 0.04025
R36526 VDD.n4210 VDD.n2551 0.04025
R36527 VDD.n4214 VDD.n2551 0.04025
R36528 VDD.n4215 VDD.n4214 0.04025
R36529 VDD.n4216 VDD.n4215 0.04025
R36530 VDD.n4216 VDD.n2549 0.04025
R36531 VDD.n4220 VDD.n2549 0.04025
R36532 VDD.n4221 VDD.n4220 0.04025
R36533 VDD.n4222 VDD.n4221 0.04025
R36534 VDD.n4222 VDD.n2547 0.04025
R36535 VDD.n4226 VDD.n2547 0.04025
R36536 VDD.n4227 VDD.n4226 0.04025
R36537 VDD.n4228 VDD.n4227 0.04025
R36538 VDD.n4228 VDD.n2545 0.04025
R36539 VDD.n4232 VDD.n2545 0.04025
R36540 VDD.n4233 VDD.n4232 0.04025
R36541 VDD.n4234 VDD.n4233 0.04025
R36542 VDD.n4234 VDD.n2543 0.04025
R36543 VDD.n4238 VDD.n2543 0.04025
R36544 VDD.n4239 VDD.n4238 0.04025
R36545 VDD.n4240 VDD.n4239 0.04025
R36546 VDD.n4240 VDD.n2541 0.04025
R36547 VDD.n4244 VDD.n2541 0.04025
R36548 VDD.n4245 VDD.n4244 0.04025
R36549 VDD.n4246 VDD.n4245 0.04025
R36550 VDD.n4246 VDD.n2539 0.04025
R36551 VDD.n4250 VDD.n2539 0.04025
R36552 VDD.n4251 VDD.n4250 0.04025
R36553 VDD.n4252 VDD.n4251 0.04025
R36554 VDD.n4252 VDD.n2537 0.04025
R36555 VDD.n4256 VDD.n2537 0.04025
R36556 VDD.n4257 VDD.n4256 0.04025
R36557 VDD.n4258 VDD.n4257 0.04025
R36558 VDD.n4258 VDD.n2535 0.04025
R36559 VDD.n4262 VDD.n2535 0.04025
R36560 VDD.n4263 VDD.n4262 0.04025
R36561 VDD.n4264 VDD.n4263 0.04025
R36562 VDD.n4264 VDD.n2533 0.04025
R36563 VDD.n4268 VDD.n2533 0.04025
R36564 VDD.n4269 VDD.n4268 0.04025
R36565 VDD.n4270 VDD.n4269 0.04025
R36566 VDD.n4270 VDD.n2531 0.04025
R36567 VDD.n4274 VDD.n2531 0.04025
R36568 VDD.n4275 VDD.n4274 0.04025
R36569 VDD.n4276 VDD.n4275 0.04025
R36570 VDD.n4276 VDD.n2529 0.04025
R36571 VDD.n4280 VDD.n2529 0.04025
R36572 VDD.n4281 VDD.n4280 0.04025
R36573 VDD.n4282 VDD.n4281 0.04025
R36574 VDD.n4282 VDD.n2527 0.04025
R36575 VDD.n4286 VDD.n2527 0.04025
R36576 VDD.n4287 VDD.n4286 0.04025
R36577 VDD.n4288 VDD.n4287 0.04025
R36578 VDD.n4288 VDD.n2525 0.04025
R36579 VDD.n4292 VDD.n2525 0.04025
R36580 VDD.n4293 VDD.n4292 0.04025
R36581 VDD.n4294 VDD.n4293 0.04025
R36582 VDD.n4294 VDD.n2523 0.04025
R36583 VDD.n4298 VDD.n2523 0.04025
R36584 VDD.n4299 VDD.n4298 0.04025
R36585 VDD.n4300 VDD.n4299 0.04025
R36586 VDD.n4300 VDD.n2521 0.04025
R36587 VDD.n4304 VDD.n2521 0.04025
R36588 VDD.n4305 VDD.n4304 0.04025
R36589 VDD.n4306 VDD.n4305 0.04025
R36590 VDD.n4306 VDD.n2519 0.04025
R36591 VDD.n4310 VDD.n2519 0.04025
R36592 VDD.n4311 VDD.n4310 0.04025
R36593 VDD.n4312 VDD.n4311 0.04025
R36594 VDD.n4312 VDD.n2517 0.04025
R36595 VDD.n4316 VDD.n2517 0.04025
R36596 VDD.n4317 VDD.n4316 0.04025
R36597 VDD.n4318 VDD.n4317 0.04025
R36598 VDD.n4318 VDD.n2515 0.04025
R36599 VDD.n4322 VDD.n2515 0.04025
R36600 VDD.n4323 VDD.n4322 0.04025
R36601 VDD.n4324 VDD.n4323 0.04025
R36602 VDD.n4324 VDD.n2513 0.04025
R36603 VDD.n4328 VDD.n2513 0.04025
R36604 VDD.n4329 VDD.n4328 0.04025
R36605 VDD.n4330 VDD.n4329 0.04025
R36606 VDD.n4330 VDD.n2511 0.04025
R36607 VDD.n4334 VDD.n2511 0.04025
R36608 VDD.n4335 VDD.n4334 0.04025
R36609 VDD.n4336 VDD.n4335 0.04025
R36610 VDD.n4336 VDD.n2509 0.04025
R36611 VDD.n4340 VDD.n2509 0.04025
R36612 VDD.n4341 VDD.n4340 0.04025
R36613 VDD.n4342 VDD.n4341 0.04025
R36614 VDD.n4342 VDD.n2507 0.04025
R36615 VDD.n4346 VDD.n2507 0.04025
R36616 VDD.n4347 VDD.n4346 0.04025
R36617 VDD.n4348 VDD.n4347 0.04025
R36618 VDD.n4348 VDD.n2505 0.04025
R36619 VDD.n4352 VDD.n2505 0.04025
R36620 VDD.n4353 VDD.n4352 0.04025
R36621 VDD.n4354 VDD.n4353 0.04025
R36622 VDD.n4354 VDD.n2503 0.04025
R36623 VDD.n4358 VDD.n2503 0.04025
R36624 VDD.n4359 VDD.n4358 0.04025
R36625 VDD.n4360 VDD.n4359 0.04025
R36626 VDD.n4360 VDD.n2501 0.04025
R36627 VDD.n4364 VDD.n2501 0.04025
R36628 VDD.n4365 VDD.n4364 0.04025
R36629 VDD.n4366 VDD.n4365 0.04025
R36630 VDD.n4366 VDD.n2499 0.04025
R36631 VDD.n4370 VDD.n2499 0.04025
R36632 VDD.n4371 VDD.n4370 0.04025
R36633 VDD.n4372 VDD.n4371 0.04025
R36634 VDD.n4372 VDD.n2497 0.04025
R36635 VDD.n4376 VDD.n2497 0.04025
R36636 VDD.n4377 VDD.n4376 0.04025
R36637 VDD.n4378 VDD.n4377 0.04025
R36638 VDD.n4378 VDD.n2495 0.04025
R36639 VDD.n4382 VDD.n2495 0.04025
R36640 VDD.n4383 VDD.n4382 0.04025
R36641 VDD.n4384 VDD.n4383 0.04025
R36642 VDD.n4384 VDD.n2493 0.04025
R36643 VDD.n4388 VDD.n2493 0.04025
R36644 VDD.n4389 VDD.n4388 0.04025
R36645 VDD.n4390 VDD.n4389 0.04025
R36646 VDD.n4390 VDD.n2491 0.04025
R36647 VDD.n4394 VDD.n2491 0.04025
R36648 VDD.n4395 VDD.n4394 0.04025
R36649 VDD.n4396 VDD.n4395 0.04025
R36650 VDD.n4396 VDD.n2489 0.04025
R36651 VDD.n4400 VDD.n2489 0.04025
R36652 VDD.n4401 VDD.n4400 0.04025
R36653 VDD.n4402 VDD.n4401 0.04025
R36654 VDD.n4402 VDD.n2487 0.04025
R36655 VDD.n4406 VDD.n2487 0.04025
R36656 VDD.n4407 VDD.n4406 0.04025
R36657 VDD.n4408 VDD.n4407 0.04025
R36658 VDD.n4408 VDD.n2485 0.04025
R36659 VDD.n4412 VDD.n2485 0.04025
R36660 VDD.n4413 VDD.n4412 0.04025
R36661 VDD.n4414 VDD.n4413 0.04025
R36662 VDD.n4414 VDD.n2483 0.04025
R36663 VDD.n4418 VDD.n2483 0.04025
R36664 VDD.n4419 VDD.n4418 0.04025
R36665 VDD.n4420 VDD.n4419 0.04025
R36666 VDD.n4420 VDD.n2481 0.04025
R36667 VDD.n4424 VDD.n2481 0.04025
R36668 VDD.n4425 VDD.n4424 0.04025
R36669 VDD.n4426 VDD.n4425 0.04025
R36670 VDD.n4426 VDD.n2479 0.04025
R36671 VDD.n4430 VDD.n2479 0.04025
R36672 VDD.n4431 VDD.n4430 0.04025
R36673 VDD.n4432 VDD.n4431 0.04025
R36674 VDD.n4432 VDD.n2477 0.04025
R36675 VDD.n4436 VDD.n2477 0.04025
R36676 VDD.n4437 VDD.n4436 0.04025
R36677 VDD.n4438 VDD.n4437 0.04025
R36678 VDD.n4438 VDD.n2475 0.04025
R36679 VDD.n4442 VDD.n2475 0.04025
R36680 VDD.n4443 VDD.n4442 0.04025
R36681 VDD.n4444 VDD.n4443 0.04025
R36682 VDD.n4444 VDD.n2473 0.04025
R36683 VDD.n4448 VDD.n2473 0.04025
R36684 VDD.n4449 VDD.n4448 0.04025
R36685 VDD.n4450 VDD.n4449 0.04025
R36686 VDD.n4450 VDD.n2471 0.04025
R36687 VDD.n4454 VDD.n2471 0.04025
R36688 VDD.n4455 VDD.n4454 0.04025
R36689 VDD.n4456 VDD.n4455 0.04025
R36690 VDD.n4456 VDD.n2469 0.04025
R36691 VDD.n4460 VDD.n2469 0.04025
R36692 VDD.n4461 VDD.n4460 0.04025
R36693 VDD.n4462 VDD.n4461 0.04025
R36694 VDD.n4462 VDD.n2467 0.04025
R36695 VDD.n4466 VDD.n2467 0.04025
R36696 VDD.n4467 VDD.n4466 0.04025
R36697 VDD.n4468 VDD.n4467 0.04025
R36698 VDD.n4468 VDD.n2465 0.04025
R36699 VDD.n4472 VDD.n2465 0.04025
R36700 VDD.n4473 VDD.n4472 0.04025
R36701 VDD.n4474 VDD.n4473 0.04025
R36702 VDD.n4474 VDD.n2463 0.04025
R36703 VDD.n4478 VDD.n2463 0.04025
R36704 VDD.n4479 VDD.n4478 0.04025
R36705 VDD.n4480 VDD.n4479 0.04025
R36706 VDD.n4480 VDD.n2461 0.04025
R36707 VDD.n4484 VDD.n2461 0.04025
R36708 VDD.n4485 VDD.n4484 0.04025
R36709 VDD.n4486 VDD.n4485 0.04025
R36710 VDD.n4486 VDD.n2459 0.04025
R36711 VDD.n4490 VDD.n2459 0.04025
R36712 VDD.n4491 VDD.n4490 0.04025
R36713 VDD.n4492 VDD.n4491 0.04025
R36714 VDD.n4492 VDD.n2457 0.04025
R36715 VDD.n4496 VDD.n2457 0.04025
R36716 VDD.n4497 VDD.n4496 0.04025
R36717 VDD.n4498 VDD.n4497 0.04025
R36718 VDD.n4498 VDD.n2455 0.04025
R36719 VDD.n4502 VDD.n2455 0.04025
R36720 VDD.n4503 VDD.n4502 0.04025
R36721 VDD.n4504 VDD.n4503 0.04025
R36722 VDD.n4504 VDD.n2453 0.04025
R36723 VDD.n4508 VDD.n2453 0.04025
R36724 VDD.n4509 VDD.n4508 0.04025
R36725 VDD.n4510 VDD.n4509 0.04025
R36726 VDD.n4510 VDD.n2451 0.04025
R36727 VDD.n4514 VDD.n2451 0.04025
R36728 VDD.n4515 VDD.n4514 0.04025
R36729 VDD.n4516 VDD.n4515 0.04025
R36730 VDD.n4516 VDD.n2449 0.04025
R36731 VDD.n4520 VDD.n2449 0.04025
R36732 VDD.n4521 VDD.n4520 0.04025
R36733 VDD.n4522 VDD.n4521 0.04025
R36734 VDD.n4522 VDD.n2447 0.04025
R36735 VDD.n4526 VDD.n2447 0.04025
R36736 VDD.n4527 VDD.n4526 0.04025
R36737 VDD.n4528 VDD.n4527 0.04025
R36738 VDD.n4528 VDD.n2445 0.04025
R36739 VDD.n4532 VDD.n2445 0.04025
R36740 VDD.n4533 VDD.n4532 0.04025
R36741 VDD.n4534 VDD.n4533 0.04025
R36742 VDD.n4534 VDD.n2443 0.04025
R36743 VDD.n4538 VDD.n2443 0.04025
R36744 VDD.n4539 VDD.n4538 0.04025
R36745 VDD.n4540 VDD.n4539 0.04025
R36746 VDD.n4540 VDD.n2441 0.04025
R36747 VDD.n4544 VDD.n2441 0.04025
R36748 VDD.n4545 VDD.n4544 0.04025
R36749 VDD.n4546 VDD.n4545 0.04025
R36750 VDD.n4546 VDD.n2439 0.04025
R36751 VDD.n4550 VDD.n2439 0.04025
R36752 VDD.n4551 VDD.n4550 0.04025
R36753 VDD.n4552 VDD.n4551 0.04025
R36754 VDD.n4552 VDD.n2437 0.04025
R36755 VDD.n4556 VDD.n2437 0.04025
R36756 VDD.n4557 VDD.n4556 0.04025
R36757 VDD.n4558 VDD.n4557 0.04025
R36758 VDD.n4558 VDD.n2435 0.04025
R36759 VDD.n4562 VDD.n2435 0.04025
R36760 VDD.n4563 VDD.n4562 0.04025
R36761 VDD.n4564 VDD.n4563 0.04025
R36762 VDD.n4564 VDD.n2433 0.04025
R36763 VDD.n4568 VDD.n2433 0.04025
R36764 VDD.n4569 VDD.n4568 0.04025
R36765 VDD.n4570 VDD.n4569 0.04025
R36766 VDD.n4570 VDD.n2431 0.04025
R36767 VDD.n4574 VDD.n2431 0.04025
R36768 VDD.n4575 VDD.n4574 0.04025
R36769 VDD.n4576 VDD.n4575 0.04025
R36770 VDD.n4576 VDD.n2429 0.04025
R36771 VDD.n4580 VDD.n2429 0.04025
R36772 VDD.n4581 VDD.n4580 0.04025
R36773 VDD.n4582 VDD.n4581 0.04025
R36774 VDD.n4582 VDD.n2427 0.04025
R36775 VDD.n4586 VDD.n2427 0.04025
R36776 VDD.n4587 VDD.n4586 0.04025
R36777 VDD.n4588 VDD.n4587 0.04025
R36778 VDD.n4588 VDD.n2425 0.04025
R36779 VDD.n4593 VDD.n4592 0.04025
R36780 VDD.n4595 VDD.n4594 0.04025
R36781 VDD.n5219 VDD.n4595 0.04025
R36782 VDD.n5219 VDD.n5204 0.04025
R36783 VDD.n5199 VDD.n4599 0.04025
R36784 VDD.n5199 VDD.n5198 0.04025
R36785 VDD.n5198 VDD.n5197 0.04025
R36786 VDD.n5197 VDD.n4600 0.04025
R36787 VDD.n5193 VDD.n4600 0.04025
R36788 VDD.n5193 VDD.n5192 0.04025
R36789 VDD.n5192 VDD.n5191 0.04025
R36790 VDD.n5191 VDD.n4602 0.04025
R36791 VDD.n5187 VDD.n4602 0.04025
R36792 VDD.n5187 VDD.n5186 0.04025
R36793 VDD.n5186 VDD.n5185 0.04025
R36794 VDD.n5185 VDD.n4604 0.04025
R36795 VDD.n5181 VDD.n4604 0.04025
R36796 VDD.n5181 VDD.n5180 0.04025
R36797 VDD.n5180 VDD.n5179 0.04025
R36798 VDD.n5179 VDD.n4606 0.04025
R36799 VDD.n5175 VDD.n4606 0.04025
R36800 VDD.n5175 VDD.n5174 0.04025
R36801 VDD.n5174 VDD.n5173 0.04025
R36802 VDD.n5173 VDD.n4608 0.04025
R36803 VDD.n5169 VDD.n4608 0.04025
R36804 VDD.n5169 VDD.n5168 0.04025
R36805 VDD.n5168 VDD.n5167 0.04025
R36806 VDD.n5167 VDD.n4610 0.04025
R36807 VDD.n5163 VDD.n4610 0.04025
R36808 VDD.n5163 VDD.n5162 0.04025
R36809 VDD.n5162 VDD.n5161 0.04025
R36810 VDD.n5161 VDD.n4612 0.04025
R36811 VDD.n5157 VDD.n4612 0.04025
R36812 VDD.n5157 VDD.n5156 0.04025
R36813 VDD.n5156 VDD.n5155 0.04025
R36814 VDD.n5155 VDD.n4614 0.04025
R36815 VDD.n5151 VDD.n4614 0.04025
R36816 VDD.n5151 VDD.n5150 0.04025
R36817 VDD.n5150 VDD.n5149 0.04025
R36818 VDD.n5149 VDD.n4616 0.04025
R36819 VDD.n5145 VDD.n4616 0.04025
R36820 VDD.n5145 VDD.n5144 0.04025
R36821 VDD.n5144 VDD.n5143 0.04025
R36822 VDD.n5143 VDD.n4618 0.04025
R36823 VDD.n5139 VDD.n4618 0.04025
R36824 VDD.n5139 VDD.n5138 0.04025
R36825 VDD.n5138 VDD.n5137 0.04025
R36826 VDD.n5137 VDD.n4620 0.04025
R36827 VDD.n5133 VDD.n4620 0.04025
R36828 VDD.n5133 VDD.n5132 0.04025
R36829 VDD.n5132 VDD.n5131 0.04025
R36830 VDD.n5131 VDD.n4622 0.04025
R36831 VDD.n5127 VDD.n4622 0.04025
R36832 VDD.n5127 VDD.n5126 0.04025
R36833 VDD.n5126 VDD.n5125 0.04025
R36834 VDD.n5125 VDD.n4624 0.04025
R36835 VDD.n5121 VDD.n4624 0.04025
R36836 VDD.n5121 VDD.n5120 0.04025
R36837 VDD.n5120 VDD.n5119 0.04025
R36838 VDD.n5119 VDD.n4626 0.04025
R36839 VDD.n5115 VDD.n4626 0.04025
R36840 VDD.n5115 VDD.n5114 0.04025
R36841 VDD.n5114 VDD.n5113 0.04025
R36842 VDD.n5113 VDD.n4628 0.04025
R36843 VDD.n5109 VDD.n4628 0.04025
R36844 VDD.n5109 VDD.n5108 0.04025
R36845 VDD.n5108 VDD.n5107 0.04025
R36846 VDD.n5107 VDD.n4630 0.04025
R36847 VDD.n5103 VDD.n4630 0.04025
R36848 VDD.n5103 VDD.n5102 0.04025
R36849 VDD.n5102 VDD.n5101 0.04025
R36850 VDD.n5101 VDD.n4632 0.04025
R36851 VDD.n5097 VDD.n4632 0.04025
R36852 VDD.n5097 VDD.n5096 0.04025
R36853 VDD.n5096 VDD.n5095 0.04025
R36854 VDD.n5095 VDD.n4634 0.04025
R36855 VDD.n5091 VDD.n4634 0.04025
R36856 VDD.n5091 VDD.n5090 0.04025
R36857 VDD.n5090 VDD.n5089 0.04025
R36858 VDD.n5089 VDD.n4636 0.04025
R36859 VDD.n5085 VDD.n4636 0.04025
R36860 VDD.n5085 VDD.n5084 0.04025
R36861 VDD.n5084 VDD.n5083 0.04025
R36862 VDD.n5083 VDD.n4638 0.04025
R36863 VDD.n5079 VDD.n4638 0.04025
R36864 VDD.n5079 VDD.n5078 0.04025
R36865 VDD.n5078 VDD.n5077 0.04025
R36866 VDD.n5077 VDD.n4640 0.04025
R36867 VDD.n5073 VDD.n4640 0.04025
R36868 VDD.n5073 VDD.n5072 0.04025
R36869 VDD.n5072 VDD.n5071 0.04025
R36870 VDD.n5071 VDD.n4642 0.04025
R36871 VDD.n5067 VDD.n4642 0.04025
R36872 VDD.n5067 VDD.n5066 0.04025
R36873 VDD.n5066 VDD.n5065 0.04025
R36874 VDD.n5065 VDD.n4644 0.04025
R36875 VDD.n5061 VDD.n4644 0.04025
R36876 VDD.n5061 VDD.n5060 0.04025
R36877 VDD.n5060 VDD.n5059 0.04025
R36878 VDD.n5059 VDD.n4646 0.04025
R36879 VDD.n5055 VDD.n4646 0.04025
R36880 VDD.n5055 VDD.n5054 0.04025
R36881 VDD.n5054 VDD.n5053 0.04025
R36882 VDD.n5053 VDD.n4648 0.04025
R36883 VDD.n5049 VDD.n4648 0.04025
R36884 VDD.n5049 VDD.n5048 0.04025
R36885 VDD.n5048 VDD.n5047 0.04025
R36886 VDD.n5047 VDD.n4650 0.04025
R36887 VDD.n5043 VDD.n4650 0.04025
R36888 VDD.n5043 VDD.n5042 0.04025
R36889 VDD.n5042 VDD.n5041 0.04025
R36890 VDD.n5041 VDD.n4652 0.04025
R36891 VDD.n5037 VDD.n4652 0.04025
R36892 VDD.n5037 VDD.n5036 0.04025
R36893 VDD.n5036 VDD.n5035 0.04025
R36894 VDD.n5035 VDD.n4654 0.04025
R36895 VDD.n5031 VDD.n4654 0.04025
R36896 VDD.n5031 VDD.n5030 0.04025
R36897 VDD.n5030 VDD.n5029 0.04025
R36898 VDD.n5029 VDD.n4656 0.04025
R36899 VDD.n5025 VDD.n4656 0.04025
R36900 VDD.n5025 VDD.n5024 0.04025
R36901 VDD.n5024 VDD.n5023 0.04025
R36902 VDD.n5023 VDD.n4658 0.04025
R36903 VDD.n5019 VDD.n4658 0.04025
R36904 VDD.n5019 VDD.n5018 0.04025
R36905 VDD.n5018 VDD.n5017 0.04025
R36906 VDD.n5017 VDD.n4660 0.04025
R36907 VDD.n5013 VDD.n4660 0.04025
R36908 VDD.n5013 VDD.n5012 0.04025
R36909 VDD.n5012 VDD.n5011 0.04025
R36910 VDD.n5011 VDD.n4662 0.04025
R36911 VDD.n5007 VDD.n4662 0.04025
R36912 VDD.n5007 VDD.n5006 0.04025
R36913 VDD.n5006 VDD.n5005 0.04025
R36914 VDD.n5005 VDD.n4664 0.04025
R36915 VDD.n5001 VDD.n4664 0.04025
R36916 VDD.n5001 VDD.n5000 0.04025
R36917 VDD.n5000 VDD.n4999 0.04025
R36918 VDD.n4999 VDD.n4666 0.04025
R36919 VDD.n4995 VDD.n4666 0.04025
R36920 VDD.n4995 VDD.n4994 0.04025
R36921 VDD.n4994 VDD.n4993 0.04025
R36922 VDD.n4993 VDD.n4668 0.04025
R36923 VDD.n4989 VDD.n4668 0.04025
R36924 VDD.n4989 VDD.n4988 0.04025
R36925 VDD.n4988 VDD.n4987 0.04025
R36926 VDD.n4987 VDD.n4670 0.04025
R36927 VDD.n4983 VDD.n4670 0.04025
R36928 VDD.n4983 VDD.n4982 0.04025
R36929 VDD.n4982 VDD.n4981 0.04025
R36930 VDD.n4981 VDD.n4672 0.04025
R36931 VDD.n4977 VDD.n4672 0.04025
R36932 VDD.n4977 VDD.n4976 0.04025
R36933 VDD.n4976 VDD.n4975 0.04025
R36934 VDD.n4975 VDD.n4674 0.04025
R36935 VDD.n4971 VDD.n4674 0.04025
R36936 VDD.n4971 VDD.n4970 0.04025
R36937 VDD.n4970 VDD.n4969 0.04025
R36938 VDD.n4969 VDD.n4676 0.04025
R36939 VDD.n4965 VDD.n4676 0.04025
R36940 VDD.n4965 VDD.n4964 0.04025
R36941 VDD.n4964 VDD.n4963 0.04025
R36942 VDD.n4963 VDD.n4678 0.04025
R36943 VDD.n4959 VDD.n4678 0.04025
R36944 VDD.n4959 VDD.n4958 0.04025
R36945 VDD.n4958 VDD.n4957 0.04025
R36946 VDD.n4957 VDD.n4680 0.04025
R36947 VDD.n4953 VDD.n4680 0.04025
R36948 VDD.n4953 VDD.n4952 0.04025
R36949 VDD.n4952 VDD.n4951 0.04025
R36950 VDD.n4951 VDD.n4682 0.04025
R36951 VDD.n4947 VDD.n4682 0.04025
R36952 VDD.n4947 VDD.n4946 0.04025
R36953 VDD.n4946 VDD.n4945 0.04025
R36954 VDD.n4945 VDD.n4684 0.04025
R36955 VDD.n4941 VDD.n4684 0.04025
R36956 VDD.n4941 VDD.n4940 0.04025
R36957 VDD.n4940 VDD.n4939 0.04025
R36958 VDD.n4939 VDD.n4686 0.04025
R36959 VDD.n4935 VDD.n4686 0.04025
R36960 VDD.n4935 VDD.n4934 0.04025
R36961 VDD.n4934 VDD.n4933 0.04025
R36962 VDD.n4933 VDD.n4688 0.04025
R36963 VDD.n4929 VDD.n4688 0.04025
R36964 VDD.n4929 VDD.n4928 0.04025
R36965 VDD.n4928 VDD.n4927 0.04025
R36966 VDD.n4927 VDD.n4690 0.04025
R36967 VDD.n4923 VDD.n4690 0.04025
R36968 VDD.n4923 VDD.n4922 0.04025
R36969 VDD.n4922 VDD.n4921 0.04025
R36970 VDD.n4921 VDD.n4692 0.04025
R36971 VDD.n4917 VDD.n4692 0.04025
R36972 VDD.n4917 VDD.n4916 0.04025
R36973 VDD.n4916 VDD.n4915 0.04025
R36974 VDD.n4915 VDD.n4694 0.04025
R36975 VDD.n4911 VDD.n4694 0.04025
R36976 VDD.n4911 VDD.n4910 0.04025
R36977 VDD.n4910 VDD.n4909 0.04025
R36978 VDD.n4909 VDD.n4696 0.04025
R36979 VDD.n4905 VDD.n4696 0.04025
R36980 VDD.n3628 VDD.n3627 0.04025
R36981 VDD.n3627 VDD.n3626 0.04025
R36982 VDD.n3626 VDD.n2747 0.04025
R36983 VDD.n3622 VDD.n2747 0.04025
R36984 VDD.n3622 VDD.n3621 0.04025
R36985 VDD.n3621 VDD.n3620 0.04025
R36986 VDD.n3620 VDD.n2749 0.04025
R36987 VDD.n3616 VDD.n2749 0.04025
R36988 VDD.n3616 VDD.n3615 0.04025
R36989 VDD.n3615 VDD.n3614 0.04025
R36990 VDD.n3614 VDD.n2751 0.04025
R36991 VDD.n3610 VDD.n2751 0.04025
R36992 VDD.n3610 VDD.n3609 0.04025
R36993 VDD.n3609 VDD.n3608 0.04025
R36994 VDD.n3608 VDD.n2753 0.04025
R36995 VDD.n3604 VDD.n2753 0.04025
R36996 VDD.n3604 VDD.n3603 0.04025
R36997 VDD.n3603 VDD.n3602 0.04025
R36998 VDD.n3602 VDD.n2755 0.04025
R36999 VDD.n3598 VDD.n2755 0.04025
R37000 VDD.n3598 VDD.n3597 0.04025
R37001 VDD.n3597 VDD.n3596 0.04025
R37002 VDD.n3596 VDD.n2757 0.04025
R37003 VDD.n3592 VDD.n2757 0.04025
R37004 VDD.n3592 VDD.n3591 0.04025
R37005 VDD.n3591 VDD.n3590 0.04025
R37006 VDD.n3590 VDD.n2759 0.04025
R37007 VDD.n3586 VDD.n2759 0.04025
R37008 VDD.n3586 VDD.n3585 0.04025
R37009 VDD.n3585 VDD.n3584 0.04025
R37010 VDD.n3584 VDD.n2761 0.04025
R37011 VDD.n3580 VDD.n2761 0.04025
R37012 VDD.n3580 VDD.n3579 0.04025
R37013 VDD.n3579 VDD.n3578 0.04025
R37014 VDD.n3578 VDD.n2763 0.04025
R37015 VDD.n3574 VDD.n2763 0.04025
R37016 VDD.n3574 VDD.n3573 0.04025
R37017 VDD.n3573 VDD.n3572 0.04025
R37018 VDD.n3572 VDD.n2765 0.04025
R37019 VDD.n3568 VDD.n2765 0.04025
R37020 VDD.n3568 VDD.n3567 0.04025
R37021 VDD.n3567 VDD.n3566 0.04025
R37022 VDD.n3566 VDD.n2767 0.04025
R37023 VDD.n3562 VDD.n2767 0.04025
R37024 VDD.n3562 VDD.n3561 0.04025
R37025 VDD.n3561 VDD.n3560 0.04025
R37026 VDD.n3560 VDD.n2769 0.04025
R37027 VDD.n3556 VDD.n2769 0.04025
R37028 VDD.n3556 VDD.n3555 0.04025
R37029 VDD.n3555 VDD.n3554 0.04025
R37030 VDD.n3554 VDD.n2771 0.04025
R37031 VDD.n3550 VDD.n2771 0.04025
R37032 VDD.n3550 VDD.n3549 0.04025
R37033 VDD.n3549 VDD.n3548 0.04025
R37034 VDD.n3548 VDD.n2773 0.04025
R37035 VDD.n3544 VDD.n2773 0.04025
R37036 VDD.n3544 VDD.n3543 0.04025
R37037 VDD.n3543 VDD.n3542 0.04025
R37038 VDD.n3542 VDD.n2775 0.04025
R37039 VDD.n3538 VDD.n2775 0.04025
R37040 VDD.n3538 VDD.n3537 0.04025
R37041 VDD.n3537 VDD.n3536 0.04025
R37042 VDD.n3536 VDD.n2777 0.04025
R37043 VDD.n3532 VDD.n2777 0.04025
R37044 VDD.n3532 VDD.n3531 0.04025
R37045 VDD.n3531 VDD.n3530 0.04025
R37046 VDD.n3530 VDD.n2779 0.04025
R37047 VDD.n3526 VDD.n2779 0.04025
R37048 VDD.n3526 VDD.n3525 0.04025
R37049 VDD.n3525 VDD.n3524 0.04025
R37050 VDD.n3524 VDD.n2781 0.04025
R37051 VDD.n3520 VDD.n2781 0.04025
R37052 VDD.n3520 VDD.n3519 0.04025
R37053 VDD.n3519 VDD.n3518 0.04025
R37054 VDD.n3518 VDD.n2783 0.04025
R37055 VDD.n3514 VDD.n2783 0.04025
R37056 VDD.n3514 VDD.n3513 0.04025
R37057 VDD.n3513 VDD.n3512 0.04025
R37058 VDD.n3512 VDD.n2785 0.04025
R37059 VDD.n3508 VDD.n2785 0.04025
R37060 VDD.n3508 VDD.n3507 0.04025
R37061 VDD.n3507 VDD.n3506 0.04025
R37062 VDD.n3506 VDD.n2787 0.04025
R37063 VDD.n3502 VDD.n2787 0.04025
R37064 VDD.n3502 VDD.n3501 0.04025
R37065 VDD.n3501 VDD.n3500 0.04025
R37066 VDD.n3500 VDD.n2789 0.04025
R37067 VDD.n3496 VDD.n2789 0.04025
R37068 VDD.n3496 VDD.n3495 0.04025
R37069 VDD.n3495 VDD.n3494 0.04025
R37070 VDD.n3494 VDD.n2791 0.04025
R37071 VDD.n3490 VDD.n2791 0.04025
R37072 VDD.n3490 VDD.n3489 0.04025
R37073 VDD.n3489 VDD.n3488 0.04025
R37074 VDD.n3488 VDD.n2793 0.04025
R37075 VDD.n3484 VDD.n2793 0.04025
R37076 VDD.n3484 VDD.n3483 0.04025
R37077 VDD.n3483 VDD.n3482 0.04025
R37078 VDD.n3482 VDD.n2795 0.04025
R37079 VDD.n3478 VDD.n2795 0.04025
R37080 VDD.n3478 VDD.n3477 0.04025
R37081 VDD.n3477 VDD.n3476 0.04025
R37082 VDD.n3476 VDD.n2797 0.04025
R37083 VDD.n3472 VDD.n2797 0.04025
R37084 VDD.n3472 VDD.n3471 0.04025
R37085 VDD.n3471 VDD.n3470 0.04025
R37086 VDD.n3470 VDD.n2799 0.04025
R37087 VDD.n3466 VDD.n2799 0.04025
R37088 VDD.n3466 VDD.n3465 0.04025
R37089 VDD.n3465 VDD.n3464 0.04025
R37090 VDD.n3464 VDD.n2801 0.04025
R37091 VDD.n3460 VDD.n2801 0.04025
R37092 VDD.n3460 VDD.n3459 0.04025
R37093 VDD.n3459 VDD.n3458 0.04025
R37094 VDD.n3458 VDD.n2803 0.04025
R37095 VDD.n3454 VDD.n2803 0.04025
R37096 VDD.n3454 VDD.n3453 0.04025
R37097 VDD.n3453 VDD.n3452 0.04025
R37098 VDD.n3452 VDD.n2805 0.04025
R37099 VDD.n3448 VDD.n2805 0.04025
R37100 VDD.n3448 VDD.n3447 0.04025
R37101 VDD.n3447 VDD.n3446 0.04025
R37102 VDD.n3446 VDD.n2807 0.04025
R37103 VDD.n3442 VDD.n2807 0.04025
R37104 VDD.n3442 VDD.n3441 0.04025
R37105 VDD.n3441 VDD.n3440 0.04025
R37106 VDD.n3440 VDD.n2809 0.04025
R37107 VDD.n3436 VDD.n2809 0.04025
R37108 VDD.n3436 VDD.n3435 0.04025
R37109 VDD.n3435 VDD.n3434 0.04025
R37110 VDD.n3434 VDD.n2811 0.04025
R37111 VDD.n3430 VDD.n2811 0.04025
R37112 VDD.n3430 VDD.n3429 0.04025
R37113 VDD.n3429 VDD.n3428 0.04025
R37114 VDD.n3428 VDD.n2813 0.04025
R37115 VDD.n3424 VDD.n2813 0.04025
R37116 VDD.n3424 VDD.n3423 0.04025
R37117 VDD.n3423 VDD.n3422 0.04025
R37118 VDD.n3422 VDD.n2815 0.04025
R37119 VDD.n3418 VDD.n2815 0.04025
R37120 VDD.n3418 VDD.n3417 0.04025
R37121 VDD.n3417 VDD.n3416 0.04025
R37122 VDD.n3416 VDD.n2817 0.04025
R37123 VDD.n3412 VDD.n2817 0.04025
R37124 VDD.n3412 VDD.n3411 0.04025
R37125 VDD.n3411 VDD.n3410 0.04025
R37126 VDD.n3410 VDD.n2819 0.04025
R37127 VDD.n3406 VDD.n2819 0.04025
R37128 VDD.n3406 VDD.n3405 0.04025
R37129 VDD.n3405 VDD.n3404 0.04025
R37130 VDD.n3404 VDD.n2821 0.04025
R37131 VDD.n3400 VDD.n2821 0.04025
R37132 VDD.n3400 VDD.n3399 0.04025
R37133 VDD.n3399 VDD.n3398 0.04025
R37134 VDD.n3398 VDD.n2823 0.04025
R37135 VDD.n3394 VDD.n2823 0.04025
R37136 VDD.n3394 VDD.n3393 0.04025
R37137 VDD.n3393 VDD.n3392 0.04025
R37138 VDD.n3392 VDD.n2825 0.04025
R37139 VDD.n3388 VDD.n2825 0.04025
R37140 VDD.n3388 VDD.n3387 0.04025
R37141 VDD.n3387 VDD.n3386 0.04025
R37142 VDD.n3386 VDD.n2827 0.04025
R37143 VDD.n3382 VDD.n2827 0.04025
R37144 VDD.n3382 VDD.n3381 0.04025
R37145 VDD.n3381 VDD.n3380 0.04025
R37146 VDD.n3380 VDD.n2829 0.04025
R37147 VDD.n3376 VDD.n2829 0.04025
R37148 VDD.n3376 VDD.n3375 0.04025
R37149 VDD.n3375 VDD.n3374 0.04025
R37150 VDD.n3374 VDD.n2831 0.04025
R37151 VDD.n3370 VDD.n2831 0.04025
R37152 VDD.n3370 VDD.n3369 0.04025
R37153 VDD.n3369 VDD.n3368 0.04025
R37154 VDD.n3368 VDD.n2833 0.04025
R37155 VDD.n3364 VDD.n2833 0.04025
R37156 VDD.n3364 VDD.n3363 0.04025
R37157 VDD.n3363 VDD.n3362 0.04025
R37158 VDD.n3362 VDD.n2835 0.04025
R37159 VDD.n3358 VDD.n2835 0.04025
R37160 VDD.n3358 VDD.n3357 0.04025
R37161 VDD.n3357 VDD.n3356 0.04025
R37162 VDD.n3356 VDD.n2837 0.04025
R37163 VDD.n3352 VDD.n2837 0.04025
R37164 VDD.n3352 VDD.n3351 0.04025
R37165 VDD.n3351 VDD.n3350 0.04025
R37166 VDD.n3350 VDD.n2839 0.04025
R37167 VDD.n3346 VDD.n2839 0.04025
R37168 VDD.n3346 VDD.n3345 0.04025
R37169 VDD.n3345 VDD.n3344 0.04025
R37170 VDD.n3344 VDD.n2841 0.04025
R37171 VDD.n3340 VDD.n2841 0.04025
R37172 VDD.n3340 VDD.n3339 0.04025
R37173 VDD.n3339 VDD.n3338 0.04025
R37174 VDD.n3338 VDD.n2843 0.04025
R37175 VDD.n3334 VDD.n2843 0.04025
R37176 VDD.n3334 VDD.n3333 0.04025
R37177 VDD.n3333 VDD.n3332 0.04025
R37178 VDD.n3332 VDD.n2845 0.04025
R37179 VDD.n3328 VDD.n2845 0.04025
R37180 VDD.n3328 VDD.n3327 0.04025
R37181 VDD.n3327 VDD.n3326 0.04025
R37182 VDD.n3326 VDD.n2847 0.04025
R37183 VDD.n3322 VDD.n2847 0.04025
R37184 VDD.n3322 VDD.n3321 0.04025
R37185 VDD.n3321 VDD.n3320 0.04025
R37186 VDD.n3320 VDD.n2849 0.04025
R37187 VDD.n3316 VDD.n2849 0.04025
R37188 VDD.n3316 VDD.n3315 0.04025
R37189 VDD.n3315 VDD.n3314 0.04025
R37190 VDD.n3314 VDD.n2851 0.04025
R37191 VDD.n3310 VDD.n2851 0.04025
R37192 VDD.n3310 VDD.n3309 0.04025
R37193 VDD.n3309 VDD.n3308 0.04025
R37194 VDD.n3308 VDD.n2853 0.04025
R37195 VDD.n3304 VDD.n2853 0.04025
R37196 VDD.n3304 VDD.n3303 0.04025
R37197 VDD.n3303 VDD.n3302 0.04025
R37198 VDD.n3302 VDD.n2855 0.04025
R37199 VDD.n3298 VDD.n2855 0.04025
R37200 VDD.n3298 VDD.n3297 0.04025
R37201 VDD.n3297 VDD.n3296 0.04025
R37202 VDD.n3296 VDD.n2857 0.04025
R37203 VDD.n3292 VDD.n2857 0.04025
R37204 VDD.n3292 VDD.n3291 0.04025
R37205 VDD.n3291 VDD.n3290 0.04025
R37206 VDD.n3290 VDD.n2859 0.04025
R37207 VDD.n3286 VDD.n2859 0.04025
R37208 VDD.n3286 VDD.n3285 0.04025
R37209 VDD.n3285 VDD.n3284 0.04025
R37210 VDD.n3284 VDD.n2861 0.04025
R37211 VDD.n3280 VDD.n2861 0.04025
R37212 VDD.n3280 VDD.n3279 0.04025
R37213 VDD.n3279 VDD.n3278 0.04025
R37214 VDD.n3278 VDD.n2863 0.04025
R37215 VDD.n3274 VDD.n2863 0.04025
R37216 VDD.n3274 VDD.n3273 0.04025
R37217 VDD.n3273 VDD.n3272 0.04025
R37218 VDD.n3272 VDD.n2865 0.04025
R37219 VDD.n3268 VDD.n2865 0.04025
R37220 VDD.n3268 VDD.n3267 0.04025
R37221 VDD.n3267 VDD.n3266 0.04025
R37222 VDD.n3266 VDD.n2867 0.04025
R37223 VDD.n3262 VDD.n2867 0.04025
R37224 VDD.n3262 VDD.n3261 0.04025
R37225 VDD.n3261 VDD.n3260 0.04025
R37226 VDD.n3260 VDD.n2869 0.04025
R37227 VDD.n3256 VDD.n2869 0.04025
R37228 VDD.n3256 VDD.n3255 0.04025
R37229 VDD.n3255 VDD.n3254 0.04025
R37230 VDD.n3254 VDD.n2871 0.04025
R37231 VDD.n3250 VDD.n2871 0.04025
R37232 VDD.n3250 VDD.n3249 0.04025
R37233 VDD.n3249 VDD.n3248 0.04025
R37234 VDD.n3248 VDD.n2873 0.04025
R37235 VDD.n3244 VDD.n2873 0.04025
R37236 VDD.n3244 VDD.n3243 0.04025
R37237 VDD.n3243 VDD.n3242 0.04025
R37238 VDD.n3242 VDD.n2875 0.04025
R37239 VDD.n3238 VDD.n2875 0.04025
R37240 VDD.n3238 VDD.n3237 0.04025
R37241 VDD.n3237 VDD.n3236 0.04025
R37242 VDD.n3236 VDD.n2877 0.04025
R37243 VDD.n3232 VDD.n2877 0.04025
R37244 VDD.n3232 VDD.n3231 0.04025
R37245 VDD.n3231 VDD.n3230 0.04025
R37246 VDD.n3230 VDD.n2879 0.04025
R37247 VDD.n3226 VDD.n2879 0.04025
R37248 VDD.n3226 VDD.n3225 0.04025
R37249 VDD.n3225 VDD.n3224 0.04025
R37250 VDD.n3224 VDD.n2881 0.04025
R37251 VDD.n3220 VDD.n2881 0.04025
R37252 VDD.n3220 VDD.n3219 0.04025
R37253 VDD.n3219 VDD.n3218 0.04025
R37254 VDD.n3218 VDD.n2883 0.04025
R37255 VDD.n3214 VDD.n2883 0.04025
R37256 VDD.n3214 VDD.n3213 0.04025
R37257 VDD.n3213 VDD.n3212 0.04025
R37258 VDD.n3212 VDD.n2885 0.04025
R37259 VDD.n3208 VDD.n2885 0.04025
R37260 VDD.n3208 VDD.n3207 0.04025
R37261 VDD.n3207 VDD.n3206 0.04025
R37262 VDD.n3206 VDD.n2887 0.04025
R37263 VDD.n3202 VDD.n2887 0.04025
R37264 VDD.n3202 VDD.n3201 0.04025
R37265 VDD.n3201 VDD.n3200 0.04025
R37266 VDD.n3200 VDD.n2889 0.04025
R37267 VDD.n3196 VDD.n2889 0.04025
R37268 VDD.n3196 VDD.n3195 0.04025
R37269 VDD.n3195 VDD.n3194 0.04025
R37270 VDD.n3194 VDD.n2891 0.04025
R37271 VDD.n3190 VDD.n2891 0.04025
R37272 VDD.n3190 VDD.n3189 0.04025
R37273 VDD.n3189 VDD.n3188 0.04025
R37274 VDD.n3188 VDD.n2893 0.04025
R37275 VDD.n3184 VDD.n2893 0.04025
R37276 VDD.n3184 VDD.n3183 0.04025
R37277 VDD.n3183 VDD.n3182 0.04025
R37278 VDD.n3182 VDD.n2895 0.04025
R37279 VDD.n3178 VDD.n2895 0.04025
R37280 VDD.n3178 VDD.n3177 0.04025
R37281 VDD.n3177 VDD.n3176 0.04025
R37282 VDD.n3176 VDD.n2897 0.04025
R37283 VDD.n3172 VDD.n2897 0.04025
R37284 VDD.n3172 VDD.n3171 0.04025
R37285 VDD.n3171 VDD.n3170 0.04025
R37286 VDD.n3170 VDD.n2899 0.04025
R37287 VDD.n3166 VDD.n2899 0.04025
R37288 VDD.n3166 VDD.n3165 0.04025
R37289 VDD.n3165 VDD.n3164 0.04025
R37290 VDD.n3164 VDD.n2901 0.04025
R37291 VDD.n3160 VDD.n2901 0.04025
R37292 VDD.n3160 VDD.n3159 0.04025
R37293 VDD.n3159 VDD.n3158 0.04025
R37294 VDD.n3158 VDD.n2903 0.04025
R37295 VDD.n3154 VDD.n2903 0.04025
R37296 VDD.n3154 VDD.n3153 0.04025
R37297 VDD.n3153 VDD.n3152 0.04025
R37298 VDD.n3152 VDD.n2905 0.04025
R37299 VDD.n3148 VDD.n2905 0.04025
R37300 VDD.n3148 VDD.n3147 0.04025
R37301 VDD.n3147 VDD.n3146 0.04025
R37302 VDD.n3146 VDD.n2907 0.04025
R37303 VDD.n3142 VDD.n2907 0.04025
R37304 VDD.n3142 VDD.n3141 0.04025
R37305 VDD.n3141 VDD.n3140 0.04025
R37306 VDD.n3140 VDD.n2909 0.04025
R37307 VDD.n3136 VDD.n2909 0.04025
R37308 VDD.n3136 VDD.n3135 0.04025
R37309 VDD.n3135 VDD.n3134 0.04025
R37310 VDD.n3134 VDD.n2911 0.04025
R37311 VDD.n3130 VDD.n2911 0.04025
R37312 VDD.n3130 VDD.n3129 0.04025
R37313 VDD.n3129 VDD.n3128 0.04025
R37314 VDD.n3128 VDD.n2913 0.04025
R37315 VDD.n3124 VDD.n2913 0.04025
R37316 VDD.n3124 VDD.n3123 0.04025
R37317 VDD.n3123 VDD.n3122 0.04025
R37318 VDD.n3122 VDD.n2915 0.04025
R37319 VDD.n3118 VDD.n2915 0.04025
R37320 VDD.n3118 VDD.n3117 0.04025
R37321 VDD.n3117 VDD.n3116 0.04025
R37322 VDD.n3116 VDD.n2917 0.04025
R37323 VDD.n3112 VDD.n2917 0.04025
R37324 VDD.n3112 VDD.n3111 0.04025
R37325 VDD.n3111 VDD.n3110 0.04025
R37326 VDD.n3110 VDD.n2919 0.04025
R37327 VDD.n3106 VDD.n2919 0.04025
R37328 VDD.n3106 VDD.n3105 0.04025
R37329 VDD.n3105 VDD.n3104 0.04025
R37330 VDD.n3104 VDD.n2921 0.04025
R37331 VDD.n3100 VDD.n2921 0.04025
R37332 VDD.n3100 VDD.n3099 0.04025
R37333 VDD.n3099 VDD.n3098 0.04025
R37334 VDD.n3098 VDD.n2923 0.04025
R37335 VDD.n3094 VDD.n2923 0.04025
R37336 VDD.n3094 VDD.n3093 0.04025
R37337 VDD.n3093 VDD.n3092 0.04025
R37338 VDD.n3092 VDD.n2925 0.04025
R37339 VDD.n3088 VDD.n2925 0.04025
R37340 VDD.n3088 VDD.n3087 0.04025
R37341 VDD.n3087 VDD.n3086 0.04025
R37342 VDD.n3086 VDD.n2927 0.04025
R37343 VDD.n3082 VDD.n2927 0.04025
R37344 VDD.n3082 VDD.n3081 0.04025
R37345 VDD.n3081 VDD.n3080 0.04025
R37346 VDD.n3080 VDD.n2929 0.04025
R37347 VDD.n3076 VDD.n2929 0.04025
R37348 VDD.n3076 VDD.n3075 0.04025
R37349 VDD.n3075 VDD.n3074 0.04025
R37350 VDD.n3074 VDD.n2931 0.04025
R37351 VDD.n3070 VDD.n2931 0.04025
R37352 VDD.n3070 VDD.n3069 0.04025
R37353 VDD.n3069 VDD.n3068 0.04025
R37354 VDD.n3068 VDD.n2933 0.04025
R37355 VDD.n3064 VDD.n2933 0.04025
R37356 VDD.n3064 VDD.n3063 0.04025
R37357 VDD.n3063 VDD.n3062 0.04025
R37358 VDD.n3062 VDD.n2935 0.04025
R37359 VDD.n3058 VDD.n2935 0.04025
R37360 VDD.n3058 VDD.n3057 0.04025
R37361 VDD.n3057 VDD.n3056 0.04025
R37362 VDD.n3056 VDD.n2937 0.04025
R37363 VDD.n3052 VDD.n2937 0.04025
R37364 VDD.n3052 VDD.n3051 0.04025
R37365 VDD.n3051 VDD.n3050 0.04025
R37366 VDD.n3050 VDD.n2939 0.04025
R37367 VDD.n3046 VDD.n2939 0.04025
R37368 VDD.n3046 VDD.n3045 0.04025
R37369 VDD.n3045 VDD.n3044 0.04025
R37370 VDD.n3044 VDD.n2941 0.04025
R37371 VDD.n3040 VDD.n2941 0.04025
R37372 VDD.n3040 VDD.n3039 0.04025
R37373 VDD.n3039 VDD.n3038 0.04025
R37374 VDD.n3038 VDD.n2943 0.04025
R37375 VDD.n3034 VDD.n2943 0.04025
R37376 VDD.n3034 VDD.n3033 0.04025
R37377 VDD.n3033 VDD.n3032 0.04025
R37378 VDD.n3032 VDD.n2945 0.04025
R37379 VDD.n3028 VDD.n2945 0.04025
R37380 VDD.n3028 VDD.n3027 0.04025
R37381 VDD.n3027 VDD.n3026 0.04025
R37382 VDD.n3026 VDD.n2947 0.04025
R37383 VDD.n3022 VDD.n2947 0.04025
R37384 VDD.n3022 VDD.n3021 0.04025
R37385 VDD.n3021 VDD.n3020 0.04025
R37386 VDD.n3020 VDD.n2949 0.04025
R37387 VDD.n3016 VDD.n2949 0.04025
R37388 VDD.n3016 VDD.n3015 0.04025
R37389 VDD.n3015 VDD.n3014 0.04025
R37390 VDD.n3014 VDD.n2951 0.04025
R37391 VDD.n3010 VDD.n2951 0.04025
R37392 VDD.n3010 VDD.n3009 0.04025
R37393 VDD.n3009 VDD.n3008 0.04025
R37394 VDD.n3008 VDD.n2953 0.04025
R37395 VDD.n3004 VDD.n2953 0.04025
R37396 VDD.n3004 VDD.n3003 0.04025
R37397 VDD.n3003 VDD.n3002 0.04025
R37398 VDD.n3002 VDD.n2955 0.04025
R37399 VDD.n2998 VDD.n2955 0.04025
R37400 VDD.n2998 VDD.n2997 0.04025
R37401 VDD.n2997 VDD.n2996 0.04025
R37402 VDD.n2996 VDD.n2957 0.04025
R37403 VDD.n2992 VDD.n2957 0.04025
R37404 VDD.n2992 VDD.n2991 0.04025
R37405 VDD.n2991 VDD.n2990 0.04025
R37406 VDD.n2990 VDD.n2959 0.04025
R37407 VDD.n2986 VDD.n2959 0.04025
R37408 VDD.n2986 VDD.n2985 0.04025
R37409 VDD.n2985 VDD.n2984 0.04025
R37410 VDD.n2984 VDD.n2961 0.04025
R37411 VDD.n2980 VDD.n2961 0.04025
R37412 VDD.n2980 VDD.n2979 0.04025
R37413 VDD.n2979 VDD.n2978 0.04025
R37414 VDD.n2978 VDD.n2963 0.04025
R37415 VDD.n2974 VDD.n2963 0.04025
R37416 VDD.n2974 VDD.n2973 0.04025
R37417 VDD.n2973 VDD.n2972 0.04025
R37418 VDD.n2972 VDD.n2965 0.04025
R37419 VDD.n2968 VDD.n2965 0.04025
R37420 VDD.n2968 VDD.n2967 0.04025
R37421 VDD.n2967 VDD.n1767 0.04025
R37422 VDD.n11039 VDD.n1767 0.04025
R37423 VDD.n11042 VDD.n11039 0.04025
R37424 VDD.n11042 VDD.n11041 0.04025
R37425 VDD.n11041 VDD.n11040 0.04025
R37426 VDD.n11040 VDD.n668 0.04025
R37427 VDD.n11051 VDD.n668 0.04025
R37428 VDD.n11052 VDD.n11051 0.04025
R37429 VDD.n11053 VDD.n11052 0.04025
R37430 VDD.n11053 VDD.n666 0.04025
R37431 VDD.n11059 VDD.n666 0.04025
R37432 VDD.n11060 VDD.n11059 0.04025
R37433 VDD.n11061 VDD.n11060 0.04025
R37434 VDD.n11061 VDD.n664 0.04025
R37435 VDD.n11066 VDD.n664 0.04025
R37436 VDD.n11067 VDD.n11066 0.04025
R37437 VDD.n11068 VDD.n11067 0.04025
R37438 VDD.n11068 VDD.n662 0.04025
R37439 VDD.n11072 VDD.n662 0.04025
R37440 VDD.n11073 VDD.n11072 0.04025
R37441 VDD.n11073 VDD.n660 0.04025
R37442 VDD.n11079 VDD.n660 0.04025
R37443 VDD.n11080 VDD.n11079 0.04025
R37444 VDD.n11081 VDD.n11080 0.04025
R37445 VDD.n11081 VDD.n658 0.04025
R37446 VDD.n11085 VDD.n658 0.04025
R37447 VDD.n11086 VDD.n11085 0.04025
R37448 VDD.n11086 VDD.n656 0.04025
R37449 VDD.n11092 VDD.n656 0.04025
R37450 VDD.n11093 VDD.n11092 0.04025
R37451 VDD.n11094 VDD.n11093 0.04025
R37452 VDD.n11094 VDD.n654 0.04025
R37453 VDD.n11099 VDD.n654 0.04025
R37454 VDD.n11100 VDD.n11099 0.04025
R37455 VDD.n11101 VDD.n11100 0.04025
R37456 VDD.n11101 VDD.n652 0.04025
R37457 VDD.n11105 VDD.n652 0.04025
R37458 VDD.n11106 VDD.n11105 0.04025
R37459 VDD.n11106 VDD.n650 0.04025
R37460 VDD.n11110 VDD.n650 0.04025
R37461 VDD.n11111 VDD.n11110 0.04025
R37462 VDD.n11111 VDD.n647 0.04025
R37463 VDD.n11115 VDD.n647 0.04025
R37464 VDD.n11116 VDD.n11115 0.04025
R37465 VDD.n11117 VDD.n11116 0.04025
R37466 VDD.n11117 VDD.n645 0.04025
R37467 VDD.n11122 VDD.n645 0.04025
R37468 VDD.n11124 VDD.n11122 0.04025
R37469 VDD.n11125 VDD.n11124 0.04025
R37470 VDD.n11125 VDD.n632 0.04025
R37471 VDD.n11132 VDD.n632 0.04025
R37472 VDD.n11133 VDD.n11132 0.04025
R37473 VDD.n11134 VDD.n11133 0.04025
R37474 VDD.n11134 VDD.n630 0.04025
R37475 VDD.n11138 VDD.n630 0.04025
R37476 VDD.n11139 VDD.n11138 0.04025
R37477 VDD.n11140 VDD.n11139 0.04025
R37478 VDD.n11140 VDD.n628 0.04025
R37479 VDD.n11144 VDD.n628 0.04025
R37480 VDD.n11145 VDD.n11144 0.04025
R37481 VDD.n11146 VDD.n11145 0.04025
R37482 VDD.n11146 VDD.n626 0.04025
R37483 VDD.n11150 VDD.n626 0.04025
R37484 VDD.n11151 VDD.n11150 0.04025
R37485 VDD.n11152 VDD.n11151 0.04025
R37486 VDD.n11152 VDD.n624 0.04025
R37487 VDD.n11156 VDD.n624 0.04025
R37488 VDD.n11157 VDD.n11156 0.04025
R37489 VDD.n11158 VDD.n11157 0.04025
R37490 VDD.n11158 VDD.n622 0.04025
R37491 VDD.n11162 VDD.n622 0.04025
R37492 VDD.n11163 VDD.n11162 0.04025
R37493 VDD.n11164 VDD.n11163 0.04025
R37494 VDD.n11164 VDD.n620 0.04025
R37495 VDD.n11168 VDD.n620 0.04025
R37496 VDD.n11169 VDD.n11168 0.04025
R37497 VDD.n11170 VDD.n11169 0.04025
R37498 VDD.n11170 VDD.n618 0.04025
R37499 VDD.n11174 VDD.n618 0.04025
R37500 VDD.n11175 VDD.n11174 0.04025
R37501 VDD.n11176 VDD.n11175 0.04025
R37502 VDD.n11176 VDD.n616 0.04025
R37503 VDD.n11180 VDD.n616 0.04025
R37504 VDD.n11181 VDD.n11180 0.04025
R37505 VDD.n11182 VDD.n11181 0.04025
R37506 VDD.n11182 VDD.n614 0.04025
R37507 VDD.n11186 VDD.n614 0.04025
R37508 VDD.n11187 VDD.n11186 0.04025
R37509 VDD.n11188 VDD.n11187 0.04025
R37510 VDD.n11188 VDD.n612 0.04025
R37511 VDD.n11192 VDD.n612 0.04025
R37512 VDD.n11193 VDD.n11192 0.04025
R37513 VDD.n11194 VDD.n11193 0.04025
R37514 VDD.n11194 VDD.n610 0.04025
R37515 VDD.n11198 VDD.n610 0.04025
R37516 VDD.n11199 VDD.n11198 0.04025
R37517 VDD.n11200 VDD.n11199 0.04025
R37518 VDD.n11200 VDD.n608 0.04025
R37519 VDD.n11204 VDD.n608 0.04025
R37520 VDD.n11205 VDD.n11204 0.04025
R37521 VDD.n11206 VDD.n11205 0.04025
R37522 VDD.n11206 VDD.n606 0.04025
R37523 VDD.n11210 VDD.n606 0.04025
R37524 VDD.n11211 VDD.n11210 0.04025
R37525 VDD.n11212 VDD.n11211 0.04025
R37526 VDD.n11212 VDD.n604 0.04025
R37527 VDD.n11216 VDD.n604 0.04025
R37528 VDD.n11217 VDD.n11216 0.04025
R37529 VDD.n11218 VDD.n11217 0.04025
R37530 VDD.n11218 VDD.n602 0.04025
R37531 VDD.n11222 VDD.n602 0.04025
R37532 VDD.n11223 VDD.n11222 0.04025
R37533 VDD.n11224 VDD.n11223 0.04025
R37534 VDD.n11224 VDD.n600 0.04025
R37535 VDD.n11228 VDD.n600 0.04025
R37536 VDD.n11229 VDD.n11228 0.04025
R37537 VDD.n11230 VDD.n11229 0.04025
R37538 VDD.n11230 VDD.n598 0.04025
R37539 VDD.n11234 VDD.n598 0.04025
R37540 VDD.n11235 VDD.n11234 0.04025
R37541 VDD.n11236 VDD.n11235 0.04025
R37542 VDD.n11236 VDD.n596 0.04025
R37543 VDD.n11240 VDD.n596 0.04025
R37544 VDD.n11241 VDD.n11240 0.04025
R37545 VDD.n11242 VDD.n11241 0.04025
R37546 VDD.n11242 VDD.n594 0.04025
R37547 VDD.n11246 VDD.n594 0.04025
R37548 VDD.n11247 VDD.n11246 0.04025
R37549 VDD.n11248 VDD.n11247 0.04025
R37550 VDD.n11248 VDD.n592 0.04025
R37551 VDD.n11252 VDD.n592 0.04025
R37552 VDD.n11253 VDD.n11252 0.04025
R37553 VDD.n11254 VDD.n11253 0.04025
R37554 VDD.n11254 VDD.n590 0.04025
R37555 VDD.n11258 VDD.n590 0.04025
R37556 VDD.n11259 VDD.n11258 0.04025
R37557 VDD.n11260 VDD.n11259 0.04025
R37558 VDD.n11260 VDD.n588 0.04025
R37559 VDD.n11264 VDD.n588 0.04025
R37560 VDD.n11265 VDD.n11264 0.04025
R37561 VDD.n11266 VDD.n11265 0.04025
R37562 VDD.n11266 VDD.n586 0.04025
R37563 VDD.n11270 VDD.n586 0.04025
R37564 VDD.n11271 VDD.n11270 0.04025
R37565 VDD.n11272 VDD.n11271 0.04025
R37566 VDD.n11272 VDD.n584 0.04025
R37567 VDD.n11276 VDD.n584 0.04025
R37568 VDD.n11277 VDD.n11276 0.04025
R37569 VDD.n11278 VDD.n11277 0.04025
R37570 VDD.n11278 VDD.n582 0.04025
R37571 VDD.n11282 VDD.n582 0.04025
R37572 VDD.n11283 VDD.n11282 0.04025
R37573 VDD.n11284 VDD.n11283 0.04025
R37574 VDD.n11284 VDD.n580 0.04025
R37575 VDD.n11288 VDD.n580 0.04025
R37576 VDD.n11289 VDD.n11288 0.04025
R37577 VDD.n11290 VDD.n11289 0.04025
R37578 VDD.n11290 VDD.n578 0.04025
R37579 VDD.n11294 VDD.n578 0.04025
R37580 VDD.n11295 VDD.n11294 0.04025
R37581 VDD.n11296 VDD.n11295 0.04025
R37582 VDD.n11296 VDD.n576 0.04025
R37583 VDD.n11300 VDD.n576 0.04025
R37584 VDD.n11301 VDD.n11300 0.04025
R37585 VDD.n11302 VDD.n11301 0.04025
R37586 VDD.n11302 VDD.n574 0.04025
R37587 VDD.n11306 VDD.n574 0.04025
R37588 VDD.n11307 VDD.n11306 0.04025
R37589 VDD.n11308 VDD.n11307 0.04025
R37590 VDD.n11308 VDD.n572 0.04025
R37591 VDD.n11312 VDD.n572 0.04025
R37592 VDD.n11313 VDD.n11312 0.04025
R37593 VDD.n11314 VDD.n11313 0.04025
R37594 VDD.n11314 VDD.n570 0.04025
R37595 VDD.n11318 VDD.n570 0.04025
R37596 VDD.n11319 VDD.n11318 0.04025
R37597 VDD.n11320 VDD.n11319 0.04025
R37598 VDD.n11320 VDD.n568 0.04025
R37599 VDD.n11324 VDD.n568 0.04025
R37600 VDD.n11325 VDD.n11324 0.04025
R37601 VDD.n11326 VDD.n11325 0.04025
R37602 VDD.n11326 VDD.n566 0.04025
R37603 VDD.n11330 VDD.n566 0.04025
R37604 VDD.n11331 VDD.n11330 0.04025
R37605 VDD.n11332 VDD.n11331 0.04025
R37606 VDD.n11332 VDD.n564 0.04025
R37607 VDD.n11336 VDD.n564 0.04025
R37608 VDD.n11337 VDD.n11336 0.04025
R37609 VDD.n11338 VDD.n11337 0.04025
R37610 VDD.n11338 VDD.n562 0.04025
R37611 VDD.n11342 VDD.n562 0.04025
R37612 VDD.n11343 VDD.n11342 0.04025
R37613 VDD.n11344 VDD.n11343 0.04025
R37614 VDD.n11344 VDD.n560 0.04025
R37615 VDD.n11348 VDD.n560 0.04025
R37616 VDD.n11349 VDD.n11348 0.04025
R37617 VDD.n11350 VDD.n11349 0.04025
R37618 VDD.n11350 VDD.n558 0.04025
R37619 VDD.n11354 VDD.n558 0.04025
R37620 VDD.n11355 VDD.n11354 0.04025
R37621 VDD.n11356 VDD.n11355 0.04025
R37622 VDD.n11356 VDD.n556 0.04025
R37623 VDD.n11360 VDD.n556 0.04025
R37624 VDD.n11361 VDD.n11360 0.04025
R37625 VDD.n11362 VDD.n11361 0.04025
R37626 VDD.n11362 VDD.n554 0.04025
R37627 VDD.n11366 VDD.n554 0.04025
R37628 VDD.n11367 VDD.n11366 0.04025
R37629 VDD.n11368 VDD.n11367 0.04025
R37630 VDD.n11368 VDD.n552 0.04025
R37631 VDD.n11372 VDD.n552 0.04025
R37632 VDD.n11373 VDD.n11372 0.04025
R37633 VDD.n11374 VDD.n11373 0.04025
R37634 VDD.n11374 VDD.n550 0.04025
R37635 VDD.n11378 VDD.n550 0.04025
R37636 VDD.n11379 VDD.n11378 0.04025
R37637 VDD.n11380 VDD.n11379 0.04025
R37638 VDD.n11380 VDD.n548 0.04025
R37639 VDD.n11384 VDD.n548 0.04025
R37640 VDD.n11385 VDD.n11384 0.04025
R37641 VDD.n11386 VDD.n11385 0.04025
R37642 VDD.n11386 VDD.n546 0.04025
R37643 VDD.n11390 VDD.n546 0.04025
R37644 VDD.n11391 VDD.n11390 0.04025
R37645 VDD.n11392 VDD.n11391 0.04025
R37646 VDD.n11392 VDD.n544 0.04025
R37647 VDD.n11396 VDD.n544 0.04025
R37648 VDD.n11397 VDD.n11396 0.04025
R37649 VDD.n11398 VDD.n11397 0.04025
R37650 VDD.n11398 VDD.n542 0.04025
R37651 VDD.n11402 VDD.n542 0.04025
R37652 VDD.n11403 VDD.n11402 0.04025
R37653 VDD.n11404 VDD.n11403 0.04025
R37654 VDD.n11404 VDD.n540 0.04025
R37655 VDD.n11408 VDD.n540 0.04025
R37656 VDD.n11409 VDD.n11408 0.04025
R37657 VDD.n11410 VDD.n11409 0.04025
R37658 VDD.n11410 VDD.n538 0.04025
R37659 VDD.n11414 VDD.n538 0.04025
R37660 VDD.n11415 VDD.n11414 0.04025
R37661 VDD.n11416 VDD.n11415 0.04025
R37662 VDD.n11416 VDD.n536 0.04025
R37663 VDD.n11420 VDD.n536 0.04025
R37664 VDD.n11421 VDD.n11420 0.04025
R37665 VDD.n11422 VDD.n11421 0.04025
R37666 VDD.n11422 VDD.n534 0.04025
R37667 VDD.n11426 VDD.n534 0.04025
R37668 VDD.n11427 VDD.n11426 0.04025
R37669 VDD.n11428 VDD.n11427 0.04025
R37670 VDD.n11428 VDD.n532 0.04025
R37671 VDD.n11432 VDD.n532 0.04025
R37672 VDD.n11433 VDD.n11432 0.04025
R37673 VDD.n11434 VDD.n11433 0.04025
R37674 VDD.n11434 VDD.n530 0.04025
R37675 VDD.n11438 VDD.n530 0.04025
R37676 VDD.n11439 VDD.n11438 0.04025
R37677 VDD.n11440 VDD.n11439 0.04025
R37678 VDD.n11440 VDD.n528 0.04025
R37679 VDD.n11444 VDD.n528 0.04025
R37680 VDD.n11445 VDD.n11444 0.04025
R37681 VDD.n11446 VDD.n11445 0.04025
R37682 VDD.n11446 VDD.n526 0.04025
R37683 VDD.n11450 VDD.n526 0.04025
R37684 VDD.n11451 VDD.n11450 0.04025
R37685 VDD.n11452 VDD.n11451 0.04025
R37686 VDD.n11452 VDD.n524 0.04025
R37687 VDD.n11456 VDD.n524 0.04025
R37688 VDD.n11457 VDD.n11456 0.04025
R37689 VDD.n11458 VDD.n11457 0.04025
R37690 VDD.n11458 VDD.n522 0.04025
R37691 VDD.n11462 VDD.n522 0.04025
R37692 VDD.n11463 VDD.n11462 0.04025
R37693 VDD.n11464 VDD.n11463 0.04025
R37694 VDD.n11464 VDD.n520 0.04025
R37695 VDD.n11468 VDD.n520 0.04025
R37696 VDD.n11469 VDD.n11468 0.04025
R37697 VDD.n11470 VDD.n11469 0.04025
R37698 VDD.n11470 VDD.n518 0.04025
R37699 VDD.n11474 VDD.n518 0.04025
R37700 VDD.n11475 VDD.n11474 0.04025
R37701 VDD.n11476 VDD.n11475 0.04025
R37702 VDD.n11476 VDD.n516 0.04025
R37703 VDD.n11480 VDD.n516 0.04025
R37704 VDD.n11481 VDD.n11480 0.04025
R37705 VDD.n11482 VDD.n11481 0.04025
R37706 VDD.n11482 VDD.n514 0.04025
R37707 VDD.n11486 VDD.n514 0.04025
R37708 VDD.n11487 VDD.n11486 0.04025
R37709 VDD.n11488 VDD.n11487 0.04025
R37710 VDD.n11488 VDD.n512 0.04025
R37711 VDD.n11492 VDD.n512 0.04025
R37712 VDD.n11493 VDD.n11492 0.04025
R37713 VDD.n11494 VDD.n11493 0.04025
R37714 VDD.n11494 VDD.n510 0.04025
R37715 VDD.n11498 VDD.n510 0.04025
R37716 VDD.n11499 VDD.n11498 0.04025
R37717 VDD.n11500 VDD.n11499 0.04025
R37718 VDD.n11500 VDD.n508 0.04025
R37719 VDD.n11504 VDD.n508 0.04025
R37720 VDD.n11505 VDD.n11504 0.04025
R37721 VDD.n11506 VDD.n11505 0.04025
R37722 VDD.n11506 VDD.n506 0.04025
R37723 VDD.n11510 VDD.n506 0.04025
R37724 VDD.n11511 VDD.n11510 0.04025
R37725 VDD.n11512 VDD.n11511 0.04025
R37726 VDD.n11512 VDD.n504 0.04025
R37727 VDD.n11516 VDD.n504 0.04025
R37728 VDD.n11517 VDD.n11516 0.04025
R37729 VDD.n11518 VDD.n11517 0.04025
R37730 VDD.n11518 VDD.n502 0.04025
R37731 VDD.n11522 VDD.n502 0.04025
R37732 VDD.n11523 VDD.n11522 0.04025
R37733 VDD.n11524 VDD.n11523 0.04025
R37734 VDD.n11524 VDD.n500 0.04025
R37735 VDD.n11528 VDD.n500 0.04025
R37736 VDD.n11529 VDD.n11528 0.04025
R37737 VDD.n11530 VDD.n11529 0.04025
R37738 VDD.n11530 VDD.n498 0.04025
R37739 VDD.n11534 VDD.n498 0.04025
R37740 VDD.n11535 VDD.n11534 0.04025
R37741 VDD.n11536 VDD.n11535 0.04025
R37742 VDD.n11536 VDD.n496 0.04025
R37743 VDD.n11540 VDD.n496 0.04025
R37744 VDD.n11541 VDD.n11540 0.04025
R37745 VDD.n11542 VDD.n11541 0.04025
R37746 VDD.n11542 VDD.n494 0.04025
R37747 VDD.n11546 VDD.n494 0.04025
R37748 VDD.n11547 VDD.n11546 0.04025
R37749 VDD.n11548 VDD.n11547 0.04025
R37750 VDD.n11548 VDD.n492 0.04025
R37751 VDD.n11552 VDD.n492 0.04025
R37752 VDD.n11553 VDD.n11552 0.04025
R37753 VDD.n11554 VDD.n11553 0.04025
R37754 VDD.n11554 VDD.n490 0.04025
R37755 VDD.n11558 VDD.n490 0.04025
R37756 VDD.n11559 VDD.n11558 0.04025
R37757 VDD.n11560 VDD.n11559 0.04025
R37758 VDD.n11560 VDD.n488 0.04025
R37759 VDD.n11564 VDD.n488 0.04025
R37760 VDD.n11565 VDD.n11564 0.04025
R37761 VDD.n11566 VDD.n11565 0.04025
R37762 VDD.n11566 VDD.n486 0.04025
R37763 VDD.n11570 VDD.n486 0.04025
R37764 VDD.n11571 VDD.n11570 0.04025
R37765 VDD.n11572 VDD.n11571 0.04025
R37766 VDD.n11572 VDD.n484 0.04025
R37767 VDD.n11576 VDD.n484 0.04025
R37768 VDD.n11577 VDD.n11576 0.04025
R37769 VDD.n11578 VDD.n11577 0.04025
R37770 VDD.n11578 VDD.n482 0.04025
R37771 VDD.n11582 VDD.n482 0.04025
R37772 VDD.n11583 VDD.n11582 0.04025
R37773 VDD.n11584 VDD.n11583 0.04025
R37774 VDD.n11584 VDD.n480 0.04025
R37775 VDD.n11588 VDD.n480 0.04025
R37776 VDD.n11589 VDD.n11588 0.04025
R37777 VDD.n11590 VDD.n11589 0.04025
R37778 VDD.n11590 VDD.n478 0.04025
R37779 VDD.n11594 VDD.n478 0.04025
R37780 VDD.n11595 VDD.n11594 0.04025
R37781 VDD.n11596 VDD.n11595 0.04025
R37782 VDD.n11596 VDD.n476 0.04025
R37783 VDD.n11600 VDD.n476 0.04025
R37784 VDD.n11601 VDD.n11600 0.04025
R37785 VDD.n11602 VDD.n11601 0.04025
R37786 VDD.n11602 VDD.n474 0.04025
R37787 VDD.n11606 VDD.n474 0.04025
R37788 VDD.n11607 VDD.n11606 0.04025
R37789 VDD.n11608 VDD.n11607 0.04025
R37790 VDD.n11608 VDD.n472 0.04025
R37791 VDD.n11612 VDD.n472 0.04025
R37792 VDD.n11613 VDD.n11612 0.04025
R37793 VDD.n11614 VDD.n11613 0.04025
R37794 VDD.n11614 VDD.n470 0.04025
R37795 VDD.n11618 VDD.n470 0.04025
R37796 VDD.n11619 VDD.n11618 0.04025
R37797 VDD.n11620 VDD.n11619 0.04025
R37798 VDD.n11620 VDD.n468 0.04025
R37799 VDD.n11624 VDD.n468 0.04025
R37800 VDD.n11625 VDD.n11624 0.04025
R37801 VDD.n11626 VDD.n11625 0.04025
R37802 VDD.n11626 VDD.n466 0.04025
R37803 VDD.n11630 VDD.n466 0.04025
R37804 VDD.n11631 VDD.n11630 0.04025
R37805 VDD.n11632 VDD.n11631 0.04025
R37806 VDD.n11632 VDD.n464 0.04025
R37807 VDD.n11636 VDD.n464 0.04025
R37808 VDD.n11637 VDD.n11636 0.04025
R37809 VDD.n11638 VDD.n11637 0.04025
R37810 VDD.n11638 VDD.n462 0.04025
R37811 VDD.n11642 VDD.n462 0.04025
R37812 VDD.n11643 VDD.n11642 0.04025
R37813 VDD.n11644 VDD.n11643 0.04025
R37814 VDD.n11644 VDD.n460 0.04025
R37815 VDD.n11648 VDD.n460 0.04025
R37816 VDD.n11649 VDD.n11648 0.04025
R37817 VDD.n11650 VDD.n11649 0.04025
R37818 VDD.n11650 VDD.n458 0.04025
R37819 VDD.n11654 VDD.n458 0.04025
R37820 VDD.n11655 VDD.n11654 0.04025
R37821 VDD.n11656 VDD.n11655 0.04025
R37822 VDD.n11656 VDD.n456 0.04025
R37823 VDD.n11660 VDD.n456 0.04025
R37824 VDD.n11661 VDD.n11660 0.04025
R37825 VDD.n11662 VDD.n11661 0.04025
R37826 VDD.n11662 VDD.n454 0.04025
R37827 VDD.n11666 VDD.n454 0.04025
R37828 VDD.n11667 VDD.n11666 0.04025
R37829 VDD.n11668 VDD.n11667 0.04025
R37830 VDD.n11668 VDD.n452 0.04025
R37831 VDD.n11672 VDD.n452 0.04025
R37832 VDD.n11673 VDD.n11672 0.04025
R37833 VDD.n11674 VDD.n11673 0.04025
R37834 VDD.n11674 VDD.n450 0.04025
R37835 VDD.n11678 VDD.n450 0.04025
R37836 VDD.n11679 VDD.n11678 0.04025
R37837 VDD.n11680 VDD.n11679 0.04025
R37838 VDD.n11680 VDD.n448 0.04025
R37839 VDD.n11684 VDD.n448 0.04025
R37840 VDD.n11685 VDD.n11684 0.04025
R37841 VDD.n11686 VDD.n11685 0.04025
R37842 VDD.n11686 VDD.n446 0.04025
R37843 VDD.n11690 VDD.n446 0.04025
R37844 VDD.n11691 VDD.n11690 0.04025
R37845 VDD.n11692 VDD.n11691 0.04025
R37846 VDD.n11692 VDD.n444 0.04025
R37847 VDD.n11696 VDD.n444 0.04025
R37848 VDD.n11697 VDD.n11696 0.04025
R37849 VDD.n11698 VDD.n11697 0.04025
R37850 VDD.n11698 VDD.n442 0.04025
R37851 VDD.n11702 VDD.n442 0.04025
R37852 VDD.n11703 VDD.n11702 0.04025
R37853 VDD.n11704 VDD.n11703 0.04025
R37854 VDD.n11704 VDD.n440 0.04025
R37855 VDD.n11708 VDD.n440 0.04025
R37856 VDD.n11709 VDD.n11708 0.04025
R37857 VDD.n11710 VDD.n11709 0.04025
R37858 VDD.n11710 VDD.n438 0.04025
R37859 VDD.n11714 VDD.n438 0.04025
R37860 VDD.n11715 VDD.n11714 0.04025
R37861 VDD.n11716 VDD.n11715 0.04025
R37862 VDD.n11716 VDD.n436 0.04025
R37863 VDD.n11720 VDD.n436 0.04025
R37864 VDD.n11721 VDD.n11720 0.04025
R37865 VDD.n11722 VDD.n11721 0.04025
R37866 VDD.n11722 VDD.n434 0.04025
R37867 VDD.n11726 VDD.n434 0.04025
R37868 VDD.n11727 VDD.n11726 0.04025
R37869 VDD.n11728 VDD.n11727 0.04025
R37870 VDD.n11728 VDD.n432 0.04025
R37871 VDD.n11732 VDD.n432 0.04025
R37872 VDD.n11733 VDD.n11732 0.04025
R37873 VDD.n11734 VDD.n11733 0.04025
R37874 VDD.n11734 VDD.n430 0.04025
R37875 VDD.n11738 VDD.n430 0.04025
R37876 VDD.n11739 VDD.n11738 0.04025
R37877 VDD.n11740 VDD.n11739 0.04025
R37878 VDD.n11740 VDD.n428 0.04025
R37879 VDD.n11744 VDD.n428 0.04025
R37880 VDD.n11745 VDD.n11744 0.04025
R37881 VDD.n11746 VDD.n11745 0.04025
R37882 VDD.n11746 VDD.n426 0.04025
R37883 VDD.n11750 VDD.n426 0.04025
R37884 VDD.n11751 VDD.n11750 0.04025
R37885 VDD.n11752 VDD.n11751 0.04025
R37886 VDD.n11752 VDD.n424 0.04025
R37887 VDD.n11756 VDD.n424 0.04025
R37888 VDD.n11757 VDD.n11756 0.04025
R37889 VDD.n11758 VDD.n11757 0.04025
R37890 VDD.n11758 VDD.n422 0.04025
R37891 VDD.n11762 VDD.n422 0.04025
R37892 VDD.n11763 VDD.n11762 0.04025
R37893 VDD.n11764 VDD.n11763 0.04025
R37894 VDD.n11764 VDD.n420 0.04025
R37895 VDD.n11768 VDD.n420 0.04025
R37896 VDD.n11769 VDD.n11768 0.04025
R37897 VDD.n11770 VDD.n11769 0.04025
R37898 VDD.n11770 VDD.n418 0.04025
R37899 VDD.n11774 VDD.n418 0.04025
R37900 VDD.n11775 VDD.n11774 0.04025
R37901 VDD.n11776 VDD.n11775 0.04025
R37902 VDD.n11776 VDD.n416 0.04025
R37903 VDD.n11780 VDD.n416 0.04025
R37904 VDD.n11781 VDD.n11780 0.04025
R37905 VDD.n11782 VDD.n11781 0.04025
R37906 VDD.n11782 VDD.n414 0.04025
R37907 VDD.n11786 VDD.n414 0.04025
R37908 VDD.n11787 VDD.n11786 0.04025
R37909 VDD.n11788 VDD.n11787 0.04025
R37910 VDD.n11788 VDD.n412 0.04025
R37911 VDD.n11792 VDD.n412 0.04025
R37912 VDD.n11793 VDD.n11792 0.04025
R37913 VDD.n11794 VDD.n11793 0.04025
R37914 VDD.n11794 VDD.n410 0.04025
R37915 VDD.n11798 VDD.n410 0.04025
R37916 VDD.n11799 VDD.n11798 0.04025
R37917 VDD.n11800 VDD.n11799 0.04025
R37918 VDD.n11800 VDD.n408 0.04025
R37919 VDD.n11804 VDD.n408 0.04025
R37920 VDD.n11805 VDD.n11804 0.04025
R37921 VDD.n11806 VDD.n11805 0.04025
R37922 VDD.n11806 VDD.n406 0.04025
R37923 VDD.n11810 VDD.n406 0.04025
R37924 VDD.n11811 VDD.n11810 0.04025
R37925 VDD.n11812 VDD.n404 0.04025
R37926 VDD.n11816 VDD.n404 0.04025
R37927 VDD.n11817 VDD.n11816 0.04025
R37928 VDD.n11818 VDD.n11817 0.04025
R37929 VDD.n11818 VDD.n402 0.04025
R37930 VDD.n11822 VDD.n402 0.04025
R37931 VDD.n11823 VDD.n11822 0.04025
R37932 VDD.n11824 VDD.n11823 0.04025
R37933 VDD.n11824 VDD.n400 0.04025
R37934 VDD.n11828 VDD.n400 0.04025
R37935 VDD.n11829 VDD.n11828 0.04025
R37936 VDD.n11830 VDD.n11829 0.04025
R37937 VDD.n11830 VDD.n398 0.04025
R37938 VDD.n11834 VDD.n398 0.04025
R37939 VDD.n11835 VDD.n11834 0.04025
R37940 VDD.n11836 VDD.n11835 0.04025
R37941 VDD.n11836 VDD.n396 0.04025
R37942 VDD.n11840 VDD.n396 0.04025
R37943 VDD.n11841 VDD.n11840 0.04025
R37944 VDD.n11842 VDD.n11841 0.04025
R37945 VDD.n11842 VDD.n394 0.04025
R37946 VDD.n11846 VDD.n394 0.04025
R37947 VDD.n11847 VDD.n11846 0.04025
R37948 VDD.n11848 VDD.n11847 0.04025
R37949 VDD.n11848 VDD.n392 0.04025
R37950 VDD.n11852 VDD.n392 0.04025
R37951 VDD.n11853 VDD.n11852 0.04025
R37952 VDD.n11854 VDD.n11853 0.04025
R37953 VDD.n11854 VDD.n390 0.04025
R37954 VDD.n11858 VDD.n390 0.04025
R37955 VDD.n11859 VDD.n11858 0.04025
R37956 VDD.n11860 VDD.n11859 0.04025
R37957 VDD.n11860 VDD.n388 0.04025
R37958 VDD.n11864 VDD.n388 0.04025
R37959 VDD.n11865 VDD.n11864 0.04025
R37960 VDD.n11866 VDD.n11865 0.04025
R37961 VDD.n11866 VDD.n386 0.04025
R37962 VDD.n11870 VDD.n386 0.04025
R37963 VDD.n11871 VDD.n11870 0.04025
R37964 VDD.n11873 VDD.n11871 0.04025
R37965 VDD.n11877 VDD.n384 0.04025
R37966 VDD.n11878 VDD.n11877 0.04025
R37967 VDD.n11879 VDD.n11878 0.04025
R37968 VDD.n11879 VDD.n382 0.04025
R37969 VDD.n11883 VDD.n382 0.04025
R37970 VDD.n11884 VDD.n11883 0.04025
R37971 VDD.n11885 VDD.n11884 0.04025
R37972 VDD.n11885 VDD.n380 0.04025
R37973 VDD.n11889 VDD.n380 0.04025
R37974 VDD.n11890 VDD.n11889 0.04025
R37975 VDD.n11891 VDD.n11890 0.04025
R37976 VDD.n11891 VDD.n378 0.04025
R37977 VDD.n11895 VDD.n378 0.04025
R37978 VDD.n11896 VDD.n11895 0.04025
R37979 VDD.n11897 VDD.n11896 0.04025
R37980 VDD.n11897 VDD.n376 0.04025
R37981 VDD.n11901 VDD.n376 0.04025
R37982 VDD.n11902 VDD.n11901 0.04025
R37983 VDD.n11903 VDD.n11902 0.04025
R37984 VDD.n11903 VDD.n374 0.04025
R37985 VDD.n11907 VDD.n374 0.04025
R37986 VDD.n11908 VDD.n11907 0.04025
R37987 VDD.n11909 VDD.n11908 0.04025
R37988 VDD.n11909 VDD.n372 0.04025
R37989 VDD.n11913 VDD.n372 0.04025
R37990 VDD.n11914 VDD.n11913 0.04025
R37991 VDD.n11915 VDD.n11914 0.04025
R37992 VDD.n11915 VDD.n370 0.04025
R37993 VDD.n11919 VDD.n370 0.04025
R37994 VDD.n11920 VDD.n11919 0.04025
R37995 VDD.n11921 VDD.n11920 0.04025
R37996 VDD.n11921 VDD.n368 0.04025
R37997 VDD.n11925 VDD.n368 0.04025
R37998 VDD.n11926 VDD.n11925 0.04025
R37999 VDD.n11927 VDD.n11926 0.04025
R38000 VDD.n11927 VDD.n366 0.04025
R38001 VDD.n11931 VDD.n366 0.04025
R38002 VDD.n11932 VDD.n11931 0.04025
R38003 VDD.n11933 VDD.n11932 0.04025
R38004 VDD.n11933 VDD.n364 0.04025
R38005 VDD.n11937 VDD.n364 0.04025
R38006 VDD.n11938 VDD.n11937 0.04025
R38007 VDD.n11939 VDD.n11938 0.04025
R38008 VDD.n11939 VDD.n362 0.04025
R38009 VDD.n11943 VDD.n362 0.04025
R38010 VDD.n11944 VDD.n11943 0.04025
R38011 VDD.n11945 VDD.n11944 0.04025
R38012 VDD.n11945 VDD.n360 0.04025
R38013 VDD.n11949 VDD.n360 0.04025
R38014 VDD.n11950 VDD.n11949 0.04025
R38015 VDD.n11951 VDD.n11950 0.04025
R38016 VDD.n11951 VDD.n358 0.04025
R38017 VDD.n11955 VDD.n358 0.04025
R38018 VDD.n11956 VDD.n11955 0.04025
R38019 VDD.n11957 VDD.n11956 0.04025
R38020 VDD.n11957 VDD.n356 0.04025
R38021 VDD.n11961 VDD.n356 0.04025
R38022 VDD.n11962 VDD.n11961 0.04025
R38023 VDD.n11963 VDD.n11962 0.04025
R38024 VDD.n11963 VDD.n354 0.04025
R38025 VDD.n11967 VDD.n354 0.04025
R38026 VDD.n11968 VDD.n11967 0.04025
R38027 VDD.n11969 VDD.n11968 0.04025
R38028 VDD.n11969 VDD.n352 0.04025
R38029 VDD.n11973 VDD.n352 0.04025
R38030 VDD.n11974 VDD.n11973 0.04025
R38031 VDD.n11975 VDD.n11974 0.04025
R38032 VDD.n11975 VDD.n350 0.04025
R38033 VDD.n11979 VDD.n350 0.04025
R38034 VDD.n11980 VDD.n11979 0.04025
R38035 VDD.n11981 VDD.n11980 0.04025
R38036 VDD.n11981 VDD.n348 0.04025
R38037 VDD.n11985 VDD.n348 0.04025
R38038 VDD.n11986 VDD.n11985 0.04025
R38039 VDD.n11987 VDD.n11986 0.04025
R38040 VDD.n11987 VDD.n346 0.04025
R38041 VDD.n11991 VDD.n346 0.04025
R38042 VDD.n11992 VDD.n11991 0.04025
R38043 VDD.n11993 VDD.n11992 0.04025
R38044 VDD.n11993 VDD.n344 0.04025
R38045 VDD.n11997 VDD.n344 0.04025
R38046 VDD.n11998 VDD.n11997 0.04025
R38047 VDD.n11999 VDD.n11998 0.04025
R38048 VDD.n11999 VDD.n342 0.04025
R38049 VDD.n12003 VDD.n342 0.04025
R38050 VDD.n12004 VDD.n12003 0.04025
R38051 VDD.n12005 VDD.n12004 0.04025
R38052 VDD.n12005 VDD.n340 0.04025
R38053 VDD.n12009 VDD.n340 0.04025
R38054 VDD.n12010 VDD.n12009 0.04025
R38055 VDD.n12011 VDD.n12010 0.04025
R38056 VDD.n12011 VDD.n338 0.04025
R38057 VDD.n12015 VDD.n338 0.04025
R38058 VDD.n12016 VDD.n12015 0.04025
R38059 VDD.n12017 VDD.n12016 0.04025
R38060 VDD.n12017 VDD.n336 0.04025
R38061 VDD.n12021 VDD.n336 0.04025
R38062 VDD.n12022 VDD.n12021 0.04025
R38063 VDD.n12023 VDD.n12022 0.04025
R38064 VDD.n12023 VDD.n334 0.04025
R38065 VDD.n12027 VDD.n334 0.04025
R38066 VDD.n12028 VDD.n12027 0.04025
R38067 VDD.n12029 VDD.n12028 0.04025
R38068 VDD.n12029 VDD.n332 0.04025
R38069 VDD.n12033 VDD.n332 0.04025
R38070 VDD.n12034 VDD.n12033 0.04025
R38071 VDD.n12035 VDD.n12034 0.04025
R38072 VDD.n12035 VDD.n330 0.04025
R38073 VDD.n12039 VDD.n330 0.04025
R38074 VDD.n12040 VDD.n12039 0.04025
R38075 VDD.n12041 VDD.n12040 0.04025
R38076 VDD.n12041 VDD.n328 0.04025
R38077 VDD.n12045 VDD.n328 0.04025
R38078 VDD.n12046 VDD.n12045 0.04025
R38079 VDD.n12047 VDD.n12046 0.04025
R38080 VDD.n12047 VDD.n326 0.04025
R38081 VDD.n12051 VDD.n326 0.04025
R38082 VDD.n12052 VDD.n12051 0.04025
R38083 VDD.n12053 VDD.n12052 0.04025
R38084 VDD.n12053 VDD.n324 0.04025
R38085 VDD.n12057 VDD.n324 0.04025
R38086 VDD.n12058 VDD.n12057 0.04025
R38087 VDD.n12059 VDD.n12058 0.04025
R38088 VDD.n12059 VDD.n322 0.04025
R38089 VDD.n12063 VDD.n322 0.04025
R38090 VDD.n12064 VDD.n12063 0.04025
R38091 VDD.n12065 VDD.n12064 0.04025
R38092 VDD.n12065 VDD.n320 0.04025
R38093 VDD.n12069 VDD.n320 0.04025
R38094 VDD.n12070 VDD.n12069 0.04025
R38095 VDD.n12071 VDD.n12070 0.04025
R38096 VDD.n12071 VDD.n318 0.04025
R38097 VDD.n12075 VDD.n318 0.04025
R38098 VDD.n12076 VDD.n12075 0.04025
R38099 VDD.n12077 VDD.n12076 0.04025
R38100 VDD.n12077 VDD.n316 0.04025
R38101 VDD.n12081 VDD.n316 0.04025
R38102 VDD.n12082 VDD.n12081 0.04025
R38103 VDD.n12083 VDD.n12082 0.04025
R38104 VDD.n12083 VDD.n314 0.04025
R38105 VDD.n12087 VDD.n314 0.04025
R38106 VDD.n12088 VDD.n12087 0.04025
R38107 VDD.n12089 VDD.n12088 0.04025
R38108 VDD.n12089 VDD.n312 0.04025
R38109 VDD.n12093 VDD.n312 0.04025
R38110 VDD.n12094 VDD.n12093 0.04025
R38111 VDD.n12095 VDD.n12094 0.04025
R38112 VDD.n12095 VDD.n310 0.04025
R38113 VDD.n12099 VDD.n310 0.04025
R38114 VDD.n12100 VDD.n12099 0.04025
R38115 VDD.n12101 VDD.n12100 0.04025
R38116 VDD.n12101 VDD.n308 0.04025
R38117 VDD.n12105 VDD.n308 0.04025
R38118 VDD.n12106 VDD.n12105 0.04025
R38119 VDD.n12107 VDD.n12106 0.04025
R38120 VDD.n12107 VDD.n306 0.04025
R38121 VDD.n12111 VDD.n306 0.04025
R38122 VDD.n12112 VDD.n12111 0.04025
R38123 VDD.n12113 VDD.n12112 0.04025
R38124 VDD.n12113 VDD.n304 0.04025
R38125 VDD.n12117 VDD.n304 0.04025
R38126 VDD.n12118 VDD.n12117 0.04025
R38127 VDD.n12119 VDD.n12118 0.04025
R38128 VDD.n12119 VDD.n302 0.04025
R38129 VDD.n12123 VDD.n302 0.04025
R38130 VDD.n12124 VDD.n12123 0.04025
R38131 VDD.n12125 VDD.n12124 0.04025
R38132 VDD.n12125 VDD.n300 0.04025
R38133 VDD.n12129 VDD.n300 0.04025
R38134 VDD.n12130 VDD.n12129 0.04025
R38135 VDD.n12131 VDD.n12130 0.04025
R38136 VDD.n12131 VDD.n298 0.04025
R38137 VDD.n12135 VDD.n298 0.04025
R38138 VDD.n12136 VDD.n12135 0.04025
R38139 VDD.n12137 VDD.n12136 0.04025
R38140 VDD.n12137 VDD.n296 0.04025
R38141 VDD.n12141 VDD.n296 0.04025
R38142 VDD.n12142 VDD.n12141 0.04025
R38143 VDD.n12143 VDD.n12142 0.04025
R38144 VDD.n12143 VDD.n294 0.04025
R38145 VDD.n12147 VDD.n294 0.04025
R38146 VDD.n12148 VDD.n12147 0.04025
R38147 VDD.n12149 VDD.n12148 0.04025
R38148 VDD.n12149 VDD.n292 0.04025
R38149 VDD.n12153 VDD.n292 0.04025
R38150 VDD.n12154 VDD.n12153 0.04025
R38151 VDD.n12155 VDD.n12154 0.04025
R38152 VDD.n12155 VDD.n290 0.04025
R38153 VDD.n12159 VDD.n290 0.04025
R38154 VDD.n12160 VDD.n12159 0.04025
R38155 VDD.n12161 VDD.n12160 0.04025
R38156 VDD.n12161 VDD.n288 0.04025
R38157 VDD.n12165 VDD.n288 0.04025
R38158 VDD.n12166 VDD.n12165 0.04025
R38159 VDD.n12167 VDD.n12166 0.04025
R38160 VDD.n12167 VDD.n286 0.04025
R38161 VDD.n12171 VDD.n286 0.04025
R38162 VDD.n12172 VDD.n12171 0.04025
R38163 VDD.n12173 VDD.n12172 0.04025
R38164 VDD.n12173 VDD.n284 0.04025
R38165 VDD.n12177 VDD.n284 0.04025
R38166 VDD.n12178 VDD.n12177 0.04025
R38167 VDD.n12179 VDD.n12178 0.04025
R38168 VDD.n12179 VDD.n282 0.04025
R38169 VDD.n12183 VDD.n282 0.04025
R38170 VDD.n12184 VDD.n12183 0.04025
R38171 VDD.n12185 VDD.n12184 0.04025
R38172 VDD.n12185 VDD.n280 0.04025
R38173 VDD.n12189 VDD.n280 0.04025
R38174 VDD.n12190 VDD.n12189 0.04025
R38175 VDD.n12191 VDD.n12190 0.04025
R38176 VDD.n12191 VDD.n278 0.04025
R38177 VDD.n12195 VDD.n278 0.04025
R38178 VDD.n12196 VDD.n12195 0.04025
R38179 VDD.n12197 VDD.n12196 0.04025
R38180 VDD.n12197 VDD.n276 0.04025
R38181 VDD.n12201 VDD.n276 0.04025
R38182 VDD.n12202 VDD.n12201 0.04025
R38183 VDD.n12203 VDD.n12202 0.04025
R38184 VDD.n12203 VDD.n274 0.04025
R38185 VDD.n12207 VDD.n274 0.04025
R38186 VDD.n12208 VDD.n12207 0.04025
R38187 VDD.n12209 VDD.n12208 0.04025
R38188 VDD.n12209 VDD.n272 0.04025
R38189 VDD.n12213 VDD.n272 0.04025
R38190 VDD.n12214 VDD.n12213 0.04025
R38191 VDD.n12215 VDD.n12214 0.04025
R38192 VDD.n12215 VDD.n270 0.04025
R38193 VDD.n12219 VDD.n270 0.04025
R38194 VDD.n12220 VDD.n12219 0.04025
R38195 VDD.n12221 VDD.n12220 0.04025
R38196 VDD.n12221 VDD.n268 0.04025
R38197 VDD.n12225 VDD.n268 0.04025
R38198 VDD.n12226 VDD.n12225 0.04025
R38199 VDD.n12227 VDD.n12226 0.04025
R38200 VDD.n12227 VDD.n266 0.04025
R38201 VDD.n12231 VDD.n266 0.04025
R38202 VDD.n12232 VDD.n12231 0.04025
R38203 VDD.n12233 VDD.n12232 0.04025
R38204 VDD.n12233 VDD.n264 0.04025
R38205 VDD.n12237 VDD.n264 0.04025
R38206 VDD.n12238 VDD.n12237 0.04025
R38207 VDD.n12239 VDD.n12238 0.04025
R38208 VDD.n12239 VDD.n262 0.04025
R38209 VDD.n12243 VDD.n262 0.04025
R38210 VDD.n12244 VDD.n12243 0.04025
R38211 VDD.n12245 VDD.n12244 0.04025
R38212 VDD.n12245 VDD.n260 0.04025
R38213 VDD.n12249 VDD.n260 0.04025
R38214 VDD.n12250 VDD.n12249 0.04025
R38215 VDD.n12251 VDD.n12250 0.04025
R38216 VDD.n12251 VDD.n258 0.04025
R38217 VDD.n12255 VDD.n258 0.04025
R38218 VDD.n12256 VDD.n12255 0.04025
R38219 VDD.n12257 VDD.n12256 0.04025
R38220 VDD.n12257 VDD.n256 0.04025
R38221 VDD.n12261 VDD.n256 0.04025
R38222 VDD.n12262 VDD.n12261 0.04025
R38223 VDD.n12263 VDD.n12262 0.04025
R38224 VDD.n12263 VDD.n254 0.04025
R38225 VDD.n12267 VDD.n254 0.04025
R38226 VDD.n12268 VDD.n12267 0.04025
R38227 VDD.n12269 VDD.n12268 0.04025
R38228 VDD.n12269 VDD.n252 0.04025
R38229 VDD.n12273 VDD.n252 0.04025
R38230 VDD.n12274 VDD.n12273 0.04025
R38231 VDD.n12275 VDD.n12274 0.04025
R38232 VDD.n12275 VDD.n250 0.04025
R38233 VDD.n12279 VDD.n250 0.04025
R38234 VDD.n12280 VDD.n12279 0.04025
R38235 VDD.n12281 VDD.n12280 0.04025
R38236 VDD.n12281 VDD.n248 0.04025
R38237 VDD.n12285 VDD.n248 0.04025
R38238 VDD.n12286 VDD.n12285 0.04025
R38239 VDD.n12287 VDD.n12286 0.04025
R38240 VDD.n12287 VDD.n246 0.04025
R38241 VDD.n12291 VDD.n246 0.04025
R38242 VDD.n12292 VDD.n12291 0.04025
R38243 VDD.n12293 VDD.n12292 0.04025
R38244 VDD.n12293 VDD.n244 0.04025
R38245 VDD.n12297 VDD.n244 0.04025
R38246 VDD.n12298 VDD.n12297 0.04025
R38247 VDD.n12299 VDD.n12298 0.04025
R38248 VDD.n12299 VDD.n242 0.04025
R38249 VDD.n12303 VDD.n242 0.04025
R38250 VDD.n12304 VDD.n12303 0.04025
R38251 VDD.n12305 VDD.n12304 0.04025
R38252 VDD.n12305 VDD.n240 0.04025
R38253 VDD.n12309 VDD.n240 0.04025
R38254 VDD.n12310 VDD.n12309 0.04025
R38255 VDD.n12311 VDD.n12310 0.04025
R38256 VDD.n12311 VDD.n238 0.04025
R38257 VDD.n12315 VDD.n238 0.04025
R38258 VDD.n12316 VDD.n12315 0.04025
R38259 VDD.n12317 VDD.n12316 0.04025
R38260 VDD.n12317 VDD.n236 0.04025
R38261 VDD.n12321 VDD.n236 0.04025
R38262 VDD.n12322 VDD.n12321 0.04025
R38263 VDD.n12323 VDD.n12322 0.04025
R38264 VDD.n12323 VDD.n234 0.04025
R38265 VDD.n12327 VDD.n234 0.04025
R38266 VDD.n12328 VDD.n12327 0.04025
R38267 VDD.n12329 VDD.n12328 0.04025
R38268 VDD.n12329 VDD.n232 0.04025
R38269 VDD.n12333 VDD.n232 0.04025
R38270 VDD.n12334 VDD.n12333 0.04025
R38271 VDD.n12335 VDD.n12334 0.04025
R38272 VDD.n12335 VDD.n230 0.04025
R38273 VDD.n12339 VDD.n230 0.04025
R38274 VDD.n12340 VDD.n12339 0.04025
R38275 VDD.n12341 VDD.n12340 0.04025
R38276 VDD.n12341 VDD.n228 0.04025
R38277 VDD.n12345 VDD.n228 0.04025
R38278 VDD.n12346 VDD.n12345 0.04025
R38279 VDD.n12347 VDD.n12346 0.04025
R38280 VDD.n12347 VDD.n226 0.04025
R38281 VDD.n12351 VDD.n226 0.04025
R38282 VDD.n12352 VDD.n12351 0.04025
R38283 VDD.n12353 VDD.n12352 0.04025
R38284 VDD.n12353 VDD.n224 0.04025
R38285 VDD.n12357 VDD.n224 0.04025
R38286 VDD.n12358 VDD.n12357 0.04025
R38287 VDD.n12359 VDD.n12358 0.04025
R38288 VDD.n12359 VDD.n222 0.04025
R38289 VDD.n12363 VDD.n222 0.04025
R38290 VDD.n12364 VDD.n12363 0.04025
R38291 VDD.n12365 VDD.n12364 0.04025
R38292 VDD.n12365 VDD.n220 0.04025
R38293 VDD.n12369 VDD.n220 0.04025
R38294 VDD.n12370 VDD.n12369 0.04025
R38295 VDD.n12371 VDD.n12370 0.04025
R38296 VDD.n12371 VDD.n218 0.04025
R38297 VDD.n12375 VDD.n218 0.04025
R38298 VDD.n12376 VDD.n12375 0.04025
R38299 VDD.n12377 VDD.n12376 0.04025
R38300 VDD.n12377 VDD.n216 0.04025
R38301 VDD.n12381 VDD.n216 0.04025
R38302 VDD.n12382 VDD.n12381 0.04025
R38303 VDD.n12383 VDD.n12382 0.04025
R38304 VDD.n12383 VDD.n214 0.04025
R38305 VDD.n12387 VDD.n214 0.04025
R38306 VDD.n12388 VDD.n12387 0.04025
R38307 VDD.n12389 VDD.n12388 0.04025
R38308 VDD.n12389 VDD.n212 0.04025
R38309 VDD.n12393 VDD.n212 0.04025
R38310 VDD.n12394 VDD.n12393 0.04025
R38311 VDD.n12395 VDD.n12394 0.04025
R38312 VDD.n12395 VDD.n210 0.04025
R38313 VDD.n12399 VDD.n210 0.04025
R38314 VDD.n12400 VDD.n12399 0.04025
R38315 VDD.n12401 VDD.n12400 0.04025
R38316 VDD.n12401 VDD.n208 0.04025
R38317 VDD.n12405 VDD.n208 0.04025
R38318 VDD.n12406 VDD.n12405 0.04025
R38319 VDD.n12407 VDD.n12406 0.04025
R38320 VDD.n12407 VDD.n206 0.04025
R38321 VDD.n12411 VDD.n206 0.04025
R38322 VDD.n12412 VDD.n12411 0.04025
R38323 VDD.n12413 VDD.n12412 0.04025
R38324 VDD.n12413 VDD.n204 0.04025
R38325 VDD.n12417 VDD.n204 0.04025
R38326 VDD.n12418 VDD.n12417 0.04025
R38327 VDD.n12419 VDD.n12418 0.04025
R38328 VDD.n12419 VDD.n202 0.04025
R38329 VDD.n12423 VDD.n202 0.04025
R38330 VDD.n12424 VDD.n12423 0.04025
R38331 VDD.n12425 VDD.n12424 0.04025
R38332 VDD.n12425 VDD.n200 0.04025
R38333 VDD.n12429 VDD.n200 0.04025
R38334 VDD.n12430 VDD.n12429 0.04025
R38335 VDD.n12431 VDD.n12430 0.04025
R38336 VDD.n12431 VDD.n198 0.04025
R38337 VDD.n12435 VDD.n198 0.04025
R38338 VDD.n12436 VDD.n12435 0.04025
R38339 VDD.n12437 VDD.n12436 0.04025
R38340 VDD.n12437 VDD.n196 0.04025
R38341 VDD.n12441 VDD.n196 0.04025
R38342 VDD.n12447 VDD.n12441 0.04025
R38343 VDD.n9437 VDD.n194 0.04025
R38344 VDD.n9438 VDD.n9437 0.04025
R38345 VDD.n9438 VDD.n9435 0.04025
R38346 VDD.n9442 VDD.n9435 0.04025
R38347 VDD.n9443 VDD.n9442 0.04025
R38348 VDD.n9444 VDD.n9443 0.04025
R38349 VDD.n9444 VDD.n9433 0.04025
R38350 VDD.n9448 VDD.n9433 0.04025
R38351 VDD.n9449 VDD.n9448 0.04025
R38352 VDD.n9450 VDD.n9449 0.04025
R38353 VDD.n9450 VDD.n9431 0.04025
R38354 VDD.n9454 VDD.n9431 0.04025
R38355 VDD.n9455 VDD.n9454 0.04025
R38356 VDD.n9456 VDD.n9455 0.04025
R38357 VDD.n9456 VDD.n9429 0.04025
R38358 VDD.n9460 VDD.n9429 0.04025
R38359 VDD.n9461 VDD.n9460 0.04025
R38360 VDD.n9462 VDD.n9461 0.04025
R38361 VDD.n9462 VDD.n9427 0.04025
R38362 VDD.n9466 VDD.n9427 0.04025
R38363 VDD.n9467 VDD.n9466 0.04025
R38364 VDD.n9468 VDD.n9467 0.04025
R38365 VDD.n9468 VDD.n9425 0.04025
R38366 VDD.n9472 VDD.n9425 0.04025
R38367 VDD.n9473 VDD.n9472 0.04025
R38368 VDD.n9474 VDD.n9473 0.04025
R38369 VDD.n9474 VDD.n9423 0.04025
R38370 VDD.n9478 VDD.n9423 0.04025
R38371 VDD.n9479 VDD.n9478 0.04025
R38372 VDD.n9480 VDD.n9479 0.04025
R38373 VDD.n9480 VDD.n9421 0.04025
R38374 VDD.n9484 VDD.n9421 0.04025
R38375 VDD.n9485 VDD.n9484 0.04025
R38376 VDD.n9486 VDD.n9485 0.04025
R38377 VDD.n9486 VDD.n9419 0.04025
R38378 VDD.n9490 VDD.n9419 0.04025
R38379 VDD.n9491 VDD.n9490 0.04025
R38380 VDD.n9492 VDD.n9491 0.04025
R38381 VDD.n9492 VDD.n9417 0.04025
R38382 VDD.n9496 VDD.n9417 0.04025
R38383 VDD.n9497 VDD.n9496 0.04025
R38384 VDD.n9498 VDD.n9497 0.04025
R38385 VDD.n9498 VDD.n9415 0.04025
R38386 VDD.n9502 VDD.n9415 0.04025
R38387 VDD.n9503 VDD.n9502 0.04025
R38388 VDD.n9504 VDD.n9503 0.04025
R38389 VDD.n9504 VDD.n9413 0.04025
R38390 VDD.n9508 VDD.n9413 0.04025
R38391 VDD.n9509 VDD.n9508 0.04025
R38392 VDD.n9510 VDD.n9509 0.04025
R38393 VDD.n9510 VDD.n9411 0.04025
R38394 VDD.n9514 VDD.n9411 0.04025
R38395 VDD.n9515 VDD.n9514 0.04025
R38396 VDD.n9516 VDD.n9515 0.04025
R38397 VDD.n9516 VDD.n9409 0.04025
R38398 VDD.n9520 VDD.n9409 0.04025
R38399 VDD.n9521 VDD.n9520 0.04025
R38400 VDD.n9522 VDD.n9521 0.04025
R38401 VDD.n9522 VDD.n9407 0.04025
R38402 VDD.n9526 VDD.n9407 0.04025
R38403 VDD.n9527 VDD.n9526 0.04025
R38404 VDD.n9528 VDD.n9527 0.04025
R38405 VDD.n9528 VDD.n9405 0.04025
R38406 VDD.n9532 VDD.n9405 0.04025
R38407 VDD.n9533 VDD.n9532 0.04025
R38408 VDD.n9534 VDD.n9533 0.04025
R38409 VDD.n9534 VDD.n9403 0.04025
R38410 VDD.n9538 VDD.n9403 0.04025
R38411 VDD.n9539 VDD.n9538 0.04025
R38412 VDD.n9540 VDD.n9539 0.04025
R38413 VDD.n9540 VDD.n9401 0.04025
R38414 VDD.n9544 VDD.n9401 0.04025
R38415 VDD.n9545 VDD.n9544 0.04025
R38416 VDD.n9546 VDD.n9545 0.04025
R38417 VDD.n9546 VDD.n9399 0.04025
R38418 VDD.n9550 VDD.n9399 0.04025
R38419 VDD.n9551 VDD.n9550 0.04025
R38420 VDD.n9552 VDD.n9551 0.04025
R38421 VDD.n9552 VDD.n9397 0.04025
R38422 VDD.n9556 VDD.n9397 0.04025
R38423 VDD.n9557 VDD.n9556 0.04025
R38424 VDD.n9558 VDD.n9557 0.04025
R38425 VDD.n9558 VDD.n9395 0.04025
R38426 VDD.n9562 VDD.n9395 0.04025
R38427 VDD.n9563 VDD.n9562 0.04025
R38428 VDD.n9564 VDD.n9563 0.04025
R38429 VDD.n9564 VDD.n9393 0.04025
R38430 VDD.n9568 VDD.n9393 0.04025
R38431 VDD.n9569 VDD.n9568 0.04025
R38432 VDD.n9570 VDD.n9569 0.04025
R38433 VDD.n9570 VDD.n9391 0.04025
R38434 VDD.n9574 VDD.n9391 0.04025
R38435 VDD.n9575 VDD.n9574 0.04025
R38436 VDD.n9576 VDD.n9575 0.04025
R38437 VDD.n9576 VDD.n9389 0.04025
R38438 VDD.n9580 VDD.n9389 0.04025
R38439 VDD.n9581 VDD.n9580 0.04025
R38440 VDD.n9582 VDD.n9581 0.04025
R38441 VDD.n9582 VDD.n9387 0.04025
R38442 VDD.n9586 VDD.n9387 0.04025
R38443 VDD.n9587 VDD.n9586 0.04025
R38444 VDD.n9588 VDD.n9587 0.04025
R38445 VDD.n9588 VDD.n9385 0.04025
R38446 VDD.n9592 VDD.n9385 0.04025
R38447 VDD.n9593 VDD.n9592 0.04025
R38448 VDD.n9594 VDD.n9593 0.04025
R38449 VDD.n9594 VDD.n9383 0.04025
R38450 VDD.n9598 VDD.n9383 0.04025
R38451 VDD.n9599 VDD.n9598 0.04025
R38452 VDD.n9600 VDD.n9599 0.04025
R38453 VDD.n9600 VDD.n9381 0.04025
R38454 VDD.n9604 VDD.n9381 0.04025
R38455 VDD.n9605 VDD.n9604 0.04025
R38456 VDD.n9606 VDD.n9605 0.04025
R38457 VDD.n9606 VDD.n9379 0.04025
R38458 VDD.n9610 VDD.n9379 0.04025
R38459 VDD.n9611 VDD.n9610 0.04025
R38460 VDD.n9612 VDD.n9611 0.04025
R38461 VDD.n9612 VDD.n9377 0.04025
R38462 VDD.n9616 VDD.n9377 0.04025
R38463 VDD.n9617 VDD.n9616 0.04025
R38464 VDD.n9618 VDD.n9617 0.04025
R38465 VDD.n9618 VDD.n9375 0.04025
R38466 VDD.n9622 VDD.n9375 0.04025
R38467 VDD.n9623 VDD.n9622 0.04025
R38468 VDD.n9624 VDD.n9623 0.04025
R38469 VDD.n9624 VDD.n9373 0.04025
R38470 VDD.n9628 VDD.n9373 0.04025
R38471 VDD.n9629 VDD.n9628 0.04025
R38472 VDD.n9630 VDD.n9629 0.04025
R38473 VDD.n9630 VDD.n9371 0.04025
R38474 VDD.n9634 VDD.n9371 0.04025
R38475 VDD.n9635 VDD.n9634 0.04025
R38476 VDD.n9636 VDD.n9635 0.04025
R38477 VDD.n9636 VDD.n9369 0.04025
R38478 VDD.n9640 VDD.n9369 0.04025
R38479 VDD.n9641 VDD.n9640 0.04025
R38480 VDD.n9642 VDD.n9641 0.04025
R38481 VDD.n9642 VDD.n9367 0.04025
R38482 VDD.n9646 VDD.n9367 0.04025
R38483 VDD.n9647 VDD.n9646 0.04025
R38484 VDD.n9648 VDD.n9647 0.04025
R38485 VDD.n9648 VDD.n9365 0.04025
R38486 VDD.n9652 VDD.n9365 0.04025
R38487 VDD.n9653 VDD.n9652 0.04025
R38488 VDD.n9654 VDD.n9653 0.04025
R38489 VDD.n9654 VDD.n9363 0.04025
R38490 VDD.n9658 VDD.n9363 0.04025
R38491 VDD.n9659 VDD.n9658 0.04025
R38492 VDD.n9660 VDD.n9659 0.04025
R38493 VDD.n9660 VDD.n9361 0.04025
R38494 VDD.n9664 VDD.n9361 0.04025
R38495 VDD.n9665 VDD.n9664 0.04025
R38496 VDD.n9666 VDD.n9665 0.04025
R38497 VDD.n9666 VDD.n9359 0.04025
R38498 VDD.n9670 VDD.n9359 0.04025
R38499 VDD.n9671 VDD.n9670 0.04025
R38500 VDD.n9672 VDD.n9671 0.04025
R38501 VDD.n9672 VDD.n9357 0.04025
R38502 VDD.n9676 VDD.n9357 0.04025
R38503 VDD.n9677 VDD.n9676 0.04025
R38504 VDD.n9678 VDD.n9677 0.04025
R38505 VDD.n9678 VDD.n9355 0.04025
R38506 VDD.n9682 VDD.n9355 0.04025
R38507 VDD.n9683 VDD.n9682 0.04025
R38508 VDD.n9684 VDD.n9683 0.04025
R38509 VDD.n9684 VDD.n9353 0.04025
R38510 VDD.n9688 VDD.n9353 0.04025
R38511 VDD.n9689 VDD.n9688 0.04025
R38512 VDD.n9690 VDD.n9689 0.04025
R38513 VDD.n9690 VDD.n9351 0.04025
R38514 VDD.n9694 VDD.n9351 0.04025
R38515 VDD.n9695 VDD.n9694 0.04025
R38516 VDD.n9696 VDD.n9695 0.04025
R38517 VDD.n9696 VDD.n9349 0.04025
R38518 VDD.n9700 VDD.n9349 0.04025
R38519 VDD.n9701 VDD.n9700 0.04025
R38520 VDD.n9702 VDD.n9701 0.04025
R38521 VDD.n9702 VDD.n9347 0.04025
R38522 VDD.n9706 VDD.n9347 0.04025
R38523 VDD.n9707 VDD.n9706 0.04025
R38524 VDD.n9708 VDD.n9707 0.04025
R38525 VDD.n9708 VDD.n9345 0.04025
R38526 VDD.n9712 VDD.n9345 0.04025
R38527 VDD.n9713 VDD.n9712 0.04025
R38528 VDD.n9714 VDD.n9713 0.04025
R38529 VDD.n9714 VDD.n9343 0.04025
R38530 VDD.n9718 VDD.n9343 0.04025
R38531 VDD.n9719 VDD.n9718 0.04025
R38532 VDD.n9720 VDD.n9719 0.04025
R38533 VDD.n9720 VDD.n9341 0.04025
R38534 VDD.n9724 VDD.n9341 0.04025
R38535 VDD.n9725 VDD.n9724 0.04025
R38536 VDD.n9726 VDD.n9725 0.04025
R38537 VDD.n9726 VDD.n9339 0.04025
R38538 VDD.n9730 VDD.n9339 0.04025
R38539 VDD.n9731 VDD.n9730 0.04025
R38540 VDD.n9732 VDD.n9731 0.04025
R38541 VDD.n9732 VDD.n9337 0.04025
R38542 VDD.n9736 VDD.n9337 0.04025
R38543 VDD.n9737 VDD.n9736 0.04025
R38544 VDD.n9738 VDD.n9737 0.04025
R38545 VDD.n9738 VDD.n9335 0.04025
R38546 VDD.n9742 VDD.n9335 0.04025
R38547 VDD.n9743 VDD.n9742 0.04025
R38548 VDD.n9744 VDD.n9743 0.04025
R38549 VDD.n9744 VDD.n9333 0.04025
R38550 VDD.n9748 VDD.n9333 0.04025
R38551 VDD.n9749 VDD.n9748 0.04025
R38552 VDD.n9750 VDD.n9749 0.04025
R38553 VDD.n9750 VDD.n9331 0.04025
R38554 VDD.n9754 VDD.n9331 0.04025
R38555 VDD.n9755 VDD.n9754 0.04025
R38556 VDD.n9756 VDD.n9755 0.04025
R38557 VDD.n9756 VDD.n9329 0.04025
R38558 VDD.n9760 VDD.n9329 0.04025
R38559 VDD.n9761 VDD.n9760 0.04025
R38560 VDD.n9762 VDD.n9761 0.04025
R38561 VDD.n9762 VDD.n9327 0.04025
R38562 VDD.n9766 VDD.n9327 0.04025
R38563 VDD.n9767 VDD.n9766 0.04025
R38564 VDD.n9768 VDD.n9767 0.04025
R38565 VDD.n9768 VDD.n9325 0.04025
R38566 VDD.n9772 VDD.n9325 0.04025
R38567 VDD.n9773 VDD.n9772 0.04025
R38568 VDD.n9774 VDD.n9773 0.04025
R38569 VDD.n9774 VDD.n9323 0.04025
R38570 VDD.n9778 VDD.n9323 0.04025
R38571 VDD.n9779 VDD.n9778 0.04025
R38572 VDD.n9780 VDD.n9779 0.04025
R38573 VDD.n9780 VDD.n9321 0.04025
R38574 VDD.n9784 VDD.n9321 0.04025
R38575 VDD.n9785 VDD.n9784 0.04025
R38576 VDD.n9786 VDD.n9785 0.04025
R38577 VDD.n9786 VDD.n9319 0.04025
R38578 VDD.n9790 VDD.n9319 0.04025
R38579 VDD.n9791 VDD.n9790 0.04025
R38580 VDD.n9792 VDD.n9791 0.04025
R38581 VDD.n9792 VDD.n9317 0.04025
R38582 VDD.n9796 VDD.n9317 0.04025
R38583 VDD.n9797 VDD.n9796 0.04025
R38584 VDD.n9798 VDD.n9797 0.04025
R38585 VDD.n9798 VDD.n9315 0.04025
R38586 VDD.n9802 VDD.n9315 0.04025
R38587 VDD.n9803 VDD.n9802 0.04025
R38588 VDD.n9804 VDD.n9803 0.04025
R38589 VDD.n9804 VDD.n9313 0.04025
R38590 VDD.n9808 VDD.n9313 0.04025
R38591 VDD.n9809 VDD.n9808 0.04025
R38592 VDD.n9810 VDD.n9809 0.04025
R38593 VDD.n9810 VDD.n9311 0.04025
R38594 VDD.n9814 VDD.n9311 0.04025
R38595 VDD.n9815 VDD.n9814 0.04025
R38596 VDD.n9816 VDD.n9815 0.04025
R38597 VDD.n9816 VDD.n9309 0.04025
R38598 VDD.n9820 VDD.n9309 0.04025
R38599 VDD.n9821 VDD.n9820 0.04025
R38600 VDD.n9822 VDD.n9821 0.04025
R38601 VDD.n9822 VDD.n9307 0.04025
R38602 VDD.n9826 VDD.n9307 0.04025
R38603 VDD.n9827 VDD.n9826 0.04025
R38604 VDD.n9828 VDD.n9827 0.04025
R38605 VDD.n9828 VDD.n9305 0.04025
R38606 VDD.n9832 VDD.n9305 0.04025
R38607 VDD.n9833 VDD.n9832 0.04025
R38608 VDD.n9834 VDD.n9833 0.04025
R38609 VDD.n9834 VDD.n9303 0.04025
R38610 VDD.n9838 VDD.n9303 0.04025
R38611 VDD.n9839 VDD.n9838 0.04025
R38612 VDD.n9840 VDD.n9839 0.04025
R38613 VDD.n9840 VDD.n9301 0.04025
R38614 VDD.n9844 VDD.n9301 0.04025
R38615 VDD.n9845 VDD.n9844 0.04025
R38616 VDD.n9846 VDD.n9845 0.04025
R38617 VDD.n9846 VDD.n9299 0.04025
R38618 VDD.n9850 VDD.n9299 0.04025
R38619 VDD.n9851 VDD.n9850 0.04025
R38620 VDD.n9852 VDD.n9851 0.04025
R38621 VDD.n9852 VDD.n9297 0.04025
R38622 VDD.n9856 VDD.n9297 0.04025
R38623 VDD.n9857 VDD.n9856 0.04025
R38624 VDD.n9858 VDD.n9857 0.04025
R38625 VDD.n9858 VDD.n9295 0.04025
R38626 VDD.n9862 VDD.n9295 0.04025
R38627 VDD.n9863 VDD.n9862 0.04025
R38628 VDD.n9864 VDD.n9863 0.04025
R38629 VDD.n9864 VDD.n9293 0.04025
R38630 VDD.n9868 VDD.n9293 0.04025
R38631 VDD.n9869 VDD.n9868 0.04025
R38632 VDD.n9870 VDD.n9869 0.04025
R38633 VDD.n9870 VDD.n9291 0.04025
R38634 VDD.n9874 VDD.n9291 0.04025
R38635 VDD.n9875 VDD.n9874 0.04025
R38636 VDD.n9876 VDD.n9875 0.04025
R38637 VDD.n9876 VDD.n9289 0.04025
R38638 VDD.n9880 VDD.n9289 0.04025
R38639 VDD.n9881 VDD.n9880 0.04025
R38640 VDD.n9882 VDD.n9881 0.04025
R38641 VDD.n9882 VDD.n9287 0.04025
R38642 VDD.n9886 VDD.n9287 0.04025
R38643 VDD.n9887 VDD.n9886 0.04025
R38644 VDD.n9888 VDD.n9887 0.04025
R38645 VDD.n9888 VDD.n9285 0.04025
R38646 VDD.n9892 VDD.n9285 0.04025
R38647 VDD.n9893 VDD.n9892 0.04025
R38648 VDD.n9894 VDD.n9893 0.04025
R38649 VDD.n9894 VDD.n9283 0.04025
R38650 VDD.n9898 VDD.n9283 0.04025
R38651 VDD.n9899 VDD.n9898 0.04025
R38652 VDD.n9900 VDD.n9899 0.04025
R38653 VDD.n9900 VDD.n9281 0.04025
R38654 VDD.n9904 VDD.n9281 0.04025
R38655 VDD.n9905 VDD.n9904 0.04025
R38656 VDD.n9906 VDD.n9905 0.04025
R38657 VDD.n9906 VDD.n9279 0.04025
R38658 VDD.n9910 VDD.n9279 0.04025
R38659 VDD.n9911 VDD.n9910 0.04025
R38660 VDD.n9912 VDD.n9911 0.04025
R38661 VDD.n9912 VDD.n9277 0.04025
R38662 VDD.n9916 VDD.n9277 0.04025
R38663 VDD.n9917 VDD.n9916 0.04025
R38664 VDD.n9918 VDD.n9917 0.04025
R38665 VDD.n9918 VDD.n9275 0.04025
R38666 VDD.n9922 VDD.n9275 0.04025
R38667 VDD.n9923 VDD.n9922 0.04025
R38668 VDD.n9924 VDD.n9923 0.04025
R38669 VDD.n9924 VDD.n9273 0.04025
R38670 VDD.n9928 VDD.n9273 0.04025
R38671 VDD.n9929 VDD.n9928 0.04025
R38672 VDD.n9930 VDD.n9929 0.04025
R38673 VDD.n9930 VDD.n9271 0.04025
R38674 VDD.n9934 VDD.n9271 0.04025
R38675 VDD.n9935 VDD.n9934 0.04025
R38676 VDD.n9936 VDD.n9935 0.04025
R38677 VDD.n9936 VDD.n9269 0.04025
R38678 VDD.n9940 VDD.n9269 0.04025
R38679 VDD.n9941 VDD.n9940 0.04025
R38680 VDD.n9942 VDD.n9941 0.04025
R38681 VDD.n9942 VDD.n9267 0.04025
R38682 VDD.n9946 VDD.n9267 0.04025
R38683 VDD.n9947 VDD.n9946 0.04025
R38684 VDD.n9948 VDD.n9947 0.04025
R38685 VDD.n9948 VDD.n9265 0.04025
R38686 VDD.n9952 VDD.n9265 0.04025
R38687 VDD.n9953 VDD.n9952 0.04025
R38688 VDD.n9954 VDD.n9953 0.04025
R38689 VDD.n9954 VDD.n9263 0.04025
R38690 VDD.n9958 VDD.n9263 0.04025
R38691 VDD.n9959 VDD.n9958 0.04025
R38692 VDD.n9960 VDD.n9959 0.04025
R38693 VDD.n9960 VDD.n9261 0.04025
R38694 VDD.n9964 VDD.n9261 0.04025
R38695 VDD.n9965 VDD.n9964 0.04025
R38696 VDD.n9966 VDD.n9965 0.04025
R38697 VDD.n9966 VDD.n9259 0.04025
R38698 VDD.n9970 VDD.n9259 0.04025
R38699 VDD.n9971 VDD.n9970 0.04025
R38700 VDD.n9972 VDD.n9971 0.04025
R38701 VDD.n9972 VDD.n9257 0.04025
R38702 VDD.n9976 VDD.n9257 0.04025
R38703 VDD.n9977 VDD.n9976 0.04025
R38704 VDD.n9978 VDD.n9977 0.04025
R38705 VDD.n9978 VDD.n9255 0.04025
R38706 VDD.n9982 VDD.n9255 0.04025
R38707 VDD.n9983 VDD.n9982 0.04025
R38708 VDD.n9984 VDD.n9983 0.04025
R38709 VDD.n9984 VDD.n9253 0.04025
R38710 VDD.n9988 VDD.n9253 0.04025
R38711 VDD.n9989 VDD.n9988 0.04025
R38712 VDD.n9990 VDD.n9989 0.04025
R38713 VDD.n9990 VDD.n9251 0.04025
R38714 VDD.n9994 VDD.n9251 0.04025
R38715 VDD.n9995 VDD.n9994 0.04025
R38716 VDD.n9996 VDD.n9995 0.04025
R38717 VDD.n9996 VDD.n9249 0.04025
R38718 VDD.n10000 VDD.n9249 0.04025
R38719 VDD.n10001 VDD.n10000 0.04025
R38720 VDD.n10002 VDD.n10001 0.04025
R38721 VDD.n10002 VDD.n9247 0.04025
R38722 VDD.n10006 VDD.n9247 0.04025
R38723 VDD.n10007 VDD.n10006 0.04025
R38724 VDD.n10008 VDD.n10007 0.04025
R38725 VDD.n10008 VDD.n9245 0.04025
R38726 VDD.n10012 VDD.n9245 0.04025
R38727 VDD.n10013 VDD.n10012 0.04025
R38728 VDD.n10014 VDD.n10013 0.04025
R38729 VDD.n10014 VDD.n9243 0.04025
R38730 VDD.n10018 VDD.n9243 0.04025
R38731 VDD.n10019 VDD.n10018 0.04025
R38732 VDD.n10020 VDD.n10019 0.04025
R38733 VDD.n10020 VDD.n9241 0.04025
R38734 VDD.n10024 VDD.n9241 0.04025
R38735 VDD.n10025 VDD.n10024 0.04025
R38736 VDD.n10026 VDD.n10025 0.04025
R38737 VDD.n10026 VDD.n9239 0.04025
R38738 VDD.n10030 VDD.n9239 0.04025
R38739 VDD.n10031 VDD.n10030 0.04025
R38740 VDD.n10032 VDD.n10031 0.04025
R38741 VDD.n10032 VDD.n9237 0.04025
R38742 VDD.n10036 VDD.n9237 0.04025
R38743 VDD.n10037 VDD.n10036 0.04025
R38744 VDD.n10038 VDD.n10037 0.04025
R38745 VDD.n10038 VDD.n9235 0.04025
R38746 VDD.n10042 VDD.n9235 0.04025
R38747 VDD.n10043 VDD.n10042 0.04025
R38748 VDD.n10044 VDD.n10043 0.04025
R38749 VDD.n10044 VDD.n9233 0.04025
R38750 VDD.n10048 VDD.n9233 0.04025
R38751 VDD.n10049 VDD.n10048 0.04025
R38752 VDD.n10050 VDD.n10049 0.04025
R38753 VDD.n10050 VDD.n9231 0.04025
R38754 VDD.n10054 VDD.n9231 0.04025
R38755 VDD.n10055 VDD.n10054 0.04025
R38756 VDD.n10056 VDD.n10055 0.04025
R38757 VDD.n10056 VDD.n9229 0.04025
R38758 VDD.n10060 VDD.n9229 0.04025
R38759 VDD.n10061 VDD.n10060 0.04025
R38760 VDD.n10062 VDD.n10061 0.04025
R38761 VDD.n10062 VDD.n9227 0.04025
R38762 VDD.n10066 VDD.n9227 0.04025
R38763 VDD.n10067 VDD.n10066 0.04025
R38764 VDD.n10068 VDD.n10067 0.04025
R38765 VDD.n10068 VDD.n9225 0.04025
R38766 VDD.n10072 VDD.n9225 0.04025
R38767 VDD.n10073 VDD.n10072 0.04025
R38768 VDD.n10074 VDD.n10073 0.04025
R38769 VDD.n10074 VDD.n9223 0.04025
R38770 VDD.n10078 VDD.n9223 0.04025
R38771 VDD.n10079 VDD.n10078 0.04025
R38772 VDD.n10080 VDD.n10079 0.04025
R38773 VDD.n10080 VDD.n9221 0.04025
R38774 VDD.n10084 VDD.n9221 0.04025
R38775 VDD.n10085 VDD.n10084 0.04025
R38776 VDD.n10086 VDD.n10085 0.04025
R38777 VDD.n10086 VDD.n9219 0.04025
R38778 VDD.n10090 VDD.n9219 0.04025
R38779 VDD.n10091 VDD.n10090 0.04025
R38780 VDD.n10092 VDD.n10091 0.04025
R38781 VDD.n10092 VDD.n9217 0.04025
R38782 VDD.n10096 VDD.n9217 0.04025
R38783 VDD.n10097 VDD.n10096 0.04025
R38784 VDD.n10098 VDD.n10097 0.04025
R38785 VDD.n10098 VDD.n9215 0.04025
R38786 VDD.n10102 VDD.n9215 0.04025
R38787 VDD.n4904 VDD.n4903 0.04025
R38788 VDD.n4903 VDD.n4698 0.04025
R38789 VDD.n4899 VDD.n4698 0.04025
R38790 VDD.n4899 VDD.n4898 0.04025
R38791 VDD.n4898 VDD.n4897 0.04025
R38792 VDD.n4897 VDD.n4700 0.04025
R38793 VDD.n4893 VDD.n4700 0.04025
R38794 VDD.n4893 VDD.n4892 0.04025
R38795 VDD.n4892 VDD.n4891 0.04025
R38796 VDD.n4891 VDD.n4702 0.04025
R38797 VDD.n4887 VDD.n4702 0.04025
R38798 VDD.n4887 VDD.n4886 0.04025
R38799 VDD.n4886 VDD.n4885 0.04025
R38800 VDD.n4885 VDD.n4704 0.04025
R38801 VDD.n4881 VDD.n4704 0.04025
R38802 VDD.n4881 VDD.n4880 0.04025
R38803 VDD.n4880 VDD.n4879 0.04025
R38804 VDD.n4879 VDD.n4706 0.04025
R38805 VDD.n4875 VDD.n4706 0.04025
R38806 VDD.n4875 VDD.n4874 0.04025
R38807 VDD.n4874 VDD.n4873 0.04025
R38808 VDD.n4873 VDD.n4708 0.04025
R38809 VDD.n4869 VDD.n4708 0.04025
R38810 VDD.n4869 VDD.n4868 0.04025
R38811 VDD.n4868 VDD.n4867 0.04025
R38812 VDD.n4867 VDD.n4710 0.04025
R38813 VDD.n4863 VDD.n4710 0.04025
R38814 VDD.n4863 VDD.n4862 0.04025
R38815 VDD.n4862 VDD.n4861 0.04025
R38816 VDD.n4861 VDD.n4712 0.04025
R38817 VDD.n4857 VDD.n4712 0.04025
R38818 VDD.n4857 VDD.n4856 0.04025
R38819 VDD.n4856 VDD.n4855 0.04025
R38820 VDD.n4855 VDD.n4714 0.04025
R38821 VDD.n4851 VDD.n4714 0.04025
R38822 VDD.n4851 VDD.n4850 0.04025
R38823 VDD.n4850 VDD.n4849 0.04025
R38824 VDD.n4849 VDD.n4716 0.04025
R38825 VDD.n4845 VDD.n4716 0.04025
R38826 VDD.n4845 VDD.n4844 0.04025
R38827 VDD.n4844 VDD.n4843 0.04025
R38828 VDD.n4843 VDD.n4718 0.04025
R38829 VDD.n4839 VDD.n4718 0.04025
R38830 VDD.n4839 VDD.n4838 0.04025
R38831 VDD.n4838 VDD.n4837 0.04025
R38832 VDD.n4837 VDD.n4720 0.04025
R38833 VDD.n4833 VDD.n4720 0.04025
R38834 VDD.n4833 VDD.n4832 0.04025
R38835 VDD.n4832 VDD.n4831 0.04025
R38836 VDD.n4831 VDD.n4722 0.04025
R38837 VDD.n4827 VDD.n4722 0.04025
R38838 VDD.n4827 VDD.n4826 0.04025
R38839 VDD.n4826 VDD.n4825 0.04025
R38840 VDD.n4825 VDD.n4724 0.04025
R38841 VDD.n4821 VDD.n4724 0.04025
R38842 VDD.n4821 VDD.n4820 0.04025
R38843 VDD.n4820 VDD.n4819 0.04025
R38844 VDD.n4819 VDD.n4726 0.04025
R38845 VDD.n4815 VDD.n4726 0.04025
R38846 VDD.n4815 VDD.n4814 0.04025
R38847 VDD.n4814 VDD.n4813 0.04025
R38848 VDD.n4813 VDD.n4728 0.04025
R38849 VDD.n4809 VDD.n4728 0.04025
R38850 VDD.n4809 VDD.n4808 0.04025
R38851 VDD.n4808 VDD.n4807 0.04025
R38852 VDD.n4807 VDD.n4730 0.04025
R38853 VDD.n4803 VDD.n4730 0.04025
R38854 VDD.n4803 VDD.n4802 0.04025
R38855 VDD.n4802 VDD.n4801 0.04025
R38856 VDD.n4801 VDD.n4732 0.04025
R38857 VDD.n4797 VDD.n4732 0.04025
R38858 VDD.n4797 VDD.n4796 0.04025
R38859 VDD.n4796 VDD.n4795 0.04025
R38860 VDD.n4795 VDD.n4734 0.04025
R38861 VDD.n4791 VDD.n4734 0.04025
R38862 VDD.n4791 VDD.n4790 0.04025
R38863 VDD.n4790 VDD.n4789 0.04025
R38864 VDD.n4789 VDD.n4736 0.04025
R38865 VDD.n4785 VDD.n4736 0.04025
R38866 VDD.n4785 VDD.n4784 0.04025
R38867 VDD.n4784 VDD.n4783 0.04025
R38868 VDD.n4783 VDD.n4738 0.04025
R38869 VDD.n4779 VDD.n4738 0.04025
R38870 VDD.n4779 VDD.n4778 0.04025
R38871 VDD.n4778 VDD.n4777 0.04025
R38872 VDD.n4777 VDD.n4740 0.04025
R38873 VDD.n4773 VDD.n4740 0.04025
R38874 VDD.n4773 VDD.n4772 0.04025
R38875 VDD.n4772 VDD.n4771 0.04025
R38876 VDD.n4771 VDD.n4742 0.04025
R38877 VDD.n4767 VDD.n4742 0.04025
R38878 VDD.n4767 VDD.n4766 0.04025
R38879 VDD.n4766 VDD.n4765 0.04025
R38880 VDD.n4765 VDD.n4744 0.04025
R38881 VDD.n4761 VDD.n4744 0.04025
R38882 VDD.n4761 VDD.n4760 0.04025
R38883 VDD.n4760 VDD.n4759 0.04025
R38884 VDD.n4759 VDD.n4746 0.04025
R38885 VDD.n4755 VDD.n4746 0.04025
R38886 VDD.n4755 VDD.n4754 0.04025
R38887 VDD.n4754 VDD.n4753 0.04025
R38888 VDD.n4753 VDD.n4748 0.04025
R38889 VDD.n4749 VDD.n4748 0.04025
R38890 VDD.n4749 VDD.n2244 0.04025
R38891 VDD.n7819 VDD.n2244 0.04025
R38892 VDD.n7819 VDD.n7818 0.04025
R38893 VDD.n7818 VDD.n7817 0.04025
R38894 VDD.n7817 VDD.n2245 0.04025
R38895 VDD.n7813 VDD.n2245 0.04025
R38896 VDD.n7813 VDD.n7812 0.04025
R38897 VDD.n7812 VDD.n7811 0.04025
R38898 VDD.n7811 VDD.n2247 0.04025
R38899 VDD.n7806 VDD.n2247 0.04025
R38900 VDD.n7806 VDD.n7805 0.04025
R38901 VDD.n7805 VDD.n7804 0.04025
R38902 VDD.n7804 VDD.n2249 0.04025
R38903 VDD.n7800 VDD.n2249 0.04025
R38904 VDD.n7800 VDD.n7799 0.04025
R38905 VDD.n7799 VDD.n2251 0.04025
R38906 VDD.n7795 VDD.n2251 0.04025
R38907 VDD.n7795 VDD.n7794 0.04025
R38908 VDD.n7794 VDD.n2253 0.04025
R38909 VDD.n7790 VDD.n2253 0.04025
R38910 VDD.n7790 VDD.n7789 0.04025
R38911 VDD.n7789 VDD.n7788 0.04025
R38912 VDD.n7788 VDD.n2255 0.04025
R38913 VDD.n7784 VDD.n2255 0.04025
R38914 VDD.n7784 VDD.n7783 0.04025
R38915 VDD.n7783 VDD.n7782 0.04025
R38916 VDD.n7782 VDD.n2257 0.04025
R38917 VDD.n7777 VDD.n2257 0.04025
R38918 VDD.n7777 VDD.n7776 0.04025
R38919 VDD.n7776 VDD.n7775 0.04025
R38920 VDD.n7775 VDD.n2259 0.04025
R38921 VDD.n7771 VDD.n2259 0.04025
R38922 VDD.n7771 VDD.n7770 0.04025
R38923 VDD.n7770 VDD.n7769 0.04025
R38924 VDD.n7769 VDD.n2262 0.04025
R38925 VDD.n7765 VDD.n2262 0.04025
R38926 VDD.n7765 VDD.n7764 0.04025
R38927 VDD.n7764 VDD.n7763 0.04025
R38928 VDD.n7763 VDD.n2264 0.04025
R38929 VDD.n7758 VDD.n2264 0.04025
R38930 VDD.n7758 VDD.n7757 0.04025
R38931 VDD.n7757 VDD.n7756 0.04025
R38932 VDD.n7756 VDD.n2267 0.04025
R38933 VDD.n7752 VDD.n2267 0.04025
R38934 VDD.n7752 VDD.n7751 0.04025
R38935 VDD.n7751 VDD.n7750 0.04025
R38936 VDD.n7750 VDD.n2269 0.04025
R38937 VDD.n7746 VDD.n2269 0.04025
R38938 VDD.n7746 VDD.n7745 0.04025
R38939 VDD.n7745 VDD.n2271 0.04025
R38940 VDD.n7741 VDD.n2271 0.04025
R38941 VDD.n7741 VDD.n7740 0.04025
R38942 VDD.n7740 VDD.n2273 0.04025
R38943 VDD.n7736 VDD.n2273 0.04025
R38944 VDD.n7736 VDD.n7735 0.04025
R38945 VDD.n7735 VDD.n7734 0.04025
R38946 VDD.n7734 VDD.n2275 0.04025
R38947 VDD.n7730 VDD.n2275 0.04025
R38948 VDD.n7730 VDD.n7729 0.04025
R38949 VDD.n7729 VDD.n7728 0.04025
R38950 VDD.n7728 VDD.n2277 0.04025
R38951 VDD.n7723 VDD.n2277 0.04025
R38952 VDD.n7723 VDD.n7722 0.04025
R38953 VDD.n7722 VDD.n7721 0.04025
R38954 VDD.n7721 VDD.n2279 0.04025
R38955 VDD.n7716 VDD.n2279 0.04025
R38956 VDD.n7716 VDD.n7715 0.04025
R38957 VDD.n7715 VDD.n7714 0.04025
R38958 VDD.n7714 VDD.n2281 0.04025
R38959 VDD.n7710 VDD.n2281 0.04025
R38960 VDD.n7710 VDD.n7709 0.04025
R38961 VDD.n7709 VDD.n2284 0.04025
R38962 VDD.n7705 VDD.n2284 0.04025
R38963 VDD.n7705 VDD.n7704 0.04025
R38964 VDD.n7704 VDD.n7703 0.04025
R38965 VDD.n7703 VDD.n2286 0.04025
R38966 VDD.n7698 VDD.n2286 0.04025
R38967 VDD.n7698 VDD.n7697 0.04025
R38968 VDD.n7697 VDD.n7696 0.04025
R38969 VDD.n7696 VDD.n2288 0.04025
R38970 VDD.n7692 VDD.n2288 0.04025
R38971 VDD.n7692 VDD.n7691 0.04025
R38972 VDD.n7691 VDD.n7690 0.04025
R38973 VDD.n7690 VDD.n2290 0.04025
R38974 VDD.n7686 VDD.n2290 0.04025
R38975 VDD.n7686 VDD.n7685 0.04025
R38976 VDD.n7685 VDD.n2293 0.04025
R38977 VDD.n7680 VDD.n2293 0.04025
R38978 VDD.n7680 VDD.n7679 0.04025
R38979 VDD.n7679 VDD.n7678 0.04025
R38980 VDD.n7678 VDD.n7179 0.04025
R38981 VDD.n7674 VDD.n7179 0.04025
R38982 VDD.n7674 VDD.n7673 0.04025
R38983 VDD.n7673 VDD.n7672 0.04025
R38984 VDD.n7672 VDD.n7181 0.04025
R38985 VDD.n7668 VDD.n7181 0.04025
R38986 VDD.n7668 VDD.n7667 0.04025
R38987 VDD.n7667 VDD.n7666 0.04025
R38988 VDD.n7666 VDD.n7183 0.04025
R38989 VDD.n7662 VDD.n7183 0.04025
R38990 VDD.n7662 VDD.n7661 0.04025
R38991 VDD.n7661 VDD.n7660 0.04025
R38992 VDD.n7660 VDD.n7185 0.04025
R38993 VDD.n7656 VDD.n7185 0.04025
R38994 VDD.n7656 VDD.n7655 0.04025
R38995 VDD.n7655 VDD.n7654 0.04025
R38996 VDD.n7654 VDD.n7187 0.04025
R38997 VDD.n7650 VDD.n7187 0.04025
R38998 VDD.n7650 VDD.n7649 0.04025
R38999 VDD.n7649 VDD.n7648 0.04025
R39000 VDD.n7648 VDD.n7189 0.04025
R39001 VDD.n7644 VDD.n7189 0.04025
R39002 VDD.n7644 VDD.n7643 0.04025
R39003 VDD.n7643 VDD.n7642 0.04025
R39004 VDD.n7642 VDD.n7191 0.04025
R39005 VDD.n7638 VDD.n7191 0.04025
R39006 VDD.n7638 VDD.n7637 0.04025
R39007 VDD.n7637 VDD.n7636 0.04025
R39008 VDD.n7636 VDD.n7193 0.04025
R39009 VDD.n7632 VDD.n7193 0.04025
R39010 VDD.n7632 VDD.n7631 0.04025
R39011 VDD.n7631 VDD.n7630 0.04025
R39012 VDD.n7630 VDD.n7195 0.04025
R39013 VDD.n7626 VDD.n7195 0.04025
R39014 VDD.n7626 VDD.n7625 0.04025
R39015 VDD.n7625 VDD.n7624 0.04025
R39016 VDD.n7624 VDD.n7197 0.04025
R39017 VDD.n7620 VDD.n7197 0.04025
R39018 VDD.n7620 VDD.n7619 0.04025
R39019 VDD.n7619 VDD.n7618 0.04025
R39020 VDD.n7618 VDD.n7199 0.04025
R39021 VDD.n7614 VDD.n7199 0.04025
R39022 VDD.n7614 VDD.n7613 0.04025
R39023 VDD.n7613 VDD.n7612 0.04025
R39024 VDD.n7612 VDD.n7201 0.04025
R39025 VDD.n7608 VDD.n7201 0.04025
R39026 VDD.n7608 VDD.n7607 0.04025
R39027 VDD.n7607 VDD.n7606 0.04025
R39028 VDD.n7606 VDD.n7203 0.04025
R39029 VDD.n7602 VDD.n7203 0.04025
R39030 VDD.n7602 VDD.n7601 0.04025
R39031 VDD.n7601 VDD.n7600 0.04025
R39032 VDD.n7600 VDD.n7205 0.04025
R39033 VDD.n7596 VDD.n7205 0.04025
R39034 VDD.n7596 VDD.n7595 0.04025
R39035 VDD.n7595 VDD.n7594 0.04025
R39036 VDD.n7594 VDD.n7207 0.04025
R39037 VDD.n7590 VDD.n7207 0.04025
R39038 VDD.n7590 VDD.n7589 0.04025
R39039 VDD.n7589 VDD.n7588 0.04025
R39040 VDD.n7588 VDD.n7209 0.04025
R39041 VDD.n7584 VDD.n7209 0.04025
R39042 VDD.n7584 VDD.n7583 0.04025
R39043 VDD.n7583 VDD.n7582 0.04025
R39044 VDD.n7582 VDD.n7211 0.04025
R39045 VDD.n7578 VDD.n7211 0.04025
R39046 VDD.n7578 VDD.n7577 0.04025
R39047 VDD.n7577 VDD.n7576 0.04025
R39048 VDD.n7576 VDD.n7213 0.04025
R39049 VDD.n7572 VDD.n7213 0.04025
R39050 VDD.n7572 VDD.n7571 0.04025
R39051 VDD.n7571 VDD.n7570 0.04025
R39052 VDD.n7570 VDD.n7215 0.04025
R39053 VDD.n7566 VDD.n7215 0.04025
R39054 VDD.n7566 VDD.n7565 0.04025
R39055 VDD.n7565 VDD.n7564 0.04025
R39056 VDD.n7564 VDD.n7217 0.04025
R39057 VDD.n7560 VDD.n7217 0.04025
R39058 VDD.n7560 VDD.n7559 0.04025
R39059 VDD.n7559 VDD.n7558 0.04025
R39060 VDD.n7558 VDD.n7219 0.04025
R39061 VDD.n7554 VDD.n7219 0.04025
R39062 VDD.n7554 VDD.n7553 0.04025
R39063 VDD.n7553 VDD.n7552 0.04025
R39064 VDD.n7552 VDD.n7221 0.04025
R39065 VDD.n7548 VDD.n7221 0.04025
R39066 VDD.n7548 VDD.n7547 0.04025
R39067 VDD.n7547 VDD.n7546 0.04025
R39068 VDD.n7546 VDD.n7223 0.04025
R39069 VDD.n7542 VDD.n7223 0.04025
R39070 VDD.n7542 VDD.n7541 0.04025
R39071 VDD.n7541 VDD.n7540 0.04025
R39072 VDD.n7540 VDD.n7225 0.04025
R39073 VDD.n7536 VDD.n7225 0.04025
R39074 VDD.n7536 VDD.n7535 0.04025
R39075 VDD.n7535 VDD.n7534 0.04025
R39076 VDD.n7534 VDD.n7227 0.04025
R39077 VDD.n7530 VDD.n7227 0.04025
R39078 VDD.n7530 VDD.n7529 0.04025
R39079 VDD.n7529 VDD.n7528 0.04025
R39080 VDD.n7528 VDD.n7229 0.04025
R39081 VDD.n7524 VDD.n7229 0.04025
R39082 VDD.n7524 VDD.n7523 0.04025
R39083 VDD.n7523 VDD.n7522 0.04025
R39084 VDD.n7522 VDD.n7231 0.04025
R39085 VDD.n7518 VDD.n7231 0.04025
R39086 VDD.n7518 VDD.n7517 0.04025
R39087 VDD.n7517 VDD.n7516 0.04025
R39088 VDD.n7516 VDD.n7233 0.04025
R39089 VDD.n7512 VDD.n7233 0.04025
R39090 VDD.n7512 VDD.n7511 0.04025
R39091 VDD.n7511 VDD.n7510 0.04025
R39092 VDD.n7510 VDD.n7235 0.04025
R39093 VDD.n7506 VDD.n7235 0.04025
R39094 VDD.n7506 VDD.n7505 0.04025
R39095 VDD.n7505 VDD.n7504 0.04025
R39096 VDD.n7504 VDD.n7237 0.04025
R39097 VDD.n7500 VDD.n7237 0.04025
R39098 VDD.n7500 VDD.n7499 0.04025
R39099 VDD.n7499 VDD.n7498 0.04025
R39100 VDD.n7498 VDD.n7239 0.04025
R39101 VDD.n7494 VDD.n7239 0.04025
R39102 VDD.n7494 VDD.n7493 0.04025
R39103 VDD.n7493 VDD.n7492 0.04025
R39104 VDD.n7492 VDD.n7241 0.04025
R39105 VDD.n7488 VDD.n7241 0.04025
R39106 VDD.n7488 VDD.n7487 0.04025
R39107 VDD.n7487 VDD.n7486 0.04025
R39108 VDD.n7486 VDD.n7243 0.04025
R39109 VDD.n7482 VDD.n7243 0.04025
R39110 VDD.n7482 VDD.n7481 0.04025
R39111 VDD.n7481 VDD.n7480 0.04025
R39112 VDD.n7480 VDD.n7245 0.04025
R39113 VDD.n7476 VDD.n7245 0.04025
R39114 VDD.n7476 VDD.n7475 0.04025
R39115 VDD.n7475 VDD.n7474 0.04025
R39116 VDD.n7474 VDD.n7247 0.04025
R39117 VDD.n7470 VDD.n7247 0.04025
R39118 VDD.n7470 VDD.n7469 0.04025
R39119 VDD.n7469 VDD.n7468 0.04025
R39120 VDD.n7468 VDD.n7249 0.04025
R39121 VDD.n7464 VDD.n7249 0.04025
R39122 VDD.n7464 VDD.n7463 0.04025
R39123 VDD.n7463 VDD.n7462 0.04025
R39124 VDD.n7462 VDD.n7251 0.04025
R39125 VDD.n7458 VDD.n7251 0.04025
R39126 VDD.n7458 VDD.n7457 0.04025
R39127 VDD.n7457 VDD.n7456 0.04025
R39128 VDD.n7456 VDD.n7253 0.04025
R39129 VDD.n7452 VDD.n7253 0.04025
R39130 VDD.n7452 VDD.n7451 0.04025
R39131 VDD.n7451 VDD.n7450 0.04025
R39132 VDD.n7450 VDD.n7255 0.04025
R39133 VDD.n7446 VDD.n7255 0.04025
R39134 VDD.n7446 VDD.n7445 0.04025
R39135 VDD.n7445 VDD.n7444 0.04025
R39136 VDD.n7444 VDD.n7257 0.04025
R39137 VDD.n7440 VDD.n7257 0.04025
R39138 VDD.n7440 VDD.n7439 0.04025
R39139 VDD.n7439 VDD.n7438 0.04025
R39140 VDD.n7438 VDD.n7259 0.04025
R39141 VDD.n7434 VDD.n7259 0.04025
R39142 VDD.n7434 VDD.n7433 0.04025
R39143 VDD.n7433 VDD.n7432 0.04025
R39144 VDD.n7432 VDD.n7261 0.04025
R39145 VDD.n7428 VDD.n7261 0.04025
R39146 VDD.n7428 VDD.n7427 0.04025
R39147 VDD.n7427 VDD.n7426 0.04025
R39148 VDD.n7426 VDD.n7263 0.04025
R39149 VDD.n7422 VDD.n7263 0.04025
R39150 VDD.n7422 VDD.n7421 0.04025
R39151 VDD.n7421 VDD.n7420 0.04025
R39152 VDD.n7420 VDD.n7265 0.04025
R39153 VDD.n7416 VDD.n7265 0.04025
R39154 VDD.n7416 VDD.n7415 0.04025
R39155 VDD.n7415 VDD.n7414 0.04025
R39156 VDD.n7414 VDD.n7267 0.04025
R39157 VDD.n7410 VDD.n7267 0.04025
R39158 VDD.n7410 VDD.n7409 0.04025
R39159 VDD.n7409 VDD.n7408 0.04025
R39160 VDD.n7408 VDD.n7269 0.04025
R39161 VDD.n7404 VDD.n7269 0.04025
R39162 VDD.n7404 VDD.n7403 0.04025
R39163 VDD.n7403 VDD.n7402 0.04025
R39164 VDD.n7402 VDD.n7271 0.04025
R39165 VDD.n7398 VDD.n7271 0.04025
R39166 VDD.n7398 VDD.n7397 0.04025
R39167 VDD.n7397 VDD.n7396 0.04025
R39168 VDD.n7396 VDD.n7273 0.04025
R39169 VDD.n7392 VDD.n7273 0.04025
R39170 VDD.n7392 VDD.n7391 0.04025
R39171 VDD.n7391 VDD.n7390 0.04025
R39172 VDD.n7390 VDD.n7275 0.04025
R39173 VDD.n7386 VDD.n7275 0.04025
R39174 VDD.n7386 VDD.n7385 0.04025
R39175 VDD.n7385 VDD.n7384 0.04025
R39176 VDD.n7384 VDD.n7277 0.04025
R39177 VDD.n7380 VDD.n7277 0.04025
R39178 VDD.n7380 VDD.n7379 0.04025
R39179 VDD.n7379 VDD.n7378 0.04025
R39180 VDD.n7378 VDD.n7279 0.04025
R39181 VDD.n7374 VDD.n7279 0.04025
R39182 VDD.n7374 VDD.n7373 0.04025
R39183 VDD.n7373 VDD.n7372 0.04025
R39184 VDD.n7372 VDD.n7281 0.04025
R39185 VDD.n7368 VDD.n7281 0.04025
R39186 VDD.n7368 VDD.n7367 0.04025
R39187 VDD.n7367 VDD.n7366 0.04025
R39188 VDD.n7366 VDD.n7283 0.04025
R39189 VDD.n7362 VDD.n7283 0.04025
R39190 VDD.n7362 VDD.n7361 0.04025
R39191 VDD.n7361 VDD.n7360 0.04025
R39192 VDD.n7360 VDD.n7285 0.04025
R39193 VDD.n7356 VDD.n7285 0.04025
R39194 VDD.n7356 VDD.n7355 0.04025
R39195 VDD.n7355 VDD.n7354 0.04025
R39196 VDD.n7354 VDD.n7287 0.04025
R39197 VDD.n7350 VDD.n7287 0.04025
R39198 VDD.n7350 VDD.n7349 0.04025
R39199 VDD.n7349 VDD.n7348 0.04025
R39200 VDD.n7348 VDD.n7289 0.04025
R39201 VDD.n7344 VDD.n7289 0.04025
R39202 VDD.n7344 VDD.n7343 0.04025
R39203 VDD.n7343 VDD.n7342 0.04025
R39204 VDD.n7342 VDD.n7291 0.04025
R39205 VDD.n7338 VDD.n7291 0.04025
R39206 VDD.n7338 VDD.n7337 0.04025
R39207 VDD.n7337 VDD.n7336 0.04025
R39208 VDD.n7336 VDD.n7293 0.04025
R39209 VDD.n7332 VDD.n7293 0.04025
R39210 VDD.n7332 VDD.n7331 0.04025
R39211 VDD.n7331 VDD.n7330 0.04025
R39212 VDD.n7330 VDD.n7295 0.04025
R39213 VDD.n7326 VDD.n7295 0.04025
R39214 VDD.n7326 VDD.n7325 0.04025
R39215 VDD.n7325 VDD.n7324 0.04025
R39216 VDD.n7324 VDD.n7297 0.04025
R39217 VDD.n7320 VDD.n7297 0.04025
R39218 VDD.n7320 VDD.n7319 0.04025
R39219 VDD.n7319 VDD.n7318 0.04025
R39220 VDD.n7318 VDD.n7299 0.04025
R39221 VDD.n7314 VDD.n7299 0.04025
R39222 VDD.n7314 VDD.n7313 0.04025
R39223 VDD.n7313 VDD.n7312 0.04025
R39224 VDD.n7312 VDD.n7301 0.04025
R39225 VDD.n7308 VDD.n7301 0.04025
R39226 VDD.n7308 VDD.n7307 0.04025
R39227 VDD.n7307 VDD.n7306 0.04025
R39228 VDD.n7306 VDD.n7303 0.04025
R39229 VDD.n7303 VDD.n2087 0.04025
R39230 VDD.n8169 VDD.n2087 0.04025
R39231 VDD.n8170 VDD.n8169 0.04025
R39232 VDD.n8171 VDD.n8170 0.04025
R39233 VDD.n8171 VDD.n2085 0.04025
R39234 VDD.n8176 VDD.n2085 0.04025
R39235 VDD.n8177 VDD.n8176 0.04025
R39236 VDD.n8178 VDD.n8177 0.04025
R39237 VDD.n8178 VDD.n2083 0.04025
R39238 VDD.n8184 VDD.n2083 0.04025
R39239 VDD.n8185 VDD.n8184 0.04025
R39240 VDD.n8186 VDD.n8185 0.04025
R39241 VDD.n8186 VDD.n2081 0.04025
R39242 VDD.n8191 VDD.n2081 0.04025
R39243 VDD.n8192 VDD.n8191 0.04025
R39244 VDD.n8193 VDD.n8192 0.04025
R39245 VDD.n8193 VDD.n2079 0.04025
R39246 VDD.n8197 VDD.n2079 0.04025
R39247 VDD.n8198 VDD.n8197 0.04025
R39248 VDD.n8198 VDD.n2077 0.04025
R39249 VDD.n8204 VDD.n2077 0.04025
R39250 VDD.n8205 VDD.n8204 0.04025
R39251 VDD.n8206 VDD.n8205 0.04025
R39252 VDD.n8206 VDD.n2075 0.04025
R39253 VDD.n8210 VDD.n2075 0.04025
R39254 VDD.n8211 VDD.n8210 0.04025
R39255 VDD.n8211 VDD.n2073 0.04025
R39256 VDD.n8217 VDD.n2073 0.04025
R39257 VDD.n8218 VDD.n8217 0.04025
R39258 VDD.n8219 VDD.n8218 0.04025
R39259 VDD.n8219 VDD.n2071 0.04025
R39260 VDD.n8224 VDD.n2071 0.04025
R39261 VDD.n8225 VDD.n8224 0.04025
R39262 VDD.n8226 VDD.n8225 0.04025
R39263 VDD.n8226 VDD.n2069 0.04025
R39264 VDD.n8231 VDD.n2069 0.04025
R39265 VDD.n8232 VDD.n8231 0.04025
R39266 VDD.n8233 VDD.n8232 0.04025
R39267 VDD.n8233 VDD.n2067 0.04025
R39268 VDD.n8239 VDD.n2067 0.04025
R39269 VDD.n8240 VDD.n8239 0.04025
R39270 VDD.n8241 VDD.n8240 0.04025
R39271 VDD.n8241 VDD.n2065 0.04025
R39272 VDD.n8245 VDD.n2065 0.04025
R39273 VDD.n8246 VDD.n8245 0.04025
R39274 VDD.n8246 VDD.n2063 0.04025
R39275 VDD.n8252 VDD.n2063 0.04025
R39276 VDD.n8253 VDD.n8252 0.04025
R39277 VDD.n10764 VDD.n8253 0.04025
R39278 VDD.n10764 VDD.n10763 0.04025
R39279 VDD.n10763 VDD.n10762 0.04025
R39280 VDD.n10762 VDD.n8254 0.04025
R39281 VDD.n10758 VDD.n8254 0.04025
R39282 VDD.n10758 VDD.n10757 0.04025
R39283 VDD.n10757 VDD.n10756 0.04025
R39284 VDD.n10756 VDD.n8256 0.04025
R39285 VDD.n10752 VDD.n8256 0.04025
R39286 VDD.n10752 VDD.n10751 0.04025
R39287 VDD.n10751 VDD.n10750 0.04025
R39288 VDD.n10750 VDD.n8258 0.04025
R39289 VDD.n10746 VDD.n8258 0.04025
R39290 VDD.n10746 VDD.n10745 0.04025
R39291 VDD.n10745 VDD.n10744 0.04025
R39292 VDD.n10744 VDD.n8260 0.04025
R39293 VDD.n10740 VDD.n8260 0.04025
R39294 VDD.n10740 VDD.n10739 0.04025
R39295 VDD.n10739 VDD.n10738 0.04025
R39296 VDD.n10738 VDD.n8262 0.04025
R39297 VDD.n10734 VDD.n8262 0.04025
R39298 VDD.n10734 VDD.n10733 0.04025
R39299 VDD.n10733 VDD.n10732 0.04025
R39300 VDD.n10732 VDD.n8264 0.04025
R39301 VDD.n10728 VDD.n8264 0.04025
R39302 VDD.n10728 VDD.n10727 0.04025
R39303 VDD.n10727 VDD.n10726 0.04025
R39304 VDD.n10726 VDD.n8266 0.04025
R39305 VDD.n10722 VDD.n8266 0.04025
R39306 VDD.n10722 VDD.n10721 0.04025
R39307 VDD.n10721 VDD.n10720 0.04025
R39308 VDD.n10720 VDD.n8268 0.04025
R39309 VDD.n10716 VDD.n8268 0.04025
R39310 VDD.n10716 VDD.n10715 0.04025
R39311 VDD.n10715 VDD.n10714 0.04025
R39312 VDD.n10714 VDD.n8270 0.04025
R39313 VDD.n10710 VDD.n8270 0.04025
R39314 VDD.n10710 VDD.n10709 0.04025
R39315 VDD.n10709 VDD.n10708 0.04025
R39316 VDD.n10708 VDD.n8272 0.04025
R39317 VDD.n10704 VDD.n8272 0.04025
R39318 VDD.n10704 VDD.n10703 0.04025
R39319 VDD.n10703 VDD.n10702 0.04025
R39320 VDD.n10702 VDD.n8274 0.04025
R39321 VDD.n10698 VDD.n8274 0.04025
R39322 VDD.n10698 VDD.n10697 0.04025
R39323 VDD.n10697 VDD.n10696 0.04025
R39324 VDD.n10696 VDD.n8276 0.04025
R39325 VDD.n10692 VDD.n8276 0.04025
R39326 VDD.n10692 VDD.n10691 0.04025
R39327 VDD.n10691 VDD.n10690 0.04025
R39328 VDD.n10690 VDD.n8278 0.04025
R39329 VDD.n10686 VDD.n8278 0.04025
R39330 VDD.n10686 VDD.n10685 0.04025
R39331 VDD.n10685 VDD.n10684 0.04025
R39332 VDD.n10684 VDD.n8280 0.04025
R39333 VDD.n10680 VDD.n8280 0.04025
R39334 VDD.n10680 VDD.n10679 0.04025
R39335 VDD.n10679 VDD.n10678 0.04025
R39336 VDD.n10678 VDD.n8282 0.04025
R39337 VDD.n10674 VDD.n8282 0.04025
R39338 VDD.n10674 VDD.n10673 0.04025
R39339 VDD.n10673 VDD.n10672 0.04025
R39340 VDD.n10672 VDD.n8284 0.04025
R39341 VDD.n10668 VDD.n8284 0.04025
R39342 VDD.n10668 VDD.n10667 0.04025
R39343 VDD.n10667 VDD.n10666 0.04025
R39344 VDD.n10666 VDD.n8286 0.04025
R39345 VDD.n10662 VDD.n8286 0.04025
R39346 VDD.n10662 VDD.n10661 0.04025
R39347 VDD.n10661 VDD.n10660 0.04025
R39348 VDD.n10660 VDD.n8288 0.04025
R39349 VDD.n10656 VDD.n8288 0.04025
R39350 VDD.n10656 VDD.n10655 0.04025
R39351 VDD.n10655 VDD.n10654 0.04025
R39352 VDD.n10654 VDD.n8290 0.04025
R39353 VDD.n10650 VDD.n8290 0.04025
R39354 VDD.n10650 VDD.n10649 0.04025
R39355 VDD.n10649 VDD.n10648 0.04025
R39356 VDD.n10648 VDD.n8292 0.04025
R39357 VDD.n10644 VDD.n8292 0.04025
R39358 VDD.n10644 VDD.n10643 0.04025
R39359 VDD.n10643 VDD.n10642 0.04025
R39360 VDD.n10642 VDD.n8294 0.04025
R39361 VDD.n10638 VDD.n8294 0.04025
R39362 VDD.n10638 VDD.n10637 0.04025
R39363 VDD.n10637 VDD.n10636 0.04025
R39364 VDD.n10636 VDD.n8296 0.04025
R39365 VDD.n10632 VDD.n8296 0.04025
R39366 VDD.n10632 VDD.n10631 0.04025
R39367 VDD.n10631 VDD.n10630 0.04025
R39368 VDD.n10630 VDD.n8298 0.04025
R39369 VDD.n10626 VDD.n8298 0.04025
R39370 VDD.n10626 VDD.n10625 0.04025
R39371 VDD.n10625 VDD.n10624 0.04025
R39372 VDD.n10624 VDD.n8300 0.04025
R39373 VDD.n10620 VDD.n8300 0.04025
R39374 VDD.n10620 VDD.n10619 0.04025
R39375 VDD.n10619 VDD.n10618 0.04025
R39376 VDD.n10618 VDD.n8302 0.04025
R39377 VDD.n10614 VDD.n8302 0.04025
R39378 VDD.n10614 VDD.n10613 0.04025
R39379 VDD.n10613 VDD.n10612 0.04025
R39380 VDD.n10612 VDD.n8304 0.04025
R39381 VDD.n10608 VDD.n8304 0.04025
R39382 VDD.n10608 VDD.n10607 0.04025
R39383 VDD.n10607 VDD.n10606 0.04025
R39384 VDD.n10606 VDD.n8306 0.04025
R39385 VDD.n10602 VDD.n8306 0.04025
R39386 VDD.n10602 VDD.n10601 0.04025
R39387 VDD.n10601 VDD.n10600 0.04025
R39388 VDD.n10600 VDD.n8308 0.04025
R39389 VDD.n10596 VDD.n8308 0.04025
R39390 VDD.n10596 VDD.n10595 0.04025
R39391 VDD.n10595 VDD.n10594 0.04025
R39392 VDD.n10594 VDD.n8310 0.04025
R39393 VDD.n10590 VDD.n8310 0.04025
R39394 VDD.n10590 VDD.n10589 0.04025
R39395 VDD.n10589 VDD.n10588 0.04025
R39396 VDD.n10588 VDD.n8312 0.04025
R39397 VDD.n10584 VDD.n8312 0.04025
R39398 VDD.n10584 VDD.n10583 0.04025
R39399 VDD.n10583 VDD.n10582 0.04025
R39400 VDD.n10582 VDD.n8314 0.04025
R39401 VDD.n10578 VDD.n8314 0.04025
R39402 VDD.n10578 VDD.n10577 0.04025
R39403 VDD.n10577 VDD.n10576 0.04025
R39404 VDD.n10576 VDD.n8316 0.04025
R39405 VDD.n10572 VDD.n8316 0.04025
R39406 VDD.n10572 VDD.n10571 0.04025
R39407 VDD.n10571 VDD.n10570 0.04025
R39408 VDD.n10570 VDD.n8318 0.04025
R39409 VDD.n10566 VDD.n8318 0.04025
R39410 VDD.n10566 VDD.n10565 0.04025
R39411 VDD.n10565 VDD.n10564 0.04025
R39412 VDD.n10564 VDD.n8320 0.04025
R39413 VDD.n10560 VDD.n8320 0.04025
R39414 VDD.n10560 VDD.n10559 0.04025
R39415 VDD.n10559 VDD.n10558 0.04025
R39416 VDD.n10558 VDD.n8322 0.04025
R39417 VDD.n10554 VDD.n8322 0.04025
R39418 VDD.n10554 VDD.n10553 0.04025
R39419 VDD.n10553 VDD.n10552 0.04025
R39420 VDD.n10552 VDD.n8324 0.04025
R39421 VDD.n10548 VDD.n8324 0.04025
R39422 VDD.n10548 VDD.n10547 0.04025
R39423 VDD.n10547 VDD.n10546 0.04025
R39424 VDD.n10546 VDD.n8326 0.04025
R39425 VDD.n10542 VDD.n8326 0.04025
R39426 VDD.n10542 VDD.n10541 0.04025
R39427 VDD.n10541 VDD.n10540 0.04025
R39428 VDD.n10540 VDD.n8328 0.04025
R39429 VDD.n10536 VDD.n8328 0.04025
R39430 VDD.n10536 VDD.n10535 0.04025
R39431 VDD.n10535 VDD.n10534 0.04025
R39432 VDD.n10534 VDD.n8330 0.04025
R39433 VDD.n10530 VDD.n8330 0.04025
R39434 VDD.n10530 VDD.n10529 0.04025
R39435 VDD.n10529 VDD.n10528 0.04025
R39436 VDD.n10528 VDD.n8332 0.04025
R39437 VDD.n10524 VDD.n8332 0.04025
R39438 VDD.n10524 VDD.n10523 0.04025
R39439 VDD.n10523 VDD.n10522 0.04025
R39440 VDD.n10522 VDD.n8334 0.04025
R39441 VDD.n10518 VDD.n8334 0.04025
R39442 VDD.n10518 VDD.n10517 0.04025
R39443 VDD.n10517 VDD.n10516 0.04025
R39444 VDD.n10516 VDD.n8336 0.04025
R39445 VDD.n10512 VDD.n8336 0.04025
R39446 VDD.n10512 VDD.n10511 0.04025
R39447 VDD.n10511 VDD.n10510 0.04025
R39448 VDD.n10510 VDD.n8338 0.04025
R39449 VDD.n10506 VDD.n8338 0.04025
R39450 VDD.n10506 VDD.n10505 0.04025
R39451 VDD.n10505 VDD.n10504 0.04025
R39452 VDD.n10504 VDD.n8340 0.04025
R39453 VDD.n10500 VDD.n8340 0.04025
R39454 VDD.n10500 VDD.n10499 0.04025
R39455 VDD.n10499 VDD.n10498 0.04025
R39456 VDD.n10498 VDD.n8342 0.04025
R39457 VDD.n10494 VDD.n8342 0.04025
R39458 VDD.n10494 VDD.n10493 0.04025
R39459 VDD.n10493 VDD.n10492 0.04025
R39460 VDD.n10492 VDD.n8344 0.04025
R39461 VDD.n10488 VDD.n8344 0.04025
R39462 VDD.n10488 VDD.n10487 0.04025
R39463 VDD.n10487 VDD.n10486 0.04025
R39464 VDD.n10486 VDD.n8346 0.04025
R39465 VDD.n10482 VDD.n8346 0.04025
R39466 VDD.n10482 VDD.n10481 0.04025
R39467 VDD.n10481 VDD.n10480 0.04025
R39468 VDD.n10480 VDD.n8348 0.04025
R39469 VDD.n10476 VDD.n8348 0.04025
R39470 VDD.n10476 VDD.n10475 0.04025
R39471 VDD.n10475 VDD.n10474 0.04025
R39472 VDD.n10474 VDD.n8350 0.04025
R39473 VDD.n10470 VDD.n8350 0.04025
R39474 VDD.n10470 VDD.n10469 0.04025
R39475 VDD.n10469 VDD.n10468 0.04025
R39476 VDD.n10468 VDD.n8352 0.04025
R39477 VDD.n10464 VDD.n8352 0.04025
R39478 VDD.n10464 VDD.n10463 0.04025
R39479 VDD.n10463 VDD.n10462 0.04025
R39480 VDD.n10462 VDD.n8354 0.04025
R39481 VDD.n10458 VDD.n8354 0.04025
R39482 VDD.n10458 VDD.n10457 0.04025
R39483 VDD.n10457 VDD.n10456 0.04025
R39484 VDD.n10456 VDD.n8356 0.04025
R39485 VDD.n10452 VDD.n8356 0.04025
R39486 VDD.n10452 VDD.n10451 0.04025
R39487 VDD.n10451 VDD.n10450 0.04025
R39488 VDD.n10450 VDD.n8358 0.04025
R39489 VDD.n10446 VDD.n8358 0.04025
R39490 VDD.n10446 VDD.n10445 0.04025
R39491 VDD.n10445 VDD.n10444 0.04025
R39492 VDD.n10444 VDD.n8360 0.04025
R39493 VDD.n10440 VDD.n8360 0.04025
R39494 VDD.n10440 VDD.n10439 0.04025
R39495 VDD.n10439 VDD.n10438 0.04025
R39496 VDD.n10438 VDD.n8362 0.04025
R39497 VDD.n10434 VDD.n8362 0.04025
R39498 VDD.n10434 VDD.n10433 0.04025
R39499 VDD.n10433 VDD.n10432 0.04025
R39500 VDD.n10432 VDD.n8364 0.04025
R39501 VDD.n10428 VDD.n8364 0.04025
R39502 VDD.n10428 VDD.n10427 0.04025
R39503 VDD.n10427 VDD.n10426 0.04025
R39504 VDD.n10426 VDD.n8366 0.04025
R39505 VDD.n10422 VDD.n8366 0.04025
R39506 VDD.n10422 VDD.n10421 0.04025
R39507 VDD.n10421 VDD.n10420 0.04025
R39508 VDD.n10420 VDD.n8368 0.04025
R39509 VDD.n10416 VDD.n8368 0.04025
R39510 VDD.n10416 VDD.n10415 0.04025
R39511 VDD.n10415 VDD.n10414 0.04025
R39512 VDD.n10414 VDD.n8370 0.04025
R39513 VDD.n10410 VDD.n8370 0.04025
R39514 VDD.n10410 VDD.n10409 0.04025
R39515 VDD.n10409 VDD.n10408 0.04025
R39516 VDD.n10408 VDD.n8372 0.04025
R39517 VDD.n10404 VDD.n8372 0.04025
R39518 VDD.n10404 VDD.n10403 0.04025
R39519 VDD.n10403 VDD.n10402 0.04025
R39520 VDD.n10402 VDD.n8374 0.04025
R39521 VDD.n10398 VDD.n8374 0.04025
R39522 VDD.n10398 VDD.n10397 0.04025
R39523 VDD.n10397 VDD.n10396 0.04025
R39524 VDD.n10396 VDD.n8376 0.04025
R39525 VDD.n10392 VDD.n8376 0.04025
R39526 VDD.n10392 VDD.n10391 0.04025
R39527 VDD.n10391 VDD.n10390 0.04025
R39528 VDD.n10390 VDD.n8378 0.04025
R39529 VDD.n10386 VDD.n8378 0.04025
R39530 VDD.n10386 VDD.n10385 0.04025
R39531 VDD.n10385 VDD.n10384 0.04025
R39532 VDD.n10384 VDD.n8380 0.04025
R39533 VDD.n10380 VDD.n8380 0.04025
R39534 VDD.n10380 VDD.n10379 0.04025
R39535 VDD.n10379 VDD.n10378 0.04025
R39536 VDD.n10378 VDD.n8382 0.04025
R39537 VDD.n10374 VDD.n8382 0.04025
R39538 VDD.n10374 VDD.n10373 0.04025
R39539 VDD.n10373 VDD.n10372 0.04025
R39540 VDD.n10372 VDD.n8384 0.04025
R39541 VDD.n10368 VDD.n8384 0.04025
R39542 VDD.n10368 VDD.n10367 0.04025
R39543 VDD.n10367 VDD.n10366 0.04025
R39544 VDD.n10366 VDD.n8386 0.04025
R39545 VDD.n10362 VDD.n8386 0.04025
R39546 VDD.n10362 VDD.n10361 0.04025
R39547 VDD.n10361 VDD.n10360 0.04025
R39548 VDD.n10360 VDD.n8388 0.04025
R39549 VDD.n10356 VDD.n8388 0.04025
R39550 VDD.n10356 VDD.n10355 0.04025
R39551 VDD.n10355 VDD.n10354 0.04025
R39552 VDD.n10354 VDD.n8390 0.04025
R39553 VDD.n10350 VDD.n8390 0.04025
R39554 VDD.n10350 VDD.n10349 0.04025
R39555 VDD.n10349 VDD.n10348 0.04025
R39556 VDD.n10348 VDD.n8392 0.04025
R39557 VDD.n10344 VDD.n8392 0.04025
R39558 VDD.n10344 VDD.n10343 0.04025
R39559 VDD.n10343 VDD.n10342 0.04025
R39560 VDD.n10342 VDD.n8394 0.04025
R39561 VDD.n10338 VDD.n8394 0.04025
R39562 VDD.n10338 VDD.n10337 0.04025
R39563 VDD.n10337 VDD.n10336 0.04025
R39564 VDD.n10336 VDD.n8396 0.04025
R39565 VDD.n10332 VDD.n8396 0.04025
R39566 VDD.n10332 VDD.n10331 0.04025
R39567 VDD.n10331 VDD.n10330 0.04025
R39568 VDD.n10330 VDD.n8398 0.04025
R39569 VDD.n10326 VDD.n8398 0.04025
R39570 VDD.n10326 VDD.n10325 0.04025
R39571 VDD.n10325 VDD.n10324 0.04025
R39572 VDD.n10324 VDD.n8400 0.04025
R39573 VDD.n10320 VDD.n8400 0.04025
R39574 VDD.n10320 VDD.n10319 0.04025
R39575 VDD.n10319 VDD.n10318 0.04025
R39576 VDD.n10318 VDD.n8402 0.04025
R39577 VDD.n10314 VDD.n8402 0.04025
R39578 VDD.n10314 VDD.n10313 0.04025
R39579 VDD.n10313 VDD.n10312 0.04025
R39580 VDD.n10312 VDD.n8404 0.04025
R39581 VDD.n10308 VDD.n8404 0.04025
R39582 VDD.n10308 VDD.n10307 0.04025
R39583 VDD.n10307 VDD.n10306 0.04025
R39584 VDD.n10306 VDD.n8406 0.04025
R39585 VDD.n10302 VDD.n8406 0.04025
R39586 VDD.n10302 VDD.n10301 0.04025
R39587 VDD.n10301 VDD.n10300 0.04025
R39588 VDD.n10300 VDD.n8408 0.04025
R39589 VDD.n10296 VDD.n8408 0.04025
R39590 VDD.n10296 VDD.n10295 0.04025
R39591 VDD.n10295 VDD.n10294 0.04025
R39592 VDD.n10294 VDD.n8410 0.04025
R39593 VDD.n10290 VDD.n8410 0.04025
R39594 VDD.n10290 VDD.n10289 0.04025
R39595 VDD.n10289 VDD.n10288 0.04025
R39596 VDD.n10288 VDD.n8412 0.04025
R39597 VDD.n10284 VDD.n8412 0.04025
R39598 VDD.n10284 VDD.n10283 0.04025
R39599 VDD.n10283 VDD.n10282 0.04025
R39600 VDD.n10282 VDD.n8414 0.04025
R39601 VDD.n10278 VDD.n8414 0.04025
R39602 VDD.n10278 VDD.n10277 0.04025
R39603 VDD.n10277 VDD.n10276 0.04025
R39604 VDD.n10276 VDD.n8416 0.04025
R39605 VDD.n10272 VDD.n8416 0.04025
R39606 VDD.n10272 VDD.n10271 0.04025
R39607 VDD.n10271 VDD.n10270 0.04025
R39608 VDD.n10270 VDD.n8418 0.04025
R39609 VDD.n10266 VDD.n8418 0.04025
R39610 VDD.n10266 VDD.n10265 0.04025
R39611 VDD.n10265 VDD.n10264 0.04025
R39612 VDD.n10264 VDD.n8420 0.04025
R39613 VDD.n10260 VDD.n8420 0.04025
R39614 VDD.n10260 VDD.n10259 0.04025
R39615 VDD.n10259 VDD.n10258 0.04025
R39616 VDD.n10258 VDD.n8422 0.04025
R39617 VDD.n10254 VDD.n8422 0.04025
R39618 VDD.n10254 VDD.n10253 0.04025
R39619 VDD.n10253 VDD.n10252 0.04025
R39620 VDD.n10252 VDD.n8424 0.04025
R39621 VDD.n10248 VDD.n8424 0.04025
R39622 VDD.n10248 VDD.n10247 0.04025
R39623 VDD.n10247 VDD.n10246 0.04025
R39624 VDD.n10246 VDD.n8426 0.04025
R39625 VDD.n10242 VDD.n8426 0.04025
R39626 VDD.n10242 VDD.n10241 0.04025
R39627 VDD.n10241 VDD.n10240 0.04025
R39628 VDD.n10240 VDD.n8428 0.04025
R39629 VDD.n10236 VDD.n8428 0.04025
R39630 VDD.n10236 VDD.n10235 0.04025
R39631 VDD.n10235 VDD.n10234 0.04025
R39632 VDD.n10234 VDD.n8430 0.04025
R39633 VDD.n10230 VDD.n8430 0.04025
R39634 VDD.n10230 VDD.n10229 0.04025
R39635 VDD.n10229 VDD.n10228 0.04025
R39636 VDD.n10228 VDD.n8432 0.04025
R39637 VDD.n10224 VDD.n8432 0.04025
R39638 VDD.n10224 VDD.n10223 0.04025
R39639 VDD.n10223 VDD.n10222 0.04025
R39640 VDD.n10222 VDD.n8434 0.04025
R39641 VDD.n10218 VDD.n8434 0.04025
R39642 VDD.n10218 VDD.n10217 0.04025
R39643 VDD.n10217 VDD.n10216 0.04025
R39644 VDD.n10216 VDD.n8436 0.04025
R39645 VDD.n10212 VDD.n8436 0.04025
R39646 VDD.n10212 VDD.n10211 0.04025
R39647 VDD.n10211 VDD.n10210 0.04025
R39648 VDD.n10210 VDD.n8438 0.04025
R39649 VDD.n10206 VDD.n8438 0.04025
R39650 VDD.n10206 VDD.n10205 0.04025
R39651 VDD.n10205 VDD.n10204 0.04025
R39652 VDD.n10204 VDD.n8440 0.04025
R39653 VDD.n10200 VDD.n8440 0.04025
R39654 VDD.n10200 VDD.n10199 0.04025
R39655 VDD.n10199 VDD.n10198 0.04025
R39656 VDD.n10198 VDD.n8442 0.04025
R39657 VDD.n10194 VDD.n8442 0.04025
R39658 VDD.n10194 VDD.n10193 0.04025
R39659 VDD.n10193 VDD.n10192 0.04025
R39660 VDD.n10192 VDD.n8444 0.04025
R39661 VDD.n10188 VDD.n8444 0.04025
R39662 VDD.n10188 VDD.n10187 0.04025
R39663 VDD.n10187 VDD.n10186 0.04025
R39664 VDD.n10186 VDD.n8446 0.04025
R39665 VDD.n10182 VDD.n8446 0.04025
R39666 VDD.n10182 VDD.n10181 0.04025
R39667 VDD.n10181 VDD.n10180 0.04025
R39668 VDD.n10180 VDD.n8448 0.04025
R39669 VDD.n10176 VDD.n8448 0.04025
R39670 VDD.n10176 VDD.n10175 0.04025
R39671 VDD.n10175 VDD.n10174 0.04025
R39672 VDD.n10174 VDD.n8450 0.04025
R39673 VDD.n10170 VDD.n8450 0.04025
R39674 VDD.n10170 VDD.n10169 0.04025
R39675 VDD.n10169 VDD.n10168 0.04025
R39676 VDD.n10168 VDD.n8452 0.04025
R39677 VDD.n10164 VDD.n8452 0.04025
R39678 VDD.n10164 VDD.n10163 0.04025
R39679 VDD.n10163 VDD.n10162 0.04025
R39680 VDD.n10162 VDD.n8454 0.04025
R39681 VDD.n10158 VDD.n8454 0.04025
R39682 VDD.n10158 VDD.n10157 0.04025
R39683 VDD.n10157 VDD.n10156 0.04025
R39684 VDD.n10156 VDD.n8456 0.04025
R39685 VDD.n10152 VDD.n8456 0.04025
R39686 VDD.n10152 VDD.n10151 0.04025
R39687 VDD.n10151 VDD.n10150 0.04025
R39688 VDD.n10150 VDD.n8458 0.04025
R39689 VDD.n10146 VDD.n9200 0.04025
R39690 VDD.n10146 VDD.n10145 0.04025
R39691 VDD.n10145 VDD.n10144 0.04025
R39692 VDD.n10144 VDD.n9201 0.04025
R39693 VDD.n10140 VDD.n9201 0.04025
R39694 VDD.n10140 VDD.n10139 0.04025
R39695 VDD.n10139 VDD.n10138 0.04025
R39696 VDD.n10138 VDD.n9203 0.04025
R39697 VDD.n10134 VDD.n9203 0.04025
R39698 VDD.n10134 VDD.n10133 0.04025
R39699 VDD.n10133 VDD.n10132 0.04025
R39700 VDD.n10132 VDD.n9205 0.04025
R39701 VDD.n10128 VDD.n9205 0.04025
R39702 VDD.n10128 VDD.n10127 0.04025
R39703 VDD.n10127 VDD.n10126 0.04025
R39704 VDD.n10126 VDD.n9207 0.04025
R39705 VDD.n10122 VDD.n9207 0.04025
R39706 VDD.n10122 VDD.n10121 0.04025
R39707 VDD.n10121 VDD.n10120 0.04025
R39708 VDD.n10120 VDD.n9209 0.04025
R39709 VDD.n10116 VDD.n9209 0.04025
R39710 VDD.n10116 VDD.n10115 0.04025
R39711 VDD.n10115 VDD.n10114 0.04025
R39712 VDD.n10114 VDD.n9211 0.04025
R39713 VDD.n10110 VDD.n9211 0.04025
R39714 VDD.n10110 VDD.n10109 0.04025
R39715 VDD.n10109 VDD.n10108 0.04025
R39716 VDD.n10108 VDD.n9213 0.04025
R39717 VDD.n10104 VDD.n9213 0.04025
R39718 VDD.n10104 VDD.n10103 0.04025
R39719 VDD.n10147 VDD.n9186 0.04025
R39720 VDD.n10143 VDD.n9186 0.04025
R39721 VDD.n10143 VDD.n10142 0.04025
R39722 VDD.n10142 VDD.n10141 0.04025
R39723 VDD.n10141 VDD.n9202 0.04025
R39724 VDD.n10137 VDD.n9202 0.04025
R39725 VDD.n10137 VDD.n10136 0.04025
R39726 VDD.n10136 VDD.n10135 0.04025
R39727 VDD.n10135 VDD.n9204 0.04025
R39728 VDD.n10131 VDD.n9204 0.04025
R39729 VDD.n10131 VDD.n10130 0.04025
R39730 VDD.n10130 VDD.n10129 0.04025
R39731 VDD.n10129 VDD.n9206 0.04025
R39732 VDD.n10125 VDD.n9206 0.04025
R39733 VDD.n10125 VDD.n10124 0.04025
R39734 VDD.n10124 VDD.n10123 0.04025
R39735 VDD.n10123 VDD.n9208 0.04025
R39736 VDD.n10119 VDD.n9208 0.04025
R39737 VDD.n10119 VDD.n10118 0.04025
R39738 VDD.n10118 VDD.n10117 0.04025
R39739 VDD.n10117 VDD.n9210 0.04025
R39740 VDD.n10113 VDD.n9210 0.04025
R39741 VDD.n10113 VDD.n10112 0.04025
R39742 VDD.n10112 VDD.n10111 0.04025
R39743 VDD.n10111 VDD.n9212 0.04025
R39744 VDD.n10107 VDD.n9212 0.04025
R39745 VDD.n10107 VDD.n10106 0.04025
R39746 VDD.n10106 VDD.n10105 0.04025
R39747 VDD.n10105 VDD.n9214 0.04025
R39748 VDD.n9439 VDD.n9436 0.04025
R39749 VDD.n9440 VDD.n9439 0.04025
R39750 VDD.n9441 VDD.n9440 0.04025
R39751 VDD.n9441 VDD.n9434 0.04025
R39752 VDD.n9445 VDD.n9434 0.04025
R39753 VDD.n9446 VDD.n9445 0.04025
R39754 VDD.n9447 VDD.n9446 0.04025
R39755 VDD.n9447 VDD.n9432 0.04025
R39756 VDD.n9451 VDD.n9432 0.04025
R39757 VDD.n9452 VDD.n9451 0.04025
R39758 VDD.n9453 VDD.n9452 0.04025
R39759 VDD.n9453 VDD.n9430 0.04025
R39760 VDD.n9457 VDD.n9430 0.04025
R39761 VDD.n9458 VDD.n9457 0.04025
R39762 VDD.n9459 VDD.n9458 0.04025
R39763 VDD.n9459 VDD.n9428 0.04025
R39764 VDD.n9463 VDD.n9428 0.04025
R39765 VDD.n9464 VDD.n9463 0.04025
R39766 VDD.n9465 VDD.n9464 0.04025
R39767 VDD.n9465 VDD.n9426 0.04025
R39768 VDD.n9469 VDD.n9426 0.04025
R39769 VDD.n9470 VDD.n9469 0.04025
R39770 VDD.n9471 VDD.n9470 0.04025
R39771 VDD.n9471 VDD.n9424 0.04025
R39772 VDD.n9475 VDD.n9424 0.04025
R39773 VDD.n9476 VDD.n9475 0.04025
R39774 VDD.n9477 VDD.n9476 0.04025
R39775 VDD.n9477 VDD.n9422 0.04025
R39776 VDD.n9481 VDD.n9422 0.04025
R39777 VDD.n9482 VDD.n9481 0.04025
R39778 VDD.n9483 VDD.n9482 0.04025
R39779 VDD.n9483 VDD.n9420 0.04025
R39780 VDD.n9487 VDD.n9420 0.04025
R39781 VDD.n9488 VDD.n9487 0.04025
R39782 VDD.n9489 VDD.n9488 0.04025
R39783 VDD.n9489 VDD.n9418 0.04025
R39784 VDD.n9493 VDD.n9418 0.04025
R39785 VDD.n9494 VDD.n9493 0.04025
R39786 VDD.n9495 VDD.n9494 0.04025
R39787 VDD.n9495 VDD.n9416 0.04025
R39788 VDD.n9499 VDD.n9416 0.04025
R39789 VDD.n9500 VDD.n9499 0.04025
R39790 VDD.n9501 VDD.n9500 0.04025
R39791 VDD.n9501 VDD.n9414 0.04025
R39792 VDD.n9505 VDD.n9414 0.04025
R39793 VDD.n9506 VDD.n9505 0.04025
R39794 VDD.n9507 VDD.n9506 0.04025
R39795 VDD.n9507 VDD.n9412 0.04025
R39796 VDD.n9511 VDD.n9412 0.04025
R39797 VDD.n9512 VDD.n9511 0.04025
R39798 VDD.n9513 VDD.n9512 0.04025
R39799 VDD.n9513 VDD.n9410 0.04025
R39800 VDD.n9517 VDD.n9410 0.04025
R39801 VDD.n9518 VDD.n9517 0.04025
R39802 VDD.n9519 VDD.n9518 0.04025
R39803 VDD.n9519 VDD.n9408 0.04025
R39804 VDD.n9523 VDD.n9408 0.04025
R39805 VDD.n9524 VDD.n9523 0.04025
R39806 VDD.n9525 VDD.n9524 0.04025
R39807 VDD.n9525 VDD.n9406 0.04025
R39808 VDD.n9529 VDD.n9406 0.04025
R39809 VDD.n9530 VDD.n9529 0.04025
R39810 VDD.n9531 VDD.n9530 0.04025
R39811 VDD.n9531 VDD.n9404 0.04025
R39812 VDD.n9535 VDD.n9404 0.04025
R39813 VDD.n9536 VDD.n9535 0.04025
R39814 VDD.n9537 VDD.n9536 0.04025
R39815 VDD.n9537 VDD.n9402 0.04025
R39816 VDD.n9541 VDD.n9402 0.04025
R39817 VDD.n9542 VDD.n9541 0.04025
R39818 VDD.n9543 VDD.n9542 0.04025
R39819 VDD.n9543 VDD.n9400 0.04025
R39820 VDD.n9547 VDD.n9400 0.04025
R39821 VDD.n9548 VDD.n9547 0.04025
R39822 VDD.n9549 VDD.n9548 0.04025
R39823 VDD.n9549 VDD.n9398 0.04025
R39824 VDD.n9553 VDD.n9398 0.04025
R39825 VDD.n9554 VDD.n9553 0.04025
R39826 VDD.n9555 VDD.n9554 0.04025
R39827 VDD.n9555 VDD.n9396 0.04025
R39828 VDD.n9559 VDD.n9396 0.04025
R39829 VDD.n9560 VDD.n9559 0.04025
R39830 VDD.n9561 VDD.n9560 0.04025
R39831 VDD.n9561 VDD.n9394 0.04025
R39832 VDD.n9565 VDD.n9394 0.04025
R39833 VDD.n9566 VDD.n9565 0.04025
R39834 VDD.n9567 VDD.n9566 0.04025
R39835 VDD.n9567 VDD.n9392 0.04025
R39836 VDD.n9571 VDD.n9392 0.04025
R39837 VDD.n9572 VDD.n9571 0.04025
R39838 VDD.n9573 VDD.n9572 0.04025
R39839 VDD.n9573 VDD.n9390 0.04025
R39840 VDD.n9577 VDD.n9390 0.04025
R39841 VDD.n9578 VDD.n9577 0.04025
R39842 VDD.n9579 VDD.n9578 0.04025
R39843 VDD.n9579 VDD.n9388 0.04025
R39844 VDD.n9583 VDD.n9388 0.04025
R39845 VDD.n9584 VDD.n9583 0.04025
R39846 VDD.n9585 VDD.n9584 0.04025
R39847 VDD.n9585 VDD.n9386 0.04025
R39848 VDD.n9589 VDD.n9386 0.04025
R39849 VDD.n9590 VDD.n9589 0.04025
R39850 VDD.n9591 VDD.n9590 0.04025
R39851 VDD.n9591 VDD.n9384 0.04025
R39852 VDD.n9595 VDD.n9384 0.04025
R39853 VDD.n9596 VDD.n9595 0.04025
R39854 VDD.n9597 VDD.n9596 0.04025
R39855 VDD.n9597 VDD.n9382 0.04025
R39856 VDD.n9601 VDD.n9382 0.04025
R39857 VDD.n9602 VDD.n9601 0.04025
R39858 VDD.n9603 VDD.n9602 0.04025
R39859 VDD.n9603 VDD.n9380 0.04025
R39860 VDD.n9607 VDD.n9380 0.04025
R39861 VDD.n9608 VDD.n9607 0.04025
R39862 VDD.n9609 VDD.n9608 0.04025
R39863 VDD.n9609 VDD.n9378 0.04025
R39864 VDD.n9613 VDD.n9378 0.04025
R39865 VDD.n9614 VDD.n9613 0.04025
R39866 VDD.n9615 VDD.n9614 0.04025
R39867 VDD.n9615 VDD.n9376 0.04025
R39868 VDD.n9619 VDD.n9376 0.04025
R39869 VDD.n9620 VDD.n9619 0.04025
R39870 VDD.n9621 VDD.n9620 0.04025
R39871 VDD.n9621 VDD.n9374 0.04025
R39872 VDD.n9625 VDD.n9374 0.04025
R39873 VDD.n9626 VDD.n9625 0.04025
R39874 VDD.n9627 VDD.n9626 0.04025
R39875 VDD.n9627 VDD.n9372 0.04025
R39876 VDD.n9631 VDD.n9372 0.04025
R39877 VDD.n9632 VDD.n9631 0.04025
R39878 VDD.n9633 VDD.n9632 0.04025
R39879 VDD.n9633 VDD.n9370 0.04025
R39880 VDD.n9637 VDD.n9370 0.04025
R39881 VDD.n9638 VDD.n9637 0.04025
R39882 VDD.n9639 VDD.n9638 0.04025
R39883 VDD.n9639 VDD.n9368 0.04025
R39884 VDD.n9643 VDD.n9368 0.04025
R39885 VDD.n9644 VDD.n9643 0.04025
R39886 VDD.n9645 VDD.n9644 0.04025
R39887 VDD.n9645 VDD.n9366 0.04025
R39888 VDD.n9649 VDD.n9366 0.04025
R39889 VDD.n9650 VDD.n9649 0.04025
R39890 VDD.n9651 VDD.n9650 0.04025
R39891 VDD.n9651 VDD.n9364 0.04025
R39892 VDD.n9655 VDD.n9364 0.04025
R39893 VDD.n9656 VDD.n9655 0.04025
R39894 VDD.n9657 VDD.n9656 0.04025
R39895 VDD.n9657 VDD.n9362 0.04025
R39896 VDD.n9661 VDD.n9362 0.04025
R39897 VDD.n9662 VDD.n9661 0.04025
R39898 VDD.n9663 VDD.n9662 0.04025
R39899 VDD.n9663 VDD.n9360 0.04025
R39900 VDD.n9667 VDD.n9360 0.04025
R39901 VDD.n9668 VDD.n9667 0.04025
R39902 VDD.n9669 VDD.n9668 0.04025
R39903 VDD.n9669 VDD.n9358 0.04025
R39904 VDD.n9673 VDD.n9358 0.04025
R39905 VDD.n9674 VDD.n9673 0.04025
R39906 VDD.n9675 VDD.n9674 0.04025
R39907 VDD.n9675 VDD.n9356 0.04025
R39908 VDD.n9679 VDD.n9356 0.04025
R39909 VDD.n9680 VDD.n9679 0.04025
R39910 VDD.n9681 VDD.n9680 0.04025
R39911 VDD.n9681 VDD.n9354 0.04025
R39912 VDD.n9685 VDD.n9354 0.04025
R39913 VDD.n9686 VDD.n9685 0.04025
R39914 VDD.n9687 VDD.n9686 0.04025
R39915 VDD.n9687 VDD.n9352 0.04025
R39916 VDD.n9691 VDD.n9352 0.04025
R39917 VDD.n9692 VDD.n9691 0.04025
R39918 VDD.n9693 VDD.n9692 0.04025
R39919 VDD.n9693 VDD.n9350 0.04025
R39920 VDD.n9697 VDD.n9350 0.04025
R39921 VDD.n9698 VDD.n9697 0.04025
R39922 VDD.n9699 VDD.n9698 0.04025
R39923 VDD.n9699 VDD.n9348 0.04025
R39924 VDD.n9703 VDD.n9348 0.04025
R39925 VDD.n9704 VDD.n9703 0.04025
R39926 VDD.n9705 VDD.n9704 0.04025
R39927 VDD.n9705 VDD.n9346 0.04025
R39928 VDD.n9709 VDD.n9346 0.04025
R39929 VDD.n9710 VDD.n9709 0.04025
R39930 VDD.n9711 VDD.n9710 0.04025
R39931 VDD.n9711 VDD.n9344 0.04025
R39932 VDD.n9715 VDD.n9344 0.04025
R39933 VDD.n9716 VDD.n9715 0.04025
R39934 VDD.n9717 VDD.n9716 0.04025
R39935 VDD.n9717 VDD.n9342 0.04025
R39936 VDD.n9721 VDD.n9342 0.04025
R39937 VDD.n9722 VDD.n9721 0.04025
R39938 VDD.n9723 VDD.n9722 0.04025
R39939 VDD.n9723 VDD.n9340 0.04025
R39940 VDD.n9727 VDD.n9340 0.04025
R39941 VDD.n9728 VDD.n9727 0.04025
R39942 VDD.n9729 VDD.n9728 0.04025
R39943 VDD.n9729 VDD.n9338 0.04025
R39944 VDD.n9733 VDD.n9338 0.04025
R39945 VDD.n9734 VDD.n9733 0.04025
R39946 VDD.n9735 VDD.n9734 0.04025
R39947 VDD.n9735 VDD.n9336 0.04025
R39948 VDD.n9739 VDD.n9336 0.04025
R39949 VDD.n9740 VDD.n9739 0.04025
R39950 VDD.n9741 VDD.n9740 0.04025
R39951 VDD.n9741 VDD.n9334 0.04025
R39952 VDD.n9745 VDD.n9334 0.04025
R39953 VDD.n9746 VDD.n9745 0.04025
R39954 VDD.n9747 VDD.n9746 0.04025
R39955 VDD.n9747 VDD.n9332 0.04025
R39956 VDD.n9751 VDD.n9332 0.04025
R39957 VDD.n9752 VDD.n9751 0.04025
R39958 VDD.n9753 VDD.n9752 0.04025
R39959 VDD.n9753 VDD.n9330 0.04025
R39960 VDD.n9757 VDD.n9330 0.04025
R39961 VDD.n9758 VDD.n9757 0.04025
R39962 VDD.n9759 VDD.n9758 0.04025
R39963 VDD.n9759 VDD.n9328 0.04025
R39964 VDD.n9763 VDD.n9328 0.04025
R39965 VDD.n9764 VDD.n9763 0.04025
R39966 VDD.n9765 VDD.n9764 0.04025
R39967 VDD.n9765 VDD.n9326 0.04025
R39968 VDD.n9769 VDD.n9326 0.04025
R39969 VDD.n9770 VDD.n9769 0.04025
R39970 VDD.n9771 VDD.n9770 0.04025
R39971 VDD.n9771 VDD.n9324 0.04025
R39972 VDD.n9775 VDD.n9324 0.04025
R39973 VDD.n9776 VDD.n9775 0.04025
R39974 VDD.n9777 VDD.n9776 0.04025
R39975 VDD.n9777 VDD.n9322 0.04025
R39976 VDD.n9781 VDD.n9322 0.04025
R39977 VDD.n9782 VDD.n9781 0.04025
R39978 VDD.n9783 VDD.n9782 0.04025
R39979 VDD.n9783 VDD.n9320 0.04025
R39980 VDD.n9787 VDD.n9320 0.04025
R39981 VDD.n9788 VDD.n9787 0.04025
R39982 VDD.n9789 VDD.n9788 0.04025
R39983 VDD.n9789 VDD.n9318 0.04025
R39984 VDD.n9793 VDD.n9318 0.04025
R39985 VDD.n9794 VDD.n9793 0.04025
R39986 VDD.n9795 VDD.n9794 0.04025
R39987 VDD.n9795 VDD.n9316 0.04025
R39988 VDD.n9799 VDD.n9316 0.04025
R39989 VDD.n9800 VDD.n9799 0.04025
R39990 VDD.n9801 VDD.n9800 0.04025
R39991 VDD.n9801 VDD.n9314 0.04025
R39992 VDD.n9805 VDD.n9314 0.04025
R39993 VDD.n9806 VDD.n9805 0.04025
R39994 VDD.n9807 VDD.n9806 0.04025
R39995 VDD.n9807 VDD.n9312 0.04025
R39996 VDD.n9811 VDD.n9312 0.04025
R39997 VDD.n9812 VDD.n9811 0.04025
R39998 VDD.n9813 VDD.n9812 0.04025
R39999 VDD.n9813 VDD.n9310 0.04025
R40000 VDD.n9817 VDD.n9310 0.04025
R40001 VDD.n9818 VDD.n9817 0.04025
R40002 VDD.n9819 VDD.n9818 0.04025
R40003 VDD.n9819 VDD.n9308 0.04025
R40004 VDD.n9823 VDD.n9308 0.04025
R40005 VDD.n9824 VDD.n9823 0.04025
R40006 VDD.n9825 VDD.n9824 0.04025
R40007 VDD.n9825 VDD.n9306 0.04025
R40008 VDD.n9829 VDD.n9306 0.04025
R40009 VDD.n9830 VDD.n9829 0.04025
R40010 VDD.n9831 VDD.n9830 0.04025
R40011 VDD.n9831 VDD.n9304 0.04025
R40012 VDD.n9835 VDD.n9304 0.04025
R40013 VDD.n9836 VDD.n9835 0.04025
R40014 VDD.n9837 VDD.n9836 0.04025
R40015 VDD.n9837 VDD.n9302 0.04025
R40016 VDD.n9841 VDD.n9302 0.04025
R40017 VDD.n9842 VDD.n9841 0.04025
R40018 VDD.n9843 VDD.n9842 0.04025
R40019 VDD.n9843 VDD.n9300 0.04025
R40020 VDD.n9847 VDD.n9300 0.04025
R40021 VDD.n9848 VDD.n9847 0.04025
R40022 VDD.n9849 VDD.n9848 0.04025
R40023 VDD.n9849 VDD.n9298 0.04025
R40024 VDD.n9853 VDD.n9298 0.04025
R40025 VDD.n9854 VDD.n9853 0.04025
R40026 VDD.n9855 VDD.n9854 0.04025
R40027 VDD.n9855 VDD.n9296 0.04025
R40028 VDD.n9859 VDD.n9296 0.04025
R40029 VDD.n9860 VDD.n9859 0.04025
R40030 VDD.n9861 VDD.n9860 0.04025
R40031 VDD.n9861 VDD.n9294 0.04025
R40032 VDD.n9865 VDD.n9294 0.04025
R40033 VDD.n9866 VDD.n9865 0.04025
R40034 VDD.n9867 VDD.n9866 0.04025
R40035 VDD.n9867 VDD.n9292 0.04025
R40036 VDD.n9871 VDD.n9292 0.04025
R40037 VDD.n9872 VDD.n9871 0.04025
R40038 VDD.n9873 VDD.n9872 0.04025
R40039 VDD.n9873 VDD.n9290 0.04025
R40040 VDD.n9877 VDD.n9290 0.04025
R40041 VDD.n9878 VDD.n9877 0.04025
R40042 VDD.n9879 VDD.n9878 0.04025
R40043 VDD.n9879 VDD.n9288 0.04025
R40044 VDD.n9883 VDD.n9288 0.04025
R40045 VDD.n9884 VDD.n9883 0.04025
R40046 VDD.n9885 VDD.n9884 0.04025
R40047 VDD.n9885 VDD.n9286 0.04025
R40048 VDD.n9889 VDD.n9286 0.04025
R40049 VDD.n9890 VDD.n9889 0.04025
R40050 VDD.n9891 VDD.n9890 0.04025
R40051 VDD.n9891 VDD.n9284 0.04025
R40052 VDD.n9895 VDD.n9284 0.04025
R40053 VDD.n9896 VDD.n9895 0.04025
R40054 VDD.n9897 VDD.n9896 0.04025
R40055 VDD.n9897 VDD.n9282 0.04025
R40056 VDD.n9901 VDD.n9282 0.04025
R40057 VDD.n9902 VDD.n9901 0.04025
R40058 VDD.n9903 VDD.n9902 0.04025
R40059 VDD.n9903 VDD.n9280 0.04025
R40060 VDD.n9907 VDD.n9280 0.04025
R40061 VDD.n9908 VDD.n9907 0.04025
R40062 VDD.n9909 VDD.n9908 0.04025
R40063 VDD.n9909 VDD.n9278 0.04025
R40064 VDD.n9913 VDD.n9278 0.04025
R40065 VDD.n9914 VDD.n9913 0.04025
R40066 VDD.n9915 VDD.n9914 0.04025
R40067 VDD.n9915 VDD.n9276 0.04025
R40068 VDD.n9919 VDD.n9276 0.04025
R40069 VDD.n9920 VDD.n9919 0.04025
R40070 VDD.n9921 VDD.n9920 0.04025
R40071 VDD.n9921 VDD.n9274 0.04025
R40072 VDD.n9925 VDD.n9274 0.04025
R40073 VDD.n9926 VDD.n9925 0.04025
R40074 VDD.n9927 VDD.n9926 0.04025
R40075 VDD.n9927 VDD.n9272 0.04025
R40076 VDD.n9931 VDD.n9272 0.04025
R40077 VDD.n9932 VDD.n9931 0.04025
R40078 VDD.n9933 VDD.n9932 0.04025
R40079 VDD.n9933 VDD.n9270 0.04025
R40080 VDD.n9937 VDD.n9270 0.04025
R40081 VDD.n9938 VDD.n9937 0.04025
R40082 VDD.n9939 VDD.n9938 0.04025
R40083 VDD.n9939 VDD.n9268 0.04025
R40084 VDD.n9943 VDD.n9268 0.04025
R40085 VDD.n9944 VDD.n9943 0.04025
R40086 VDD.n9945 VDD.n9944 0.04025
R40087 VDD.n9945 VDD.n9266 0.04025
R40088 VDD.n9949 VDD.n9266 0.04025
R40089 VDD.n9950 VDD.n9949 0.04025
R40090 VDD.n9951 VDD.n9950 0.04025
R40091 VDD.n9951 VDD.n9264 0.04025
R40092 VDD.n9955 VDD.n9264 0.04025
R40093 VDD.n9956 VDD.n9955 0.04025
R40094 VDD.n9957 VDD.n9956 0.04025
R40095 VDD.n9957 VDD.n9262 0.04025
R40096 VDD.n9961 VDD.n9262 0.04025
R40097 VDD.n9962 VDD.n9961 0.04025
R40098 VDD.n9963 VDD.n9962 0.04025
R40099 VDD.n9963 VDD.n9260 0.04025
R40100 VDD.n9967 VDD.n9260 0.04025
R40101 VDD.n9968 VDD.n9967 0.04025
R40102 VDD.n9969 VDD.n9968 0.04025
R40103 VDD.n9969 VDD.n9258 0.04025
R40104 VDD.n9973 VDD.n9258 0.04025
R40105 VDD.n9974 VDD.n9973 0.04025
R40106 VDD.n9975 VDD.n9974 0.04025
R40107 VDD.n9975 VDD.n9256 0.04025
R40108 VDD.n9979 VDD.n9256 0.04025
R40109 VDD.n9980 VDD.n9979 0.04025
R40110 VDD.n9981 VDD.n9980 0.04025
R40111 VDD.n9981 VDD.n9254 0.04025
R40112 VDD.n9985 VDD.n9254 0.04025
R40113 VDD.n9986 VDD.n9985 0.04025
R40114 VDD.n9987 VDD.n9986 0.04025
R40115 VDD.n9987 VDD.n9252 0.04025
R40116 VDD.n9991 VDD.n9252 0.04025
R40117 VDD.n9992 VDD.n9991 0.04025
R40118 VDD.n9993 VDD.n9992 0.04025
R40119 VDD.n9993 VDD.n9250 0.04025
R40120 VDD.n9997 VDD.n9250 0.04025
R40121 VDD.n9998 VDD.n9997 0.04025
R40122 VDD.n9999 VDD.n9998 0.04025
R40123 VDD.n9999 VDD.n9248 0.04025
R40124 VDD.n10003 VDD.n9248 0.04025
R40125 VDD.n10004 VDD.n10003 0.04025
R40126 VDD.n10005 VDD.n10004 0.04025
R40127 VDD.n10005 VDD.n9246 0.04025
R40128 VDD.n10009 VDD.n9246 0.04025
R40129 VDD.n10010 VDD.n10009 0.04025
R40130 VDD.n10011 VDD.n10010 0.04025
R40131 VDD.n10011 VDD.n9244 0.04025
R40132 VDD.n10015 VDD.n9244 0.04025
R40133 VDD.n10016 VDD.n10015 0.04025
R40134 VDD.n10017 VDD.n10016 0.04025
R40135 VDD.n10017 VDD.n9242 0.04025
R40136 VDD.n10021 VDD.n9242 0.04025
R40137 VDD.n10022 VDD.n10021 0.04025
R40138 VDD.n10023 VDD.n10022 0.04025
R40139 VDD.n10023 VDD.n9240 0.04025
R40140 VDD.n10027 VDD.n9240 0.04025
R40141 VDD.n10028 VDD.n10027 0.04025
R40142 VDD.n10029 VDD.n10028 0.04025
R40143 VDD.n10029 VDD.n9238 0.04025
R40144 VDD.n10033 VDD.n9238 0.04025
R40145 VDD.n10034 VDD.n10033 0.04025
R40146 VDD.n10035 VDD.n10034 0.04025
R40147 VDD.n10035 VDD.n9236 0.04025
R40148 VDD.n10039 VDD.n9236 0.04025
R40149 VDD.n10040 VDD.n10039 0.04025
R40150 VDD.n10041 VDD.n10040 0.04025
R40151 VDD.n10041 VDD.n9234 0.04025
R40152 VDD.n10045 VDD.n9234 0.04025
R40153 VDD.n10046 VDD.n10045 0.04025
R40154 VDD.n10047 VDD.n10046 0.04025
R40155 VDD.n10047 VDD.n9232 0.04025
R40156 VDD.n10051 VDD.n9232 0.04025
R40157 VDD.n10052 VDD.n10051 0.04025
R40158 VDD.n10053 VDD.n10052 0.04025
R40159 VDD.n10053 VDD.n9230 0.04025
R40160 VDD.n10057 VDD.n9230 0.04025
R40161 VDD.n10058 VDD.n10057 0.04025
R40162 VDD.n10059 VDD.n10058 0.04025
R40163 VDD.n10059 VDD.n9228 0.04025
R40164 VDD.n10063 VDD.n9228 0.04025
R40165 VDD.n10064 VDD.n10063 0.04025
R40166 VDD.n10065 VDD.n10064 0.04025
R40167 VDD.n10065 VDD.n9226 0.04025
R40168 VDD.n10069 VDD.n9226 0.04025
R40169 VDD.n10070 VDD.n10069 0.04025
R40170 VDD.n10071 VDD.n10070 0.04025
R40171 VDD.n10071 VDD.n9224 0.04025
R40172 VDD.n10075 VDD.n9224 0.04025
R40173 VDD.n10076 VDD.n10075 0.04025
R40174 VDD.n10077 VDD.n10076 0.04025
R40175 VDD.n10077 VDD.n9222 0.04025
R40176 VDD.n10081 VDD.n9222 0.04025
R40177 VDD.n10082 VDD.n10081 0.04025
R40178 VDD.n10083 VDD.n10082 0.04025
R40179 VDD.n10083 VDD.n9220 0.04025
R40180 VDD.n10087 VDD.n9220 0.04025
R40181 VDD.n10088 VDD.n10087 0.04025
R40182 VDD.n10089 VDD.n10088 0.04025
R40183 VDD.n10089 VDD.n9218 0.04025
R40184 VDD.n10093 VDD.n9218 0.04025
R40185 VDD.n10094 VDD.n10093 0.04025
R40186 VDD.n10095 VDD.n10094 0.04025
R40187 VDD.n10095 VDD.n9216 0.04025
R40188 VDD.n10099 VDD.n9216 0.04025
R40189 VDD.n10100 VDD.n10099 0.04025
R40190 VDD.n10101 VDD.n10100 0.04025
R40191 VDD.n11814 VDD.n11813 0.04025
R40192 VDD.n11815 VDD.n11814 0.04025
R40193 VDD.n11815 VDD.n403 0.04025
R40194 VDD.n11819 VDD.n403 0.04025
R40195 VDD.n11820 VDD.n11819 0.04025
R40196 VDD.n11821 VDD.n11820 0.04025
R40197 VDD.n11821 VDD.n401 0.04025
R40198 VDD.n11825 VDD.n401 0.04025
R40199 VDD.n11826 VDD.n11825 0.04025
R40200 VDD.n11827 VDD.n11826 0.04025
R40201 VDD.n11827 VDD.n399 0.04025
R40202 VDD.n11831 VDD.n399 0.04025
R40203 VDD.n11832 VDD.n11831 0.04025
R40204 VDD.n11833 VDD.n11832 0.04025
R40205 VDD.n11833 VDD.n397 0.04025
R40206 VDD.n11837 VDD.n397 0.04025
R40207 VDD.n11838 VDD.n11837 0.04025
R40208 VDD.n11839 VDD.n11838 0.04025
R40209 VDD.n11839 VDD.n395 0.04025
R40210 VDD.n11843 VDD.n395 0.04025
R40211 VDD.n11844 VDD.n11843 0.04025
R40212 VDD.n11845 VDD.n11844 0.04025
R40213 VDD.n11845 VDD.n393 0.04025
R40214 VDD.n11849 VDD.n393 0.04025
R40215 VDD.n11850 VDD.n11849 0.04025
R40216 VDD.n11851 VDD.n11850 0.04025
R40217 VDD.n11851 VDD.n391 0.04025
R40218 VDD.n11855 VDD.n391 0.04025
R40219 VDD.n11856 VDD.n11855 0.04025
R40220 VDD.n11857 VDD.n11856 0.04025
R40221 VDD.n11857 VDD.n389 0.04025
R40222 VDD.n11861 VDD.n389 0.04025
R40223 VDD.n11862 VDD.n11861 0.04025
R40224 VDD.n11863 VDD.n11862 0.04025
R40225 VDD.n11863 VDD.n387 0.04025
R40226 VDD.n11867 VDD.n387 0.04025
R40227 VDD.n11868 VDD.n11867 0.04025
R40228 VDD.n11869 VDD.n11868 0.04025
R40229 VDD.n11869 VDD.n385 0.04025
R40230 VDD.n11874 VDD.n385 0.04025
R40231 VDD.n11875 VDD.n11874 0.04025
R40232 VDD.n11876 VDD.n11875 0.04025
R40233 VDD.n11876 VDD.n383 0.04025
R40234 VDD.n11880 VDD.n383 0.04025
R40235 VDD.n11881 VDD.n11880 0.04025
R40236 VDD.n11882 VDD.n11881 0.04025
R40237 VDD.n11882 VDD.n381 0.04025
R40238 VDD.n11886 VDD.n381 0.04025
R40239 VDD.n11887 VDD.n11886 0.04025
R40240 VDD.n11888 VDD.n11887 0.04025
R40241 VDD.n11888 VDD.n379 0.04025
R40242 VDD.n11892 VDD.n379 0.04025
R40243 VDD.n11893 VDD.n11892 0.04025
R40244 VDD.n11894 VDD.n11893 0.04025
R40245 VDD.n11894 VDD.n377 0.04025
R40246 VDD.n11898 VDD.n377 0.04025
R40247 VDD.n11899 VDD.n11898 0.04025
R40248 VDD.n11900 VDD.n11899 0.04025
R40249 VDD.n11900 VDD.n375 0.04025
R40250 VDD.n11904 VDD.n375 0.04025
R40251 VDD.n11905 VDD.n11904 0.04025
R40252 VDD.n11906 VDD.n11905 0.04025
R40253 VDD.n11906 VDD.n373 0.04025
R40254 VDD.n11910 VDD.n373 0.04025
R40255 VDD.n11911 VDD.n11910 0.04025
R40256 VDD.n11912 VDD.n11911 0.04025
R40257 VDD.n11912 VDD.n371 0.04025
R40258 VDD.n11916 VDD.n371 0.04025
R40259 VDD.n11917 VDD.n11916 0.04025
R40260 VDD.n11918 VDD.n11917 0.04025
R40261 VDD.n11918 VDD.n369 0.04025
R40262 VDD.n11922 VDD.n369 0.04025
R40263 VDD.n11923 VDD.n11922 0.04025
R40264 VDD.n11924 VDD.n11923 0.04025
R40265 VDD.n11924 VDD.n367 0.04025
R40266 VDD.n11928 VDD.n367 0.04025
R40267 VDD.n11929 VDD.n11928 0.04025
R40268 VDD.n11930 VDD.n11929 0.04025
R40269 VDD.n11930 VDD.n365 0.04025
R40270 VDD.n11934 VDD.n365 0.04025
R40271 VDD.n11935 VDD.n11934 0.04025
R40272 VDD.n11936 VDD.n11935 0.04025
R40273 VDD.n11936 VDD.n363 0.04025
R40274 VDD.n11940 VDD.n363 0.04025
R40275 VDD.n11941 VDD.n11940 0.04025
R40276 VDD.n11942 VDD.n11941 0.04025
R40277 VDD.n11942 VDD.n361 0.04025
R40278 VDD.n11946 VDD.n361 0.04025
R40279 VDD.n11947 VDD.n11946 0.04025
R40280 VDD.n11948 VDD.n11947 0.04025
R40281 VDD.n11948 VDD.n359 0.04025
R40282 VDD.n11952 VDD.n359 0.04025
R40283 VDD.n11953 VDD.n11952 0.04025
R40284 VDD.n11954 VDD.n11953 0.04025
R40285 VDD.n11954 VDD.n357 0.04025
R40286 VDD.n11958 VDD.n357 0.04025
R40287 VDD.n11959 VDD.n11958 0.04025
R40288 VDD.n11960 VDD.n11959 0.04025
R40289 VDD.n11960 VDD.n355 0.04025
R40290 VDD.n11964 VDD.n355 0.04025
R40291 VDD.n11965 VDD.n11964 0.04025
R40292 VDD.n11966 VDD.n11965 0.04025
R40293 VDD.n11966 VDD.n353 0.04025
R40294 VDD.n11970 VDD.n353 0.04025
R40295 VDD.n11971 VDD.n11970 0.04025
R40296 VDD.n11972 VDD.n11971 0.04025
R40297 VDD.n11972 VDD.n351 0.04025
R40298 VDD.n11976 VDD.n351 0.04025
R40299 VDD.n11977 VDD.n11976 0.04025
R40300 VDD.n11978 VDD.n11977 0.04025
R40301 VDD.n11978 VDD.n349 0.04025
R40302 VDD.n11982 VDD.n349 0.04025
R40303 VDD.n11983 VDD.n11982 0.04025
R40304 VDD.n11984 VDD.n11983 0.04025
R40305 VDD.n11984 VDD.n347 0.04025
R40306 VDD.n11988 VDD.n347 0.04025
R40307 VDD.n11989 VDD.n11988 0.04025
R40308 VDD.n11990 VDD.n11989 0.04025
R40309 VDD.n11990 VDD.n345 0.04025
R40310 VDD.n11994 VDD.n345 0.04025
R40311 VDD.n11995 VDD.n11994 0.04025
R40312 VDD.n11996 VDD.n11995 0.04025
R40313 VDD.n11996 VDD.n343 0.04025
R40314 VDD.n12000 VDD.n343 0.04025
R40315 VDD.n12001 VDD.n12000 0.04025
R40316 VDD.n12002 VDD.n12001 0.04025
R40317 VDD.n12002 VDD.n341 0.04025
R40318 VDD.n12006 VDD.n341 0.04025
R40319 VDD.n12007 VDD.n12006 0.04025
R40320 VDD.n12008 VDD.n12007 0.04025
R40321 VDD.n12008 VDD.n339 0.04025
R40322 VDD.n12012 VDD.n339 0.04025
R40323 VDD.n12013 VDD.n12012 0.04025
R40324 VDD.n12014 VDD.n12013 0.04025
R40325 VDD.n12014 VDD.n337 0.04025
R40326 VDD.n12018 VDD.n337 0.04025
R40327 VDD.n12019 VDD.n12018 0.04025
R40328 VDD.n12020 VDD.n12019 0.04025
R40329 VDD.n12020 VDD.n335 0.04025
R40330 VDD.n12024 VDD.n335 0.04025
R40331 VDD.n12025 VDD.n12024 0.04025
R40332 VDD.n12026 VDD.n12025 0.04025
R40333 VDD.n12026 VDD.n333 0.04025
R40334 VDD.n12030 VDD.n333 0.04025
R40335 VDD.n12031 VDD.n12030 0.04025
R40336 VDD.n12032 VDD.n12031 0.04025
R40337 VDD.n12032 VDD.n331 0.04025
R40338 VDD.n12036 VDD.n331 0.04025
R40339 VDD.n12037 VDD.n12036 0.04025
R40340 VDD.n12038 VDD.n12037 0.04025
R40341 VDD.n12038 VDD.n329 0.04025
R40342 VDD.n12042 VDD.n329 0.04025
R40343 VDD.n12043 VDD.n12042 0.04025
R40344 VDD.n12044 VDD.n12043 0.04025
R40345 VDD.n12044 VDD.n327 0.04025
R40346 VDD.n12048 VDD.n327 0.04025
R40347 VDD.n12049 VDD.n12048 0.04025
R40348 VDD.n12050 VDD.n12049 0.04025
R40349 VDD.n12050 VDD.n325 0.04025
R40350 VDD.n12054 VDD.n325 0.04025
R40351 VDD.n12055 VDD.n12054 0.04025
R40352 VDD.n12056 VDD.n12055 0.04025
R40353 VDD.n12056 VDD.n323 0.04025
R40354 VDD.n12060 VDD.n323 0.04025
R40355 VDD.n12061 VDD.n12060 0.04025
R40356 VDD.n12062 VDD.n12061 0.04025
R40357 VDD.n12062 VDD.n321 0.04025
R40358 VDD.n12066 VDD.n321 0.04025
R40359 VDD.n12067 VDD.n12066 0.04025
R40360 VDD.n12068 VDD.n12067 0.04025
R40361 VDD.n12068 VDD.n319 0.04025
R40362 VDD.n12072 VDD.n319 0.04025
R40363 VDD.n12073 VDD.n12072 0.04025
R40364 VDD.n12074 VDD.n12073 0.04025
R40365 VDD.n12074 VDD.n317 0.04025
R40366 VDD.n12078 VDD.n317 0.04025
R40367 VDD.n12079 VDD.n12078 0.04025
R40368 VDD.n12080 VDD.n12079 0.04025
R40369 VDD.n12080 VDD.n315 0.04025
R40370 VDD.n12084 VDD.n315 0.04025
R40371 VDD.n12085 VDD.n12084 0.04025
R40372 VDD.n12086 VDD.n12085 0.04025
R40373 VDD.n12086 VDD.n313 0.04025
R40374 VDD.n12090 VDD.n313 0.04025
R40375 VDD.n12091 VDD.n12090 0.04025
R40376 VDD.n12092 VDD.n12091 0.04025
R40377 VDD.n12092 VDD.n311 0.04025
R40378 VDD.n12096 VDD.n311 0.04025
R40379 VDD.n12097 VDD.n12096 0.04025
R40380 VDD.n12098 VDD.n12097 0.04025
R40381 VDD.n12098 VDD.n309 0.04025
R40382 VDD.n12102 VDD.n309 0.04025
R40383 VDD.n12103 VDD.n12102 0.04025
R40384 VDD.n12104 VDD.n12103 0.04025
R40385 VDD.n12104 VDD.n307 0.04025
R40386 VDD.n12108 VDD.n307 0.04025
R40387 VDD.n12109 VDD.n12108 0.04025
R40388 VDD.n12110 VDD.n12109 0.04025
R40389 VDD.n12110 VDD.n305 0.04025
R40390 VDD.n12114 VDD.n305 0.04025
R40391 VDD.n12115 VDD.n12114 0.04025
R40392 VDD.n12116 VDD.n12115 0.04025
R40393 VDD.n12116 VDD.n303 0.04025
R40394 VDD.n12120 VDD.n303 0.04025
R40395 VDD.n12121 VDD.n12120 0.04025
R40396 VDD.n12122 VDD.n12121 0.04025
R40397 VDD.n12122 VDD.n301 0.04025
R40398 VDD.n12126 VDD.n301 0.04025
R40399 VDD.n12127 VDD.n12126 0.04025
R40400 VDD.n12128 VDD.n12127 0.04025
R40401 VDD.n12128 VDD.n299 0.04025
R40402 VDD.n12132 VDD.n299 0.04025
R40403 VDD.n12133 VDD.n12132 0.04025
R40404 VDD.n12134 VDD.n12133 0.04025
R40405 VDD.n12134 VDD.n297 0.04025
R40406 VDD.n12138 VDD.n297 0.04025
R40407 VDD.n12139 VDD.n12138 0.04025
R40408 VDD.n12140 VDD.n12139 0.04025
R40409 VDD.n12140 VDD.n295 0.04025
R40410 VDD.n12144 VDD.n295 0.04025
R40411 VDD.n12145 VDD.n12144 0.04025
R40412 VDD.n12146 VDD.n12145 0.04025
R40413 VDD.n12146 VDD.n293 0.04025
R40414 VDD.n12150 VDD.n293 0.04025
R40415 VDD.n12151 VDD.n12150 0.04025
R40416 VDD.n12152 VDD.n12151 0.04025
R40417 VDD.n12152 VDD.n291 0.04025
R40418 VDD.n12156 VDD.n291 0.04025
R40419 VDD.n12157 VDD.n12156 0.04025
R40420 VDD.n12158 VDD.n12157 0.04025
R40421 VDD.n12158 VDD.n289 0.04025
R40422 VDD.n12162 VDD.n289 0.04025
R40423 VDD.n12163 VDD.n12162 0.04025
R40424 VDD.n12164 VDD.n12163 0.04025
R40425 VDD.n12164 VDD.n287 0.04025
R40426 VDD.n12168 VDD.n287 0.04025
R40427 VDD.n12169 VDD.n12168 0.04025
R40428 VDD.n12170 VDD.n12169 0.04025
R40429 VDD.n12170 VDD.n285 0.04025
R40430 VDD.n12174 VDD.n285 0.04025
R40431 VDD.n12175 VDD.n12174 0.04025
R40432 VDD.n12176 VDD.n12175 0.04025
R40433 VDD.n12176 VDD.n283 0.04025
R40434 VDD.n12180 VDD.n283 0.04025
R40435 VDD.n12181 VDD.n12180 0.04025
R40436 VDD.n12182 VDD.n12181 0.04025
R40437 VDD.n12182 VDD.n281 0.04025
R40438 VDD.n12186 VDD.n281 0.04025
R40439 VDD.n12187 VDD.n12186 0.04025
R40440 VDD.n12188 VDD.n12187 0.04025
R40441 VDD.n12188 VDD.n279 0.04025
R40442 VDD.n12192 VDD.n279 0.04025
R40443 VDD.n12193 VDD.n12192 0.04025
R40444 VDD.n12194 VDD.n12193 0.04025
R40445 VDD.n12194 VDD.n277 0.04025
R40446 VDD.n12198 VDD.n277 0.04025
R40447 VDD.n12199 VDD.n12198 0.04025
R40448 VDD.n12200 VDD.n12199 0.04025
R40449 VDD.n12200 VDD.n275 0.04025
R40450 VDD.n12204 VDD.n275 0.04025
R40451 VDD.n12205 VDD.n12204 0.04025
R40452 VDD.n12206 VDD.n12205 0.04025
R40453 VDD.n12206 VDD.n273 0.04025
R40454 VDD.n12210 VDD.n273 0.04025
R40455 VDD.n12211 VDD.n12210 0.04025
R40456 VDD.n12212 VDD.n12211 0.04025
R40457 VDD.n12212 VDD.n271 0.04025
R40458 VDD.n12216 VDD.n271 0.04025
R40459 VDD.n12217 VDD.n12216 0.04025
R40460 VDD.n12218 VDD.n12217 0.04025
R40461 VDD.n12218 VDD.n269 0.04025
R40462 VDD.n12222 VDD.n269 0.04025
R40463 VDD.n12223 VDD.n12222 0.04025
R40464 VDD.n12224 VDD.n12223 0.04025
R40465 VDD.n12224 VDD.n267 0.04025
R40466 VDD.n12228 VDD.n267 0.04025
R40467 VDD.n12229 VDD.n12228 0.04025
R40468 VDD.n12230 VDD.n12229 0.04025
R40469 VDD.n12230 VDD.n265 0.04025
R40470 VDD.n12234 VDD.n265 0.04025
R40471 VDD.n12235 VDD.n12234 0.04025
R40472 VDD.n12236 VDD.n12235 0.04025
R40473 VDD.n12236 VDD.n263 0.04025
R40474 VDD.n12240 VDD.n263 0.04025
R40475 VDD.n12241 VDD.n12240 0.04025
R40476 VDD.n12242 VDD.n12241 0.04025
R40477 VDD.n12242 VDD.n261 0.04025
R40478 VDD.n12246 VDD.n261 0.04025
R40479 VDD.n12247 VDD.n12246 0.04025
R40480 VDD.n12248 VDD.n12247 0.04025
R40481 VDD.n12248 VDD.n259 0.04025
R40482 VDD.n12252 VDD.n259 0.04025
R40483 VDD.n12253 VDD.n12252 0.04025
R40484 VDD.n12254 VDD.n12253 0.04025
R40485 VDD.n12254 VDD.n257 0.04025
R40486 VDD.n12258 VDD.n257 0.04025
R40487 VDD.n12259 VDD.n12258 0.04025
R40488 VDD.n12260 VDD.n12259 0.04025
R40489 VDD.n12260 VDD.n255 0.04025
R40490 VDD.n12264 VDD.n255 0.04025
R40491 VDD.n12265 VDD.n12264 0.04025
R40492 VDD.n12266 VDD.n12265 0.04025
R40493 VDD.n12266 VDD.n253 0.04025
R40494 VDD.n12270 VDD.n253 0.04025
R40495 VDD.n12271 VDD.n12270 0.04025
R40496 VDD.n12272 VDD.n12271 0.04025
R40497 VDD.n12272 VDD.n251 0.04025
R40498 VDD.n12276 VDD.n251 0.04025
R40499 VDD.n12277 VDD.n12276 0.04025
R40500 VDD.n12278 VDD.n12277 0.04025
R40501 VDD.n12278 VDD.n249 0.04025
R40502 VDD.n12282 VDD.n249 0.04025
R40503 VDD.n12283 VDD.n12282 0.04025
R40504 VDD.n12284 VDD.n12283 0.04025
R40505 VDD.n12284 VDD.n247 0.04025
R40506 VDD.n12288 VDD.n247 0.04025
R40507 VDD.n12289 VDD.n12288 0.04025
R40508 VDD.n12290 VDD.n12289 0.04025
R40509 VDD.n12290 VDD.n245 0.04025
R40510 VDD.n12294 VDD.n245 0.04025
R40511 VDD.n12295 VDD.n12294 0.04025
R40512 VDD.n12296 VDD.n12295 0.04025
R40513 VDD.n12296 VDD.n243 0.04025
R40514 VDD.n12300 VDD.n243 0.04025
R40515 VDD.n12301 VDD.n12300 0.04025
R40516 VDD.n12302 VDD.n12301 0.04025
R40517 VDD.n12302 VDD.n241 0.04025
R40518 VDD.n12306 VDD.n241 0.04025
R40519 VDD.n12307 VDD.n12306 0.04025
R40520 VDD.n12308 VDD.n12307 0.04025
R40521 VDD.n12308 VDD.n239 0.04025
R40522 VDD.n12312 VDD.n239 0.04025
R40523 VDD.n12313 VDD.n12312 0.04025
R40524 VDD.n12314 VDD.n12313 0.04025
R40525 VDD.n12314 VDD.n237 0.04025
R40526 VDD.n12318 VDD.n237 0.04025
R40527 VDD.n12319 VDD.n12318 0.04025
R40528 VDD.n12320 VDD.n12319 0.04025
R40529 VDD.n12320 VDD.n235 0.04025
R40530 VDD.n12324 VDD.n235 0.04025
R40531 VDD.n12325 VDD.n12324 0.04025
R40532 VDD.n12326 VDD.n12325 0.04025
R40533 VDD.n12326 VDD.n233 0.04025
R40534 VDD.n12330 VDD.n233 0.04025
R40535 VDD.n12331 VDD.n12330 0.04025
R40536 VDD.n12332 VDD.n12331 0.04025
R40537 VDD.n12332 VDD.n231 0.04025
R40538 VDD.n12336 VDD.n231 0.04025
R40539 VDD.n12337 VDD.n12336 0.04025
R40540 VDD.n12338 VDD.n12337 0.04025
R40541 VDD.n12338 VDD.n229 0.04025
R40542 VDD.n12342 VDD.n229 0.04025
R40543 VDD.n12343 VDD.n12342 0.04025
R40544 VDD.n12344 VDD.n12343 0.04025
R40545 VDD.n12344 VDD.n227 0.04025
R40546 VDD.n12348 VDD.n227 0.04025
R40547 VDD.n12349 VDD.n12348 0.04025
R40548 VDD.n12350 VDD.n12349 0.04025
R40549 VDD.n12350 VDD.n225 0.04025
R40550 VDD.n12354 VDD.n225 0.04025
R40551 VDD.n12355 VDD.n12354 0.04025
R40552 VDD.n12356 VDD.n12355 0.04025
R40553 VDD.n12356 VDD.n223 0.04025
R40554 VDD.n12360 VDD.n223 0.04025
R40555 VDD.n12361 VDD.n12360 0.04025
R40556 VDD.n12362 VDD.n12361 0.04025
R40557 VDD.n12362 VDD.n221 0.04025
R40558 VDD.n12366 VDD.n221 0.04025
R40559 VDD.n12367 VDD.n12366 0.04025
R40560 VDD.n12368 VDD.n12367 0.04025
R40561 VDD.n12368 VDD.n219 0.04025
R40562 VDD.n12372 VDD.n219 0.04025
R40563 VDD.n12373 VDD.n12372 0.04025
R40564 VDD.n12374 VDD.n12373 0.04025
R40565 VDD.n12374 VDD.n217 0.04025
R40566 VDD.n12378 VDD.n217 0.04025
R40567 VDD.n12379 VDD.n12378 0.04025
R40568 VDD.n12380 VDD.n12379 0.04025
R40569 VDD.n12380 VDD.n215 0.04025
R40570 VDD.n12384 VDD.n215 0.04025
R40571 VDD.n12385 VDD.n12384 0.04025
R40572 VDD.n12386 VDD.n12385 0.04025
R40573 VDD.n12386 VDD.n213 0.04025
R40574 VDD.n12390 VDD.n213 0.04025
R40575 VDD.n12391 VDD.n12390 0.04025
R40576 VDD.n12392 VDD.n12391 0.04025
R40577 VDD.n12392 VDD.n211 0.04025
R40578 VDD.n12396 VDD.n211 0.04025
R40579 VDD.n12397 VDD.n12396 0.04025
R40580 VDD.n12398 VDD.n12397 0.04025
R40581 VDD.n12398 VDD.n209 0.04025
R40582 VDD.n12402 VDD.n209 0.04025
R40583 VDD.n12403 VDD.n12402 0.04025
R40584 VDD.n12404 VDD.n12403 0.04025
R40585 VDD.n12404 VDD.n207 0.04025
R40586 VDD.n12408 VDD.n207 0.04025
R40587 VDD.n12409 VDD.n12408 0.04025
R40588 VDD.n12410 VDD.n12409 0.04025
R40589 VDD.n12410 VDD.n205 0.04025
R40590 VDD.n12414 VDD.n205 0.04025
R40591 VDD.n12415 VDD.n12414 0.04025
R40592 VDD.n12416 VDD.n12415 0.04025
R40593 VDD.n12416 VDD.n203 0.04025
R40594 VDD.n12420 VDD.n203 0.04025
R40595 VDD.n12421 VDD.n12420 0.04025
R40596 VDD.n12422 VDD.n12421 0.04025
R40597 VDD.n12422 VDD.n201 0.04025
R40598 VDD.n12426 VDD.n201 0.04025
R40599 VDD.n12427 VDD.n12426 0.04025
R40600 VDD.n12428 VDD.n12427 0.04025
R40601 VDD.n12428 VDD.n199 0.04025
R40602 VDD.n12432 VDD.n199 0.04025
R40603 VDD.n12433 VDD.n12432 0.04025
R40604 VDD.n12434 VDD.n12433 0.04025
R40605 VDD.n12434 VDD.n197 0.04025
R40606 VDD.n12438 VDD.n197 0.04025
R40607 VDD.n12439 VDD.n12438 0.04025
R40608 VDD.n12440 VDD.n12439 0.04025
R40609 VDD.n7843 VDD.n7842 0.0395167
R40610 VDD.n2173 VDD.n2172 0.0394276
R40611 VDD.n6875 VDD.n2390 0.0392688
R40612 VDD.n8052 VDD.n8051 0.0387235
R40613 VDD.n8048 VDD.n8047 0.0383
R40614 VDD.n9137 VDD.n9136 0.0382419
R40615 VDD.n9126 VDD.n9125 0.0382419
R40616 VDD.n12565 VDD.n12563 0.0382419
R40617 VDD.n12577 VDD.n12576 0.0382419
R40618 VDD.n10148 VDD.n10147 0.037625
R40619 VDD.n8052 VDD.n2148 0.0373471
R40620 VDD.n7942 VDD.n7854 0.0371353
R40621 VDD.n1564 VDD.n1563 0.0370902
R40622 VDD.n1542 VDD.n1541 0.0370902
R40623 VDD.n1640 VDD.n771 0.0370902
R40624 VDD.n1529 VDD.n1528 0.0370902
R40625 VDD.n7912 VDD.n7911 0.0369637
R40626 VDD.n7943 VDD.n7942 0.0369235
R40627 VDD.n7912 VDD.n7863 0.0367529
R40628 VDD.n12567 VDD.n12566 0.0364748
R40629 VDD.n12574 VDD.n12573 0.0364748
R40630 VDD.n9184 VDD.n9183 0.0363759
R40631 VDD.n5369 VDD.n5368 0.0360345
R40632 VDD.n6372 VDD.n5375 0.0360345
R40633 VDD.n6368 VDD.n6367 0.0360345
R40634 VDD.n5944 VDD.n5943 0.0360345
R40635 VDD.n2366 VDD.n2365 0.0360345
R40636 VDD.n7135 VDD.n2316 0.0360345
R40637 VDD.n7131 VDD.n7130 0.0360345
R40638 VDD.n7044 VDD.n7043 0.0360345
R40639 VDD.n7864 VDD.n2146 0.0359624
R40640 VDD.n12641 VDD.n12638 0.0359286
R40641 VDD.n1003 VDD.n957 0.0359286
R40642 VDD.n1755 VDD.n1754 0.0359286
R40643 VDD.n9135 VDD.n9134 0.0357174
R40644 VDD.n6024 VDD.n5299 0.0347688
R40645 VDD.n6174 VDD.n6171 0.0347688
R40646 VDD.n6412 VDD.n5299 0.0347688
R40647 VDD.n8011 VDD.n8010 0.0347688
R40648 VDD.n2403 VDD.n2402 0.0347688
R40649 VDD.n2402 VDD.n2396 0.0347688
R40650 VDD.n8133 VDD.n8132 0.0346711
R40651 VDD.n8134 VDD.n8133 0.0346711
R40652 VDD.n8134 VDD.n2090 0.0346711
R40653 VDD.n8136 VDD.n2090 0.0346711
R40654 VDD.n8139 VDD.n8138 0.0346711
R40655 VDD.n8162 VDD.n8139 0.0346711
R40656 VDD.n8112 VDD.n8111 0.0346711
R40657 VDD.n8113 VDD.n8112 0.0346711
R40658 VDD.n8113 VDD.n2092 0.0346711
R40659 VDD.n8115 VDD.n2092 0.0346711
R40660 VDD.n8118 VDD.n8117 0.0346711
R40661 VDD.n8119 VDD.n8118 0.0346711
R40662 VDD.n8119 VDD.n2091 0.0346711
R40663 VDD.n8121 VDD.n2091 0.0346711
R40664 VDD.n8100 VDD.n8099 0.0346711
R40665 VDD.n8101 VDD.n8100 0.0346711
R40666 VDD.n8101 VDD.n2103 0.0346711
R40667 VDD.n8103 VDD.n2103 0.0346711
R40668 VDD.n8106 VDD.n8105 0.0346711
R40669 VDD.n8107 VDD.n8106 0.0346711
R40670 VDD.n8107 VDD.n2102 0.0346711
R40671 VDD.n8109 VDD.n2102 0.0346711
R40672 VDD.n5584 VDD.n5551 0.0346711
R40673 VDD.n5582 VDD.n5551 0.0346711
R40674 VDD.n5582 VDD.n5581 0.0346711
R40675 VDD.n5581 VDD.n5580 0.0346711
R40676 VDD.n5578 VDD.n5552 0.0346711
R40677 VDD.n5576 VDD.n5552 0.0346711
R40678 VDD.n5605 VDD.n5549 0.0346711
R40679 VDD.n5603 VDD.n5549 0.0346711
R40680 VDD.n5603 VDD.n5602 0.0346711
R40681 VDD.n5602 VDD.n5601 0.0346711
R40682 VDD.n5599 VDD.n5550 0.0346711
R40683 VDD.n5597 VDD.n5550 0.0346711
R40684 VDD.n5597 VDD.n5596 0.0346711
R40685 VDD.n5596 VDD.n5595 0.0346711
R40686 VDD.n5626 VDD.n5547 0.0346711
R40687 VDD.n5624 VDD.n5547 0.0346711
R40688 VDD.n5624 VDD.n5623 0.0346711
R40689 VDD.n5623 VDD.n5622 0.0346711
R40690 VDD.n5620 VDD.n5548 0.0346711
R40691 VDD.n5618 VDD.n5548 0.0346711
R40692 VDD.n5618 VDD.n5617 0.0346711
R40693 VDD.n5617 VDD.n5616 0.0346711
R40694 VDD.n5666 VDD.n5542 0.0346711
R40695 VDD.n5664 VDD.n5542 0.0346711
R40696 VDD.n5664 VDD.n5663 0.0346711
R40697 VDD.n5663 VDD.n5662 0.0346711
R40698 VDD.n5660 VDD.n5543 0.0346711
R40699 VDD.n5658 VDD.n5543 0.0346711
R40700 VDD.n5867 VDD.n5866 0.0346711
R40701 VDD.n5868 VDD.n5867 0.0346711
R40702 VDD.n5868 VDD.n5668 0.0346711
R40703 VDD.n5870 VDD.n5668 0.0346711
R40704 VDD.n5873 VDD.n5872 0.0346711
R40705 VDD.n5874 VDD.n5873 0.0346711
R40706 VDD.n5874 VDD.n5667 0.0346711
R40707 VDD.n5876 VDD.n5667 0.0346711
R40708 VDD.n5855 VDD.n5854 0.0346711
R40709 VDD.n5856 VDD.n5855 0.0346711
R40710 VDD.n5856 VDD.n5679 0.0346711
R40711 VDD.n5858 VDD.n5679 0.0346711
R40712 VDD.n5861 VDD.n5860 0.0346711
R40713 VDD.n5862 VDD.n5861 0.0346711
R40714 VDD.n5862 VDD.n5678 0.0346711
R40715 VDD.n5864 VDD.n5678 0.0346711
R40716 VDD.n5812 VDD.n5811 0.0346711
R40717 VDD.n5813 VDD.n5812 0.0346711
R40718 VDD.n5813 VDD.n5681 0.0346711
R40719 VDD.n5815 VDD.n5681 0.0346711
R40720 VDD.n5818 VDD.n5817 0.0346711
R40721 VDD.n5841 VDD.n5818 0.0346711
R40722 VDD.n5800 VDD.n5799 0.0346711
R40723 VDD.n5801 VDD.n5800 0.0346711
R40724 VDD.n5801 VDD.n5692 0.0346711
R40725 VDD.n5803 VDD.n5692 0.0346711
R40726 VDD.n5806 VDD.n5805 0.0346711
R40727 VDD.n5807 VDD.n5806 0.0346711
R40728 VDD.n5807 VDD.n5691 0.0346711
R40729 VDD.n5809 VDD.n5691 0.0346711
R40730 VDD.n5779 VDD.n5778 0.0346711
R40731 VDD.n5780 VDD.n5779 0.0346711
R40732 VDD.n5780 VDD.n5694 0.0346711
R40733 VDD.n5782 VDD.n5694 0.0346711
R40734 VDD.n5785 VDD.n5784 0.0346711
R40735 VDD.n5786 VDD.n5785 0.0346711
R40736 VDD.n5786 VDD.n5693 0.0346711
R40737 VDD.n5788 VDD.n5693 0.0346711
R40738 VDD.n5745 VDD.n5744 0.0346711
R40739 VDD.n5746 VDD.n5745 0.0346711
R40740 VDD.n5746 VDD.n5705 0.0346711
R40741 VDD.n5748 VDD.n5705 0.0346711
R40742 VDD.n5751 VDD.n5750 0.0346711
R40743 VDD.n5774 VDD.n5751 0.0346711
R40744 VDD.n5724 VDD.n5723 0.0346711
R40745 VDD.n5725 VDD.n5724 0.0346711
R40746 VDD.n5725 VDD.n5707 0.0346711
R40747 VDD.n5727 VDD.n5707 0.0346711
R40748 VDD.n5730 VDD.n5729 0.0346711
R40749 VDD.n5731 VDD.n5730 0.0346711
R40750 VDD.n5731 VDD.n5706 0.0346711
R40751 VDD.n5733 VDD.n5706 0.0346711
R40752 VDD.n11036 VDD.n1769 0.0346711
R40753 VDD.n11034 VDD.n1769 0.0346711
R40754 VDD.n11034 VDD.n11033 0.0346711
R40755 VDD.n11033 VDD.n11032 0.0346711
R40756 VDD.n5718 VDD.n1770 0.0346711
R40757 VDD.n5719 VDD.n5718 0.0346711
R40758 VDD.n5719 VDD.n5717 0.0346711
R40759 VDD.n5721 VDD.n5717 0.0346711
R40760 VDD.n8975 VDD.n8971 0.0346711
R40761 VDD.n8973 VDD.n8971 0.0346711
R40762 VDD.n8973 VDD.n8972 0.0346711
R40763 VDD.n8972 VDD.n8490 0.0346711
R40764 VDD.n9039 VDD.n9038 0.0346711
R40765 VDD.n9040 VDD.n9039 0.0346711
R40766 VDD.n9040 VDD.n8489 0.0346711
R40767 VDD.n9042 VDD.n8489 0.0346711
R40768 VDD.n8948 VDD.n8947 0.0346711
R40769 VDD.n8949 VDD.n8948 0.0346711
R40770 VDD.n8949 VDD.n8502 0.0346711
R40771 VDD.n8951 VDD.n8502 0.0346711
R40772 VDD.n9007 VDD.n8952 0.0346711
R40773 VDD.n9005 VDD.n8952 0.0346711
R40774 VDD.n8848 VDD.n8844 0.0346711
R40775 VDD.n8846 VDD.n8844 0.0346711
R40776 VDD.n8846 VDD.n8845 0.0346711
R40777 VDD.n8845 VDD.n8507 0.0346711
R40778 VDD.n8942 VDD.n8941 0.0346711
R40779 VDD.n8943 VDD.n8942 0.0346711
R40780 VDD.n8943 VDD.n8506 0.0346711
R40781 VDD.n8945 VDD.n8506 0.0346711
R40782 VDD.n8839 VDD.n8838 0.0346711
R40783 VDD.n8840 VDD.n8839 0.0346711
R40784 VDD.n8840 VDD.n8521 0.0346711
R40785 VDD.n8842 VDD.n8521 0.0346711
R40786 VDD.n8876 VDD.n8843 0.0346711
R40787 VDD.n8874 VDD.n8843 0.0346711
R40788 VDD.n8874 VDD.n8873 0.0346711
R40789 VDD.n8873 VDD.n8872 0.0346711
R40790 VDD.n8547 VDD.n8543 0.0346711
R40791 VDD.n8545 VDD.n8543 0.0346711
R40792 VDD.n8545 VDD.n8544 0.0346711
R40793 VDD.n8544 VDD.n8526 0.0346711
R40794 VDD.n8811 VDD.n8810 0.0346711
R40795 VDD.n8834 VDD.n8811 0.0346711
R40796 VDD.n8550 VDD.n184 0.0346711
R40797 VDD.n8551 VDD.n8550 0.0346711
R40798 VDD.n8551 VDD.n8549 0.0346711
R40799 VDD.n8553 VDD.n8549 0.0346711
R40800 VDD.n8556 VDD.n8555 0.0346711
R40801 VDD.n8557 VDD.n8556 0.0346711
R40802 VDD.n8557 VDD.n8548 0.0346711
R40803 VDD.n8559 VDD.n8548 0.0346711
R40804 VDD.n171 VDD.n170 0.0346711
R40805 VDD.n172 VDD.n171 0.0346711
R40806 VDD.n172 VDD.n125 0.0346711
R40807 VDD.n174 VDD.n125 0.0346711
R40808 VDD.n187 VDD.n186 0.0346711
R40809 VDD.n188 VDD.n187 0.0346711
R40810 VDD.n188 VDD.n185 0.0346711
R40811 VDD.n190 VDD.n185 0.0346711
R40812 VDD.n9092 VDD.n8470 0.0346711
R40813 VDD.n9093 VDD.n9092 0.0346711
R40814 VDD.n9093 VDD.n9091 0.0346711
R40815 VDD.n9095 VDD.n9091 0.0346711
R40816 VDD.n9098 VDD.n9097 0.0346711
R40817 VDD.n9121 VDD.n9098 0.0346711
R40818 VDD.n8488 VDD.n8484 0.0346711
R40819 VDD.n8486 VDD.n8484 0.0346711
R40820 VDD.n8486 VDD.n8485 0.0346711
R40821 VDD.n8485 VDD.n8472 0.0346711
R40822 VDD.n9163 VDD.n9162 0.0346711
R40823 VDD.n9164 VDD.n9163 0.0346711
R40824 VDD.n9164 VDD.n8471 0.0346711
R40825 VDD.n9166 VDD.n8471 0.0346711
R40826 VDD.n137 VDD.n106 0.0346711
R40827 VDD.n138 VDD.n137 0.0346711
R40828 VDD.n138 VDD.n136 0.0346711
R40829 VDD.n140 VDD.n136 0.0346711
R40830 VDD.n143 VDD.n142 0.0346711
R40831 VDD.n166 VDD.n143 0.0346711
R40832 VDD.n12498 VDD.n104 0.0346711
R40833 VDD.n12496 VDD.n104 0.0346711
R40834 VDD.n12496 VDD.n12495 0.0346711
R40835 VDD.n12495 VDD.n12494 0.0346711
R40836 VDD.n12492 VDD.n105 0.0346711
R40837 VDD.n12490 VDD.n105 0.0346711
R40838 VDD.n12490 VDD.n12489 0.0346711
R40839 VDD.n12489 VDD.n12488 0.0346711
R40840 VDD.n91 VDD.n90 0.0346711
R40841 VDD.n92 VDD.n91 0.0346711
R40842 VDD.n92 VDD.n45 0.0346711
R40843 VDD.n94 VDD.n45 0.0346711
R40844 VDD.n12501 VDD.n12500 0.0346711
R40845 VDD.n12502 VDD.n12501 0.0346711
R40846 VDD.n12502 VDD.n12499 0.0346711
R40847 VDD.n12504 VDD.n12499 0.0346711
R40848 VDD.n48 VDD.n26 0.0346711
R40849 VDD.n49 VDD.n48 0.0346711
R40850 VDD.n49 VDD.n47 0.0346711
R40851 VDD.n51 VDD.n47 0.0346711
R40852 VDD.n54 VDD.n53 0.0346711
R40853 VDD.n77 VDD.n54 0.0346711
R40854 VDD.n12554 VDD.n24 0.0346711
R40855 VDD.n12552 VDD.n24 0.0346711
R40856 VDD.n12552 VDD.n12551 0.0346711
R40857 VDD.n12551 VDD.n12550 0.0346711
R40858 VDD.n12548 VDD.n25 0.0346711
R40859 VDD.n12546 VDD.n25 0.0346711
R40860 VDD.n12546 VDD.n12545 0.0346711
R40861 VDD.n12545 VDD.n12544 0.0346711
R40862 VDD.n12588 VDD.n12587 0.0346711
R40863 VDD.n12589 VDD.n12588 0.0346711
R40864 VDD.n12589 VDD.n12556 0.0346711
R40865 VDD.n12591 VDD.n12556 0.0346711
R40866 VDD.n12595 VDD.n12594 0.0346711
R40867 VDD.n12596 VDD.n12595 0.0346711
R40868 VDD.n12596 VDD.n12555 0.0346711
R40869 VDD.n12598 VDD.n12555 0.0346711
R40870 VDD.n12580 VDD.n12579 0.0345
R40871 VDD.n11129 VDD.n638 0.0345
R40872 VDD.n1763 VDD.n674 0.0345
R40873 VDD.n6325 VDD.n6324 0.0345
R40874 VDD.n6014 VDD.n6011 0.0345
R40875 VDD.n5538 VDD.n5537 0.0345
R40876 VDD.n5886 VDD.n5880 0.0345
R40877 VDD.n5911 VDD.n5910 0.0345
R40878 VDD.n8088 VDD.n1996 0.0345
R40879 VDD.n8090 VDD.n2118 0.0345
R40880 VDD.n12632 VDD.n12631 0.0345
R40881 VDD.n12635 VDD.n3 0.0345
R40882 VDD.n1000 VDD.n953 0.0345
R40883 VDD.n1760 VDD.n1759 0.0345
R40884 VDD.n6024 VDD.n6022 0.0341759
R40885 VDD.n6036 VDD.n6023 0.0341759
R40886 VDD.n6033 VDD.n6023 0.0341759
R40887 VDD.n6033 VDD.n6032 0.0341759
R40888 VDD.n6032 VDD.n6031 0.0341759
R40889 VDD.n6031 VDD.n6025 0.0341759
R40890 VDD.n6029 VDD.n6025 0.0341759
R40891 VDD.n6028 VDD.n6026 0.0341759
R40892 VDD.n6026 VDD.n5283 0.0341759
R40893 VDD.n6574 VDD.n6573 0.0341759
R40894 VDD.n6573 VDD.n5284 0.0341759
R40895 VDD.n6571 VDD.n5284 0.0341759
R40896 VDD.n6570 VDD.n5285 0.0341759
R40897 VDD.n6568 VDD.n5285 0.0341759
R40898 VDD.n6568 VDD.n6567 0.0341759
R40899 VDD.n6567 VDD.n6566 0.0341759
R40900 VDD.n6566 VDD.n5286 0.0341759
R40901 VDD.n6563 VDD.n5286 0.0341759
R40902 VDD.n6171 VDD.n6018 0.0341759
R40903 VDD.n6169 VDD.n6168 0.0341759
R40904 VDD.n6168 VDD.n6167 0.0341759
R40905 VDD.n6167 VDD.n6158 0.0341759
R40906 VDD.n6164 VDD.n6158 0.0341759
R40907 VDD.n6164 VDD.n6163 0.0341759
R40908 VDD.n6163 VDD.n6162 0.0341759
R40909 VDD.n6161 VDD.n6159 0.0341759
R40910 VDD.n6159 VDD.n5302 0.0341759
R40911 VDD.n6400 VDD.n6399 0.0341759
R40912 VDD.n6400 VDD.n5301 0.0341759
R40913 VDD.n6402 VDD.n5301 0.0341759
R40914 VDD.n6404 VDD.n6403 0.0341759
R40915 VDD.n6405 VDD.n6404 0.0341759
R40916 VDD.n6405 VDD.n5300 0.0341759
R40917 VDD.n6408 VDD.n5300 0.0341759
R40918 VDD.n6409 VDD.n6408 0.0341759
R40919 VDD.n6410 VDD.n6409 0.0341759
R40920 VDD.n8010 VDD.n2166 0.0341759
R40921 VDD.n8008 VDD.n2166 0.0341759
R40922 VDD.n8008 VDD.n8007 0.0341759
R40923 VDD.n8007 VDD.n8006 0.0341759
R40924 VDD.n8006 VDD.n2167 0.0341759
R40925 VDD.n8003 VDD.n2167 0.0341759
R40926 VDD.n8003 VDD.n8002 0.0341759
R40927 VDD.n8002 VDD.n8001 0.0341759
R40928 VDD.n8000 VDD.n2168 0.0341759
R40929 VDD.n7998 VDD.n2168 0.0341759
R40930 VDD.n2186 VDD.n2185 0.0341759
R40931 VDD.n2185 VDD.n2169 0.0341759
R40932 VDD.n2183 VDD.n2169 0.0341759
R40933 VDD.n2182 VDD.n2170 0.0341759
R40934 VDD.n2180 VDD.n2170 0.0341759
R40935 VDD.n2180 VDD.n2179 0.0341759
R40936 VDD.n2179 VDD.n2178 0.0341759
R40937 VDD.n2178 VDD.n2171 0.0341759
R40938 VDD.n2175 VDD.n2171 0.0341759
R40939 VDD.n2175 VDD.n2174 0.0341759
R40940 VDD.n2174 VDD.n2173 0.0341759
R40941 VDD.n2404 VDD.n2403 0.0341759
R40942 VDD.n6850 VDD.n2395 0.0341759
R40943 VDD.n6853 VDD.n2395 0.0341759
R40944 VDD.n6854 VDD.n6853 0.0341759
R40945 VDD.n6855 VDD.n6854 0.0341759
R40946 VDD.n6855 VDD.n2394 0.0341759
R40947 VDD.n6857 VDD.n2394 0.0341759
R40948 VDD.n6858 VDD.n2393 0.0341759
R40949 VDD.n6860 VDD.n2393 0.0341759
R40950 VDD.n6863 VDD.n6862 0.0341759
R40951 VDD.n6863 VDD.n2392 0.0341759
R40952 VDD.n6865 VDD.n2392 0.0341759
R40953 VDD.n6867 VDD.n6866 0.0341759
R40954 VDD.n6868 VDD.n6867 0.0341759
R40955 VDD.n6868 VDD.n2391 0.0341759
R40956 VDD.n6871 VDD.n2391 0.0341759
R40957 VDD.n6872 VDD.n6871 0.0341759
R40958 VDD.n6873 VDD.n6872 0.0341759
R40959 VDD.n6726 VDD.n2407 0.0341759
R40960 VDD.n6723 VDD.n2407 0.0341759
R40961 VDD.n6723 VDD.n6722 0.0341759
R40962 VDD.n6722 VDD.n6721 0.0341759
R40963 VDD.n6721 VDD.n6715 0.0341759
R40964 VDD.n6719 VDD.n6715 0.0341759
R40965 VDD.n6718 VDD.n6716 0.0341759
R40966 VDD.n6716 VDD.n2370 0.0341759
R40967 VDD.n7037 VDD.n7036 0.0341759
R40968 VDD.n7036 VDD.n2371 0.0341759
R40969 VDD.n7034 VDD.n2371 0.0341759
R40970 VDD.n7033 VDD.n2372 0.0341759
R40971 VDD.n7031 VDD.n2372 0.0341759
R40972 VDD.n7031 VDD.n7030 0.0341759
R40973 VDD.n7030 VDD.n7029 0.0341759
R40974 VDD.n7029 VDD.n2373 0.0341759
R40975 VDD.n7026 VDD.n2373 0.0341759
R40976 VDD.n5950 VDD.n5936 0.0337609
R40977 VDD.n6624 VDD.n6593 0.0337609
R40978 VDD.n5980 VDD.n5978 0.0337609
R40979 VDD.n5951 VDD.n5950 0.0337609
R40980 VDD.n6624 VDD.n6623 0.0337609
R40981 VDD.n5936 VDD.n5922 0.0331854
R40982 VDD.n5934 VDD.n5922 0.0331854
R40983 VDD.n5934 VDD.n5933 0.0331854
R40984 VDD.n5933 VDD.n5932 0.0331854
R40985 VDD.n5932 VDD.n5923 0.0331854
R40986 VDD.n5929 VDD.n5923 0.0331854
R40987 VDD.n5929 VDD.n5928 0.0331854
R40988 VDD.n5928 VDD.n5927 0.0331854
R40989 VDD.n5926 VDD.n5924 0.0331854
R40990 VDD.n5924 VDD.n5274 0.0331854
R40991 VDD.n6581 VDD.n6580 0.0331854
R40992 VDD.n6581 VDD.n5273 0.0331854
R40993 VDD.n6583 VDD.n5273 0.0331854
R40994 VDD.n6585 VDD.n6584 0.0331854
R40995 VDD.n6586 VDD.n6585 0.0331854
R40996 VDD.n6586 VDD.n5272 0.0331854
R40997 VDD.n6589 VDD.n5272 0.0331854
R40998 VDD.n6590 VDD.n6589 0.0331854
R40999 VDD.n6591 VDD.n6590 0.0331854
R41000 VDD.n6591 VDD.n5271 0.0331854
R41001 VDD.n6593 VDD.n5271 0.0331854
R41002 VDD.n5978 VDD.n5916 0.0331854
R41003 VDD.n5976 VDD.n5916 0.0331854
R41004 VDD.n5976 VDD.n5975 0.0331854
R41005 VDD.n5975 VDD.n5974 0.0331854
R41006 VDD.n5974 VDD.n5917 0.0331854
R41007 VDD.n5971 VDD.n5917 0.0331854
R41008 VDD.n5971 VDD.n5970 0.0331854
R41009 VDD.n5970 VDD.n5969 0.0331854
R41010 VDD.n5968 VDD.n5918 0.0331854
R41011 VDD.n5966 VDD.n5918 0.0331854
R41012 VDD.n5964 VDD.n5963 0.0331854
R41013 VDD.n5963 VDD.n5919 0.0331854
R41014 VDD.n5961 VDD.n5919 0.0331854
R41015 VDD.n5960 VDD.n5920 0.0331854
R41016 VDD.n5958 VDD.n5920 0.0331854
R41017 VDD.n5958 VDD.n5957 0.0331854
R41018 VDD.n5957 VDD.n5956 0.0331854
R41019 VDD.n5956 VDD.n5921 0.0331854
R41020 VDD.n5953 VDD.n5921 0.0331854
R41021 VDD.n5953 VDD.n5952 0.0331854
R41022 VDD.n5952 VDD.n5951 0.0331854
R41023 VDD.n6623 VDD.n6594 0.0331854
R41024 VDD.n6621 VDD.n6594 0.0331854
R41025 VDD.n6621 VDD.n6620 0.0331854
R41026 VDD.n6620 VDD.n6619 0.0331854
R41027 VDD.n6619 VDD.n6595 0.0331854
R41028 VDD.n6616 VDD.n6595 0.0331854
R41029 VDD.n6616 VDD.n6615 0.0331854
R41030 VDD.n6615 VDD.n6614 0.0331854
R41031 VDD.n6613 VDD.n6596 0.0331854
R41032 VDD.n6611 VDD.n6596 0.0331854
R41033 VDD.n6609 VDD.n6608 0.0331854
R41034 VDD.n6608 VDD.n6597 0.0331854
R41035 VDD.n6606 VDD.n6597 0.0331854
R41036 VDD.n6605 VDD.n6598 0.0331854
R41037 VDD.n6603 VDD.n6598 0.0331854
R41038 VDD.n6603 VDD.n6602 0.0331854
R41039 VDD.n6602 VDD.n6601 0.0331854
R41040 VDD.n7845 VDD.n2208 0.0331854
R41041 VDD.n7845 VDD.n7844 0.0331854
R41042 VDD.n7844 VDD.n7843 0.0331854
R41043 VDD.n1664 VDD.n1663 0.0331792
R41044 VDD.n1571 VDD.n1570 0.0331792
R41045 VDD.n1573 VDD.n1572 0.0331792
R41046 VDD.n1575 VDD.n1574 0.0331792
R41047 VDD.n1590 VDD.n1589 0.0331792
R41048 VDD.n1588 VDD.n1587 0.0331792
R41049 VDD.n1586 VDD.n1585 0.0331792
R41050 VDD.n1584 VDD.n1583 0.0331792
R41051 VDD.n1670 VDD.n1669 0.0331792
R41052 VDD.n1668 VDD.n1667 0.0331792
R41053 VDD.n1666 VDD.n1665 0.0331792
R41054 VDD.n7683 VDD.n7177 0.0328372
R41055 VDD.n6303 VDD.n6302 0.0325255
R41056 VDD.n6307 VDD.n6306 0.0325255
R41057 VDD.n5986 VDD.n5985 0.0325255
R41058 VDD.n6316 VDD.n6315 0.0325255
R41059 VDD.n6193 VDD.n6192 0.0325255
R41060 VDD.n6198 VDD.n6197 0.0325255
R41061 VDD.n6183 VDD.n6182 0.0325255
R41062 VDD.n6188 VDD.n6187 0.0325255
R41063 VDD.n6029 VDD.n6028 0.0325158
R41064 VDD.n6571 VDD.n6570 0.0325158
R41065 VDD.n6162 VDD.n6161 0.0325158
R41066 VDD.n6403 VDD.n6402 0.0325158
R41067 VDD.n8001 VDD.n8000 0.0325158
R41068 VDD.n2183 VDD.n2182 0.0325158
R41069 VDD.n6858 VDD.n6857 0.0325158
R41070 VDD.n6866 VDD.n6865 0.0325158
R41071 VDD.n6719 VDD.n6718 0.0325158
R41072 VDD.n7034 VDD.n7033 0.0325158
R41073 VDD.n1660 VDD.n1659 0.0324891
R41074 VDD.n1645 VDD.n1644 0.0324891
R41075 VDD.n7946 VDD.n7945 0.0320529
R41076 VDD.n7944 VDD.n7943 0.0320529
R41077 VDD.n7887 VDD.n7854 0.0320529
R41078 VDD.n7888 VDD.n2148 0.0320529
R41079 VDD.n8051 VDD.n8050 0.0320529
R41080 VDD.n8049 VDD.n8048 0.0320529
R41081 VDD.n2172 VDD.n2149 0.0320529
R41082 VDD.n1663 VDD.n753 0.0320159
R41083 VDD.n1662 VDD.n753 0.0320159
R41084 VDD.n1569 VDD.n1509 0.0320159
R41085 VDD.n1570 VDD.n1509 0.0320159
R41086 VDD.n1571 VDD.n1508 0.0320159
R41087 VDD.n1572 VDD.n1508 0.0320159
R41088 VDD.n1575 VDD.n1505 0.0320159
R41089 VDD.n1576 VDD.n1505 0.0320159
R41090 VDD.n1591 VDD.n1577 0.0320159
R41091 VDD.n1590 VDD.n1577 0.0320159
R41092 VDD.n1589 VDD.n1578 0.0320159
R41093 VDD.n1588 VDD.n1578 0.0320159
R41094 VDD.n1587 VDD.n1579 0.0320159
R41095 VDD.n1586 VDD.n1579 0.0320159
R41096 VDD.n1585 VDD.n1580 0.0320159
R41097 VDD.n1584 VDD.n1580 0.0320159
R41098 VDD.n1583 VDD.n1581 0.0320159
R41099 VDD.n1582 VDD.n1581 0.0320159
R41100 VDD.n1671 VDD.n748 0.0320159
R41101 VDD.n1670 VDD.n748 0.0320159
R41102 VDD.n1669 VDD.n749 0.0320159
R41103 VDD.n1668 VDD.n749 0.0320159
R41104 VDD.n1667 VDD.n750 0.0320159
R41105 VDD.n1666 VDD.n750 0.0320159
R41106 VDD.n6686 VDD.n6685 0.0319413
R41107 VDD.n6685 VDD.n6641 0.0319104
R41108 VDD.n7861 VDD.n2204 0.0319052
R41109 VDD.n7863 VDD.n7862 0.0319052
R41110 VDD.n7911 VDD.n7910 0.0319052
R41111 VDD.n7177 VDD.n7176 0.031686
R41112 VDD.n2296 VDD.n2295 0.031686
R41113 VDD.n2294 VDD.n2209 0.031686
R41114 VDD.n7838 VDD.n7837 0.031686
R41115 VDD.n7840 VDD.n7839 0.031686
R41116 VDD.n7842 VDD.n7841 0.031686
R41117 VDD.n2390 VDD.n2389 0.031686
R41118 VDD.n2388 VDD.n2387 0.031686
R41119 VDD.n2386 VDD.n2239 0.031686
R41120 VDD.n7831 VDD.n7830 0.031686
R41121 VDD.n7829 VDD.n7828 0.031686
R41122 VDD.n7826 VDD.n7825 0.031686
R41123 VDD.n7824 VDD.n7823 0.031686
R41124 VDD.n9134 VDD.n9127 0.0316781
R41125 VDD.n5927 VDD.n5926 0.0315742
R41126 VDD.n6584 VDD.n6583 0.0315742
R41127 VDD.n5969 VDD.n5968 0.0315742
R41128 VDD.n5961 VDD.n5960 0.0315742
R41129 VDD.n6614 VDD.n6613 0.0315742
R41130 VDD.n6606 VDD.n6605 0.0315742
R41131 VDD.n6711 VDD.n6710 0.0315707
R41132 VDD.n6702 VDD.n6701 0.0315707
R41133 VDD.n6697 VDD.n6696 0.0315707
R41134 VDD.n6688 VDD.n6687 0.0315707
R41135 VDD.n6640 VDD.n6639 0.0315707
R41136 VDD.n5437 VDD.n5436 0.0315707
R41137 VDD.n5442 VDD.n5441 0.0315707
R41138 VDD.n6627 VDD.n6626 0.0315707
R41139 VDD.n5368 VDD.n5367 0.0313793
R41140 VDD.n6373 VDD.n6372 0.0313793
R41141 VDD.n6368 VDD.n5377 0.0313793
R41142 VDD.n5943 VDD.n5941 0.0313793
R41143 VDD.n2366 VDD.n2360 0.0313793
R41144 VDD.n7136 VDD.n7135 0.0313793
R41145 VDD.n7131 VDD.n2320 0.0313793
R41146 VDD.n7043 VDD.n2347 0.0313793
R41147 VDD.n7309 VDD.n7302 0.0312734
R41148 VDD.n2208 VDD.n2206 0.0311937
R41149 VDD.n9124 VDD.n9123 0.0308128
R41150 VDD.n9139 VDD.n9138 0.0307932
R41151 VDD.n2970 VDD.n2969 0.0305815
R41152 VDD.n6575 VDD.n5283 0.0303814
R41153 VDD.n6398 VDD.n5302 0.0303814
R41154 VDD.n6861 VDD.n6860 0.0303814
R41155 VDD.n7038 VDD.n2370 0.0303814
R41156 VDD.n5288 VDD.n2410 0.0302628
R41157 VDD.n6413 VDD.n6412 0.0302628
R41158 VDD.n6876 VDD.n6875 0.0302628
R41159 VDD.n2396 VDD.n2375 0.0302628
R41160 VDD.n8162 VDD.n8161 0.0302193
R41161 VDD.n5576 VDD.n5575 0.0302193
R41162 VDD.n5658 VDD.n5657 0.0302193
R41163 VDD.n5841 VDD.n5840 0.0302193
R41164 VDD.n5774 VDD.n5773 0.0302193
R41165 VDD.n9005 VDD.n9004 0.0302193
R41166 VDD.n8834 VDD.n8833 0.0302193
R41167 VDD.n9121 VDD.n9120 0.0302193
R41168 VDD.n166 VDD.n165 0.0302193
R41169 VDD.n77 VDD.n76 0.0302193
R41170 VDD.n7998 VDD.n7997 0.0295514
R41171 VDD.n6579 VDD.n5274 0.0295026
R41172 VDD.n5966 VDD.n5965 0.0295026
R41173 VDD.n6611 VDD.n6610 0.0295026
R41174 VDD.n2056 VDD.n2055 0.0293162
R41175 VDD.n2057 VDD.n2056 0.0293162
R41176 VDD.n2057 VDD.n2026 0.0293162
R41177 VDD.n2059 VDD.n2026 0.0293162
R41178 VDD.n10771 VDD.n2060 0.0293162
R41179 VDD.n10769 VDD.n2060 0.0293162
R41180 VDD.n10769 VDD.n10768 0.0293162
R41181 VDD.n10768 VDD.n10767 0.0293162
R41182 VDD.n2045 VDD.n2044 0.0293162
R41183 VDD.n2045 VDD.n2037 0.0293162
R41184 VDD.n2047 VDD.n2037 0.0293162
R41185 VDD.n2050 VDD.n2049 0.0293162
R41186 VDD.n2051 VDD.n2050 0.0293162
R41187 VDD.n2051 VDD.n2036 0.0293162
R41188 VDD.n2053 VDD.n2036 0.0293162
R41189 VDD.n10808 VDD.n2005 0.0293162
R41190 VDD.n10806 VDD.n2005 0.0293162
R41191 VDD.n10806 VDD.n10805 0.0293162
R41192 VDD.n10805 VDD.n10804 0.0293162
R41193 VDD.n10802 VDD.n2006 0.0293162
R41194 VDD.n10800 VDD.n2006 0.0293162
R41195 VDD.n10800 VDD.n10799 0.0293162
R41196 VDD.n10799 VDD.n10798 0.0293162
R41197 VDD.n1983 VDD.n1982 0.0293162
R41198 VDD.n1984 VDD.n1983 0.0293162
R41199 VDD.n1984 VDD.n1953 0.0293162
R41200 VDD.n1986 VDD.n1953 0.0293162
R41201 VDD.n10811 VDD.n10810 0.0293162
R41202 VDD.n10812 VDD.n10811 0.0293162
R41203 VDD.n10812 VDD.n10809 0.0293162
R41204 VDD.n10814 VDD.n10809 0.0293162
R41205 VDD.n1963 VDD.n1962 0.0293162
R41206 VDD.n1963 VDD.n1955 0.0293162
R41207 VDD.n1965 VDD.n1955 0.0293162
R41208 VDD.n1968 VDD.n1967 0.0293162
R41209 VDD.n1969 VDD.n1968 0.0293162
R41210 VDD.n1969 VDD.n1954 0.0293162
R41211 VDD.n1971 VDD.n1954 0.0293162
R41212 VDD.n10866 VDD.n1932 0.0293162
R41213 VDD.n10864 VDD.n1932 0.0293162
R41214 VDD.n10864 VDD.n10863 0.0293162
R41215 VDD.n10863 VDD.n10862 0.0293162
R41216 VDD.n10860 VDD.n1933 0.0293162
R41217 VDD.n10858 VDD.n1933 0.0293162
R41218 VDD.n10858 VDD.n10857 0.0293162
R41219 VDD.n10857 VDD.n10856 0.0293162
R41220 VDD.n5509 VDD.n5504 0.0293162
R41221 VDD.n5507 VDD.n5504 0.0293162
R41222 VDD.n5507 VDD.n5506 0.0293162
R41223 VDD.n5506 VDD.n5505 0.0293162
R41224 VDD.n10869 VDD.n10868 0.0293162
R41225 VDD.n10870 VDD.n10869 0.0293162
R41226 VDD.n10870 VDD.n10867 0.0293162
R41227 VDD.n10872 VDD.n10867 0.0293162
R41228 VDD.n5519 VDD.n5518 0.0293162
R41229 VDD.n5519 VDD.n5511 0.0293162
R41230 VDD.n5521 VDD.n5511 0.0293162
R41231 VDD.n5524 VDD.n5523 0.0293162
R41232 VDD.n5525 VDD.n5524 0.0293162
R41233 VDD.n5525 VDD.n5510 0.0293162
R41234 VDD.n5527 VDD.n5510 0.0293162
R41235 VDD.n10921 VDD.n1905 0.0293162
R41236 VDD.n10919 VDD.n1905 0.0293162
R41237 VDD.n10919 VDD.n10918 0.0293162
R41238 VDD.n10918 VDD.n10917 0.0293162
R41239 VDD.n10915 VDD.n1906 0.0293162
R41240 VDD.n10913 VDD.n1906 0.0293162
R41241 VDD.n10913 VDD.n10912 0.0293162
R41242 VDD.n10912 VDD.n10911 0.0293162
R41243 VDD.n1891 VDD.n1890 0.0293162
R41244 VDD.n1892 VDD.n1891 0.0293162
R41245 VDD.n1892 VDD.n1861 0.0293162
R41246 VDD.n1894 VDD.n1861 0.0293162
R41247 VDD.n10924 VDD.n10923 0.0293162
R41248 VDD.n10925 VDD.n10924 0.0293162
R41249 VDD.n10925 VDD.n10922 0.0293162
R41250 VDD.n10927 VDD.n10922 0.0293162
R41251 VDD.n1871 VDD.n1870 0.0293162
R41252 VDD.n1871 VDD.n1863 0.0293162
R41253 VDD.n1873 VDD.n1863 0.0293162
R41254 VDD.n1876 VDD.n1875 0.0293162
R41255 VDD.n1877 VDD.n1876 0.0293162
R41256 VDD.n1877 VDD.n1862 0.0293162
R41257 VDD.n1879 VDD.n1862 0.0293162
R41258 VDD.n10976 VDD.n1840 0.0293162
R41259 VDD.n10974 VDD.n1840 0.0293162
R41260 VDD.n10974 VDD.n10973 0.0293162
R41261 VDD.n10973 VDD.n10972 0.0293162
R41262 VDD.n10970 VDD.n1841 0.0293162
R41263 VDD.n10968 VDD.n1841 0.0293162
R41264 VDD.n10968 VDD.n10967 0.0293162
R41265 VDD.n10967 VDD.n10966 0.0293162
R41266 VDD.n1826 VDD.n1825 0.0293162
R41267 VDD.n1827 VDD.n1826 0.0293162
R41268 VDD.n1827 VDD.n1796 0.0293162
R41269 VDD.n1829 VDD.n1796 0.0293162
R41270 VDD.n10979 VDD.n10978 0.0293162
R41271 VDD.n10980 VDD.n10979 0.0293162
R41272 VDD.n10980 VDD.n10977 0.0293162
R41273 VDD.n10982 VDD.n10977 0.0293162
R41274 VDD.n1815 VDD.n1814 0.0293162
R41275 VDD.n1815 VDD.n1807 0.0293162
R41276 VDD.n1817 VDD.n1807 0.0293162
R41277 VDD.n1820 VDD.n1819 0.0293162
R41278 VDD.n1821 VDD.n1820 0.0293162
R41279 VDD.n1821 VDD.n1806 0.0293162
R41280 VDD.n1823 VDD.n1806 0.0293162
R41281 VDD.n1775 VDD.n1774 0.0293162
R41282 VDD.n1776 VDD.n1775 0.0293162
R41283 VDD.n1776 VDD.n1773 0.0293162
R41284 VDD.n1778 VDD.n1773 0.0293162
R41285 VDD.n11025 VDD.n1779 0.0293162
R41286 VDD.n11023 VDD.n1779 0.0293162
R41287 VDD.n11023 VDD.n11022 0.0293162
R41288 VDD.n11022 VDD.n11021 0.0293162
R41289 VDD.n9071 VDD.n9070 0.0293162
R41290 VDD.n9071 VDD.n8474 0.0293162
R41291 VDD.n9073 VDD.n8474 0.0293162
R41292 VDD.n9155 VDD.n9074 0.0293162
R41293 VDD.n9153 VDD.n9074 0.0293162
R41294 VDD.n9153 VDD.n9152 0.0293162
R41295 VDD.n9152 VDD.n9151 0.0293162
R41296 VDD.n9023 VDD.n9022 0.0293162
R41297 VDD.n9024 VDD.n9023 0.0293162
R41298 VDD.n9024 VDD.n8494 0.0293162
R41299 VDD.n9026 VDD.n8494 0.0293162
R41300 VDD.n9031 VDD.n9027 0.0293162
R41301 VDD.n9029 VDD.n9027 0.0293162
R41302 VDD.n9029 VDD.n9028 0.0293162
R41303 VDD.n9028 VDD.n8476 0.0293162
R41304 VDD.n8906 VDD.n8902 0.0293162
R41305 VDD.n8904 VDD.n8902 0.0293162
R41306 VDD.n8904 VDD.n8903 0.0293162
R41307 VDD.n8903 VDD.n8499 0.0293162
R41308 VDD.n9017 VDD.n9016 0.0293162
R41309 VDD.n9018 VDD.n9017 0.0293162
R41310 VDD.n9018 VDD.n8498 0.0293162
R41311 VDD.n9020 VDD.n8498 0.0293162
R41312 VDD.n8898 VDD.n8897 0.0293162
R41313 VDD.n8898 VDD.n8512 0.0293162
R41314 VDD.n8900 VDD.n8512 0.0293162
R41315 VDD.n8934 VDD.n8901 0.0293162
R41316 VDD.n8932 VDD.n8901 0.0293162
R41317 VDD.n8932 VDD.n8931 0.0293162
R41318 VDD.n8931 VDD.n8930 0.0293162
R41319 VDD.n8775 VDD.n8771 0.0293162
R41320 VDD.n8773 VDD.n8771 0.0293162
R41321 VDD.n8773 VDD.n8772 0.0293162
R41322 VDD.n8772 VDD.n8518 0.0293162
R41323 VDD.n8886 VDD.n8885 0.0293162
R41324 VDD.n8887 VDD.n8886 0.0293162
R41325 VDD.n8887 VDD.n8517 0.0293162
R41326 VDD.n8889 VDD.n8517 0.0293162
R41327 VDD.n8766 VDD.n8765 0.0293162
R41328 VDD.n8767 VDD.n8766 0.0293162
R41329 VDD.n8767 VDD.n8531 0.0293162
R41330 VDD.n8769 VDD.n8531 0.0293162
R41331 VDD.n8803 VDD.n8770 0.0293162
R41332 VDD.n8801 VDD.n8770 0.0293162
R41333 VDD.n8801 VDD.n8800 0.0293162
R41334 VDD.n8800 VDD.n8799 0.0293162
R41335 VDD.n8755 VDD.n8754 0.0293162
R41336 VDD.n8755 VDD.n8581 0.0293162
R41337 VDD.n8757 VDD.n8581 0.0293162
R41338 VDD.n8760 VDD.n8759 0.0293162
R41339 VDD.n8761 VDD.n8760 0.0293162
R41340 VDD.n8761 VDD.n8580 0.0293162
R41341 VDD.n8763 VDD.n8580 0.0293162
R41342 VDD.n9149 VDD.n9084 0.0293162
R41343 VDD.n9147 VDD.n9084 0.0293162
R41344 VDD.n9147 VDD.n9146 0.0293162
R41345 VDD.n9146 VDD.n9145 0.0293162
R41346 VDD.n9143 VDD.n9085 0.0293162
R41347 VDD.n9141 VDD.n9085 0.0293162
R41348 VDD.n9141 VDD.n9140 0.0293162
R41349 VDD.n9140 VDD.n9139 0.0293162
R41350 VDD.n8737 VDD.n8736 0.0293162
R41351 VDD.n8738 VDD.n8737 0.0293162
R41352 VDD.n8738 VDD.n8593 0.0293162
R41353 VDD.n8740 VDD.n8593 0.0293162
R41354 VDD.n8743 VDD.n8742 0.0293162
R41355 VDD.n8744 VDD.n8743 0.0293162
R41356 VDD.n8744 VDD.n8592 0.0293162
R41357 VDD.n8746 VDD.n8592 0.0293162
R41358 VDD.n8716 VDD.n8715 0.0293162
R41359 VDD.n8717 VDD.n8716 0.0293162
R41360 VDD.n8717 VDD.n8595 0.0293162
R41361 VDD.n8719 VDD.n8595 0.0293162
R41362 VDD.n8722 VDD.n8721 0.0293162
R41363 VDD.n8723 VDD.n8722 0.0293162
R41364 VDD.n8723 VDD.n8594 0.0293162
R41365 VDD.n8725 VDD.n8594 0.0293162
R41366 VDD.n8705 VDD.n8704 0.0293162
R41367 VDD.n8705 VDD.n8606 0.0293162
R41368 VDD.n8707 VDD.n8606 0.0293162
R41369 VDD.n8710 VDD.n8709 0.0293162
R41370 VDD.n8711 VDD.n8710 0.0293162
R41371 VDD.n8711 VDD.n8605 0.0293162
R41372 VDD.n8713 VDD.n8605 0.0293162
R41373 VDD.n8678 VDD.n8677 0.0293162
R41374 VDD.n8679 VDD.n8678 0.0293162
R41375 VDD.n8679 VDD.n8609 0.0293162
R41376 VDD.n8681 VDD.n8609 0.0293162
R41377 VDD.n8684 VDD.n8683 0.0293162
R41378 VDD.n8685 VDD.n8684 0.0293162
R41379 VDD.n8685 VDD.n8608 0.0293162
R41380 VDD.n8687 VDD.n8608 0.0293162
R41381 VDD.n8666 VDD.n8665 0.0293162
R41382 VDD.n8667 VDD.n8666 0.0293162
R41383 VDD.n8667 VDD.n8620 0.0293162
R41384 VDD.n8669 VDD.n8620 0.0293162
R41385 VDD.n8672 VDD.n8671 0.0293162
R41386 VDD.n8673 VDD.n8672 0.0293162
R41387 VDD.n8673 VDD.n8619 0.0293162
R41388 VDD.n8675 VDD.n8619 0.0293162
R41389 VDD.n8646 VDD.n8645 0.0293162
R41390 VDD.n8646 VDD.n8622 0.0293162
R41391 VDD.n8648 VDD.n8622 0.0293162
R41392 VDD.n8651 VDD.n8650 0.0293162
R41393 VDD.n8652 VDD.n8651 0.0293162
R41394 VDD.n8652 VDD.n8621 0.0293162
R41395 VDD.n8654 VDD.n8621 0.0293162
R41396 VDD.n12620 VDD.n11 0.0293162
R41397 VDD.n12618 VDD.n11 0.0293162
R41398 VDD.n12618 VDD.n12617 0.0293162
R41399 VDD.n12617 VDD.n12616 0.0293162
R41400 VDD.n8634 VDD.n12 0.0293162
R41401 VDD.n8635 VDD.n8634 0.0293162
R41402 VDD.n8635 VDD.n8633 0.0293162
R41403 VDD.n8637 VDD.n8633 0.0293162
R41404 VDD.n7683 VDD.n7682 0.029
R41405 VDD.n2139 VDD.n2138 0.0289485
R41406 VDD.n1177 VDD.n1176 0.0287717
R41407 VDD.n1206 VDD.n1188 0.0287717
R41408 VDD.n1164 VDD.n1163 0.0287717
R41409 VDD.n1176 VDD.n1175 0.0287717
R41410 VDD.n1336 VDD.n1318 0.0287717
R41411 VDD.n1305 VDD.n1304 0.0287717
R41412 VDD.n1337 VDD.n1336 0.0287717
R41413 VDD.n1383 VDD.n1364 0.0287717
R41414 VDD.n1304 VDD.n1286 0.0287717
R41415 VDD.n1073 VDD.n1072 0.0287717
R41416 VDD.n1384 VDD.n1383 0.0287717
R41417 VDD.n1269 VDD.n1250 0.0287717
R41418 VDD.n1237 VDD.n1236 0.0287717
R41419 VDD.n1270 VDD.n1269 0.0287717
R41420 VDD.n1207 VDD.n1206 0.0287717
R41421 VDD.n1236 VDD.n1218 0.0287717
R41422 VDD.n1060 VDD.n1059 0.0287717
R41423 VDD.n1072 VDD.n1071 0.0287717
R41424 VDD.n905 VDD.n0 0.0287717
R41425 VDD.n1059 VDD.n916 0.0287717
R41426 VDD.n1751 VDD.n1750 0.0287717
R41427 VDD.n1163 VDD.n1162 0.0287717
R41428 VDD.n8132 VDD.n8131 0.0284144
R41429 VDD.n8165 VDD.n8164 0.0284144
R41430 VDD.n8111 VDD.n8110 0.0284144
R41431 VDD.n8131 VDD.n8121 0.0284144
R41432 VDD.n8099 VDD.n8098 0.0284144
R41433 VDD.n8110 VDD.n8109 0.0284144
R41434 VDD.n5594 VDD.n5584 0.0284144
R41435 VDD.n8098 VDD.n2104 0.0284144
R41436 VDD.n5615 VDD.n5605 0.0284144
R41437 VDD.n5595 VDD.n5594 0.0284144
R41438 VDD.n5636 VDD.n5626 0.0284144
R41439 VDD.n5616 VDD.n5615 0.0284144
R41440 VDD.n5900 VDD.n5666 0.0284144
R41441 VDD.n5637 VDD.n5636 0.0284144
R41442 VDD.n5866 VDD.n5865 0.0284144
R41443 VDD.n5900 VDD.n5876 0.0284144
R41444 VDD.n5854 VDD.n5853 0.0284144
R41445 VDD.n5865 VDD.n5864 0.0284144
R41446 VDD.n5811 VDD.n5810 0.0284144
R41447 VDD.n5853 VDD.n5843 0.0284144
R41448 VDD.n5799 VDD.n5798 0.0284144
R41449 VDD.n5810 VDD.n5809 0.0284144
R41450 VDD.n5778 VDD.n5777 0.0284144
R41451 VDD.n5798 VDD.n5788 0.0284144
R41452 VDD.n5744 VDD.n5743 0.0284144
R41453 VDD.n5777 VDD.n5776 0.0284144
R41454 VDD.n5723 VDD.n5722 0.0284144
R41455 VDD.n5743 VDD.n5733 0.0284144
R41456 VDD.n11037 VDD.n11036 0.0284144
R41457 VDD.n5722 VDD.n5721 0.0284144
R41458 VDD.n8998 VDD.n8975 0.0284144
R41459 VDD.n9043 VDD.n9042 0.0284144
R41460 VDD.n8947 VDD.n8946 0.0284144
R41461 VDD.n8999 VDD.n8998 0.0284144
R41462 VDD.n8871 VDD.n8848 0.0284144
R41463 VDD.n8946 VDD.n8945 0.0284144
R41464 VDD.n8838 VDD.n8837 0.0284144
R41465 VDD.n8872 VDD.n8871 0.0284144
R41466 VDD.n8560 VDD.n8547 0.0284144
R41467 VDD.n8837 VDD.n8836 0.0284144
R41468 VDD.n12449 VDD.n184 0.0284144
R41469 VDD.n8560 VDD.n8559 0.0284144
R41470 VDD.n170 VDD.n169 0.0284144
R41471 VDD.n12449 VDD.n190 0.0284144
R41472 VDD.n9167 VDD.n8470 0.0284144
R41473 VDD.n9043 VDD.n8488 0.0284144
R41474 VDD.n9167 VDD.n9166 0.0284144
R41475 VDD.n12487 VDD.n106 0.0284144
R41476 VDD.n169 VDD.n168 0.0284144
R41477 VDD.n12505 VDD.n12498 0.0284144
R41478 VDD.n12488 VDD.n12487 0.0284144
R41479 VDD.n90 VDD.n89 0.0284144
R41480 VDD.n12505 VDD.n12504 0.0284144
R41481 VDD.n12543 VDD.n26 0.0284144
R41482 VDD.n89 VDD.n79 0.0284144
R41483 VDD.n12599 VDD.n12554 0.0284144
R41484 VDD.n12544 VDD.n12543 0.0284144
R41485 VDD.n12587 VDD.n12586 0.0284144
R41486 VDD.n12599 VDD.n12598 0.0284144
R41487 VDD.n6713 VDD.n5220 0.0282968
R41488 VDD.n1177 VDD.n1117 0.0282826
R41489 VDD.n1178 VDD.n1117 0.0282826
R41490 VDD.n1179 VDD.n1116 0.0282826
R41491 VDD.n1181 VDD.n1116 0.0282826
R41492 VDD.n1182 VDD.n1181 0.0282826
R41493 VDD.n1184 VDD.n1115 0.0282826
R41494 VDD.n1186 VDD.n1115 0.0282826
R41495 VDD.n1187 VDD.n1114 0.0282826
R41496 VDD.n1188 VDD.n1114 0.0282826
R41497 VDD.n1164 VDD.n1138 0.0282826
R41498 VDD.n1165 VDD.n1138 0.0282826
R41499 VDD.n1166 VDD.n1137 0.0282826
R41500 VDD.n1168 VDD.n1137 0.0282826
R41501 VDD.n1169 VDD.n1168 0.0282826
R41502 VDD.n1171 VDD.n1136 0.0282826
R41503 VDD.n1173 VDD.n1136 0.0282826
R41504 VDD.n1174 VDD.n1135 0.0282826
R41505 VDD.n1175 VDD.n1135 0.0282826
R41506 VDD.n1318 VDD.n1312 0.0282826
R41507 VDD.n1317 VDD.n1312 0.0282826
R41508 VDD.n1316 VDD.n1313 0.0282826
R41509 VDD.n1314 VDD.n1313 0.0282826
R41510 VDD.n1314 VDD.n757 0.0282826
R41511 VDD.n1655 VDD.n756 0.0282826
R41512 VDD.n1657 VDD.n756 0.0282826
R41513 VDD.n1658 VDD.n755 0.0282826
R41514 VDD.n1659 VDD.n755 0.0282826
R41515 VDD.n1660 VDD.n754 0.0282826
R41516 VDD.n1305 VDD.n1280 0.0282826
R41517 VDD.n1306 VDD.n1280 0.0282826
R41518 VDD.n1308 VDD.n1307 0.0282826
R41519 VDD.n1309 VDD.n1308 0.0282826
R41520 VDD.n1309 VDD.n1278 0.0282826
R41521 VDD.n1341 VDD.n1279 0.0282826
R41522 VDD.n1339 VDD.n1279 0.0282826
R41523 VDD.n1338 VDD.n1311 0.0282826
R41524 VDD.n1337 VDD.n1311 0.0282826
R41525 VDD.n1364 VDD.n1080 0.0282826
R41526 VDD.n1363 VDD.n1080 0.0282826
R41527 VDD.n1362 VDD.n1081 0.0282826
R41528 VDD.n1360 VDD.n1081 0.0282826
R41529 VDD.n1360 VDD.n1359 0.0282826
R41530 VDD.n1282 VDD.n1082 0.0282826
R41531 VDD.n1284 VDD.n1282 0.0282826
R41532 VDD.n1285 VDD.n1281 0.0282826
R41533 VDD.n1286 VDD.n1281 0.0282826
R41534 VDD.n1073 VDD.n878 0.0282826
R41535 VDD.n1074 VDD.n878 0.0282826
R41536 VDD.n1076 VDD.n1075 0.0282826
R41537 VDD.n1077 VDD.n1076 0.0282826
R41538 VDD.n1077 VDD.n876 0.0282826
R41539 VDD.n1388 VDD.n877 0.0282826
R41540 VDD.n1386 VDD.n877 0.0282826
R41541 VDD.n1385 VDD.n1079 0.0282826
R41542 VDD.n1384 VDD.n1079 0.0282826
R41543 VDD.n1250 VDD.n1244 0.0282826
R41544 VDD.n1249 VDD.n1244 0.0282826
R41545 VDD.n1248 VDD.n1245 0.0282826
R41546 VDD.n1246 VDD.n1245 0.0282826
R41547 VDD.n1246 VDD.n765 0.0282826
R41548 VDD.n1649 VDD.n766 0.0282826
R41549 VDD.n1647 VDD.n766 0.0282826
R41550 VDD.n1646 VDD.n767 0.0282826
R41551 VDD.n1645 VDD.n767 0.0282826
R41552 VDD.n1644 VDD.n768 0.0282826
R41553 VDD.n1237 VDD.n1109 0.0282826
R41554 VDD.n1238 VDD.n1109 0.0282826
R41555 VDD.n1240 VDD.n1239 0.0282826
R41556 VDD.n1241 VDD.n1240 0.0282826
R41557 VDD.n1241 VDD.n1107 0.0282826
R41558 VDD.n1274 VDD.n1108 0.0282826
R41559 VDD.n1272 VDD.n1108 0.0282826
R41560 VDD.n1271 VDD.n1243 0.0282826
R41561 VDD.n1270 VDD.n1243 0.0282826
R41562 VDD.n1207 VDD.n1113 0.0282826
R41563 VDD.n1208 VDD.n1113 0.0282826
R41564 VDD.n1209 VDD.n1112 0.0282826
R41565 VDD.n1211 VDD.n1112 0.0282826
R41566 VDD.n1212 VDD.n1211 0.0282826
R41567 VDD.n1214 VDD.n1111 0.0282826
R41568 VDD.n1216 VDD.n1111 0.0282826
R41569 VDD.n1217 VDD.n1110 0.0282826
R41570 VDD.n1218 VDD.n1110 0.0282826
R41571 VDD.n1060 VDD.n900 0.0282826
R41572 VDD.n1061 VDD.n900 0.0282826
R41573 VDD.n1062 VDD.n899 0.0282826
R41574 VDD.n1064 VDD.n899 0.0282826
R41575 VDD.n1065 VDD.n1064 0.0282826
R41576 VDD.n1067 VDD.n898 0.0282826
R41577 VDD.n1069 VDD.n898 0.0282826
R41578 VDD.n1070 VDD.n897 0.0282826
R41579 VDD.n1071 VDD.n897 0.0282826
R41580 VDD.n905 VDD.n904 0.0282826
R41581 VDD.n906 VDD.n904 0.0282826
R41582 VDD.n907 VDD.n903 0.0282826
R41583 VDD.n909 VDD.n903 0.0282826
R41584 VDD.n910 VDD.n909 0.0282826
R41585 VDD.n912 VDD.n902 0.0282826
R41586 VDD.n914 VDD.n902 0.0282826
R41587 VDD.n915 VDD.n901 0.0282826
R41588 VDD.n916 VDD.n901 0.0282826
R41589 VDD.n1750 VDD.n683 0.0282826
R41590 VDD.n1749 VDD.n683 0.0282826
R41591 VDD.n1748 VDD.n684 0.0282826
R41592 VDD.n1746 VDD.n684 0.0282826
R41593 VDD.n1746 VDD.n1745 0.0282826
R41594 VDD.n1158 VDD.n685 0.0282826
R41595 VDD.n1160 VDD.n1158 0.0282826
R41596 VDD.n1161 VDD.n1157 0.0282826
R41597 VDD.n1162 VDD.n1157 0.0282826
R41598 VDD.n11873 VDD.n11872 0.027875
R41599 VDD.n8086 VDD.n2120 0.027874
R41600 VDD.n72 VDD.n56 0.0271036
R41601 VDD.n161 VDD.n145 0.0271036
R41602 VDD.n5771 VDD.n5755 0.0271036
R41603 VDD.n5838 VDD.n5822 0.0271036
R41604 VDD.n5655 VDD.n5639 0.0271036
R41605 VDD.n5573 VDD.n5557 0.0271036
R41606 VDD.n8159 VDD.n8143 0.0271036
R41607 VDD.n9116 VDD.n9100 0.0271036
R41608 VDD.n8829 VDD.n8813 0.0271036
R41609 VDD.n9000 VDD.n8969 0.0271036
R41610 VDD.n12572 VDD.n12570 0.0270708
R41611 VDD.n1179 VDD.n1178 0.026913
R41612 VDD.n1184 VDD.n1183 0.026913
R41613 VDD.n1187 VDD.n1186 0.026913
R41614 VDD.n1166 VDD.n1165 0.026913
R41615 VDD.n1171 VDD.n1170 0.026913
R41616 VDD.n1174 VDD.n1173 0.026913
R41617 VDD.n1317 VDD.n1316 0.026913
R41618 VDD.n1655 VDD.n1654 0.026913
R41619 VDD.n1658 VDD.n1657 0.026913
R41620 VDD.n1307 VDD.n1306 0.026913
R41621 VDD.n1342 VDD.n1341 0.026913
R41622 VDD.n1339 VDD.n1338 0.026913
R41623 VDD.n1363 VDD.n1362 0.026913
R41624 VDD.n1358 VDD.n1082 0.026913
R41625 VDD.n1285 VDD.n1284 0.026913
R41626 VDD.n1075 VDD.n1074 0.026913
R41627 VDD.n1389 VDD.n1388 0.026913
R41628 VDD.n1386 VDD.n1385 0.026913
R41629 VDD.n1249 VDD.n1248 0.026913
R41630 VDD.n1650 VDD.n1649 0.026913
R41631 VDD.n1647 VDD.n1646 0.026913
R41632 VDD.n1239 VDD.n1238 0.026913
R41633 VDD.n1275 VDD.n1274 0.026913
R41634 VDD.n1272 VDD.n1271 0.026913
R41635 VDD.n1209 VDD.n1208 0.026913
R41636 VDD.n1214 VDD.n1213 0.026913
R41637 VDD.n1217 VDD.n1216 0.026913
R41638 VDD.n1062 VDD.n1061 0.026913
R41639 VDD.n1067 VDD.n1066 0.026913
R41640 VDD.n1070 VDD.n1069 0.026913
R41641 VDD.n907 VDD.n906 0.026913
R41642 VDD.n912 VDD.n911 0.026913
R41643 VDD.n915 VDD.n914 0.026913
R41644 VDD.n1749 VDD.n1748 0.026913
R41645 VDD.n1744 VDD.n685 0.026913
R41646 VDD.n1161 VDD.n1160 0.026913
R41647 VDD.n1531 VDD.n1530 0.0266202
R41648 VDD.n1544 VDD.n1543 0.0266202
R41649 VDD.n8079 VDD.n2122 0.0261926
R41650 VDD.n9436 VDD.n195 0.026
R41651 VDD.n8075 VDD.n2125 0.0259774
R41652 VDD.n5201 VDD.n5200 0.025625
R41653 VDD.n6302 VDD.n6301 0.0249708
R41654 VDD.n6304 VDD.n6303 0.0249708
R41655 VDD.n6308 VDD.n6307 0.0249708
R41656 VDD.n6306 VDD.n6305 0.0249708
R41657 VDD.n5985 VDD.n5984 0.0249708
R41658 VDD.n5987 VDD.n5986 0.0249708
R41659 VDD.n6315 VDD.n6314 0.0249708
R41660 VDD.n6317 VDD.n6316 0.0249708
R41661 VDD.n6192 VDD.n6191 0.0249708
R41662 VDD.n6194 VDD.n6193 0.0249708
R41663 VDD.n6197 VDD.n6196 0.0249708
R41664 VDD.n6199 VDD.n6198 0.0249708
R41665 VDD.n6182 VDD.n6181 0.0249708
R41666 VDD.n6184 VDD.n6183 0.0249708
R41667 VDD.n6187 VDD.n6186 0.0249708
R41668 VDD.n6189 VDD.n6188 0.0249708
R41669 VDD.n8080 VDD.n2119 0.0242213
R41670 VDD.n8164 VDD.n2089 0.0240829
R41671 VDD.n5556 VDD.n2104 0.0240829
R41672 VDD.n5638 VDD.n5637 0.0240829
R41673 VDD.n5843 VDD.n5680 0.0240829
R41674 VDD.n5776 VDD.n5704 0.0240829
R41675 VDD.n9001 VDD.n8999 0.0240829
R41676 VDD.n8836 VDD.n8525 0.0240829
R41677 VDD.n9123 VDD.n9090 0.0240829
R41678 VDD.n168 VDD.n135 0.0240829
R41679 VDD.n79 VDD.n46 0.0240829
R41680 VDD.n2055 VDD.n2054 0.02404
R41681 VDD.n10767 VDD.n10766 0.02404
R41682 VDD.n2054 VDD.n2053 0.02404
R41683 VDD.n10815 VDD.n10808 0.02404
R41684 VDD.n10798 VDD.n10797 0.02404
R41685 VDD.n1982 VDD.n1981 0.02404
R41686 VDD.n10815 VDD.n10814 0.02404
R41687 VDD.n1981 VDD.n1971 0.02404
R41688 VDD.n10873 VDD.n10866 0.02404
R41689 VDD.n10856 VDD.n10855 0.02404
R41690 VDD.n5528 VDD.n5509 0.02404
R41691 VDD.n10873 VDD.n10872 0.02404
R41692 VDD.n5528 VDD.n5527 0.02404
R41693 VDD.n10928 VDD.n10921 0.02404
R41694 VDD.n10911 VDD.n10910 0.02404
R41695 VDD.n1890 VDD.n1889 0.02404
R41696 VDD.n10928 VDD.n10927 0.02404
R41697 VDD.n1889 VDD.n1879 0.02404
R41698 VDD.n10983 VDD.n10976 0.02404
R41699 VDD.n10966 VDD.n10965 0.02404
R41700 VDD.n1825 VDD.n1824 0.02404
R41701 VDD.n10983 VDD.n10982 0.02404
R41702 VDD.n1824 VDD.n1823 0.02404
R41703 VDD.n1774 VDD.n644 0.02404
R41704 VDD.n11021 VDD.n11020 0.02404
R41705 VDD.n9151 VDD.n9150 0.02404
R41706 VDD.n9022 VDD.n9021 0.02404
R41707 VDD.n9063 VDD.n8476 0.02404
R41708 VDD.n8929 VDD.n8906 0.02404
R41709 VDD.n9021 VDD.n9020 0.02404
R41710 VDD.n8930 VDD.n8929 0.02404
R41711 VDD.n8798 VDD.n8775 0.02404
R41712 VDD.n8890 VDD.n8889 0.02404
R41713 VDD.n8765 VDD.n8764 0.02404
R41714 VDD.n8799 VDD.n8798 0.02404
R41715 VDD.n8764 VDD.n8763 0.02404
R41716 VDD.n9150 VDD.n9149 0.02404
R41717 VDD.n8736 VDD.n8735 0.02404
R41718 VDD.n8747 VDD.n8746 0.02404
R41719 VDD.n8715 VDD.n8714 0.02404
R41720 VDD.n8735 VDD.n8725 0.02404
R41721 VDD.n8714 VDD.n8713 0.02404
R41722 VDD.n8677 VDD.n8676 0.02404
R41723 VDD.n8697 VDD.n8687 0.02404
R41724 VDD.n8665 VDD.n8664 0.02404
R41725 VDD.n8676 VDD.n8675 0.02404
R41726 VDD.n8664 VDD.n8654 0.02404
R41727 VDD.n12621 VDD.n12620 0.02404
R41728 VDD.n8638 VDD.n8637 0.02404
R41729 VDD.n2142 VDD.n2141 0.0234742
R41730 VDD.n2140 VDD.n2139 0.0234742
R41731 VDD.n6713 VDD.n6712 0.0232316
R41732 VDD.n2044 VDD.n2043 0.0232283
R41733 VDD.n1962 VDD.n1961 0.0232283
R41734 VDD.n5518 VDD.n5517 0.0232283
R41735 VDD.n1870 VDD.n1869 0.0232283
R41736 VDD.n1814 VDD.n1813 0.0232283
R41737 VDD.n9070 VDD.n9069 0.0232283
R41738 VDD.n8897 VDD.n8896 0.0232283
R41739 VDD.n8754 VDD.n8753 0.0232283
R41740 VDD.n8704 VDD.n8703 0.0232283
R41741 VDD.n8645 VDD.n8644 0.0232283
R41742 VDD.n6379 VDD.n5374 0.0228966
R41743 VDD.n6362 VDD.n6361 0.0228966
R41744 VDD.n7142 VDD.n2311 0.0228966
R41745 VDD.n7125 VDD.n7124 0.0228966
R41746 VDD.n6379 VDD.n6378 0.0228448
R41747 VDD.n6361 VDD.n5473 0.0228448
R41748 VDD.n7142 VDD.n7141 0.0228448
R41749 VDD.n7124 VDD.n2323 0.0228448
R41750 VDD.n1204 VDD.n1203 0.0225862
R41751 VDD.n1133 VDD.n1132 0.0225862
R41752 VDD.n1334 VDD.n1333 0.0225862
R41753 VDD.n1381 VDD.n1380 0.0225862
R41754 VDD.n1267 VDD.n1266 0.0225862
R41755 VDD.n1234 VDD.n1233 0.0225862
R41756 VDD.n1302 VDD.n1301 0.0225862
R41757 VDD.n895 VDD.n894 0.0225862
R41758 VDD.n1057 VDD.n1056 0.0225862
R41759 VDD.n1155 VDD.n1154 0.0225862
R41760 VDD.n2132 VDD.n2131 0.0224615
R41761 VDD.n12570 VDD.n12569 0.0222742
R41762 VDD.n1642 VDD.n769 0.0221383
R41763 VDD.n6706 VDD.n6705 0.0217183
R41764 VDD.n6692 VDD.n6691 0.0217183
R41765 VDD.n6635 VDD.n5267 0.0217183
R41766 VDD.n6631 VDD.n6630 0.0217183
R41767 VDD.n2120 VDD.n2119 0.021485
R41768 VDD.n4591 VDD.n4590 0.0214211
R41769 VDD.n4590 VDD.n2409 0.0214211
R41770 VDD.n2425 VDD.n2424 0.0207876
R41771 VDD.n5217 VDD.n4593 0.0207876
R41772 VDD.n5204 VDD.n5203 0.0207876
R41773 VDD.n4592 VDD.n2424 0.0207876
R41774 VDD.n5205 VDD.n4594 0.0207876
R41775 VDD.n4599 VDD.n4597 0.0207876
R41776 VDD.n12444 VDD.n194 0.0207876
R41777 VDD.n9200 VDD.n9199 0.0207876
R41778 VDD.n9187 VDD.n8458 0.0207876
R41779 VDD.n12447 VDD.n12446 0.0207876
R41780 VDD.n5366 VDD.n5365 0.0206724
R41781 VDD.n5371 VDD.n5370 0.0206724
R41782 VDD.n6375 VDD.n6374 0.0206724
R41783 VDD.n6217 VDD.n6216 0.0206724
R41784 VDD.n6264 VDD.n6263 0.0206724
R41785 VDD.n6366 VDD.n6365 0.0206724
R41786 VDD.n5940 VDD.n5939 0.0206724
R41787 VDD.n5946 VDD.n5945 0.0206724
R41788 VDD.n2359 VDD.n2358 0.0206724
R41789 VDD.n2364 VDD.n2363 0.0206724
R41790 VDD.n7138 VDD.n7137 0.0206724
R41791 VDD.n2315 VDD.n2314 0.0206724
R41792 VDD.n2398 VDD.n2397 0.0206724
R41793 VDD.n7129 VDD.n7128 0.0206724
R41794 VDD.n2346 VDD.n2345 0.0206724
R41795 VDD.n7046 VDD.n7045 0.0206724
R41796 VDD.n1708 VDD.n728 0.0206207
R41797 VDD.n1610 VDD.n802 0.0206207
R41798 VDD.n1442 VDD.n839 0.0206207
R41799 VDD.n1480 VDD.n1476 0.0206207
R41800 VDD.n1708 VDD.n1707 0.0206207
R41801 VDD.n1732 VDD.n699 0.0206207
R41802 VDD.n1732 VDD.n1731 0.0206207
R41803 VDD.n6563 VDD.n6562 0.0204161
R41804 VDD.n6410 VDD.n5297 0.0204161
R41805 VDD.n6873 VDD.n2384 0.0204161
R41806 VDD.n7026 VDD.n7025 0.0204161
R41807 VDD.n1533 VDD.n1532 0.0203361
R41808 VDD.n1546 VDD.n1545 0.0203361
R41809 VDD.n75 VDD.n72 0.0199738
R41810 VDD.n164 VDD.n161 0.0199738
R41811 VDD.n5772 VDD.n5771 0.0199738
R41812 VDD.n5839 VDD.n5838 0.0199738
R41813 VDD.n5656 VDD.n5655 0.0199738
R41814 VDD.n5574 VDD.n5573 0.0199738
R41815 VDD.n8160 VDD.n8159 0.0199738
R41816 VDD.n9119 VDD.n9116 0.0199738
R41817 VDD.n8832 VDD.n8829 0.0199738
R41818 VDD.n9003 VDD.n8969 0.0199738
R41819 VDD.n6037 VDD.n6022 0.019782
R41820 VDD.n6157 VDD.n6018 0.019782
R41821 VDD.n6849 VDD.n2404 0.019782
R41822 VDD.n6727 VDD.n2406 0.019782
R41823 VDD.n6009 VDD.n6007 0.0196477
R41824 VDD.n6331 VDD.n6330 0.0196477
R41825 VDD.n7173 VDD.n7172 0.0196477
R41826 VDD.n7096 VDD.n7095 0.0196477
R41827 VDD.n9138 VDD.n9137 0.0193079
R41828 VDD.n9136 VDD.n9135 0.0193079
R41829 VDD.n9127 VDD.n9126 0.0193079
R41830 VDD.n9125 VDD.n9124 0.0193079
R41831 VDD.n12566 VDD.n12565 0.0193079
R41832 VDD.n12569 VDD.n12567 0.0193079
R41833 VDD.n12573 VDD.n12572 0.0193079
R41834 VDD.n12576 VDD.n12574 0.0193079
R41835 VDD.n8128 VDD.n8127 0.0192265
R41836 VDD.n2032 VDD.n2031 0.0192265
R41837 VDD.n2099 VDD.n2098 0.0192265
R41838 VDD.n10793 VDD.n10792 0.0192265
R41839 VDD.n5591 VDD.n5590 0.0192265
R41840 VDD.n1977 VDD.n1976 0.0192265
R41841 VDD.n5612 VDD.n5611 0.0192265
R41842 VDD.n10851 VDD.n10850 0.0192265
R41843 VDD.n5897 VDD.n5896 0.0192265
R41844 VDD.n5499 VDD.n5498 0.0192265
R41845 VDD.n5675 VDD.n5674 0.0192265
R41846 VDD.n10906 VDD.n10905 0.0192265
R41847 VDD.n5688 VDD.n5687 0.0192265
R41848 VDD.n1885 VDD.n1884 0.0192265
R41849 VDD.n5795 VDD.n5794 0.0192265
R41850 VDD.n10961 VDD.n10960 0.0192265
R41851 VDD.n5740 VDD.n5739 0.0192265
R41852 VDD.n1802 VDD.n1801 0.0192265
R41853 VDD.n5714 VDD.n5713 0.0192265
R41854 VDD.n11016 VDD.n11015 0.0192265
R41855 VDD.n9060 VDD.n9059 0.0192265
R41856 VDD.n9048 VDD.n9046 0.0192265
R41857 VDD.n8926 VDD.n8925 0.0192265
R41858 VDD.n8914 VDD.n8912 0.0192265
R41859 VDD.n8852 VDD.n8849 0.0192265
R41860 VDD.n8867 VDD.n8866 0.0192265
R41861 VDD.n8577 VDD.n8576 0.0192265
R41862 VDD.n8565 VDD.n8563 0.0192265
R41863 VDD.n9081 VDD.n9080 0.0192265
R41864 VDD.n9172 VDD.n9170 0.0192265
R41865 VDD.n8589 VDD.n8588 0.0192265
R41866 VDD.n12454 VDD.n12452 0.0192265
R41867 VDD.n8602 VDD.n8601 0.0192265
R41868 VDD.n12483 VDD.n12482 0.0192265
R41869 VDD.n8694 VDD.n8693 0.0192265
R41870 VDD.n12510 VDD.n12508 0.0192265
R41871 VDD.n8661 VDD.n8660 0.0192265
R41872 VDD.n12539 VDD.n12538 0.0192265
R41873 VDD.n8630 VDD.n8629 0.0192265
R41874 VDD.n12604 VDD.n12602 0.0192265
R41875 VDD.n8086 VDD.n8085 0.019179
R41876 VDD.n2116 VDD.n2115 0.0190522
R41877 VDD.n10823 VDD.n10821 0.0190522
R41878 VDD.n5633 VDD.n5632 0.0190522
R41879 VDD.n10878 VDD.n10876 0.0190522
R41880 VDD.n5850 VDD.n5849 0.0190522
R41881 VDD.n10933 VDD.n10931 0.0190522
R41882 VDD.n5701 VDD.n5700 0.0190522
R41883 VDD.n10988 VDD.n10986 0.0190522
R41884 VDD.n8979 VDD.n8976 0.0190522
R41885 VDD.n8994 VDD.n8993 0.0190522
R41886 VDD.n8795 VDD.n8794 0.0190522
R41887 VDD.n8783 VDD.n8781 0.0190522
R41888 VDD.n8732 VDD.n8731 0.0190522
R41889 VDD.n131 VDD.n130 0.0190522
R41890 VDD.n8616 VDD.n8615 0.0190522
R41891 VDD.n85 VDD.n84 0.0190522
R41892 VDD.n6707 VDD.n6706 0.0189386
R41893 VDD.n6693 VDD.n6692 0.0189386
R41894 VDD.n6636 VDD.n6635 0.0189386
R41895 VDD.n6631 VDD.n5269 0.0189386
R41896 VDD.n12562 VDD.n12559 0.0186448
R41897 VDD.n12578 VDD.n12559 0.0186448
R41898 VDD.n643 VDD.n637 0.0186448
R41899 VDD.n639 VDD.n637 0.0186448
R41900 VDD.n11128 VDD.n636 0.0186448
R41901 VDD.n675 VDD.n672 0.0186448
R41902 VDD.n675 VDD.n671 0.0186448
R41903 VDD.n674 VDD.n670 0.0186448
R41904 VDD.n6322 VDD.n6321 0.0186448
R41905 VDD.n5982 VDD.n5913 0.0186448
R41906 VDD.n6324 VDD.n5915 0.0186448
R41907 VDD.n6321 VDD.n5983 0.0186448
R41908 VDD.n5983 VDD.n5982 0.0186448
R41909 VDD.n5981 VDD.n5915 0.0186448
R41910 VDD.n6176 VDD.n6015 0.0186448
R41911 VDD.n6178 VDD.n6017 0.0186448
R41912 VDD.n6172 VDD.n6012 0.0186448
R41913 VDD.n6176 VDD.n6012 0.0186448
R41914 VDD.n6017 VDD.n6011 0.0186448
R41915 VDD.n5532 VDD.n5531 0.0186448
R41916 VDD.n5531 VDD.n5530 0.0186448
R41917 VDD.n5536 VDD.n5535 0.0186448
R41918 VDD.n5882 VDD.n5881 0.0186448
R41919 VDD.n5887 VDD.n5881 0.0186448
R41920 VDD.n5885 VDD.n5884 0.0186448
R41921 VDD.n5906 VDD.n5904 0.0186448
R41922 VDD.n5903 VDD.n5540 0.0186448
R41923 VDD.n5909 VDD.n5908 0.0186448
R41924 VDD.n10816 VDD.n1997 0.0186448
R41925 VDD.n2003 VDD.n1997 0.0186448
R41926 VDD.n10818 VDD.n1996 0.0186448
R41927 VDD.n8093 VDD.n2110 0.0186448
R41928 VDD.n2110 VDD.n2107 0.0186448
R41929 VDD.n2118 VDD.n2117 0.0186448
R41930 VDD.n10816 VDD.n2001 0.0186448
R41931 VDD.n10819 VDD.n10818 0.0186448
R41932 VDD.n8094 VDD.n8093 0.0186448
R41933 VDD.n8091 VDD.n2107 0.0186448
R41934 VDD.n2117 VDD.n2109 0.0186448
R41935 VDD.n2003 VDD.n2002 0.0186448
R41936 VDD.n5533 VDD.n5532 0.0186448
R41937 VDD.n5883 VDD.n5882 0.0186448
R41938 VDD.n5904 VDD.n5903 0.0186448
R41939 VDD.n5530 VDD.n5489 0.0186448
R41940 VDD.n5910 VDD.n5909 0.0186448
R41941 VDD.n5884 VDD.n5880 0.0186448
R41942 VDD.n5888 VDD.n5887 0.0186448
R41943 VDD.n5537 VDD.n5536 0.0186448
R41944 VDD.n1764 VDD.n671 0.0186448
R41945 VDD.n11045 VDD.n670 0.0186448
R41946 VDD.n11047 VDD.n672 0.0186448
R41947 VDD.n11129 VDD.n11128 0.0186448
R41948 VDD.n639 VDD.n634 0.0186448
R41949 VDD.n643 VDD.n635 0.0186448
R41950 VDD.n12578 VDD.n12561 0.0186448
R41951 VDD.n12580 VDD.n12560 0.0186448
R41952 VDD.n12584 VDD.n12562 0.0186448
R41953 VDD.n12628 VDD.n12627 0.0186448
R41954 VDD.n12622 VDD.n8 0.0186448
R41955 VDD.n12631 VDD.n10 0.0186448
R41956 VDD.n12629 VDD.n10 0.0186448
R41957 VDD.n12627 VDD.n12623 0.0186448
R41958 VDD.n12623 VDD.n12622 0.0186448
R41959 VDD.n12638 VDD.n12637 0.0186448
R41960 VDD.n4 VDD.n3 0.0186448
R41961 VDD.n1001 VDD.n955 0.0186448
R41962 VDD.n999 VDD.n953 0.0186448
R41963 VDD.n1754 VDD.n1753 0.0186448
R41964 VDD.n1758 VDD.n1757 0.0186448
R41965 VDD.n1753 VDD.n677 0.0186448
R41966 VDD.n1759 VDD.n1758 0.0186448
R41967 VDD.n999 VDD.n954 0.0186448
R41968 VDD.n957 VDD.n955 0.0186448
R41969 VDD.n5 VDD.n4 0.0186448
R41970 VDD.n12637 VDD.n12636 0.0186448
R41971 VDD.n10772 VDD.n2059 0.0185609
R41972 VDD.n2048 VDD.n2047 0.0185609
R41973 VDD.n10804 VDD.n10803 0.0185609
R41974 VDD.n1987 VDD.n1986 0.0185609
R41975 VDD.n1966 VDD.n1965 0.0185609
R41976 VDD.n10862 VDD.n10861 0.0185609
R41977 VDD.n5505 VDD.n1922 0.0185609
R41978 VDD.n5522 VDD.n5521 0.0185609
R41979 VDD.n10917 VDD.n10916 0.0185609
R41980 VDD.n1895 VDD.n1894 0.0185609
R41981 VDD.n1874 VDD.n1873 0.0185609
R41982 VDD.n10972 VDD.n10971 0.0185609
R41983 VDD.n1830 VDD.n1829 0.0185609
R41984 VDD.n1818 VDD.n1817 0.0185609
R41985 VDD.n11026 VDD.n1778 0.0185609
R41986 VDD.n9156 VDD.n9073 0.0185609
R41987 VDD.n9032 VDD.n9026 0.0185609
R41988 VDD.n9015 VDD.n8499 0.0185609
R41989 VDD.n8935 VDD.n8900 0.0185609
R41990 VDD.n8884 VDD.n8518 0.0185609
R41991 VDD.n8804 VDD.n8769 0.0185609
R41992 VDD.n8758 VDD.n8757 0.0185609
R41993 VDD.n9145 VDD.n9144 0.0185609
R41994 VDD.n8741 VDD.n8740 0.0185609
R41995 VDD.n8720 VDD.n8719 0.0185609
R41996 VDD.n8708 VDD.n8707 0.0185609
R41997 VDD.n8682 VDD.n8681 0.0185609
R41998 VDD.n8670 VDD.n8669 0.0185609
R41999 VDD.n8649 VDD.n8648 0.0185609
R42000 VDD.n12616 VDD.n12615 0.0185609
R42001 VDD.n8065 VDD.n8064 0.0185
R42002 VDD.n8125 VDD.n8124 0.0183497
R42003 VDD.n2028 VDD.n2027 0.0183497
R42004 VDD.n2096 VDD.n2095 0.0183497
R42005 VDD.n10789 VDD.n10788 0.0183497
R42006 VDD.n5588 VDD.n5587 0.0183497
R42007 VDD.n1973 VDD.n1972 0.0183497
R42008 VDD.n5609 VDD.n5608 0.0183497
R42009 VDD.n10847 VDD.n10846 0.0183497
R42010 VDD.n5894 VDD.n5893 0.0183497
R42011 VDD.n5495 VDD.n5494 0.0183497
R42012 VDD.n5672 VDD.n5671 0.0183497
R42013 VDD.n10902 VDD.n10901 0.0183497
R42014 VDD.n5685 VDD.n5684 0.0183497
R42015 VDD.n1881 VDD.n1880 0.0183497
R42016 VDD.n5792 VDD.n5791 0.0183497
R42017 VDD.n10957 VDD.n10956 0.0183497
R42018 VDD.n5737 VDD.n5736 0.0183497
R42019 VDD.n1798 VDD.n1797 0.0183497
R42020 VDD.n5711 VDD.n5710 0.0183497
R42021 VDD.n11012 VDD.n11011 0.0183497
R42022 VDD.n9057 VDD.n9056 0.0183497
R42023 VDD.n9050 VDD.n9049 0.0183497
R42024 VDD.n8923 VDD.n8922 0.0183497
R42025 VDD.n8916 VDD.n8915 0.0183497
R42026 VDD.n8854 VDD.n8853 0.0183497
R42027 VDD.n8863 VDD.n8862 0.0183497
R42028 VDD.n8574 VDD.n8573 0.0183497
R42029 VDD.n8567 VDD.n8566 0.0183497
R42030 VDD.n9078 VDD.n9077 0.0183497
R42031 VDD.n9174 VDD.n9173 0.0183497
R42032 VDD.n8586 VDD.n8585 0.0183497
R42033 VDD.n12456 VDD.n12455 0.0183497
R42034 VDD.n8599 VDD.n8598 0.0183497
R42035 VDD.n12479 VDD.n12478 0.0183497
R42036 VDD.n8691 VDD.n8690 0.0183497
R42037 VDD.n12512 VDD.n12511 0.0183497
R42038 VDD.n8658 VDD.n8657 0.0183497
R42039 VDD.n12535 VDD.n12534 0.0183497
R42040 VDD.n8627 VDD.n8626 0.0183497
R42041 VDD.n12606 VDD.n12605 0.0183497
R42042 VDD.n2113 VDD.n2112 0.0181836
R42043 VDD.n10825 VDD.n10824 0.0181836
R42044 VDD.n5630 VDD.n5629 0.0181836
R42045 VDD.n10880 VDD.n10879 0.0181836
R42046 VDD.n5847 VDD.n5846 0.0181836
R42047 VDD.n10935 VDD.n10934 0.0181836
R42048 VDD.n5698 VDD.n5697 0.0181836
R42049 VDD.n10990 VDD.n10989 0.0181836
R42050 VDD.n8981 VDD.n8980 0.0181836
R42051 VDD.n8990 VDD.n8989 0.0181836
R42052 VDD.n8792 VDD.n8791 0.0181836
R42053 VDD.n8785 VDD.n8784 0.0181836
R42054 VDD.n8729 VDD.n8728 0.0181836
R42055 VDD.n127 VDD.n126 0.0181836
R42056 VDD.n8613 VDD.n8612 0.0181836
R42057 VDD.n81 VDD.n80 0.0181836
R42058 VDD.n9130 VDD.n9128 0.0181276
R42059 VDD.n9132 VDD.n9128 0.0181276
R42060 VDD.n9133 VDD.n8459 0.0181276
R42061 VDD.n8081 VDD.n8079 0.0179831
R42062 VDD.n8075 VDD.n8074 0.0178367
R42063 VDD.n6037 VDD.n6036 0.0177463
R42064 VDD.n6169 VDD.n6157 0.0177463
R42065 VDD.n6850 VDD.n6849 0.0177463
R42066 VDD.n6727 VDD.n6726 0.0177463
R42067 VDD.n12563 VDD.n9 0.0176669
R42068 VDD.n8138 VDD.n8137 0.0175856
R42069 VDD.n8117 VDD.n8116 0.0175856
R42070 VDD.n8105 VDD.n8104 0.0175856
R42071 VDD.n5579 VDD.n5578 0.0175856
R42072 VDD.n5600 VDD.n5599 0.0175856
R42073 VDD.n5621 VDD.n5620 0.0175856
R42074 VDD.n5661 VDD.n5660 0.0175856
R42075 VDD.n5872 VDD.n5871 0.0175856
R42076 VDD.n5860 VDD.n5859 0.0175856
R42077 VDD.n5817 VDD.n5816 0.0175856
R42078 VDD.n5805 VDD.n5804 0.0175856
R42079 VDD.n5784 VDD.n5783 0.0175856
R42080 VDD.n5750 VDD.n5749 0.0175856
R42081 VDD.n5729 VDD.n5728 0.0175856
R42082 VDD.n11031 VDD.n1770 0.0175856
R42083 VDD.n9038 VDD.n9037 0.0175856
R42084 VDD.n9008 VDD.n9007 0.0175856
R42085 VDD.n8941 VDD.n8940 0.0175856
R42086 VDD.n8877 VDD.n8876 0.0175856
R42087 VDD.n8810 VDD.n8809 0.0175856
R42088 VDD.n8555 VDD.n8554 0.0175856
R42089 VDD.n186 VDD.n175 0.0175856
R42090 VDD.n9097 VDD.n9096 0.0175856
R42091 VDD.n9162 VDD.n9161 0.0175856
R42092 VDD.n142 VDD.n141 0.0175856
R42093 VDD.n12493 VDD.n12492 0.0175856
R42094 VDD.n12500 VDD.n95 0.0175856
R42095 VDD.n53 VDD.n52 0.0175856
R42096 VDD.n12549 VDD.n12548 0.0175856
R42097 VDD.n12594 VDD.n12593 0.0175856
R42098 VDD.n10797 VDD.n2007 0.0175462
R42099 VDD.n10855 VDD.n1934 0.0175462
R42100 VDD.n10910 VDD.n1907 0.0175462
R42101 VDD.n10965 VDD.n1842 0.0175462
R42102 VDD.n11020 VDD.n1780 0.0175462
R42103 VDD.n9064 VDD.n9063 0.0175462
R42104 VDD.n8891 VDD.n8890 0.0175462
R42105 VDD.n8748 VDD.n8747 0.0175462
R42106 VDD.n8698 VDD.n8697 0.0175462
R42107 VDD.n8639 VDD.n8638 0.0175462
R42108 VDD.n6699 VDD.n5262 0.0174226
R42109 VDD.n7124 VDD.n2322 0.0174226
R42110 VDD.n6361 VDD.n5472 0.0174226
R42111 VDD.n5445 VDD.n5444 0.0174226
R42112 VDD.n6379 VDD.n5361 0.0174226
R42113 VDD.n6699 VDD.n5263 0.0174226
R42114 VDD.n6380 VDD.n6379 0.0174226
R42115 VDD.n6361 VDD.n6360 0.0174226
R42116 VDD.n7143 VDD.n7142 0.0174226
R42117 VDD.n5444 VDD.n5433 0.0174226
R42118 VDD.n7142 VDD.n2310 0.0174226
R42119 VDD.n7124 VDD.n7123 0.0174226
R42120 VDD.n12440 VDD.n195 0.017375
R42121 VDD.n1664 VDD.n752 0.0172098
R42122 VDD.n1573 VDD.n1507 0.0172098
R42123 VDD.n1574 VDD.n1507 0.0172098
R42124 VDD.n1665 VDD.n752 0.0172098
R42125 VDD.n5262 VDD.n5222 0.0171298
R42126 VDD.n5260 VDD.n5222 0.0171298
R42127 VDD.n5260 VDD.n5259 0.0171298
R42128 VDD.n5259 VDD.n5258 0.0171298
R42129 VDD.n5258 VDD.n5225 0.0171298
R42130 VDD.n5255 VDD.n5225 0.0171298
R42131 VDD.n5255 VDD.n5254 0.0171298
R42132 VDD.n5254 VDD.n5253 0.0171298
R42133 VDD.n5252 VDD.n5227 0.0171298
R42134 VDD.n5250 VDD.n5227 0.0171298
R42135 VDD.n5248 VDD.n5247 0.0171298
R42136 VDD.n5247 VDD.n5230 0.0171298
R42137 VDD.n5245 VDD.n5230 0.0171298
R42138 VDD.n5244 VDD.n5231 0.0171298
R42139 VDD.n5242 VDD.n5231 0.0171298
R42140 VDD.n5242 VDD.n5241 0.0171298
R42141 VDD.n5241 VDD.n5240 0.0171298
R42142 VDD.n5240 VDD.n5234 0.0171298
R42143 VDD.n5237 VDD.n5234 0.0171298
R42144 VDD.n5237 VDD.n5236 0.0171298
R42145 VDD.n5236 VDD.n2322 0.0171298
R42146 VDD.n5472 VDD.n5379 0.0171298
R42147 VDD.n5470 VDD.n5379 0.0171298
R42148 VDD.n5470 VDD.n5469 0.0171298
R42149 VDD.n5469 VDD.n5468 0.0171298
R42150 VDD.n5468 VDD.n5382 0.0171298
R42151 VDD.n5465 VDD.n5382 0.0171298
R42152 VDD.n5465 VDD.n5464 0.0171298
R42153 VDD.n5464 VDD.n5463 0.0171298
R42154 VDD.n5462 VDD.n5384 0.0171298
R42155 VDD.n5460 VDD.n5384 0.0171298
R42156 VDD.n5458 VDD.n5457 0.0171298
R42157 VDD.n5457 VDD.n5387 0.0171298
R42158 VDD.n5455 VDD.n5387 0.0171298
R42159 VDD.n5454 VDD.n5388 0.0171298
R42160 VDD.n5452 VDD.n5388 0.0171298
R42161 VDD.n5452 VDD.n5451 0.0171298
R42162 VDD.n5451 VDD.n5450 0.0171298
R42163 VDD.n5450 VDD.n5391 0.0171298
R42164 VDD.n5447 VDD.n5391 0.0171298
R42165 VDD.n5447 VDD.n5446 0.0171298
R42166 VDD.n5446 VDD.n5445 0.0171298
R42167 VDD.n5361 VDD.n5321 0.0171298
R42168 VDD.n5359 VDD.n5321 0.0171298
R42169 VDD.n5359 VDD.n5358 0.0171298
R42170 VDD.n5358 VDD.n5357 0.0171298
R42171 VDD.n5357 VDD.n5324 0.0171298
R42172 VDD.n5354 VDD.n5324 0.0171298
R42173 VDD.n5354 VDD.n5353 0.0171298
R42174 VDD.n5353 VDD.n5352 0.0171298
R42175 VDD.n5351 VDD.n5326 0.0171298
R42176 VDD.n5349 VDD.n5326 0.0171298
R42177 VDD.n5347 VDD.n5346 0.0171298
R42178 VDD.n5346 VDD.n5329 0.0171298
R42179 VDD.n5344 VDD.n5329 0.0171298
R42180 VDD.n5343 VDD.n5330 0.0171298
R42181 VDD.n5341 VDD.n5330 0.0171298
R42182 VDD.n5341 VDD.n5340 0.0171298
R42183 VDD.n5340 VDD.n5339 0.0171298
R42184 VDD.n5339 VDD.n5333 0.0171298
R42185 VDD.n5336 VDD.n5333 0.0171298
R42186 VDD.n5336 VDD.n5335 0.0171298
R42187 VDD.n5335 VDD.n5263 0.0171298
R42188 VDD.n6010 VDD.n6009 0.0171298
R42189 VDD.n6007 VDD.n5989 0.0171298
R42190 VDD.n6005 VDD.n5989 0.0171298
R42191 VDD.n6005 VDD.n6004 0.0171298
R42192 VDD.n6004 VDD.n6003 0.0171298
R42193 VDD.n6003 VDD.n5992 0.0171298
R42194 VDD.n6000 VDD.n5992 0.0171298
R42195 VDD.n6000 VDD.n5999 0.0171298
R42196 VDD.n5999 VDD.n5998 0.0171298
R42197 VDD.n5997 VDD.n5995 0.0171298
R42198 VDD.n5995 VDD.n5313 0.0171298
R42199 VDD.n6393 VDD.n6392 0.0171298
R42200 VDD.n6392 VDD.n5315 0.0171298
R42201 VDD.n6390 VDD.n5315 0.0171298
R42202 VDD.n6389 VDD.n5316 0.0171298
R42203 VDD.n6387 VDD.n5316 0.0171298
R42204 VDD.n6387 VDD.n6386 0.0171298
R42205 VDD.n6386 VDD.n6385 0.0171298
R42206 VDD.n6385 VDD.n5319 0.0171298
R42207 VDD.n6382 VDD.n5319 0.0171298
R42208 VDD.n6382 VDD.n6381 0.0171298
R42209 VDD.n6381 VDD.n6380 0.0171298
R42210 VDD.n6330 VDD.n5486 0.0171298
R42211 VDD.n6331 VDD.n5485 0.0171298
R42212 VDD.n6333 VDD.n5485 0.0171298
R42213 VDD.n6333 VDD.n5484 0.0171298
R42214 VDD.n6336 VDD.n5484 0.0171298
R42215 VDD.n6336 VDD.n5483 0.0171298
R42216 VDD.n6339 VDD.n5483 0.0171298
R42217 VDD.n6339 VDD.n5482 0.0171298
R42218 VDD.n6341 VDD.n5482 0.0171298
R42219 VDD.n6342 VDD.n5480 0.0171298
R42220 VDD.n6344 VDD.n5480 0.0171298
R42221 VDD.n6347 VDD.n5479 0.0171298
R42222 VDD.n6347 VDD.n5478 0.0171298
R42223 VDD.n6349 VDD.n5478 0.0171298
R42224 VDD.n6350 VDD.n5477 0.0171298
R42225 VDD.n6352 VDD.n5477 0.0171298
R42226 VDD.n6352 VDD.n5476 0.0171298
R42227 VDD.n6355 VDD.n5476 0.0171298
R42228 VDD.n6355 VDD.n5475 0.0171298
R42229 VDD.n6358 VDD.n5475 0.0171298
R42230 VDD.n6358 VDD.n5474 0.0171298
R42231 VDD.n6360 VDD.n5474 0.0171298
R42232 VDD.n7143 VDD.n2309 0.0171298
R42233 VDD.n7145 VDD.n2309 0.0171298
R42234 VDD.n7145 VDD.n2308 0.0171298
R42235 VDD.n7148 VDD.n2308 0.0171298
R42236 VDD.n7148 VDD.n2307 0.0171298
R42237 VDD.n7151 VDD.n2307 0.0171298
R42238 VDD.n7151 VDD.n2306 0.0171298
R42239 VDD.n7153 VDD.n2306 0.0171298
R42240 VDD.n7154 VDD.n2304 0.0171298
R42241 VDD.n7156 VDD.n2304 0.0171298
R42242 VDD.n7159 VDD.n2303 0.0171298
R42243 VDD.n7159 VDD.n2302 0.0171298
R42244 VDD.n7161 VDD.n2302 0.0171298
R42245 VDD.n7162 VDD.n2301 0.0171298
R42246 VDD.n7164 VDD.n2301 0.0171298
R42247 VDD.n7164 VDD.n2300 0.0171298
R42248 VDD.n7167 VDD.n2300 0.0171298
R42249 VDD.n7167 VDD.n2299 0.0171298
R42250 VDD.n7170 VDD.n2299 0.0171298
R42251 VDD.n7170 VDD.n2298 0.0171298
R42252 VDD.n7172 VDD.n2298 0.0171298
R42253 VDD.n7173 VDD.n2297 0.0171298
R42254 VDD.n5433 VDD.n5393 0.0171298
R42255 VDD.n5431 VDD.n5393 0.0171298
R42256 VDD.n5431 VDD.n5430 0.0171298
R42257 VDD.n5430 VDD.n5429 0.0171298
R42258 VDD.n5429 VDD.n5396 0.0171298
R42259 VDD.n5426 VDD.n5396 0.0171298
R42260 VDD.n5426 VDD.n5425 0.0171298
R42261 VDD.n5425 VDD.n5424 0.0171298
R42262 VDD.n5423 VDD.n5398 0.0171298
R42263 VDD.n5421 VDD.n5398 0.0171298
R42264 VDD.n5419 VDD.n5418 0.0171298
R42265 VDD.n5418 VDD.n5401 0.0171298
R42266 VDD.n5416 VDD.n5401 0.0171298
R42267 VDD.n5415 VDD.n5402 0.0171298
R42268 VDD.n5413 VDD.n5402 0.0171298
R42269 VDD.n5413 VDD.n5412 0.0171298
R42270 VDD.n5412 VDD.n5411 0.0171298
R42271 VDD.n5411 VDD.n5405 0.0171298
R42272 VDD.n5408 VDD.n5405 0.0171298
R42273 VDD.n5408 VDD.n5407 0.0171298
R42274 VDD.n5407 VDD.n2310 0.0171298
R42275 VDD.n7123 VDD.n2324 0.0171298
R42276 VDD.n7121 VDD.n2324 0.0171298
R42277 VDD.n7121 VDD.n7120 0.0171298
R42278 VDD.n7120 VDD.n7119 0.0171298
R42279 VDD.n7119 VDD.n2327 0.0171298
R42280 VDD.n7116 VDD.n2327 0.0171298
R42281 VDD.n7116 VDD.n7115 0.0171298
R42282 VDD.n7115 VDD.n7114 0.0171298
R42283 VDD.n7113 VDD.n2329 0.0171298
R42284 VDD.n7111 VDD.n2329 0.0171298
R42285 VDD.n7109 VDD.n7108 0.0171298
R42286 VDD.n7108 VDD.n7089 0.0171298
R42287 VDD.n7106 VDD.n7089 0.0171298
R42288 VDD.n7105 VDD.n7090 0.0171298
R42289 VDD.n7103 VDD.n7090 0.0171298
R42290 VDD.n7103 VDD.n7102 0.0171298
R42291 VDD.n7102 VDD.n7101 0.0171298
R42292 VDD.n7101 VDD.n7093 0.0171298
R42293 VDD.n7098 VDD.n7093 0.0171298
R42294 VDD.n7098 VDD.n7097 0.0171298
R42295 VDD.n7097 VDD.n7096 0.0171298
R42296 VDD.n7095 VDD.n2240 0.0171298
R42297 VDD.n1530 VDD.n1523 0.0167842
R42298 VDD.n1531 VDD.n1522 0.0167842
R42299 VDD.n1532 VDD.n1522 0.0167842
R42300 VDD.n1547 VDD.n1546 0.0167842
R42301 VDD.n1545 VDD.n1534 0.0167842
R42302 VDD.n1544 VDD.n1534 0.0167842
R42303 VDD.n1543 VDD.n1535 0.0167842
R42304 VDD.n1672 VDD.n1671 0.016681
R42305 VDD.n4590 VDD.n4589 0.016625
R42306 VDD.n1582 VDD.n747 0.0165752
R42307 VDD.n1202 VDD.n1201 0.0164828
R42308 VDD.n1200 VDD.n1199 0.0164828
R42309 VDD.n1198 VDD.n1197 0.0164828
R42310 VDD.n1196 VDD.n1195 0.0164828
R42311 VDD.n1434 VDD.n1433 0.0164828
R42312 VDD.n1436 VDD.n1435 0.0164828
R42313 VDD.n1438 VDD.n1437 0.0164828
R42314 VDD.n1440 VDD.n1439 0.0164828
R42315 VDD.n1131 VDD.n1130 0.0164828
R42316 VDD.n1129 VDD.n1128 0.0164828
R42317 VDD.n1127 VDD.n1126 0.0164828
R42318 VDD.n1125 VDD.n1124 0.0164828
R42319 VDD.n872 VDD.n871 0.0164828
R42320 VDD.n870 VDD.n869 0.0164828
R42321 VDD.n868 VDD.n867 0.0164828
R42322 VDD.n866 VDD.n865 0.0164828
R42323 VDD.n801 VDD.n800 0.0164828
R42324 VDD.n799 VDD.n798 0.0164828
R42325 VDD.n797 VDD.n796 0.0164828
R42326 VDD.n795 VDD.n794 0.0164828
R42327 VDD.n1326 VDD.n1325 0.0164828
R42328 VDD.n1328 VDD.n1327 0.0164828
R42329 VDD.n1330 VDD.n1329 0.0164828
R42330 VDD.n1332 VDD.n1331 0.0164828
R42331 VDD.n838 VDD.n837 0.0164828
R42332 VDD.n836 VDD.n835 0.0164828
R42333 VDD.n834 VDD.n833 0.0164828
R42334 VDD.n832 VDD.n831 0.0164828
R42335 VDD.n1373 VDD.n1372 0.0164828
R42336 VDD.n1375 VDD.n1374 0.0164828
R42337 VDD.n1377 VDD.n1376 0.0164828
R42338 VDD.n1379 VDD.n1378 0.0164828
R42339 VDD.n1265 VDD.n1264 0.0164828
R42340 VDD.n1263 VDD.n1262 0.0164828
R42341 VDD.n1261 VDD.n1260 0.0164828
R42342 VDD.n1259 VDD.n1258 0.0164828
R42343 VDD.n1617 VDD.n1616 0.0164828
R42344 VDD.n1615 VDD.n1614 0.0164828
R42345 VDD.n1613 VDD.n1612 0.0164828
R42346 VDD.n1232 VDD.n1231 0.0164828
R42347 VDD.n1230 VDD.n1229 0.0164828
R42348 VDD.n1228 VDD.n1227 0.0164828
R42349 VDD.n1226 VDD.n1225 0.0164828
R42350 VDD.n1099 VDD.n1098 0.0164828
R42351 VDD.n1097 VDD.n1096 0.0164828
R42352 VDD.n1095 VDD.n813 0.0164828
R42353 VDD.n1475 VDD.n1474 0.0164828
R42354 VDD.n1473 VDD.n1472 0.0164828
R42355 VDD.n1471 VDD.n1470 0.0164828
R42356 VDD.n1469 VDD.n1468 0.0164828
R42357 VDD.n1294 VDD.n1293 0.0164828
R42358 VDD.n1296 VDD.n1295 0.0164828
R42359 VDD.n1298 VDD.n1297 0.0164828
R42360 VDD.n1300 VDD.n1299 0.0164828
R42361 VDD.n1706 VDD.n1705 0.0164828
R42362 VDD.n1704 VDD.n1703 0.0164828
R42363 VDD.n1702 VDD.n1701 0.0164828
R42364 VDD.n1700 VDD.n1699 0.0164828
R42365 VDD.n887 VDD.n886 0.0164828
R42366 VDD.n889 VDD.n888 0.0164828
R42367 VDD.n891 VDD.n890 0.0164828
R42368 VDD.n893 VDD.n892 0.0164828
R42369 VDD.n929 VDD.n928 0.0164828
R42370 VDD.n931 VDD.n930 0.0164828
R42371 VDD.n933 VDD.n932 0.0164828
R42372 VDD.n935 VDD.n934 0.0164828
R42373 VDD.n1049 VDD.n1048 0.0164828
R42374 VDD.n1051 VDD.n1050 0.0164828
R42375 VDD.n1053 VDD.n1052 0.0164828
R42376 VDD.n1055 VDD.n1054 0.0164828
R42377 VDD.n1153 VDD.n1152 0.0164828
R42378 VDD.n1151 VDD.n1150 0.0164828
R42379 VDD.n1149 VDD.n1148 0.0164828
R42380 VDD.n1147 VDD.n1146 0.0164828
R42381 VDD.n1724 VDD.n1723 0.0164828
R42382 VDD.n1726 VDD.n1725 0.0164828
R42383 VDD.n1728 VDD.n1727 0.0164828
R42384 VDD.n1730 VDD.n1729 0.0164828
R42385 VDD.n2136 VDD.n2135 0.0163144
R42386 VDD.n5253 VDD.n5252 0.01631
R42387 VDD.n5245 VDD.n5244 0.01631
R42388 VDD.n5463 VDD.n5462 0.01631
R42389 VDD.n5455 VDD.n5454 0.01631
R42390 VDD.n5352 VDD.n5351 0.01631
R42391 VDD.n5344 VDD.n5343 0.01631
R42392 VDD.n5998 VDD.n5997 0.01631
R42393 VDD.n6390 VDD.n6389 0.01631
R42394 VDD.n6342 VDD.n6341 0.01631
R42395 VDD.n6350 VDD.n6349 0.01631
R42396 VDD.n7154 VDD.n7153 0.01631
R42397 VDD.n7162 VDD.n7161 0.01631
R42398 VDD.n5424 VDD.n5423 0.01631
R42399 VDD.n5416 VDD.n5415 0.01631
R42400 VDD.n7114 VDD.n7113 0.01631
R42401 VDD.n7106 VDD.n7105 0.01631
R42402 VDD.n6562 VDD.n5287 0.0162238
R42403 VDD.n5298 VDD.n5297 0.0162238
R42404 VDD.n2385 VDD.n2384 0.0162238
R42405 VDD.n7025 VDD.n2374 0.0162238
R42406 VDD.n5363 VDD.n5362 0.0159138
R42407 VDD.n5365 VDD.n5364 0.0159138
R42408 VDD.n5367 VDD.n5366 0.0159138
R42409 VDD.n5370 VDD.n5369 0.0159138
R42410 VDD.n5372 VDD.n5371 0.0159138
R42411 VDD.n5374 VDD.n5373 0.0159138
R42412 VDD.n6378 VDD.n6377 0.0159138
R42413 VDD.n6376 VDD.n6375 0.0159138
R42414 VDD.n6374 VDD.n6373 0.0159138
R42415 VDD.n6216 VDD.n5375 0.0159138
R42416 VDD.n6218 VDD.n6217 0.0159138
R42417 VDD.n6265 VDD.n6264 0.0159138
R42418 VDD.n6263 VDD.n5377 0.0159138
R42419 VDD.n6367 VDD.n6366 0.0159138
R42420 VDD.n6365 VDD.n6364 0.0159138
R42421 VDD.n6363 VDD.n6362 0.0159138
R42422 VDD.n5937 VDD.n5473 0.0159138
R42423 VDD.n5939 VDD.n5938 0.0159138
R42424 VDD.n5941 VDD.n5940 0.0159138
R42425 VDD.n5945 VDD.n5944 0.0159138
R42426 VDD.n5947 VDD.n5946 0.0159138
R42427 VDD.n5949 VDD.n5948 0.0159138
R42428 VDD.n2358 VDD.n2341 0.0159138
R42429 VDD.n2360 VDD.n2359 0.0159138
R42430 VDD.n2365 VDD.n2364 0.0159138
R42431 VDD.n2363 VDD.n2362 0.0159138
R42432 VDD.n2361 VDD.n2311 0.0159138
R42433 VDD.n7141 VDD.n7140 0.0159138
R42434 VDD.n7139 VDD.n7138 0.0159138
R42435 VDD.n7137 VDD.n7136 0.0159138
R42436 VDD.n2316 VDD.n2315 0.0159138
R42437 VDD.n2314 VDD.n2313 0.0159138
R42438 VDD.n2401 VDD.n2400 0.0159138
R42439 VDD.n2399 VDD.n2398 0.0159138
R42440 VDD.n2397 VDD.n2320 0.0159138
R42441 VDD.n7130 VDD.n7129 0.0159138
R42442 VDD.n7128 VDD.n7127 0.0159138
R42443 VDD.n7126 VDD.n7125 0.0159138
R42444 VDD.n2343 VDD.n2323 0.0159138
R42445 VDD.n2345 VDD.n2344 0.0159138
R42446 VDD.n2347 VDD.n2346 0.0159138
R42447 VDD.n7045 VDD.n7044 0.0159138
R42448 VDD.n7047 VDD.n7046 0.0159138
R42449 VDD.n1205 VDD.n1204 0.0159138
R42450 VDD.n1203 VDD.n1190 0.0159138
R42451 VDD.n1202 VDD.n1190 0.0159138
R42452 VDD.n1201 VDD.n1191 0.0159138
R42453 VDD.n1200 VDD.n1191 0.0159138
R42454 VDD.n1199 VDD.n1192 0.0159138
R42455 VDD.n1198 VDD.n1192 0.0159138
R42456 VDD.n1197 VDD.n1193 0.0159138
R42457 VDD.n1196 VDD.n1193 0.0159138
R42458 VDD.n1195 VDD.n1194 0.0159138
R42459 VDD.n1194 VDD.n851 0.0159138
R42460 VDD.n1432 VDD.n843 0.0159138
R42461 VDD.n1433 VDD.n843 0.0159138
R42462 VDD.n1434 VDD.n842 0.0159138
R42463 VDD.n1435 VDD.n842 0.0159138
R42464 VDD.n1436 VDD.n841 0.0159138
R42465 VDD.n1437 VDD.n841 0.0159138
R42466 VDD.n1438 VDD.n840 0.0159138
R42467 VDD.n1439 VDD.n840 0.0159138
R42468 VDD.n1134 VDD.n1133 0.0159138
R42469 VDD.n1132 VDD.n1119 0.0159138
R42470 VDD.n1131 VDD.n1119 0.0159138
R42471 VDD.n1130 VDD.n1120 0.0159138
R42472 VDD.n1129 VDD.n1120 0.0159138
R42473 VDD.n1128 VDD.n1121 0.0159138
R42474 VDD.n1127 VDD.n1121 0.0159138
R42475 VDD.n1126 VDD.n1122 0.0159138
R42476 VDD.n1125 VDD.n1122 0.0159138
R42477 VDD.n1124 VDD.n1123 0.0159138
R42478 VDD.n1123 VDD.n852 0.0159138
R42479 VDD.n873 VDD.n860 0.0159138
R42480 VDD.n872 VDD.n860 0.0159138
R42481 VDD.n871 VDD.n861 0.0159138
R42482 VDD.n870 VDD.n861 0.0159138
R42483 VDD.n869 VDD.n862 0.0159138
R42484 VDD.n868 VDD.n862 0.0159138
R42485 VDD.n867 VDD.n863 0.0159138
R42486 VDD.n866 VDD.n863 0.0159138
R42487 VDD.n865 VDD.n864 0.0159138
R42488 VDD.n864 VDD.n728 0.0159138
R42489 VDD.n802 VDD.n788 0.0159138
R42490 VDD.n801 VDD.n788 0.0159138
R42491 VDD.n800 VDD.n789 0.0159138
R42492 VDD.n799 VDD.n789 0.0159138
R42493 VDD.n798 VDD.n790 0.0159138
R42494 VDD.n797 VDD.n790 0.0159138
R42495 VDD.n796 VDD.n791 0.0159138
R42496 VDD.n795 VDD.n791 0.0159138
R42497 VDD.n794 VDD.n792 0.0159138
R42498 VDD.n793 VDD.n792 0.0159138
R42499 VDD.n1324 VDD.n745 0.0159138
R42500 VDD.n1325 VDD.n1324 0.0159138
R42501 VDD.n1326 VDD.n1323 0.0159138
R42502 VDD.n1327 VDD.n1323 0.0159138
R42503 VDD.n1328 VDD.n1322 0.0159138
R42504 VDD.n1329 VDD.n1322 0.0159138
R42505 VDD.n1330 VDD.n1321 0.0159138
R42506 VDD.n1331 VDD.n1321 0.0159138
R42507 VDD.n1332 VDD.n1320 0.0159138
R42508 VDD.n1333 VDD.n1320 0.0159138
R42509 VDD.n1334 VDD.n1319 0.0159138
R42510 VDD.n839 VDD.n825 0.0159138
R42511 VDD.n838 VDD.n825 0.0159138
R42512 VDD.n837 VDD.n826 0.0159138
R42513 VDD.n836 VDD.n826 0.0159138
R42514 VDD.n835 VDD.n827 0.0159138
R42515 VDD.n834 VDD.n827 0.0159138
R42516 VDD.n833 VDD.n828 0.0159138
R42517 VDD.n832 VDD.n828 0.0159138
R42518 VDD.n831 VDD.n829 0.0159138
R42519 VDD.n830 VDD.n829 0.0159138
R42520 VDD.n1371 VDD.n1370 0.0159138
R42521 VDD.n1372 VDD.n1370 0.0159138
R42522 VDD.n1373 VDD.n1369 0.0159138
R42523 VDD.n1374 VDD.n1369 0.0159138
R42524 VDD.n1375 VDD.n1368 0.0159138
R42525 VDD.n1376 VDD.n1368 0.0159138
R42526 VDD.n1377 VDD.n1367 0.0159138
R42527 VDD.n1378 VDD.n1367 0.0159138
R42528 VDD.n1379 VDD.n1366 0.0159138
R42529 VDD.n1380 VDD.n1366 0.0159138
R42530 VDD.n1381 VDD.n1365 0.0159138
R42531 VDD.n1268 VDD.n1267 0.0159138
R42532 VDD.n1266 VDD.n1252 0.0159138
R42533 VDD.n1265 VDD.n1252 0.0159138
R42534 VDD.n1264 VDD.n1253 0.0159138
R42535 VDD.n1263 VDD.n1253 0.0159138
R42536 VDD.n1262 VDD.n1254 0.0159138
R42537 VDD.n1261 VDD.n1254 0.0159138
R42538 VDD.n1260 VDD.n1255 0.0159138
R42539 VDD.n1259 VDD.n1255 0.0159138
R42540 VDD.n1258 VDD.n1256 0.0159138
R42541 VDD.n1257 VDD.n1256 0.0159138
R42542 VDD.n1618 VDD.n785 0.0159138
R42543 VDD.n1617 VDD.n785 0.0159138
R42544 VDD.n1616 VDD.n786 0.0159138
R42545 VDD.n1615 VDD.n786 0.0159138
R42546 VDD.n1614 VDD.n787 0.0159138
R42547 VDD.n1613 VDD.n787 0.0159138
R42548 VDD.n1235 VDD.n1234 0.0159138
R42549 VDD.n1233 VDD.n1220 0.0159138
R42550 VDD.n1232 VDD.n1220 0.0159138
R42551 VDD.n1231 VDD.n1221 0.0159138
R42552 VDD.n1230 VDD.n1221 0.0159138
R42553 VDD.n1229 VDD.n1222 0.0159138
R42554 VDD.n1228 VDD.n1222 0.0159138
R42555 VDD.n1227 VDD.n1223 0.0159138
R42556 VDD.n1226 VDD.n1223 0.0159138
R42557 VDD.n1225 VDD.n1224 0.0159138
R42558 VDD.n1224 VDD.n1085 0.0159138
R42559 VDD.n1100 VDD.n1092 0.0159138
R42560 VDD.n1099 VDD.n1092 0.0159138
R42561 VDD.n1098 VDD.n1093 0.0159138
R42562 VDD.n1097 VDD.n1093 0.0159138
R42563 VDD.n1096 VDD.n1094 0.0159138
R42564 VDD.n1095 VDD.n1094 0.0159138
R42565 VDD.n1476 VDD.n1462 0.0159138
R42566 VDD.n1475 VDD.n1462 0.0159138
R42567 VDD.n1474 VDD.n1463 0.0159138
R42568 VDD.n1473 VDD.n1463 0.0159138
R42569 VDD.n1472 VDD.n1464 0.0159138
R42570 VDD.n1471 VDD.n1464 0.0159138
R42571 VDD.n1470 VDD.n1465 0.0159138
R42572 VDD.n1469 VDD.n1465 0.0159138
R42573 VDD.n1468 VDD.n1466 0.0159138
R42574 VDD.n1467 VDD.n1466 0.0159138
R42575 VDD.n1292 VDD.n742 0.0159138
R42576 VDD.n1293 VDD.n1292 0.0159138
R42577 VDD.n1294 VDD.n1291 0.0159138
R42578 VDD.n1295 VDD.n1291 0.0159138
R42579 VDD.n1296 VDD.n1290 0.0159138
R42580 VDD.n1297 VDD.n1290 0.0159138
R42581 VDD.n1298 VDD.n1289 0.0159138
R42582 VDD.n1299 VDD.n1289 0.0159138
R42583 VDD.n1300 VDD.n1288 0.0159138
R42584 VDD.n1301 VDD.n1288 0.0159138
R42585 VDD.n1302 VDD.n1287 0.0159138
R42586 VDD.n1707 VDD.n730 0.0159138
R42587 VDD.n1706 VDD.n730 0.0159138
R42588 VDD.n1705 VDD.n731 0.0159138
R42589 VDD.n1704 VDD.n731 0.0159138
R42590 VDD.n1703 VDD.n732 0.0159138
R42591 VDD.n1702 VDD.n732 0.0159138
R42592 VDD.n1701 VDD.n733 0.0159138
R42593 VDD.n1700 VDD.n733 0.0159138
R42594 VDD.n1699 VDD.n734 0.0159138
R42595 VDD.n1698 VDD.n734 0.0159138
R42596 VDD.n885 VDD.n884 0.0159138
R42597 VDD.n886 VDD.n884 0.0159138
R42598 VDD.n887 VDD.n883 0.0159138
R42599 VDD.n888 VDD.n883 0.0159138
R42600 VDD.n889 VDD.n882 0.0159138
R42601 VDD.n890 VDD.n882 0.0159138
R42602 VDD.n891 VDD.n881 0.0159138
R42603 VDD.n892 VDD.n881 0.0159138
R42604 VDD.n893 VDD.n880 0.0159138
R42605 VDD.n894 VDD.n880 0.0159138
R42606 VDD.n895 VDD.n879 0.0159138
R42607 VDD.n927 VDD.n699 0.0159138
R42608 VDD.n928 VDD.n927 0.0159138
R42609 VDD.n929 VDD.n926 0.0159138
R42610 VDD.n930 VDD.n926 0.0159138
R42611 VDD.n931 VDD.n925 0.0159138
R42612 VDD.n932 VDD.n925 0.0159138
R42613 VDD.n933 VDD.n924 0.0159138
R42614 VDD.n934 VDD.n924 0.0159138
R42615 VDD.n935 VDD.n923 0.0159138
R42616 VDD.n936 VDD.n923 0.0159138
R42617 VDD.n1047 VDD.n922 0.0159138
R42618 VDD.n1048 VDD.n922 0.0159138
R42619 VDD.n1049 VDD.n921 0.0159138
R42620 VDD.n1050 VDD.n921 0.0159138
R42621 VDD.n1051 VDD.n920 0.0159138
R42622 VDD.n1052 VDD.n920 0.0159138
R42623 VDD.n1053 VDD.n919 0.0159138
R42624 VDD.n1054 VDD.n919 0.0159138
R42625 VDD.n1055 VDD.n918 0.0159138
R42626 VDD.n1056 VDD.n918 0.0159138
R42627 VDD.n1057 VDD.n917 0.0159138
R42628 VDD.n1156 VDD.n1155 0.0159138
R42629 VDD.n1154 VDD.n1140 0.0159138
R42630 VDD.n1153 VDD.n1140 0.0159138
R42631 VDD.n1152 VDD.n1141 0.0159138
R42632 VDD.n1151 VDD.n1141 0.0159138
R42633 VDD.n1150 VDD.n1142 0.0159138
R42634 VDD.n1149 VDD.n1142 0.0159138
R42635 VDD.n1148 VDD.n1143 0.0159138
R42636 VDD.n1147 VDD.n1143 0.0159138
R42637 VDD.n1146 VDD.n1144 0.0159138
R42638 VDD.n1145 VDD.n1144 0.0159138
R42639 VDD.n1722 VDD.n705 0.0159138
R42640 VDD.n1723 VDD.n705 0.0159138
R42641 VDD.n1724 VDD.n704 0.0159138
R42642 VDD.n1725 VDD.n704 0.0159138
R42643 VDD.n1726 VDD.n703 0.0159138
R42644 VDD.n1727 VDD.n703 0.0159138
R42645 VDD.n1728 VDD.n702 0.0159138
R42646 VDD.n1729 VDD.n702 0.0159138
R42647 VDD.n1730 VDD.n701 0.0159138
R42648 VDD.n1731 VDD.n701 0.0159138
R42649 VDD.n8137 VDD.n8136 0.0159011
R42650 VDD.n8116 VDD.n8115 0.0159011
R42651 VDD.n8104 VDD.n8103 0.0159011
R42652 VDD.n5580 VDD.n5579 0.0159011
R42653 VDD.n5601 VDD.n5600 0.0159011
R42654 VDD.n5622 VDD.n5621 0.0159011
R42655 VDD.n5662 VDD.n5661 0.0159011
R42656 VDD.n5871 VDD.n5870 0.0159011
R42657 VDD.n5859 VDD.n5858 0.0159011
R42658 VDD.n5816 VDD.n5815 0.0159011
R42659 VDD.n5804 VDD.n5803 0.0159011
R42660 VDD.n5783 VDD.n5782 0.0159011
R42661 VDD.n5749 VDD.n5748 0.0159011
R42662 VDD.n5728 VDD.n5727 0.0159011
R42663 VDD.n11032 VDD.n11031 0.0159011
R42664 VDD.n9037 VDD.n8490 0.0159011
R42665 VDD.n9008 VDD.n8951 0.0159011
R42666 VDD.n8940 VDD.n8507 0.0159011
R42667 VDD.n8877 VDD.n8842 0.0159011
R42668 VDD.n8809 VDD.n8526 0.0159011
R42669 VDD.n8554 VDD.n8553 0.0159011
R42670 VDD.n175 VDD.n174 0.0159011
R42671 VDD.n9096 VDD.n9095 0.0159011
R42672 VDD.n9161 VDD.n8472 0.0159011
R42673 VDD.n141 VDD.n140 0.0159011
R42674 VDD.n12494 VDD.n12493 0.0159011
R42675 VDD.n95 VDD.n94 0.0159011
R42676 VDD.n52 VDD.n51 0.0159011
R42677 VDD.n12550 VDD.n12549 0.0159011
R42678 VDD.n12593 VDD.n12591 0.0159011
R42679 VDD.n10149 VDD.n10148 0.015875
R42680 VDD.n2134 VDD.n2133 0.0156839
R42681 VDD.n2137 VDD.n2136 0.0154737
R42682 VDD.n6180 VDD.n6179 0.0154453
R42683 VDD.n6320 VDD.n6318 0.0153631
R42684 VDD.n5250 VDD.n5249 0.015256
R42685 VDD.n5460 VDD.n5459 0.015256
R42686 VDD.n5349 VDD.n5348 0.015256
R42687 VDD.n6394 VDD.n5313 0.015256
R42688 VDD.n6344 VDD.n5481 0.015256
R42689 VDD.n7156 VDD.n2305 0.015256
R42690 VDD.n5421 VDD.n5420 0.015256
R42691 VDD.n7111 VDD.n7110 0.015256
R42692 VDD.n2163 VDD.n2162 0.0148793
R42693 VDD.n1548 VDD.n1533 0.014653
R42694 VDD.n1495 VDD.n1494 0.0142459
R42695 VDD.n1607 VDD.n1606 0.0142459
R42696 VDD.n1595 VDD.n1594 0.0142459
R42697 VDD.n1711 VDD.n1710 0.0142459
R42698 VDD.n1398 VDD.n1397 0.0142459
R42699 VDD.n1407 VDD.n1406 0.0142459
R42700 VDD.n1445 VDD.n1444 0.0142459
R42701 VDD.n1460 VDD.n1459 0.0142459
R42702 VDD.n1483 VDD.n1482 0.0142459
R42703 VDD.n1735 VDD.n1734 0.0142459
R42704 VDD.n720 VDD.n719 0.0142459
R42705 VDD.n2161 VDD.n2160 0.0142069
R42706 VDD.n6714 VDD.n2406 0.0141364
R42707 VDD.n6700 VDD.n6699 0.0138734
R42708 VDD.n5444 VDD.n5438 0.0138734
R42709 VDD.n8015 VDD.n8014 0.0138448
R42710 VDD.n6699 VDD.n6698 0.0138425
R42711 VDD.n5444 VDD.n5443 0.0138425
R42712 VDD.n1559 VDD.n1558 0.0137787
R42713 VDD.n1554 VDD.n1517 0.0137787
R42714 VDD.n6190 VDD.n6010 0.0137336
R42715 VDD.n5487 VDD.n5486 0.0137336
R42716 VDD.n10777 VDD.n2020 0.0136837
R42717 VDD.n10784 VDD.n2010 0.0136837
R42718 VDD.n10835 VDD.n1947 0.0136837
R42719 VDD.n10842 VDD.n1937 0.0136837
R42720 VDD.n10897 VDD.n1910 0.0136837
R42721 VDD.n10945 VDD.n1855 0.0136837
R42722 VDD.n10952 VDD.n1845 0.0136837
R42723 VDD.n11000 VDD.n1790 0.0136837
R42724 VDD.n11007 VDD.n1783 0.0136837
R42725 VDD.n9053 VDD.n9052 0.0136837
R42726 VDD.n8919 VDD.n8918 0.0136837
R42727 VDD.n8861 VDD.n8858 0.0136837
R42728 VDD.n8570 VDD.n8569 0.0136837
R42729 VDD.n9177 VDD.n9176 0.0136837
R42730 VDD.n12459 VDD.n12458 0.0136837
R42731 VDD.n12477 VDD.n12474 0.0136837
R42732 VDD.n12515 VDD.n12514 0.0136837
R42733 VDD.n12533 VDD.n12530 0.0136837
R42734 VDD.n12609 VDD.n12608 0.0136837
R42735 VDD.n10828 VDD.n1993 0.013561
R42736 VDD.n10883 VDD.n1928 0.013561
R42737 VDD.n10938 VDD.n1901 0.013561
R42738 VDD.n10993 VDD.n1836 0.013561
R42739 VDD.n8988 VDD.n8985 0.013561
R42740 VDD.n8788 VDD.n8787 0.013561
R42741 VDD.n12467 VDD.n122 0.013561
R42742 VDD.n12523 VDD.n42 0.013561
R42743 VDD.n1537 VDD.n1512 0.0133852
R42744 VDD.n1553 VDD.n1518 0.0133852
R42745 VDD.n1752 VDD.n682 0.0131331
R42746 VDD.n996 VDD.n995 0.0131331
R42747 VDD.n1007 VDD.n1006 0.0131331
R42748 VDD.n7822 VDD.n2242 0.012875
R42749 VDD.n11872 VDD.n384 0.012875
R42750 VDD.n6601 VDD.n6599 0.012725
R42751 VDD.n952 VDD.n951 0.0126485
R42752 VDD.n6709 VDD.n6708 0.0125453
R42753 VDD.n6704 VDD.n6703 0.0125453
R42754 VDD.n6695 VDD.n6694 0.0125453
R42755 VDD.n6690 VDD.n6689 0.0125453
R42756 VDD.n6638 VDD.n6637 0.0125453
R42757 VDD.n5435 VDD.n5434 0.0125453
R42758 VDD.n5440 VDD.n5439 0.0125453
R42759 VDD.n6629 VDD.n6628 0.0125453
R42760 VDD.n1495 VDD.n805 0.0124383
R42761 VDD.n1496 VDD.n805 0.0124383
R42762 VDD.n1608 VDD.n1497 0.0124383
R42763 VDD.n1607 VDD.n1497 0.0124383
R42764 VDD.n1606 VDD.n1498 0.0124383
R42765 VDD.n1605 VDD.n1498 0.0124383
R42766 VDD.n1604 VDD.n1499 0.0124383
R42767 VDD.n1602 VDD.n1499 0.0124383
R42768 VDD.n1602 VDD.n1601 0.0124383
R42769 VDD.n1599 VDD.n1502 0.0124383
R42770 VDD.n1597 VDD.n1502 0.0124383
R42771 VDD.n1596 VDD.n1503 0.0124383
R42772 VDD.n1595 VDD.n1503 0.0124383
R42773 VDD.n1594 VDD.n1504 0.0124383
R42774 VDD.n1710 VDD.n727 0.0124383
R42775 VDD.n1709 VDD.n727 0.0124383
R42776 VDD.n1396 VDD.n729 0.0124383
R42777 VDD.n1397 VDD.n1396 0.0124383
R42778 VDD.n1398 VDD.n1395 0.0124383
R42779 VDD.n1399 VDD.n1395 0.0124383
R42780 VDD.n1400 VDD.n1394 0.0124383
R42781 VDD.n1402 VDD.n1394 0.0124383
R42782 VDD.n1402 VDD.n1391 0.0124383
R42783 VDD.n1411 VDD.n1393 0.0124383
R42784 VDD.n1409 VDD.n1393 0.0124383
R42785 VDD.n1408 VDD.n1404 0.0124383
R42786 VDD.n1407 VDD.n1404 0.0124383
R42787 VDD.n1406 VDD.n1405 0.0124383
R42788 VDD.n1405 VDD.n824 0.0124383
R42789 VDD.n1443 VDD.n822 0.0124383
R42790 VDD.n1444 VDD.n822 0.0124383
R42791 VDD.n1446 VDD.n1445 0.0124383
R42792 VDD.n1450 VDD.n819 0.0124383
R42793 VDD.n1452 VDD.n819 0.0124383
R42794 VDD.n1452 VDD.n820 0.0124383
R42795 VDD.n1455 VDD.n817 0.0124383
R42796 VDD.n1457 VDD.n817 0.0124383
R42797 VDD.n1458 VDD.n816 0.0124383
R42798 VDD.n1459 VDD.n816 0.0124383
R42799 VDD.n1460 VDD.n815 0.0124383
R42800 VDD.n1461 VDD.n815 0.0124383
R42801 VDD.n1481 VDD.n812 0.0124383
R42802 VDD.n1482 VDD.n812 0.0124383
R42803 VDD.n1483 VDD.n811 0.0124383
R42804 VDD.n1484 VDD.n811 0.0124383
R42805 VDD.n1485 VDD.n809 0.0124383
R42806 VDD.n1487 VDD.n809 0.0124383
R42807 VDD.n1487 VDD.n810 0.0124383
R42808 VDD.n1490 VDD.n807 0.0124383
R42809 VDD.n1492 VDD.n807 0.0124383
R42810 VDD.n1493 VDD.n806 0.0124383
R42811 VDD.n1494 VDD.n806 0.0124383
R42812 VDD.n951 VDD.n943 0.0124383
R42813 VDD.n950 VDD.n943 0.0124383
R42814 VDD.n948 VDD.n944 0.0124383
R42815 VDD.n946 VDD.n944 0.0124383
R42816 VDD.n946 VDD.n693 0.0124383
R42817 VDD.n1739 VDD.n695 0.0124383
R42818 VDD.n1737 VDD.n695 0.0124383
R42819 VDD.n1735 VDD.n697 0.0124383
R42820 VDD.n1734 VDD.n698 0.0124383
R42821 VDD.n1733 VDD.n698 0.0124383
R42822 VDD.n718 VDD.n700 0.0124383
R42823 VDD.n719 VDD.n718 0.0124383
R42824 VDD.n720 VDD.n717 0.0124383
R42825 VDD.n721 VDD.n717 0.0124383
R42826 VDD.n722 VDD.n716 0.0124383
R42827 VDD.n724 VDD.n716 0.0124383
R42828 VDD.n724 VDD.n713 0.0124383
R42829 VDD.n1715 VDD.n715 0.0124383
R42830 VDD.n1713 VDD.n715 0.0124383
R42831 VDD.n1712 VDD.n726 0.0124383
R42832 VDD.n1711 VDD.n726 0.0124383
R42833 VDD.n9183 VDD.n8459 0.0123552
R42834 VDD.n1005 VDD.n1004 0.0120089
R42835 VDD.n2138 VDD.n2137 0.0119536
R42836 VDD.n2135 VDD.n2134 0.0119536
R42837 VDD.n2133 VDD.n2132 0.0119536
R42838 VDD.n1605 VDD.n1604 0.0118498
R42839 VDD.n1600 VDD.n1599 0.0118498
R42840 VDD.n1597 VDD.n1596 0.0118498
R42841 VDD.n1400 VDD.n1399 0.0118498
R42842 VDD.n1412 VDD.n1411 0.0118498
R42843 VDD.n1409 VDD.n1408 0.0118498
R42844 VDD.n1455 VDD.n818 0.0118498
R42845 VDD.n1458 VDD.n1457 0.0118498
R42846 VDD.n1485 VDD.n1484 0.0118498
R42847 VDD.n1490 VDD.n808 0.0118498
R42848 VDD.n1493 VDD.n1492 0.0118498
R42849 VDD.n1740 VDD.n1739 0.0118498
R42850 VDD.n1737 VDD.n1736 0.0118498
R42851 VDD.n722 VDD.n721 0.0118498
R42852 VDD.n1716 VDD.n1715 0.0118498
R42853 VDD.n1713 VDD.n1712 0.0118498
R42854 VDD.n8067 VDD.n8066 0.0117759
R42855 VDD.n2156 VDD.n2147 0.0117759
R42856 VDD.n2165 VDD.n2164 0.0117759
R42857 VDD.n8016 VDD.n8015 0.0117759
R42858 VDD.n2130 VDD.n2129 0.0116909
R42859 VDD.n1610 VDD.n1496 0.0115976
R42860 VDD.n1610 VDD.n1608 0.0115976
R42861 VDD.n1709 VDD.n1708 0.0115976
R42862 VDD.n1708 VDD.n729 0.0115976
R42863 VDD.n1442 VDD.n824 0.0115976
R42864 VDD.n1443 VDD.n1442 0.0115976
R42865 VDD.n1480 VDD.n1461 0.0115976
R42866 VDD.n1481 VDD.n1480 0.0115976
R42867 VDD.n1733 VDD.n1732 0.0115976
R42868 VDD.n1732 VDD.n700 0.0115976
R42869 VDD.n9134 VDD.n9133 0.0114862
R42870 VDD.n1022 VDD.n1 0.0114467
R42871 VDD.n6297 VDD.n6296 0.0113718
R42872 VDD.n6269 VDD.n6268 0.0113718
R42873 VDD.n6261 VDD.n6260 0.0113718
R42874 VDD.n6657 VDD.n6656 0.0113718
R42875 VDD.n7051 VDD.n7050 0.0113718
R42876 VDD.n10777 VDD.n2023 0.0113038
R42877 VDD.n10787 VDD.n10784 0.0113038
R42878 VDD.n10835 VDD.n1950 0.0113038
R42879 VDD.n10845 VDD.n10842 0.0113038
R42880 VDD.n10900 VDD.n10897 0.0113038
R42881 VDD.n10945 VDD.n1858 0.0113038
R42882 VDD.n10955 VDD.n10952 0.0113038
R42883 VDD.n11000 VDD.n1793 0.0113038
R42884 VDD.n11010 VDD.n11007 0.0113038
R42885 VDD.n9055 VDD.n9053 0.0113038
R42886 VDD.n8921 VDD.n8919 0.0113038
R42887 VDD.n8858 VDD.n8857 0.0113038
R42888 VDD.n8572 VDD.n8570 0.0113038
R42889 VDD.n9177 VDD.n8465 0.0113038
R42890 VDD.n12459 VDD.n180 0.0113038
R42891 VDD.n12474 VDD.n109 0.0113038
R42892 VDD.n12515 VDD.n100 0.0113038
R42893 VDD.n12530 VDD.n29 0.0113038
R42894 VDD.n12609 VDD.n20 0.0113038
R42895 VDD.n10828 VDD.n10827 0.0112032
R42896 VDD.n10883 VDD.n10882 0.0112032
R42897 VDD.n10938 VDD.n10937 0.0112032
R42898 VDD.n10993 VDD.n10992 0.0112032
R42899 VDD.n8985 VDD.n8984 0.0112032
R42900 VDD.n8790 VDD.n8788 0.0112032
R42901 VDD.n12467 VDD.n119 0.0112032
R42902 VDD.n12523 VDD.n39 0.0112032
R42903 VDD.n2158 VDD.n2157 0.0111034
R42904 VDD.n8142 VDD.n8141 0.0109679
R42905 VDD.n5555 VDD.n5554 0.0109679
R42906 VDD.n5546 VDD.n5545 0.0109679
R42907 VDD.n5821 VDD.n5820 0.0109679
R42908 VDD.n5754 VDD.n5753 0.0109679
R42909 VDD.n9002 VDD.n8970 0.0109679
R42910 VDD.n8831 VDD.n8830 0.0109679
R42911 VDD.n9118 VDD.n9117 0.0109679
R42912 VDD.n163 VDD.n162 0.0109679
R42913 VDD.n74 VDD.n73 0.0109679
R42914 VDD.n5202 VDD.n5201 0.0109148
R42915 VDD.n5201 VDD.n2408 0.0109148
R42916 VDD.n1569 VDD.n1568 0.0108543
R42917 VDD.n7175 VDD.n7174 0.0108058
R42918 VDD.n7827 VDD.n2241 0.0108058
R42919 VDD.n1661 VDD.n754 0.0106739
R42920 VDD.n1643 VDD.n768 0.0106739
R42921 VDD.n1447 VDD.n1446 0.0102524
R42922 VDD.n6685 VDD.n5265 0.0101084
R42923 VDD.n6685 VDD.n6684 0.0101084
R42924 VDD.n7760 VDD.n2265 0.0101084
R42925 VDD.n6297 VDD.n6200 0.00994219
R42926 VDD.n6296 VDD.n6201 0.00994219
R42927 VDD.n6294 VDD.n6201 0.00994219
R42928 VDD.n6294 VDD.n6293 0.00994219
R42929 VDD.n6293 VDD.n6292 0.00994219
R42930 VDD.n6292 VDD.n6204 0.00994219
R42931 VDD.n6289 VDD.n6204 0.00994219
R42932 VDD.n6289 VDD.n6288 0.00994219
R42933 VDD.n6288 VDD.n6287 0.00994219
R42934 VDD.n6286 VDD.n6206 0.00994219
R42935 VDD.n6284 VDD.n6206 0.00994219
R42936 VDD.n6282 VDD.n6281 0.00994219
R42937 VDD.n6281 VDD.n6209 0.00994219
R42938 VDD.n6279 VDD.n6209 0.00994219
R42939 VDD.n6278 VDD.n6210 0.00994219
R42940 VDD.n6276 VDD.n6210 0.00994219
R42941 VDD.n6276 VDD.n6275 0.00994219
R42942 VDD.n6275 VDD.n6274 0.00994219
R42943 VDD.n6274 VDD.n6213 0.00994219
R42944 VDD.n6271 VDD.n6213 0.00994219
R42945 VDD.n6271 VDD.n6270 0.00994219
R42946 VDD.n6270 VDD.n6269 0.00994219
R42947 VDD.n6268 VDD.n6215 0.00994219
R42948 VDD.n6267 VDD.n6215 0.00994219
R42949 VDD.n6262 VDD.n6219 0.00994219
R42950 VDD.n6261 VDD.n6219 0.00994219
R42951 VDD.n6260 VDD.n6220 0.00994219
R42952 VDD.n6258 VDD.n6220 0.00994219
R42953 VDD.n6258 VDD.n6257 0.00994219
R42954 VDD.n6257 VDD.n6256 0.00994219
R42955 VDD.n6256 VDD.n6223 0.00994219
R42956 VDD.n6253 VDD.n6223 0.00994219
R42957 VDD.n6253 VDD.n6252 0.00994219
R42958 VDD.n6252 VDD.n6251 0.00994219
R42959 VDD.n6250 VDD.n6225 0.00994219
R42960 VDD.n6248 VDD.n6225 0.00994219
R42961 VDD.n6246 VDD.n6245 0.00994219
R42962 VDD.n6245 VDD.n6228 0.00994219
R42963 VDD.n6243 VDD.n6228 0.00994219
R42964 VDD.n6242 VDD.n6229 0.00994219
R42965 VDD.n6240 VDD.n6229 0.00994219
R42966 VDD.n6240 VDD.n6239 0.00994219
R42967 VDD.n6239 VDD.n6238 0.00994219
R42968 VDD.n6238 VDD.n6232 0.00994219
R42969 VDD.n6235 VDD.n6232 0.00994219
R42970 VDD.n6235 VDD.n6234 0.00994219
R42971 VDD.n6234 VDD.n5265 0.00994219
R42972 VDD.n6684 VDD.n6642 0.00994219
R42973 VDD.n6682 VDD.n6642 0.00994219
R42974 VDD.n6682 VDD.n6681 0.00994219
R42975 VDD.n6681 VDD.n6680 0.00994219
R42976 VDD.n6680 VDD.n6645 0.00994219
R42977 VDD.n6677 VDD.n6645 0.00994219
R42978 VDD.n6677 VDD.n6676 0.00994219
R42979 VDD.n6676 VDD.n6675 0.00994219
R42980 VDD.n6674 VDD.n6647 0.00994219
R42981 VDD.n6672 VDD.n6647 0.00994219
R42982 VDD.n6669 VDD.n6648 0.00994219
R42983 VDD.n6669 VDD.n6649 0.00994219
R42984 VDD.n6667 VDD.n6649 0.00994219
R42985 VDD.n6666 VDD.n6650 0.00994219
R42986 VDD.n6664 VDD.n6650 0.00994219
R42987 VDD.n6664 VDD.n6663 0.00994219
R42988 VDD.n6663 VDD.n6662 0.00994219
R42989 VDD.n6662 VDD.n6653 0.00994219
R42990 VDD.n6659 VDD.n6653 0.00994219
R42991 VDD.n6659 VDD.n6658 0.00994219
R42992 VDD.n6658 VDD.n6657 0.00994219
R42993 VDD.n6656 VDD.n6655 0.00994219
R42994 VDD.n6655 VDD.n2342 0.00994219
R42995 VDD.n7049 VDD.n2340 0.00994219
R42996 VDD.n7050 VDD.n2340 0.00994219
R42997 VDD.n7051 VDD.n2339 0.00994219
R42998 VDD.n7053 VDD.n2339 0.00994219
R42999 VDD.n7053 VDD.n2338 0.00994219
R43000 VDD.n7056 VDD.n2338 0.00994219
R43001 VDD.n7056 VDD.n2337 0.00994219
R43002 VDD.n7059 VDD.n2337 0.00994219
R43003 VDD.n7059 VDD.n2336 0.00994219
R43004 VDD.n7061 VDD.n2336 0.00994219
R43005 VDD.n7064 VDD.n7063 0.00994219
R43006 VDD.n7063 VDD.n2333 0.00994219
R43007 VDD.n7083 VDD.n7082 0.00994219
R43008 VDD.n7082 VDD.n2335 0.00994219
R43009 VDD.n7080 VDD.n2335 0.00994219
R43010 VDD.n7079 VDD.n7066 0.00994219
R43011 VDD.n7077 VDD.n7066 0.00994219
R43012 VDD.n7077 VDD.n7076 0.00994219
R43013 VDD.n7076 VDD.n7075 0.00994219
R43014 VDD.n7075 VDD.n7069 0.00994219
R43015 VDD.n7072 VDD.n7069 0.00994219
R43016 VDD.n7072 VDD.n7071 0.00994219
R43017 VDD.n7071 VDD.n2265 0.00994219
R43018 VDD.n10772 VDD.n10771 0.00983484
R43019 VDD.n2049 VDD.n2048 0.00983484
R43020 VDD.n10803 VDD.n10802 0.00983484
R43021 VDD.n10810 VDD.n1987 0.00983484
R43022 VDD.n1967 VDD.n1966 0.00983484
R43023 VDD.n10861 VDD.n10860 0.00983484
R43024 VDD.n10868 VDD.n1922 0.00983484
R43025 VDD.n5523 VDD.n5522 0.00983484
R43026 VDD.n10916 VDD.n10915 0.00983484
R43027 VDD.n10923 VDD.n1895 0.00983484
R43028 VDD.n1875 VDD.n1874 0.00983484
R43029 VDD.n10971 VDD.n10970 0.00983484
R43030 VDD.n10978 VDD.n1830 0.00983484
R43031 VDD.n1819 VDD.n1818 0.00983484
R43032 VDD.n11026 VDD.n11025 0.00983484
R43033 VDD.n9156 VDD.n9155 0.00983484
R43034 VDD.n9032 VDD.n9031 0.00983484
R43035 VDD.n9016 VDD.n9015 0.00983484
R43036 VDD.n8935 VDD.n8934 0.00983484
R43037 VDD.n8885 VDD.n8884 0.00983484
R43038 VDD.n8804 VDD.n8803 0.00983484
R43039 VDD.n8759 VDD.n8758 0.00983484
R43040 VDD.n9144 VDD.n9143 0.00983484
R43041 VDD.n8742 VDD.n8741 0.00983484
R43042 VDD.n8721 VDD.n8720 0.00983484
R43043 VDD.n8709 VDD.n8708 0.00983484
R43044 VDD.n8683 VDD.n8682 0.00983484
R43045 VDD.n8671 VDD.n8670 0.00983484
R43046 VDD.n8650 VDD.n8649 0.00983484
R43047 VDD.n12615 VDD.n12 0.00983484
R43048 VDD.n8130 VDD.n8128 0.00983194
R43049 VDD.n8127 VDD.n8125 0.00983194
R43050 VDD.n8124 VDD.n2020 0.00983194
R43051 VDD.n2027 VDD.n2023 0.00983194
R43052 VDD.n2031 VDD.n2028 0.00983194
R43053 VDD.n2035 VDD.n2032 0.00983194
R43054 VDD.n2101 VDD.n2099 0.00983194
R43055 VDD.n2098 VDD.n2096 0.00983194
R43056 VDD.n2095 VDD.n2010 0.00983194
R43057 VDD.n10788 VDD.n10787 0.00983194
R43058 VDD.n10792 VDD.n10789 0.00983194
R43059 VDD.n10796 VDD.n10793 0.00983194
R43060 VDD.n5593 VDD.n5591 0.00983194
R43061 VDD.n5590 VDD.n5588 0.00983194
R43062 VDD.n5587 VDD.n1947 0.00983194
R43063 VDD.n1972 VDD.n1950 0.00983194
R43064 VDD.n1976 VDD.n1973 0.00983194
R43065 VDD.n1980 VDD.n1977 0.00983194
R43066 VDD.n5614 VDD.n5612 0.00983194
R43067 VDD.n5611 VDD.n5609 0.00983194
R43068 VDD.n5608 VDD.n1937 0.00983194
R43069 VDD.n10846 VDD.n10845 0.00983194
R43070 VDD.n10850 VDD.n10847 0.00983194
R43071 VDD.n10854 VDD.n10851 0.00983194
R43072 VDD.n5899 VDD.n5897 0.00983194
R43073 VDD.n5896 VDD.n5894 0.00983194
R43074 VDD.n5893 VDD.n5892 0.00983194
R43075 VDD.n5494 VDD.n5493 0.00983194
R43076 VDD.n5498 VDD.n5495 0.00983194
R43077 VDD.n5502 VDD.n5499 0.00983194
R43078 VDD.n5677 VDD.n5675 0.00983194
R43079 VDD.n5674 VDD.n5672 0.00983194
R43080 VDD.n5671 VDD.n1910 0.00983194
R43081 VDD.n10901 VDD.n10900 0.00983194
R43082 VDD.n10905 VDD.n10902 0.00983194
R43083 VDD.n10909 VDD.n10906 0.00983194
R43084 VDD.n5690 VDD.n5688 0.00983194
R43085 VDD.n5687 VDD.n5685 0.00983194
R43086 VDD.n5684 VDD.n1855 0.00983194
R43087 VDD.n1880 VDD.n1858 0.00983194
R43088 VDD.n1884 VDD.n1881 0.00983194
R43089 VDD.n1888 VDD.n1885 0.00983194
R43090 VDD.n5797 VDD.n5795 0.00983194
R43091 VDD.n5794 VDD.n5792 0.00983194
R43092 VDD.n5791 VDD.n1845 0.00983194
R43093 VDD.n10956 VDD.n10955 0.00983194
R43094 VDD.n10960 VDD.n10957 0.00983194
R43095 VDD.n10964 VDD.n10961 0.00983194
R43096 VDD.n5742 VDD.n5740 0.00983194
R43097 VDD.n5739 VDD.n5737 0.00983194
R43098 VDD.n5736 VDD.n1790 0.00983194
R43099 VDD.n1797 VDD.n1793 0.00983194
R43100 VDD.n1801 VDD.n1798 0.00983194
R43101 VDD.n1805 VDD.n1802 0.00983194
R43102 VDD.n5716 VDD.n5714 0.00983194
R43103 VDD.n5713 VDD.n5711 0.00983194
R43104 VDD.n5710 VDD.n1783 0.00983194
R43105 VDD.n11011 VDD.n11010 0.00983194
R43106 VDD.n11015 VDD.n11012 0.00983194
R43107 VDD.n11019 VDD.n11016 0.00983194
R43108 VDD.n9062 VDD.n9060 0.00983194
R43109 VDD.n9059 VDD.n9057 0.00983194
R43110 VDD.n9056 VDD.n9055 0.00983194
R43111 VDD.n9052 VDD.n9050 0.00983194
R43112 VDD.n9049 VDD.n9048 0.00983194
R43113 VDD.n9046 VDD.n9045 0.00983194
R43114 VDD.n8928 VDD.n8926 0.00983194
R43115 VDD.n8925 VDD.n8923 0.00983194
R43116 VDD.n8922 VDD.n8921 0.00983194
R43117 VDD.n8918 VDD.n8916 0.00983194
R43118 VDD.n8915 VDD.n8914 0.00983194
R43119 VDD.n8912 VDD.n8505 0.00983194
R43120 VDD.n8849 VDD.n8516 0.00983194
R43121 VDD.n8853 VDD.n8852 0.00983194
R43122 VDD.n8857 VDD.n8854 0.00983194
R43123 VDD.n8862 VDD.n8861 0.00983194
R43124 VDD.n8866 VDD.n8863 0.00983194
R43125 VDD.n8870 VDD.n8867 0.00983194
R43126 VDD.n8579 VDD.n8577 0.00983194
R43127 VDD.n8576 VDD.n8574 0.00983194
R43128 VDD.n8573 VDD.n8572 0.00983194
R43129 VDD.n8569 VDD.n8567 0.00983194
R43130 VDD.n8566 VDD.n8565 0.00983194
R43131 VDD.n8563 VDD.n8562 0.00983194
R43132 VDD.n9083 VDD.n9081 0.00983194
R43133 VDD.n9080 VDD.n9078 0.00983194
R43134 VDD.n9077 VDD.n8465 0.00983194
R43135 VDD.n9176 VDD.n9174 0.00983194
R43136 VDD.n9173 VDD.n9172 0.00983194
R43137 VDD.n9170 VDD.n9169 0.00983194
R43138 VDD.n8591 VDD.n8589 0.00983194
R43139 VDD.n8588 VDD.n8586 0.00983194
R43140 VDD.n8585 VDD.n180 0.00983194
R43141 VDD.n12458 VDD.n12456 0.00983194
R43142 VDD.n12455 VDD.n12454 0.00983194
R43143 VDD.n12452 VDD.n12451 0.00983194
R43144 VDD.n8604 VDD.n8602 0.00983194
R43145 VDD.n8601 VDD.n8599 0.00983194
R43146 VDD.n8598 VDD.n109 0.00983194
R43147 VDD.n12478 VDD.n12477 0.00983194
R43148 VDD.n12482 VDD.n12479 0.00983194
R43149 VDD.n12486 VDD.n12483 0.00983194
R43150 VDD.n8696 VDD.n8694 0.00983194
R43151 VDD.n8693 VDD.n8691 0.00983194
R43152 VDD.n8690 VDD.n100 0.00983194
R43153 VDD.n12514 VDD.n12512 0.00983194
R43154 VDD.n12511 VDD.n12510 0.00983194
R43155 VDD.n12508 VDD.n12507 0.00983194
R43156 VDD.n8663 VDD.n8661 0.00983194
R43157 VDD.n8660 VDD.n8658 0.00983194
R43158 VDD.n8657 VDD.n29 0.00983194
R43159 VDD.n12534 VDD.n12533 0.00983194
R43160 VDD.n12538 VDD.n12535 0.00983194
R43161 VDD.n12542 VDD.n12539 0.00983194
R43162 VDD.n8632 VDD.n8630 0.00983194
R43163 VDD.n8629 VDD.n8627 0.00983194
R43164 VDD.n8626 VDD.n20 0.00983194
R43165 VDD.n12608 VDD.n12606 0.00983194
R43166 VDD.n12605 VDD.n12604 0.00983194
R43167 VDD.n12602 VDD.n12601 0.00983194
R43168 VDD.n2115 VDD.n2113 0.00974509
R43169 VDD.n2112 VDD.n1993 0.00974509
R43170 VDD.n10827 VDD.n10825 0.00974509
R43171 VDD.n10824 VDD.n10823 0.00974509
R43172 VDD.n5635 VDD.n5633 0.00974509
R43173 VDD.n5632 VDD.n5630 0.00974509
R43174 VDD.n5629 VDD.n1928 0.00974509
R43175 VDD.n10882 VDD.n10880 0.00974509
R43176 VDD.n10879 VDD.n10878 0.00974509
R43177 VDD.n10876 VDD.n10875 0.00974509
R43178 VDD.n5852 VDD.n5850 0.00974509
R43179 VDD.n5849 VDD.n5847 0.00974509
R43180 VDD.n5846 VDD.n1901 0.00974509
R43181 VDD.n10937 VDD.n10935 0.00974509
R43182 VDD.n10934 VDD.n10933 0.00974509
R43183 VDD.n10931 VDD.n10930 0.00974509
R43184 VDD.n5703 VDD.n5701 0.00974509
R43185 VDD.n5700 VDD.n5698 0.00974509
R43186 VDD.n5697 VDD.n1836 0.00974509
R43187 VDD.n10992 VDD.n10990 0.00974509
R43188 VDD.n10989 VDD.n10988 0.00974509
R43189 VDD.n10986 VDD.n10985 0.00974509
R43190 VDD.n8976 VDD.n8497 0.00974509
R43191 VDD.n8980 VDD.n8979 0.00974509
R43192 VDD.n8984 VDD.n8981 0.00974509
R43193 VDD.n8989 VDD.n8988 0.00974509
R43194 VDD.n8993 VDD.n8990 0.00974509
R43195 VDD.n8997 VDD.n8994 0.00974509
R43196 VDD.n8797 VDD.n8795 0.00974509
R43197 VDD.n8794 VDD.n8792 0.00974509
R43198 VDD.n8791 VDD.n8790 0.00974509
R43199 VDD.n8787 VDD.n8785 0.00974509
R43200 VDD.n8784 VDD.n8783 0.00974509
R43201 VDD.n8781 VDD.n8524 0.00974509
R43202 VDD.n8734 VDD.n8732 0.00974509
R43203 VDD.n8731 VDD.n8729 0.00974509
R43204 VDD.n8728 VDD.n119 0.00974509
R43205 VDD.n126 VDD.n122 0.00974509
R43206 VDD.n130 VDD.n127 0.00974509
R43207 VDD.n134 VDD.n131 0.00974509
R43208 VDD.n8618 VDD.n8616 0.00974509
R43209 VDD.n8615 VDD.n8613 0.00974509
R43210 VDD.n8612 VDD.n39 0.00974509
R43211 VDD.n80 VDD.n42 0.00974509
R43212 VDD.n84 VDD.n81 0.00974509
R43213 VDD.n88 VDD.n85 0.00974509
R43214 VDD.n6712 VDD.n6711 0.00970384
R43215 VDD.n6710 VDD.n6709 0.00970384
R43216 VDD.n6708 VDD.n6707 0.00970384
R43217 VDD.n6705 VDD.n6704 0.00970384
R43218 VDD.n6703 VDD.n6702 0.00970384
R43219 VDD.n6701 VDD.n6700 0.00970384
R43220 VDD.n6698 VDD.n6697 0.00970384
R43221 VDD.n6696 VDD.n6695 0.00970384
R43222 VDD.n6694 VDD.n6693 0.00970384
R43223 VDD.n6691 VDD.n6690 0.00970384
R43224 VDD.n6689 VDD.n6688 0.00970384
R43225 VDD.n6687 VDD.n6686 0.00970384
R43226 VDD.n6641 VDD.n6640 0.00970384
R43227 VDD.n6639 VDD.n6638 0.00970384
R43228 VDD.n6637 VDD.n6636 0.00970384
R43229 VDD.n5434 VDD.n5267 0.00970384
R43230 VDD.n5436 VDD.n5435 0.00970384
R43231 VDD.n5438 VDD.n5437 0.00970384
R43232 VDD.n5443 VDD.n5442 0.00970384
R43233 VDD.n5441 VDD.n5440 0.00970384
R43234 VDD.n5439 VDD.n5269 0.00970384
R43235 VDD.n6630 VDD.n6629 0.00970384
R43236 VDD.n6628 VDD.n6627 0.00970384
R43237 VDD.n6626 VDD.n6625 0.00970384
R43238 VDD.n950 VDD.n949 0.00969752
R43239 VDD.n970 VDD.n969 0.00964201
R43240 VDD.n972 VDD.n971 0.00964201
R43241 VDD.n974 VDD.n973 0.00964201
R43242 VDD.n976 VDD.n975 0.00964201
R43243 VDD.n988 VDD.n987 0.00964201
R43244 VDD.n990 VDD.n989 0.00964201
R43245 VDD.n992 VDD.n991 0.00964201
R43246 VDD.n994 VDD.n993 0.00964201
R43247 VDD.n1009 VDD.n1008 0.00964201
R43248 VDD.n1011 VDD.n1010 0.00964201
R43249 VDD.n1013 VDD.n1012 0.00964201
R43250 VDD.n1015 VDD.n1014 0.00964201
R43251 VDD.n1030 VDD.n1029 0.00964201
R43252 VDD.n1028 VDD.n1027 0.00964201
R43253 VDD.n1026 VDD.n1025 0.00964201
R43254 VDD.n1024 VDD.n1023 0.00964201
R43255 VDD.n1206 VDD.n1189 0.0095
R43256 VDD.n1176 VDD.n1118 0.0095
R43257 VDD.n1336 VDD.n1335 0.0095
R43258 VDD.n1383 VDD.n1382 0.0095
R43259 VDD.n1269 VDD.n1251 0.0095
R43260 VDD.n1236 VDD.n1219 0.0095
R43261 VDD.n1304 VDD.n1303 0.0095
R43262 VDD.n1072 VDD.n896 0.0095
R43263 VDD.n1059 VDD.n1058 0.0095
R43264 VDD.n1163 VDD.n1139 0.0095
R43265 VDD.n6287 VDD.n6286 0.00947673
R43266 VDD.n6279 VDD.n6278 0.00947673
R43267 VDD.n6251 VDD.n6250 0.00947673
R43268 VDD.n6243 VDD.n6242 0.00947673
R43269 VDD.n6675 VDD.n6674 0.00947673
R43270 VDD.n6667 VDD.n6666 0.00947673
R43271 VDD.n7064 VDD.n7061 0.00947673
R43272 VDD.n7080 VDD.n7079 0.00947673
R43273 VDD.n5892 VDD.n5890 0.00945616
R43274 VDD.n8017 VDD.n8016 0.00944828
R43275 VDD.n968 VDD.n682 0.00931657
R43276 VDD.n969 VDD.n968 0.00931657
R43277 VDD.n970 VDD.n967 0.00931657
R43278 VDD.n971 VDD.n967 0.00931657
R43279 VDD.n972 VDD.n966 0.00931657
R43280 VDD.n973 VDD.n966 0.00931657
R43281 VDD.n974 VDD.n965 0.00931657
R43282 VDD.n975 VDD.n965 0.00931657
R43283 VDD.n976 VDD.n964 0.00931657
R43284 VDD.n977 VDD.n964 0.00931657
R43285 VDD.n986 VDD.n963 0.00931657
R43286 VDD.n987 VDD.n963 0.00931657
R43287 VDD.n988 VDD.n962 0.00931657
R43288 VDD.n989 VDD.n962 0.00931657
R43289 VDD.n990 VDD.n961 0.00931657
R43290 VDD.n991 VDD.n961 0.00931657
R43291 VDD.n992 VDD.n960 0.00931657
R43292 VDD.n993 VDD.n960 0.00931657
R43293 VDD.n994 VDD.n959 0.00931657
R43294 VDD.n995 VDD.n959 0.00931657
R43295 VDD.n996 VDD.n958 0.00931657
R43296 VDD.n997 VDD.n958 0.00931657
R43297 VDD.n1005 VDD.n942 0.00931657
R43298 VDD.n1006 VDD.n942 0.00931657
R43299 VDD.n1007 VDD.n941 0.00931657
R43300 VDD.n1008 VDD.n941 0.00931657
R43301 VDD.n1009 VDD.n940 0.00931657
R43302 VDD.n1010 VDD.n940 0.00931657
R43303 VDD.n1011 VDD.n939 0.00931657
R43304 VDD.n1012 VDD.n939 0.00931657
R43305 VDD.n1013 VDD.n938 0.00931657
R43306 VDD.n1014 VDD.n938 0.00931657
R43307 VDD.n1015 VDD.n937 0.00931657
R43308 VDD.n1016 VDD.n937 0.00931657
R43309 VDD.n1031 VDD.n1017 0.00931657
R43310 VDD.n1030 VDD.n1017 0.00931657
R43311 VDD.n1029 VDD.n1018 0.00931657
R43312 VDD.n1028 VDD.n1018 0.00931657
R43313 VDD.n1027 VDD.n1019 0.00931657
R43314 VDD.n1026 VDD.n1019 0.00931657
R43315 VDD.n1025 VDD.n1020 0.00931657
R43316 VDD.n1024 VDD.n1020 0.00931657
R43317 VDD.n1023 VDD.n1021 0.00931657
R43318 VDD.n1022 VDD.n1021 0.00931657
R43319 VDD.n6267 VDD.n6266 0.00927724
R43320 VDD.n6266 VDD.n6262 0.00927724
R43321 VDD.n7048 VDD.n2342 0.00927724
R43322 VDD.n7049 VDD.n7048 0.00927724
R43323 VDD.n6284 VDD.n6283 0.00887828
R43324 VDD.n6248 VDD.n6247 0.00887828
R43325 VDD.n6672 VDD.n2350 0.00887828
R43326 VDD.n7084 VDD.n2333 0.00887828
R43327 VDD.n1450 VDD.n1449 0.00882321
R43328 VDD.n8014 VDD.n8013 0.00877586
R43329 VDD.n1612 VDD.n1610 0.00867241
R43330 VDD.n1480 VDD.n813 0.00867241
R43331 VDD.n5493 VDD.n1919 0.00864196
R43332 VDD.n1418 VDD.n852 0.00841379
R43333 VDD.n1678 VDD.n745 0.00841379
R43334 VDD.n1619 VDD.n1618 0.00841379
R43335 VDD.n1106 VDD.n1100 0.00841379
R43336 VDD.n1684 VDD.n742 0.00841379
R43337 VDD.n1698 VDD.n1697 0.00841379
R43338 VDD.n1045 VDD.n936 0.00841379
R43339 VDD.n1145 VDD.n706 0.00841379
R43340 VDD.n12583 VDD.n12577 0.0083892
R43341 VDD.n1426 VDD.n851 0.00836207
R43342 VDD.n1432 VDD.n1431 0.00836207
R43343 VDD.n1417 VDD.n873 0.00836207
R43344 VDD.n793 VDD.n744 0.00836207
R43345 VDD.n830 VDD.n738 0.00836207
R43346 VDD.n1371 VDD.n739 0.00836207
R43347 VDD.n1257 VDD.n783 0.00836207
R43348 VDD.n1352 VDD.n1085 0.00836207
R43349 VDD.n1467 VDD.n741 0.00836207
R43350 VDD.n885 VDD.n736 0.00836207
R43351 VDD.n1047 VDD.n1046 0.00836207
R43352 VDD.n1722 VDD.n1721 0.00836207
R43353 VDD.n1002 VDD.n997 0.00831065
R43354 VDD.n1637 VDD.n773 0.00808484
R43355 VDD.n1593 VDD.n1592 0.00806656
R43356 VDD.n6300 VDD.n6200 0.00801385
R43357 VDD.n1567 VDD.n1566 0.00800848
R43358 VDD.n697 VDD.n696 0.00797611
R43359 VDD.n7890 VDD.n7889 0.00791176
R43360 VDD.n7909 VDD.n7864 0.00787705
R43361 VDD.n8013 VDD.n8012 0.00763793
R43362 VDD.n1636 VDD.n774 0.0076267
R43363 VDD.n776 VDD.n775 0.0076267
R43364 VDD.n1635 VDD.n1634 0.0076267
R43365 VDD.n7983 VDD.n7982 0.0073513
R43366 VDD.n2196 VDD.n2195 0.0073513
R43367 VDD.n2191 VDD.n2190 0.0073513
R43368 VDD.n7989 VDD.n2192 0.0073513
R43369 VDD.n7988 VDD.n7987 0.0073513
R43370 VDD.n2221 VDD.n2220 0.0073513
R43371 VDD.n2224 VDD.n2223 0.0073513
R43372 VDD.n2231 VDD.n2212 0.0073513
R43373 VDD.n2214 VDD.n2213 0.0073513
R43374 VDD.n2228 VDD.n2227 0.0073513
R43375 VDD.n1542 VDD.n1535 0.00716667
R43376 VDD.n9134 VDD.n9132 0.00714138
R43377 VDD.n7986 VDD.n2193 0.00713029
R43378 VDD.n2219 VDD.n2218 0.00713029
R43379 VDD.n1529 VDD.n1523 0.00711202
R43380 VDD.n7980 VDD.n2197 0.0070075
R43381 VDD.n7979 VDD.n2194 0.0070075
R43382 VDD.n2217 VDD.n2216 0.0070075
R43383 VDD.n2215 VDD.n2207 0.0070075
R43384 VDD.n2038 VDD.n2007 0.0069938
R43385 VDD.n1956 VDD.n1934 0.0069938
R43386 VDD.n5512 VDD.n1907 0.0069938
R43387 VDD.n1864 VDD.n1842 0.0069938
R43388 VDD.n1808 VDD.n1780 0.0069938
R43389 VDD.n9064 VDD.n8475 0.0069938
R43390 VDD.n8891 VDD.n8513 0.0069938
R43391 VDD.n8748 VDD.n8582 0.0069938
R43392 VDD.n8698 VDD.n8607 0.0069938
R43393 VDD.n8639 VDD.n8623 0.0069938
R43394 VDD.n2160 VDD.n2159 0.00696552
R43395 VDD.n7962 VDD.n7961 0.00693383
R43396 VDD.n7965 VDD.n2202 0.00693383
R43397 VDD.n7968 VDD.n7966 0.00693383
R43398 VDD.n7967 VDD.n2200 0.00693383
R43399 VDD.n7970 VDD.n7969 0.00693383
R43400 VDD.n1206 VDD.n1205 0.00691379
R43401 VDD.n1176 VDD.n1134 0.00691379
R43402 VDD.n1336 VDD.n1319 0.00691379
R43403 VDD.n1383 VDD.n1365 0.00691379
R43404 VDD.n1269 VDD.n1268 0.00691379
R43405 VDD.n1236 VDD.n1235 0.00691379
R43406 VDD.n1304 VDD.n1287 0.00691379
R43407 VDD.n1072 VDD.n879 0.00691379
R43408 VDD.n1059 VDD.n917 0.00691379
R43409 VDD.n1163 VDD.n1156 0.00691379
R43410 VDD.n7175 VDD.n2297 0.00682401
R43411 VDD.n7827 VDD.n2240 0.00682401
R43412 VDD.n10821 VDD.n10820 0.00664271
R43413 VDD.n2043 VDD.n2038 0.00658794
R43414 VDD.n1961 VDD.n1956 0.00658794
R43415 VDD.n5517 VDD.n5512 0.00658794
R43416 VDD.n1869 VDD.n1864 0.00658794
R43417 VDD.n1813 VDD.n1808 0.00658794
R43418 VDD.n9069 VDD.n8475 0.00658794
R43419 VDD.n8896 VDD.n8513 0.00658794
R43420 VDD.n8753 VDD.n8582 0.00658794
R43421 VDD.n8703 VDD.n8607 0.00658794
R43422 VDD.n8644 VDD.n8623 0.00658794
R43423 VDD.n2233 VDD.n2211 0.00656548
R43424 VDD.n7993 VDD.n2189 0.00651637
R43425 VDD.n8017 VDD.n2165 0.0065
R43426 VDD.n2201 VDD.n2199 0.0064427
R43427 VDD.n10760 VDD.n10759 0.00633837
R43428 VDD.n1633 VDD.n777 0.00625226
R43429 VDD.n1519 VDD.n778 0.00625226
R43430 VDD.n1632 VDD.n1631 0.00625226
R43431 VDD.n8092 VDD.n2116 0.00617735
R43432 VDD.n12448 VDD.n195 0.00617182
R43433 VDD.n12445 VDD.n195 0.00617182
R43434 VDD.n12626 VDD.n12621 0.00599088
R43435 VDD.n1736 VDD.n696 0.00595628
R43436 VDD.n7975 VDD.n7973 0.00595157
R43437 VDD.n7974 VDD.n2198 0.00595157
R43438 VDD.n7977 VDD.n7976 0.00595157
R43439 VDD.n7850 VDD.n7849 0.00595157
R43440 VDD.n7851 VDD.n2206 0.00595157
R43441 VDD.n12630 VDD.n12625 0.00580154
R43442 VDD.n6320 VDD.n6319 0.00551189
R43443 VDD.n6319 VDD.n5914 0.00551189
R43444 VDD.n6177 VDD.n6016 0.00551189
R43445 VDD.n6179 VDD.n6016 0.00551189
R43446 VDD.n6174 VDD.n6173 0.00550912
R43447 VDD.n2159 VDD.n2158 0.00531034
R43448 VDD.n5768 VDD.n5763 0.00523684
R43449 VDD.n5759 VDD.n5758 0.00523684
R43450 VDD.n5835 VDD.n5830 0.00523684
R43451 VDD.n5826 VDD.n5825 0.00523684
R43452 VDD.n5652 VDD.n5647 0.00523684
R43453 VDD.n5643 VDD.n5642 0.00523684
R43454 VDD.n5570 VDD.n5565 0.00523684
R43455 VDD.n5561 VDD.n5560 0.00523684
R43456 VDD.n8156 VDD.n8151 0.00523684
R43457 VDD.n8147 VDD.n8146 0.00523684
R43458 VDD.n7997 VDD.n2186 0.00512451
R43459 VDD.n1442 VDD.n823 0.00510675
R43460 VDD.n1440 VDD.n823 0.00506157
R43461 VDD.n1756 VDD.n1752 0.00505621
R43462 VDD.n984 VDD.n977 0.00502663
R43463 VDD.n1033 VDD.n1016 0.00502663
R43464 VDD.n5980 VDD.n5979 0.00501642
R43465 VDD.n7305 VDD.n7302 0.00500851
R43466 VDD.n7305 VDD.n7304 0.00500851
R43467 VDD.n7304 VDD.n2088 0.00500851
R43468 VDD.n8168 VDD.n2086 0.00500851
R43469 VDD.n8172 VDD.n2086 0.00500851
R43470 VDD.n8175 VDD.n8174 0.00500851
R43471 VDD.n8175 VDD.n2084 0.00500851
R43472 VDD.n8179 VDD.n2084 0.00500851
R43473 VDD.n8180 VDD.n8179 0.00500851
R43474 VDD.n8183 VDD.n8180 0.00500851
R43475 VDD.n8187 VDD.n2082 0.00500851
R43476 VDD.n8190 VDD.n8189 0.00500851
R43477 VDD.n8190 VDD.n2080 0.00500851
R43478 VDD.n8194 VDD.n2080 0.00500851
R43479 VDD.n8195 VDD.n8194 0.00500851
R43480 VDD.n8196 VDD.n8195 0.00500851
R43481 VDD.n8200 VDD.n8199 0.00500851
R43482 VDD.n8203 VDD.n8200 0.00500851
R43483 VDD.n8207 VDD.n2076 0.00500851
R43484 VDD.n8208 VDD.n8207 0.00500851
R43485 VDD.n8209 VDD.n8208 0.00500851
R43486 VDD.n8213 VDD.n8212 0.00500851
R43487 VDD.n8216 VDD.n8213 0.00500851
R43488 VDD.n8220 VDD.n2072 0.00500851
R43489 VDD.n8221 VDD.n8220 0.00500851
R43490 VDD.n8223 VDD.n2070 0.00500851
R43491 VDD.n8227 VDD.n2070 0.00500851
R43492 VDD.n8228 VDD.n8227 0.00500851
R43493 VDD.n8230 VDD.n8228 0.00500851
R43494 VDD.n8234 VDD.n2068 0.00500851
R43495 VDD.n8235 VDD.n8234 0.00500851
R43496 VDD.n8238 VDD.n2066 0.00500851
R43497 VDD.n8242 VDD.n2066 0.00500851
R43498 VDD.n8243 VDD.n8242 0.00500851
R43499 VDD.n8244 VDD.n8243 0.00500851
R43500 VDD.n8248 VDD.n8247 0.00500851
R43501 VDD.n8251 VDD.n8248 0.00500851
R43502 VDD.n10765 VDD.n2062 0.00500851
R43503 VDD.n10761 VDD.n2062 0.00500851
R43504 VDD.n10761 VDD.n10760 0.00500851
R43505 VDD.n986 VDD.n985 0.00499704
R43506 VDD.n1032 VDD.n1031 0.00499704
R43507 VDD.n1564 VDD.n1510 0.00497964
R43508 VDD.n7960 VDD.n2203 0.00489563
R43509 VDD.n1630 VDD.n779 0.00487783
R43510 VDD.n781 VDD.n780 0.00487783
R43511 VDD.n1629 VDD.n1628 0.00487783
R43512 VDD.n1592 VDD.n1504 0.00487179
R43513 VDD.n2157 VDD.n2156 0.00484483
R43514 VDD.n8141 VDD.n8140 0.00483155
R43515 VDD.n5554 VDD.n5553 0.00483155
R43516 VDD.n5545 VDD.n5544 0.00483155
R43517 VDD.n5820 VDD.n5819 0.00483155
R43518 VDD.n5753 VDD.n5752 0.00483155
R43519 VDD.n8970 VDD.n8953 0.00483155
R43520 VDD.n8830 VDD.n8812 0.00483155
R43521 VDD.n9117 VDD.n9099 0.00483155
R43522 VDD.n162 VDD.n144 0.00483155
R43523 VDD.n73 VDD.n55 0.00483155
R43524 VDD.n8244 VDD.n2064 0.00479584
R43525 VDD.n8212 VDD.n2074 0.00475331
R43526 VDD.n8182 VDD.n2082 0.00462571
R43527 VDD.n8202 VDD.n2076 0.00462571
R43528 VDD.n8188 VDD.n8187 0.00454064
R43529 VDD.n770 VDD.n769 0.00452149
R43530 VDD.n12640 VDD.n12639 0.00449408
R43531 VDD.n12581 VDD.n12558 0.00447616
R43532 VDD.n12582 VDD.n12581 0.00446857
R43533 VDD.n12583 VDD.n12582 0.00446857
R43534 VDD VDD.n0 0.0044645
R43535 VDD.n8223 VDD.n8222 0.00445558
R43536 VDD.n6323 VDD.n5980 0.00444161
R43537 VDD.n5288 VDD.n5287 0.00441304
R43538 VDD.n6413 VDD.n5298 0.00441304
R43539 VDD.n6876 VDD.n2385 0.00441304
R43540 VDD.n2375 VDD.n2374 0.00441304
R43541 VDD.n1628 VDD.n1627 0.00436878
R43542 VDD.n1639 VDD.n1638 0.00434333
R43543 VDD.n773 VDD.n772 0.00434333
R43544 VDD.n1626 VDD.n782 0.00431787
R43545 VDD.n6575 VDD.n6574 0.00429447
R43546 VDD.n6399 VDD.n6398 0.00429447
R43547 VDD.n6862 VDD.n6861 0.00429447
R43548 VDD.n7038 VDD.n7037 0.00429447
R43549 VDD.n1638 VDD.n772 0.00424152
R43550 VDD.n6580 VDD.n6579 0.00418286
R43551 VDD.n5965 VDD.n5964 0.00418286
R43552 VDD.n6610 VDD.n6609 0.00418286
R43553 VDD.n12639 VDD.n0 0.00416864
R43554 VDD.n1641 VDD.n770 0.00406335
R43555 VDD.n60 VDD.n59 0.00405263
R43556 VDD.n69 VDD.n68 0.00405263
R43557 VDD.n149 VDD.n148 0.00405263
R43558 VDD.n158 VDD.n157 0.00405263
R43559 VDD.n9104 VDD.n9103 0.00405263
R43560 VDD.n9113 VDD.n9112 0.00405263
R43561 VDD.n8817 VDD.n8816 0.00405263
R43562 VDD.n8826 VDD.n8825 0.00405263
R43563 VDD.n8957 VDD.n8956 0.00405263
R43564 VDD.n8966 VDD.n8965 0.00405263
R43565 VDD.n6175 VDD.n6174 0.00403102
R43566 VDD.n10766 VDD.n2061 0.00403025
R43567 VDD.n1631 VDD.n1630 0.00398699
R43568 VDD.n8251 VDD.n8250 0.00394518
R43569 VDD.n2054 VDD.n2035 0.00388205
R43570 VDD.n10797 VDD.n10796 0.00388205
R43571 VDD.n1981 VDD.n1980 0.00388205
R43572 VDD.n10855 VDD.n10854 0.00388205
R43573 VDD.n10910 VDD.n10909 0.00388205
R43574 VDD.n1889 VDD.n1888 0.00388205
R43575 VDD.n10965 VDD.n10964 0.00388205
R43576 VDD.n1824 VDD.n1805 0.00388205
R43577 VDD.n11020 VDD.n11019 0.00388205
R43578 VDD.n9063 VDD.n9062 0.00385073
R43579 VDD.n8929 VDD.n8928 0.00385073
R43580 VDD.n8890 VDD.n8516 0.00385073
R43581 VDD.n8764 VDD.n8579 0.00385073
R43582 VDD.n9150 VDD.n9083 0.00385073
R43583 VDD.n8747 VDD.n8591 0.00385073
R43584 VDD.n8714 VDD.n8604 0.00385073
R43585 VDD.n8697 VDD.n8696 0.00385073
R43586 VDD.n8664 VDD.n8663 0.00385073
R43587 VDD.n8638 VDD.n8632 0.00385073
R43588 VDD.n10875 VDD.n10873 0.00385057
R43589 VDD.n10930 VDD.n10928 0.00385057
R43590 VDD.n10985 VDD.n10983 0.00385057
R43591 VDD.n9021 VDD.n8497 0.00381954
R43592 VDD.n8798 VDD.n8797 0.00381954
R43593 VDD.n8735 VDD.n8734 0.00381954
R43594 VDD.n8676 VDD.n8618 0.00381954
R43595 VDD.n10148 VDD.n9184 0.00378966
R43596 VDD.n10148 VDD.n9185 0.00378966
R43597 VDD.n8199 VDD.n2078 0.00377505
R43598 VDD.n11136 VDD.n11135 0.00372459
R43599 VDD.n6190 VDD.n5988 0.0037107
R43600 VDD.n6328 VDD.n5487 0.00371011
R43601 VDD.n780 VDD.n779 0.00370701
R43602 VDD.n1629 VDD.n781 0.00370701
R43603 VDD.n949 VDD.n948 0.00364636
R43604 VDD.n8215 VDD.n2072 0.00360491
R43605 VDD.n8238 VDD.n8237 0.00360491
R43606 VDD.n10820 VDD.n2000 0.00360238
R43607 VDD.n1640 VDD.n1639 0.00357975
R43608 VDD.n8064 VDD.n2147 0.00355172
R43609 VDD.n10815 VDD.n2004 0.00354033
R43610 VDD.n1565 VDD.n1564 0.00352885
R43611 VDD.n1449 VDD.n821 0.00352662
R43612 VDD.n7853 VDD.n7852 0.00342224
R43613 VDD.n5950 VDD.n5949 0.00334483
R43614 VDD.n10890 VDD.n1919 0.0031618
R43615 VDD.n7853 VDD.n2205 0.00302933
R43616 VDD.n8174 VDD.n8173 0.00300945
R43617 VDD.n12586 VDD.n12558 0.00289832
R43618 VDD.n8012 VDD.n8011 0.00277586
R43619 VDD.n8230 VDD.n8229 0.00275425
R43620 VDD.n8229 VDD.n2068 0.00275425
R43621 VDD.n680 VDD.n679 0.00274852
R43622 VDD.n5362 VDD.n5299 0.00272414
R43623 VDD.n2402 VDD.n2401 0.00272414
R43624 VDD.n5902 VDD.n5541 0.00272168
R43625 VDD.n5905 VDD.n5901 0.00272168
R43626 VDD.n5889 VDD.n1918 0.00272168
R43627 VDD.n5534 VDD.n5490 0.00272168
R43628 VDD.n5907 VDD.n5541 0.00272168
R43629 VDD.n5905 VDD.n5902 0.00272168
R43630 VDD.n5529 VDD.n5490 0.00272168
R43631 VDD.n5890 VDD.n5889 0.00272168
R43632 VDD.n8092 VDD.n2108 0.00270566
R43633 VDD.n8095 VDD.n2108 0.00270566
R43634 VDD.n1447 VDD.n821 0.00268589
R43635 VDD.n8068 VDD.n8067 0.00267241
R43636 VDD.n5529 VDD.n5528 0.00266075
R43637 VDD.n5220 VDD.n2411 0.00263633
R43638 VDD.n5218 VDD.n2411 0.00263633
R43639 VDD.n1548 VDD.n1547 0.00263115
R43640 VDD.n1756 VDD.n681 0.00262663
R43641 VDD.n998 VDD.n956 0.00262663
R43642 VDD.n12640 VDD.n2 0.00262663
R43643 VDD.n681 VDD.n678 0.00262663
R43644 VDD.n1002 VDD.n998 0.00262663
R43645 VDD.n12642 VDD.n2 0.00262663
R43646 VDD.n1634 VDD.n1633 0.00261256
R43647 VDD.n5503 VDD.n5502 0.00259812
R43648 VDD.n8098 VDD.n2105 0.00257859
R43649 VDD.n6300 VDD.n6299 0.00254425
R43650 VDD.n7963 VDD.n7960 0.0025382
R43651 VDD.n8173 VDD.n8172 0.00249905
R43652 VDD.n5249 VDD.n5248 0.00237378
R43653 VDD.n5459 VDD.n5458 0.00237378
R43654 VDD.n5348 VDD.n5347 0.00237378
R43655 VDD.n6394 VDD.n6393 0.00237378
R43656 VDD.n5481 VDD.n5479 0.00237378
R43657 VDD.n2305 VDD.n2303 0.00237378
R43658 VDD.n5420 VDD.n5419 0.00237378
R43659 VDD.n7110 VDD.n7109 0.00237378
R43660 VDD.n956 VDD.n952 0.00236391
R43661 VDD.n8011 VDD.n2121 0.00236207
R43662 VDD.n7820 VDD.n2243 0.00235027
R43663 VDD.n7816 VDD.n2243 0.00235027
R43664 VDD.n7816 VDD.n7815 0.00235027
R43665 VDD.n7815 VDD.n7814 0.00235027
R43666 VDD.n7814 VDD.n2246 0.00235027
R43667 VDD.n7810 VDD.n2246 0.00235027
R43668 VDD.n7808 VDD.n7807 0.00235027
R43669 VDD.n7807 VDD.n2248 0.00235027
R43670 VDD.n7803 VDD.n2248 0.00235027
R43671 VDD.n7803 VDD.n7802 0.00235027
R43672 VDD.n7802 VDD.n7801 0.00235027
R43673 VDD.n7798 VDD.n7797 0.00235027
R43674 VDD.n7797 VDD.n7796 0.00235027
R43675 VDD.n7793 VDD.n7792 0.00235027
R43676 VDD.n7792 VDD.n7791 0.00235027
R43677 VDD.n7791 VDD.n2254 0.00235027
R43678 VDD.n7787 VDD.n2254 0.00235027
R43679 VDD.n7787 VDD.n7786 0.00235027
R43680 VDD.n7786 VDD.n7785 0.00235027
R43681 VDD.n7785 VDD.n2256 0.00235027
R43682 VDD.n7781 VDD.n2256 0.00235027
R43683 VDD.n7779 VDD.n7778 0.00235027
R43684 VDD.n7778 VDD.n2258 0.00235027
R43685 VDD.n7774 VDD.n7773 0.00235027
R43686 VDD.n7773 VDD.n7772 0.00235027
R43687 VDD.n7772 VDD.n2261 0.00235027
R43688 VDD.n7768 VDD.n2261 0.00235027
R43689 VDD.n7768 VDD.n7767 0.00235027
R43690 VDD.n7767 VDD.n7766 0.00235027
R43691 VDD.n7766 VDD.n2263 0.00235027
R43692 VDD.n7762 VDD.n2263 0.00235027
R43693 VDD.n7762 VDD.n7761 0.00235027
R43694 VDD.n7759 VDD.n2266 0.00235027
R43695 VDD.n7755 VDD.n2266 0.00235027
R43696 VDD.n7755 VDD.n7754 0.00235027
R43697 VDD.n7754 VDD.n7753 0.00235027
R43698 VDD.n7753 VDD.n2268 0.00235027
R43699 VDD.n7749 VDD.n2268 0.00235027
R43700 VDD.n7749 VDD.n7748 0.00235027
R43701 VDD.n7748 VDD.n7747 0.00235027
R43702 VDD.n7744 VDD.n7743 0.00235027
R43703 VDD.n7743 VDD.n7742 0.00235027
R43704 VDD.n7739 VDD.n7738 0.00235027
R43705 VDD.n7738 VDD.n7737 0.00235027
R43706 VDD.n7737 VDD.n2274 0.00235027
R43707 VDD.n7733 VDD.n2274 0.00235027
R43708 VDD.n7733 VDD.n7732 0.00235027
R43709 VDD.n7732 VDD.n7731 0.00235027
R43710 VDD.n7731 VDD.n2276 0.00235027
R43711 VDD.n7727 VDD.n2276 0.00235027
R43712 VDD.n7727 VDD.n7726 0.00235027
R43713 VDD.n7724 VDD.n2278 0.00235027
R43714 VDD.n7720 VDD.n2278 0.00235027
R43715 VDD.n7718 VDD.n7717 0.00235027
R43716 VDD.n7717 VDD.n2280 0.00235027
R43717 VDD.n7713 VDD.n7712 0.00235027
R43718 VDD.n7712 VDD.n7711 0.00235027
R43719 VDD.n7708 VDD.n7707 0.00235027
R43720 VDD.n7707 VDD.n7706 0.00235027
R43721 VDD.n7706 VDD.n2285 0.00235027
R43722 VDD.n7702 VDD.n2285 0.00235027
R43723 VDD.n7702 VDD.n7701 0.00235027
R43724 VDD.n7699 VDD.n2287 0.00235027
R43725 VDD.n7695 VDD.n2287 0.00235027
R43726 VDD.n7695 VDD.n7694 0.00235027
R43727 VDD.n7694 VDD.n7693 0.00235027
R43728 VDD.n7693 VDD.n2289 0.00235027
R43729 VDD.n7689 VDD.n7688 0.00235027
R43730 VDD.n7688 VDD.n7687 0.00235027
R43731 VDD.n7747 VDD.n2270 0.00233282
R43732 VDD.n1632 VDD.n778 0.00233258
R43733 VDD.n7781 VDD.n7780 0.00231536
R43734 VDD.n2969 VDD.n2966 0.00229222
R43735 VDD.n2966 VDD.n1768 0.00229222
R43736 VDD.n11038 VDD.n1768 0.00229222
R43737 VDD.n11050 VDD.n11049 0.00229222
R43738 VDD.n11050 VDD.n667 0.00229222
R43739 VDD.n11054 VDD.n667 0.00229222
R43740 VDD.n11055 VDD.n11054 0.00229222
R43741 VDD.n11058 VDD.n11055 0.00229222
R43742 VDD.n11062 VDD.n665 0.00229222
R43743 VDD.n11065 VDD.n11064 0.00229222
R43744 VDD.n11065 VDD.n663 0.00229222
R43745 VDD.n11069 VDD.n663 0.00229222
R43746 VDD.n11070 VDD.n11069 0.00229222
R43747 VDD.n11071 VDD.n11070 0.00229222
R43748 VDD.n11075 VDD.n11074 0.00229222
R43749 VDD.n11078 VDD.n11075 0.00229222
R43750 VDD.n11082 VDD.n659 0.00229222
R43751 VDD.n11083 VDD.n11082 0.00229222
R43752 VDD.n11084 VDD.n11083 0.00229222
R43753 VDD.n11088 VDD.n11087 0.00229222
R43754 VDD.n11091 VDD.n11088 0.00229222
R43755 VDD.n11095 VDD.n655 0.00229222
R43756 VDD.n11096 VDD.n11095 0.00229222
R43757 VDD.n11098 VDD.n653 0.00229222
R43758 VDD.n11102 VDD.n653 0.00229222
R43759 VDD.n11103 VDD.n11102 0.00229222
R43760 VDD.n11104 VDD.n11103 0.00229222
R43761 VDD.n11108 VDD.n11107 0.00229222
R43762 VDD.n11109 VDD.n11108 0.00229222
R43763 VDD.n11113 VDD.n11112 0.00229222
R43764 VDD.n11114 VDD.n11113 0.00229222
R43765 VDD.n11114 VDD.n646 0.00229222
R43766 VDD.n11118 VDD.n646 0.00229222
R43767 VDD.n11121 VDD.n11120 0.00229222
R43768 VDD.n11131 VDD.n631 0.00229222
R43769 VDD.n11135 VDD.n631 0.00229222
R43770 VDD.n11131 VDD.n11130 0.00225841
R43771 VDD.n11119 VDD.n11118 0.00220768
R43772 VDD.n6625 VDD.n6624 0.0021987
R43773 VDD.n11087 VDD.n657 0.00219078
R43774 VDD.n11121 VDD.n640 0.00219078
R43775 VDD.n12643 VDD.n1 0.00218639
R43776 VDD.n8168 VDD.n8167 0.00215879
R43777 VDD.n7719 VDD.n7718 0.00215826
R43778 VDD.n12625 VDD.n9 0.00214095
R43779 VDD.n11057 VDD.n665 0.00214005
R43780 VDD.n11077 VDD.n659 0.00214005
R43781 VDD.n8167 VDD.n8165 0.00211626
R43782 VDD.n11063 VDD.n11062 0.00210624
R43783 VDD.n7966 VDD.n7965 0.00209618
R43784 VDD.n11098 VDD.n11097 0.00207242
R43785 VDD.n12643 VDD.n12642 0.00206805
R43786 VDD.n7975 VDD.n7974 0.00202251
R43787 VDD.n7977 VDD.n2198 0.00202251
R43788 VDD.n7976 VDD.n2197 0.00202251
R43789 VDD.n7850 VDD.n2207 0.00202251
R43790 VDD.n7849 VDD.n2205 0.00202251
R43791 VDD.n7852 VDD.n7851 0.00202251
R43792 VDD.n7809 VDD.n7808 0.00200116
R43793 VDD.n7742 VDD.n2272 0.00198371
R43794 VDD.n5901 VDD.n5900 0.00197182
R43795 VDD.n2260 VDD.n2258 0.00196625
R43796 VDD.n12630 VDD.n12621 0.00195161
R43797 VDD.n2282 VDD.n2280 0.0019488
R43798 VDD.n7700 VDD.n7699 0.00193134
R43799 VDD.n12579 VDD.n12561 0.00192857
R43800 VDD.n638 VDD.n634 0.00192857
R43801 VDD.n1764 VDD.n1763 0.00192857
R43802 VDD.n6325 VDD.n5913 0.00192857
R43803 VDD.n6015 VDD.n6014 0.00192857
R43804 VDD.n5538 VDD.n5489 0.00192857
R43805 VDD.n5888 VDD.n5886 0.00192857
R43806 VDD.n5911 VDD.n5540 0.00192857
R43807 VDD.n8088 VDD.n2002 0.00192857
R43808 VDD.n8091 VDD.n8090 0.00192857
R43809 VDD.n12632 VDD.n8 0.00192857
R43810 VDD.n12636 VDD.n12635 0.00192857
R43811 VDD.n1001 VDD.n1000 0.00192857
R43812 VDD.n1760 VDD.n677 0.00192857
R43813 VDD.n1751 VDD.n680 0.00192012
R43814 VDD.n8216 VDD.n8215 0.00190359
R43815 VDD.n8237 VDD.n8235 0.00190359
R43816 VDD.n11126 VDD.n644 0.00190334
R43817 VDD.n8068 VDD.n2146 0.00189655
R43818 VDD.n1004 VDD.n952 0.00189053
R43819 VDD.n1183 VDD.n1182 0.00186957
R43820 VDD.n1170 VDD.n1169 0.00186957
R43821 VDD.n1654 VDD.n757 0.00186957
R43822 VDD.n1342 VDD.n1278 0.00186957
R43823 VDD.n1359 VDD.n1358 0.00186957
R43824 VDD.n1389 VDD.n876 0.00186957
R43825 VDD.n1650 VDD.n765 0.00186957
R43826 VDD.n1275 VDD.n1107 0.00186957
R43827 VDD.n1213 VDD.n1212 0.00186957
R43828 VDD.n1066 VDD.n1065 0.00186957
R43829 VDD.n911 VDD.n910 0.00186957
R43830 VDD.n1745 VDD.n1744 0.00186957
R43831 VDD.n11123 VDD.n642 0.00186953
R43832 VDD.n7725 VDD.n7724 0.00180915
R43833 VDD.n2291 VDD.n2289 0.00180915
R43834 VDD.n11074 VDD.n661 0.0018019
R43835 VDD.n5528 VDD.n5503 0.00178392
R43836 VDD.n7801 VDD.n2250 0.00175679
R43837 VDD.n11090 VDD.n655 0.00173427
R43838 VDD.n11112 VDD.n649 0.00173427
R43839 VDD.n8165 VDD.n2088 0.00173346
R43840 VDD.n8196 VDD.n2078 0.00173346
R43841 VDD.n8131 VDD.n8130 0.00168998
R43842 VDD.n8110 VDD.n2101 0.00168998
R43843 VDD.n5594 VDD.n5593 0.00168998
R43844 VDD.n5615 VDD.n5614 0.00168998
R43845 VDD.n5900 VDD.n5899 0.00168998
R43846 VDD.n5865 VDD.n5677 0.00168998
R43847 VDD.n5810 VDD.n5690 0.00168998
R43848 VDD.n5798 VDD.n5797 0.00168998
R43849 VDD.n5743 VDD.n5742 0.00168998
R43850 VDD.n5722 VDD.n5716 0.00168998
R43851 VDD.n9045 VDD.n9043 0.00168998
R43852 VDD.n8946 VDD.n8505 0.00168998
R43853 VDD.n8871 VDD.n8870 0.00168998
R43854 VDD.n8562 VDD.n8560 0.00168998
R43855 VDD.n9169 VDD.n9167 0.00168998
R43856 VDD.n12451 VDD.n12449 0.00168998
R43857 VDD.n12487 VDD.n12486 0.00168998
R43858 VDD.n12507 VDD.n12505 0.00168998
R43859 VDD.n12543 VDD.n12542 0.00168998
R43860 VDD.n12601 VDD.n12599 0.00168998
R43861 VDD.n2164 VDD.n2163 0.00168966
R43862 VDD.n6744 VDD.n6741 0.00168421
R43863 VDD.n6753 VDD.n6751 0.00168421
R43864 VDD.n6756 VDD.n6748 0.00168421
R43865 VDD.n6997 VDD.n6996 0.00168421
R43866 VDD.n6992 VDD.n6991 0.00168421
R43867 VDD.n6987 VDD.n6986 0.00168421
R43868 VDD.n6982 VDD.n6981 0.00168421
R43869 VDD.n6900 VDD.n6899 0.00168421
R43870 VDD.n6895 VDD.n6894 0.00168421
R43871 VDD.n6890 VDD.n6889 0.00168421
R43872 VDD.n6949 VDD.n6948 0.00168421
R43873 VDD.n6944 VDD.n6943 0.00168421
R43874 VDD.n6939 VDD.n6938 0.00168421
R43875 VDD.n6934 VDD.n6933 0.00168421
R43876 VDD.n6919 VDD.n6918 0.00168421
R43877 VDD.n6914 VDD.n6913 0.00168421
R43878 VDD.n6909 VDD.n6908 0.00168421
R43879 VDD.n6524 VDD.n6446 0.00168421
R43880 VDD.n6527 VDD.n6443 0.00168421
R43881 VDD.n6530 VDD.n6440 0.00168421
R43882 VDD.n6533 VDD.n6437 0.00168421
R43883 VDD.n6433 VDD.n6432 0.00168421
R43884 VDD.n6428 VDD.n6427 0.00168421
R43885 VDD.n6423 VDD.n6422 0.00168421
R43886 VDD.n6484 VDD.n6483 0.00168421
R43887 VDD.n6487 VDD.n6480 0.00168421
R43888 VDD.n6490 VDD.n6477 0.00168421
R43889 VDD.n6493 VDD.n6474 0.00168421
R43890 VDD.n6470 VDD.n6469 0.00168421
R43891 VDD.n6465 VDD.n6464 0.00168421
R43892 VDD.n6460 VDD.n6459 0.00168421
R43893 VDD.n6071 VDD.n6068 0.00168421
R43894 VDD.n6065 VDD.n6064 0.00168421
R43895 VDD.n6060 VDD.n6059 0.00168421
R43896 VDD.n6114 VDD.n6111 0.00168421
R43897 VDD.n6108 VDD.n6107 0.00168421
R43898 VDD.n6103 VDD.n6102 0.00168421
R43899 VDD.n7940 VDD.n7939 0.00168421
R43900 VDD.n7935 VDD.n7934 0.00168421
R43901 VDD.n7930 VDD.n7929 0.00168421
R43902 VDD.n7925 VDD.n7924 0.00168421
R43903 VDD.n7921 VDD.n7920 0.00168421
R43904 VDD.n7916 VDD.n7915 0.00168421
R43905 VDD.n7892 VDD.n7885 0.00168421
R43906 VDD.n7895 VDD.n7881 0.00168421
R43907 VDD.n7898 VDD.n7877 0.00168421
R43908 VDD.n7901 VDD.n7874 0.00168421
R43909 VDD.n7904 VDD.n7871 0.00168421
R43910 VDD.n7907 VDD.n7867 0.00168421
R43911 VDD.n8045 VDD.n8044 0.00168421
R43912 VDD.n8040 VDD.n8039 0.00168421
R43913 VDD.n8035 VDD.n8034 0.00168421
R43914 VDD.n8030 VDD.n8029 0.00168421
R43915 VDD.n8026 VDD.n8025 0.00168421
R43916 VDD.n8021 VDD.n8020 0.00168421
R43917 VDD.n6738 VDD.n6735 0.00168421
R43918 VDD.n6802 VDD.n6733 0.00168421
R43919 VDD.n6805 VDD.n6730 0.00168421
R43920 VDD.n6329 VDD.n6328 0.00168023
R43921 VDD.n6008 VDD.n5988 0.00167963
R43922 VDD.n8098 VDD.n8097 0.0016789
R43923 VDD.n5636 VDD.n5635 0.0016789
R43924 VDD.n5853 VDD.n5852 0.0016789
R43925 VDD.n5777 VDD.n5703 0.0016789
R43926 VDD.n8998 VDD.n8997 0.0016789
R43927 VDD.n8837 VDD.n8524 0.0016789
R43928 VDD.n169 VDD.n134 0.0016789
R43929 VDD.n89 VDD.n88 0.0016789
R43930 VDD.n7760 VDD.n7759 0.00161715
R43931 VDD.n7711 VDD.n2283 0.00159969
R43932 VDD.n6283 VDD.n6282 0.00156391
R43933 VDD.n6247 VDD.n6246 0.00156391
R43934 VDD.n6648 VDD.n2350 0.00156391
R43935 VDD.n7084 VDD.n7083 0.00156391
R43936 VDD.n8250 VDD.n2061 0.00156333
R43937 VDD.n2162 VDD.n2161 0.00153448
R43938 VDD.n7973 VDD.n2199 0.00153138
R43939 VDD.n11044 VDD.n673 0.00153137
R43940 VDD.n679 VDD.n678 0.00150592
R43941 VDD.n1520 VDD.n1519 0.00149265
R43942 VDD.n10766 VDD.n10765 0.00147826
R43943 VDD.n11046 VDD.n676 0.00146374
R43944 VDD.n7687 VDD.n2292 0.00146005
R43945 VDD.n7793 VDD.n2252 0.00144259
R43946 VDD.n1641 VDD.n1640 0.00144174
R43947 VDD.n7796 VDD.n2252 0.00140768
R43948 VDD.n11049 VDD.n11048 0.00139611
R43949 VDD.n11104 VDD.n651 0.00139611
R43950 VDD.n11107 VDD.n651 0.00139611
R43951 VDD.n7684 VDD.n2292 0.00139023
R43952 VDD.n6299 VDD.n6298 0.00138218
R43953 VDD.n1520 VDD.n777 0.00133993
R43954 VDD.n7993 VDD.n7992 0.00133493
R43955 VDD.n11046 VDD.n673 0.00132848
R43956 VDD.n676 VDD.n669 0.00129466
R43957 VDD.n2233 VDD.n2232 0.00128581
R43958 VDD.n10890 VDD.n1918 0.00128288
R43959 VDD.n11044 VDD.n11043 0.00126085
R43960 VDD.n7708 VDD.n2283 0.00125058
R43961 VDD.n1637 VDD.n1636 0.00123812
R43962 VDD.n7822 VDD.n7821 0.00123313
R43963 VDD.n7761 VDD.n7760 0.00123313
R43964 VDD.n11043 VDD.n1766 0.0011594
R43965 VDD.n11037 VDD.n1766 0.0011425
R43966 VDD.n7798 VDD.n2250 0.00109348
R43967 VDD.n1601 VDD.n1600 0.00108851
R43968 VDD.n1412 VDD.n1391 0.00108851
R43969 VDD.n820 VDD.n818 0.00108851
R43970 VDD.n810 VDD.n808 0.00108851
R43971 VDD.n1740 VDD.n693 0.00108851
R43972 VDD.n1716 VDD.n713 0.00108851
R43973 VDD.n5979 VDD.n5914 0.00107482
R43974 VDD.n8066 VDD.n8065 0.00106897
R43975 VDD.n12586 VDD.n12585 0.00106802
R43976 VDD.n11091 VDD.n11090 0.00105796
R43977 VDD.n11109 VDD.n649 0.00105796
R43978 VDD.n8222 VDD.n8221 0.00105293
R43979 VDD.n7821 VDD.n7820 0.00104112
R43980 VDD.n7726 VDD.n7725 0.00104112
R43981 VDD.n7689 VDD.n2291 0.00104112
R43982 VDD.n6599 VDD.n2203 0.00104025
R43983 VDD.n7963 VDD.n7962 0.00104025
R43984 VDD.n7961 VDD.n2202 0.00104025
R43985 VDD.n7968 VDD.n7967 0.00104025
R43986 VDD.n7970 VDD.n2200 0.00104025
R43987 VDD.n7969 VDD.n2201 0.00104025
R43988 VDD.n7684 VDD.n7683 0.00102366
R43989 VDD.n6177 VDD.n6175 0.000992701
R43990 VDD.n11038 VDD.n11037 0.000990325
R43991 VDD.n11071 VDD.n661 0.000990325
R43992 VDD.n8189 VDD.n8188 0.000967864
R43993 VDD.n7980 VDD.n7979 0.000966576
R43994 VDD.n2216 VDD.n2215 0.000966576
R43995 VDD.n775 VDD.n774 0.000958145
R43996 VDD.n1635 VDD.n776 0.000958145
R43997 VDD.n1672 VDD.n747 0.000923032
R43998 VDD.n7701 VDD.n7700 0.000918929
R43999 VDD.n7713 VDD.n2282 0.000901474
R44000 VDD.n1558 VDD.n1512 0.000893443
R44001 VDD.n1554 VDD.n1553 0.000893443
R44002 VDD.n11127 VDD.n642 0.000888878
R44003 VDD.n644 VDD.n633 0.000888878
R44004 VDD.n7774 VDD.n2260 0.000884019
R44005 VDD.n8183 VDD.n8182 0.000882798
R44006 VDD.n8203 VDD.n8202 0.000882798
R44007 VDD.n10817 VDD.n10815 0.000872285
R44008 VDD.n7739 VDD.n2272 0.000866563
R44009 VDD.n7810 VDD.n7809 0.000849108
R44010 VDD.n2004 VDD.n2000 0.000810238
R44011 VDD.n2131 VDD.n2130 0.000762697
R44012 VDD.n8209 VDD.n2074 0.000755198
R44013 VDD.n2218 VDD.n2193 0.00072101
R44014 VDD.n11097 VDD.n11096 0.000719801
R44015 VDD.n8247 VDD.n2064 0.000712665
R44016 VDD.n1418 VDD.n1417 0.000706897
R44017 VDD.n1678 VDD.n744 0.000706897
R44018 VDD.n1619 VDD.n783 0.000706897
R44019 VDD.n1352 VDD.n1106 0.000706897
R44020 VDD.n1684 VDD.n741 0.000706897
R44021 VDD.n1697 VDD.n736 0.000706897
R44022 VDD.n1046 VDD.n1045 0.000706897
R44023 VDD.n1721 VDD.n706 0.000706897
R44024 VDD.n7720 VDD.n7719 0.000692009
R44025 VDD.n11064 VDD.n11063 0.000685985
R44026 VDD.n1425 VDD.n844 0.000655172
R44027 VDD.n1691 VDD.n1690 0.000655172
R44028 VDD.n8097 VDD.n8095 0.000655119
R44029 VDD.n11058 VDD.n11057 0.00065217
R44030 VDD.n11078 VDD.n11077 0.00065217
R44031 VDD.n7983 VDD.n2194 0.000622783
R44032 VDD.n7982 VDD.n2196 0.000622783
R44033 VDD.n2195 VDD.n2189 0.000622783
R44034 VDD.n7992 VDD.n2190 0.000622783
R44035 VDD.n2192 VDD.n2191 0.000622783
R44036 VDD.n7989 VDD.n7988 0.000622783
R44037 VDD.n7987 VDD.n7986 0.000622783
R44038 VDD.n2220 VDD.n2219 0.000622783
R44039 VDD.n2223 VDD.n2221 0.000622783
R44040 VDD.n2224 VDD.n2211 0.000622783
R44041 VDD.n2232 VDD.n2231 0.000622783
R44042 VDD.n2213 VDD.n2212 0.000622783
R44043 VDD.n2228 VDD.n2214 0.000622783
R44044 VDD.n2227 VDD.n2217 0.000622783
R44045 VDD.n8161 VDD.n8140 0.000620321
R44046 VDD.n8142 VDD.n2089 0.000620321
R44047 VDD.n5575 VDD.n5553 0.000620321
R44048 VDD.n5556 VDD.n5555 0.000620321
R44049 VDD.n5657 VDD.n5544 0.000620321
R44050 VDD.n5638 VDD.n5546 0.000620321
R44051 VDD.n5840 VDD.n5819 0.000620321
R44052 VDD.n5821 VDD.n5680 0.000620321
R44053 VDD.n5773 VDD.n5752 0.000620321
R44054 VDD.n5754 VDD.n5704 0.000620321
R44055 VDD.n9004 VDD.n8953 0.000620321
R44056 VDD.n9002 VDD.n9001 0.000620321
R44057 VDD.n8833 VDD.n8812 0.000620321
R44058 VDD.n8831 VDD.n8525 0.000620321
R44059 VDD.n9120 VDD.n9099 0.000620321
R44060 VDD.n9118 VDD.n9090 0.000620321
R44061 VDD.n165 VDD.n144 0.000620321
R44062 VDD.n163 VDD.n135 0.000620321
R44063 VDD.n76 VDD.n55 0.000620321
R44064 VDD.n74 VDD.n46 0.000620321
R44065 VDD.n985 VDD.n984 0.000618343
R44066 VDD.n1033 VDD.n1032 0.000618343
R44067 VDD.n1627 VDD.n1626 0.00060181
R44068 VDD.n11048 VDD.n669 0.000601447
R44069 VDD.n11084 VDD.n657 0.000601447
R44070 VDD.n11123 VDD.n640 0.000601447
R44071 VDD.n11120 VDD.n11119 0.000584539
R44072 VDD.n1567 VDD.n782 0.000576357
R44073 VDD.n1566 VDD.n1565 0.000576357
R44074 VDD.n1568 VDD.n1510 0.000576357
R44075 VDD.n1426 VDD.n1425 0.000551724
R44076 VDD.n1431 VDD.n844 0.000551724
R44077 VDD.n1691 VDD.n738 0.000551724
R44078 VDD.n1690 VDD.n739 0.000551724
R44079 VDD.n7780 VDD.n7779 0.000534911
R44080 VDD.n11127 VDD.n11126 0.000533816
R44081 VDD.n11130 VDD.n633 0.000533816
R44082 VDD.n7744 VDD.n2270 0.000517455
R44083 a_52635_49681.n19 a_52635_49681.n17 7.94229
R44084 a_52635_49681.n193 a_52635_49681.n190 7.94229
R44085 a_52635_49681.n147 a_52635_49681.t81 6.58663
R44086 a_52635_49681.n103 a_52635_49681.t2 6.58663
R44087 a_52635_49681.n148 a_52635_49681.n145 5.95439
R44088 a_52635_49681.n104 a_52635_49681.n101 5.95439
R44089 a_52635_49681.n16 a_52635_49681.t111 5.69423
R44090 a_52635_49681.n20 a_52635_49681.t175 5.69423
R44091 a_52635_49681.n192 a_52635_49681.t151 5.69423
R44092 a_52635_49681.n188 a_52635_49681.t120 5.69423
R44093 a_52635_49681.n16 a_52635_49681.n15 5.49558
R44094 a_52635_49681.n192 a_52635_49681.n191 5.49558
R44095 a_52635_49681.n145 a_52635_49681.t9 5.31528
R44096 a_52635_49681.n101 a_52635_49681.t17 5.31528
R44097 a_52635_49681.n0 a_52635_49681.n12 4.22068
R44098 a_52635_49681.n1 a_52635_49681.t126 5.69068
R44099 a_52635_49681.n2 a_52635_49681.n57 4.22068
R44100 a_52635_49681.n3 a_52635_49681.t100 5.69068
R44101 a_52635_49681.n4 a_52635_49681.n56 4.22068
R44102 a_52635_49681.n6 a_52635_49681.n64 3.84173
R44103 a_52635_49681.n9 a_52635_49681.n60 3.84173
R44104 a_52635_49681.n11 a_52635_49681.n197 4.22067
R44105 a_52635_49681.n5 a_52635_49681.t31 5.31173
R44106 a_52635_49681.n7 a_52635_49681.t57 5.31173
R44107 a_52635_49681.n8 a_52635_49681.t27 5.31173
R44108 a_52635_49681.n10 a_52635_49681.t46 5.31173
R44109 a_52635_49681.n144 a_52635_49681.n142 4.50663
R44110 a_52635_49681.n100 a_52635_49681.n59 4.50663
R44111 a_52635_49681.n65 a_52635_49681.n7 4.46113
R44112 a_52635_49681.n19 a_52635_49681.n18 4.22423
R44113 a_52635_49681.n190 a_52635_49681.n189 4.22423
R44114 a_52635_49681.n26 a_52635_49681.t156 4.05054
R44115 a_52635_49681.n31 a_52635_49681.t150 4.05054
R44116 a_52635_49681.n33 a_52635_49681.t147 4.05054
R44117 a_52635_49681.n40 a_52635_49681.t138 4.05054
R44118 a_52635_49681.n42 a_52635_49681.t144 4.05054
R44119 a_52635_49681.n48 a_52635_49681.t142 4.05054
R44120 a_52635_49681.n50 a_52635_49681.t116 4.05054
R44121 a_52635_49681.n21 a_52635_49681.t140 4.05054
R44122 a_52635_49681.n159 a_52635_49681.t131 4.05054
R44123 a_52635_49681.n164 a_52635_49681.t127 4.05054
R44124 a_52635_49681.n166 a_52635_49681.t123 4.05054
R44125 a_52635_49681.n173 a_52635_49681.t105 4.05054
R44126 a_52635_49681.n175 a_52635_49681.t117 4.05054
R44127 a_52635_49681.n181 a_52635_49681.t114 4.05054
R44128 a_52635_49681.n183 a_52635_49681.t94 4.05054
R44129 a_52635_49681.n154 a_52635_49681.t107 4.05054
R44130 a_52635_49681.n150 a_52635_49681.n55 3.97558
R44131 a_52635_49681.n26 a_52635_49681.t135 3.87765
R44132 a_52635_49681.n31 a_52635_49681.t133 3.87765
R44133 a_52635_49681.n33 a_52635_49681.t129 3.87765
R44134 a_52635_49681.n40 a_52635_49681.t109 3.87765
R44135 a_52635_49681.n42 a_52635_49681.t124 3.87765
R44136 a_52635_49681.n48 a_52635_49681.t119 3.87765
R44137 a_52635_49681.n50 a_52635_49681.t98 3.87765
R44138 a_52635_49681.n21 a_52635_49681.t113 3.87765
R44139 a_52635_49681.n159 a_52635_49681.t173 3.87765
R44140 a_52635_49681.n164 a_52635_49681.t169 3.87765
R44141 a_52635_49681.n166 a_52635_49681.t168 3.87765
R44142 a_52635_49681.n173 a_52635_49681.t149 3.87765
R44143 a_52635_49681.n175 a_52635_49681.t164 3.87765
R44144 a_52635_49681.n181 a_52635_49681.t162 3.87765
R44145 a_52635_49681.n183 a_52635_49681.t137 3.87765
R44146 a_52635_49681.n154 a_52635_49681.t154 3.87765
R44147 a_52635_49681.n147 a_52635_49681.n146 3.84528
R44148 a_52635_49681.n144 a_52635_49681.n143 3.84528
R44149 a_52635_49681.n103 a_52635_49681.n102 3.84528
R44150 a_52635_49681.n100 a_52635_49681.n99 3.84528
R44151 a_52635_49681.n136 a_52635_49681.n132 3.79678
R44152 a_52635_49681.n119 a_52635_49681.n115 3.79678
R44153 a_52635_49681.n77 a_52635_49681.n73 3.79678
R44154 a_52635_49681.n92 a_52635_49681.n88 3.79678
R44155 a_52635_49681.n108 a_52635_49681.n10 3.87644
R44156 a_52635_49681.n128 a_52635_49681.n124 3.73034
R44157 a_52635_49681.n97 a_52635_49681.n81 3.73034
R44158 a_52635_49681.n53 a_52635_49681.n20 3.25667
R44159 a_52635_49681.n153 a_52635_49681.n4 3.15553
R44160 a_52635_49681.n54 a_52635_49681.n11 3.15589
R44161 a_52635_49681.n148 a_52635_49681.n147 3.00663
R44162 a_52635_49681.n104 a_52635_49681.n103 3.00663
R44163 a_52635_49681.n111 a_52635_49681.n109 2.7866
R44164 a_52635_49681.n114 a_52635_49681.n112 2.7866
R44165 a_52635_49681.n118 a_52635_49681.n116 2.7866
R44166 a_52635_49681.n122 a_52635_49681.n120 2.7866
R44167 a_52635_49681.n127 a_52635_49681.n125 2.7866
R44168 a_52635_49681.n131 a_52635_49681.n129 2.7866
R44169 a_52635_49681.n135 a_52635_49681.n133 2.7866
R44170 a_52635_49681.n139 a_52635_49681.n137 2.7866
R44171 a_52635_49681.n84 a_52635_49681.n82 2.7866
R44172 a_52635_49681.n87 a_52635_49681.n85 2.7866
R44173 a_52635_49681.n91 a_52635_49681.n89 2.7866
R44174 a_52635_49681.n95 a_52635_49681.n93 2.7866
R44175 a_52635_49681.n80 a_52635_49681.n78 2.7866
R44176 a_52635_49681.n76 a_52635_49681.n74 2.7866
R44177 a_52635_49681.n72 a_52635_49681.n70 2.7866
R44178 a_52635_49681.n68 a_52635_49681.n66 2.7866
R44179 a_52635_49681.n25 a_52635_49681.n21 2.73714
R44180 a_52635_49681.n158 a_52635_49681.n154 2.73714
R44181 a_52635_49681.n30 a_52635_49681.n26 2.73672
R44182 a_52635_49681.n163 a_52635_49681.n159 2.73672
R44183 a_52635_49681.n115 a_52635_49681.n111 2.73672
R44184 a_52635_49681.n88 a_52635_49681.n84 2.73672
R44185 a_52635_49681.n43 a_52635_49681.n41 2.60203
R44186 a_52635_49681.n176 a_52635_49681.n174 2.60203
R44187 a_52635_49681.n29 a_52635_49681.n28 2.58054
R44188 a_52635_49681.n38 a_52635_49681.n37 2.58054
R44189 a_52635_49681.n46 a_52635_49681.n45 2.58054
R44190 a_52635_49681.n24 a_52635_49681.n23 2.58054
R44191 a_52635_49681.n162 a_52635_49681.n161 2.58054
R44192 a_52635_49681.n171 a_52635_49681.n170 2.58054
R44193 a_52635_49681.n179 a_52635_49681.n178 2.58054
R44194 a_52635_49681.n157 a_52635_49681.n156 2.58054
R44195 a_52635_49681.n51 a_52635_49681.n49 2.53418
R44196 a_52635_49681.n34 a_52635_49681.n32 2.53418
R44197 a_52635_49681.n184 a_52635_49681.n182 2.53418
R44198 a_52635_49681.n167 a_52635_49681.n165 2.53418
R44199 a_52635_49681.n188 a_52635_49681.n187 2.51873
R44200 a_52635_49681.n29 a_52635_49681.n27 2.40765
R44201 a_52635_49681.n38 a_52635_49681.n36 2.40765
R44202 a_52635_49681.n46 a_52635_49681.n44 2.40765
R44203 a_52635_49681.n24 a_52635_49681.n22 2.40765
R44204 a_52635_49681.n162 a_52635_49681.n160 2.40765
R44205 a_52635_49681.n171 a_52635_49681.n169 2.40765
R44206 a_52635_49681.n179 a_52635_49681.n177 2.40765
R44207 a_52635_49681.n157 a_52635_49681.n155 2.40765
R44208 a_52635_49681.n107 a_52635_49681.n8 2.37644
R44209 a_52635_49681.n63 a_52635_49681.n5 2.37644
R44210 a_52635_49681.n17 a_52635_49681.n13 2.23844
R44211 a_52635_49681.n111 a_52635_49681.n110 2.2016
R44212 a_52635_49681.n114 a_52635_49681.n113 2.2016
R44213 a_52635_49681.n118 a_52635_49681.n117 2.2016
R44214 a_52635_49681.n122 a_52635_49681.n121 2.2016
R44215 a_52635_49681.n127 a_52635_49681.n126 2.2016
R44216 a_52635_49681.n131 a_52635_49681.n130 2.2016
R44217 a_52635_49681.n135 a_52635_49681.n134 2.2016
R44218 a_52635_49681.n139 a_52635_49681.n138 2.2016
R44219 a_52635_49681.n84 a_52635_49681.n83 2.2016
R44220 a_52635_49681.n87 a_52635_49681.n86 2.2016
R44221 a_52635_49681.n91 a_52635_49681.n90 2.2016
R44222 a_52635_49681.n95 a_52635_49681.n94 2.2016
R44223 a_52635_49681.n80 a_52635_49681.n79 2.2016
R44224 a_52635_49681.n76 a_52635_49681.n75 2.2016
R44225 a_52635_49681.n72 a_52635_49681.n71 2.2016
R44226 a_52635_49681.n68 a_52635_49681.n67 2.2016
R44227 a_52635_49681.n98 a_52635_49681.n63 2.0852
R44228 a_52635_49681.n142 a_52635_49681.n55 1.85726
R44229 a_52635_49681.n151 a_52635_49681.n150 1.83738
R44230 a_52635_49681.n141 a_52635_49681.n140 1.65018
R44231 a_52635_49681.n69 a_52635_49681.n65 1.65018
R44232 a_52635_49681.n152 a_52635_49681.n2 1.65553
R44233 a_52635_49681.n196 a_52635_49681.n0 1.65553
R44234 a_52635_49681.n186 a_52635_49681.n185 1.5005
R44235 a_52635_49681.n53 a_52635_49681.n52 1.5005
R44236 a_52635_49681.n105 a_52635_49681.n104 1.5005
R44237 a_52635_49681.n107 a_52635_49681.n106 1.5005
R44238 a_52635_49681.n149 a_52635_49681.n148 1.5005
R44239 a_52635_49681.n98 a_52635_49681.n97 1.5005
R44240 a_52635_49681.n124 a_52635_49681.n58 1.5005
R44241 a_52635_49681.n152 a_52635_49681.n151 1.5005
R44242 a_52635_49681.n168 a_52635_49681.n14 1.5005
R44243 a_52635_49681.n194 a_52635_49681.n193 1.5005
R44244 a_52635_49681.n35 a_52635_49681.n13 1.5005
R44245 a_52635_49681.n196 a_52635_49681.n195 1.5005
R44246 a_52635_49681.n12 a_52635_49681.t121 1.4705
R44247 a_52635_49681.n12 a_52635_49681.t93 1.4705
R44248 a_52635_49681.n15 a_52635_49681.t88 1.4705
R44249 a_52635_49681.n15 a_52635_49681.t128 1.4705
R44250 a_52635_49681.n18 a_52635_49681.t170 1.4705
R44251 a_52635_49681.n18 a_52635_49681.t115 1.4705
R44252 a_52635_49681.n27 a_52635_49681.t91 1.4705
R44253 a_52635_49681.n27 a_52635_49681.t166 1.4705
R44254 a_52635_49681.n28 a_52635_49681.t108 1.4705
R44255 a_52635_49681.n28 a_52635_49681.t97 1.4705
R44256 a_52635_49681.n36 a_52635_49681.t155 1.4705
R44257 a_52635_49681.n36 a_52635_49681.t125 1.4705
R44258 a_52635_49681.n37 a_52635_49681.t89 1.4705
R44259 a_52635_49681.n37 a_52635_49681.t145 1.4705
R44260 a_52635_49681.n44 a_52635_49681.t163 1.4705
R44261 a_52635_49681.n44 a_52635_49681.t134 1.4705
R44262 a_52635_49681.n45 a_52635_49681.t96 1.4705
R44263 a_52635_49681.n45 a_52635_49681.t153 1.4705
R44264 a_52635_49681.n22 a_52635_49681.t143 1.4705
R44265 a_52635_49681.n22 a_52635_49681.t112 1.4705
R44266 a_52635_49681.n23 a_52635_49681.t171 1.4705
R44267 a_52635_49681.n23 a_52635_49681.t139 1.4705
R44268 a_52635_49681.n191 a_52635_49681.t122 1.4705
R44269 a_52635_49681.n191 a_52635_49681.t167 1.4705
R44270 a_52635_49681.n189 a_52635_49681.t110 1.4705
R44271 a_52635_49681.n189 a_52635_49681.t157 1.4705
R44272 a_52635_49681.n160 a_52635_49681.t132 1.4705
R44273 a_52635_49681.n160 a_52635_49681.t104 1.4705
R44274 a_52635_49681.n161 a_52635_49681.t90 1.4705
R44275 a_52635_49681.n161 a_52635_49681.t161 1.4705
R44276 a_52635_49681.n169 a_52635_49681.t101 1.4705
R44277 a_52635_49681.n169 a_52635_49681.t165 1.4705
R44278 a_52635_49681.n170 a_52635_49681.t148 1.4705
R44279 a_52635_49681.n170 a_52635_49681.t118 1.4705
R44280 a_52635_49681.n177 a_52635_49681.t103 1.4705
R44281 a_52635_49681.n177 a_52635_49681.t172 1.4705
R44282 a_52635_49681.n178 a_52635_49681.t160 1.4705
R44283 a_52635_49681.n178 a_52635_49681.t130 1.4705
R44284 a_52635_49681.n155 a_52635_49681.t95 1.4705
R44285 a_52635_49681.n155 a_52635_49681.t152 1.4705
R44286 a_52635_49681.n156 a_52635_49681.t141 1.4705
R44287 a_52635_49681.n156 a_52635_49681.t106 1.4705
R44288 a_52635_49681.n57 a_52635_49681.t99 1.4705
R44289 a_52635_49681.n57 a_52635_49681.t159 1.4705
R44290 a_52635_49681.n56 a_52635_49681.t158 1.4705
R44291 a_52635_49681.n56 a_52635_49681.t146 1.4705
R44292 a_52635_49681.n62 a_52635_49681.t55 1.4705
R44293 a_52635_49681.n62 a_52635_49681.t26 1.4705
R44294 a_52635_49681.n64 a_52635_49681.t62 1.4705
R44295 a_52635_49681.n64 a_52635_49681.t29 1.4705
R44296 a_52635_49681.n109 a_52635_49681.t48 1.4705
R44297 a_52635_49681.n109 a_52635_49681.t70 1.4705
R44298 a_52635_49681.n110 a_52635_49681.t43 1.4705
R44299 a_52635_49681.n110 a_52635_49681.t66 1.4705
R44300 a_52635_49681.n112 a_52635_49681.t74 1.4705
R44301 a_52635_49681.n112 a_52635_49681.t35 1.4705
R44302 a_52635_49681.n113 a_52635_49681.t68 1.4705
R44303 a_52635_49681.n113 a_52635_49681.t30 1.4705
R44304 a_52635_49681.n116 a_52635_49681.t84 1.4705
R44305 a_52635_49681.n116 a_52635_49681.t78 1.4705
R44306 a_52635_49681.n117 a_52635_49681.t72 1.4705
R44307 a_52635_49681.n117 a_52635_49681.t69 1.4705
R44308 a_52635_49681.n120 a_52635_49681.t16 1.4705
R44309 a_52635_49681.n120 a_52635_49681.t58 1.4705
R44310 a_52635_49681.n121 a_52635_49681.t7 1.4705
R44311 a_52635_49681.n121 a_52635_49681.t50 1.4705
R44312 a_52635_49681.n125 a_52635_49681.t71 1.4705
R44313 a_52635_49681.n125 a_52635_49681.t85 1.4705
R44314 a_52635_49681.n126 a_52635_49681.t67 1.4705
R44315 a_52635_49681.n126 a_52635_49681.t73 1.4705
R44316 a_52635_49681.n129 a_52635_49681.t3 1.4705
R44317 a_52635_49681.n129 a_52635_49681.t49 1.4705
R44318 a_52635_49681.n130 a_52635_49681.t80 1.4705
R44319 a_52635_49681.n130 a_52635_49681.t44 1.4705
R44320 a_52635_49681.n133 a_52635_49681.t13 1.4705
R44321 a_52635_49681.n133 a_52635_49681.t32 1.4705
R44322 a_52635_49681.n134 a_52635_49681.t1 1.4705
R44323 a_52635_49681.n134 a_52635_49681.t28 1.4705
R44324 a_52635_49681.n137 a_52635_49681.t12 1.4705
R44325 a_52635_49681.n137 a_52635_49681.t63 1.4705
R44326 a_52635_49681.n138 a_52635_49681.t0 1.4705
R44327 a_52635_49681.n138 a_52635_49681.t59 1.4705
R44328 a_52635_49681.n82 a_52635_49681.t54 1.4705
R44329 a_52635_49681.n82 a_52635_49681.t77 1.4705
R44330 a_52635_49681.n83 a_52635_49681.t51 1.4705
R44331 a_52635_49681.n83 a_52635_49681.t75 1.4705
R44332 a_52635_49681.n85 a_52635_49681.t83 1.4705
R44333 a_52635_49681.n85 a_52635_49681.t37 1.4705
R44334 a_52635_49681.n86 a_52635_49681.t82 1.4705
R44335 a_52635_49681.n86 a_52635_49681.t36 1.4705
R44336 a_52635_49681.n89 a_52635_49681.t6 1.4705
R44337 a_52635_49681.n89 a_52635_49681.t87 1.4705
R44338 a_52635_49681.n90 a_52635_49681.t4 1.4705
R44339 a_52635_49681.n90 a_52635_49681.t86 1.4705
R44340 a_52635_49681.n93 a_52635_49681.t24 1.4705
R44341 a_52635_49681.n93 a_52635_49681.t61 1.4705
R44342 a_52635_49681.n94 a_52635_49681.t23 1.4705
R44343 a_52635_49681.n94 a_52635_49681.t60 1.4705
R44344 a_52635_49681.n78 a_52635_49681.t79 1.4705
R44345 a_52635_49681.n78 a_52635_49681.t8 1.4705
R44346 a_52635_49681.n79 a_52635_49681.t76 1.4705
R44347 a_52635_49681.n79 a_52635_49681.t5 1.4705
R44348 a_52635_49681.n74 a_52635_49681.t11 1.4705
R44349 a_52635_49681.n74 a_52635_49681.t56 1.4705
R44350 a_52635_49681.n75 a_52635_49681.t10 1.4705
R44351 a_52635_49681.n75 a_52635_49681.t53 1.4705
R44352 a_52635_49681.n70 a_52635_49681.t21 1.4705
R44353 a_52635_49681.n70 a_52635_49681.t34 1.4705
R44354 a_52635_49681.n71 a_52635_49681.t19 1.4705
R44355 a_52635_49681.n71 a_52635_49681.t33 1.4705
R44356 a_52635_49681.n66 a_52635_49681.t20 1.4705
R44357 a_52635_49681.n66 a_52635_49681.t65 1.4705
R44358 a_52635_49681.n67 a_52635_49681.t18 1.4705
R44359 a_52635_49681.n67 a_52635_49681.t64 1.4705
R44360 a_52635_49681.n146 a_52635_49681.t14 1.4705
R44361 a_52635_49681.n146 a_52635_49681.t38 1.4705
R44362 a_52635_49681.n143 a_52635_49681.t39 1.4705
R44363 a_52635_49681.n143 a_52635_49681.t42 1.4705
R44364 a_52635_49681.n61 a_52635_49681.t45 1.4705
R44365 a_52635_49681.n61 a_52635_49681.t15 1.4705
R44366 a_52635_49681.n60 a_52635_49681.t52 1.4705
R44367 a_52635_49681.n60 a_52635_49681.t25 1.4705
R44368 a_52635_49681.n102 a_52635_49681.t22 1.4705
R44369 a_52635_49681.n102 a_52635_49681.t40 1.4705
R44370 a_52635_49681.n99 a_52635_49681.t41 1.4705
R44371 a_52635_49681.n99 a_52635_49681.t47 1.4705
R44372 a_52635_49681.n197 a_52635_49681.t92 1.4705
R44373 a_52635_49681.t174 a_52635_49681.n197 1.4705
R44374 a_52635_49681.n30 a_52635_49681.n29 1.46537
R44375 a_52635_49681.n32 a_52635_49681.n31 1.46537
R44376 a_52635_49681.n39 a_52635_49681.n38 1.46537
R44377 a_52635_49681.n41 a_52635_49681.n40 1.46537
R44378 a_52635_49681.n43 a_52635_49681.n42 1.46537
R44379 a_52635_49681.n47 a_52635_49681.n46 1.46537
R44380 a_52635_49681.n49 a_52635_49681.n48 1.46537
R44381 a_52635_49681.n25 a_52635_49681.n24 1.46537
R44382 a_52635_49681.n163 a_52635_49681.n162 1.46537
R44383 a_52635_49681.n165 a_52635_49681.n164 1.46537
R44384 a_52635_49681.n172 a_52635_49681.n171 1.46537
R44385 a_52635_49681.n174 a_52635_49681.n173 1.46537
R44386 a_52635_49681.n176 a_52635_49681.n175 1.46537
R44387 a_52635_49681.n180 a_52635_49681.n179 1.46537
R44388 a_52635_49681.n182 a_52635_49681.n181 1.46537
R44389 a_52635_49681.n158 a_52635_49681.n157 1.46537
R44390 a_52635_49681.n115 a_52635_49681.n114 1.46537
R44391 a_52635_49681.n119 a_52635_49681.n118 1.46537
R44392 a_52635_49681.n123 a_52635_49681.n122 1.46537
R44393 a_52635_49681.n128 a_52635_49681.n127 1.46537
R44394 a_52635_49681.n132 a_52635_49681.n131 1.46537
R44395 a_52635_49681.n136 a_52635_49681.n135 1.46537
R44396 a_52635_49681.n140 a_52635_49681.n139 1.46537
R44397 a_52635_49681.n88 a_52635_49681.n87 1.46537
R44398 a_52635_49681.n92 a_52635_49681.n91 1.46537
R44399 a_52635_49681.n96 a_52635_49681.n95 1.46537
R44400 a_52635_49681.n81 a_52635_49681.n80 1.46537
R44401 a_52635_49681.n77 a_52635_49681.n76 1.46537
R44402 a_52635_49681.n73 a_52635_49681.n72 1.46537
R44403 a_52635_49681.n69 a_52635_49681.n68 1.46537
R44404 a_52635_49681.n34 a_52635_49681.n33 1.46535
R44405 a_52635_49681.n51 a_52635_49681.n50 1.46535
R44406 a_52635_49681.n167 a_52635_49681.n166 1.46535
R44407 a_52635_49681.n184 a_52635_49681.n183 1.46535
R44408 a_52635_49681.n20 a_52635_49681.n19 1.27228
R44409 a_52635_49681.n49 a_52635_49681.n47 1.27228
R44410 a_52635_49681.n47 a_52635_49681.n43 1.27228
R44411 a_52635_49681.n41 a_52635_49681.n39 1.27228
R44412 a_52635_49681.n32 a_52635_49681.n30 1.27228
R44413 a_52635_49681.n190 a_52635_49681.n188 1.27228
R44414 a_52635_49681.n182 a_52635_49681.n180 1.27228
R44415 a_52635_49681.n180 a_52635_49681.n176 1.27228
R44416 a_52635_49681.n174 a_52635_49681.n172 1.27228
R44417 a_52635_49681.n165 a_52635_49681.n163 1.27228
R44418 a_52635_49681.n140 a_52635_49681.n136 1.27228
R44419 a_52635_49681.n132 a_52635_49681.n128 1.27228
R44420 a_52635_49681.n123 a_52635_49681.n119 1.27228
R44421 a_52635_49681.n73 a_52635_49681.n69 1.27228
R44422 a_52635_49681.n81 a_52635_49681.n77 1.27228
R44423 a_52635_49681.n96 a_52635_49681.n92 1.27228
R44424 a_52635_49681.n145 a_52635_49681.n144 1.27228
R44425 a_52635_49681.n101 a_52635_49681.n100 1.27228
R44426 a_52635_49681.n150 a_52635_49681.n149 1.25341
R44427 a_52635_49681.n153 a_52635_49681.n55 1.23151
R44428 a_52635_49681.n17 a_52635_49681.n16 1.01873
R44429 a_52635_49681.n193 a_52635_49681.n192 1.01873
R44430 a_52635_49681.n54 a_52635_49681.n53 0.778574
R44431 a_52635_49681.n186 a_52635_49681.n153 0.778574
R44432 a_52635_49681.n195 a_52635_49681.n13 0.778574
R44433 a_52635_49681.n151 a_52635_49681.n14 0.778574
R44434 a_52635_49681.n187 a_52635_49681.n186 0.738439
R44435 a_52635_49681.n194 a_52635_49681.n14 0.738439
R44436 a_52635_49681.n142 a_52635_49681.n141 0.737223
R44437 a_52635_49681.n65 a_52635_49681.n59 0.737223
R44438 a_52635_49681.n149 a_52635_49681.n58 0.737223
R44439 a_52635_49681.n105 a_52635_49681.n98 0.737223
R44440 a_52635_49681.n108 a_52635_49681.n59 0.725061
R44441 a_52635_49681.n106 a_52635_49681.n105 0.725061
R44442 a_52635_49681.n52 a_52635_49681.n51 0.699581
R44443 a_52635_49681.n35 a_52635_49681.n34 0.699581
R44444 a_52635_49681.n185 a_52635_49681.n184 0.699581
R44445 a_52635_49681.n168 a_52635_49681.n167 0.699581
R44446 a_52635_49681.n141 a_52635_49681.n108 0.585196
R44447 a_52635_49681.n106 a_52635_49681.n58 0.585196
R44448 a_52635_49681.n52 a_52635_49681.n25 0.557791
R44449 a_52635_49681.n39 a_52635_49681.n35 0.557791
R44450 a_52635_49681.n185 a_52635_49681.n158 0.557791
R44451 a_52635_49681.n172 a_52635_49681.n168 0.557791
R44452 a_52635_49681.n187 a_52635_49681.n54 0.530466
R44453 a_52635_49681.n195 a_52635_49681.n194 0.530466
R44454 a_52635_49681.n124 a_52635_49681.n123 0.150184
R44455 a_52635_49681.n97 a_52635_49681.n96 0.150184
R44456 a_52635_49681.n3 a_52635_49681.n4 1.27228
R44457 a_52635_49681.n152 a_52635_49681.n3 7.30549
R44458 a_52635_49681.t102 a_52635_49681.n2 6.96214
R44459 a_52635_49681.n9 a_52635_49681.n10 1.26457
R44460 a_52635_49681.n107 a_52635_49681.n9 6.59229
R44461 a_52635_49681.n61 a_52635_49681.n8 5.10549
R44462 a_52635_49681.n6 a_52635_49681.n7 1.26457
R44463 a_52635_49681.n63 a_52635_49681.n6 6.59229
R44464 a_52635_49681.n62 a_52635_49681.n5 5.10549
R44465 a_52635_49681.n11 a_52635_49681.n1 1.27192
R44466 a_52635_49681.n196 a_52635_49681.n1 7.30549
R44467 a_52635_49681.t136 a_52635_49681.n0 6.96214
R44468 a_57977_n12421.t0 a_57977_n12421.t1 93.1589
R44469 a_57977_n12421.t0 a_57977_n12421.t2 24.9014
R44470 a_100820_11614.n2 a_100820_11614.t19 12.8637
R44471 a_100820_11614.n1 a_100820_11614.t3 10.7018
R44472 a_100820_11614.n1 a_100820_11614.t6 10.1659
R44473 a_100820_11614.n1 a_100820_11614.t5 9.64387
R44474 a_100820_11614.n1 a_100820_11614.t2 9.27665
R44475 a_100820_11614.n1 a_100820_11614.n2 8.75198
R44476 a_100820_11614.n2 a_100820_11614.t14 8.14051
R44477 a_100820_11614.n2 a_100820_11614.t10 8.14051
R44478 a_100820_11614.n2 a_100820_11614.t8 8.14051
R44479 a_100820_11614.n2 a_100820_11614.t17 8.14051
R44480 a_100820_11614.n2 a_100820_11614.t21 8.06917
R44481 a_100820_11614.n2 a_100820_11614.t18 8.06917
R44482 a_100820_11614.n2 a_100820_11614.t11 8.06917
R44483 a_100820_11614.n2 a_100820_11614.t15 8.06917
R44484 a_100820_11614.n2 a_100820_11614.t13 8.06917
R44485 a_100820_11614.n2 a_100820_11614.t23 8.06917
R44486 a_100820_11614.n2 a_100820_11614.t9 8.06917
R44487 a_100820_11614.n0 a_100820_11614.t7 7.94068
R44488 a_100820_11614.t0 a_100820_11614.n1 7.72524
R44489 a_100820_11614.n0 a_100820_11614.t4 7.22855
R44490 a_100820_11614.n1 a_100820_11614.t1 7.17942
R44491 a_100820_11614.t16 a_100820_11614.n2 8.33649
R44492 a_100820_11614.n2 a_100820_11614.t20 8.33649
R44493 a_100820_11614.t22 a_100820_11614.n2 8.33556
R44494 a_100820_11614.n2 a_100820_11614.t12 8.33556
R44495 a_100820_11614.n1 a_100820_11614.n0 7.46075
R44496 a_30324_4421.t2 a_30324_4421.t0 21.6693
R44497 a_30324_4421.t1 a_30324_4421.t0 15.3476
R44498 a_31284_4481.t0 a_31284_4481.t2 41.3314
R44499 a_31284_4481.t2 a_31284_4481.t1 15.0742
R44500 a_100820_10448.n0 a_100820_10448.t7 10.2828
R44501 a_100820_10448.t0 a_100820_10448.t5 10.2828
R44502 a_100820_10448.n0 a_100820_10448.t17 10.2828
R44503 a_100820_10448.n0 a_100820_10448.t13 10.2828
R44504 a_100820_10448.n0 a_100820_10448.t20 10.1333
R44505 a_100820_10448.t0 a_100820_10448.t21 10.1333
R44506 a_100820_10448.n0 a_100820_10448.t3 10.1333
R44507 a_100820_10448.n0 a_100820_10448.t9 10.1333
R44508 a_100820_10448.n0 a_100820_10448.t16 9.57156
R44509 a_100820_10448.n0 a_100820_10448.t14 9.57156
R44510 a_100820_10448.t0 a_100820_10448.t15 9.57156
R44511 a_100820_10448.n0 a_100820_10448.t11 9.57156
R44512 a_100820_10448.n0 a_100820_10448.t22 9.57156
R44513 a_100820_10448.n0 a_100820_10448.t18 9.57156
R44514 a_100820_10448.t0 a_100820_10448.t19 9.57156
R44515 a_100820_10448.n0 a_100820_10448.t12 9.57156
R44516 a_100820_10448.t0 a_100820_10448.n1 8.94763
R44517 a_100820_10448.t0 a_100820_10448.t2 8.02945
R44518 a_100820_10448.t0 a_100820_10448.t1 8.02708
R44519 a_100820_10448.t0 a_100820_10448.t8 7.90829
R44520 a_100820_10448.n1 a_100820_10448.t6 7.90829
R44521 a_100820_10448.n1 a_100820_10448.t10 7.41776
R44522 a_100820_10448.t4 a_100820_10448.t0 7.41776
R44523 a_100820_10448.t0 a_100820_10448.n0 7.31642
R44524 a_53829_n36382.n5 a_53829_n36382.n1 10.2377
R44525 a_53829_n36382.n4 a_53829_n36382.t0 10.2105
R44526 a_53829_n36382.n4 a_53829_n36382.t1 9.99998
R44527 a_53829_n36382.n5 a_53829_n36382.t7 9.80532
R44528 a_53829_n36382.n5 a_53829_n36382.t5 9.55206
R44529 a_53829_n36382.n0 a_53829_n36382.t9 8.17385
R44530 a_53829_n36382.n3 a_53829_n36382.t21 8.17299
R44531 a_53829_n36382.n3 a_53829_n36382.t10 8.17134
R44532 a_53829_n36382.n0 a_53829_n36382.t23 8.16754
R44533 a_53829_n36382.n1 a_53829_n36382.t17 8.10567
R44534 a_53829_n36382.n1 a_53829_n36382.t20 8.10567
R44535 a_53829_n36382.n3 a_53829_n36382.t16 8.10567
R44536 a_53829_n36382.n3 a_53829_n36382.t11 8.10567
R44537 a_53829_n36382.n1 a_53829_n36382.t18 8.10567
R44538 a_53829_n36382.n1 a_53829_n36382.t19 8.10567
R44539 a_53829_n36382.n0 a_53829_n36382.t15 8.10567
R44540 a_53829_n36382.n0 a_53829_n36382.t14 8.10567
R44541 a_53829_n36382.n6 a_53829_n36382.t3 7.74888
R44542 a_53829_n36382.n7 a_53829_n36382.t6 7.73141
R44543 a_53829_n36382.n6 a_53829_n36382.t2 7.46359
R44544 a_53829_n36382.t4 a_53829_n36382.n7 7.13081
R44545 a_53829_n36382.n4 a_53829_n36382.n6 2.2505
R44546 a_53829_n36382.n7 a_53829_n36382.n5 2.2505
R44547 a_53829_n36382.t8 a_53829_n36382.n1 8.35729
R44548 a_53829_n36382.n1 a_53829_n36382.t22 8.37586
R44549 a_53829_n36382.n0 a_53829_n36382.t12 8.38104
R44550 a_53829_n36382.n1 a_53829_n36382.n0 4.35658
R44551 a_53829_n36382.n5 a_53829_n36382.n4 2.96863
R44552 a_53829_n36382.n2 a_53829_n36382.n1 1.08819
R44553 a_53829_n36382.n2 a_53829_n36382.n3 1.08408
R44554 a_53829_n36382.n2 a_53829_n36382.t13 8.6675
R44555 a_36032_n36322.n1 a_36032_n36322.n0 26.5241
R44556 a_36032_n36322.n0 a_36032_n36322.t3 11.5094
R44557 a_36032_n36322.t0 a_36032_n36322.n1 10.937
R44558 a_36032_n36322.n1 a_36032_n36322.t1 9.33982
R44559 a_36032_n36322.n0 a_36032_n36322.t2 9.24966
R44560 a_35502_25545.n345 a_35502_25545.t22 10.621
R44561 a_35502_25545.n349 a_35502_25545.t71 10.621
R44562 a_35502_25545.n342 a_35502_25545.n326 10.3121
R44563 a_35502_25545.n347 a_35502_25545.t91 10.3044
R44564 a_35502_25545.n351 a_35502_25545.t20 10.3044
R44565 a_35502_25545.n346 a_35502_25545.t48 9.9994
R44566 a_35502_25545.n350 a_35502_25545.t26 9.9994
R44567 a_35502_25545.n345 a_35502_25545.t24 9.999
R44568 a_35502_25545.n349 a_35502_25545.t62 9.999
R44569 a_35502_25545.n224 a_35502_25545.t39 8.33806
R44570 a_35502_25545.n319 a_35502_25545.t64 8.3366
R44571 a_35502_25545.n278 a_35502_25545.t35 8.26493
R44572 a_35502_25545.n96 a_35502_25545.t69 8.35715
R44573 a_35502_25545.n43 a_35502_25545.t81 8.06917
R44574 a_35502_25545.n55 a_35502_25545.t77 8.06917
R44575 a_35502_25545.n122 a_35502_25545.t102 8.06917
R44576 a_35502_25545.n31 a_35502_25545.t85 8.06917
R44577 a_35502_25545.n132 a_35502_25545.t30 8.06917
R44578 a_35502_25545.n50 a_35502_25545.t47 8.06917
R44579 a_35502_25545.n57 a_35502_25545.t51 8.06917
R44580 a_35502_25545.n17 a_35502_25545.t80 8.06917
R44581 a_35502_25545.n78 a_35502_25545.t100 8.06917
R44582 a_35502_25545.n28 a_35502_25545.t45 8.06917
R44583 a_35502_25545.n133 a_35502_25545.t72 8.06917
R44584 a_35502_25545.n9 a_35502_25545.t29 8.06917
R44585 a_35502_25545.n8 a_35502_25545.t59 8.06917
R44586 a_35502_25545.n170 a_35502_25545.t56 8.06917
R44587 a_35502_25545.n6 a_35502_25545.t57 8.06917
R44588 a_35502_25545.n5 a_35502_25545.t86 8.06917
R44589 a_35502_25545.n175 a_35502_25545.t83 8.06917
R44590 a_35502_25545.n40 a_35502_25545.t76 8.06917
R44591 a_35502_25545.n93 a_35502_25545.t44 8.06917
R44592 a_35502_25545.n75 a_35502_25545.t78 8.06917
R44593 a_35502_25545.n61 a_35502_25545.t103 8.06917
R44594 a_35502_25545.n34 a_35502_25545.t41 8.06917
R44595 a_35502_25545.n90 a_35502_25545.t49 8.06917
R44596 a_35502_25545.n2 a_35502_25545.t75 8.06917
R44597 a_35502_25545.n86 a_35502_25545.t95 8.06917
R44598 a_35502_25545.n71 a_35502_25545.t40 8.06917
R44599 a_35502_25545.n65 a_35502_25545.t68 8.06917
R44600 a_35502_25545.n125 a_35502_25545.t28 8.06917
R44601 a_35502_25545.n23 a_35502_25545.t54 8.06917
R44602 a_35502_25545.n163 a_35502_25545.t52 8.06917
R44603 a_35502_25545.n128 a_35502_25545.t53 8.06917
R44604 a_35502_25545.n20 a_35502_25545.t82 8.06917
R44605 a_35502_25545.n152 a_35502_25545.t79 8.06917
R44606 a_35502_25545.n82 a_35502_25545.t73 8.06917
R44607 a_35502_25545.n68 a_35502_25545.t96 8.06917
R44608 a_35502_25545.n108 a_35502_25545.t66 8.06917
R44609 a_35502_25545.n97 a_35502_25545.t74 8.06917
R44610 a_35502_25545.n259 a_35502_25545.t97 8.06917
R44611 a_35502_25545.n248 a_35502_25545.t36 8.06917
R44612 a_35502_25545.n247 a_35502_25545.t42 8.06917
R44613 a_35502_25545.n246 a_35502_25545.t88 8.06917
R44614 a_35502_25545.n95 a_35502_25545.t101 8.06917
R44615 a_35502_25545.n239 a_35502_25545.t46 8.06917
R44616 a_35502_25545.n112 a_35502_25545.t98 8.06917
R44617 a_35502_25545.n225 a_35502_25545.t94 8.06917
R44618 a_35502_25545.n231 a_35502_25545.t63 8.06917
R44619 a_35502_25545.n232 a_35502_25545.t67 8.06917
R44620 a_35502_25545.n233 a_35502_25545.t38 8.06917
R44621 a_35502_25545.n109 a_35502_25545.t37 8.06917
R44622 a_35502_25545.n100 a_35502_25545.t65 8.06917
R44623 a_35502_25545.n267 a_35502_25545.t89 8.06917
R44624 a_35502_25545.n318 a_35502_25545.t99 8.06917
R44625 a_35502_25545.n118 a_35502_25545.t43 8.06917
R44626 a_35502_25545.n316 a_35502_25545.t84 8.06917
R44627 a_35502_25545.n315 a_35502_25545.t33 8.06917
R44628 a_35502_25545.n314 a_35502_25545.t31 8.06917
R44629 a_35502_25545.n312 a_35502_25545.t61 8.06917
R44630 a_35502_25545.n305 a_35502_25545.t70 8.06917
R44631 a_35502_25545.n115 a_35502_25545.t92 8.06917
R44632 a_35502_25545.n300 a_35502_25545.t34 8.06917
R44633 a_35502_25545.n101 a_35502_25545.t60 8.06917
R44634 a_35502_25545.n119 a_35502_25545.t87 8.06917
R44635 a_35502_25545.n289 a_35502_25545.t32 8.06917
R44636 a_35502_25545.n288 a_35502_25545.t58 8.06917
R44637 a_35502_25545.n287 a_35502_25545.t55 8.06917
R44638 a_35502_25545.n274 a_35502_25545.t93 8.06917
R44639 a_35502_25545.n277 a_35502_25545.t90 8.06917
R44640 a_35502_25545.n330 a_35502_25545.t5 6.49245
R44641 a_35502_25545.n327 a_35502_25545.t17 6.49245
R44642 a_35502_25545.n138 a_35502_25545.t2 6.50349
R44643 a_35502_25545.n343 a_35502_25545.t23 5.70664
R44644 a_35502_25545.n353 a_35502_25545.t21 5.23357
R44645 a_35502_25545.n328 a_35502_25545.t19 5.22068
R44646 a_35502_25545.t27 a_35502_25545.n353 5.15077
R44647 a_35502_25545.n343 a_35502_25545.t25 4.6582
R44648 a_35502_25545.n84 a_35502_25545.n69 2.0194
R44649 a_35502_25545.n178 a_35502_25545.n123 2.42484
R44650 a_35502_25545.n123 a_35502_25545.n177 2.4256
R44651 a_35502_25545.n110 a_35502_25545.n109 2.25048
R44652 a_35502_25545.n115 a_35502_25545.n113 2.25048
R44653 a_35502_25545.n134 a_35502_25545.t4 5.23239
R44654 a_35502_25545.n135 a_35502_25545.t12 5.23239
R44655 a_35502_25545.n339 a_35502_25545.n338 4.60825
R44656 a_35502_25545.t8 a_35502_25545.n138 5.23239
R44657 a_35502_25545.n10 a_35502_25545.n9 1.44552
R44658 a_35502_25545.n7 a_35502_25545.n6 1.44552
R44659 a_35502_25545.n126 a_35502_25545.n125 2.22591
R44660 a_35502_25545.n129 a_35502_25545.n128 2.22591
R44661 a_35502_25545.n85 a_35502_25545.n159 4.51491
R44662 a_35502_25545.n216 a_35502_25545.n215 4.51075
R44663 a_35502_25545.n62 a_35502_25545.n61 2.21906
R44664 a_35502_25545.n66 a_35502_25545.n65 2.21906
R44665 a_35502_25545.n34 a_35502_25545.n35 2.21826
R44666 a_35502_25545.n40 a_35502_25545.n39 2.21826
R44667 a_35502_25545.n338 a_35502_25545.n334 4.50168
R44668 a_35502_25545.n12 a_35502_25545.n5 2.21666
R44669 a_35502_25545.n11 a_35502_25545.n174 4.5005
R44670 a_35502_25545.n184 a_35502_25545.n183 4.5005
R44671 a_35502_25545.n14 a_35502_25545.n8 2.21666
R44672 a_35502_25545.n13 a_35502_25545.n169 4.5005
R44673 a_35502_25545.n202 a_35502_25545.n201 4.5005
R44674 a_35502_25545.n194 a_35502_25545.n193 4.5005
R44675 a_35502_25545.n78 a_35502_25545.n79 2.21666
R44676 a_35502_25545.n191 a_35502_25545.n27 4.5005
R44677 a_35502_25545.n28 a_35502_25545.n25 2.21666
R44678 a_35502_25545.n26 a_35502_25545.n190 4.5005
R44679 a_35502_25545.n189 a_35502_25545.n133 4.5005
R44680 a_35502_25545.n188 a_35502_25545.n187 4.5005
R44681 a_35502_25545.n51 a_35502_25545.n50 2.21666
R44682 a_35502_25545.n196 a_35502_25545.n49 4.5005
R44683 a_35502_25545.n198 a_35502_25545.n197 4.5005
R44684 a_35502_25545.n58 a_35502_25545.n57 2.21666
R44685 a_35502_25545.n16 a_35502_25545.n171 4.5005
R44686 a_35502_25545.n18 a_35502_25545.n17 2.21666
R44687 a_35502_25545.n0 a_35502_25545.n1 0.0657695
R44688 a_35502_25545.n30 a_35502_25545.n206 4.5005
R44689 a_35502_25545.n32 a_35502_25545.n31 2.21666
R44690 a_35502_25545.n131 a_35502_25545.n205 4.5005
R44691 a_35502_25545.n132 a_35502_25545.n204 4.5005
R44692 a_35502_25545.n208 a_35502_25545.n203 4.5005
R44693 a_35502_25545.n44 a_35502_25545.n43 2.21666
R44694 a_35502_25545.n42 a_35502_25545.n181 4.5005
R44695 a_35502_25545.n180 a_35502_25545.n54 4.5005
R44696 a_35502_25545.n55 a_35502_25545.n52 2.21666
R44697 a_35502_25545.n53 a_35502_25545.n178 4.5005
R44698 a_35502_25545.n123 a_35502_25545.n122 0.0107891
R44699 a_35502_25545.n127 a_35502_25545.n158 4.5005
R44700 a_35502_25545.n21 a_35502_25545.n20 2.21666
R44701 a_35502_25545.n19 a_35502_25545.n151 4.5005
R44702 a_35502_25545.n157 a_35502_25545.n156 4.5005
R44703 a_35502_25545.n124 a_35502_25545.n166 4.5005
R44704 a_35502_25545.n24 a_35502_25545.n23 2.21666
R44705 a_35502_25545.n22 a_35502_25545.n162 4.5005
R44706 a_35502_25545.n165 a_35502_25545.n164 4.5005
R44707 a_35502_25545.n65 a_35502_25545.n67 2.21666
R44708 a_35502_25545.n64 a_35502_25545.n107 4.5005
R44709 a_35502_25545.n71 a_35502_25545.n73 2.21666
R44710 a_35502_25545.n70 a_35502_25545.n105 4.5005
R44711 a_35502_25545.n86 a_35502_25545.n88 2.21666
R44712 a_35502_25545.n215 a_35502_25545.n214 4.5005
R44713 a_35502_25545.n2 a_35502_25545.n3 2.21666
R44714 a_35502_25545.n90 a_35502_25545.n92 2.21666
R44715 a_35502_25545.n89 a_35502_25545.n102 4.5005
R44716 a_35502_25545.n160 a_35502_25545.n120 4.5005
R44717 a_35502_25545.n36 a_35502_25545.n34 2.21666
R44718 a_35502_25545.n61 a_35502_25545.n63 2.21666
R44719 a_35502_25545.n60 a_35502_25545.n106 4.5005
R44720 a_35502_25545.n75 a_35502_25545.n77 2.21666
R44721 a_35502_25545.n74 a_35502_25545.n104 4.5005
R44722 a_35502_25545.n68 a_35502_25545.n69 0.0231698
R44723 a_35502_25545.n82 a_35502_25545.n84 2.21666
R44724 a_35502_25545.n153 a_35502_25545.n81 4.5005
R44725 a_35502_25545.n121 a_35502_25545.n154 4.5005
R44726 a_35502_25545.n41 a_35502_25545.n40 2.21666
R44727 a_35502_25545.n83 a_35502_25545.n82 2.21666
R44728 a_35502_25545.n81 a_35502_25545.n103 4.5005
R44729 a_35502_25545.n38 a_35502_25545.n121 4.5005
R44730 a_35502_25545.n64 a_35502_25545.n219 4.5005
R44731 a_35502_25545.n72 a_35502_25545.n71 2.21666
R44732 a_35502_25545.n70 a_35502_25545.n218 4.5005
R44733 a_35502_25545.n87 a_35502_25545.n86 2.21666
R44734 a_35502_25545.n85 a_35502_25545.n217 4.5005
R44735 a_35502_25545.n2 a_35502_25545.n4 2.21666
R44736 a_35502_25545.n91 a_35502_25545.n90 2.21666
R44737 a_35502_25545.n89 a_35502_25545.n213 4.5005
R44738 a_35502_25545.n212 a_35502_25545.n120 4.5005
R44739 a_35502_25545.n60 a_35502_25545.n168 4.5005
R44740 a_35502_25545.n76 a_35502_25545.n75 2.21666
R44741 a_35502_25545.n74 a_35502_25545.n167 4.5005
R44742 a_35502_25545.n94 a_35502_25545.n93 0.023589
R44743 a_35502_25545.n56 a_35502_25545.n55 2.21666
R44744 a_35502_25545.n179 a_35502_25545.n54 4.5005
R44745 a_35502_25545.n42 a_35502_25545.n176 4.5005
R44746 a_35502_25545.n43 a_35502_25545.n45 2.21666
R44747 a_35502_25545.n53 a_35502_25545.n177 4.5005
R44748 a_35502_25545.n80 a_35502_25545.n78 2.21666
R44749 a_35502_25545.n193 a_35502_25545.n192 4.5005
R44750 a_35502_25545.n187 a_35502_25545.n186 4.5005
R44751 a_35502_25545.n185 a_35502_25545.n133 4.5005
R44752 a_35502_25545.n26 a_35502_25545.n173 4.5005
R44753 a_35502_25545.n29 a_35502_25545.n28 2.21666
R44754 a_35502_25545.n27 a_35502_25545.n172 4.5005
R44755 a_35502_25545.n57 a_35502_25545.n59 2.21666
R44756 a_35502_25545.n199 a_35502_25545.n198 4.5005
R44757 a_35502_25545.n47 a_35502_25545.n49 4.5005
R44758 a_35502_25545.n50 a_35502_25545.n48 2.21666
R44759 a_35502_25545.n17 a_35502_25545.n15 2.21666
R44760 a_35502_25545.n195 a_35502_25545.n16 4.5005
R44761 a_35502_25545.n209 a_35502_25545.n208 4.5005
R44762 a_35502_25545.n132 a_35502_25545.n130 4.5005
R44763 a_35502_25545.n131 a_35502_25545.n207 4.5005
R44764 a_35502_25545.n33 a_35502_25545.n31 2.21666
R44765 a_35502_25545.n30 a_35502_25545.n0 0.0743189
R44766 a_35502_25545.n299 a_35502_25545.n148 4.5005
R44767 a_35502_25545.n279 a_35502_25545.n276 4.5005
R44768 a_35502_25545.n281 a_35502_25545.n280 4.5005
R44769 a_35502_25545.n282 a_35502_25545.n275 4.5005
R44770 a_35502_25545.n284 a_35502_25545.n283 4.5005
R44771 a_35502_25545.n286 a_35502_25545.n285 4.5005
R44772 a_35502_25545.n291 a_35502_25545.n290 4.5005
R44773 a_35502_25545.n119 a_35502_25545.n292 4.5005
R44774 a_35502_25545.n293 a_35502_25545.n149 4.5005
R44775 a_35502_25545.n295 a_35502_25545.n294 4.5005
R44776 a_35502_25545.n296 a_35502_25545.n101 4.5005
R44777 a_35502_25545.n298 a_35502_25545.n297 4.5005
R44778 a_35502_25545.n302 a_35502_25545.n114 4.5005
R44779 a_35502_25545.n304 a_35502_25545.n303 4.5005
R44780 a_35502_25545.n306 a_35502_25545.n147 4.5005
R44781 a_35502_25545.n308 a_35502_25545.n307 4.5005
R44782 a_35502_25545.n309 a_35502_25545.n146 4.5005
R44783 a_35502_25545.n311 a_35502_25545.n310 4.5005
R44784 a_35502_25545.n313 a_35502_25545.n145 4.5005
R44785 a_35502_25545.n323 a_35502_25545.n322 4.5005
R44786 a_35502_25545.n118 a_35502_25545.n116 4.5005
R44787 a_35502_25545.n117 a_35502_25545.n321 4.5005
R44788 a_35502_25545.n320 a_35502_25545.n317 4.5005
R44789 a_35502_25545.n230 a_35502_25545.n222 4.5005
R44790 a_35502_25545.n112 a_35502_25545.n229 4.5005
R44791 a_35502_25545.n228 a_35502_25545.n111 4.5005
R44792 a_35502_25545.n227 a_35502_25545.n226 4.5005
R44793 a_35502_25545.n270 a_35502_25545.n269 4.5005
R44794 a_35502_25545.n268 a_35502_25545.n223 4.5005
R44795 a_35502_25545.n266 a_35502_25545.n265 4.5005
R44796 a_35502_25545.n264 a_35502_25545.n98 4.5005
R44797 a_35502_25545.n263 a_35502_25545.n100 4.5005
R44798 a_35502_25545.n99 a_35502_25545.n234 4.5005
R44799 a_35502_25545.n262 a_35502_25545.n261 4.5005
R44800 a_35502_25545.n250 a_35502_25545.n249 4.5005
R44801 a_35502_25545.n108 a_35502_25545.n251 4.5005
R44802 a_35502_25545.n252 a_35502_25545.n236 4.5005
R44803 a_35502_25545.n254 a_35502_25545.n253 4.5005
R44804 a_35502_25545.n255 a_35502_25545.n97 4.5005
R44805 a_35502_25545.n257 a_35502_25545.n256 4.5005
R44806 a_35502_25545.n258 a_35502_25545.n235 4.5005
R44807 a_35502_25545.n245 a_35502_25545.n244 4.5005
R44808 a_35502_25545.n243 a_35502_25545.n237 4.5005
R44809 a_35502_25545.n242 a_35502_25545.n241 4.5005
R44810 a_35502_25545.n240 a_35502_25545.n238 4.5005
R44811 a_35502_25545.n337 a_35502_25545.n336 4.5005
R44812 a_35502_25545.n137 a_35502_25545.n136 2.24327
R44813 a_35502_25545.n141 a_35502_25545.n139 4.5005
R44814 a_35502_25545.n142 a_35502_25545.n140 2.24296
R44815 a_35502_25545.n338 a_35502_25545.t3 3.83265
R44816 a_35502_25545.n335 a_35502_25545.t10 3.82765
R44817 a_35502_25545.n142 a_35502_25545.t14 3.82673
R44818 a_35502_25545.n332 a_35502_25545.t1 3.78255
R44819 a_35502_25545.n136 a_35502_25545.t6 3.76633
R44820 a_35502_25545.n330 a_35502_25545.t13 3.75068
R44821 a_35502_25545.n327 a_35502_25545.t0 3.75068
R44822 a_35502_25545.n329 a_35502_25545.t7 3.74975
R44823 a_35502_25545.n221 a_35502_25545.n143 3.37223
R44824 a_35502_25545.n113 a_35502_25545.n301 3.02216
R44825 a_35502_25545.n217 a_35502_25545.n216 2.89625
R44826 a_35502_25545.n18 a_35502_25545.n194 2.95081
R44827 a_35502_25545.n214 a_35502_25545.n159 2.88162
R44828 a_35502_25545.n192 a_35502_25545.n15 2.95081
R44829 a_35502_25545.n344 a_35502_25545.n342 2.76066
R44830 a_35502_25545.n344 a_35502_25545.n343 2.57313
R44831 a_35502_25545.n69 a_35502_25545.n83 2.00991
R44832 a_35502_25545.n272 a_35502_25545.n271 2.30989
R44833 a_35502_25545.n325 a_35502_25545.n144 2.30989
R44834 a_35502_25545.n301 a_35502_25545.n300 2.29659
R44835 a_35502_25545.n260 a_35502_25545.n259 2.2812
R44836 a_35502_25545.n331 a_35502_25545.n329 2.24389
R44837 a_35502_25545.n200 a_35502_25545.n170 2.23529
R44838 a_35502_25545.n182 a_35502_25545.n175 2.23529
R44839 a_35502_25545.n163 a_35502_25545.n161 2.23423
R44840 a_35502_25545.n155 a_35502_25545.n152 2.23423
R44841 a_35502_25545.n285 a_35502_25545.n273 2.18975
R44842 a_35502_25545.n324 a_35502_25545.n145 2.18975
R44843 a_35502_25545.n271 a_35502_25545.n222 2.16725
R44844 a_35502_25545.n250 a_35502_25545.n144 2.16725
R44845 a_35502_25545.n221 a_35502_25545.n220 2.11247
R44846 a_35502_25545.n186 a_35502_25545.n150 2.102
R44847 a_35502_25545.n46 a_35502_25545.n209 2.102
R44848 a_35502_25545.n341 a_35502_25545.n333 2.07395
R44849 a_35502_25545.n220 a_35502_25545.n150 2.07182
R44850 a_35502_25545.n210 a_35502_25545.n46 2.07182
R44851 a_35502_25545.n37 a_35502_25545.n66 2.13751
R44852 a_35502_25545.n211 a_35502_25545.n62 2.13751
R44853 a_35502_25545.n342 a_35502_25545.n341 1.90955
R44854 a_35502_25545.n353 a_35502_25545.n352 1.71486
R44855 a_35502_25545.n210 a_35502_25545.n143 1.50911
R44856 a_35502_25545.n220 a_35502_25545.n37 1.5005
R44857 a_35502_25545.n211 a_35502_25545.n210 1.5005
R44858 a_35502_25545.n273 a_35502_25545.n272 1.5005
R44859 a_35502_25545.n325 a_35502_25545.n324 1.5005
R44860 a_35502_25545.n341 a_35502_25545.n340 1.5005
R44861 a_35502_25545.n352 a_35502_25545.n351 1.5005
R44862 a_35502_25545.n348 a_35502_25545.n347 1.5005
R44863 a_35502_25545.t10 a_35502_25545.t15 1.4705
R44864 a_35502_25545.t13 a_35502_25545.t18 1.4705
R44865 a_35502_25545.t1 a_35502_25545.t9 1.4705
R44866 a_35502_25545.t0 a_35502_25545.t16 1.4705
R44867 a_35502_25545.n279 a_35502_25545.n278 1.39514
R44868 a_35502_25545.n272 a_35502_25545.n221 1.39023
R44869 a_35502_25545.n326 a_35502_25545.n325 1.39023
R44870 a_35502_25545.n328 a_35502_25545.n327 1.27228
R44871 a_35502_25545.n314 a_35502_25545.n313 1.26997
R44872 a_35502_25545.n287 a_35502_25545.n286 1.26997
R44873 a_35502_25545.n322 a_35502_25545.n316 1.24392
R44874 a_35502_25545.n290 a_35502_25545.n289 1.24392
R44875 a_35502_25545.n249 a_35502_25545.n248 1.24204
R44876 a_35502_25545.n231 a_35502_25545.n230 1.24204
R44877 a_35502_25545.n331 a_35502_25545.n330 1.20682
R44878 a_35502_25545.n246 a_35502_25545.n245 1.20414
R44879 a_35502_25545.n269 a_35502_25545.n233 1.20414
R44880 a_35502_25545.n320 a_35502_25545.n319 1.14132
R44881 a_35502_25545.n332 a_35502_25545.n140 1.20835
R44882 a_35502_25545.n227 a_35502_25545.n224 1.13598
R44883 a_35502_25545.n339 a_35502_25545.n335 1.13573
R44884 a_35502_25545.n346 a_35502_25545.n345 0.90675
R44885 a_35502_25545.n350 a_35502_25545.n349 0.90675
R44886 a_35502_25545.n335 a_35502_25545.n135 0.939226
R44887 a_35502_25545.n291 a_35502_25545.n273 0.752
R44888 a_35502_25545.n324 a_35502_25545.n323 0.752
R44889 a_35502_25545.n271 a_35502_25545.n270 0.71825
R44890 a_35502_25545.n244 a_35502_25545.n144 0.71825
R44891 a_35502_25545.n315 a_35502_25545.n314 0.663658
R44892 a_35502_25545.n316 a_35502_25545.n315 0.663658
R44893 a_35502_25545.n288 a_35502_25545.n287 0.663658
R44894 a_35502_25545.n289 a_35502_25545.n288 0.663658
R44895 a_35502_25545.n247 a_35502_25545.n246 0.655156
R44896 a_35502_25545.n248 a_35502_25545.n247 0.655156
R44897 a_35502_25545.n233 a_35502_25545.n232 0.655156
R44898 a_35502_25545.n232 a_35502_25545.n231 0.655156
R44899 a_35502_25545.n326 a_35502_25545.n143 0.603852
R44900 a_35502_25545.n333 a_35502_25545.n332 0.596867
R44901 a_35502_25545.n96 a_35502_25545.n95 0.313126
R44902 a_35502_25545.n278 a_35502_25545.n277 0.432797
R44903 a_35502_25545.n304 a_35502_25545.n114 0.394842
R44904 a_35502_25545.n299 a_35502_25545.n298 0.394842
R44905 a_35502_25545.n117 a_35502_25545.n317 0.381816
R44906 a_35502_25545.n294 a_35502_25545.n293 0.381816
R44907 a_35502_25545.n241 a_35502_25545.n240 0.379447
R44908 a_35502_25545.n258 a_35502_25545.n257 0.379447
R44909 a_35502_25545.n253 a_35502_25545.n252 0.379447
R44910 a_35502_25545.n266 a_35502_25545.n98 0.379447
R44911 a_35502_25545.n99 a_35502_25545.n262 0.379447
R44912 a_35502_25545.n226 a_35502_25545.n111 0.379447
R44913 a_35502_25545.n178 a_35502_25545.n52 0.44431
R44914 a_35502_25545.n79 a_35502_25545.n191 0.44431
R44915 a_35502_25545.n58 a_35502_25545.n171 0.44431
R44916 a_35502_25545.n1 a_35502_25545.n206 1.94004
R44917 a_35502_25545.n88 a_35502_25545.n105 0.44431
R44918 a_35502_25545.n94 a_35502_25545.n104 1.95665
R44919 a_35502_25545.n56 a_35502_25545.n177 0.44431
R44920 a_35502_25545.n80 a_35502_25545.n172 0.44431
R44921 a_35502_25545.n59 a_35502_25545.n195 0.44431
R44922 a_35502_25545.n297 a_35502_25545.n148 0.375125
R44923 a_35502_25545.n303 a_35502_25545.n302 0.375125
R44924 a_35502_25545.n190 a_35502_25545.n25 0.431935
R44925 a_35502_25545.n32 a_35502_25545.n205 0.431935
R44926 a_35502_25545.n73 a_35502_25545.n107 0.431935
R44927 a_35502_25545.n77 a_35502_25545.n106 0.431935
R44928 a_35502_25545.n29 a_35502_25545.n173 0.431935
R44929 a_35502_25545.n207 a_35502_25545.n33 0.431935
R44930 a_35502_25545.n295 a_35502_25545.n149 0.36275
R44931 a_35502_25545.n321 a_35502_25545.n320 0.36275
R44932 a_35502_25545.n183 a_35502_25545.n174 0.3605
R44933 a_35502_25545.n201 a_35502_25545.n169 0.3605
R44934 a_35502_25545.n156 a_35502_25545.n151 0.3605
R44935 a_35502_25545.n164 a_35502_25545.n162 0.3605
R44936 a_35502_25545.n38 a_35502_25545.n103 0.3605
R44937 a_35502_25545.n219 a_35502_25545.n72 0.429685
R44938 a_35502_25545.n218 a_35502_25545.n87 0.429685
R44939 a_35502_25545.n213 a_35502_25545.n212 0.3605
R44940 a_35502_25545.n168 a_35502_25545.n76 0.429685
R44941 a_35502_25545.n167 a_35502_25545.n94 1.93517
R44942 a_35502_25545.n228 a_35502_25545.n227 0.3605
R44943 a_35502_25545.n265 a_35502_25545.n264 0.3605
R44944 a_35502_25545.n261 a_35502_25545.n234 0.3605
R44945 a_35502_25545.n256 a_35502_25545.n235 0.3605
R44946 a_35502_25545.n254 a_35502_25545.n236 0.3605
R44947 a_35502_25545.n242 a_35502_25545.n238 0.3605
R44948 a_35502_25545.n333 a_35502_25545.n328 0.339591
R44949 a_35502_25545.n319 a_35502_25545.n318 0.335806
R44950 a_35502_25545.n225 a_35502_25545.n224 0.33475
R44951 a_35502_25545.n347 a_35502_25545.n346 0.320048
R44952 a_35502_25545.n351 a_35502_25545.n350 0.320048
R44953 a_35502_25545.n307 a_35502_25545.n146 0.302474
R44954 a_35502_25545.n282 a_35502_25545.n281 0.302474
R44955 a_35502_25545.n181 a_35502_25545.n180 0.287375
R44956 a_35502_25545.n197 a_35502_25545.n196 0.287375
R44957 a_35502_25545.n154 a_35502_25545.n153 0.287375
R44958 a_35502_25545.n160 a_35502_25545.n102 0.287375
R44959 a_35502_25545.n179 a_35502_25545.n176 0.287375
R44960 a_35502_25545.n47 a_35502_25545.n199 0.287375
R44961 a_35502_25545.n280 a_35502_25545.n275 0.287375
R44962 a_35502_25545.n309 a_35502_25545.n308 0.287375
R44963 a_35502_25545.n348 a_35502_25545.n344 0.212426
R44964 a_35502_25545.n156 a_35502_25545.n155 0.208888
R44965 a_35502_25545.n164 a_35502_25545.n161 0.208888
R44966 a_35502_25545.n183 a_35502_25545.n182 0.20887
R44967 a_35502_25545.n201 a_35502_25545.n200 0.20887
R44968 a_35502_25545.n139 a_35502_25545.n331 0.208385
R44969 a_35502_25545.n301 a_35502_25545.n148 0.208099
R44970 a_35502_25545.n260 a_35502_25545.n235 0.208099
R44971 a_35502_25545.n245 a_35502_25545.n237 0.147342
R44972 a_35502_25545.n257 a_35502_25545.n97 0.147342
R44973 a_35502_25545.n252 a_35502_25545.n108 0.147342
R44974 a_35502_25545.n269 a_35502_25545.n268 0.147342
R44975 a_35502_25545.n100 a_35502_25545.n98 0.147342
R44976 a_35502_25545.n112 a_35502_25545.n111 0.147342
R44977 a_35502_25545.n307 a_35502_25545.n306 0.147342
R44978 a_35502_25545.n311 a_35502_25545.n146 0.147342
R44979 a_35502_25545.n118 a_35502_25545.n117 0.147342
R44980 a_35502_25545.n281 a_35502_25545.n276 0.147342
R44981 a_35502_25545.n283 a_35502_25545.n282 0.147342
R44982 a_35502_25545.n293 a_35502_25545.n119 0.147342
R44983 a_35502_25545.n298 a_35502_25545.n101 0.147342
R44984 a_35502_25545.n180 a_35502_25545.n52 0.209185
R44985 a_35502_25545.n181 a_35502_25545.n44 0.209185
R44986 a_35502_25545.n182 a_35502_25545.n44 0.825446
R44987 a_35502_25545.n12 a_35502_25545.n174 0.209185
R44988 a_35502_25545.n7 a_35502_25545.n12 0.565419
R44989 a_35502_25545.n188 a_35502_25545.n7 0.834884
R44990 a_35502_25545.n189 a_35502_25545.n188 0.14
R44991 a_35502_25545.n190 a_35502_25545.n189 0.14
R44992 a_35502_25545.n191 a_35502_25545.n25 0.209185
R44993 a_35502_25545.n194 a_35502_25545.n79 0.209185
R44994 a_35502_25545.n18 a_35502_25545.n171 0.209185
R44995 a_35502_25545.n197 a_35502_25545.n58 0.209185
R44996 a_35502_25545.n196 a_35502_25545.n51 0.209185
R44997 a_35502_25545.n200 a_35502_25545.n51 0.825446
R44998 a_35502_25545.n14 a_35502_25545.n169 0.209185
R44999 a_35502_25545.n10 a_35502_25545.n14 0.565419
R45000 a_35502_25545.n203 a_35502_25545.n10 0.834884
R45001 a_35502_25545.n204 a_35502_25545.n203 0.14
R45002 a_35502_25545.n205 a_35502_25545.n204 0.14
R45003 a_35502_25545.n206 a_35502_25545.n32 0.209185
R45004 a_35502_25545.n153 a_35502_25545.n84 0.209185
R45005 a_35502_25545.n154 a_35502_25545.n41 0.209185
R45006 a_35502_25545.n155 a_35502_25545.n41 0.825427
R45007 a_35502_25545.n21 a_35502_25545.n151 0.209185
R45008 a_35502_25545.n158 a_35502_25545.n21 0.429685
R45009 a_35502_25545.n158 a_35502_25545.n129 0.208907
R45010 a_35502_25545.n67 a_35502_25545.n129 0.836657
R45011 a_35502_25545.n67 a_35502_25545.n107 0.209185
R45012 a_35502_25545.n73 a_35502_25545.n105 0.209185
R45013 a_35502_25545.n88 a_35502_25545.n159 0.209185
R45014 a_35502_25545.n214 a_35502_25545.n3 0.209185
R45015 a_35502_25545.n3 a_35502_25545.n92 0.513496
R45016 a_35502_25545.n92 a_35502_25545.n102 0.209185
R45017 a_35502_25545.n36 a_35502_25545.n160 0.209185
R45018 a_35502_25545.n36 a_35502_25545.n161 0.825427
R45019 a_35502_25545.n24 a_35502_25545.n162 0.209185
R45020 a_35502_25545.n166 a_35502_25545.n24 0.429685
R45021 a_35502_25545.n166 a_35502_25545.n126 0.208907
R45022 a_35502_25545.n63 a_35502_25545.n126 0.836657
R45023 a_35502_25545.n63 a_35502_25545.n106 0.209185
R45024 a_35502_25545.n77 a_35502_25545.n104 0.209185
R45025 a_35502_25545.n83 a_35502_25545.n103 0.209185
R45026 a_35502_25545.n39 a_35502_25545.n38 0.209137
R45027 a_35502_25545.n39 a_35502_25545.n37 0.886485
R45028 a_35502_25545.n219 a_35502_25545.n66 0.209113
R45029 a_35502_25545.n218 a_35502_25545.n72 0.209185
R45030 a_35502_25545.n217 a_35502_25545.n87 0.209185
R45031 a_35502_25545.n216 a_35502_25545.n4 0.209185
R45032 a_35502_25545.n91 a_35502_25545.n4 0.498871
R45033 a_35502_25545.n213 a_35502_25545.n91 0.209185
R45034 a_35502_25545.n212 a_35502_25545.n35 0.209137
R45035 a_35502_25545.n211 a_35502_25545.n35 0.886485
R45036 a_35502_25545.n168 a_35502_25545.n62 0.209113
R45037 a_35502_25545.n167 a_35502_25545.n76 0.209185
R45038 a_35502_25545.n56 a_35502_25545.n179 0.209185
R45039 a_35502_25545.n45 a_35502_25545.n176 0.209185
R45040 a_35502_25545.n150 a_35502_25545.n45 0.908935
R45041 a_35502_25545.n186 a_35502_25545.n185 0.14
R45042 a_35502_25545.n185 a_35502_25545.n173 0.14
R45043 a_35502_25545.n29 a_35502_25545.n172 0.209185
R45044 a_35502_25545.n192 a_35502_25545.n80 0.209185
R45045 a_35502_25545.n195 a_35502_25545.n15 0.209185
R45046 a_35502_25545.n199 a_35502_25545.n59 0.209185
R45047 a_35502_25545.n48 a_35502_25545.n47 0.209185
R45048 a_35502_25545.n48 a_35502_25545.n46 0.908935
R45049 a_35502_25545.n209 a_35502_25545.n130 0.14
R45050 a_35502_25545.n207 a_35502_25545.n130 0.14
R45051 a_35502_25545.n33 a_35502_25545.n0 1.54288
R45052 a_35502_25545.n280 a_35502_25545.n279 0.14
R45053 a_35502_25545.n284 a_35502_25545.n275 0.14
R45054 a_35502_25545.n285 a_35502_25545.n284 0.14
R45055 a_35502_25545.n292 a_35502_25545.n291 0.14
R45056 a_35502_25545.n292 a_35502_25545.n149 0.14
R45057 a_35502_25545.n296 a_35502_25545.n295 0.14
R45058 a_35502_25545.n297 a_35502_25545.n296 0.14
R45059 a_35502_25545.n302 a_35502_25545.n113 0.208168
R45060 a_35502_25545.n303 a_35502_25545.n147 0.14
R45061 a_35502_25545.n308 a_35502_25545.n147 0.14
R45062 a_35502_25545.n310 a_35502_25545.n309 0.14
R45063 a_35502_25545.n310 a_35502_25545.n145 0.14
R45064 a_35502_25545.n323 a_35502_25545.n116 0.14
R45065 a_35502_25545.n321 a_35502_25545.n116 0.14
R45066 a_35502_25545.n229 a_35502_25545.n228 0.14
R45067 a_35502_25545.n229 a_35502_25545.n222 0.14
R45068 a_35502_25545.n270 a_35502_25545.n223 0.14
R45069 a_35502_25545.n265 a_35502_25545.n223 0.14
R45070 a_35502_25545.n264 a_35502_25545.n263 0.14
R45071 a_35502_25545.n263 a_35502_25545.n234 0.14
R45072 a_35502_25545.n261 a_35502_25545.n110 0.208168
R45073 a_35502_25545.n110 a_35502_25545.n260 3.03679
R45074 a_35502_25545.n256 a_35502_25545.n255 0.14
R45075 a_35502_25545.n255 a_35502_25545.n254 0.14
R45076 a_35502_25545.n251 a_35502_25545.n236 0.14
R45077 a_35502_25545.n251 a_35502_25545.n250 0.14
R45078 a_35502_25545.n244 a_35502_25545.n243 0.14
R45079 a_35502_25545.n243 a_35502_25545.n242 0.14
R45080 a_35502_25545.n96 a_35502_25545.n238 1.12911
R45081 a_35502_25545.n137 a_35502_25545.n138 1.2061
R45082 a_35502_25545.n336 a_35502_25545.n137 0.230885
R45083 a_35502_25545.n336 a_35502_25545.n334 0.14
R45084 a_35502_25545.n134 a_35502_25545.n135 1.27228
R45085 a_35502_25545.t11 a_35502_25545.n134 6.50385
R45086 a_35502_25545.n140 a_35502_25545.n139 0.230894
R45087 a_35502_25545.n142 a_35502_25545.n141 0.138586
R45088 a_35502_25545.n337 a_35502_25545.n136 0.137318
R45089 a_35502_25545.n226 a_35502_25545.n225 0.128395
R45090 a_35502_25545.n318 a_35502_25545.n317 0.128395
R45091 a_35502_25545.n241 a_35502_25545.n239 0.118921
R45092 a_35502_25545.n259 a_35502_25545.n258 0.118921
R45093 a_35502_25545.n267 a_35502_25545.n266 0.118921
R45094 a_35502_25545.n313 a_35502_25545.n312 0.114184
R45095 a_35502_25545.n286 a_35502_25545.n274 0.114184
R45096 a_35502_25545.n305 a_35502_25545.n304 0.113
R45097 a_35502_25545.n338 a_35502_25545.n337 0.110782
R45098 a_35502_25545.n141 a_35502_25545.n329 0.109514
R45099 a_35502_25545.n13 a_35502_25545.n202 0.109179
R45100 a_35502_25545.n11 a_35502_25545.n184 0.109179
R45101 a_35502_25545.n57 a_35502_25545.n16 0.107155
R45102 a_35502_25545.n78 a_35502_25545.n27 0.107155
R45103 a_35502_25545.n55 a_35502_25545.n53 0.107155
R45104 a_35502_25545.n352 a_35502_25545.n348 0.105095
R45105 a_35502_25545.n131 a_35502_25545.n31 0.103632
R45106 a_35502_25545.n28 a_35502_25545.n26 0.103632
R45107 a_35502_25545.n300 a_35502_25545.n299 0.103526
R45108 a_35502_25545.n22 a_35502_25545.n165 0.102991
R45109 a_35502_25545.n124 a_35502_25545.n23 0.102991
R45110 a_35502_25545.n19 a_35502_25545.n157 0.102991
R45111 a_35502_25545.n127 a_35502_25545.n20 0.102991
R45112 a_35502_25545.n340 a_35502_25545.n339 0.0995
R45113 a_35502_25545.n75 a_35502_25545.n60 0.0933826
R45114 a_35502_25545.n71 a_35502_25545.n64 0.0933826
R45115 a_35502_25545.n93 a_35502_25545.n74 0.092742
R45116 a_35502_25545.n90 a_35502_25545.n2 0.092742
R45117 a_35502_25545.n86 a_35502_25545.n70 0.092742
R45118 a_35502_25545.n82 a_35502_25545.n68 0.092742
R45119 a_35502_25545.n198 a_35502_25545.n49 0.0821726
R45120 a_35502_25545.n42 a_35502_25545.n54 0.0821726
R45121 a_35502_25545.n120 a_35502_25545.n89 0.0821726
R45122 a_35502_25545.n121 a_35502_25545.n81 0.0821726
R45123 a_35502_25545.n128 a_35502_25545.n127 0.0427776
R45124 a_35502_25545.n125 a_35502_25545.n124 0.0427776
R45125 a_35502_25545.n340 a_35502_25545.n334 0.041
R45126 a_35502_25545.n132 a_35502_25545.n131 0.0402153
R45127 a_35502_25545.n26 a_35502_25545.n133 0.0402153
R45128 a_35502_25545.n53 a_35502_25545.n122 0.0402153
R45129 a_35502_25545.n187 a_35502_25545.n133 0.0402153
R45130 a_35502_25545.n208 a_35502_25545.n132 0.0402153
R45131 a_35502_25545.n306 a_35502_25545.n305 0.0348421
R45132 a_35502_25545.n277 a_35502_25545.n276 0.0348421
R45133 a_35502_25545.n202 a_35502_25545.n170 0.0344623
R45134 a_35502_25545.n184 a_35502_25545.n175 0.0344623
R45135 a_35502_25545.n312 a_35502_25545.n311 0.0336579
R45136 a_35502_25545.n283 a_35502_25545.n274 0.0336579
R45137 a_35502_25545.n165 a_35502_25545.n163 0.0325285
R45138 a_35502_25545.n157 a_35502_25545.n152 0.0325285
R45139 a_35502_25545.n239 a_35502_25545.n237 0.0289211
R45140 a_35502_25545.n268 a_35502_25545.n267 0.0289211
R45141 a_35502_25545.n240 a_35502_25545.n95 0.166289
R45142 a_35502_25545.n115 a_35502_25545.n114 0.156816
R45143 a_35502_25545.n262 a_35502_25545.n109 0.156816
R45144 a_35502_25545.n9 a_35502_25545.n8 0.154009
R45145 a_35502_25545.n6 a_35502_25545.n5 0.154009
R45146 a_35502_25545.n290 a_35502_25545.n119 0.147342
R45147 a_35502_25545.n322 a_35502_25545.n118 0.147342
R45148 a_35502_25545.n230 a_35502_25545.n112 0.147342
R45149 a_35502_25545.n249 a_35502_25545.n108 0.147342
R45150 a_35502_25545.n294 a_35502_25545.n101 0.147342
R45151 a_35502_25545.n100 a_35502_25545.n99 0.147342
R45152 a_35502_25545.n253 a_35502_25545.n97 0.147342
R45153 a_35502_25545.n90 a_35502_25545.n89 0.0943434
R45154 a_35502_25545.n82 a_35502_25545.n81 0.0943434
R45155 a_35502_25545.n75 a_35502_25545.n74 0.0901797
R45156 a_35502_25545.n71 a_35502_25545.n70 0.0901797
R45157 a_35502_25545.n8 a_35502_25545.n13 0.0847264
R45158 a_35502_25545.n5 a_35502_25545.n11 0.0847264
R45159 a_35502_25545.n86 a_35502_25545.n85 0.0799306
R45160 a_35502_25545.n193 a_35502_25545.n78 0.0799306
R45161 a_35502_25545.n65 a_35502_25545.n64 0.0799306
R45162 a_35502_25545.n61 a_35502_25545.n60 0.0799306
R45163 a_35502_25545.n198 a_35502_25545.n57 0.0799306
R45164 a_35502_25545.n55 a_35502_25545.n54 0.0799306
R45165 a_35502_25545.n50 a_35502_25545.n49 0.0799306
R45166 a_35502_25545.n43 a_35502_25545.n42 0.0799306
R45167 a_35502_25545.n121 a_35502_25545.n40 0.0799306
R45168 a_35502_25545.n120 a_35502_25545.n34 0.0799306
R45169 a_35502_25545.n31 a_35502_25545.n30 0.0799306
R45170 a_35502_25545.n28 a_35502_25545.n27 0.0799306
R45171 a_35502_25545.n23 a_35502_25545.n22 0.0799306
R45172 a_35502_25545.n20 a_35502_25545.n19 0.0799306
R45173 a_35502_25545.n17 a_35502_25545.n16 0.0799306
R45174 a_35502_25545.n215 a_35502_25545.n2 0.0799306
R45175 a_35502_25545.n1 a_35502_25545.t50 8.08727
R45176 a_33249_35053.n109 a_33249_35053.n106 9.23995
R45177 a_33249_35053.n35 a_33249_35053.n33 7.94229
R45178 a_33249_35053.n80 a_33249_35053.n77 7.94229
R45179 a_33249_35053.n108 a_33249_35053.t103 6.72766
R45180 a_33249_35053.n129 a_33249_35053.n127 6.58329
R45181 a_33249_35053.n106 a_33249_35053.n14 6.01251
R45182 a_33249_35053.n126 a_33249_35053.t130 5.85326
R45183 a_33249_35053.n130 a_33249_35053.t117 5.85326
R45184 a_33249_35053.n126 a_33249_35053.n125 5.84661
R45185 a_33249_35053.n32 a_33249_35053.t50 5.69423
R45186 a_33249_35053.n36 a_33249_35053.t60 5.69423
R45187 a_33249_35053.n79 a_33249_35053.t57 5.69423
R45188 a_33249_35053.n75 a_33249_35053.t63 5.69423
R45189 a_33249_35053.n32 a_33249_35053.n31 5.49558
R45190 a_33249_35053.n79 a_33249_35053.n78 5.49558
R45191 a_33249_35053.n157 a_33249_35053.n0 4.58971
R45192 a_33249_35053.n1 a_33249_35053.t126 5.84971
R45193 a_33249_35053.n2 a_33249_35053.n132 4.58971
R45194 a_33249_35053.n3 a_33249_35053.n103 4.22068
R45195 a_33249_35053.n4 a_33249_35053.t64 5.69068
R45196 a_33249_35053.n5 a_33249_35053.n102 4.22068
R45197 a_33249_35053.n6 a_33249_35053.n72 4.22068
R45198 a_33249_35053.t61 a_33249_35053.n7 5.69068
R45199 a_33249_35053.n71 a_33249_35053.n8 4.22068
R45200 a_33249_35053.n9 a_33249_35053.t104 5.47076
R45201 a_33249_35053.n129 a_33249_35053.n128 4.59326
R45202 a_33249_35053.n109 a_33249_35053.n108 4.52463
R45203 a_33249_35053.n110 a_33249_35053.t97 4.41563
R45204 a_33249_35053.n119 a_33249_35053.t88 4.41563
R45205 a_33249_35053.n35 a_33249_35053.n34 4.22423
R45206 a_33249_35053.n77 a_33249_35053.n76 4.22423
R45207 a_33249_35053.n108 a_33249_35053.n107 4.21432
R45208 a_33249_35053.n150 a_33249_35053.t139 4.21195
R45209 a_33249_35053.n152 a_33249_35053.t134 4.21195
R45210 a_33249_35053.n137 a_33249_35053.t123 4.21195
R45211 a_33249_35053.n135 a_33249_35053.t115 4.21195
R45212 a_33249_35053.n42 a_33249_35053.t29 4.05054
R45213 a_33249_35053.n47 a_33249_35053.t7 4.05054
R45214 a_33249_35053.n49 a_33249_35053.t38 4.05054
R45215 a_33249_35053.n56 a_33249_35053.t42 4.05054
R45216 a_33249_35053.n58 a_33249_35053.t32 4.05054
R45217 a_33249_35053.n64 a_33249_35053.t36 4.05054
R45218 a_33249_35053.n66 a_33249_35053.t68 4.05054
R45219 a_33249_35053.n37 a_33249_35053.t84 4.05054
R45220 a_33249_35053.n21 a_33249_35053.t33 4.05054
R45221 a_33249_35053.n26 a_33249_35053.t18 4.05054
R45222 a_33249_35053.n28 a_33249_35053.t52 4.05054
R45223 a_33249_35053.n88 a_33249_35053.t58 4.05054
R45224 a_33249_35053.n90 a_33249_35053.t41 4.05054
R45225 a_33249_35053.n96 a_33249_35053.t46 4.05054
R45226 a_33249_35053.n98 a_33249_35053.t78 4.05054
R45227 a_33249_35053.n16 a_33249_35053.t3 4.05054
R45228 a_33249_35053.n150 a_33249_35053.t106 4.03668
R45229 a_33249_35053.n152 a_33249_35053.t137 4.03668
R45230 a_33249_35053.n137 a_33249_35053.t124 4.03668
R45231 a_33249_35053.n135 a_33249_35053.t120 4.03668
R45232 a_33249_35053.n42 a_33249_35053.t31 3.87765
R45233 a_33249_35053.n47 a_33249_35053.t12 3.87765
R45234 a_33249_35053.n49 a_33249_35053.t47 3.87765
R45235 a_33249_35053.n56 a_33249_35053.t51 3.87765
R45236 a_33249_35053.n58 a_33249_35053.t37 3.87765
R45237 a_33249_35053.n64 a_33249_35053.t40 3.87765
R45238 a_33249_35053.n66 a_33249_35053.t72 3.87765
R45239 a_33249_35053.n37 a_33249_35053.t1 3.87765
R45240 a_33249_35053.n21 a_33249_35053.t35 3.87765
R45241 a_33249_35053.n26 a_33249_35053.t20 3.87765
R45242 a_33249_35053.n28 a_33249_35053.t55 3.87765
R45243 a_33249_35053.n88 a_33249_35053.t59 3.87765
R45244 a_33249_35053.n90 a_33249_35053.t43 3.87765
R45245 a_33249_35053.n96 a_33249_35053.t48 3.87765
R45246 a_33249_35053.n98 a_33249_35053.t79 3.87765
R45247 a_33249_35053.n16 a_33249_35053.t4 3.87765
R45248 a_33249_35053.n110 a_33249_35053.t93 3.833
R45249 a_33249_35053.n119 a_33249_35053.t94 3.833
R45250 a_33249_35053.n146 a_33249_35053.n142 3.81703
R45251 a_33249_35053.n133 a_33249_35053.n2 3.95161
R45252 a_33249_35053.n118 a_33249_35053.n114 3.80578
R45253 a_33249_35053.n123 a_33249_35053.n9 3.90344
R45254 a_33249_35053.n124 a_33249_35053.n10 3.69568
R45255 a_33249_35053.n69 a_33249_35053.n36 3.25667
R45256 a_33249_35053.n113 a_33249_35053.n111 3.15563
R45257 a_33249_35053.n117 a_33249_35053.n115 3.15563
R45258 a_33249_35053.n8 a_33249_35053.n70 3.15553
R45259 a_33249_35053.n105 a_33249_35053.n5 3.15553
R45260 a_33249_35053.n149 a_33249_35053.n148 2.95195
R45261 a_33249_35053.n145 a_33249_35053.n144 2.95195
R45262 a_33249_35053.n141 a_33249_35053.n140 2.95195
R45263 a_33249_35053.n13 a_33249_35053.n12 2.95195
R45264 a_33249_35053.n149 a_33249_35053.n147 2.77668
R45265 a_33249_35053.n145 a_33249_35053.n143 2.77668
R45266 a_33249_35053.n141 a_33249_35053.n139 2.77668
R45267 a_33249_35053.n13 a_33249_35053.n11 2.77668
R45268 a_33249_35053.n41 a_33249_35053.n37 2.73714
R45269 a_33249_35053.n20 a_33249_35053.n16 2.73714
R45270 a_33249_35053.n46 a_33249_35053.n42 2.73672
R45271 a_33249_35053.n25 a_33249_35053.n21 2.73672
R45272 a_33249_35053.n151 a_33249_35053.n149 2.71872
R45273 a_33249_35053.n114 a_33249_35053.n110 2.71872
R45274 a_33249_35053.n59 a_33249_35053.n57 2.60203
R45275 a_33249_35053.n91 a_33249_35053.n89 2.60203
R45276 a_33249_35053.n131 a_33249_35053.n124 2.5825
R45277 a_33249_35053.n45 a_33249_35053.n44 2.58054
R45278 a_33249_35053.n54 a_33249_35053.n53 2.58054
R45279 a_33249_35053.n62 a_33249_35053.n61 2.58054
R45280 a_33249_35053.n40 a_33249_35053.n39 2.58054
R45281 a_33249_35053.n24 a_33249_35053.n23 2.58054
R45282 a_33249_35053.n86 a_33249_35053.n85 2.58054
R45283 a_33249_35053.n94 a_33249_35053.n93 2.58054
R45284 a_33249_35053.n19 a_33249_35053.n18 2.58054
R45285 a_33249_35053.n113 a_33249_35053.n112 2.573
R45286 a_33249_35053.n117 a_33249_35053.n116 2.573
R45287 a_33249_35053.n138 a_33249_35053.n136 2.56118
R45288 a_33249_35053.n153 a_33249_35053.n151 2.56118
R45289 a_33249_35053.n131 a_33249_35053.n130 2.54573
R45290 a_33249_35053.n67 a_33249_35053.n65 2.53418
R45291 a_33249_35053.n50 a_33249_35053.n48 2.53418
R45292 a_33249_35053.n99 a_33249_35053.n97 2.53418
R45293 a_33249_35053.n29 a_33249_35053.n27 2.53418
R45294 a_33249_35053.n75 a_33249_35053.n15 2.51873
R45295 a_33249_35053.n45 a_33249_35053.n43 2.40765
R45296 a_33249_35053.n54 a_33249_35053.n52 2.40765
R45297 a_33249_35053.n62 a_33249_35053.n60 2.40765
R45298 a_33249_35053.n40 a_33249_35053.n38 2.40765
R45299 a_33249_35053.n24 a_33249_35053.n22 2.40765
R45300 a_33249_35053.n86 a_33249_35053.n84 2.40765
R45301 a_33249_35053.n94 a_33249_35053.n92 2.40765
R45302 a_33249_35053.n19 a_33249_35053.n17 2.40765
R45303 a_33249_35053.n156 a_33249_35053.n155 2.27857
R45304 a_33249_35053.n33 a_33249_35053.n30 2.23844
R45305 a_33249_35053.n134 a_33249_35053.n13 2.00466
R45306 a_33249_35053.n121 a_33249_35053.n120 1.67718
R45307 a_33249_35053.n0 a_33249_35053.n156 1.67353
R45308 a_33249_35053.n73 a_33249_35053.n6 1.65553
R45309 a_33249_35053.n104 a_33249_35053.n3 1.65553
R45310 a_33249_35053.n101 a_33249_35053.n100 1.5005
R45311 a_33249_35053.n69 a_33249_35053.n68 1.5005
R45312 a_33249_35053.n104 a_33249_35053.n14 1.5005
R45313 a_33249_35053.n83 a_33249_35053.n82 1.5005
R45314 a_33249_35053.n81 a_33249_35053.n80 1.5005
R45315 a_33249_35053.n74 a_33249_35053.n73 1.5005
R45316 a_33249_35053.n51 a_33249_35053.n30 1.5005
R45317 a_33249_35053.n134 a_33249_35053.n133 1.5005
R45318 a_33249_35053.n155 a_33249_35053.n154 1.5005
R45319 a_33249_35053.n127 a_33249_35053.n10 1.5005
R45320 a_33249_35053.n103 a_33249_35053.t67 1.4705
R45321 a_33249_35053.n103 a_33249_35053.t9 1.4705
R45322 a_33249_35053.n102 a_33249_35053.t73 1.4705
R45323 a_33249_35053.n102 a_33249_35053.t17 1.4705
R45324 a_33249_35053.n31 a_33249_35053.t77 1.4705
R45325 a_33249_35053.n31 a_33249_35053.t28 1.4705
R45326 a_33249_35053.n34 a_33249_35053.t87 1.4705
R45327 a_33249_35053.n34 a_33249_35053.t45 1.4705
R45328 a_33249_35053.n43 a_33249_35053.t70 1.4705
R45329 a_33249_35053.n43 a_33249_35053.t13 1.4705
R45330 a_33249_35053.n44 a_33249_35053.t66 1.4705
R45331 a_33249_35053.n44 a_33249_35053.t8 1.4705
R45332 a_33249_35053.n52 a_33249_35053.t76 1.4705
R45333 a_33249_35053.n52 a_33249_35053.t22 1.4705
R45334 a_33249_35053.n53 a_33249_35053.t69 1.4705
R45335 a_33249_35053.n53 a_33249_35053.t11 1.4705
R45336 a_33249_35053.n60 a_33249_35053.t80 1.4705
R45337 a_33249_35053.n60 a_33249_35053.t10 1.4705
R45338 a_33249_35053.n61 a_33249_35053.t71 1.4705
R45339 a_33249_35053.n61 a_33249_35053.t5 1.4705
R45340 a_33249_35053.n38 a_33249_35053.t23 1.4705
R45341 a_33249_35053.n38 a_33249_35053.t49 1.4705
R45342 a_33249_35053.n39 a_33249_35053.t14 1.4705
R45343 a_33249_35053.n39 a_33249_35053.t39 1.4705
R45344 a_33249_35053.n72 a_33249_35053.t62 1.4705
R45345 a_33249_35053.n72 a_33249_35053.t0 1.4705
R45346 a_33249_35053.n71 a_33249_35053.t65 1.4705
R45347 a_33249_35053.n71 a_33249_35053.t6 1.4705
R45348 a_33249_35053.n78 a_33249_35053.t83 1.4705
R45349 a_33249_35053.n78 a_33249_35053.t30 1.4705
R45350 a_33249_35053.n76 a_33249_35053.t2 1.4705
R45351 a_33249_35053.n76 a_33249_35053.t53 1.4705
R45352 a_33249_35053.n22 a_33249_35053.t75 1.4705
R45353 a_33249_35053.n22 a_33249_35053.t21 1.4705
R45354 a_33249_35053.n23 a_33249_35053.t74 1.4705
R45355 a_33249_35053.n23 a_33249_35053.t19 1.4705
R45356 a_33249_35053.n84 a_33249_35053.t82 1.4705
R45357 a_33249_35053.n84 a_33249_35053.t26 1.4705
R45358 a_33249_35053.n85 a_33249_35053.t81 1.4705
R45359 a_33249_35053.n85 a_33249_35053.t24 1.4705
R45360 a_33249_35053.n92 a_33249_35053.t86 1.4705
R45361 a_33249_35053.n92 a_33249_35053.t16 1.4705
R45362 a_33249_35053.n93 a_33249_35053.t85 1.4705
R45363 a_33249_35053.n93 a_33249_35053.t15 1.4705
R45364 a_33249_35053.n17 a_33249_35053.t27 1.4705
R45365 a_33249_35053.n17 a_33249_35053.t56 1.4705
R45366 a_33249_35053.n18 a_33249_35053.t25 1.4705
R45367 a_33249_35053.n18 a_33249_35053.t54 1.4705
R45368 a_33249_35053.n151 a_33249_35053.n150 1.46537
R45369 a_33249_35053.n146 a_33249_35053.n145 1.46537
R45370 a_33249_35053.n142 a_33249_35053.n141 1.46537
R45371 a_33249_35053.n138 a_33249_35053.n137 1.46537
R45372 a_33249_35053.n46 a_33249_35053.n45 1.46537
R45373 a_33249_35053.n48 a_33249_35053.n47 1.46537
R45374 a_33249_35053.n55 a_33249_35053.n54 1.46537
R45375 a_33249_35053.n57 a_33249_35053.n56 1.46537
R45376 a_33249_35053.n59 a_33249_35053.n58 1.46537
R45377 a_33249_35053.n63 a_33249_35053.n62 1.46537
R45378 a_33249_35053.n65 a_33249_35053.n64 1.46537
R45379 a_33249_35053.n41 a_33249_35053.n40 1.46537
R45380 a_33249_35053.n25 a_33249_35053.n24 1.46537
R45381 a_33249_35053.n27 a_33249_35053.n26 1.46537
R45382 a_33249_35053.n87 a_33249_35053.n86 1.46537
R45383 a_33249_35053.n89 a_33249_35053.n88 1.46537
R45384 a_33249_35053.n91 a_33249_35053.n90 1.46537
R45385 a_33249_35053.n95 a_33249_35053.n94 1.46537
R45386 a_33249_35053.n97 a_33249_35053.n96 1.46537
R45387 a_33249_35053.n20 a_33249_35053.n19 1.46537
R45388 a_33249_35053.n114 a_33249_35053.n113 1.46537
R45389 a_33249_35053.n118 a_33249_35053.n117 1.46537
R45390 a_33249_35053.n120 a_33249_35053.n119 1.46537
R45391 a_33249_35053.n153 a_33249_35053.n152 1.46535
R45392 a_33249_35053.n136 a_33249_35053.n135 1.46535
R45393 a_33249_35053.n50 a_33249_35053.n49 1.46535
R45394 a_33249_35053.n67 a_33249_35053.n66 1.46535
R45395 a_33249_35053.n29 a_33249_35053.n28 1.46535
R45396 a_33249_35053.n99 a_33249_35053.n98 1.46535
R45397 a_33249_35053.n106 a_33249_35053.n105 1.43535
R45398 a_33249_35053.n124 a_33249_35053.n123 1.31908
R45399 a_33249_35053.n36 a_33249_35053.n35 1.27228
R45400 a_33249_35053.n65 a_33249_35053.n63 1.27228
R45401 a_33249_35053.n63 a_33249_35053.n59 1.27228
R45402 a_33249_35053.n57 a_33249_35053.n55 1.27228
R45403 a_33249_35053.n48 a_33249_35053.n46 1.27228
R45404 a_33249_35053.n77 a_33249_35053.n75 1.27228
R45405 a_33249_35053.n97 a_33249_35053.n95 1.27228
R45406 a_33249_35053.n95 a_33249_35053.n91 1.27228
R45407 a_33249_35053.n89 a_33249_35053.n87 1.27228
R45408 a_33249_35053.n27 a_33249_35053.n25 1.27228
R45409 a_33249_35053.n157 a_33249_35053.t127 1.2605
R45410 a_33249_35053.n157 a_33249_35053.t125 1.2605
R45411 a_33249_35053.n132 a_33249_35053.t113 1.2605
R45412 a_33249_35053.n132 a_33249_35053.t111 1.2605
R45413 a_33249_35053.n147 a_33249_35053.t118 1.2605
R45414 a_33249_35053.n147 a_33249_35053.t136 1.2605
R45415 a_33249_35053.n148 a_33249_35053.t112 1.2605
R45416 a_33249_35053.n148 a_33249_35053.t132 1.2605
R45417 a_33249_35053.n143 a_33249_35053.t121 1.2605
R45418 a_33249_35053.n143 a_33249_35053.t133 1.2605
R45419 a_33249_35053.n144 a_33249_35053.t116 1.2605
R45420 a_33249_35053.n144 a_33249_35053.t131 1.2605
R45421 a_33249_35053.n139 a_33249_35053.t138 1.2605
R45422 a_33249_35053.n139 a_33249_35053.t110 1.2605
R45423 a_33249_35053.n140 a_33249_35053.t135 1.2605
R45424 a_33249_35053.n140 a_33249_35053.t108 1.2605
R45425 a_33249_35053.n11 a_33249_35053.t109 1.2605
R45426 a_33249_35053.n11 a_33249_35053.t122 1.2605
R45427 a_33249_35053.n12 a_33249_35053.t107 1.2605
R45428 a_33249_35053.n12 a_33249_35053.t119 1.2605
R45429 a_33249_35053.n111 a_33249_35053.t101 1.2605
R45430 a_33249_35053.n111 a_33249_35053.t95 1.2605
R45431 a_33249_35053.n112 a_33249_35053.t89 1.2605
R45432 a_33249_35053.n112 a_33249_35053.t91 1.2605
R45433 a_33249_35053.n115 a_33249_35053.t102 1.2605
R45434 a_33249_35053.n115 a_33249_35053.t100 1.2605
R45435 a_33249_35053.n116 a_33249_35053.t96 1.2605
R45436 a_33249_35053.n116 a_33249_35053.t99 1.2605
R45437 a_33249_35053.n107 a_33249_35053.t98 1.2605
R45438 a_33249_35053.n107 a_33249_35053.t105 1.2605
R45439 a_33249_35053.n122 a_33249_35053.t90 1.2605
R45440 a_33249_35053.n122 a_33249_35053.t92 1.2605
R45441 a_33249_35053.n125 a_33249_35053.t128 1.2605
R45442 a_33249_35053.n125 a_33249_35053.t141 1.2605
R45443 a_33249_35053.n128 a_33249_35053.t114 1.2605
R45444 a_33249_35053.n128 a_33249_35053.t129 1.2605
R45445 a_33249_35053.n130 a_33249_35053.n129 1.25428
R45446 a_33249_35053.n142 a_33249_35053.n138 1.25428
R45447 a_33249_35053.n120 a_33249_35053.n118 1.25428
R45448 a_33249_35053.n127 a_33249_35053.n126 1.04573
R45449 a_33249_35053.n33 a_33249_35053.n32 1.01873
R45450 a_33249_35053.n80 a_33249_35053.n79 1.01873
R45451 a_33249_35053.n70 a_33249_35053.n69 0.778574
R45452 a_33249_35053.n105 a_33249_35053.n101 0.778574
R45453 a_33249_35053.n74 a_33249_35053.n30 0.778574
R45454 a_33249_35053.n82 a_33249_35053.n14 0.778574
R45455 a_33249_35053.n101 a_33249_35053.n15 0.738439
R45456 a_33249_35053.n82 a_33249_35053.n81 0.738439
R45457 a_33249_35053.n133 a_33249_35053.n131 0.738439
R45458 a_33249_35053.n155 a_33249_35053.n10 0.738439
R45459 a_33249_35053.n121 a_33249_35053.n109 0.737223
R45460 a_33249_35053.n68 a_33249_35053.n67 0.699581
R45461 a_33249_35053.n51 a_33249_35053.n50 0.699581
R45462 a_33249_35053.n100 a_33249_35053.n99 0.699581
R45463 a_33249_35053.n83 a_33249_35053.n29 0.699581
R45464 a_33249_35053.n136 a_33249_35053.n134 0.699581
R45465 a_33249_35053.n154 a_33249_35053.n153 0.699581
R45466 a_33249_35053.n123 a_33249_35053.n121 0.585196
R45467 a_33249_35053.n68 a_33249_35053.n41 0.557791
R45468 a_33249_35053.n55 a_33249_35053.n51 0.557791
R45469 a_33249_35053.n100 a_33249_35053.n20 0.557791
R45470 a_33249_35053.n87 a_33249_35053.n83 0.557791
R45471 a_33249_35053.n154 a_33249_35053.n146 0.539791
R45472 a_33249_35053.n70 a_33249_35053.n15 0.530466
R45473 a_33249_35053.n81 a_33249_35053.n74 0.530466
R45474 a_33249_35053.n7 a_33249_35053.n8 1.27228
R45475 a_33249_35053.n73 a_33249_35053.n7 7.30549
R45476 a_33249_35053.t34 a_33249_35053.n6 6.96214
R45477 a_33249_35053.n4 a_33249_35053.n5 1.27228
R45478 a_33249_35053.n104 a_33249_35053.n4 7.30549
R45479 a_33249_35053.t44 a_33249_35053.n3 6.96214
R45480 a_33249_35053.n122 a_33249_35053.n9 5.45652
R45481 a_33249_35053.n1 a_33249_35053.n2 1.25428
R45482 a_33249_35053.n1 a_33249_35053.n156 5.95549
R45483 a_33249_35053.t140 a_33249_35053.n0 7.10317
R45484 a_31953_n19727.n226 a_31953_n19727.n321 15.3954
R45485 a_31953_n19727.n321 a_31953_n19727.t73 13.6649
R45486 a_31953_n19727.n233 a_31953_n19727.t99 10.1674
R45487 a_31953_n19727.t174 a_31953_n19727.n238 10.1674
R45488 a_31953_n19727.n239 a_31953_n19727.t174 10.1674
R45489 a_31953_n19727.t159 a_31953_n19727.n242 10.1674
R45490 a_31953_n19727.n243 a_31953_n19727.t159 10.1674
R45491 a_31953_n19727.n255 a_31953_n19727.t238 10.1674
R45492 a_31953_n19727.t238 a_31953_n19727.n254 10.1674
R45493 a_31953_n19727.n251 a_31953_n19727.t311 10.1674
R45494 a_31953_n19727.t311 a_31953_n19727.n250 10.1674
R45495 a_31953_n19727.n247 a_31953_n19727.t299 10.1674
R45496 a_31953_n19727.t299 a_31953_n19727.n246 10.1674
R45497 a_31953_n19727.t78 a_31953_n19727.n263 10.1674
R45498 a_31953_n19727.n264 a_31953_n19727.t78 10.1674
R45499 a_31953_n19727.t146 a_31953_n19727.n267 10.1674
R45500 a_31953_n19727.n268 a_31953_n19727.t146 10.1674
R45501 a_31953_n19727.t128 a_31953_n19727.n271 10.1674
R45502 a_31953_n19727.n272 a_31953_n19727.t128 10.1674
R45503 a_31953_n19727.n466 a_31953_n19727.t246 10.1674
R45504 a_31953_n19727.t317 a_31953_n19727.n471 10.1674
R45505 a_31953_n19727.n472 a_31953_n19727.t317 10.1674
R45506 a_31953_n19727.t98 a_31953_n19727.n475 10.1674
R45507 a_31953_n19727.n476 a_31953_n19727.t98 10.1674
R45508 a_31953_n19727.t86 a_31953_n19727.n483 10.1674
R45509 a_31953_n19727.n484 a_31953_n19727.t86 10.1674
R45510 a_31953_n19727.t158 a_31953_n19727.n487 10.1674
R45511 a_31953_n19727.n488 a_31953_n19727.t158 10.1674
R45512 a_31953_n19727.t222 a_31953_n19727.n491 10.1674
R45513 a_31953_n19727.n492 a_31953_n19727.t222 10.1674
R45514 a_31953_n19727.n505 a_31953_n19727.t296 10.1674
R45515 a_31953_n19727.t296 a_31953_n19727.n504 10.1674
R45516 a_31953_n19727.n501 a_31953_n19727.t354 10.1674
R45517 a_31953_n19727.t354 a_31953_n19727.n500 10.1674
R45518 a_31953_n19727.n499 a_31953_n19727.t137 10.1674
R45519 a_31953_n19727.t137 a_31953_n19727.n498 10.1674
R45520 a_31953_n19727.n279 a_31953_n19727.t180 10.1674
R45521 a_31953_n19727.t255 a_31953_n19727.n284 10.1674
R45522 a_31953_n19727.n285 a_31953_n19727.t255 10.1674
R45523 a_31953_n19727.t240 a_31953_n19727.n288 10.1674
R45524 a_31953_n19727.n289 a_31953_n19727.t240 10.1674
R45525 a_31953_n19727.n301 a_31953_n19727.t312 10.1674
R45526 a_31953_n19727.t312 a_31953_n19727.n300 10.1674
R45527 a_31953_n19727.n297 a_31953_n19727.t91 10.1674
R45528 a_31953_n19727.t91 a_31953_n19727.n296 10.1674
R45529 a_31953_n19727.n293 a_31953_n19727.t81 10.1674
R45530 a_31953_n19727.t81 a_31953_n19727.n292 10.1674
R45531 a_31953_n19727.t151 a_31953_n19727.n309 10.1674
R45532 a_31953_n19727.n310 a_31953_n19727.t151 10.1674
R45533 a_31953_n19727.t231 a_31953_n19727.n313 10.1674
R45534 a_31953_n19727.n314 a_31953_n19727.t231 10.1674
R45535 a_31953_n19727.t210 a_31953_n19727.n317 10.1674
R45536 a_31953_n19727.n318 a_31953_n19727.t210 10.1674
R45537 a_31953_n19727.n364 a_31953_n19727.t126 10.1674
R45538 a_31953_n19727.n360 a_31953_n19727.t203 10.1674
R45539 a_31953_n19727.t203 a_31953_n19727.n359 10.1674
R45540 a_31953_n19727.n356 a_31953_n19727.t279 10.1674
R45541 a_31953_n19727.t279 a_31953_n19727.n355 10.1674
R45542 a_31953_n19727.t266 a_31953_n19727.n325 10.1674
R45543 a_31953_n19727.n326 a_31953_n19727.t266 10.1674
R45544 a_31953_n19727.t336 a_31953_n19727.n329 10.1674
R45545 a_31953_n19727.n330 a_31953_n19727.t336 10.1674
R45546 a_31953_n19727.t103 a_31953_n19727.n333 10.1674
R45547 a_31953_n19727.n334 a_31953_n19727.t103 10.1674
R45548 a_31953_n19727.n347 a_31953_n19727.t179 10.1674
R45549 a_31953_n19727.t179 a_31953_n19727.n346 10.1674
R45550 a_31953_n19727.n343 a_31953_n19727.t235 10.1674
R45551 a_31953_n19727.t235 a_31953_n19727.n342 10.1674
R45552 a_31953_n19727.n341 a_31953_n19727.t309 10.1674
R45553 a_31953_n19727.t309 a_31953_n19727.n340 10.1674
R45554 a_31953_n19727.n373 a_31953_n19727.t293 10.1674
R45555 a_31953_n19727.t74 a_31953_n19727.n378 10.1674
R45556 a_31953_n19727.n379 a_31953_n19727.t74 10.1674
R45557 a_31953_n19727.t356 a_31953_n19727.n382 10.1674
R45558 a_31953_n19727.n383 a_31953_n19727.t356 10.1674
R45559 a_31953_n19727.n395 a_31953_n19727.t138 10.1674
R45560 a_31953_n19727.t138 a_31953_n19727.n394 10.1674
R45561 a_31953_n19727.n391 a_31953_n19727.t215 10.1674
R45562 a_31953_n19727.t215 a_31953_n19727.n390 10.1674
R45563 a_31953_n19727.n387 a_31953_n19727.t200 10.1674
R45564 a_31953_n19727.t200 a_31953_n19727.n386 10.1674
R45565 a_31953_n19727.t278 a_31953_n19727.n403 10.1674
R45566 a_31953_n19727.n404 a_31953_n19727.t278 10.1674
R45567 a_31953_n19727.t351 a_31953_n19727.n407 10.1674
R45568 a_31953_n19727.n408 a_31953_n19727.t351 10.1674
R45569 a_31953_n19727.t318 a_31953_n19727.n411 10.1674
R45570 a_31953_n19727.n412 a_31953_n19727.t318 10.1674
R45571 a_31953_n19727.n457 a_31953_n19727.t90 10.1674
R45572 a_31953_n19727.n453 a_31953_n19727.t166 10.1674
R45573 a_31953_n19727.t166 a_31953_n19727.n452 10.1674
R45574 a_31953_n19727.n449 a_31953_n19727.t245 10.1674
R45575 a_31953_n19727.t245 a_31953_n19727.n448 10.1674
R45576 a_31953_n19727.t230 a_31953_n19727.n418 10.1674
R45577 a_31953_n19727.n419 a_31953_n19727.t230 10.1674
R45578 a_31953_n19727.t304 a_31953_n19727.n422 10.1674
R45579 a_31953_n19727.n423 a_31953_n19727.t304 10.1674
R45580 a_31953_n19727.t360 a_31953_n19727.n426 10.1674
R45581 a_31953_n19727.n427 a_31953_n19727.t360 10.1674
R45582 a_31953_n19727.n440 a_31953_n19727.t142 10.1674
R45583 a_31953_n19727.t142 a_31953_n19727.n439 10.1674
R45584 a_31953_n19727.n436 a_31953_n19727.t209 10.1674
R45585 a_31953_n19727.t209 a_31953_n19727.n435 10.1674
R45586 a_31953_n19727.n434 a_31953_n19727.t282 10.1674
R45587 a_31953_n19727.t282 a_31953_n19727.n433 10.1674
R45588 a_31953_n19727.n235 a_31953_n19727.t197 10.1674
R45589 a_31953_n19727.t276 a_31953_n19727.n240 10.1674
R45590 a_31953_n19727.n241 a_31953_n19727.t276 10.1674
R45591 a_31953_n19727.t262 a_31953_n19727.n244 10.1674
R45592 a_31953_n19727.n245 a_31953_n19727.t262 10.1674
R45593 a_31953_n19727.n257 a_31953_n19727.t333 10.1674
R45594 a_31953_n19727.t333 a_31953_n19727.n256 10.1674
R45595 a_31953_n19727.n253 a_31953_n19727.t117 10.1674
R45596 a_31953_n19727.t117 a_31953_n19727.n252 10.1674
R45597 a_31953_n19727.n249 a_31953_n19727.t102 10.1674
R45598 a_31953_n19727.t102 a_31953_n19727.n248 10.1674
R45599 a_31953_n19727.t177 a_31953_n19727.n265 10.1674
R45600 a_31953_n19727.n266 a_31953_n19727.t177 10.1674
R45601 a_31953_n19727.t253 a_31953_n19727.n269 10.1674
R45602 a_31953_n19727.n270 a_31953_n19727.t253 10.1674
R45603 a_31953_n19727.t224 a_31953_n19727.n273 10.1674
R45604 a_31953_n19727.n274 a_31953_n19727.t224 10.1674
R45605 a_31953_n19727.n468 a_31953_n19727.t290 10.1674
R45606 a_31953_n19727.t361 a_31953_n19727.n473 10.1674
R45607 a_31953_n19727.n474 a_31953_n19727.t361 10.1674
R45608 a_31953_n19727.t143 a_31953_n19727.n477 10.1674
R45609 a_31953_n19727.n478 a_31953_n19727.t143 10.1674
R45610 a_31953_n19727.t135 a_31953_n19727.n485 10.1674
R45611 a_31953_n19727.n486 a_31953_n19727.t135 10.1674
R45612 a_31953_n19727.t214 a_31953_n19727.n489 10.1674
R45613 a_31953_n19727.n490 a_31953_n19727.t214 10.1674
R45614 a_31953_n19727.t274 a_31953_n19727.n493 10.1674
R45615 a_31953_n19727.n494 a_31953_n19727.t274 10.1674
R45616 a_31953_n19727.n507 a_31953_n19727.t346 10.1674
R45617 a_31953_n19727.t346 a_31953_n19727.n506 10.1674
R45618 a_31953_n19727.n503 a_31953_n19727.t110 10.1674
R45619 a_31953_n19727.t110 a_31953_n19727.n502 10.1674
R45620 a_31953_n19727.t184 a_31953_n19727.n496 10.1674
R45621 a_31953_n19727.n497 a_31953_n19727.t184 10.1674
R45622 a_31953_n19727.n281 a_31953_n19727.t114 10.1674
R45623 a_31953_n19727.t189 a_31953_n19727.n286 10.1674
R45624 a_31953_n19727.n287 a_31953_n19727.t189 10.1674
R45625 a_31953_n19727.t172 a_31953_n19727.n290 10.1674
R45626 a_31953_n19727.n291 a_31953_n19727.t172 10.1674
R45627 a_31953_n19727.n303 a_31953_n19727.t251 10.1674
R45628 a_31953_n19727.t251 a_31953_n19727.n302 10.1674
R45629 a_31953_n19727.n299 a_31953_n19727.t320 10.1674
R45630 a_31953_n19727.t320 a_31953_n19727.n298 10.1674
R45631 a_31953_n19727.n295 a_31953_n19727.t310 10.1674
R45632 a_31953_n19727.t310 a_31953_n19727.n294 10.1674
R45633 a_31953_n19727.t89 a_31953_n19727.n311 10.1674
R45634 a_31953_n19727.n312 a_31953_n19727.t89 10.1674
R45635 a_31953_n19727.t164 a_31953_n19727.n315 10.1674
R45636 a_31953_n19727.n316 a_31953_n19727.t164 10.1674
R45637 a_31953_n19727.t139 a_31953_n19727.n319 10.1674
R45638 a_31953_n19727.n320 a_31953_n19727.t139 10.1674
R45639 a_31953_n19727.n366 a_31953_n19727.t305 10.1674
R45640 a_31953_n19727.n362 a_31953_n19727.t87 10.1674
R45641 a_31953_n19727.t87 a_31953_n19727.n361 10.1674
R45642 a_31953_n19727.n358 a_31953_n19727.t161 10.1674
R45643 a_31953_n19727.t161 a_31953_n19727.n357 10.1674
R45644 a_31953_n19727.t145 a_31953_n19727.n327 10.1674
R45645 a_31953_n19727.n328 a_31953_n19727.t145 10.1674
R45646 a_31953_n19727.t226 a_31953_n19727.n331 10.1674
R45647 a_31953_n19727.n332 a_31953_n19727.t226 10.1674
R45648 a_31953_n19727.t288 a_31953_n19727.n335 10.1674
R45649 a_31953_n19727.n336 a_31953_n19727.t288 10.1674
R45650 a_31953_n19727.n349 a_31953_n19727.t359 10.1674
R45651 a_31953_n19727.t359 a_31953_n19727.n348 10.1674
R45652 a_31953_n19727.n345 a_31953_n19727.t125 10.1674
R45653 a_31953_n19727.t125 a_31953_n19727.n344 10.1674
R45654 a_31953_n19727.t202 a_31953_n19727.n338 10.1674
R45655 a_31953_n19727.n339 a_31953_n19727.t202 10.1674
R45656 a_31953_n19727.n375 a_31953_n19727.t258 10.1674
R45657 a_31953_n19727.t326 a_31953_n19727.n380 10.1674
R45658 a_31953_n19727.n381 a_31953_n19727.t326 10.1674
R45659 a_31953_n19727.t314 a_31953_n19727.n384 10.1674
R45660 a_31953_n19727.n385 a_31953_n19727.t314 10.1674
R45661 a_31953_n19727.n397 a_31953_n19727.t94 10.1674
R45662 a_31953_n19727.t94 a_31953_n19727.n396 10.1674
R45663 a_31953_n19727.n393 a_31953_n19727.t168 10.1674
R45664 a_31953_n19727.t168 a_31953_n19727.n392 10.1674
R45665 a_31953_n19727.n389 a_31953_n19727.t155 10.1674
R45666 a_31953_n19727.t155 a_31953_n19727.n388 10.1674
R45667 a_31953_n19727.t234 a_31953_n19727.n405 10.1674
R45668 a_31953_n19727.n406 a_31953_n19727.t234 10.1674
R45669 a_31953_n19727.t308 a_31953_n19727.n409 10.1674
R45670 a_31953_n19727.n410 a_31953_n19727.t308 10.1674
R45671 a_31953_n19727.t285 a_31953_n19727.n413 10.1674
R45672 a_31953_n19727.n414 a_31953_n19727.t285 10.1674
R45673 a_31953_n19727.n459 a_31953_n19727.t193 10.1674
R45674 a_31953_n19727.n455 a_31953_n19727.t268 10.1674
R45675 a_31953_n19727.t268 a_31953_n19727.n454 10.1674
R45676 a_31953_n19727.n451 a_31953_n19727.t340 10.1674
R45677 a_31953_n19727.t340 a_31953_n19727.n450 10.1674
R45678 a_31953_n19727.t323 a_31953_n19727.n420 10.1674
R45679 a_31953_n19727.n421 a_31953_n19727.t323 10.1674
R45680 a_31953_n19727.t108 a_31953_n19727.n424 10.1674
R45681 a_31953_n19727.n425 a_31953_n19727.t108 10.1674
R45682 a_31953_n19727.t165 a_31953_n19727.n428 10.1674
R45683 a_31953_n19727.n429 a_31953_n19727.t165 10.1674
R45684 a_31953_n19727.n442 a_31953_n19727.t244 10.1674
R45685 a_31953_n19727.t244 a_31953_n19727.n441 10.1674
R45686 a_31953_n19727.n438 a_31953_n19727.t300 10.1674
R45687 a_31953_n19727.t300 a_31953_n19727.n437 10.1674
R45688 a_31953_n19727.t80 a_31953_n19727.n431 10.1674
R45689 a_31953_n19727.n432 a_31953_n19727.t80 10.1674
R45690 a_31953_n19727.t99 a_31953_n19727.n232 10.1409
R45691 a_31953_n19727.t246 a_31953_n19727.n465 10.1409
R45692 a_31953_n19727.t180 a_31953_n19727.n278 10.1409
R45693 a_31953_n19727.t126 a_31953_n19727.n363 10.1409
R45694 a_31953_n19727.t293 a_31953_n19727.n372 10.1409
R45695 a_31953_n19727.t90 a_31953_n19727.n456 10.1409
R45696 a_31953_n19727.t197 a_31953_n19727.n234 10.1409
R45697 a_31953_n19727.t290 a_31953_n19727.n467 10.1409
R45698 a_31953_n19727.t114 a_31953_n19727.n280 10.1409
R45699 a_31953_n19727.t305 a_31953_n19727.n365 10.1409
R45700 a_31953_n19727.t258 a_31953_n19727.n374 10.1409
R45701 a_31953_n19727.t193 a_31953_n19727.n458 10.1409
R45702 a_31953_n19727.t195 a_31953_n19727.n232 9.54631
R45703 a_31953_n19727.n214 a_31953_n19727.t273 9.54631
R45704 a_31953_n19727.t100 a_31953_n19727.n213 9.54631
R45705 a_31953_n19727.n234 a_31953_n19727.t208 9.54631
R45706 a_31953_n19727.t141 a_31953_n19727.n465 9.54631
R45707 a_31953_n19727.n216 a_31953_n19727.t330 9.54631
R45708 a_31953_n19727.t104 a_31953_n19727.n215 9.54631
R45709 a_31953_n19727.n467 a_31953_n19727.t358 9.54631
R45710 a_31953_n19727.t275 a_31953_n19727.n278 9.54631
R45711 a_31953_n19727.n218 a_31953_n19727.t187 9.54631
R45712 a_31953_n19727.t181 a_31953_n19727.n217 9.54631
R45713 a_31953_n19727.n280 a_31953_n19727.t286 9.54631
R45714 a_31953_n19727.t315 a_31953_n19727.n363 9.54631
R45715 a_31953_n19727.n220 a_31953_n19727.t350 9.54631
R45716 a_31953_n19727.t283 a_31953_n19727.n219 9.54631
R45717 a_31953_n19727.n365 a_31953_n19727.t243 9.54631
R45718 a_31953_n19727.t316 a_31953_n19727.n372 9.54631
R45719 a_31953_n19727.n222 a_31953_n19727.t130 9.54631
R45720 a_31953_n19727.t348 a_31953_n19727.n221 9.54631
R45721 a_31953_n19727.n374 a_31953_n19727.t132 9.54631
R45722 a_31953_n19727.t196 a_31953_n19727.n456 9.54631
R45723 a_31953_n19727.n224 a_31953_n19727.t148 9.54631
R45724 a_31953_n19727.t227 a_31953_n19727.n223 9.54631
R45725 a_31953_n19727.n458 a_31953_n19727.t123 9.54631
R45726 a_31953_n19727.n233 a_31953_n19727.t195 9.54355
R45727 a_31953_n19727.t273 a_31953_n19727.n237 9.54355
R45728 a_31953_n19727.n236 a_31953_n19727.t100 9.54355
R45729 a_31953_n19727.n235 a_31953_n19727.t208 9.54355
R45730 a_31953_n19727.n239 a_31953_n19727.t271 9.54355
R45731 a_31953_n19727.t271 a_31953_n19727.n238 9.54355
R45732 a_31953_n19727.t345 a_31953_n19727.n4 9.54355
R45733 a_31953_n19727.n1 a_31953_n19727.t345 9.54355
R45734 a_31953_n19727.n2 a_31953_n19727.t175 9.54355
R45735 a_31953_n19727.t175 a_31953_n19727.n0 9.54355
R45736 a_31953_n19727.n241 a_31953_n19727.t281 9.54355
R45737 a_31953_n19727.n240 a_31953_n19727.t281 9.54355
R45738 a_31953_n19727.n243 a_31953_n19727.t259 9.54355
R45739 a_31953_n19727.t259 a_31953_n19727.n242 9.54355
R45740 a_31953_n19727.t329 a_31953_n19727.n8 9.54355
R45741 a_31953_n19727.n6 a_31953_n19727.t329 9.54355
R45742 a_31953_n19727.n7 a_31953_n19727.t160 9.54355
R45743 a_31953_n19727.t160 a_31953_n19727.n5 9.54355
R45744 a_31953_n19727.n245 a_31953_n19727.t270 9.54355
R45745 a_31953_n19727.n244 a_31953_n19727.t270 9.54355
R45746 a_31953_n19727.t327 a_31953_n19727.n254 9.54355
R45747 a_31953_n19727.n255 a_31953_n19727.t327 9.54355
R45748 a_31953_n19727.n13 a_31953_n19727.t60 9.54355
R45749 a_31953_n19727.t60 a_31953_n19727.n11 9.54355
R45750 a_31953_n19727.t38 a_31953_n19727.n12 9.54355
R45751 a_31953_n19727.n9 a_31953_n19727.t38 9.54355
R45752 a_31953_n19727.n256 a_31953_n19727.t342 9.54355
R45753 a_31953_n19727.n257 a_31953_n19727.t342 9.54355
R45754 a_31953_n19727.t112 a_31953_n19727.n250 9.54355
R45755 a_31953_n19727.n251 a_31953_n19727.t112 9.54355
R45756 a_31953_n19727.n17 a_31953_n19727.t48 9.54355
R45757 a_31953_n19727.t48 a_31953_n19727.n15 9.54355
R45758 a_31953_n19727.t16 a_31953_n19727.n16 9.54355
R45759 a_31953_n19727.n14 a_31953_n19727.t16 9.54355
R45760 a_31953_n19727.n252 a_31953_n19727.t121 9.54355
R45761 a_31953_n19727.n253 a_31953_n19727.t121 9.54355
R45762 a_31953_n19727.t95 a_31953_n19727.n246 9.54355
R45763 a_31953_n19727.n247 a_31953_n19727.t95 9.54355
R45764 a_31953_n19727.n22 a_31953_n19727.t52 9.54355
R45765 a_31953_n19727.t52 a_31953_n19727.n20 9.54355
R45766 a_31953_n19727.t20 a_31953_n19727.n21 9.54355
R45767 a_31953_n19727.n18 a_31953_n19727.t20 9.54355
R45768 a_31953_n19727.n248 a_31953_n19727.t111 9.54355
R45769 a_31953_n19727.n249 a_31953_n19727.t111 9.54355
R45770 a_31953_n19727.n264 a_31953_n19727.t170 9.54355
R45771 a_31953_n19727.t170 a_31953_n19727.n263 9.54355
R45772 a_31953_n19727.t250 a_31953_n19727.n26 9.54355
R45773 a_31953_n19727.n24 a_31953_n19727.t250 9.54355
R45774 a_31953_n19727.n25 a_31953_n19727.t79 9.54355
R45775 a_31953_n19727.t79 a_31953_n19727.n23 9.54355
R45776 a_31953_n19727.n266 a_31953_n19727.t186 9.54355
R45777 a_31953_n19727.n265 a_31953_n19727.t186 9.54355
R45778 a_31953_n19727.n268 a_31953_n19727.t248 9.54355
R45779 a_31953_n19727.t248 a_31953_n19727.n267 9.54355
R45780 a_31953_n19727.t319 a_31953_n19727.n31 9.54355
R45781 a_31953_n19727.n28 a_31953_n19727.t319 9.54355
R45782 a_31953_n19727.n29 a_31953_n19727.t149 9.54355
R45783 a_31953_n19727.t149 a_31953_n19727.n27 9.54355
R45784 a_31953_n19727.n270 a_31953_n19727.t261 9.54355
R45785 a_31953_n19727.n269 a_31953_n19727.t261 9.54355
R45786 a_31953_n19727.n272 a_31953_n19727.t221 9.54355
R45787 a_31953_n19727.t221 a_31953_n19727.n271 9.54355
R45788 a_31953_n19727.t295 a_31953_n19727.n35 9.54355
R45789 a_31953_n19727.n33 a_31953_n19727.t295 9.54355
R45790 a_31953_n19727.n34 a_31953_n19727.t129 9.54355
R45791 a_31953_n19727.t129 a_31953_n19727.n32 9.54355
R45792 a_31953_n19727.n274 a_31953_n19727.t229 9.54355
R45793 a_31953_n19727.n273 a_31953_n19727.t229 9.54355
R45794 a_31953_n19727.n466 a_31953_n19727.t141 9.54355
R45795 a_31953_n19727.t330 a_31953_n19727.n470 9.54355
R45796 a_31953_n19727.n469 a_31953_n19727.t104 9.54355
R45797 a_31953_n19727.n468 a_31953_n19727.t358 9.54355
R45798 a_31953_n19727.n472 a_31953_n19727.t220 9.54355
R45799 a_31953_n19727.t220 a_31953_n19727.n471 9.54355
R45800 a_31953_n19727.t115 a_31953_n19727.n40 9.54355
R45801 a_31953_n19727.n37 a_31953_n19727.t115 9.54355
R45802 a_31953_n19727.n38 a_31953_n19727.t182 9.54355
R45803 a_31953_n19727.t182 a_31953_n19727.n36 9.54355
R45804 a_31953_n19727.n474 a_31953_n19727.t140 9.54355
R45805 a_31953_n19727.n473 a_31953_n19727.t140 9.54355
R45806 a_31953_n19727.n476 a_31953_n19727.t292 9.54355
R45807 a_31953_n19727.t292 a_31953_n19727.n475 9.54355
R45808 a_31953_n19727.t190 a_31953_n19727.n44 9.54355
R45809 a_31953_n19727.n42 a_31953_n19727.t190 9.54355
R45810 a_31953_n19727.n43 a_31953_n19727.t260 9.54355
R45811 a_31953_n19727.t260 a_31953_n19727.n41 9.54355
R45812 a_31953_n19727.n478 a_31953_n19727.t217 9.54355
R45813 a_31953_n19727.n477 a_31953_n19727.t217 9.54355
R45814 a_31953_n19727.n484 a_31953_n19727.t284 9.54355
R45815 a_31953_n19727.t284 a_31953_n19727.n483 9.54355
R45816 a_31953_n19727.t50 a_31953_n19727.n49 9.54355
R45817 a_31953_n19727.n46 a_31953_n19727.t50 9.54355
R45818 a_31953_n19727.n47 a_31953_n19727.t36 9.54355
R45819 a_31953_n19727.t36 a_31953_n19727.n45 9.54355
R45820 a_31953_n19727.n486 a_31953_n19727.t204 9.54355
R45821 a_31953_n19727.n485 a_31953_n19727.t204 9.54355
R45822 a_31953_n19727.n488 a_31953_n19727.t355 9.54355
R45823 a_31953_n19727.t355 a_31953_n19727.n487 9.54355
R45824 a_31953_n19727.t34 a_31953_n19727.n54 9.54355
R45825 a_31953_n19727.n51 a_31953_n19727.t34 9.54355
R45826 a_31953_n19727.n52 a_31953_n19727.t12 9.54355
R45827 a_31953_n19727.t12 a_31953_n19727.n50 9.54355
R45828 a_31953_n19727.n490 a_31953_n19727.t280 9.54355
R45829 a_31953_n19727.n489 a_31953_n19727.t280 9.54355
R45830 a_31953_n19727.n492 a_31953_n19727.t122 9.54355
R45831 a_31953_n19727.t122 a_31953_n19727.n491 9.54355
R45832 a_31953_n19727.t18 a_31953_n19727.n58 9.54355
R45833 a_31953_n19727.n56 a_31953_n19727.t18 9.54355
R45834 a_31953_n19727.n57 a_31953_n19727.t70 9.54355
R45835 a_31953_n19727.t70 a_31953_n19727.n55 9.54355
R45836 a_31953_n19727.n494 a_31953_n19727.t337 9.54355
R45837 a_31953_n19727.n493 a_31953_n19727.t337 9.54355
R45838 a_31953_n19727.t198 a_31953_n19727.n504 9.54355
R45839 a_31953_n19727.n505 a_31953_n19727.t198 9.54355
R45840 a_31953_n19727.n63 a_31953_n19727.t88 9.54355
R45841 a_31953_n19727.t88 a_31953_n19727.n61 9.54355
R45842 a_31953_n19727.t152 a_31953_n19727.n62 9.54355
R45843 a_31953_n19727.n59 a_31953_n19727.t152 9.54355
R45844 a_31953_n19727.n506 a_31953_n19727.t119 9.54355
R45845 a_31953_n19727.n507 a_31953_n19727.t119 9.54355
R45846 a_31953_n19727.t257 a_31953_n19727.n500 9.54355
R45847 a_31953_n19727.n501 a_31953_n19727.t257 9.54355
R45848 a_31953_n19727.n67 a_31953_n19727.t144 9.54355
R45849 a_31953_n19727.t144 a_31953_n19727.n65 9.54355
R45850 a_31953_n19727.t218 a_31953_n19727.n66 9.54355
R45851 a_31953_n19727.n64 a_31953_n19727.t218 9.54355
R45852 a_31953_n19727.n502 a_31953_n19727.t178 9.54355
R45853 a_31953_n19727.n503 a_31953_n19727.t178 9.54355
R45854 a_31953_n19727.t325 a_31953_n19727.n498 9.54355
R45855 a_31953_n19727.n499 a_31953_n19727.t325 9.54355
R45856 a_31953_n19727.n70 a_31953_n19727.t223 9.54355
R45857 a_31953_n19727.t223 a_31953_n19727.n68 9.54355
R45858 a_31953_n19727.n69 a_31953_n19727.t289 9.54355
R45859 a_31953_n19727.n495 a_31953_n19727.t289 9.54355
R45860 a_31953_n19727.n497 a_31953_n19727.t254 9.54355
R45861 a_31953_n19727.n496 a_31953_n19727.t254 9.54355
R45862 a_31953_n19727.n279 a_31953_n19727.t275 9.54355
R45863 a_31953_n19727.t187 a_31953_n19727.n283 9.54355
R45864 a_31953_n19727.n282 a_31953_n19727.t181 9.54355
R45865 a_31953_n19727.n281 a_31953_n19727.t286 9.54355
R45866 a_31953_n19727.n285 a_31953_n19727.t347 9.54355
R45867 a_31953_n19727.t347 a_31953_n19727.n284 9.54355
R45868 a_31953_n19727.t264 a_31953_n19727.n75 9.54355
R45869 a_31953_n19727.n72 a_31953_n19727.t264 9.54355
R45870 a_31953_n19727.n73 a_31953_n19727.t256 9.54355
R45871 a_31953_n19727.t256 a_31953_n19727.n71 9.54355
R45872 a_31953_n19727.n287 a_31953_n19727.t357 9.54355
R45873 a_31953_n19727.n286 a_31953_n19727.t357 9.54355
R45874 a_31953_n19727.n289 a_31953_n19727.t331 9.54355
R45875 a_31953_n19727.t331 a_31953_n19727.n288 9.54355
R45876 a_31953_n19727.t249 a_31953_n19727.n79 9.54355
R45877 a_31953_n19727.n77 a_31953_n19727.t249 9.54355
R45878 a_31953_n19727.n78 a_31953_n19727.t242 9.54355
R45879 a_31953_n19727.t242 a_31953_n19727.n76 9.54355
R45880 a_31953_n19727.n291 a_31953_n19727.t343 9.54355
R45881 a_31953_n19727.n290 a_31953_n19727.t343 9.54355
R45882 a_31953_n19727.t116 a_31953_n19727.n300 9.54355
R45883 a_31953_n19727.n301 a_31953_n19727.t116 9.54355
R45884 a_31953_n19727.n84 a_31953_n19727.t10 9.54355
R45885 a_31953_n19727.t10 a_31953_n19727.n82 9.54355
R45886 a_31953_n19727.t14 a_31953_n19727.n83 9.54355
R45887 a_31953_n19727.n80 a_31953_n19727.t14 9.54355
R45888 a_31953_n19727.n302 a_31953_n19727.t124 9.54355
R45889 a_31953_n19727.n303 a_31953_n19727.t124 9.54355
R45890 a_31953_n19727.t191 a_31953_n19727.n296 9.54355
R45891 a_31953_n19727.n297 a_31953_n19727.t191 9.54355
R45892 a_31953_n19727.n88 a_31953_n19727.t62 9.54355
R45893 a_31953_n19727.t62 a_31953_n19727.n86 9.54355
R45894 a_31953_n19727.t64 a_31953_n19727.n87 9.54355
R45895 a_31953_n19727.n85 a_31953_n19727.t64 9.54355
R45896 a_31953_n19727.n298 a_31953_n19727.t201 9.54355
R45897 a_31953_n19727.n299 a_31953_n19727.t201 9.54355
R45898 a_31953_n19727.t173 a_31953_n19727.n292 9.54355
R45899 a_31953_n19727.n293 a_31953_n19727.t173 9.54355
R45900 a_31953_n19727.n93 a_31953_n19727.t66 9.54355
R45901 a_31953_n19727.t66 a_31953_n19727.n91 9.54355
R45902 a_31953_n19727.t68 a_31953_n19727.n92 9.54355
R45903 a_31953_n19727.n89 a_31953_n19727.t68 9.54355
R45904 a_31953_n19727.n294 a_31953_n19727.t188 9.54355
R45905 a_31953_n19727.n295 a_31953_n19727.t188 9.54355
R45906 a_31953_n19727.n310 a_31953_n19727.t252 9.54355
R45907 a_31953_n19727.t252 a_31953_n19727.n309 9.54355
R45908 a_31953_n19727.t163 a_31953_n19727.n97 9.54355
R45909 a_31953_n19727.n95 a_31953_n19727.t163 9.54355
R45910 a_31953_n19727.n96 a_31953_n19727.t153 9.54355
R45911 a_31953_n19727.t153 a_31953_n19727.n94 9.54355
R45912 a_31953_n19727.n312 a_31953_n19727.t265 9.54355
R45913 a_31953_n19727.n311 a_31953_n19727.t265 9.54355
R45914 a_31953_n19727.n314 a_31953_n19727.t321 9.54355
R45915 a_31953_n19727.t321 a_31953_n19727.n313 9.54355
R45916 a_31953_n19727.t241 a_31953_n19727.n102 9.54355
R45917 a_31953_n19727.n99 a_31953_n19727.t241 9.54355
R45918 a_31953_n19727.n100 a_31953_n19727.t232 9.54355
R45919 a_31953_n19727.t232 a_31953_n19727.n98 9.54355
R45920 a_31953_n19727.n316 a_31953_n19727.t335 9.54355
R45921 a_31953_n19727.n315 a_31953_n19727.t335 9.54355
R45922 a_31953_n19727.n318 a_31953_n19727.t297 9.54355
R45923 a_31953_n19727.t297 a_31953_n19727.n317 9.54355
R45924 a_31953_n19727.t216 a_31953_n19727.n106 9.54355
R45925 a_31953_n19727.n104 a_31953_n19727.t216 9.54355
R45926 a_31953_n19727.n105 a_31953_n19727.t211 9.54355
R45927 a_31953_n19727.t211 a_31953_n19727.n103 9.54355
R45928 a_31953_n19727.n320 a_31953_n19727.t306 9.54355
R45929 a_31953_n19727.n319 a_31953_n19727.t306 9.54355
R45930 a_31953_n19727.n364 a_31953_n19727.t315 9.54355
R45931 a_31953_n19727.t350 a_31953_n19727.n368 9.54355
R45932 a_31953_n19727.n367 a_31953_n19727.t283 9.54355
R45933 a_31953_n19727.n366 a_31953_n19727.t243 9.54355
R45934 a_31953_n19727.t96 a_31953_n19727.n359 9.54355
R45935 a_31953_n19727.n360 a_31953_n19727.t96 9.54355
R45936 a_31953_n19727.n111 a_31953_n19727.t131 9.54355
R45937 a_31953_n19727.t131 a_31953_n19727.n109 9.54355
R45938 a_31953_n19727.t353 a_31953_n19727.n110 9.54355
R45939 a_31953_n19727.n107 a_31953_n19727.t353 9.54355
R45940 a_31953_n19727.n361 a_31953_n19727.t313 9.54355
R45941 a_31953_n19727.n362 a_31953_n19727.t313 9.54355
R45942 a_31953_n19727.t171 a_31953_n19727.n355 9.54355
R45943 a_31953_n19727.n356 a_31953_n19727.t171 9.54355
R45944 a_31953_n19727.n116 a_31953_n19727.t206 9.54355
R45945 a_31953_n19727.t206 a_31953_n19727.n114 9.54355
R45946 a_31953_n19727.t136 a_31953_n19727.n115 9.54355
R45947 a_31953_n19727.n112 a_31953_n19727.t136 9.54355
R45948 a_31953_n19727.n357 a_31953_n19727.t92 9.54355
R45949 a_31953_n19727.n358 a_31953_n19727.t92 9.54355
R45950 a_31953_n19727.n326 a_31953_n19727.t156 9.54355
R45951 a_31953_n19727.t156 a_31953_n19727.n325 9.54355
R45952 a_31953_n19727.t44 a_31953_n19727.n120 9.54355
R45953 a_31953_n19727.n118 a_31953_n19727.t44 9.54355
R45954 a_31953_n19727.n119 a_31953_n19727.t58 9.54355
R45955 a_31953_n19727.t58 a_31953_n19727.n117 9.54355
R45956 a_31953_n19727.n328 a_31953_n19727.t82 9.54355
R45957 a_31953_n19727.n327 a_31953_n19727.t82 9.54355
R45958 a_31953_n19727.n330 a_31953_n19727.t236 9.54355
R45959 a_31953_n19727.t236 a_31953_n19727.n329 9.54355
R45960 a_31953_n19727.t24 a_31953_n19727.n125 9.54355
R45961 a_31953_n19727.n122 a_31953_n19727.t24 9.54355
R45962 a_31953_n19727.n123 a_31953_n19727.t42 9.54355
R45963 a_31953_n19727.t42 a_31953_n19727.n121 9.54355
R45964 a_31953_n19727.n332 a_31953_n19727.t154 9.54355
R45965 a_31953_n19727.n331 a_31953_n19727.t154 9.54355
R45966 a_31953_n19727.n334 a_31953_n19727.t294 9.54355
R45967 a_31953_n19727.t294 a_31953_n19727.n333 9.54355
R45968 a_31953_n19727.t8 a_31953_n19727.n129 9.54355
R45969 a_31953_n19727.n127 a_31953_n19727.t8 9.54355
R45970 a_31953_n19727.n128 a_31953_n19727.t30 9.54355
R45971 a_31953_n19727.t30 a_31953_n19727.n126 9.54355
R45972 a_31953_n19727.n336 a_31953_n19727.t219 9.54355
R45973 a_31953_n19727.n335 a_31953_n19727.t219 9.54355
R45974 a_31953_n19727.t75 a_31953_n19727.n346 9.54355
R45975 a_31953_n19727.n347 a_31953_n19727.t75 9.54355
R45976 a_31953_n19727.n134 a_31953_n19727.t105 9.54355
R45977 a_31953_n19727.t105 a_31953_n19727.n132 9.54355
R45978 a_31953_n19727.t332 a_31953_n19727.n133 9.54355
R45979 a_31953_n19727.n130 a_31953_n19727.t332 9.54355
R45980 a_31953_n19727.n348 a_31953_n19727.t291 9.54355
R45981 a_31953_n19727.n349 a_31953_n19727.t291 9.54355
R45982 a_31953_n19727.t134 a_31953_n19727.n342 9.54355
R45983 a_31953_n19727.n343 a_31953_n19727.t134 9.54355
R45984 a_31953_n19727.n138 a_31953_n19727.t162 9.54355
R45985 a_31953_n19727.t162 a_31953_n19727.n136 9.54355
R45986 a_31953_n19727.t93 a_31953_n19727.n137 9.54355
R45987 a_31953_n19727.n135 a_31953_n19727.t93 9.54355
R45988 a_31953_n19727.n344 a_31953_n19727.t352 9.54355
R45989 a_31953_n19727.n345 a_31953_n19727.t352 9.54355
R45990 a_31953_n19727.t213 a_31953_n19727.n340 9.54355
R45991 a_31953_n19727.n341 a_31953_n19727.t213 9.54355
R45992 a_31953_n19727.n141 a_31953_n19727.t239 9.54355
R45993 a_31953_n19727.t239 a_31953_n19727.n139 9.54355
R45994 a_31953_n19727.n140 a_31953_n19727.t167 9.54355
R45995 a_31953_n19727.n337 a_31953_n19727.t167 9.54355
R45996 a_31953_n19727.n339 a_31953_n19727.t133 9.54355
R45997 a_31953_n19727.n338 a_31953_n19727.t133 9.54355
R45998 a_31953_n19727.n373 a_31953_n19727.t316 9.54355
R45999 a_31953_n19727.t130 a_31953_n19727.n377 9.54355
R46000 a_31953_n19727.n376 a_31953_n19727.t348 9.54355
R46001 a_31953_n19727.n375 a_31953_n19727.t132 9.54355
R46002 a_31953_n19727.n379 a_31953_n19727.t97 9.54355
R46003 a_31953_n19727.t97 a_31953_n19727.n378 9.54355
R46004 a_31953_n19727.t205 a_31953_n19727.n146 9.54355
R46005 a_31953_n19727.n143 a_31953_n19727.t205 9.54355
R46006 a_31953_n19727.n144 a_31953_n19727.t127 9.54355
R46007 a_31953_n19727.t127 a_31953_n19727.n142 9.54355
R46008 a_31953_n19727.n381 a_31953_n19727.t207 9.54355
R46009 a_31953_n19727.n380 a_31953_n19727.t207 9.54355
R46010 a_31953_n19727.n383 a_31953_n19727.t85 9.54355
R46011 a_31953_n19727.t85 a_31953_n19727.n382 9.54355
R46012 a_31953_n19727.t192 a_31953_n19727.n150 9.54355
R46013 a_31953_n19727.n148 a_31953_n19727.t192 9.54355
R46014 a_31953_n19727.n149 a_31953_n19727.t118 9.54355
R46015 a_31953_n19727.t118 a_31953_n19727.n147 9.54355
R46016 a_31953_n19727.n385 a_31953_n19727.t194 9.54355
R46017 a_31953_n19727.n384 a_31953_n19727.t194 9.54355
R46018 a_31953_n19727.t157 a_31953_n19727.n394 9.54355
R46019 a_31953_n19727.n395 a_31953_n19727.t157 9.54355
R46020 a_31953_n19727.n155 a_31953_n19727.t26 9.54355
R46021 a_31953_n19727.t26 a_31953_n19727.n153 9.54355
R46022 a_31953_n19727.t46 a_31953_n19727.n154 9.54355
R46023 a_31953_n19727.n151 a_31953_n19727.t46 9.54355
R46024 a_31953_n19727.n396 a_31953_n19727.t269 9.54355
R46025 a_31953_n19727.n397 a_31953_n19727.t269 9.54355
R46026 a_31953_n19727.t237 a_31953_n19727.n390 9.54355
R46027 a_31953_n19727.n391 a_31953_n19727.t237 9.54355
R46028 a_31953_n19727.n159 a_31953_n19727.t4 9.54355
R46029 a_31953_n19727.t4 a_31953_n19727.n157 9.54355
R46030 a_31953_n19727.t28 a_31953_n19727.n158 9.54355
R46031 a_31953_n19727.n156 a_31953_n19727.t28 9.54355
R46032 a_31953_n19727.n392 a_31953_n19727.t341 9.54355
R46033 a_31953_n19727.n393 a_31953_n19727.t341 9.54355
R46034 a_31953_n19727.t225 a_31953_n19727.n386 9.54355
R46035 a_31953_n19727.n387 a_31953_n19727.t225 9.54355
R46036 a_31953_n19727.n164 a_31953_n19727.t6 9.54355
R46037 a_31953_n19727.t6 a_31953_n19727.n162 9.54355
R46038 a_31953_n19727.t32 a_31953_n19727.n163 9.54355
R46039 a_31953_n19727.n160 a_31953_n19727.t32 9.54355
R46040 a_31953_n19727.n388 a_31953_n19727.t324 9.54355
R46041 a_31953_n19727.n389 a_31953_n19727.t324 9.54355
R46042 a_31953_n19727.n404 a_31953_n19727.t298 9.54355
R46043 a_31953_n19727.t298 a_31953_n19727.n403 9.54355
R46044 a_31953_n19727.t107 a_31953_n19727.n168 9.54355
R46045 a_31953_n19727.n166 a_31953_n19727.t107 9.54355
R46046 a_31953_n19727.n167 a_31953_n19727.t322 9.54355
R46047 a_31953_n19727.t322 a_31953_n19727.n165 9.54355
R46048 a_31953_n19727.n406 a_31953_n19727.t109 9.54355
R46049 a_31953_n19727.n405 a_31953_n19727.t109 9.54355
R46050 a_31953_n19727.n408 a_31953_n19727.t77 9.54355
R46051 a_31953_n19727.t77 a_31953_n19727.n407 9.54355
R46052 a_31953_n19727.t183 a_31953_n19727.n173 9.54355
R46053 a_31953_n19727.n170 a_31953_n19727.t183 9.54355
R46054 a_31953_n19727.n171 a_31953_n19727.t106 9.54355
R46055 a_31953_n19727.t106 a_31953_n19727.n169 9.54355
R46056 a_31953_n19727.n410 a_31953_n19727.t185 9.54355
R46057 a_31953_n19727.n409 a_31953_n19727.t185 9.54355
R46058 a_31953_n19727.n412 a_31953_n19727.t349 9.54355
R46059 a_31953_n19727.t349 a_31953_n19727.n411 9.54355
R46060 a_31953_n19727.t147 a_31953_n19727.n177 9.54355
R46061 a_31953_n19727.n175 a_31953_n19727.t147 9.54355
R46062 a_31953_n19727.n176 a_31953_n19727.t76 9.54355
R46063 a_31953_n19727.t76 a_31953_n19727.n174 9.54355
R46064 a_31953_n19727.n414 a_31953_n19727.t150 9.54355
R46065 a_31953_n19727.n413 a_31953_n19727.t150 9.54355
R46066 a_31953_n19727.n457 a_31953_n19727.t196 9.54355
R46067 a_31953_n19727.t148 a_31953_n19727.n461 9.54355
R46068 a_31953_n19727.n460 a_31953_n19727.t227 9.54355
R46069 a_31953_n19727.n459 a_31953_n19727.t123 9.54355
R46070 a_31953_n19727.t272 a_31953_n19727.n452 9.54355
R46071 a_31953_n19727.n453 a_31953_n19727.t272 9.54355
R46072 a_31953_n19727.n182 a_31953_n19727.t228 9.54355
R46073 a_31953_n19727.t228 a_31953_n19727.n180 9.54355
R46074 a_31953_n19727.t301 a_31953_n19727.n181 9.54355
R46075 a_31953_n19727.n178 a_31953_n19727.t301 9.54355
R46076 a_31953_n19727.n454 a_31953_n19727.t199 9.54355
R46077 a_31953_n19727.n455 a_31953_n19727.t199 9.54355
R46078 a_31953_n19727.t344 a_31953_n19727.n448 9.54355
R46079 a_31953_n19727.n449 a_31953_n19727.t344 9.54355
R46080 a_31953_n19727.n187 a_31953_n19727.t302 9.54355
R46081 a_31953_n19727.t302 a_31953_n19727.n185 9.54355
R46082 a_31953_n19727.t83 a_31953_n19727.n186 9.54355
R46083 a_31953_n19727.n183 a_31953_n19727.t83 9.54355
R46084 a_31953_n19727.n450 a_31953_n19727.t277 9.54355
R46085 a_31953_n19727.n451 a_31953_n19727.t277 9.54355
R46086 a_31953_n19727.n419 a_31953_n19727.t328 9.54355
R46087 a_31953_n19727.t328 a_31953_n19727.n418 9.54355
R46088 a_31953_n19727.t22 a_31953_n19727.n191 9.54355
R46089 a_31953_n19727.n189 a_31953_n19727.t22 9.54355
R46090 a_31953_n19727.n190 a_31953_n19727.t2 9.54355
R46091 a_31953_n19727.t2 a_31953_n19727.n188 9.54355
R46092 a_31953_n19727.n421 a_31953_n19727.t263 9.54355
R46093 a_31953_n19727.n420 a_31953_n19727.t263 9.54355
R46094 a_31953_n19727.n423 a_31953_n19727.t113 9.54355
R46095 a_31953_n19727.t113 a_31953_n19727.n422 9.54355
R46096 a_31953_n19727.t0 a_31953_n19727.n196 9.54355
R46097 a_31953_n19727.n193 a_31953_n19727.t0 9.54355
R46098 a_31953_n19727.n194 a_31953_n19727.t54 9.54355
R46099 a_31953_n19727.t54 a_31953_n19727.n192 9.54355
R46100 a_31953_n19727.n425 a_31953_n19727.t334 9.54355
R46101 a_31953_n19727.n424 a_31953_n19727.t334 9.54355
R46102 a_31953_n19727.n427 a_31953_n19727.t169 9.54355
R46103 a_31953_n19727.t169 a_31953_n19727.n426 9.54355
R46104 a_31953_n19727.t56 a_31953_n19727.n200 9.54355
R46105 a_31953_n19727.n198 a_31953_n19727.t56 9.54355
R46106 a_31953_n19727.n199 a_31953_n19727.t40 9.54355
R46107 a_31953_n19727.t40 a_31953_n19727.n197 9.54355
R46108 a_31953_n19727.n429 a_31953_n19727.t101 9.54355
R46109 a_31953_n19727.n428 a_31953_n19727.t101 9.54355
R46110 a_31953_n19727.t247 a_31953_n19727.n439 9.54355
R46111 a_31953_n19727.n440 a_31953_n19727.t247 9.54355
R46112 a_31953_n19727.n205 a_31953_n19727.t212 9.54355
R46113 a_31953_n19727.t212 a_31953_n19727.n203 9.54355
R46114 a_31953_n19727.t287 a_31953_n19727.n204 9.54355
R46115 a_31953_n19727.n201 a_31953_n19727.t287 9.54355
R46116 a_31953_n19727.n441 a_31953_n19727.t176 9.54355
R46117 a_31953_n19727.n442 a_31953_n19727.t176 9.54355
R46118 a_31953_n19727.t303 a_31953_n19727.n435 9.54355
R46119 a_31953_n19727.n436 a_31953_n19727.t303 9.54355
R46120 a_31953_n19727.n209 a_31953_n19727.t267 9.54355
R46121 a_31953_n19727.t267 a_31953_n19727.n207 9.54355
R46122 a_31953_n19727.t338 a_31953_n19727.n208 9.54355
R46123 a_31953_n19727.n206 a_31953_n19727.t338 9.54355
R46124 a_31953_n19727.n437 a_31953_n19727.t233 9.54355
R46125 a_31953_n19727.n438 a_31953_n19727.t233 9.54355
R46126 a_31953_n19727.t84 a_31953_n19727.n433 9.54355
R46127 a_31953_n19727.n434 a_31953_n19727.t84 9.54355
R46128 a_31953_n19727.n212 a_31953_n19727.t339 9.54355
R46129 a_31953_n19727.t339 a_31953_n19727.n210 9.54355
R46130 a_31953_n19727.n211 a_31953_n19727.t120 9.54355
R46131 a_31953_n19727.n430 a_31953_n19727.t120 9.54355
R46132 a_31953_n19727.n432 a_31953_n19727.t307 9.54355
R46133 a_31953_n19727.n431 a_31953_n19727.t307 9.54355
R46134 a_31953_n19727.n321 a_31953_n19727.t72 6.62729
R46135 a_31953_n19727.n464 a_31953_n19727.n463 3.90251
R46136 a_31953_n19727.n463 a_31953_n19727.n225 3.89899
R46137 a_31953_n19727.n479 a_31953_n19727.t37 3.3605
R46138 a_31953_n19727.n227 a_31953_n19727.t13 3.3605
R46139 a_31953_n19727.n231 a_31953_n19727.t39 3.3605
R46140 a_31953_n19727.n230 a_31953_n19727.t17 3.3605
R46141 a_31953_n19727.n229 a_31953_n19727.t21 3.3605
R46142 a_31953_n19727.n259 a_31953_n19727.t61 3.3605
R46143 a_31953_n19727.n260 a_31953_n19727.t49 3.3605
R46144 a_31953_n19727.n261 a_31953_n19727.t53 3.3605
R46145 a_31953_n19727.n277 a_31953_n19727.t15 3.3605
R46146 a_31953_n19727.n276 a_31953_n19727.t65 3.3605
R46147 a_31953_n19727.n275 a_31953_n19727.t69 3.3605
R46148 a_31953_n19727.n305 a_31953_n19727.t11 3.3605
R46149 a_31953_n19727.n306 a_31953_n19727.t63 3.3605
R46150 a_31953_n19727.n307 a_31953_n19727.t67 3.3605
R46151 a_31953_n19727.n322 a_31953_n19727.t59 3.3605
R46152 a_31953_n19727.n323 a_31953_n19727.t43 3.3605
R46153 a_31953_n19727.n324 a_31953_n19727.t31 3.3605
R46154 a_31953_n19727.n353 a_31953_n19727.t45 3.3605
R46155 a_31953_n19727.n352 a_31953_n19727.t25 3.3605
R46156 a_31953_n19727.n351 a_31953_n19727.t9 3.3605
R46157 a_31953_n19727.n371 a_31953_n19727.t47 3.3605
R46158 a_31953_n19727.n370 a_31953_n19727.t29 3.3605
R46159 a_31953_n19727.n369 a_31953_n19727.t33 3.3605
R46160 a_31953_n19727.n399 a_31953_n19727.t27 3.3605
R46161 a_31953_n19727.n400 a_31953_n19727.t5 3.3605
R46162 a_31953_n19727.n401 a_31953_n19727.t7 3.3605
R46163 a_31953_n19727.n415 a_31953_n19727.t3 3.3605
R46164 a_31953_n19727.n416 a_31953_n19727.t55 3.3605
R46165 a_31953_n19727.n417 a_31953_n19727.t41 3.3605
R46166 a_31953_n19727.n446 a_31953_n19727.t23 3.3605
R46167 a_31953_n19727.n445 a_31953_n19727.t1 3.3605
R46168 a_31953_n19727.n444 a_31953_n19727.t57 3.3605
R46169 a_31953_n19727.n481 a_31953_n19727.t51 3.3605
R46170 a_31953_n19727.n480 a_31953_n19727.t35 3.3605
R46171 a_31953_n19727.n228 a_31953_n19727.t19 3.3605
R46172 a_31953_n19727.t71 a_31953_n19727.n509 3.3605
R46173 a_31953_n19727.n258 a_31953_n19727.n231 2.59662
R46174 a_31953_n19727.n304 a_31953_n19727.n277 2.59662
R46175 a_31953_n19727.n354 a_31953_n19727.n322 2.59662
R46176 a_31953_n19727.n398 a_31953_n19727.n371 2.59662
R46177 a_31953_n19727.n447 a_31953_n19727.n415 2.59662
R46178 a_31953_n19727.n482 a_31953_n19727.n479 2.59562
R46179 a_31953_n19727.n262 a_31953_n19727.n229 2.59544
R46180 a_31953_n19727.n308 a_31953_n19727.n275 2.59544
R46181 a_31953_n19727.n350 a_31953_n19727.n324 2.59544
R46182 a_31953_n19727.n402 a_31953_n19727.n369 2.59544
R46183 a_31953_n19727.n443 a_31953_n19727.n417 2.59544
R46184 a_31953_n19727.n509 a_31953_n19727.n508 2.59544
R46185 a_31953_n19727.n259 a_31953_n19727.n258 2.58354
R46186 a_31953_n19727.n305 a_31953_n19727.n304 2.58354
R46187 a_31953_n19727.n354 a_31953_n19727.n353 2.58354
R46188 a_31953_n19727.n399 a_31953_n19727.n398 2.58354
R46189 a_31953_n19727.n447 a_31953_n19727.n446 2.58354
R46190 a_31953_n19727.n482 a_31953_n19727.n481 2.58354
R46191 a_31953_n19727.n262 a_31953_n19727.n261 2.58235
R46192 a_31953_n19727.n308 a_31953_n19727.n307 2.58235
R46193 a_31953_n19727.n351 a_31953_n19727.n350 2.58235
R46194 a_31953_n19727.n402 a_31953_n19727.n401 2.58235
R46195 a_31953_n19727.n444 a_31953_n19727.n443 2.58235
R46196 a_31953_n19727.n508 a_31953_n19727.n228 2.58235
R46197 a_31953_n19727.n225 a_31953_n19727.n226 0.0196917
R46198 a_31953_n19727.n131 a_31953_n19727.n139 1.6805
R46199 a_31953_n19727.n202 a_31953_n19727.n210 1.6805
R46200 a_31953_n19727.n60 a_31953_n19727.n68 1.6805
R46201 a_31953_n19727.n74 a_31953_n19727.n218 1.59324
R46202 a_31953_n19727.n145 a_31953_n19727.n222 1.59324
R46203 a_31953_n19727.n3 a_31953_n19727.n214 1.59324
R46204 a_31953_n19727.n350 a_31953_n19727.n131 1.5005
R46205 a_31953_n19727.n113 a_31953_n19727.n354 1.5005
R46206 a_31953_n19727.n90 a_31953_n19727.n308 1.5005
R46207 a_31953_n19727.n304 a_31953_n19727.n74 1.5005
R46208 a_31953_n19727.n131 a_31953_n19727.n141 1.5005
R46209 a_31953_n19727.n131 a_31953_n19727.n138 1.5005
R46210 a_31953_n19727.n136 a_31953_n19727.n131 1.5005
R46211 a_31953_n19727.n131 a_31953_n19727.n134 1.5005
R46212 a_31953_n19727.n132 a_31953_n19727.n131 1.5005
R46213 a_31953_n19727.n129 a_31953_n19727.n124 1.5005
R46214 a_31953_n19727.n131 a_31953_n19727.n127 1.5005
R46215 a_31953_n19727.n125 a_31953_n19727.n124 1.5005
R46216 a_31953_n19727.n124 a_31953_n19727.n122 1.5005
R46217 a_31953_n19727.n120 a_31953_n19727.n113 1.5005
R46218 a_31953_n19727.n124 a_31953_n19727.n118 1.5005
R46219 a_31953_n19727.n108 a_31953_n19727.n116 1.5005
R46220 a_31953_n19727.n114 a_31953_n19727.n113 1.5005
R46221 a_31953_n19727.n108 a_31953_n19727.n111 1.5005
R46222 a_31953_n19727.n109 a_31953_n19727.n108 1.5005
R46223 a_31953_n19727.n108 a_31953_n19727.n220 1.5005
R46224 a_31953_n19727.n106 a_31953_n19727.n101 1.5005
R46225 a_31953_n19727.n101 a_31953_n19727.n104 1.5005
R46226 a_31953_n19727.n102 a_31953_n19727.n101 1.5005
R46227 a_31953_n19727.n101 a_31953_n19727.n99 1.5005
R46228 a_31953_n19727.n97 a_31953_n19727.n90 1.5005
R46229 a_31953_n19727.n101 a_31953_n19727.n95 1.5005
R46230 a_31953_n19727.n81 a_31953_n19727.n93 1.5005
R46231 a_31953_n19727.n91 a_31953_n19727.n90 1.5005
R46232 a_31953_n19727.n81 a_31953_n19727.n88 1.5005
R46233 a_31953_n19727.n86 a_31953_n19727.n81 1.5005
R46234 a_31953_n19727.n74 a_31953_n19727.n84 1.5005
R46235 a_31953_n19727.n82 a_31953_n19727.n81 1.5005
R46236 a_31953_n19727.n79 a_31953_n19727.n74 1.5005
R46237 a_31953_n19727.n74 a_31953_n19727.n77 1.5005
R46238 a_31953_n19727.n75 a_31953_n19727.n74 1.5005
R46239 a_31953_n19727.n74 a_31953_n19727.n72 1.5005
R46240 a_31953_n19727.n443 a_31953_n19727.n202 1.5005
R46241 a_31953_n19727.n184 a_31953_n19727.n447 1.5005
R46242 a_31953_n19727.n161 a_31953_n19727.n402 1.5005
R46243 a_31953_n19727.n398 a_31953_n19727.n145 1.5005
R46244 a_31953_n19727.n202 a_31953_n19727.n212 1.5005
R46245 a_31953_n19727.n202 a_31953_n19727.n209 1.5005
R46246 a_31953_n19727.n207 a_31953_n19727.n202 1.5005
R46247 a_31953_n19727.n202 a_31953_n19727.n205 1.5005
R46248 a_31953_n19727.n203 a_31953_n19727.n202 1.5005
R46249 a_31953_n19727.n200 a_31953_n19727.n195 1.5005
R46250 a_31953_n19727.n202 a_31953_n19727.n198 1.5005
R46251 a_31953_n19727.n196 a_31953_n19727.n195 1.5005
R46252 a_31953_n19727.n195 a_31953_n19727.n193 1.5005
R46253 a_31953_n19727.n191 a_31953_n19727.n184 1.5005
R46254 a_31953_n19727.n195 a_31953_n19727.n189 1.5005
R46255 a_31953_n19727.n179 a_31953_n19727.n187 1.5005
R46256 a_31953_n19727.n185 a_31953_n19727.n184 1.5005
R46257 a_31953_n19727.n179 a_31953_n19727.n182 1.5005
R46258 a_31953_n19727.n180 a_31953_n19727.n179 1.5005
R46259 a_31953_n19727.n179 a_31953_n19727.n224 1.5005
R46260 a_31953_n19727.n177 a_31953_n19727.n172 1.5005
R46261 a_31953_n19727.n172 a_31953_n19727.n175 1.5005
R46262 a_31953_n19727.n173 a_31953_n19727.n172 1.5005
R46263 a_31953_n19727.n172 a_31953_n19727.n170 1.5005
R46264 a_31953_n19727.n168 a_31953_n19727.n161 1.5005
R46265 a_31953_n19727.n172 a_31953_n19727.n166 1.5005
R46266 a_31953_n19727.n152 a_31953_n19727.n164 1.5005
R46267 a_31953_n19727.n162 a_31953_n19727.n161 1.5005
R46268 a_31953_n19727.n152 a_31953_n19727.n159 1.5005
R46269 a_31953_n19727.n157 a_31953_n19727.n152 1.5005
R46270 a_31953_n19727.n145 a_31953_n19727.n155 1.5005
R46271 a_31953_n19727.n153 a_31953_n19727.n152 1.5005
R46272 a_31953_n19727.n150 a_31953_n19727.n145 1.5005
R46273 a_31953_n19727.n145 a_31953_n19727.n148 1.5005
R46274 a_31953_n19727.n146 a_31953_n19727.n145 1.5005
R46275 a_31953_n19727.n145 a_31953_n19727.n143 1.5005
R46276 a_31953_n19727.n48 a_31953_n19727.n482 1.5005
R46277 a_31953_n19727.n19 a_31953_n19727.n262 1.5005
R46278 a_31953_n19727.n258 a_31953_n19727.n3 1.5005
R46279 a_31953_n19727.n60 a_31953_n19727.n70 1.5005
R46280 a_31953_n19727.n60 a_31953_n19727.n67 1.5005
R46281 a_31953_n19727.n65 a_31953_n19727.n60 1.5005
R46282 a_31953_n19727.n60 a_31953_n19727.n63 1.5005
R46283 a_31953_n19727.n61 a_31953_n19727.n60 1.5005
R46284 a_31953_n19727.n58 a_31953_n19727.n53 1.5005
R46285 a_31953_n19727.n60 a_31953_n19727.n56 1.5005
R46286 a_31953_n19727.n54 a_31953_n19727.n53 1.5005
R46287 a_31953_n19727.n53 a_31953_n19727.n51 1.5005
R46288 a_31953_n19727.n49 a_31953_n19727.n48 1.5005
R46289 a_31953_n19727.n53 a_31953_n19727.n46 1.5005
R46290 a_31953_n19727.n44 a_31953_n19727.n39 1.5005
R46291 a_31953_n19727.n48 a_31953_n19727.n42 1.5005
R46292 a_31953_n19727.n40 a_31953_n19727.n39 1.5005
R46293 a_31953_n19727.n39 a_31953_n19727.n37 1.5005
R46294 a_31953_n19727.n39 a_31953_n19727.n216 1.5005
R46295 a_31953_n19727.n35 a_31953_n19727.n30 1.5005
R46296 a_31953_n19727.n30 a_31953_n19727.n33 1.5005
R46297 a_31953_n19727.n31 a_31953_n19727.n30 1.5005
R46298 a_31953_n19727.n30 a_31953_n19727.n28 1.5005
R46299 a_31953_n19727.n26 a_31953_n19727.n19 1.5005
R46300 a_31953_n19727.n30 a_31953_n19727.n24 1.5005
R46301 a_31953_n19727.n10 a_31953_n19727.n22 1.5005
R46302 a_31953_n19727.n20 a_31953_n19727.n19 1.5005
R46303 a_31953_n19727.n10 a_31953_n19727.n17 1.5005
R46304 a_31953_n19727.n15 a_31953_n19727.n10 1.5005
R46305 a_31953_n19727.n3 a_31953_n19727.n13 1.5005
R46306 a_31953_n19727.n11 a_31953_n19727.n10 1.5005
R46307 a_31953_n19727.n8 a_31953_n19727.n3 1.5005
R46308 a_31953_n19727.n3 a_31953_n19727.n6 1.5005
R46309 a_31953_n19727.n4 a_31953_n19727.n3 1.5005
R46310 a_31953_n19727.n3 a_31953_n19727.n1 1.5005
R46311 a_31953_n19727.n508 a_31953_n19727.n60 1.5005
R46312 a_31953_n19727.n260 a_31953_n19727.n259 1.06274
R46313 a_31953_n19727.n261 a_31953_n19727.n260 1.06274
R46314 a_31953_n19727.n231 a_31953_n19727.n230 1.06274
R46315 a_31953_n19727.n230 a_31953_n19727.n229 1.06274
R46316 a_31953_n19727.n306 a_31953_n19727.n305 1.06274
R46317 a_31953_n19727.n307 a_31953_n19727.n306 1.06274
R46318 a_31953_n19727.n277 a_31953_n19727.n276 1.06274
R46319 a_31953_n19727.n276 a_31953_n19727.n275 1.06274
R46320 a_31953_n19727.n353 a_31953_n19727.n352 1.06274
R46321 a_31953_n19727.n352 a_31953_n19727.n351 1.06274
R46322 a_31953_n19727.n323 a_31953_n19727.n322 1.06274
R46323 a_31953_n19727.n324 a_31953_n19727.n323 1.06274
R46324 a_31953_n19727.n400 a_31953_n19727.n399 1.06274
R46325 a_31953_n19727.n401 a_31953_n19727.n400 1.06274
R46326 a_31953_n19727.n371 a_31953_n19727.n370 1.06274
R46327 a_31953_n19727.n370 a_31953_n19727.n369 1.06274
R46328 a_31953_n19727.n446 a_31953_n19727.n445 1.06274
R46329 a_31953_n19727.n445 a_31953_n19727.n444 1.06274
R46330 a_31953_n19727.n416 a_31953_n19727.n415 1.06274
R46331 a_31953_n19727.n417 a_31953_n19727.n416 1.06274
R46332 a_31953_n19727.n481 a_31953_n19727.n480 1.06274
R46333 a_31953_n19727.n480 a_31953_n19727.n228 1.06274
R46334 a_31953_n19727.n479 a_31953_n19727.n227 1.06274
R46335 a_31953_n19727.n509 a_31953_n19727.n227 1.06274
R46336 a_31953_n19727.n236 a_31953_n19727.n235 0.97759
R46337 a_31953_n19727.n237 a_31953_n19727.n233 0.97759
R46338 a_31953_n19727.n240 a_31953_n19727.n0 0.97759
R46339 a_31953_n19727.n1 a_31953_n19727.n238 0.97759
R46340 a_31953_n19727.n2 a_31953_n19727.n241 0.97759
R46341 a_31953_n19727.n4 a_31953_n19727.n239 0.97759
R46342 a_31953_n19727.n244 a_31953_n19727.n5 0.97759
R46343 a_31953_n19727.n6 a_31953_n19727.n242 0.97759
R46344 a_31953_n19727.n7 a_31953_n19727.n245 0.97759
R46345 a_31953_n19727.n8 a_31953_n19727.n243 0.97759
R46346 a_31953_n19727.n9 a_31953_n19727.n257 0.97759
R46347 a_31953_n19727.n11 a_31953_n19727.n255 0.97759
R46348 a_31953_n19727.n256 a_31953_n19727.n12 0.97759
R46349 a_31953_n19727.n13 a_31953_n19727.n254 0.97759
R46350 a_31953_n19727.n14 a_31953_n19727.n253 0.97759
R46351 a_31953_n19727.n15 a_31953_n19727.n251 0.97759
R46352 a_31953_n19727.n252 a_31953_n19727.n16 0.97759
R46353 a_31953_n19727.n17 a_31953_n19727.n250 0.97759
R46354 a_31953_n19727.n18 a_31953_n19727.n249 0.97759
R46355 a_31953_n19727.n20 a_31953_n19727.n247 0.97759
R46356 a_31953_n19727.n248 a_31953_n19727.n21 0.97759
R46357 a_31953_n19727.n22 a_31953_n19727.n246 0.97759
R46358 a_31953_n19727.n265 a_31953_n19727.n23 0.97759
R46359 a_31953_n19727.n24 a_31953_n19727.n263 0.97759
R46360 a_31953_n19727.n25 a_31953_n19727.n266 0.97759
R46361 a_31953_n19727.n26 a_31953_n19727.n264 0.97759
R46362 a_31953_n19727.n269 a_31953_n19727.n27 0.97759
R46363 a_31953_n19727.n28 a_31953_n19727.n267 0.97759
R46364 a_31953_n19727.n29 a_31953_n19727.n270 0.97759
R46365 a_31953_n19727.n31 a_31953_n19727.n268 0.97759
R46366 a_31953_n19727.n273 a_31953_n19727.n32 0.97759
R46367 a_31953_n19727.n33 a_31953_n19727.n271 0.97759
R46368 a_31953_n19727.n34 a_31953_n19727.n274 0.97759
R46369 a_31953_n19727.n35 a_31953_n19727.n272 0.97759
R46370 a_31953_n19727.n469 a_31953_n19727.n468 0.97759
R46371 a_31953_n19727.n470 a_31953_n19727.n466 0.97759
R46372 a_31953_n19727.n473 a_31953_n19727.n36 0.97759
R46373 a_31953_n19727.n37 a_31953_n19727.n471 0.97759
R46374 a_31953_n19727.n38 a_31953_n19727.n474 0.97759
R46375 a_31953_n19727.n40 a_31953_n19727.n472 0.97759
R46376 a_31953_n19727.n477 a_31953_n19727.n41 0.97759
R46377 a_31953_n19727.n42 a_31953_n19727.n475 0.97759
R46378 a_31953_n19727.n43 a_31953_n19727.n478 0.97759
R46379 a_31953_n19727.n44 a_31953_n19727.n476 0.97759
R46380 a_31953_n19727.n485 a_31953_n19727.n45 0.97759
R46381 a_31953_n19727.n46 a_31953_n19727.n483 0.97759
R46382 a_31953_n19727.n47 a_31953_n19727.n486 0.97759
R46383 a_31953_n19727.n49 a_31953_n19727.n484 0.97759
R46384 a_31953_n19727.n489 a_31953_n19727.n50 0.97759
R46385 a_31953_n19727.n51 a_31953_n19727.n487 0.97759
R46386 a_31953_n19727.n52 a_31953_n19727.n490 0.97759
R46387 a_31953_n19727.n54 a_31953_n19727.n488 0.97759
R46388 a_31953_n19727.n493 a_31953_n19727.n55 0.97759
R46389 a_31953_n19727.n56 a_31953_n19727.n491 0.97759
R46390 a_31953_n19727.n57 a_31953_n19727.n494 0.97759
R46391 a_31953_n19727.n58 a_31953_n19727.n492 0.97759
R46392 a_31953_n19727.n59 a_31953_n19727.n507 0.97759
R46393 a_31953_n19727.n61 a_31953_n19727.n505 0.97759
R46394 a_31953_n19727.n506 a_31953_n19727.n62 0.97759
R46395 a_31953_n19727.n63 a_31953_n19727.n504 0.97759
R46396 a_31953_n19727.n64 a_31953_n19727.n503 0.97759
R46397 a_31953_n19727.n65 a_31953_n19727.n501 0.97759
R46398 a_31953_n19727.n502 a_31953_n19727.n66 0.97759
R46399 a_31953_n19727.n67 a_31953_n19727.n500 0.97759
R46400 a_31953_n19727.n496 a_31953_n19727.n495 0.97759
R46401 a_31953_n19727.n68 a_31953_n19727.n499 0.97759
R46402 a_31953_n19727.n69 a_31953_n19727.n497 0.97759
R46403 a_31953_n19727.n70 a_31953_n19727.n498 0.97759
R46404 a_31953_n19727.n282 a_31953_n19727.n281 0.97759
R46405 a_31953_n19727.n283 a_31953_n19727.n279 0.97759
R46406 a_31953_n19727.n286 a_31953_n19727.n71 0.97759
R46407 a_31953_n19727.n72 a_31953_n19727.n284 0.97759
R46408 a_31953_n19727.n73 a_31953_n19727.n287 0.97759
R46409 a_31953_n19727.n75 a_31953_n19727.n285 0.97759
R46410 a_31953_n19727.n290 a_31953_n19727.n76 0.97759
R46411 a_31953_n19727.n77 a_31953_n19727.n288 0.97759
R46412 a_31953_n19727.n78 a_31953_n19727.n291 0.97759
R46413 a_31953_n19727.n79 a_31953_n19727.n289 0.97759
R46414 a_31953_n19727.n80 a_31953_n19727.n303 0.97759
R46415 a_31953_n19727.n82 a_31953_n19727.n301 0.97759
R46416 a_31953_n19727.n302 a_31953_n19727.n83 0.97759
R46417 a_31953_n19727.n84 a_31953_n19727.n300 0.97759
R46418 a_31953_n19727.n85 a_31953_n19727.n299 0.97759
R46419 a_31953_n19727.n86 a_31953_n19727.n297 0.97759
R46420 a_31953_n19727.n298 a_31953_n19727.n87 0.97759
R46421 a_31953_n19727.n88 a_31953_n19727.n296 0.97759
R46422 a_31953_n19727.n89 a_31953_n19727.n295 0.97759
R46423 a_31953_n19727.n91 a_31953_n19727.n293 0.97759
R46424 a_31953_n19727.n294 a_31953_n19727.n92 0.97759
R46425 a_31953_n19727.n93 a_31953_n19727.n292 0.97759
R46426 a_31953_n19727.n311 a_31953_n19727.n94 0.97759
R46427 a_31953_n19727.n95 a_31953_n19727.n309 0.97759
R46428 a_31953_n19727.n96 a_31953_n19727.n312 0.97759
R46429 a_31953_n19727.n97 a_31953_n19727.n310 0.97759
R46430 a_31953_n19727.n315 a_31953_n19727.n98 0.97759
R46431 a_31953_n19727.n99 a_31953_n19727.n313 0.97759
R46432 a_31953_n19727.n100 a_31953_n19727.n316 0.97759
R46433 a_31953_n19727.n102 a_31953_n19727.n314 0.97759
R46434 a_31953_n19727.n319 a_31953_n19727.n103 0.97759
R46435 a_31953_n19727.n104 a_31953_n19727.n317 0.97759
R46436 a_31953_n19727.n105 a_31953_n19727.n320 0.97759
R46437 a_31953_n19727.n106 a_31953_n19727.n318 0.97759
R46438 a_31953_n19727.n367 a_31953_n19727.n366 0.97759
R46439 a_31953_n19727.n368 a_31953_n19727.n364 0.97759
R46440 a_31953_n19727.n107 a_31953_n19727.n362 0.97759
R46441 a_31953_n19727.n109 a_31953_n19727.n360 0.97759
R46442 a_31953_n19727.n361 a_31953_n19727.n110 0.97759
R46443 a_31953_n19727.n111 a_31953_n19727.n359 0.97759
R46444 a_31953_n19727.n112 a_31953_n19727.n358 0.97759
R46445 a_31953_n19727.n114 a_31953_n19727.n356 0.97759
R46446 a_31953_n19727.n357 a_31953_n19727.n115 0.97759
R46447 a_31953_n19727.n116 a_31953_n19727.n355 0.97759
R46448 a_31953_n19727.n327 a_31953_n19727.n117 0.97759
R46449 a_31953_n19727.n118 a_31953_n19727.n325 0.97759
R46450 a_31953_n19727.n119 a_31953_n19727.n328 0.97759
R46451 a_31953_n19727.n120 a_31953_n19727.n326 0.97759
R46452 a_31953_n19727.n331 a_31953_n19727.n121 0.97759
R46453 a_31953_n19727.n122 a_31953_n19727.n329 0.97759
R46454 a_31953_n19727.n123 a_31953_n19727.n332 0.97759
R46455 a_31953_n19727.n125 a_31953_n19727.n330 0.97759
R46456 a_31953_n19727.n335 a_31953_n19727.n126 0.97759
R46457 a_31953_n19727.n127 a_31953_n19727.n333 0.97759
R46458 a_31953_n19727.n128 a_31953_n19727.n336 0.97759
R46459 a_31953_n19727.n129 a_31953_n19727.n334 0.97759
R46460 a_31953_n19727.n130 a_31953_n19727.n349 0.97759
R46461 a_31953_n19727.n132 a_31953_n19727.n347 0.97759
R46462 a_31953_n19727.n348 a_31953_n19727.n133 0.97759
R46463 a_31953_n19727.n134 a_31953_n19727.n346 0.97759
R46464 a_31953_n19727.n135 a_31953_n19727.n345 0.97759
R46465 a_31953_n19727.n136 a_31953_n19727.n343 0.97759
R46466 a_31953_n19727.n344 a_31953_n19727.n137 0.97759
R46467 a_31953_n19727.n138 a_31953_n19727.n342 0.97759
R46468 a_31953_n19727.n338 a_31953_n19727.n337 0.97759
R46469 a_31953_n19727.n139 a_31953_n19727.n341 0.97759
R46470 a_31953_n19727.n140 a_31953_n19727.n339 0.97759
R46471 a_31953_n19727.n141 a_31953_n19727.n340 0.97759
R46472 a_31953_n19727.n376 a_31953_n19727.n375 0.97759
R46473 a_31953_n19727.n377 a_31953_n19727.n373 0.97759
R46474 a_31953_n19727.n380 a_31953_n19727.n142 0.97759
R46475 a_31953_n19727.n143 a_31953_n19727.n378 0.97759
R46476 a_31953_n19727.n144 a_31953_n19727.n381 0.97759
R46477 a_31953_n19727.n146 a_31953_n19727.n379 0.97759
R46478 a_31953_n19727.n384 a_31953_n19727.n147 0.97759
R46479 a_31953_n19727.n148 a_31953_n19727.n382 0.97759
R46480 a_31953_n19727.n149 a_31953_n19727.n385 0.97759
R46481 a_31953_n19727.n150 a_31953_n19727.n383 0.97759
R46482 a_31953_n19727.n151 a_31953_n19727.n397 0.97759
R46483 a_31953_n19727.n153 a_31953_n19727.n395 0.97759
R46484 a_31953_n19727.n396 a_31953_n19727.n154 0.97759
R46485 a_31953_n19727.n155 a_31953_n19727.n394 0.97759
R46486 a_31953_n19727.n156 a_31953_n19727.n393 0.97759
R46487 a_31953_n19727.n157 a_31953_n19727.n391 0.97759
R46488 a_31953_n19727.n392 a_31953_n19727.n158 0.97759
R46489 a_31953_n19727.n159 a_31953_n19727.n390 0.97759
R46490 a_31953_n19727.n160 a_31953_n19727.n389 0.97759
R46491 a_31953_n19727.n162 a_31953_n19727.n387 0.97759
R46492 a_31953_n19727.n388 a_31953_n19727.n163 0.97759
R46493 a_31953_n19727.n164 a_31953_n19727.n386 0.97759
R46494 a_31953_n19727.n405 a_31953_n19727.n165 0.97759
R46495 a_31953_n19727.n166 a_31953_n19727.n403 0.97759
R46496 a_31953_n19727.n167 a_31953_n19727.n406 0.97759
R46497 a_31953_n19727.n168 a_31953_n19727.n404 0.97759
R46498 a_31953_n19727.n409 a_31953_n19727.n169 0.97759
R46499 a_31953_n19727.n170 a_31953_n19727.n407 0.97759
R46500 a_31953_n19727.n171 a_31953_n19727.n410 0.97759
R46501 a_31953_n19727.n173 a_31953_n19727.n408 0.97759
R46502 a_31953_n19727.n413 a_31953_n19727.n174 0.97759
R46503 a_31953_n19727.n175 a_31953_n19727.n411 0.97759
R46504 a_31953_n19727.n176 a_31953_n19727.n414 0.97759
R46505 a_31953_n19727.n177 a_31953_n19727.n412 0.97759
R46506 a_31953_n19727.n460 a_31953_n19727.n459 0.97759
R46507 a_31953_n19727.n461 a_31953_n19727.n457 0.97759
R46508 a_31953_n19727.n178 a_31953_n19727.n455 0.97759
R46509 a_31953_n19727.n180 a_31953_n19727.n453 0.97759
R46510 a_31953_n19727.n454 a_31953_n19727.n181 0.97759
R46511 a_31953_n19727.n182 a_31953_n19727.n452 0.97759
R46512 a_31953_n19727.n183 a_31953_n19727.n451 0.97759
R46513 a_31953_n19727.n185 a_31953_n19727.n449 0.97759
R46514 a_31953_n19727.n450 a_31953_n19727.n186 0.97759
R46515 a_31953_n19727.n187 a_31953_n19727.n448 0.97759
R46516 a_31953_n19727.n420 a_31953_n19727.n188 0.97759
R46517 a_31953_n19727.n189 a_31953_n19727.n418 0.97759
R46518 a_31953_n19727.n190 a_31953_n19727.n421 0.97759
R46519 a_31953_n19727.n191 a_31953_n19727.n419 0.97759
R46520 a_31953_n19727.n424 a_31953_n19727.n192 0.97759
R46521 a_31953_n19727.n193 a_31953_n19727.n422 0.97759
R46522 a_31953_n19727.n194 a_31953_n19727.n425 0.97759
R46523 a_31953_n19727.n196 a_31953_n19727.n423 0.97759
R46524 a_31953_n19727.n428 a_31953_n19727.n197 0.97759
R46525 a_31953_n19727.n198 a_31953_n19727.n426 0.97759
R46526 a_31953_n19727.n199 a_31953_n19727.n429 0.97759
R46527 a_31953_n19727.n200 a_31953_n19727.n427 0.97759
R46528 a_31953_n19727.n201 a_31953_n19727.n442 0.97759
R46529 a_31953_n19727.n203 a_31953_n19727.n440 0.97759
R46530 a_31953_n19727.n441 a_31953_n19727.n204 0.97759
R46531 a_31953_n19727.n205 a_31953_n19727.n439 0.97759
R46532 a_31953_n19727.n206 a_31953_n19727.n438 0.97759
R46533 a_31953_n19727.n207 a_31953_n19727.n436 0.97759
R46534 a_31953_n19727.n437 a_31953_n19727.n208 0.97759
R46535 a_31953_n19727.n209 a_31953_n19727.n435 0.97759
R46536 a_31953_n19727.n431 a_31953_n19727.n430 0.97759
R46537 a_31953_n19727.n210 a_31953_n19727.n434 0.97759
R46538 a_31953_n19727.n211 a_31953_n19727.n432 0.97759
R46539 a_31953_n19727.n212 a_31953_n19727.n433 0.97759
R46540 a_31953_n19727.n234 a_31953_n19727.n213 0.931516
R46541 a_31953_n19727.n214 a_31953_n19727.n232 0.931516
R46542 a_31953_n19727.n467 a_31953_n19727.n215 0.931516
R46543 a_31953_n19727.n216 a_31953_n19727.n465 0.931516
R46544 a_31953_n19727.n280 a_31953_n19727.n217 0.931516
R46545 a_31953_n19727.n218 a_31953_n19727.n278 0.931516
R46546 a_31953_n19727.n365 a_31953_n19727.n219 0.931516
R46547 a_31953_n19727.n220 a_31953_n19727.n363 0.931516
R46548 a_31953_n19727.n374 a_31953_n19727.n221 0.931516
R46549 a_31953_n19727.n222 a_31953_n19727.n372 0.931516
R46550 a_31953_n19727.n458 a_31953_n19727.n223 0.931516
R46551 a_31953_n19727.n224 a_31953_n19727.n456 0.931516
R46552 a_31953_n19727.n74 a_31953_n19727.n81 0.82023
R46553 a_31953_n19727.n145 a_31953_n19727.n152 0.82023
R46554 a_31953_n19727.n3 a_31953_n19727.n10 0.82023
R46555 a_31953_n19727.n131 a_31953_n19727.n124 0.818405
R46556 a_31953_n19727.n202 a_31953_n19727.n195 0.818405
R46557 a_31953_n19727.n60 a_31953_n19727.n53 0.818405
R46558 a_31953_n19727.n463 a_31953_n19727.n462 0.7505
R46559 a_31953_n19727.n462 a_31953_n19727.n172 0.717155
R46560 a_31953_n19727.n464 a_31953_n19727.n30 0.717155
R46561 a_31953_n19727.n226 a_31953_n19727.n101 0.711725
R46562 a_31953_n19727.n108 a_31953_n19727.n113 0.639622
R46563 a_31953_n19727.n179 a_31953_n19727.n184 0.639622
R46564 a_31953_n19727.n48 a_31953_n19727.n39 0.639622
R46565 a_31953_n19727.n237 a_31953_n19727.n236 0.62434
R46566 a_31953_n19727.n470 a_31953_n19727.n469 0.62434
R46567 a_31953_n19727.n283 a_31953_n19727.n282 0.62434
R46568 a_31953_n19727.n368 a_31953_n19727.n367 0.62434
R46569 a_31953_n19727.n377 a_31953_n19727.n376 0.62434
R46570 a_31953_n19727.n461 a_31953_n19727.n460 0.62434
R46571 a_31953_n19727.n212 a_31953_n19727.n211 0.62434
R46572 a_31953_n19727.n430 a_31953_n19727.n210 0.62434
R46573 a_31953_n19727.n209 a_31953_n19727.n208 0.62434
R46574 a_31953_n19727.n207 a_31953_n19727.n206 0.62434
R46575 a_31953_n19727.n205 a_31953_n19727.n204 0.62434
R46576 a_31953_n19727.n203 a_31953_n19727.n201 0.62434
R46577 a_31953_n19727.n200 a_31953_n19727.n199 0.62434
R46578 a_31953_n19727.n198 a_31953_n19727.n197 0.62434
R46579 a_31953_n19727.n196 a_31953_n19727.n194 0.62434
R46580 a_31953_n19727.n193 a_31953_n19727.n192 0.62434
R46581 a_31953_n19727.n191 a_31953_n19727.n190 0.62434
R46582 a_31953_n19727.n189 a_31953_n19727.n188 0.62434
R46583 a_31953_n19727.n187 a_31953_n19727.n186 0.62434
R46584 a_31953_n19727.n185 a_31953_n19727.n183 0.62434
R46585 a_31953_n19727.n182 a_31953_n19727.n181 0.62434
R46586 a_31953_n19727.n180 a_31953_n19727.n178 0.62434
R46587 a_31953_n19727.n177 a_31953_n19727.n176 0.62434
R46588 a_31953_n19727.n175 a_31953_n19727.n174 0.62434
R46589 a_31953_n19727.n173 a_31953_n19727.n171 0.62434
R46590 a_31953_n19727.n170 a_31953_n19727.n169 0.62434
R46591 a_31953_n19727.n168 a_31953_n19727.n167 0.62434
R46592 a_31953_n19727.n166 a_31953_n19727.n165 0.62434
R46593 a_31953_n19727.n164 a_31953_n19727.n163 0.62434
R46594 a_31953_n19727.n162 a_31953_n19727.n160 0.62434
R46595 a_31953_n19727.n159 a_31953_n19727.n158 0.62434
R46596 a_31953_n19727.n157 a_31953_n19727.n156 0.62434
R46597 a_31953_n19727.n155 a_31953_n19727.n154 0.62434
R46598 a_31953_n19727.n153 a_31953_n19727.n151 0.62434
R46599 a_31953_n19727.n150 a_31953_n19727.n149 0.62434
R46600 a_31953_n19727.n148 a_31953_n19727.n147 0.62434
R46601 a_31953_n19727.n146 a_31953_n19727.n144 0.62434
R46602 a_31953_n19727.n143 a_31953_n19727.n142 0.62434
R46603 a_31953_n19727.n141 a_31953_n19727.n140 0.62434
R46604 a_31953_n19727.n337 a_31953_n19727.n139 0.62434
R46605 a_31953_n19727.n138 a_31953_n19727.n137 0.62434
R46606 a_31953_n19727.n136 a_31953_n19727.n135 0.62434
R46607 a_31953_n19727.n134 a_31953_n19727.n133 0.62434
R46608 a_31953_n19727.n132 a_31953_n19727.n130 0.62434
R46609 a_31953_n19727.n129 a_31953_n19727.n128 0.62434
R46610 a_31953_n19727.n127 a_31953_n19727.n126 0.62434
R46611 a_31953_n19727.n125 a_31953_n19727.n123 0.62434
R46612 a_31953_n19727.n122 a_31953_n19727.n121 0.62434
R46613 a_31953_n19727.n120 a_31953_n19727.n119 0.62434
R46614 a_31953_n19727.n118 a_31953_n19727.n117 0.62434
R46615 a_31953_n19727.n116 a_31953_n19727.n115 0.62434
R46616 a_31953_n19727.n114 a_31953_n19727.n112 0.62434
R46617 a_31953_n19727.n111 a_31953_n19727.n110 0.62434
R46618 a_31953_n19727.n109 a_31953_n19727.n107 0.62434
R46619 a_31953_n19727.n106 a_31953_n19727.n105 0.62434
R46620 a_31953_n19727.n104 a_31953_n19727.n103 0.62434
R46621 a_31953_n19727.n102 a_31953_n19727.n100 0.62434
R46622 a_31953_n19727.n99 a_31953_n19727.n98 0.62434
R46623 a_31953_n19727.n97 a_31953_n19727.n96 0.62434
R46624 a_31953_n19727.n95 a_31953_n19727.n94 0.62434
R46625 a_31953_n19727.n93 a_31953_n19727.n92 0.62434
R46626 a_31953_n19727.n91 a_31953_n19727.n89 0.62434
R46627 a_31953_n19727.n88 a_31953_n19727.n87 0.62434
R46628 a_31953_n19727.n86 a_31953_n19727.n85 0.62434
R46629 a_31953_n19727.n84 a_31953_n19727.n83 0.62434
R46630 a_31953_n19727.n82 a_31953_n19727.n80 0.62434
R46631 a_31953_n19727.n79 a_31953_n19727.n78 0.62434
R46632 a_31953_n19727.n77 a_31953_n19727.n76 0.62434
R46633 a_31953_n19727.n75 a_31953_n19727.n73 0.62434
R46634 a_31953_n19727.n72 a_31953_n19727.n71 0.62434
R46635 a_31953_n19727.n70 a_31953_n19727.n69 0.62434
R46636 a_31953_n19727.n495 a_31953_n19727.n68 0.62434
R46637 a_31953_n19727.n67 a_31953_n19727.n66 0.62434
R46638 a_31953_n19727.n65 a_31953_n19727.n64 0.62434
R46639 a_31953_n19727.n63 a_31953_n19727.n62 0.62434
R46640 a_31953_n19727.n61 a_31953_n19727.n59 0.62434
R46641 a_31953_n19727.n58 a_31953_n19727.n57 0.62434
R46642 a_31953_n19727.n56 a_31953_n19727.n55 0.62434
R46643 a_31953_n19727.n54 a_31953_n19727.n52 0.62434
R46644 a_31953_n19727.n51 a_31953_n19727.n50 0.62434
R46645 a_31953_n19727.n49 a_31953_n19727.n47 0.62434
R46646 a_31953_n19727.n46 a_31953_n19727.n45 0.62434
R46647 a_31953_n19727.n44 a_31953_n19727.n43 0.62434
R46648 a_31953_n19727.n42 a_31953_n19727.n41 0.62434
R46649 a_31953_n19727.n40 a_31953_n19727.n38 0.62434
R46650 a_31953_n19727.n37 a_31953_n19727.n36 0.62434
R46651 a_31953_n19727.n35 a_31953_n19727.n34 0.62434
R46652 a_31953_n19727.n33 a_31953_n19727.n32 0.62434
R46653 a_31953_n19727.n31 a_31953_n19727.n29 0.62434
R46654 a_31953_n19727.n28 a_31953_n19727.n27 0.62434
R46655 a_31953_n19727.n26 a_31953_n19727.n25 0.62434
R46656 a_31953_n19727.n24 a_31953_n19727.n23 0.62434
R46657 a_31953_n19727.n22 a_31953_n19727.n21 0.62434
R46658 a_31953_n19727.n20 a_31953_n19727.n18 0.62434
R46659 a_31953_n19727.n17 a_31953_n19727.n16 0.62434
R46660 a_31953_n19727.n15 a_31953_n19727.n14 0.62434
R46661 a_31953_n19727.n13 a_31953_n19727.n12 0.62434
R46662 a_31953_n19727.n11 a_31953_n19727.n9 0.62434
R46663 a_31953_n19727.n8 a_31953_n19727.n7 0.62434
R46664 a_31953_n19727.n6 a_31953_n19727.n5 0.62434
R46665 a_31953_n19727.n4 a_31953_n19727.n2 0.62434
R46666 a_31953_n19727.n1 a_31953_n19727.n0 0.62434
R46667 a_31953_n19727.n462 a_31953_n19727.n179 0.617426
R46668 a_31953_n19727.n39 a_31953_n19727.n464 0.617426
R46669 a_31953_n19727.n225 a_31953_n19727.n108 0.604351
R46670 a_31953_n19727.n224 a_31953_n19727.n223 0.595087
R46671 a_31953_n19727.n222 a_31953_n19727.n221 0.595087
R46672 a_31953_n19727.n220 a_31953_n19727.n219 0.595087
R46673 a_31953_n19727.n218 a_31953_n19727.n217 0.595087
R46674 a_31953_n19727.n216 a_31953_n19727.n215 0.595087
R46675 a_31953_n19727.n214 a_31953_n19727.n213 0.595087
R46676 a_31953_n19727.n124 a_31953_n19727.n113 0.545973
R46677 a_31953_n19727.n195 a_31953_n19727.n184 0.545973
R46678 a_31953_n19727.n53 a_31953_n19727.n48 0.545973
R46679 a_31953_n19727.n81 a_31953_n19727.n90 0.545365
R46680 a_31953_n19727.n152 a_31953_n19727.n161 0.545365
R46681 a_31953_n19727.n10 a_31953_n19727.n19 0.545365
R46682 a_31953_n19727.n30 a_31953_n19727.n19 0.452324
R46683 a_31953_n19727.n172 a_31953_n19727.n161 0.452324
R46684 a_31953_n19727.n101 a_31953_n19727.n90 0.452324
R46685 a_31699_20742.n388 a_31699_20742.n313 16.7377
R46686 a_31699_20742.n314 a_31699_20742.t1 10.214
R46687 a_31699_20742.n324 a_31699_20742.t131 10.214
R46688 a_31699_20742.n335 a_31699_20742.t220 10.214
R46689 a_31699_20742.n346 a_31699_20742.t60 10.214
R46690 a_31699_20742.n356 a_31699_20742.t141 10.214
R46691 a_31699_20742.n320 a_31699_20742.t27 10.2117
R46692 a_31699_20742.n330 a_31699_20742.t213 10.2117
R46693 a_31699_20742.n341 a_31699_20742.t81 10.2117
R46694 a_31699_20742.n352 a_31699_20742.t143 10.2117
R46695 a_31699_20742.n362 a_31699_20742.t224 10.2117
R46696 a_31699_20742.n317 a_31699_20742.t185 9.58832
R46697 a_31699_20742.n327 a_31699_20742.t52 9.58832
R46698 a_31699_20742.n338 a_31699_20742.t23 9.58832
R46699 a_31699_20742.n370 a_31699_20742.t144 9.58832
R46700 a_31699_20742.n349 a_31699_20742.t17 9.58832
R46701 a_31699_20742.n359 a_31699_20742.t62 9.58832
R46702 a_31699_20742.n319 a_31699_20742.t89 9.58085
R46703 a_31699_20742.n329 a_31699_20742.t172 9.58085
R46704 a_31699_20742.n340 a_31699_20742.t3 9.58085
R46705 a_31699_20742.n372 a_31699_20742.t45 9.58085
R46706 a_31699_20742.n351 a_31699_20742.t29 9.58085
R46707 a_31699_20742.n361 a_31699_20742.t184 9.58085
R46708 a_31699_20742.n318 a_31699_20742.t256 9.58045
R46709 a_31699_20742.n316 a_31699_20742.t37 9.58045
R46710 a_31699_20742.n315 a_31699_20742.t7 9.58045
R46711 a_31699_20742.n328 a_31699_20742.t127 9.58045
R46712 a_31699_20742.n326 a_31699_20742.t153 9.58045
R46713 a_31699_20742.n325 a_31699_20742.t108 9.58045
R46714 a_31699_20742.n339 a_31699_20742.t13 9.58045
R46715 a_31699_20742.n337 a_31699_20742.t244 9.58045
R46716 a_31699_20742.n336 a_31699_20742.t199 9.58045
R46717 a_31699_20742.n371 a_31699_20742.t219 9.58045
R46718 a_31699_20742.n350 a_31699_20742.t39 9.58045
R46719 a_31699_20742.n348 a_31699_20742.t85 9.58045
R46720 a_31699_20742.n347 a_31699_20742.t255 9.58045
R46721 a_31699_20742.n360 a_31699_20742.t134 9.58045
R46722 a_31699_20742.n358 a_31699_20742.t164 9.58045
R46723 a_31699_20742.n357 a_31699_20742.t118 9.58045
R46724 a_31699_20742.n314 a_31699_20742.t33 9.58005
R46725 a_31699_20742.n324 a_31699_20742.t180 9.58005
R46726 a_31699_20742.n335 a_31699_20742.t46 9.58005
R46727 a_31699_20742.n346 a_31699_20742.t111 9.58005
R46728 a_31699_20742.n356 a_31699_20742.t192 9.58005
R46729 a_31699_20742.n320 a_31699_20742.t41 9.57886
R46730 a_31699_20742.n321 a_31699_20742.t15 9.57886
R46731 a_31699_20742.n322 a_31699_20742.t25 9.57886
R46732 a_31699_20742.n330 a_31699_20742.t138 9.57886
R46733 a_31699_20742.n331 a_31699_20742.t72 9.57886
R46734 a_31699_20742.n332 a_31699_20742.t218 9.57886
R46735 a_31699_20742.n341 a_31699_20742.t234 9.57886
R46736 a_31699_20742.n342 a_31699_20742.t163 9.57886
R46737 a_31699_20742.n343 a_31699_20742.t92 9.57886
R46738 a_31699_20742.n352 a_31699_20742.t71 9.57886
R46739 a_31699_20742.n353 a_31699_20742.t226 9.57886
R46740 a_31699_20742.n354 a_31699_20742.t150 9.57886
R46741 a_31699_20742.n362 a_31699_20742.t149 9.57886
R46742 a_31699_20742.n363 a_31699_20742.t82 9.57886
R46743 a_31699_20742.n364 a_31699_20742.t235 9.57886
R46744 a_31699_20742.n376 a_31699_20742.t35 8.38951
R46745 a_31699_20742.n389 a_31699_20742.t0 8.38805
R46746 a_31699_20742.n367 a_31699_20742.t11 8.38752
R46747 a_31699_20742.n268 a_31699_20742.t142 8.38704
R46748 a_31699_20742.n262 a_31699_20742.t207 8.38704
R46749 a_31699_20742.n211 a_31699_20742.t242 8.46135
R46750 a_31699_20742.n213 a_31699_20742.t148 8.46135
R46751 a_31699_20742.n193 a_31699_20742.t69 8.48081
R46752 a_31699_20742.n188 a_31699_20742.t228 8.48081
R46753 a_31699_20742.n168 a_31699_20742.t156 8.10567
R46754 a_31699_20742.n130 a_31699_20742.t51 8.10567
R46755 a_31699_20742.n130 a_31699_20742.t223 8.10567
R46756 a_31699_20742.n131 a_31699_20742.t147 8.10567
R46757 a_31699_20742.n131 a_31699_20742.t222 8.10567
R46758 a_31699_20742.n113 a_31699_20742.t87 8.10567
R46759 a_31699_20742.n113 a_31699_20742.t237 8.10567
R46760 a_31699_20742.n127 a_31699_20742.t162 8.10567
R46761 a_31699_20742.n127 a_31699_20742.t94 8.10567
R46762 a_31699_20742.n110 a_31699_20742.t70 8.10567
R46763 a_31699_20742.n110 a_31699_20742.t217 8.10567
R46764 a_31699_20742.n124 a_31699_20742.t166 8.10567
R46765 a_31699_20742.n124 a_31699_20742.t75 8.10567
R46766 a_31699_20742.n173 a_31699_20742.t73 8.10567
R46767 a_31699_20742.n173 a_31699_20742.t201 8.10567
R46768 a_31699_20742.n219 a_31699_20742.t128 8.10567
R46769 a_31699_20742.n176 a_31699_20742.t124 8.10567
R46770 a_31699_20742.n176 a_31699_20742.t221 8.10567
R46771 a_31699_20742.n175 a_31699_20742.t146 8.10567
R46772 a_31699_20742.n168 a_31699_20742.t90 8.10567
R46773 a_31699_20742.n136 a_31699_20742.t238 8.10567
R46774 a_31699_20742.n136 a_31699_20742.t187 8.10567
R46775 a_31699_20742.n90 a_31699_20742.t145 8.10567
R46776 a_31699_20742.n158 a_31699_20742.t258 8.10567
R46777 a_31699_20742.n158 a_31699_20742.t216 8.10567
R46778 a_31699_20742.n159 a_31699_20742.t139 8.10567
R46779 a_31699_20742.n159 a_31699_20742.t214 8.10567
R46780 a_31699_20742.n83 a_31699_20742.t76 8.10567
R46781 a_31699_20742.n83 a_31699_20742.t227 8.10567
R46782 a_31699_20742.n162 a_31699_20742.t151 8.10567
R46783 a_31699_20742.n162 a_31699_20742.t84 8.10567
R46784 a_31699_20742.n87 a_31699_20742.t59 8.10567
R46785 a_31699_20742.n87 a_31699_20742.t209 8.10567
R46786 a_31699_20742.n86 a_31699_20742.t161 8.10567
R46787 a_31699_20742.n86 a_31699_20742.t66 8.10567
R46788 a_31699_20742.n198 a_31699_20742.t247 8.10567
R46789 a_31699_20742.n198 a_31699_20742.t154 8.10567
R46790 a_31699_20742.n226 a_31699_20742.t78 8.10567
R46791 a_31699_20742.n201 a_31699_20742.t74 8.10567
R46792 a_31699_20742.n201 a_31699_20742.t174 8.10567
R46793 a_31699_20742.n200 a_31699_20742.t100 8.10567
R46794 a_31699_20742.n90 a_31699_20742.t77 8.10567
R46795 a_31699_20742.n90 a_31699_20742.t230 8.10567
R46796 a_31699_20742.n90 a_31699_20742.t181 8.10567
R46797 a_31699_20742.n165 a_31699_20742.t93 8.10567
R46798 a_31699_20742.n120 a_31699_20742.t205 8.10567
R46799 a_31699_20742.n120 a_31699_20742.t159 8.10567
R46800 a_31699_20742.n121 a_31699_20742.t86 8.10567
R46801 a_31699_20742.n121 a_31699_20742.t158 8.10567
R46802 a_31699_20742.n107 a_31699_20742.t243 8.10567
R46803 a_31699_20742.n107 a_31699_20742.t168 8.10567
R46804 a_31699_20742.n106 a_31699_20742.t97 8.10567
R46805 a_31699_20742.n106 a_31699_20742.t249 8.10567
R46806 a_31699_20742.n103 a_31699_20742.t229 8.10567
R46807 a_31699_20742.n103 a_31699_20742.t152 8.10567
R46808 a_31699_20742.n102 a_31699_20742.t106 8.10567
R46809 a_31699_20742.n102 a_31699_20742.t236 8.10567
R46810 a_31699_20742.n179 a_31699_20742.t233 8.10567
R46811 a_31699_20742.n179 a_31699_20742.t136 8.10567
R46812 a_31699_20742.n178 a_31699_20742.t63 8.10567
R46813 a_31699_20742.n182 a_31699_20742.t56 8.10567
R46814 a_31699_20742.n182 a_31699_20742.t157 8.10567
R46815 a_31699_20742.n181 a_31699_20742.t83 8.10567
R46816 a_31699_20742.n165 a_31699_20742.t245 8.10567
R46817 a_31699_20742.n134 a_31699_20742.t170 8.10567
R46818 a_31699_20742.n134 a_31699_20742.t125 8.10567
R46819 a_31699_20742.n100 a_31699_20742.t54 8.10567
R46820 a_31699_20742.n214 a_31699_20742.t167 8.10567
R46821 a_31699_20742.n214 a_31699_20742.t123 8.10567
R46822 a_31699_20742.n153 a_31699_20742.t49 8.10567
R46823 a_31699_20742.n153 a_31699_20742.t122 8.10567
R46824 a_31699_20742.n93 a_31699_20742.t206 8.10567
R46825 a_31699_20742.n93 a_31699_20742.t133 8.10567
R46826 a_31699_20742.n92 a_31699_20742.t57 8.10567
R46827 a_31699_20742.n92 a_31699_20742.t215 8.10567
R46828 a_31699_20742.n97 a_31699_20742.t193 8.10567
R46829 a_31699_20742.n97 a_31699_20742.t117 8.10567
R46830 a_31699_20742.n96 a_31699_20742.t68 8.10567
R46831 a_31699_20742.n96 a_31699_20742.t200 8.10567
R46832 a_31699_20742.n204 a_31699_20742.t155 8.10567
R46833 a_31699_20742.n204 a_31699_20742.t61 8.10567
R46834 a_31699_20742.n203 a_31699_20742.t211 8.10567
R46835 a_31699_20742.n206 a_31699_20742.t203 8.10567
R46836 a_31699_20742.n206 a_31699_20742.t80 8.10567
R46837 a_31699_20742.n230 a_31699_20742.t232 8.10567
R46838 a_31699_20742.n100 a_31699_20742.t210 8.10567
R46839 a_31699_20742.n100 a_31699_20742.t135 8.10567
R46840 a_31699_20742.n100 a_31699_20742.t88 8.10567
R46841 a_31699_20742.n49 a_31699_20742.t107 8.10567
R46842 a_31699_20742.n47 a_31699_20742.t252 8.10567
R46843 a_31699_20742.n45 a_31699_20742.t182 8.10567
R46844 a_31699_20742.n260 a_31699_20742.t113 8.10567
R46845 a_31699_20742.n307 a_31699_20742.t53 8.10567
R46846 a_31699_20742.n306 a_31699_20742.t183 8.10567
R46847 a_31699_20742.n305 a_31699_20742.t110 8.10567
R46848 a_31699_20742.n192 a_31699_20742.t241 8.10567
R46849 a_31699_20742.n43 a_31699_20742.t165 8.10567
R46850 a_31699_20742.n41 a_31699_20742.t240 8.10567
R46851 a_31699_20742.n59 a_31699_20742.t176 8.10567
R46852 a_31699_20742.n57 a_31699_20742.t109 8.10567
R46853 a_31699_20742.n261 a_31699_20742.t253 8.10567
R46854 a_31699_20742.n301 a_31699_20742.t104 8.10567
R46855 a_31699_20742.n300 a_31699_20742.t202 8.10567
R46856 a_31699_20742.n299 a_31699_20742.t130 8.10567
R46857 a_31699_20742.n190 a_31699_20742.t91 8.10567
R46858 a_31699_20742.n55 a_31699_20742.t239 8.10567
R46859 a_31699_20742.n53 a_31699_20742.t188 8.10567
R46860 a_31699_20742.n52 a_31699_20742.t96 8.10567
R46861 a_31699_20742.n0 a_31699_20742.t55 8.10567
R46862 a_31699_20742.n1 a_31699_20742.t204 8.10567
R46863 a_31699_20742.n18 a_31699_20742.t132 8.10567
R46864 a_31699_20742.n144 a_31699_20742.t65 8.10567
R46865 a_31699_20742.n279 a_31699_20742.t264 8.10567
R46866 a_31699_20742.n278 a_31699_20742.t173 8.10567
R46867 a_31699_20742.n277 a_31699_20742.t99 8.10567
R46868 a_31699_20742.n210 a_31699_20742.t198 8.10567
R46869 a_31699_20742.n16 a_31699_20742.t121 8.10567
R46870 a_31699_20742.n28 a_31699_20742.t196 8.10567
R46871 a_31699_20742.n37 a_31699_20742.t129 8.10567
R46872 a_31699_20742.n5 a_31699_20742.t58 8.10567
R46873 a_31699_20742.n141 a_31699_20742.t208 8.10567
R46874 a_31699_20742.n276 a_31699_20742.t95 8.10567
R46875 a_31699_20742.n275 a_31699_20742.t195 8.10567
R46876 a_31699_20742.n274 a_31699_20742.t120 8.10567
R46877 a_31699_20742.n147 a_31699_20742.t260 8.10567
R46878 a_31699_20742.n3 a_31699_20742.t189 8.10567
R46879 a_31699_20742.n20 a_31699_20742.t140 8.10567
R46880 a_31699_20742.n30 a_31699_20742.t47 8.10567
R46881 a_31699_20742.n69 a_31699_20742.t261 8.10567
R46882 a_31699_20742.n67 a_31699_20742.t190 8.10567
R46883 a_31699_20742.n65 a_31699_20742.t115 8.10567
R46884 a_31699_20742.n286 a_31699_20742.t48 8.10567
R46885 a_31699_20742.n282 a_31699_20742.t212 8.10567
R46886 a_31699_20742.n283 a_31699_20742.t119 8.10567
R46887 a_31699_20742.n284 a_31699_20742.t263 8.10567
R46888 a_31699_20742.n189 a_31699_20742.t179 8.10567
R46889 a_31699_20742.n63 a_31699_20742.t105 8.10567
R46890 a_31699_20742.n61 a_31699_20742.t177 8.10567
R46891 a_31699_20742.n79 a_31699_20742.t112 8.10567
R46892 a_31699_20742.n77 a_31699_20742.t262 8.10567
R46893 a_31699_20742.n267 a_31699_20742.t194 8.10567
R46894 a_31699_20742.n272 a_31699_20742.t257 8.10567
R46895 a_31699_20742.n271 a_31699_20742.t137 8.10567
R46896 a_31699_20742.n270 a_31699_20742.t64 8.10567
R46897 a_31699_20742.n186 a_31699_20742.t246 8.10567
R46898 a_31699_20742.n75 a_31699_20742.t171 8.10567
R46899 a_31699_20742.n73 a_31699_20742.t126 8.10567
R46900 a_31699_20742.n71 a_31699_20742.t251 8.10567
R46901 a_31699_20742.n7 a_31699_20742.t186 8.10567
R46902 a_31699_20742.n8 a_31699_20742.t114 8.10567
R46903 a_31699_20742.n24 a_31699_20742.t259 8.10567
R46904 a_31699_20742.n142 a_31699_20742.t197 8.10567
R46905 a_31699_20742.n293 a_31699_20742.t175 8.10567
R46906 a_31699_20742.n294 a_31699_20742.t79 8.10567
R46907 a_31699_20742.n295 a_31699_20742.t231 8.10567
R46908 a_31699_20742.n212 a_31699_20742.t103 8.10567
R46909 a_31699_20742.n22 a_31699_20742.t250 8.10567
R46910 a_31699_20742.n32 a_31699_20742.t102 8.10567
R46911 a_31699_20742.n13 a_31699_20742.t254 8.10567
R46912 a_31699_20742.n14 a_31699_20742.t191 8.10567
R46913 a_31699_20742.n138 a_31699_20742.t116 8.10567
R46914 a_31699_20742.n291 a_31699_20742.t225 8.10567
R46915 a_31699_20742.n290 a_31699_20742.t101 8.10567
R46916 a_31699_20742.n289 a_31699_20742.t248 8.10567
R46917 a_31699_20742.n10 a_31699_20742.t169 8.10567
R46918 a_31699_20742.n11 a_31699_20742.t98 8.10567
R46919 a_31699_20742.n26 a_31699_20742.t50 8.10567
R46920 a_31699_20742.n34 a_31699_20742.t178 8.10567
R46921 a_31699_20742.n377 a_31699_20742.t9 8.10567
R46922 a_31699_20742.n382 a_31699_20742.t21 8.10567
R46923 a_31699_20742.n373 a_31699_20742.t31 8.10567
R46924 a_31699_20742.n184 a_31699_20742.t5 8.10567
R46925 a_31699_20742.n81 a_31699_20742.t19 8.10567
R46926 a_31699_20742.n366 a_31699_20742.t43 8.10567
R46927 a_31699_20742.n244 a_31699_20742.t2 6.61324
R46928 a_31699_20742.n241 a_31699_20742.t12 6.57135
R46929 a_31699_20742.n246 a_31699_20742.t26 5.34147
R46930 a_31699_20742.n245 a_31699_20742.t38 5.34147
R46931 a_31699_20742.n191 a_31699_20742.n190 1.45673
R46932 a_31699_20742.n187 a_31699_20742.n186 1.45673
R46933 a_31699_20742.n185 a_31699_20742.n184 1.45673
R46934 a_31699_20742.n148 a_31699_20742.n147 1.45418
R46935 a_31699_20742.n146 a_31699_20742.n10 1.45418
R46936 a_31699_20742.n145 a_31699_20742.n144 1.45392
R46937 a_31699_20742.n143 a_31699_20742.n142 1.45392
R46938 a_31699_20742.n242 a_31699_20742.n235 3.82989
R46939 a_31699_20742.n241 a_31699_20742.n391 3.82989
R46940 a_31699_20742.n234 a_31699_20742.n235 0.0670308
R46941 a_31699_20742.n233 a_31699_20742.t32 5.29989
R46942 a_31699_20742.n232 a_31699_20742.t6 5.29989
R46943 a_31699_20742.n174 a_31699_20742.n173 0.592804
R46944 a_31699_20742.n177 a_31699_20742.n176 0.592804
R46945 a_31699_20742.n180 a_31699_20742.n179 0.592804
R46946 a_31699_20742.n183 a_31699_20742.n182 0.592804
R46947 a_31699_20742.n199 a_31699_20742.n198 0.592738
R46948 a_31699_20742.n202 a_31699_20742.n201 0.592738
R46949 a_31699_20742.n205 a_31699_20742.n204 0.592738
R46950 a_31699_20742.n206 a_31699_20742.n207 0.592738
R46951 a_31699_20742.n159 a_31699_20742.n161 0.591918
R46952 a_31699_20742.n164 a_31699_20742.n162 0.591918
R46953 a_31699_20742.n157 a_31699_20742.n86 0.591918
R46954 a_31699_20742.n155 a_31699_20742.n153 0.591918
R46955 a_31699_20742.n152 a_31699_20742.n92 0.591918
R46956 a_31699_20742.n96 a_31699_20742.n150 0.591918
R46957 a_31699_20742.n83 a_31699_20742.n84 0.591886
R46958 a_31699_20742.n87 a_31699_20742.n88 0.591826
R46959 a_31699_20742.n90 a_31699_20742.n91 0.067621
R46960 a_31699_20742.n93 a_31699_20742.n94 0.591826
R46961 a_31699_20742.n98 a_31699_20742.n97 0.591886
R46962 a_31699_20742.n101 a_31699_20742.n100 0.0676312
R46963 a_31699_20742.n240 a_31699_20742.n239 1.46537
R46964 a_31699_20742.n110 a_31699_20742.n112 0.604258
R46965 a_31699_20742.n124 a_31699_20742.n125 0.591264
R46966 a_31699_20742.n113 a_31699_20742.n115 0.604258
R46967 a_31699_20742.n128 a_31699_20742.n127 0.591264
R46968 a_31699_20742.n132 a_31699_20742.n131 0.591264
R46969 a_31699_20742.n169 a_31699_20742.n168 0.604258
R46970 a_31699_20742.n136 a_31699_20742.n137 0.031901
R46971 a_31699_20742.n86 a_31699_20742.n156 0.591264
R46972 a_31699_20742.n89 a_31699_20742.n87 0.604195
R46973 a_31699_20742.n162 a_31699_20742.n163 0.591264
R46974 a_31699_20742.n83 a_31699_20742.n85 0.604258
R46975 a_31699_20742.n160 a_31699_20742.n159 0.591264
R46976 a_31699_20742.n216 a_31699_20742.n158 0.0732126
R46977 a_31699_20742.n105 a_31699_20742.n103 0.604258
R46978 a_31699_20742.n102 a_31699_20742.n116 0.591264
R46979 a_31699_20742.n109 a_31699_20742.n107 0.604258
R46980 a_31699_20742.n106 a_31699_20742.n118 0.591264
R46981 a_31699_20742.n121 a_31699_20742.n122 0.591264
R46982 a_31699_20742.n166 a_31699_20742.n165 0.604258
R46983 a_31699_20742.n134 a_31699_20742.n135 0.031901
R46984 a_31699_20742.n165 a_31699_20742.n167 0.604258
R46985 a_31699_20742.n117 a_31699_20742.n102 0.591264
R46986 a_31699_20742.n103 a_31699_20742.n104 0.604258
R46987 a_31699_20742.n119 a_31699_20742.n106 0.591264
R46988 a_31699_20742.n107 a_31699_20742.n108 0.604258
R46989 a_31699_20742.n123 a_31699_20742.n121 0.591264
R46990 a_31699_20742.n120 a_31699_20742.n171 0.0301596
R46991 a_31699_20742.n149 a_31699_20742.n96 0.591264
R46992 a_31699_20742.n97 a_31699_20742.n99 0.604258
R46993 a_31699_20742.n92 a_31699_20742.n151 0.591264
R46994 a_31699_20742.n95 a_31699_20742.n93 0.604195
R46995 a_31699_20742.n153 a_31699_20742.n154 0.591264
R46996 a_31699_20742.n214 a_31699_20742.n215 0.0732126
R46997 a_31699_20742.n168 a_31699_20742.n170 0.604258
R46998 a_31699_20742.n126 a_31699_20742.n124 0.591264
R46999 a_31699_20742.n111 a_31699_20742.n110 0.604258
R47000 a_31699_20742.n127 a_31699_20742.n129 0.591264
R47001 a_31699_20742.n114 a_31699_20742.n113 0.604258
R47002 a_31699_20742.n131 a_31699_20742.n133 0.591264
R47003 a_31699_20742.n130 a_31699_20742.n172 0.0301596
R47004 a_31699_20742.n141 a_31699_20742.n140 0.359454
R47005 a_31699_20742.n5 a_31699_20742.n6 1.44113
R47006 a_31699_20742.n37 a_31699_20742.n38 1.44113
R47007 a_31699_20742.n31 a_31699_20742.n30 1.44113
R47008 a_31699_20742.n21 a_31699_20742.n20 1.44113
R47009 a_31699_20742.n3 a_31699_20742.n4 1.44113
R47010 a_31699_20742.n18 a_31699_20742.n19 1.44113
R47011 a_31699_20742.n1 a_31699_20742.n2 1.44113
R47012 a_31699_20742.n0 a_31699_20742.n36 1.44113
R47013 a_31699_20742.n29 a_31699_20742.n28 1.44113
R47014 a_31699_20742.n17 a_31699_20742.n16 1.44113
R47015 a_31699_20742.n210 a_31699_20742.n211 0.332154
R47016 a_31699_20742.n79 a_31699_20742.n80 1.44113
R47017 a_31699_20742.n78 a_31699_20742.n77 1.44113
R47018 a_31699_20742.n269 a_31699_20742.n266 4.5005
R47019 a_31699_20742.n72 a_31699_20742.n71 1.44113
R47020 a_31699_20742.n73 a_31699_20742.n74 1.44113
R47021 a_31699_20742.n76 a_31699_20742.n75 1.44113
R47022 a_31699_20742.n70 a_31699_20742.n69 1.44113
R47023 a_31699_20742.n68 a_31699_20742.n67 1.44113
R47024 a_31699_20742.n66 a_31699_20742.n65 1.44113
R47025 a_31699_20742.n285 a_31699_20742.n273 4.5005
R47026 a_31699_20742.n61 a_31699_20742.n62 1.44113
R47027 a_31699_20742.n64 a_31699_20742.n63 1.44113
R47028 a_31699_20742.n189 a_31699_20742.n188 0.349872
R47029 a_31699_20742.n139 a_31699_20742.n138 0.359454
R47030 a_31699_20742.n15 a_31699_20742.n14 1.44113
R47031 a_31699_20742.n13 a_31699_20742.n40 1.44113
R47032 a_31699_20742.n35 a_31699_20742.n34 1.44113
R47033 a_31699_20742.n27 a_31699_20742.n26 1.44113
R47034 a_31699_20742.n11 a_31699_20742.n12 1.44113
R47035 a_31699_20742.n25 a_31699_20742.n24 1.44113
R47036 a_31699_20742.n8 a_31699_20742.n9 1.44113
R47037 a_31699_20742.n39 a_31699_20742.n7 1.44113
R47038 a_31699_20742.n32 a_31699_20742.n33 1.44113
R47039 a_31699_20742.n22 a_31699_20742.n23 1.44113
R47040 a_31699_20742.n212 a_31699_20742.n213 0.332154
R47041 a_31699_20742.n59 a_31699_20742.n60 1.44113
R47042 a_31699_20742.n57 a_31699_20742.n58 1.44113
R47043 a_31699_20742.n264 a_31699_20742.n263 4.5005
R47044 a_31699_20742.n52 a_31699_20742.n51 1.44113
R47045 a_31699_20742.n53 a_31699_20742.n54 1.44113
R47046 a_31699_20742.n56 a_31699_20742.n55 1.44113
R47047 a_31699_20742.n49 a_31699_20742.n50 1.44113
R47048 a_31699_20742.n48 a_31699_20742.n47 1.44113
R47049 a_31699_20742.n46 a_31699_20742.n45 1.44113
R47050 a_31699_20742.n304 a_31699_20742.n303 4.5005
R47051 a_31699_20742.n42 a_31699_20742.n41 1.44113
R47052 a_31699_20742.n44 a_31699_20742.n43 1.44113
R47053 a_31699_20742.n192 a_31699_20742.n193 0.349872
R47054 a_31699_20742.n369 a_31699_20742.n368 4.5005
R47055 a_31699_20742.n82 a_31699_20742.n81 1.44113
R47056 a_31699_20742.n385 a_31699_20742.n384 4.5005
R47057 a_31699_20742.n383 a_31699_20742.n374 4.5005
R47058 a_31699_20742.n382 a_31699_20742.n381 4.5005
R47059 a_31699_20742.n380 a_31699_20742.n375 4.5005
R47060 a_31699_20742.n379 a_31699_20742.n378 4.5005
R47061 a_31699_20742.n309 a_31699_20742.n252 3.97759
R47062 a_31699_20742.n244 a_31699_20742.n243 3.87147
R47063 a_31699_20742.n240 a_31699_20742.t4 3.86699
R47064 a_31699_20742.n240 a_31699_20742.t30 3.66212
R47065 a_31699_20742.n251 a_31699_20742.n239 3.08458
R47066 a_31699_20742.n239 a_31699_20742.n250 2.73715
R47067 a_31699_20742.n246 a_31699_20742.n245 2.51878
R47068 a_31699_20742.n251 a_31699_20742.n217 2.44398
R47069 a_31699_20742.n218 a_31699_20742.n247 3.87147
R47070 a_31699_20742.n250 a_31699_20742.n248 2.39895
R47071 a_31699_20742.n288 a_31699_20742.n265 2.30989
R47072 a_31699_20742.n280 a_31699_20742.n197 2.30989
R47073 a_31699_20742.n302 a_31699_20742.n260 2.25752
R47074 a_31699_20742.n287 a_31699_20742.n286 2.25752
R47075 a_31699_20742.n386 a_31699_20742.n373 2.25278
R47076 a_31699_20742.n218 a_31699_20742.n217 0.0670397
R47077 a_31699_20742.n220 a_31699_20742.n219 1.44642
R47078 a_31699_20742.n221 a_31699_20742.n175 1.44642
R47079 a_31699_20742.n222 a_31699_20742.n178 1.44642
R47080 a_31699_20742.n223 a_31699_20742.n181 1.44642
R47081 a_31699_20742.n227 a_31699_20742.n226 1.44612
R47082 a_31699_20742.n228 a_31699_20742.n200 1.44612
R47083 a_31699_20742.n229 a_31699_20742.n203 1.44612
R47084 a_31699_20742.n231 a_31699_20742.n230 1.44612
R47085 a_31699_20742.n250 a_31699_20742.n249 2.19216
R47086 a_31699_20742.n117 a_31699_20742.n255 2.49908
R47087 a_31699_20742.n224 a_31699_20742.n123 2.49908
R47088 a_31699_20742.n225 a_31699_20742.n126 2.49908
R47089 a_31699_20742.n133 a_31699_20742.n311 2.49908
R47090 a_31699_20742.n254 a_31699_20742.n237 2.07182
R47091 a_31699_20742.n256 a_31699_20742.n236 2.07182
R47092 a_31699_20742.n237 a_31699_20742.n157 2.4644
R47093 a_31699_20742.n161 a_31699_20742.n236 2.4644
R47094 a_31699_20742.n150 a_31699_20742.n257 2.4644
R47095 a_31699_20742.n238 a_31699_20742.n155 2.4644
R47096 a_31699_20742.n309 a_31699_20742.n308 2.01366
R47097 a_31699_20742.n334 a_31699_20742.n323 1.61908
R47098 a_31699_20742.n313 a_31699_20742.n312 1.53101
R47099 a_31699_20742.n310 a_31699_20742.n309 1.53101
R47100 a_31699_20742.n257 a_31699_20742.n253 1.5005
R47101 a_31699_20742.n255 a_31699_20742.n254 1.5005
R47102 a_31699_20742.n312 a_31699_20742.n225 1.5005
R47103 a_31699_20742.n311 a_31699_20742.n310 1.5005
R47104 a_31699_20742.n258 a_31699_20742.n238 1.5005
R47105 a_31699_20742.n256 a_31699_20742.n224 1.5005
R47106 a_31699_20742.n296 a_31699_20742.n196 1.5005
R47107 a_31699_20742.n288 a_31699_20742.n194 1.5005
R47108 a_31699_20742.n298 a_31699_20742.n297 1.5005
R47109 a_31699_20742.n308 a_31699_20742.n195 1.5005
R47110 a_31699_20742.n292 a_31699_20742.n259 1.5005
R47111 a_31699_20742.n281 a_31699_20742.n280 1.5005
R47112 a_31699_20742.n209 a_31699_20742.n365 1.5005
R47113 a_31699_20742.n208 a_31699_20742.n355 1.5005
R47114 a_31699_20742.n209 a_31699_20742.n387 1.5005
R47115 a_31699_20742.n345 a_31699_20742.n344 1.5005
R47116 a_31699_20742.n334 a_31699_20742.n333 1.5005
R47117 a_31699_20742.n234 a_31699_20742.n390 1.5005
R47118 a_31699_20742.n254 a_31699_20742.n253 1.47516
R47119 a_31699_20742.n258 a_31699_20742.n256 1.47516
R47120 a_31699_20742.n247 a_31699_20742.t16 1.4705
R47121 a_31699_20742.n247 a_31699_20742.t42 1.4705
R47122 a_31699_20742.n243 a_31699_20742.t34 1.4705
R47123 a_31699_20742.n243 a_31699_20742.t8 1.4705
R47124 a_31699_20742.n248 a_31699_20742.t24 1.4705
R47125 a_31699_20742.n248 a_31699_20742.t14 1.4705
R47126 a_31699_20742.n249 a_31699_20742.t18 1.4705
R47127 a_31699_20742.n249 a_31699_20742.t40 1.4705
R47128 a_31699_20742.n242 a_31699_20742.t22 1.4705
R47129 a_31699_20742.n242 a_31699_20742.t10 1.4705
R47130 a_31699_20742.t44 a_31699_20742.n391 1.4705
R47131 a_31699_20742.n391 a_31699_20742.t20 1.4705
R47132 a_31699_20742.n388 a_31699_20742.n209 1.42915
R47133 a_31699_20742.n297 a_31699_20742.n252 1.41182
R47134 a_31699_20742.n140 a_31699_20742.t160 8.49836
R47135 a_31699_20742.n139 a_31699_20742.t67 8.49836
R47136 a_31699_20742.n245 a_31699_20742.n244 1.27228
R47137 a_31699_20742.n28 a_31699_20742.n279 1.24866
R47138 a_31699_20742.n30 a_31699_20742.n276 1.24866
R47139 a_31699_20742.n293 a_31699_20742.n32 1.24866
R47140 a_31699_20742.n34 a_31699_20742.n291 1.24866
R47141 a_31699_20742.n277 a_31699_20742.n0 1.24629
R47142 a_31699_20742.n274 a_31699_20742.n37 1.24629
R47143 a_31699_20742.n7 a_31699_20742.n295 1.24629
R47144 a_31699_20742.n289 a_31699_20742.n13 1.24629
R47145 a_31699_20742.n296 a_31699_20742.n288 1.23709
R47146 a_31699_20742.n280 a_31699_20742.n259 1.23709
R47147 a_31699_20742.n305 a_31699_20742.n49 1.22261
R47148 a_31699_20742.n299 a_31699_20742.n59 1.22261
R47149 a_31699_20742.n69 a_31699_20742.n284 1.22261
R47150 a_31699_20742.n270 a_31699_20742.n79 1.22261
R47151 a_31699_20742.n41 a_31699_20742.n307 1.21313
R47152 a_31699_20742.n52 a_31699_20742.n301 1.21313
R47153 a_31699_20742.n282 a_31699_20742.n61 1.21313
R47154 a_31699_20742.n71 a_31699_20742.n272 1.21313
R47155 a_31699_20742.n217 a_31699_20742.n246 1.20609
R47156 a_31699_20742.n390 a_31699_20742.n389 1.17709
R47157 a_31699_20742.n269 a_31699_20742.n268 1.12904
R47158 a_31699_20742.n263 a_31699_20742.n262 1.12904
R47159 a_31699_20742.n368 a_31699_20742.n367 1.129
R47160 a_31699_20742.n379 a_31699_20742.n376 1.12765
R47161 a_31699_20742.n317 a_31699_20742.n316 0.915282
R47162 a_31699_20742.n327 a_31699_20742.n326 0.915282
R47163 a_31699_20742.n338 a_31699_20742.n337 0.915282
R47164 a_31699_20742.n349 a_31699_20742.n348 0.915282
R47165 a_31699_20742.n359 a_31699_20742.n358 0.915282
R47166 a_31699_20742.n390 a_31699_20742.n251 0.886209
R47167 a_31699_20742.n297 a_31699_20742.n296 0.809892
R47168 a_31699_20742.n308 a_31699_20742.n259 0.809892
R47169 a_31699_20742.n31 a_31699_20742.n265 0.888471
R47170 a_31699_20742.n197 a_31699_20742.n29 0.888471
R47171 a_31699_20742.n196 a_31699_20742.n35 0.888471
R47172 a_31699_20742.n33 a_31699_20742.n292 0.888471
R47173 a_31699_20742.n389 a_31699_20742.n388 0.741617
R47174 a_31699_20742.n194 a_31699_20742.n72 0.854361
R47175 a_31699_20742.n62 a_31699_20742.n281 0.854361
R47176 a_31699_20742.n298 a_31699_20742.n51 0.854361
R47177 a_31699_20742.n195 a_31699_20742.n42 0.854361
R47178 a_31699_20742.n323 a_31699_20742.n322 0.688348
R47179 a_31699_20742.n333 a_31699_20742.n332 0.688348
R47180 a_31699_20742.n344 a_31699_20742.n343 0.688348
R47181 a_31699_20742.n355 a_31699_20742.n354 0.688348
R47182 a_31699_20742.n365 a_31699_20742.n364 0.688348
R47183 a_31699_20742.n306 a_31699_20742.n305 0.673132
R47184 a_31699_20742.n307 a_31699_20742.n306 0.673132
R47185 a_31699_20742.n300 a_31699_20742.n299 0.673132
R47186 a_31699_20742.n301 a_31699_20742.n300 0.673132
R47187 a_31699_20742.n278 a_31699_20742.n277 0.673132
R47188 a_31699_20742.n279 a_31699_20742.n278 0.673132
R47189 a_31699_20742.n275 a_31699_20742.n274 0.673132
R47190 a_31699_20742.n276 a_31699_20742.n275 0.673132
R47191 a_31699_20742.n284 a_31699_20742.n283 0.673132
R47192 a_31699_20742.n283 a_31699_20742.n282 0.673132
R47193 a_31699_20742.n271 a_31699_20742.n270 0.673132
R47194 a_31699_20742.n272 a_31699_20742.n271 0.673132
R47195 a_31699_20742.n295 a_31699_20742.n294 0.673132
R47196 a_31699_20742.n294 a_31699_20742.n293 0.673132
R47197 a_31699_20742.n290 a_31699_20742.n289 0.673132
R47198 a_31699_20742.n291 a_31699_20742.n290 0.673132
R47199 a_31699_20742.n318 a_31699_20742.n317 0.655148
R47200 a_31699_20742.n328 a_31699_20742.n327 0.655148
R47201 a_31699_20742.n339 a_31699_20742.n338 0.655148
R47202 a_31699_20742.n371 a_31699_20742.n370 0.655148
R47203 a_31699_20742.n350 a_31699_20742.n349 0.655148
R47204 a_31699_20742.n360 a_31699_20742.n359 0.655148
R47205 a_31699_20742.n316 a_31699_20742.n315 0.63334
R47206 a_31699_20742.n322 a_31699_20742.n321 0.63334
R47207 a_31699_20742.n321 a_31699_20742.n320 0.63334
R47208 a_31699_20742.n326 a_31699_20742.n325 0.63334
R47209 a_31699_20742.n332 a_31699_20742.n331 0.63334
R47210 a_31699_20742.n331 a_31699_20742.n330 0.63334
R47211 a_31699_20742.n337 a_31699_20742.n336 0.63334
R47212 a_31699_20742.n343 a_31699_20742.n342 0.63334
R47213 a_31699_20742.n342 a_31699_20742.n341 0.63334
R47214 a_31699_20742.n348 a_31699_20742.n347 0.63334
R47215 a_31699_20742.n354 a_31699_20742.n353 0.63334
R47216 a_31699_20742.n353 a_31699_20742.n352 0.63334
R47217 a_31699_20742.n358 a_31699_20742.n357 0.63334
R47218 a_31699_20742.n364 a_31699_20742.n363 0.63334
R47219 a_31699_20742.n363 a_31699_20742.n362 0.63334
R47220 a_31699_20742.n315 a_31699_20742.n314 0.63225
R47221 a_31699_20742.n319 a_31699_20742.n318 0.63225
R47222 a_31699_20742.n325 a_31699_20742.n324 0.63225
R47223 a_31699_20742.n329 a_31699_20742.n328 0.63225
R47224 a_31699_20742.n336 a_31699_20742.n335 0.63225
R47225 a_31699_20742.n340 a_31699_20742.n339 0.63225
R47226 a_31699_20742.n372 a_31699_20742.n371 0.63225
R47227 a_31699_20742.n347 a_31699_20742.n346 0.63225
R47228 a_31699_20742.n351 a_31699_20742.n350 0.63225
R47229 a_31699_20742.n357 a_31699_20742.n356 0.63225
R47230 a_31699_20742.n361 a_31699_20742.n360 0.63225
R47231 a_31699_20742.n387 a_31699_20742.n386 0.622055
R47232 a_31699_20742.n313 a_31699_20742.n252 0.602344
R47233 a_31699_20742.n312 a_31699_20742.n253 0.571818
R47234 a_31699_20742.n310 a_31699_20742.n258 0.571818
R47235 a_31699_20742.n208 a_31699_20742.n345 0.467527
R47236 a_31699_20742.n63 a_31699_20742.n189 0.379447
R47237 a_31699_20742.n384 a_31699_20742.n383 0.379447
R47238 a_31699_20742.n378 a_31699_20742.n375 0.379447
R47239 a_31699_20742.n112 a_31699_20742.n125 1.14293
R47240 a_31699_20742.n115 a_31699_20742.n128 1.14293
R47241 a_31699_20742.n172 a_31699_20742.n132 1.74606
R47242 a_31699_20742.n105 a_31699_20742.n116 1.14293
R47243 a_31699_20742.n109 a_31699_20742.n118 1.14293
R47244 a_31699_20742.n171 a_31699_20742.n122 1.74606
R47245 a_31699_20742.n104 a_31699_20742.n117 1.14293
R47246 a_31699_20742.n108 a_31699_20742.n119 1.14293
R47247 a_31699_20742.n171 a_31699_20742.n123 1.74702
R47248 a_31699_20742.n111 a_31699_20742.n126 1.14293
R47249 a_31699_20742.n129 a_31699_20742.n114 1.14293
R47250 a_31699_20742.n172 a_31699_20742.n133 1.74702
R47251 a_31699_20742.n21 a_31699_20742.n4 0.647707
R47252 a_31699_20742.n2 a_31699_20742.n19 0.647707
R47253 a_31699_20742.n211 a_31699_20742.n17 1.34142
R47254 a_31699_20742.n12 a_31699_20742.n27 0.647707
R47255 a_31699_20742.n9 a_31699_20742.n25 0.647707
R47256 a_31699_20742.n213 a_31699_20742.n23 1.34142
R47257 a_31699_20742.n21 a_31699_20742.n31 0.635332
R47258 a_31699_20742.n145 a_31699_20742.n19 0.634233
R47259 a_31699_20742.n29 a_31699_20742.n17 0.635332
R47260 a_31699_20742.n35 a_31699_20742.n27 0.635332
R47261 a_31699_20742.n143 a_31699_20742.n25 0.634233
R47262 a_31699_20742.n23 a_31699_20742.n33 0.635332
R47263 a_31699_20742.n221 a_31699_20742.n177 0.891677
R47264 a_31699_20742.n174 a_31699_20742.n220 0.891677
R47265 a_31699_20742.n228 a_31699_20742.n202 0.891728
R47266 a_31699_20742.n199 a_31699_20742.n227 0.891728
R47267 a_31699_20742.n157 a_31699_20742.n88 1.1526
R47268 a_31699_20742.n84 a_31699_20742.n164 1.15248
R47269 a_31699_20742.n161 a_31699_20742.n216 1.74338
R47270 a_31699_20742.n223 a_31699_20742.n183 0.891677
R47271 a_31699_20742.n222 a_31699_20742.n180 0.891677
R47272 a_31699_20742.n207 a_31699_20742.n231 0.891728
R47273 a_31699_20742.n229 a_31699_20742.n205 0.891728
R47274 a_31699_20742.n98 a_31699_20742.n150 1.15284
R47275 a_31699_20742.n94 a_31699_20742.n152 1.1526
R47276 a_31699_20742.n155 a_31699_20742.n215 1.74338
R47277 a_31699_20742.n78 a_31699_20742.n269 0.496611
R47278 a_31699_20742.n66 a_31699_20742.n273 0.496611
R47279 a_31699_20742.n263 a_31699_20742.n58 0.496611
R47280 a_31699_20742.n303 a_31699_20742.n46 0.496611
R47281 a_31699_20742.n385 a_31699_20742.n374 0.3605
R47282 a_31699_20742.n380 a_31699_20742.n379 0.3605
R47283 a_31699_20742.n368 a_31699_20742.n82 0.495486
R47284 a_31699_20742.n262 a_31699_20742.n261 0.327481
R47285 a_31699_20742.n268 a_31699_20742.n267 0.327481
R47286 a_31699_20742.n367 a_31699_20742.n366 0.32675
R47287 a_31699_20742.n377 a_31699_20742.n376 0.324133
R47288 a_31699_20742.n345 a_31699_20742.n334 0.301209
R47289 a_31699_20742.n148 a_31699_20742.n4 0.558475
R47290 a_31699_20742.n36 a_31699_20742.n2 0.559597
R47291 a_31699_20742.n146 a_31699_20742.n12 0.558475
R47292 a_31699_20742.n39 a_31699_20742.n9 0.559597
R47293 a_31699_20742.n323 a_31699_20742.n319 0.254694
R47294 a_31699_20742.n333 a_31699_20742.n329 0.254694
R47295 a_31699_20742.n344 a_31699_20742.n340 0.254694
R47296 a_31699_20742.n387 a_31699_20742.n372 0.254694
R47297 a_31699_20742.n355 a_31699_20742.n351 0.254694
R47298 a_31699_20742.n365 a_31699_20742.n361 0.254694
R47299 a_31699_20742.n287 a_31699_20742.n273 0.208099
R47300 a_31699_20742.n303 a_31699_20742.n302 0.208099
R47301 a_31699_20742.n386 a_31699_20742.n385 0.208099
R47302 a_31699_20742.n384 a_31699_20742.n373 0.147342
R47303 a_31699_20742.n383 a_31699_20742.n382 0.147342
R47304 a_31699_20742.n382 a_31699_20742.n375 0.147342
R47305 a_31699_20742.n378 a_31699_20742.n377 0.147342
R47306 a_31699_20742.n369 a_31699_20742.n366 0.143789
R47307 a_31699_20742.n304 a_31699_20742.n260 0.142605
R47308 a_31699_20742.n264 a_31699_20742.n261 0.142605
R47309 a_31699_20742.n286 a_31699_20742.n285 0.142605
R47310 a_31699_20742.n267 a_31699_20742.n266 0.142605
R47311 a_31699_20742.n137 a_31699_20742.n169 1.73389
R47312 a_31699_20742.n221 a_31699_20742.n169 1.19478
R47313 a_31699_20742.n125 a_31699_20742.n177 1.49218
R47314 a_31699_20742.n128 a_31699_20742.n112 3.79267
R47315 a_31699_20742.n220 a_31699_20742.n115 1.19478
R47316 a_31699_20742.n174 a_31699_20742.n132 1.49218
R47317 a_31699_20742.n228 a_31699_20742.n91 1.6448
R47318 a_31699_20742.n156 a_31699_20742.n202 1.49177
R47319 a_31699_20742.n156 a_31699_20742.n89 1.14306
R47320 a_31699_20742.n89 a_31699_20742.n163 3.79279
R47321 a_31699_20742.n85 a_31699_20742.n163 1.14293
R47322 a_31699_20742.n227 a_31699_20742.n85 1.19475
R47323 a_31699_20742.n199 a_31699_20742.n160 1.49177
R47324 a_31699_20742.n216 a_31699_20742.n160 1.74677
R47325 a_31699_20742.n91 a_31699_20742.n237 1.65371
R47326 a_31699_20742.n164 a_31699_20742.n88 3.7612
R47327 a_31699_20742.n84 a_31699_20742.n236 1.21357
R47328 a_31699_20742.n166 a_31699_20742.n135 1.73389
R47329 a_31699_20742.n223 a_31699_20742.n166 1.19478
R47330 a_31699_20742.n116 a_31699_20742.n183 1.49218
R47331 a_31699_20742.n118 a_31699_20742.n105 3.79267
R47332 a_31699_20742.n222 a_31699_20742.n109 1.19478
R47333 a_31699_20742.n122 a_31699_20742.n180 1.49218
R47334 a_31699_20742.n135 a_31699_20742.n167 1.7332
R47335 a_31699_20742.n255 a_31699_20742.n167 1.21084
R47336 a_31699_20742.n104 a_31699_20742.n119 3.79267
R47337 a_31699_20742.n108 a_31699_20742.n224 1.21084
R47338 a_31699_20742.n231 a_31699_20742.n101 1.64472
R47339 a_31699_20742.n207 a_31699_20742.n149 1.49177
R47340 a_31699_20742.n99 a_31699_20742.n149 1.14329
R47341 a_31699_20742.n151 a_31699_20742.n99 3.79231
R47342 a_31699_20742.n95 a_31699_20742.n151 1.14306
R47343 a_31699_20742.n229 a_31699_20742.n95 1.19488
R47344 a_31699_20742.n154 a_31699_20742.n205 1.49177
R47345 a_31699_20742.n154 a_31699_20742.n215 1.74677
R47346 a_31699_20742.n257 a_31699_20742.n101 1.65364
R47347 a_31699_20742.n152 a_31699_20742.n98 3.76072
R47348 a_31699_20742.n94 a_31699_20742.n238 1.21369
R47349 a_31699_20742.n170 a_31699_20742.n137 1.7332
R47350 a_31699_20742.n170 a_31699_20742.n225 1.21084
R47351 a_31699_20742.n111 a_31699_20742.n129 3.79267
R47352 a_31699_20742.n114 a_31699_20742.n311 1.21084
R47353 a_31699_20742.n140 a_31699_20742.n6 1.34213
R47354 a_31699_20742.n38 a_31699_20742.n6 0.559597
R47355 a_31699_20742.n265 a_31699_20742.n38 2.32622
R47356 a_31699_20742.n145 a_31699_20742.n148 3.29987
R47357 a_31699_20742.n36 a_31699_20742.n197 2.32622
R47358 a_31699_20742.n80 a_31699_20742.n78 0.633082
R47359 a_31699_20742.n80 a_31699_20742.n194 2.30372
R47360 a_31699_20742.n74 a_31699_20742.n72 0.633082
R47361 a_31699_20742.n74 a_31699_20742.n76 0.633082
R47362 a_31699_20742.n76 a_31699_20742.n187 0.631741
R47363 a_31699_20742.n187 a_31699_20742.n287 3.17649
R47364 a_31699_20742.n66 a_31699_20742.n68 0.633082
R47365 a_31699_20742.n68 a_31699_20742.n70 0.633082
R47366 a_31699_20742.n70 a_31699_20742.n281 2.30372
R47367 a_31699_20742.n62 a_31699_20742.n64 0.633082
R47368 a_31699_20742.n64 a_31699_20742.n188 1.32892
R47369 a_31699_20742.n15 a_31699_20742.n139 1.34213
R47370 a_31699_20742.n40 a_31699_20742.n15 0.559597
R47371 a_31699_20742.n40 a_31699_20742.n196 2.32622
R47372 a_31699_20742.n146 a_31699_20742.n143 3.29987
R47373 a_31699_20742.n39 a_31699_20742.n292 2.32622
R47374 a_31699_20742.n60 a_31699_20742.n58 0.633082
R47375 a_31699_20742.n298 a_31699_20742.n60 2.30372
R47376 a_31699_20742.n54 a_31699_20742.n51 0.633082
R47377 a_31699_20742.n56 a_31699_20742.n54 0.633082
R47378 a_31699_20742.n191 a_31699_20742.n56 0.631741
R47379 a_31699_20742.n302 a_31699_20742.n191 3.17649
R47380 a_31699_20742.n48 a_31699_20742.n46 0.633082
R47381 a_31699_20742.n50 a_31699_20742.n48 0.633082
R47382 a_31699_20742.n50 a_31699_20742.n195 2.30372
R47383 a_31699_20742.n44 a_31699_20742.n42 0.633082
R47384 a_31699_20742.n44 a_31699_20742.n193 1.32892
R47385 a_31699_20742.n185 a_31699_20742.n82 0.631741
R47386 a_31699_20742.n370 a_31699_20742.n185 0.917116
R47387 a_31699_20742.n381 a_31699_20742.n374 0.14
R47388 a_31699_20742.n381 a_31699_20742.n380 0.14
R47389 a_31699_20742.n241 a_31699_20742.n232 1.27192
R47390 a_31699_20742.n233 a_31699_20742.n232 2.51878
R47391 a_31699_20742.n234 a_31699_20742.n233 1.2061
R47392 a_31699_20742.t36 a_31699_20742.n235 6.57099
R47393 a_31699_20742.n218 a_31699_20742.t28 6.61288
R47394 a_31699_20742.n71 a_31699_20742.n73 0.966816
R47395 a_31699_20742.n61 a_31699_20742.n63 0.966816
R47396 a_31699_20742.n53 a_31699_20742.n52 0.966816
R47397 a_31699_20742.n8 a_31699_20742.n7 0.889842
R47398 a_31699_20742.n1 a_31699_20742.n0 0.889842
R47399 a_31699_20742.n11 a_31699_20742.n10 0.771421
R47400 a_31699_20742.n147 a_31699_20742.n3 0.771421
R47401 a_31699_20742.n26 a_31699_20742.n11 0.688526
R47402 a_31699_20742.n24 a_31699_20742.n8 0.688526
R47403 a_31699_20742.n22 a_31699_20742.n212 0.688526
R47404 a_31699_20742.n3 a_31699_20742.n20 0.688526
R47405 a_31699_20742.n1 a_31699_20742.n18 0.688526
R47406 a_31699_20742.n16 a_31699_20742.n210 0.688526
R47407 a_31699_20742.n14 a_31699_20742.n138 0.688526
R47408 a_31699_20742.n5 a_31699_20742.n141 0.688526
R47409 a_31699_20742.n34 a_31699_20742.n26 0.6755
R47410 a_31699_20742.n32 a_31699_20742.n22 0.6755
R47411 a_31699_20742.n20 a_31699_20742.n30 0.6755
R47412 a_31699_20742.n28 a_31699_20742.n16 0.6755
R47413 a_31699_20742.n77 a_31699_20742.n79 0.673132
R47414 a_31699_20742.n77 a_31699_20742.n266 0.673132
R47415 a_31699_20742.n73 a_31699_20742.n75 0.673132
R47416 a_31699_20742.n67 a_31699_20742.n69 0.673132
R47417 a_31699_20742.n65 a_31699_20742.n67 0.673132
R47418 a_31699_20742.n285 a_31699_20742.n65 0.673132
R47419 a_31699_20742.n59 a_31699_20742.n57 0.673132
R47420 a_31699_20742.n57 a_31699_20742.n264 0.673132
R47421 a_31699_20742.n55 a_31699_20742.n53 0.673132
R47422 a_31699_20742.n47 a_31699_20742.n49 0.673132
R47423 a_31699_20742.n47 a_31699_20742.n45 0.673132
R47424 a_31699_20742.n45 a_31699_20742.n304 0.673132
R47425 a_31699_20742.n43 a_31699_20742.n192 0.673132
R47426 a_31699_20742.n41 a_31699_20742.n43 0.673132
R47427 a_31699_20742.n81 a_31699_20742.n369 0.671947
R47428 a_31699_20742.n127 a_31699_20742.n113 0.609682
R47429 a_31699_20742.n124 a_31699_20742.n110 0.609682
R47430 a_31699_20742.n107 a_31699_20742.n106 0.609682
R47431 a_31699_20742.n103 a_31699_20742.n102 0.609682
R47432 a_31699_20742.n97 a_31699_20742.n96 0.609682
R47433 a_31699_20742.n93 a_31699_20742.n92 0.609682
R47434 a_31699_20742.n87 a_31699_20742.n86 0.609682
R47435 a_31699_20742.n162 a_31699_20742.n83 0.609682
R47436 a_31699_20742.n14 a_31699_20742.n13 0.596158
R47437 a_31699_20742.n37 a_31699_20742.n5 0.596158
R47438 a_31699_20742.n18 a_31699_20742.n144 0.559447
R47439 a_31699_20742.n142 a_31699_20742.n24 0.559447
R47440 a_31699_20742.n190 a_31699_20742.n55 0.531026
R47441 a_31699_20742.n75 a_31699_20742.n186 0.531026
R47442 a_31699_20742.n184 a_31699_20742.n81 0.531026
R47443 a_31699_20742.n209 a_31699_20742.n208 0.427696
R47444 a_31699_20742.n182 a_31699_20742.n181 0.386311
R47445 a_31699_20742.n179 a_31699_20742.n178 0.386311
R47446 a_31699_20742.n176 a_31699_20742.n175 0.386311
R47447 a_31699_20742.n219 a_31699_20742.n173 0.386311
R47448 a_31699_20742.n131 a_31699_20742.n130 0.369148
R47449 a_31699_20742.n121 a_31699_20742.n120 0.369148
R47450 a_31699_20742.n230 a_31699_20742.n206 0.364343
R47451 a_31699_20742.n204 a_31699_20742.n203 0.364343
R47452 a_31699_20742.n201 a_31699_20742.n200 0.364343
R47453 a_31699_20742.n226 a_31699_20742.n198 0.364343
R47454 a_31699_20742.n159 a_31699_20742.n158 0.354735
R47455 a_31699_20742.n214 a_31699_20742.n153 0.354735
R47456 a_31699_20742.n168 a_31699_20742.n136 0.347689
R47457 a_31699_20742.n165 a_31699_20742.n134 0.347689
R47458 a_35502_24538.n131 a_35502_24538.n130 12.734
R47459 a_35502_24538.n57 a_35502_24538.t36 8.41809
R47460 a_35502_24538.n58 a_35502_24538.t59 8.41809
R47461 a_35502_24538.n57 a_35502_24538.t34 8.37125
R47462 a_35502_24538.n61 a_35502_24538.t41 8.37125
R47463 a_35502_24538.n58 a_35502_24538.t56 8.37125
R47464 a_35502_24538.n104 a_35502_24538.t25 8.33806
R47465 a_35502_24538.n98 a_35502_24538.t61 8.3366
R47466 a_35502_24538.n83 a_35502_24538.t47 8.26493
R47467 a_35502_24538.n117 a_35502_24538.t39 8.2602
R47468 a_35502_24538.n17 a_35502_24538.t42 8.06917
R47469 a_35502_24538.n28 a_35502_24538.t38 8.06917
R47470 a_35502_24538.n13 a_35502_24538.t50 8.06917
R47471 a_35502_24538.n13 a_35502_24538.t48 8.06917
R47472 a_35502_24538.n11 a_35502_24538.t40 8.06917
R47473 a_35502_24538.n11 a_35502_24538.t55 8.06917
R47474 a_35502_24538.n63 a_35502_24538.t26 8.06917
R47475 a_35502_24538.n17 a_35502_24538.t53 8.06917
R47476 a_35502_24538.n30 a_35502_24538.t24 8.06917
R47477 a_35502_24538.n7 a_35502_24538.t64 8.06917
R47478 a_35502_24538.n7 a_35502_24538.t37 8.06917
R47479 a_35502_24538.n32 a_35502_24538.t49 8.06917
R47480 a_35502_24538.n77 a_35502_24538.t62 8.06917
R47481 a_35502_24538.n3 a_35502_24538.t33 8.06917
R47482 a_35502_24538.n3 a_35502_24538.t31 8.06917
R47483 a_35502_24538.n21 a_35502_24538.t60 8.06917
R47484 a_35502_24538.n21 a_35502_24538.t32 8.06917
R47485 a_35502_24538.n71 a_35502_24538.t46 8.06917
R47486 a_35502_24538.n97 a_35502_24538.t29 8.06917
R47487 a_35502_24538.n0 a_35502_24538.t28 8.06917
R47488 a_35502_24538.n95 a_35502_24538.t57 8.06917
R47489 a_35502_24538.n94 a_35502_24538.t30 8.06917
R47490 a_35502_24538.n93 a_35502_24538.t45 8.06917
R47491 a_35502_24538.n91 a_35502_24538.t63 8.06917
R47492 a_35502_24538.n84 a_35502_24538.t35 8.06917
R47493 a_35502_24538.n111 a_35502_24538.t43 8.06917
R47494 a_35502_24538.n105 a_35502_24538.t54 8.06917
R47495 a_35502_24538.n113 a_35502_24538.t27 8.06917
R47496 a_35502_24538.n114 a_35502_24538.t58 8.06917
R47497 a_35502_24538.n115 a_35502_24538.t44 8.06917
R47498 a_35502_24538.n118 a_35502_24538.t52 8.06917
R47499 a_35502_24538.n124 a_35502_24538.t51 8.06917
R47500 a_35502_24538.n60 a_35502_24538.t0 6.65728
R47501 a_35502_24538.n46 a_35502_24538.t7 6.51495
R47502 a_35502_24538.n134 a_35502_24538.t15 6.40828
R47503 a_35502_24538.n43 a_35502_24538.t17 6.37877
R47504 a_35502_24538.n60 a_35502_24538.t1 5.74368
R47505 a_35502_24538.n47 a_35502_24538.t6 5.24318
R47506 a_35502_24538.n65 a_35502_24538.n31 2.4223
R47507 a_35502_24538.n72 a_35502_24538.n33 2.42484
R47508 a_35502_24538.n73 a_35502_24538.n33 2.4256
R47509 a_35502_24538.n39 a_35502_24538.n38 2.24636
R47510 a_35502_24538.t11 a_35502_24538.n35 5.26436
R47511 a_35502_24538.n54 a_35502_24538.n43 4.60825
R47512 a_35502_24538.n34 a_35502_24538.n138 3.79435
R47513 a_35502_24538.n38 a_35502_24538.n134 4.59811
R47514 a_35502_24538.n22 a_35502_24538.n21 0.592766
R47515 a_35502_24538.n12 a_35502_24538.n11 0.592803
R47516 a_35502_24538.n15 a_35502_24538.n13 0.591918
R47517 a_35502_24538.n17 a_35502_24538.n18 0.591826
R47518 a_35502_24538.n37 a_35502_24538.n36 2.24389
R47519 a_35502_24538.n50 a_35502_24538.n44 4.5005
R47520 a_35502_24538.n10 a_35502_24538.n67 4.5005
R47521 a_35502_24538.n13 a_35502_24538.n14 0.591264
R47522 a_35502_24538.n68 a_35502_24538.n24 4.5005
R47523 a_35502_24538.n31 a_35502_24538.n30 0.0133501
R47524 a_35502_24538.n16 a_35502_24538.n65 4.5005
R47525 a_35502_24538.n19 a_35502_24538.n17 0.604195
R47526 a_35502_24538.n29 a_35502_24538.n64 4.5005
R47527 a_35502_24538.n70 a_35502_24538.n69 4.5005
R47528 a_35502_24538.n28 a_35502_24538.n27 0.0143905
R47529 a_35502_24538.n20 a_35502_24538.n75 4.5005
R47530 a_35502_24538.n2 a_35502_24538.n76 4.5005
R47531 a_35502_24538.n3 a_35502_24538.n4 0.591675
R47532 a_35502_24538.n9 a_35502_24538.n7 0.604671
R47533 a_35502_24538.n6 a_35502_24538.n72 4.5005
R47534 a_35502_24538.n32 a_35502_24538.n33 0.0107891
R47535 a_35502_24538.n7 a_35502_24538.n8 0.604671
R47536 a_35502_24538.n73 a_35502_24538.n6 4.5005
R47537 a_35502_24538.n2 a_35502_24538.n23 4.5005
R47538 a_35502_24538.n5 a_35502_24538.n3 0.591675
R47539 a_35502_24538.n85 a_35502_24538.n82 4.5005
R47540 a_35502_24538.n87 a_35502_24538.n86 4.5005
R47541 a_35502_24538.n88 a_35502_24538.n81 4.5005
R47542 a_35502_24538.n90 a_35502_24538.n89 4.5005
R47543 a_35502_24538.n92 a_35502_24538.n80 4.5005
R47544 a_35502_24538.n1 a_35502_24538.n0 1.44113
R47545 a_35502_24538.n99 a_35502_24538.n96 4.5005
R47546 a_35502_24538.n112 a_35502_24538.n101 4.5005
R47547 a_35502_24538.n110 a_35502_24538.n109 4.5005
R47548 a_35502_24538.n108 a_35502_24538.n103 4.5005
R47549 a_35502_24538.n107 a_35502_24538.n106 4.5005
R47550 a_35502_24538.n127 a_35502_24538.n126 4.5005
R47551 a_35502_24538.n125 a_35502_24538.n102 4.5005
R47552 a_35502_24538.n123 a_35502_24538.n122 4.5005
R47553 a_35502_24538.n121 a_35502_24538.n116 4.5005
R47554 a_35502_24538.n120 a_35502_24538.n119 4.5005
R47555 a_35502_24538.n42 a_35502_24538.n41 2.23676
R47556 a_35502_24538.n139 a_35502_24538.n40 4.5005
R47557 a_35502_24538.n36 a_35502_24538.t9 3.79594
R47558 a_35502_24538.n41 a_35502_24538.t3 3.79475
R47559 a_35502_24538.t23 a_35502_24538.n141 3.77936
R47560 a_35502_24538.n51 a_35502_24538.t12 3.77818
R47561 a_35502_24538.n46 a_35502_24538.n45 3.77318
R47562 a_35502_24538.n137 a_35502_24538.n136 3.77081
R47563 a_35502_24538.n49 a_35502_24538.n48 3.75571
R47564 a_35502_24538.n132 a_35502_24538.n56 2.69513
R47565 a_35502_24538.n78 a_35502_24538.n76 2.4256
R47566 a_35502_24538.n23 a_35502_24538.n78 2.42484
R47567 a_35502_24538.n31 a_35502_24538.n64 2.43326
R47568 a_35502_24538.n38 a_35502_24538.n135 2.32949
R47569 a_35502_24538.n129 a_35502_24538.n100 2.30989
R47570 a_35502_24538.n54 a_35502_24538.n53 2.30818
R47571 a_35502_24538.n141 a_35502_24538.n140 2.24481
R47572 a_35502_24538.n55 a_35502_24538.n54 2.2442
R47573 a_35502_24538.n52 a_35502_24538.n51 2.24358
R47574 a_35502_24538.n74 a_35502_24538.n71 2.23529
R47575 a_35502_24538.n66 a_35502_24538.n63 2.23423
R47576 a_35502_24538.n100 a_35502_24538.n80 2.18975
R47577 a_35502_24538.n128 a_35502_24538.n101 2.16725
R47578 a_35502_24538.n26 a_35502_24538.n5 2.4981
R47579 a_35502_24538.n130 a_35502_24538.n79 2.07557
R47580 a_35502_24538.n79 a_35502_24538.n25 2.07182
R47581 a_35502_24538.n25 a_35502_24538.n15 2.4644
R47582 a_35502_24538.n61 a_35502_24538.n60 1.7613
R47583 a_35502_24538.n59 a_35502_24538.n57 1.55888
R47584 a_35502_24538.n79 a_35502_24538.n26 1.5005
R47585 a_35502_24538.n129 a_35502_24538.n128 1.5005
R47586 a_35502_24538.n59 a_35502_24538.n58 1.5005
R47587 a_35502_24538.n62 a_35502_24538.n61 1.5005
R47588 a_35502_24538.n133 a_35502_24538.n132 1.5005
R47589 a_35502_24538.n138 a_35502_24538.t21 1.4705
R47590 a_35502_24538.n138 a_35502_24538.t13 1.4705
R47591 a_35502_24538.n48 a_35502_24538.t2 1.4705
R47592 a_35502_24538.n48 a_35502_24538.t20 1.4705
R47593 a_35502_24538.n45 a_35502_24538.t22 1.4705
R47594 a_35502_24538.n45 a_35502_24538.t16 1.4705
R47595 a_35502_24538.n53 a_35502_24538.t10 1.4705
R47596 a_35502_24538.n53 a_35502_24538.t19 1.4705
R47597 a_35502_24538.n135 a_35502_24538.t8 1.4705
R47598 a_35502_24538.n135 a_35502_24538.t18 1.4705
R47599 a_35502_24538.n136 a_35502_24538.t14 1.4705
R47600 a_35502_24538.n136 a_35502_24538.t5 1.4705
R47601 a_35502_24538.n83 a_35502_24538.n82 1.39514
R47602 a_35502_24538.n120 a_35502_24538.n117 1.39105
R47603 a_35502_24538.n130 a_35502_24538.n129 1.35453
R47604 a_35502_24538.n47 a_35502_24538.n46 1.27228
R47605 a_35502_24538.n93 a_35502_24538.n92 1.26997
R47606 a_35502_24538.n0 a_35502_24538.n95 1.24392
R47607 a_35502_24538.n113 a_35502_24538.n112 1.24204
R47608 a_35502_24538.n140 a_35502_24538.n137 1.20603
R47609 a_35502_24538.n126 a_35502_24538.n115 1.20414
R47610 a_35502_24538.n99 a_35502_24538.n98 1.14132
R47611 a_35502_24538.n55 a_35502_24538.n52 1.13952
R47612 a_35502_24538.n107 a_35502_24538.n104 1.13598
R47613 a_35502_24538.n37 a_35502_24538.n49 1.20574
R47614 a_35502_24538.n42 a_35502_24538.n34 1.24017
R47615 a_35502_24538.n132 a_35502_24538.n131 0.963743
R47616 a_35502_24538.n49 a_35502_24538.n47 0.937067
R47617 a_35502_24538.n100 a_35502_24538.n1 0.888471
R47618 a_35502_24538.n128 a_35502_24538.n127 0.71825
R47619 a_35502_24538.n94 a_35502_24538.n93 0.663658
R47620 a_35502_24538.n95 a_35502_24538.n94 0.663658
R47621 a_35502_24538.n115 a_35502_24538.n114 0.655156
R47622 a_35502_24538.n114 a_35502_24538.n113 0.655156
R47623 a_35502_24538.n118 a_35502_24538.n117 0.439529
R47624 a_35502_24538.n84 a_35502_24538.n83 0.432797
R47625 a_35502_24538.n123 a_35502_24538.n116 0.379447
R47626 a_35502_24538.n106 a_35502_24538.n103 0.379447
R47627 a_35502_24538.n65 a_35502_24538.n19 0.745981
R47628 a_35502_24538.n9 a_35502_24538.n72 0.745252
R47629 a_35502_24538.n8 a_35502_24538.n73 0.745252
R47630 a_35502_24538.n1 a_35502_24538.n99 0.498861
R47631 a_35502_24538.n67 a_35502_24538.n12 0.756573
R47632 a_35502_24538.n18 a_35502_24538.n64 0.756388
R47633 a_35502_24538.n15 a_35502_24538.n70 0.756711
R47634 a_35502_24538.n75 a_35502_24538.n22 0.756011
R47635 a_35502_24538.n108 a_35502_24538.n107 0.3605
R47636 a_35502_24538.n122 a_35502_24538.n121 0.3605
R47637 a_35502_24538.n98 a_35502_24538.n97 0.335806
R47638 a_35502_24538.n105 a_35502_24538.n104 0.33475
R47639 a_35502_24538.n86 a_35502_24538.n81 0.302474
R47640 a_35502_24538.n88 a_35502_24538.n87 0.287375
R47641 a_35502_24538.n131 a_35502_24538.n62 0.277797
R47642 a_35502_24538.n67 a_35502_24538.n66 0.208888
R47643 a_35502_24538.n75 a_35502_24538.n74 0.20887
R47644 a_35502_24538.n52 a_35502_24538.n44 0.208394
R47645 a_35502_24538.n140 a_35502_24538.n139 0.208357
R47646 a_35502_24538.n62 a_35502_24538.n59 0.168946
R47647 a_35502_24538.n37 a_35502_24538.n44 0.233116
R47648 a_35502_24538.n86 a_35502_24538.n85 0.147342
R47649 a_35502_24538.n90 a_35502_24538.n81 0.147342
R47650 a_35502_24538.n126 a_35502_24538.n125 0.147342
R47651 a_35502_24538.n119 a_35502_24538.n116 0.147342
R47652 a_35502_24538.n110 a_35502_24538.n103 0.147342
R47653 a_35502_24538.n139 a_35502_24538.n42 0.211956
R47654 a_35502_24538.n41 a_35502_24538.n40 0.142388
R47655 a_35502_24538.n56 a_35502_24538.n43 0.14
R47656 a_35502_24538.n66 a_35502_24538.n19 1.12746
R47657 a_35502_24538.n14 a_35502_24538.n12 1.49123
R47658 a_35502_24538.n14 a_35502_24538.n24 0.772202
R47659 a_35502_24538.n18 a_35502_24538.n25 1.21369
R47660 a_35502_24538.n70 a_35502_24538.n27 2.42126
R47661 a_35502_24538.n74 a_35502_24538.n9 1.12837
R47662 a_35502_24538.n4 a_35502_24538.n22 1.49118
R47663 a_35502_24538.n76 a_35502_24538.n4 0.772883
R47664 a_35502_24538.n8 a_35502_24538.n26 1.21186
R47665 a_35502_24538.n5 a_35502_24538.n23 0.772883
R47666 a_35502_24538.n87 a_35502_24538.n82 0.14
R47667 a_35502_24538.n89 a_35502_24538.n88 0.14
R47668 a_35502_24538.n89 a_35502_24538.n80 0.14
R47669 a_35502_24538.n109 a_35502_24538.n108 0.14
R47670 a_35502_24538.n109 a_35502_24538.n101 0.14
R47671 a_35502_24538.n127 a_35502_24538.n102 0.14
R47672 a_35502_24538.n122 a_35502_24538.n102 0.14
R47673 a_35502_24538.n121 a_35502_24538.n120 0.14
R47674 a_35502_24538.n35 a_35502_24538.n39 1.19679
R47675 a_35502_24538.n137 a_35502_24538.n35 0.932624
R47676 a_35502_24538.t4 a_35502_24538.n34 6.53226
R47677 a_35502_24538.n112 a_35502_24538.n111 0.137868
R47678 a_35502_24538.n50 a_35502_24538.n36 0.137318
R47679 a_35502_24538.n134 a_35502_24538.n133 0.131
R47680 a_35502_24538.n97 a_35502_24538.n96 0.128395
R47681 a_35502_24538.n106 a_35502_24538.n105 0.128395
R47682 a_35502_24538.n124 a_35502_24538.n123 0.118921
R47683 a_35502_24538.n92 a_35502_24538.n91 0.114184
R47684 a_35502_24538.n51 a_35502_24538.n50 0.110782
R47685 a_35502_24538.n141 a_35502_24538.n40 0.105711
R47686 a_35502_24538.n56 a_35502_24538.n55 0.0688756
R47687 a_35502_24538.n32 a_35502_24538.n6 0.0402153
R47688 a_35502_24538.n85 a_35502_24538.n84 0.0348421
R47689 a_35502_24538.n20 a_35502_24538.n71 0.0344623
R47690 a_35502_24538.n91 a_35502_24538.n90 0.0336579
R47691 a_35502_24538.n10 a_35502_24538.n63 0.0325285
R47692 a_35502_24538.n30 a_35502_24538.n29 0.0299662
R47693 a_35502_24538.n125 a_35502_24538.n124 0.0289211
R47694 a_35502_24538.n2 a_35502_24538.n77 0.0283648
R47695 a_35502_24538.n68 a_35502_24538.n28 0.0258025
R47696 a_35502_24538.n78 a_35502_24538.n77 0.0226397
R47697 a_35502_24538.n119 a_35502_24538.n118 0.0194474
R47698 a_35502_24538.n69 a_35502_24538.n68 0.0149128
R47699 a_35502_24538.n16 a_35502_24538.n29 0.0107491
R47700 a_35502_24538.n111 a_35502_24538.n110 0.00997368
R47701 a_35502_24538.n133 a_35502_24538.n39 0.0777922
R47702 a_35502_24538.n24 a_35502_24538.n27 2.43637
R47703 a_35502_24538.n0 a_35502_24538.n96 0.6755
R47704 a_35502_24538.n3 a_35502_24538.n2 0.369148
R47705 a_35502_24538.n69 a_35502_24538.n13 0.354735
R47706 a_35502_24538.n7 a_35502_24538.n6 0.347689
R47707 a_35502_24538.n17 a_35502_24538.n16 0.347689
R47708 a_35502_24538.n21 a_35502_24538.n20 0.346915
R47709 a_35502_24538.n11 a_35502_24538.n10 0.32719
R47710 a_41891_4481.n1 a_41891_4481.t7 10.2515
R47711 a_41891_4481.n1 a_41891_4481.t9 10.2515
R47712 a_41891_4481.n1 a_41891_4481.t22 10.2515
R47713 a_41891_4481.n1 a_41891_4481.t16 10.2515
R47714 a_41891_4481.n1 a_41891_4481.t3 10.096
R47715 a_41891_4481.n1 a_41891_4481.t21 10.0935
R47716 a_41891_4481.n1 a_41891_4481.t5 10.0859
R47717 a_41891_4481.n1 a_41891_4481.t15 10.0808
R47718 a_41891_4481.n1 a_41891_4481.t18 9.53981
R47719 a_41891_4481.n1 a_41891_4481.t14 9.53981
R47720 a_41891_4481.n1 a_41891_4481.t20 9.53981
R47721 a_41891_4481.n1 a_41891_4481.t12 9.53981
R47722 a_41891_4481.n1 a_41891_4481.t17 9.53744
R47723 a_41891_4481.n1 a_41891_4481.t13 9.53744
R47724 a_41891_4481.n1 a_41891_4481.t19 9.53744
R47725 a_41891_4481.n1 a_41891_4481.t11 9.53744
R47726 a_41891_4481.n1 a_41891_4481.n0 8.41434
R47727 a_41891_4481.n1 a_41891_4481.t8 8.14082
R47728 a_41891_4481.n0 a_41891_4481.t10 8.13828
R47729 a_41891_4481.t0 a_41891_4481.t1 7.96115
R47730 a_41891_4481.t0 a_41891_4481.t2 7.94694
R47731 a_41891_4481.t0 a_41891_4481.n1 7.50666
R47732 a_41891_4481.n0 a_41891_4481.t4 7.48586
R47733 a_41891_4481.n1 a_41891_4481.t6 7.48333
R47734 a_71281_n8397.n1 a_71281_n8397.n585 13.5116
R47735 a_71281_n8397.n585 a_71281_n8397.t73 10.674
R47736 a_71281_n8397.n710 a_71281_n8397.t89 10.5154
R47737 a_71281_n8397.t89 a_71281_n8397.n705 10.5154
R47738 a_71281_n8397.n724 a_71281_n8397.t163 10.5154
R47739 a_71281_n8397.t163 a_71281_n8397.n719 10.5154
R47740 a_71281_n8397.t83 a_71281_n8397.n802 10.5154
R47741 a_71281_n8397.n806 a_71281_n8397.t83 10.5154
R47742 a_71281_n8397.t156 a_71281_n8397.n789 10.5154
R47743 a_71281_n8397.n793 a_71281_n8397.t156 10.5154
R47744 a_71281_n8397.t120 a_71281_n8397.n588 10.5154
R47745 a_71281_n8397.n592 a_71281_n8397.t120 10.5154
R47746 a_71281_n8397.t195 a_71281_n8397.n601 10.5154
R47747 a_71281_n8397.n605 a_71281_n8397.t195 10.5154
R47748 a_71281_n8397.t182 a_71281_n8397.n615 10.5154
R47749 a_71281_n8397.n619 a_71281_n8397.t182 10.5154
R47750 a_71281_n8397.t251 a_71281_n8397.n629 10.5154
R47751 a_71281_n8397.n633 a_71281_n8397.t251 10.5154
R47752 a_71281_n8397.t241 a_71281_n8397.n646 10.5154
R47753 a_71281_n8397.n650 a_71281_n8397.t241 10.5154
R47754 a_71281_n8397.t308 a_71281_n8397.n660 10.5154
R47755 a_71281_n8397.n664 a_71281_n8397.t308 10.5154
R47756 a_71281_n8397.t287 a_71281_n8397.n677 10.5154
R47757 a_71281_n8397.n681 a_71281_n8397.t287 10.5154
R47758 a_71281_n8397.t100 a_71281_n8397.n691 10.5154
R47759 a_71281_n8397.n695 a_71281_n8397.t100 10.5154
R47760 a_71281_n8397.n126 a_71281_n8397.t318 10.5154
R47761 a_71281_n8397.t318 a_71281_n8397.n121 10.5154
R47762 a_71281_n8397.n140 a_71281_n8397.t131 10.5154
R47763 a_71281_n8397.t131 a_71281_n8397.n135 10.5154
R47764 a_71281_n8397.t200 a_71281_n8397.n162 10.5154
R47765 a_71281_n8397.n166 a_71281_n8397.t200 10.5154
R47766 a_71281_n8397.t264 a_71281_n8397.n149 10.5154
R47767 a_71281_n8397.n153 a_71281_n8397.t264 10.5154
R47768 a_71281_n8397.t81 a_71281_n8397.n4 10.5154
R47769 a_71281_n8397.n8 a_71281_n8397.t81 10.5154
R47770 a_71281_n8397.t154 a_71281_n8397.n17 10.5154
R47771 a_71281_n8397.n21 a_71281_n8397.t154 10.5154
R47772 a_71281_n8397.t151 a_71281_n8397.n31 10.5154
R47773 a_71281_n8397.n35 a_71281_n8397.t151 10.5154
R47774 a_71281_n8397.t222 a_71281_n8397.n45 10.5154
R47775 a_71281_n8397.n49 a_71281_n8397.t222 10.5154
R47776 a_71281_n8397.t214 a_71281_n8397.n62 10.5154
R47777 a_71281_n8397.n66 a_71281_n8397.t214 10.5154
R47778 a_71281_n8397.t281 a_71281_n8397.n76 10.5154
R47779 a_71281_n8397.n80 a_71281_n8397.t281 10.5154
R47780 a_71281_n8397.t261 a_71281_n8397.n93 10.5154
R47781 a_71281_n8397.n97 a_71281_n8397.t261 10.5154
R47782 a_71281_n8397.t326 a_71281_n8397.n107 10.5154
R47783 a_71281_n8397.n111 a_71281_n8397.t326 10.5154
R47784 a_71281_n8397.n285 a_71281_n8397.t143 10.5154
R47785 a_71281_n8397.t143 a_71281_n8397.n280 10.5154
R47786 a_71281_n8397.n271 a_71281_n8397.t215 10.5154
R47787 a_71281_n8397.t215 a_71281_n8397.n266 10.5154
R47788 a_71281_n8397.n257 a_71281_n8397.t198 10.5154
R47789 a_71281_n8397.t198 a_71281_n8397.n252 10.5154
R47790 a_71281_n8397.n243 a_71281_n8397.t204 10.5154
R47791 a_71281_n8397.t204 a_71281_n8397.n238 10.5154
R47792 a_71281_n8397.n226 a_71281_n8397.t197 10.5154
R47793 a_71281_n8397.t197 a_71281_n8397.n221 10.5154
R47794 a_71281_n8397.n212 a_71281_n8397.t262 10.5154
R47795 a_71281_n8397.t262 a_71281_n8397.n207 10.5154
R47796 a_71281_n8397.n195 a_71281_n8397.t253 10.5154
R47797 a_71281_n8397.t253 a_71281_n8397.n190 10.5154
R47798 a_71281_n8397.n181 a_71281_n8397.t319 10.5154
R47799 a_71281_n8397.t319 a_71281_n8397.n176 10.5154
R47800 a_71281_n8397.n417 a_71281_n8397.t97 10.5154
R47801 a_71281_n8397.t97 a_71281_n8397.n412 10.5154
R47802 a_71281_n8397.n431 a_71281_n8397.t170 10.5154
R47803 a_71281_n8397.t170 a_71281_n8397.n426 10.5154
R47804 a_71281_n8397.t101 a_71281_n8397.n453 10.5154
R47805 a_71281_n8397.n457 a_71281_n8397.t101 10.5154
R47806 a_71281_n8397.t173 a_71281_n8397.n440 10.5154
R47807 a_71281_n8397.n444 a_71281_n8397.t173 10.5154
R47808 a_71281_n8397.t126 a_71281_n8397.n295 10.5154
R47809 a_71281_n8397.n299 a_71281_n8397.t126 10.5154
R47810 a_71281_n8397.t201 a_71281_n8397.n308 10.5154
R47811 a_71281_n8397.n312 a_71281_n8397.t201 10.5154
R47812 a_71281_n8397.t192 a_71281_n8397.n322 10.5154
R47813 a_71281_n8397.n326 a_71281_n8397.t192 10.5154
R47814 a_71281_n8397.t260 a_71281_n8397.n336 10.5154
R47815 a_71281_n8397.n340 a_71281_n8397.t260 10.5154
R47816 a_71281_n8397.t248 a_71281_n8397.n353 10.5154
R47817 a_71281_n8397.n357 a_71281_n8397.t248 10.5154
R47818 a_71281_n8397.t316 a_71281_n8397.n367 10.5154
R47819 a_71281_n8397.n371 a_71281_n8397.t316 10.5154
R47820 a_71281_n8397.t293 a_71281_n8397.n384 10.5154
R47821 a_71281_n8397.n388 a_71281_n8397.t293 10.5154
R47822 a_71281_n8397.t110 a_71281_n8397.n398 10.5154
R47823 a_71281_n8397.n402 a_71281_n8397.t110 10.5154
R47824 a_71281_n8397.n576 a_71281_n8397.t304 10.5154
R47825 a_71281_n8397.t304 a_71281_n8397.n571 10.5154
R47826 a_71281_n8397.n562 a_71281_n8397.t123 10.5154
R47827 a_71281_n8397.t123 a_71281_n8397.n557 10.5154
R47828 a_71281_n8397.n548 a_71281_n8397.t95 10.5154
R47829 a_71281_n8397.t95 a_71281_n8397.n543 10.5154
R47830 a_71281_n8397.n534 a_71281_n8397.t108 10.5154
R47831 a_71281_n8397.t108 a_71281_n8397.n529 10.5154
R47832 a_71281_n8397.n517 a_71281_n8397.t94 10.5154
R47833 a_71281_n8397.t94 a_71281_n8397.n512 10.5154
R47834 a_71281_n8397.n503 a_71281_n8397.t168 10.5154
R47835 a_71281_n8397.t168 a_71281_n8397.n498 10.5154
R47836 a_71281_n8397.n486 a_71281_n8397.t162 10.5154
R47837 a_71281_n8397.t162 a_71281_n8397.n481 10.5154
R47838 a_71281_n8397.n472 a_71281_n8397.t232 10.5154
R47839 a_71281_n8397.t232 a_71281_n8397.n467 10.5154
R47840 a_71281_n8397.t290 a_71281_n8397.n733 10.5154
R47841 a_71281_n8397.n737 a_71281_n8397.t290 10.5154
R47842 a_71281_n8397.t104 a_71281_n8397.n747 10.5154
R47843 a_71281_n8397.n751 a_71281_n8397.t104 10.5154
R47844 a_71281_n8397.t79 a_71281_n8397.n761 10.5154
R47845 a_71281_n8397.n765 a_71281_n8397.t79 10.5154
R47846 a_71281_n8397.t87 a_71281_n8397.n775 10.5154
R47847 a_71281_n8397.n779 a_71281_n8397.t87 10.5154
R47848 a_71281_n8397.n866 a_71281_n8397.t78 10.5154
R47849 a_71281_n8397.t78 a_71281_n8397.n861 10.5154
R47850 a_71281_n8397.n852 a_71281_n8397.t153 10.5154
R47851 a_71281_n8397.t153 a_71281_n8397.n847 10.5154
R47852 a_71281_n8397.n835 a_71281_n8397.t149 10.5154
R47853 a_71281_n8397.t149 a_71281_n8397.n830 10.5154
R47854 a_71281_n8397.n821 a_71281_n8397.t220 10.5154
R47855 a_71281_n8397.t220 a_71281_n8397.n816 10.5154
R47856 a_71281_n8397.n589 a_71281_n8397.t206 10.515
R47857 a_71281_n8397.n5 a_71281_n8397.t269 10.515
R47858 a_71281_n8397.n282 a_71281_n8397.t312 10.515
R47859 a_71281_n8397.n296 a_71281_n8397.t226 10.515
R47860 a_71281_n8397.n573 a_71281_n8397.t225 10.515
R47861 a_71281_n8397.n734 a_71281_n8397.t223 10.515
R47862 a_71281_n8397.n706 a_71281_n8397.t176 10.515
R47863 a_71281_n8397.n707 a_71281_n8397.t176 10.515
R47864 a_71281_n8397.n720 a_71281_n8397.t245 10.515
R47865 a_71281_n8397.n721 a_71281_n8397.t245 10.515
R47866 a_71281_n8397.n804 a_71281_n8397.t273 10.515
R47867 a_71281_n8397.n803 a_71281_n8397.t273 10.515
R47868 a_71281_n8397.n791 a_71281_n8397.t337 10.515
R47869 a_71281_n8397.n790 a_71281_n8397.t337 10.515
R47870 a_71281_n8397.n590 a_71281_n8397.t206 10.515
R47871 a_71281_n8397.n603 a_71281_n8397.t270 10.515
R47872 a_71281_n8397.n602 a_71281_n8397.t270 10.515
R47873 a_71281_n8397.n617 a_71281_n8397.t263 10.515
R47874 a_71281_n8397.n616 a_71281_n8397.t263 10.515
R47875 a_71281_n8397.n631 a_71281_n8397.t329 10.515
R47876 a_71281_n8397.n630 a_71281_n8397.t329 10.515
R47877 a_71281_n8397.n648 a_71281_n8397.t322 10.515
R47878 a_71281_n8397.n647 a_71281_n8397.t322 10.515
R47879 a_71281_n8397.n662 a_71281_n8397.t137 10.515
R47880 a_71281_n8397.n661 a_71281_n8397.t137 10.515
R47881 a_71281_n8397.n679 a_71281_n8397.t115 10.515
R47882 a_71281_n8397.n678 a_71281_n8397.t115 10.515
R47883 a_71281_n8397.n693 a_71281_n8397.t185 10.515
R47884 a_71281_n8397.n692 a_71281_n8397.t185 10.515
R47885 a_71281_n8397.n122 a_71281_n8397.t242 10.515
R47886 a_71281_n8397.n123 a_71281_n8397.t242 10.515
R47887 a_71281_n8397.n136 a_71281_n8397.t309 10.515
R47888 a_71281_n8397.n137 a_71281_n8397.t309 10.515
R47889 a_71281_n8397.n164 a_71281_n8397.t111 10.515
R47890 a_71281_n8397.n163 a_71281_n8397.t111 10.515
R47891 a_71281_n8397.n151 a_71281_n8397.t178 10.515
R47892 a_71281_n8397.n150 a_71281_n8397.t178 10.515
R47893 a_71281_n8397.n6 a_71281_n8397.t269 10.515
R47894 a_71281_n8397.n19 a_71281_n8397.t335 10.515
R47895 a_71281_n8397.n18 a_71281_n8397.t335 10.515
R47896 a_71281_n8397.n33 a_71281_n8397.t328 10.515
R47897 a_71281_n8397.n32 a_71281_n8397.t328 10.515
R47898 a_71281_n8397.n47 a_71281_n8397.t141 10.515
R47899 a_71281_n8397.n46 a_71281_n8397.t141 10.515
R47900 a_71281_n8397.n64 a_71281_n8397.t134 10.515
R47901 a_71281_n8397.n63 a_71281_n8397.t134 10.515
R47902 a_71281_n8397.n78 a_71281_n8397.t210 10.515
R47903 a_71281_n8397.n77 a_71281_n8397.t210 10.515
R47904 a_71281_n8397.n95 a_71281_n8397.t184 10.515
R47905 a_71281_n8397.n94 a_71281_n8397.t184 10.515
R47906 a_71281_n8397.n109 a_71281_n8397.t252 10.515
R47907 a_71281_n8397.n108 a_71281_n8397.t252 10.515
R47908 a_71281_n8397.n281 a_71281_n8397.t312 10.515
R47909 a_71281_n8397.n267 a_71281_n8397.t129 10.515
R47910 a_71281_n8397.n268 a_71281_n8397.t129 10.515
R47911 a_71281_n8397.n253 a_71281_n8397.t105 10.515
R47912 a_71281_n8397.n254 a_71281_n8397.t105 10.515
R47913 a_71281_n8397.n239 a_71281_n8397.t116 10.515
R47914 a_71281_n8397.n240 a_71281_n8397.t116 10.515
R47915 a_71281_n8397.n222 a_71281_n8397.t103 10.515
R47916 a_71281_n8397.n223 a_71281_n8397.t103 10.515
R47917 a_71281_n8397.n208 a_71281_n8397.t177 10.515
R47918 a_71281_n8397.n209 a_71281_n8397.t177 10.515
R47919 a_71281_n8397.n191 a_71281_n8397.t164 10.515
R47920 a_71281_n8397.n192 a_71281_n8397.t164 10.515
R47921 a_71281_n8397.n177 a_71281_n8397.t236 10.515
R47922 a_71281_n8397.n178 a_71281_n8397.t236 10.515
R47923 a_71281_n8397.n413 a_71281_n8397.t207 10.515
R47924 a_71281_n8397.n414 a_71281_n8397.t207 10.515
R47925 a_71281_n8397.n427 a_71281_n8397.t274 10.515
R47926 a_71281_n8397.n428 a_71281_n8397.t274 10.515
R47927 a_71281_n8397.n455 a_71281_n8397.t276 10.515
R47928 a_71281_n8397.n454 a_71281_n8397.t276 10.515
R47929 a_71281_n8397.n442 a_71281_n8397.t75 10.515
R47930 a_71281_n8397.n441 a_71281_n8397.t75 10.515
R47931 a_71281_n8397.n297 a_71281_n8397.t226 10.515
R47932 a_71281_n8397.n310 a_71281_n8397.t289 10.515
R47933 a_71281_n8397.n309 a_71281_n8397.t289 10.515
R47934 a_71281_n8397.n324 a_71281_n8397.t283 10.515
R47935 a_71281_n8397.n323 a_71281_n8397.t283 10.515
R47936 a_71281_n8397.n338 a_71281_n8397.t90 10.515
R47937 a_71281_n8397.n337 a_71281_n8397.t90 10.515
R47938 a_71281_n8397.n355 a_71281_n8397.t85 10.515
R47939 a_71281_n8397.n354 a_71281_n8397.t85 10.515
R47940 a_71281_n8397.n369 a_71281_n8397.t158 10.515
R47941 a_71281_n8397.n368 a_71281_n8397.t158 10.515
R47942 a_71281_n8397.n386 a_71281_n8397.t139 10.515
R47943 a_71281_n8397.n385 a_71281_n8397.t139 10.515
R47944 a_71281_n8397.n400 a_71281_n8397.t213 10.515
R47945 a_71281_n8397.n399 a_71281_n8397.t213 10.515
R47946 a_71281_n8397.n572 a_71281_n8397.t225 10.515
R47947 a_71281_n8397.n558 a_71281_n8397.t285 10.515
R47948 a_71281_n8397.n559 a_71281_n8397.t285 10.515
R47949 a_71281_n8397.n544 a_71281_n8397.t272 10.515
R47950 a_71281_n8397.n545 a_71281_n8397.t272 10.515
R47951 a_71281_n8397.n530 a_71281_n8397.t280 10.515
R47952 a_71281_n8397.n531 a_71281_n8397.t280 10.515
R47953 a_71281_n8397.n513 a_71281_n8397.t271 10.515
R47954 a_71281_n8397.n514 a_71281_n8397.t271 10.515
R47955 a_71281_n8397.n499 a_71281_n8397.t336 10.515
R47956 a_71281_n8397.n500 a_71281_n8397.t336 10.515
R47957 a_71281_n8397.n482 a_71281_n8397.t330 10.515
R47958 a_71281_n8397.n483 a_71281_n8397.t330 10.515
R47959 a_71281_n8397.n468 a_71281_n8397.t142 10.515
R47960 a_71281_n8397.n469 a_71281_n8397.t142 10.515
R47961 a_71281_n8397.n735 a_71281_n8397.t223 10.515
R47962 a_71281_n8397.n749 a_71281_n8397.t284 10.515
R47963 a_71281_n8397.n748 a_71281_n8397.t284 10.515
R47964 a_71281_n8397.n763 a_71281_n8397.t267 10.515
R47965 a_71281_n8397.n762 a_71281_n8397.t267 10.515
R47966 a_71281_n8397.n777 a_71281_n8397.t279 10.515
R47967 a_71281_n8397.n776 a_71281_n8397.t279 10.515
R47968 a_71281_n8397.n862 a_71281_n8397.t266 10.515
R47969 a_71281_n8397.n863 a_71281_n8397.t266 10.515
R47970 a_71281_n8397.n848 a_71281_n8397.t334 10.515
R47971 a_71281_n8397.n849 a_71281_n8397.t334 10.515
R47972 a_71281_n8397.n831 a_71281_n8397.t327 10.515
R47973 a_71281_n8397.n832 a_71281_n8397.t327 10.515
R47974 a_71281_n8397.n817 a_71281_n8397.t140 10.515
R47975 a_71281_n8397.n818 a_71281_n8397.t140 10.515
R47976 a_71281_n8397.n710 a_71281_n8397.t296 9.57886
R47977 a_71281_n8397.t296 a_71281_n8397.n705 9.57886
R47978 a_71281_n8397.n707 a_71281_n8397.t228 9.57886
R47979 a_71281_n8397.t228 a_71281_n8397.n706 9.57886
R47980 a_71281_n8397.n724 a_71281_n8397.t112 9.57886
R47981 a_71281_n8397.t112 a_71281_n8397.n719 9.57886
R47982 a_71281_n8397.n721 a_71281_n8397.t297 9.57886
R47983 a_71281_n8397.t297 a_71281_n8397.n720 9.57886
R47984 a_71281_n8397.t186 a_71281_n8397.n802 9.57886
R47985 a_71281_n8397.n806 a_71281_n8397.t186 9.57886
R47986 a_71281_n8397.t174 a_71281_n8397.n803 9.57886
R47987 a_71281_n8397.n804 a_71281_n8397.t174 9.57886
R47988 a_71281_n8397.t254 a_71281_n8397.n789 9.57886
R47989 a_71281_n8397.n793 a_71281_n8397.t254 9.57886
R47990 a_71281_n8397.t243 a_71281_n8397.n790 9.57886
R47991 a_71281_n8397.n791 a_71281_n8397.t243 9.57886
R47992 a_71281_n8397.t321 a_71281_n8397.n588 9.57886
R47993 a_71281_n8397.n592 a_71281_n8397.t321 9.57886
R47994 a_71281_n8397.t256 a_71281_n8397.n589 9.57886
R47995 a_71281_n8397.n590 a_71281_n8397.t256 9.57886
R47996 a_71281_n8397.t136 a_71281_n8397.n601 9.57886
R47997 a_71281_n8397.n605 a_71281_n8397.t136 9.57886
R47998 a_71281_n8397.t323 a_71281_n8397.n602 9.57886
R47999 a_71281_n8397.n603 a_71281_n8397.t323 9.57886
R48000 a_71281_n8397.t128 a_71281_n8397.n615 9.57886
R48001 a_71281_n8397.n619 a_71281_n8397.t128 9.57886
R48002 a_71281_n8397.t313 a_71281_n8397.n616 9.57886
R48003 a_71281_n8397.n617 a_71281_n8397.t313 9.57886
R48004 a_71281_n8397.t203 a_71281_n8397.n629 9.57886
R48005 a_71281_n8397.n633 a_71281_n8397.t203 9.57886
R48006 a_71281_n8397.t130 a_71281_n8397.n630 9.57886
R48007 a_71281_n8397.n631 a_71281_n8397.t130 9.57886
R48008 a_71281_n8397.t32 a_71281_n8397.n646 9.57886
R48009 a_71281_n8397.n650 a_71281_n8397.t32 9.57886
R48010 a_71281_n8397.t58 a_71281_n8397.n647 9.57886
R48011 a_71281_n8397.n648 a_71281_n8397.t58 9.57886
R48012 a_71281_n8397.t12 a_71281_n8397.n660 9.57886
R48013 a_71281_n8397.n664 a_71281_n8397.t12 9.57886
R48014 a_71281_n8397.t30 a_71281_n8397.n661 9.57886
R48015 a_71281_n8397.n662 a_71281_n8397.t30 9.57886
R48016 a_71281_n8397.t235 a_71281_n8397.n677 9.57886
R48017 a_71281_n8397.n681 a_71281_n8397.t235 9.57886
R48018 a_71281_n8397.t165 a_71281_n8397.n678 9.57886
R48019 a_71281_n8397.n679 a_71281_n8397.t165 9.57886
R48020 a_71281_n8397.t302 a_71281_n8397.n691 9.57886
R48021 a_71281_n8397.n695 a_71281_n8397.t302 9.57886
R48022 a_71281_n8397.t237 a_71281_n8397.n692 9.57886
R48023 a_71281_n8397.n693 a_71281_n8397.t237 9.57886
R48024 a_71281_n8397.n126 a_71281_n8397.t118 9.57886
R48025 a_71281_n8397.t118 a_71281_n8397.n121 9.57886
R48026 a_71281_n8397.n123 a_71281_n8397.t217 9.57886
R48027 a_71281_n8397.t217 a_71281_n8397.n122 9.57886
R48028 a_71281_n8397.n140 a_71281_n8397.t191 9.57886
R48029 a_71281_n8397.t191 a_71281_n8397.n135 9.57886
R48030 a_71281_n8397.n137 a_71281_n8397.t282 9.57886
R48031 a_71281_n8397.t282 a_71281_n8397.n136 9.57886
R48032 a_71281_n8397.t187 a_71281_n8397.n162 9.57886
R48033 a_71281_n8397.n166 a_71281_n8397.t187 9.57886
R48034 a_71281_n8397.t298 a_71281_n8397.n163 9.57886
R48035 a_71281_n8397.n164 a_71281_n8397.t298 9.57886
R48036 a_71281_n8397.t255 a_71281_n8397.n149 9.57886
R48037 a_71281_n8397.n153 a_71281_n8397.t255 9.57886
R48038 a_71281_n8397.t113 a_71281_n8397.n150 9.57886
R48039 a_71281_n8397.n151 a_71281_n8397.t113 9.57886
R48040 a_71281_n8397.t144 a_71281_n8397.n4 9.57886
R48041 a_71281_n8397.n8 a_71281_n8397.t144 9.57886
R48042 a_71281_n8397.t234 a_71281_n8397.n5 9.57886
R48043 a_71281_n8397.n6 a_71281_n8397.t234 9.57886
R48044 a_71281_n8397.t216 a_71281_n8397.n17 9.57886
R48045 a_71281_n8397.n21 a_71281_n8397.t216 9.57886
R48046 a_71281_n8397.t300 a_71281_n8397.n18 9.57886
R48047 a_71281_n8397.n19 a_71281_n8397.t300 9.57886
R48048 a_71281_n8397.t212 a_71281_n8397.n31 9.57886
R48049 a_71281_n8397.n35 a_71281_n8397.t212 9.57886
R48050 a_71281_n8397.t292 a_71281_n8397.n32 9.57886
R48051 a_71281_n8397.n33 a_71281_n8397.t292 9.57886
R48052 a_71281_n8397.t278 a_71281_n8397.n45 9.57886
R48053 a_71281_n8397.n49 a_71281_n8397.t278 9.57886
R48054 a_71281_n8397.t109 a_71281_n8397.n46 9.57886
R48055 a_71281_n8397.n47 a_71281_n8397.t109 9.57886
R48056 a_71281_n8397.t8 a_71281_n8397.n62 9.57886
R48057 a_71281_n8397.n66 a_71281_n8397.t8 9.57886
R48058 a_71281_n8397.t64 a_71281_n8397.n63 9.57886
R48059 a_71281_n8397.n64 a_71281_n8397.t64 9.57886
R48060 a_71281_n8397.t0 a_71281_n8397.n76 9.57886
R48061 a_71281_n8397.n80 a_71281_n8397.t0 9.57886
R48062 a_71281_n8397.t44 a_71281_n8397.n77 9.57886
R48063 a_71281_n8397.n78 a_71281_n8397.t44 9.57886
R48064 a_71281_n8397.t310 a_71281_n8397.n93 9.57886
R48065 a_71281_n8397.n97 a_71281_n8397.t310 9.57886
R48066 a_71281_n8397.t152 a_71281_n8397.n94 9.57886
R48067 a_71281_n8397.n95 a_71281_n8397.t152 9.57886
R48068 a_71281_n8397.t125 a_71281_n8397.n107 9.57886
R48069 a_71281_n8397.n111 a_71281_n8397.t125 9.57886
R48070 a_71281_n8397.t224 a_71281_n8397.n108 9.57886
R48071 a_71281_n8397.n109 a_71281_n8397.t224 9.57886
R48072 a_71281_n8397.n285 a_71281_n8397.t133 9.57886
R48073 a_71281_n8397.t133 a_71281_n8397.n280 9.57886
R48074 a_71281_n8397.n282 a_71281_n8397.t249 9.57886
R48075 a_71281_n8397.t249 a_71281_n8397.n281 9.57886
R48076 a_71281_n8397.n271 a_71281_n8397.t209 9.57886
R48077 a_71281_n8397.t209 a_71281_n8397.n266 9.57886
R48078 a_71281_n8397.n268 a_71281_n8397.t317 9.57886
R48079 a_71281_n8397.t317 a_71281_n8397.n267 9.57886
R48080 a_71281_n8397.n257 a_71281_n8397.t183 9.57886
R48081 a_71281_n8397.t183 a_71281_n8397.n252 9.57886
R48082 a_71281_n8397.n254 a_71281_n8397.t294 9.57886
R48083 a_71281_n8397.t294 a_71281_n8397.n253 9.57886
R48084 a_71281_n8397.n243 a_71281_n8397.t196 9.57886
R48085 a_71281_n8397.t196 a_71281_n8397.n238 9.57886
R48086 a_71281_n8397.n240 a_71281_n8397.t301 9.57886
R48087 a_71281_n8397.t301 a_71281_n8397.n239 9.57886
R48088 a_71281_n8397.n226 a_71281_n8397.t36 9.57886
R48089 a_71281_n8397.t36 a_71281_n8397.n221 9.57886
R48090 a_71281_n8397.n223 a_71281_n8397.t4 9.57886
R48091 a_71281_n8397.t4 a_71281_n8397.n222 9.57886
R48092 a_71281_n8397.n212 a_71281_n8397.t14 9.57886
R48093 a_71281_n8397.t14 a_71281_n8397.n207 9.57886
R48094 a_71281_n8397.n209 a_71281_n8397.t62 9.57886
R48095 a_71281_n8397.t62 a_71281_n8397.n208 9.57886
R48096 a_71281_n8397.n195 a_71281_n8397.t240 9.57886
R48097 a_71281_n8397.t240 a_71281_n8397.n190 9.57886
R48098 a_71281_n8397.n192 a_71281_n8397.t96 9.57886
R48099 a_71281_n8397.t96 a_71281_n8397.n191 9.57886
R48100 a_71281_n8397.n181 a_71281_n8397.t307 9.57886
R48101 a_71281_n8397.t307 a_71281_n8397.n176 9.57886
R48102 a_71281_n8397.n178 a_71281_n8397.t169 9.57886
R48103 a_71281_n8397.t169 a_71281_n8397.n177 9.57886
R48104 a_71281_n8397.n417 a_71281_n8397.t331 9.57886
R48105 a_71281_n8397.t331 a_71281_n8397.n412 9.57886
R48106 a_71281_n8397.n414 a_71281_n8397.t161 9.57886
R48107 a_71281_n8397.t161 a_71281_n8397.n413 9.57886
R48108 a_71281_n8397.n431 a_71281_n8397.t145 9.57886
R48109 a_71281_n8397.t145 a_71281_n8397.n426 9.57886
R48110 a_71281_n8397.n428 a_71281_n8397.t231 9.57886
R48111 a_71281_n8397.t231 a_71281_n8397.n427 9.57886
R48112 a_71281_n8397.t84 a_71281_n8397.n453 9.57886
R48113 a_71281_n8397.n457 a_71281_n8397.t84 9.57886
R48114 a_71281_n8397.t117 a_71281_n8397.n454 9.57886
R48115 a_71281_n8397.n455 a_71281_n8397.t117 9.57886
R48116 a_71281_n8397.t157 a_71281_n8397.n440 9.57886
R48117 a_71281_n8397.n444 a_71281_n8397.t157 9.57886
R48118 a_71281_n8397.t188 a_71281_n8397.n441 9.57886
R48119 a_71281_n8397.n442 a_71281_n8397.t188 9.57886
R48120 a_71281_n8397.t91 a_71281_n8397.n295 9.57886
R48121 a_71281_n8397.n299 a_71281_n8397.t91 9.57886
R48122 a_71281_n8397.t190 a_71281_n8397.n296 9.57886
R48123 a_71281_n8397.n297 a_71281_n8397.t190 9.57886
R48124 a_71281_n8397.t166 a_71281_n8397.n308 9.57886
R48125 a_71281_n8397.n312 a_71281_n8397.t166 9.57886
R48126 a_71281_n8397.t258 a_71281_n8397.n309 9.57886
R48127 a_71281_n8397.n310 a_71281_n8397.t258 9.57886
R48128 a_71281_n8397.t160 a_71281_n8397.n322 9.57886
R48129 a_71281_n8397.n326 a_71281_n8397.t160 9.57886
R48130 a_71281_n8397.t247 a_71281_n8397.n323 9.57886
R48131 a_71281_n8397.n324 a_71281_n8397.t247 9.57886
R48132 a_71281_n8397.t230 a_71281_n8397.n336 9.57886
R48133 a_71281_n8397.n340 a_71281_n8397.t230 9.57886
R48134 a_71281_n8397.t315 a_71281_n8397.n337 9.57886
R48135 a_71281_n8397.n338 a_71281_n8397.t315 9.57886
R48136 a_71281_n8397.t22 a_71281_n8397.n353 9.57886
R48137 a_71281_n8397.n357 a_71281_n8397.t22 9.57886
R48138 a_71281_n8397.t2 a_71281_n8397.n354 9.57886
R48139 a_71281_n8397.n355 a_71281_n8397.t2 9.57886
R48140 a_71281_n8397.t6 a_71281_n8397.n367 9.57886
R48141 a_71281_n8397.n371 a_71281_n8397.t6 9.57886
R48142 a_71281_n8397.t56 a_71281_n8397.n368 9.57886
R48143 a_71281_n8397.n369 a_71281_n8397.t56 9.57886
R48144 a_71281_n8397.t275 a_71281_n8397.n384 9.57886
R48145 a_71281_n8397.n388 a_71281_n8397.t275 9.57886
R48146 a_71281_n8397.t93 a_71281_n8397.n385 9.57886
R48147 a_71281_n8397.n386 a_71281_n8397.t93 9.57886
R48148 a_71281_n8397.t74 a_71281_n8397.n398 9.57886
R48149 a_71281_n8397.n402 a_71281_n8397.t74 9.57886
R48150 a_71281_n8397.t167 a_71281_n8397.n399 9.57886
R48151 a_71281_n8397.n400 a_71281_n8397.t167 9.57886
R48152 a_71281_n8397.n576 a_71281_n8397.t291 9.57886
R48153 a_71281_n8397.t291 a_71281_n8397.n571 9.57886
R48154 a_71281_n8397.n573 a_71281_n8397.t320 9.57886
R48155 a_71281_n8397.t320 a_71281_n8397.n572 9.57886
R48156 a_71281_n8397.n562 a_71281_n8397.t106 9.57886
R48157 a_71281_n8397.t106 a_71281_n8397.n557 9.57886
R48158 a_71281_n8397.n559 a_71281_n8397.t135 9.57886
R48159 a_71281_n8397.t135 a_71281_n8397.n558 9.57886
R48160 a_71281_n8397.n548 a_71281_n8397.t80 9.57886
R48161 a_71281_n8397.t80 a_71281_n8397.n543 9.57886
R48162 a_71281_n8397.n545 a_71281_n8397.t114 9.57886
R48163 a_71281_n8397.t114 a_71281_n8397.n544 9.57886
R48164 a_71281_n8397.n534 a_71281_n8397.t88 9.57886
R48165 a_71281_n8397.t88 a_71281_n8397.n529 9.57886
R48166 a_71281_n8397.n531 a_71281_n8397.t122 9.57886
R48167 a_71281_n8397.t122 a_71281_n8397.n530 9.57886
R48168 a_71281_n8397.n517 a_71281_n8397.t68 9.57886
R48169 a_71281_n8397.t68 a_71281_n8397.n512 9.57886
R48170 a_71281_n8397.n514 a_71281_n8397.t60 9.57886
R48171 a_71281_n8397.t60 a_71281_n8397.n513 9.57886
R48172 a_71281_n8397.n503 a_71281_n8397.t48 9.57886
R48173 a_71281_n8397.t48 a_71281_n8397.n498 9.57886
R48174 a_71281_n8397.n500 a_71281_n8397.t34 9.57886
R48175 a_71281_n8397.t34 a_71281_n8397.n499 9.57886
R48176 a_71281_n8397.n486 a_71281_n8397.t150 9.57886
R48177 a_71281_n8397.t150 a_71281_n8397.n481 9.57886
R48178 a_71281_n8397.n483 a_71281_n8397.t175 9.57886
R48179 a_71281_n8397.t175 a_71281_n8397.n482 9.57886
R48180 a_71281_n8397.n472 a_71281_n8397.t221 9.57886
R48181 a_71281_n8397.t221 a_71281_n8397.n467 9.57886
R48182 a_71281_n8397.n469 a_71281_n8397.t244 9.57886
R48183 a_71281_n8397.t244 a_71281_n8397.n468 9.57886
R48184 a_71281_n8397.t132 a_71281_n8397.n733 9.57886
R48185 a_71281_n8397.n737 a_71281_n8397.t132 9.57886
R48186 a_71281_n8397.t124 a_71281_n8397.n734 9.57886
R48187 a_71281_n8397.n735 a_71281_n8397.t124 9.57886
R48188 a_71281_n8397.t208 a_71281_n8397.n747 9.57886
R48189 a_71281_n8397.n751 a_71281_n8397.t208 9.57886
R48190 a_71281_n8397.t199 a_71281_n8397.n748 9.57886
R48191 a_71281_n8397.n749 a_71281_n8397.t199 9.57886
R48192 a_71281_n8397.t181 a_71281_n8397.n761 9.57886
R48193 a_71281_n8397.n765 a_71281_n8397.t181 9.57886
R48194 a_71281_n8397.t171 a_71281_n8397.n762 9.57886
R48195 a_71281_n8397.n763 a_71281_n8397.t171 9.57886
R48196 a_71281_n8397.t194 a_71281_n8397.n775 9.57886
R48197 a_71281_n8397.n779 a_71281_n8397.t194 9.57886
R48198 a_71281_n8397.t179 a_71281_n8397.n776 9.57886
R48199 a_71281_n8397.n777 a_71281_n8397.t179 9.57886
R48200 a_71281_n8397.n866 a_71281_n8397.t38 9.57886
R48201 a_71281_n8397.t38 a_71281_n8397.n861 9.57886
R48202 a_71281_n8397.n863 a_71281_n8397.t42 9.57886
R48203 a_71281_n8397.t42 a_71281_n8397.n862 9.57886
R48204 a_71281_n8397.n852 a_71281_n8397.t16 9.57886
R48205 a_71281_n8397.t16 a_71281_n8397.n847 9.57886
R48206 a_71281_n8397.n849 a_71281_n8397.t20 9.57886
R48207 a_71281_n8397.t20 a_71281_n8397.n848 9.57886
R48208 a_71281_n8397.n835 a_71281_n8397.t239 9.57886
R48209 a_71281_n8397.t239 a_71281_n8397.n830 9.57886
R48210 a_71281_n8397.n832 a_71281_n8397.t233 9.57886
R48211 a_71281_n8397.t233 a_71281_n8397.n831 9.57886
R48212 a_71281_n8397.n821 a_71281_n8397.t306 9.57886
R48213 a_71281_n8397.t306 a_71281_n8397.n816 9.57886
R48214 a_71281_n8397.n818 a_71281_n8397.t299 9.57886
R48215 a_71281_n8397.t299 a_71281_n8397.n817 9.57886
R48216 a_71281_n8397.t238 a_71281_n8397.n712 8.10567
R48217 a_71281_n8397.n713 a_71281_n8397.t238 8.10567
R48218 a_71281_n8397.t305 a_71281_n8397.n726 8.10567
R48219 a_71281_n8397.n727 a_71281_n8397.t305 8.10567
R48220 a_71281_n8397.n810 a_71281_n8397.t82 8.10567
R48221 a_71281_n8397.t82 a_71281_n8397.n809 8.10567
R48222 a_71281_n8397.n796 a_71281_n8397.t155 8.10567
R48223 a_71281_n8397.t155 a_71281_n8397.n795 8.10567
R48224 a_71281_n8397.n595 a_71281_n8397.t265 8.10567
R48225 a_71281_n8397.t265 a_71281_n8397.n594 8.10567
R48226 a_71281_n8397.n609 a_71281_n8397.t333 8.10567
R48227 a_71281_n8397.t333 a_71281_n8397.n608 8.10567
R48228 a_71281_n8397.n623 a_71281_n8397.t325 8.10567
R48229 a_71281_n8397.t325 a_71281_n8397.n622 8.10567
R48230 a_71281_n8397.n637 a_71281_n8397.t138 8.10567
R48231 a_71281_n8397.t138 a_71281_n8397.n636 8.10567
R48232 a_71281_n8397.n654 a_71281_n8397.t54 8.10567
R48233 a_71281_n8397.t54 a_71281_n8397.n653 8.10567
R48234 a_71281_n8397.n668 a_71281_n8397.t26 8.10567
R48235 a_71281_n8397.t26 a_71281_n8397.n667 8.10567
R48236 a_71281_n8397.n685 a_71281_n8397.t180 8.10567
R48237 a_71281_n8397.t180 a_71281_n8397.n684 8.10567
R48238 a_71281_n8397.n699 a_71281_n8397.t250 8.10567
R48239 a_71281_n8397.t250 a_71281_n8397.n698 8.10567
R48240 a_71281_n8397.t286 a_71281_n8397.n128 8.10567
R48241 a_71281_n8397.n129 a_71281_n8397.t286 8.10567
R48242 a_71281_n8397.t98 a_71281_n8397.n142 8.10567
R48243 a_71281_n8397.n143 a_71281_n8397.t98 8.10567
R48244 a_71281_n8397.n170 a_71281_n8397.t205 8.10567
R48245 a_71281_n8397.t205 a_71281_n8397.n169 8.10567
R48246 a_71281_n8397.n156 a_71281_n8397.t268 8.10567
R48247 a_71281_n8397.t268 a_71281_n8397.n155 8.10567
R48248 a_71281_n8397.n11 a_71281_n8397.t311 8.10567
R48249 a_71281_n8397.t311 a_71281_n8397.n10 8.10567
R48250 a_71281_n8397.n25 a_71281_n8397.t127 8.10567
R48251 a_71281_n8397.t127 a_71281_n8397.n24 8.10567
R48252 a_71281_n8397.n39 a_71281_n8397.t119 8.10567
R48253 a_71281_n8397.t119 a_71281_n8397.n38 8.10567
R48254 a_71281_n8397.n53 a_71281_n8397.t193 8.10567
R48255 a_71281_n8397.t193 a_71281_n8397.n52 8.10567
R48256 a_71281_n8397.n70 a_71281_n8397.t40 8.10567
R48257 a_71281_n8397.t40 a_71281_n8397.n69 8.10567
R48258 a_71281_n8397.n84 a_71281_n8397.t18 8.10567
R48259 a_71281_n8397.t18 a_71281_n8397.n83 8.10567
R48260 a_71281_n8397.n101 a_71281_n8397.t227 8.10567
R48261 a_71281_n8397.t227 a_71281_n8397.n100 8.10567
R48262 a_71281_n8397.n115 a_71281_n8397.t295 8.10567
R48263 a_71281_n8397.t295 a_71281_n8397.n114 8.10567
R48264 a_71281_n8397.t148 a_71281_n8397.n287 8.10567
R48265 a_71281_n8397.n288 a_71281_n8397.t148 8.10567
R48266 a_71281_n8397.t219 a_71281_n8397.n273 8.10567
R48267 a_71281_n8397.n274 a_71281_n8397.t219 8.10567
R48268 a_71281_n8397.t202 a_71281_n8397.n259 8.10567
R48269 a_71281_n8397.n260 a_71281_n8397.t202 8.10567
R48270 a_71281_n8397.t211 a_71281_n8397.n245 8.10567
R48271 a_71281_n8397.n246 a_71281_n8397.t211 8.10567
R48272 a_71281_n8397.t28 a_71281_n8397.n228 8.10567
R48273 a_71281_n8397.n229 a_71281_n8397.t28 8.10567
R48274 a_71281_n8397.t10 a_71281_n8397.n214 8.10567
R48275 a_71281_n8397.n215 a_71281_n8397.t10 8.10567
R48276 a_71281_n8397.t259 a_71281_n8397.n197 8.10567
R48277 a_71281_n8397.n198 a_71281_n8397.t259 8.10567
R48278 a_71281_n8397.t324 a_71281_n8397.n183 8.10567
R48279 a_71281_n8397.n184 a_71281_n8397.t324 8.10567
R48280 a_71281_n8397.t246 a_71281_n8397.n419 8.10567
R48281 a_71281_n8397.n420 a_71281_n8397.t246 8.10567
R48282 a_71281_n8397.t314 a_71281_n8397.n433 8.10567
R48283 a_71281_n8397.n434 a_71281_n8397.t314 8.10567
R48284 a_71281_n8397.n461 a_71281_n8397.t99 8.10567
R48285 a_71281_n8397.t99 a_71281_n8397.n460 8.10567
R48286 a_71281_n8397.n447 a_71281_n8397.t172 8.10567
R48287 a_71281_n8397.t172 a_71281_n8397.n446 8.10567
R48288 a_71281_n8397.n302 a_71281_n8397.t277 8.10567
R48289 a_71281_n8397.t277 a_71281_n8397.n301 8.10567
R48290 a_71281_n8397.n316 a_71281_n8397.t76 8.10567
R48291 a_71281_n8397.t76 a_71281_n8397.n315 8.10567
R48292 a_71281_n8397.n330 a_71281_n8397.t332 8.10567
R48293 a_71281_n8397.t332 a_71281_n8397.n329 8.10567
R48294 a_71281_n8397.n344 a_71281_n8397.t146 8.10567
R48295 a_71281_n8397.t146 a_71281_n8397.n343 8.10567
R48296 a_71281_n8397.n361 a_71281_n8397.t52 8.10567
R48297 a_71281_n8397.t52 a_71281_n8397.n360 8.10567
R48298 a_71281_n8397.n375 a_71281_n8397.t24 8.10567
R48299 a_71281_n8397.t24 a_71281_n8397.n374 8.10567
R48300 a_71281_n8397.n392 a_71281_n8397.t189 8.10567
R48301 a_71281_n8397.t189 a_71281_n8397.n391 8.10567
R48302 a_71281_n8397.n406 a_71281_n8397.t257 8.10567
R48303 a_71281_n8397.t257 a_71281_n8397.n405 8.10567
R48304 a_71281_n8397.t303 a_71281_n8397.n578 8.10567
R48305 a_71281_n8397.n579 a_71281_n8397.t303 8.10567
R48306 a_71281_n8397.t121 a_71281_n8397.n564 8.10567
R48307 a_71281_n8397.n565 a_71281_n8397.t121 8.10567
R48308 a_71281_n8397.t92 a_71281_n8397.n550 8.10567
R48309 a_71281_n8397.n551 a_71281_n8397.t92 8.10567
R48310 a_71281_n8397.t107 a_71281_n8397.n536 8.10567
R48311 a_71281_n8397.n537 a_71281_n8397.t107 8.10567
R48312 a_71281_n8397.t66 a_71281_n8397.n519 8.10567
R48313 a_71281_n8397.n520 a_71281_n8397.t66 8.10567
R48314 a_71281_n8397.t46 a_71281_n8397.n505 8.10567
R48315 a_71281_n8397.n506 a_71281_n8397.t46 8.10567
R48316 a_71281_n8397.t159 a_71281_n8397.n488 8.10567
R48317 a_71281_n8397.n489 a_71281_n8397.t159 8.10567
R48318 a_71281_n8397.t229 a_71281_n8397.n474 8.10567
R48319 a_71281_n8397.n475 a_71281_n8397.t229 8.10567
R48320 a_71281_n8397.n741 a_71281_n8397.t288 8.10567
R48321 a_71281_n8397.t288 a_71281_n8397.n740 8.10567
R48322 a_71281_n8397.n755 a_71281_n8397.t102 8.10567
R48323 a_71281_n8397.t102 a_71281_n8397.n754 8.10567
R48324 a_71281_n8397.n769 a_71281_n8397.t77 8.10567
R48325 a_71281_n8397.t77 a_71281_n8397.n768 8.10567
R48326 a_71281_n8397.n783 a_71281_n8397.t86 8.10567
R48327 a_71281_n8397.t86 a_71281_n8397.n782 8.10567
R48328 a_71281_n8397.t70 a_71281_n8397.n868 8.10567
R48329 a_71281_n8397.n869 a_71281_n8397.t70 8.10567
R48330 a_71281_n8397.t50 a_71281_n8397.n854 8.10567
R48331 a_71281_n8397.n855 a_71281_n8397.t50 8.10567
R48332 a_71281_n8397.t147 a_71281_n8397.n837 8.10567
R48333 a_71281_n8397.n838 a_71281_n8397.t147 8.10567
R48334 a_71281_n8397.t218 a_71281_n8397.n823 8.10567
R48335 a_71281_n8397.n824 a_71281_n8397.t218 8.10567
R48336 a_71281_n8397.n585 a_71281_n8397.t72 7.10686
R48337 a_71281_n8397.n673 a_71281_n8397.t13 6.12845
R48338 a_71281_n8397.n843 a_71281_n8397.t17 6.12845
R48339 a_71281_n8397.n89 a_71281_n8397.t1 6.12845
R48340 a_71281_n8397.n203 a_71281_n8397.t15 6.12845
R48341 a_71281_n8397.n380 a_71281_n8397.t7 6.12845
R48342 a_71281_n8397.n494 a_71281_n8397.t49 6.12845
R48343 a_71281_n8397.n874 a_71281_n8397.t43 6.12049
R48344 a_71281_n8397.n642 a_71281_n8397.t59 6.12049
R48345 a_71281_n8397.n58 a_71281_n8397.t65 6.12049
R48346 a_71281_n8397.n234 a_71281_n8397.t5 6.12049
R48347 a_71281_n8397.n349 a_71281_n8397.t3 6.12049
R48348 a_71281_n8397.n525 a_71281_n8397.t61 6.12049
R48349 a_71281_n8397.n712 a_71281_n8397.n708 4.64734
R48350 a_71281_n8397.n713 a_71281_n8397.n704 4.64734
R48351 a_71281_n8397.n726 a_71281_n8397.n722 4.64734
R48352 a_71281_n8397.n727 a_71281_n8397.n718 4.64734
R48353 a_71281_n8397.n810 a_71281_n8397.n801 4.64734
R48354 a_71281_n8397.n809 a_71281_n8397.n805 4.64734
R48355 a_71281_n8397.n796 a_71281_n8397.n788 4.64734
R48356 a_71281_n8397.n795 a_71281_n8397.n792 4.64734
R48357 a_71281_n8397.n595 a_71281_n8397.n587 4.64734
R48358 a_71281_n8397.n594 a_71281_n8397.n591 4.64734
R48359 a_71281_n8397.n609 a_71281_n8397.n600 4.64734
R48360 a_71281_n8397.n608 a_71281_n8397.n604 4.64734
R48361 a_71281_n8397.n623 a_71281_n8397.n614 4.64734
R48362 a_71281_n8397.n622 a_71281_n8397.n618 4.64734
R48363 a_71281_n8397.n637 a_71281_n8397.n628 4.64734
R48364 a_71281_n8397.n636 a_71281_n8397.n632 4.64734
R48365 a_71281_n8397.n654 a_71281_n8397.n645 4.64734
R48366 a_71281_n8397.n653 a_71281_n8397.n649 4.64734
R48367 a_71281_n8397.n668 a_71281_n8397.n659 4.64734
R48368 a_71281_n8397.n667 a_71281_n8397.n663 4.64734
R48369 a_71281_n8397.n685 a_71281_n8397.n676 4.64734
R48370 a_71281_n8397.n684 a_71281_n8397.n680 4.64734
R48371 a_71281_n8397.n699 a_71281_n8397.n690 4.64734
R48372 a_71281_n8397.n698 a_71281_n8397.n694 4.64734
R48373 a_71281_n8397.n128 a_71281_n8397.n124 4.64734
R48374 a_71281_n8397.n129 a_71281_n8397.n120 4.64734
R48375 a_71281_n8397.n142 a_71281_n8397.n138 4.64734
R48376 a_71281_n8397.n143 a_71281_n8397.n134 4.64734
R48377 a_71281_n8397.n170 a_71281_n8397.n161 4.64734
R48378 a_71281_n8397.n169 a_71281_n8397.n165 4.64734
R48379 a_71281_n8397.n156 a_71281_n8397.n148 4.64734
R48380 a_71281_n8397.n155 a_71281_n8397.n152 4.64734
R48381 a_71281_n8397.n11 a_71281_n8397.n3 4.64734
R48382 a_71281_n8397.n10 a_71281_n8397.n7 4.64734
R48383 a_71281_n8397.n25 a_71281_n8397.n16 4.64734
R48384 a_71281_n8397.n24 a_71281_n8397.n20 4.64734
R48385 a_71281_n8397.n39 a_71281_n8397.n30 4.64734
R48386 a_71281_n8397.n38 a_71281_n8397.n34 4.64734
R48387 a_71281_n8397.n53 a_71281_n8397.n44 4.64734
R48388 a_71281_n8397.n52 a_71281_n8397.n48 4.64734
R48389 a_71281_n8397.n70 a_71281_n8397.n61 4.64734
R48390 a_71281_n8397.n69 a_71281_n8397.n65 4.64734
R48391 a_71281_n8397.n84 a_71281_n8397.n75 4.64734
R48392 a_71281_n8397.n83 a_71281_n8397.n79 4.64734
R48393 a_71281_n8397.n101 a_71281_n8397.n92 4.64734
R48394 a_71281_n8397.n100 a_71281_n8397.n96 4.64734
R48395 a_71281_n8397.n115 a_71281_n8397.n106 4.64734
R48396 a_71281_n8397.n114 a_71281_n8397.n110 4.64734
R48397 a_71281_n8397.n287 a_71281_n8397.n283 4.64734
R48398 a_71281_n8397.n288 a_71281_n8397.n279 4.64734
R48399 a_71281_n8397.n273 a_71281_n8397.n269 4.64734
R48400 a_71281_n8397.n274 a_71281_n8397.n265 4.64734
R48401 a_71281_n8397.n259 a_71281_n8397.n255 4.64734
R48402 a_71281_n8397.n260 a_71281_n8397.n251 4.64734
R48403 a_71281_n8397.n245 a_71281_n8397.n241 4.64734
R48404 a_71281_n8397.n246 a_71281_n8397.n237 4.64734
R48405 a_71281_n8397.n228 a_71281_n8397.n224 4.64734
R48406 a_71281_n8397.n229 a_71281_n8397.n220 4.64734
R48407 a_71281_n8397.n214 a_71281_n8397.n210 4.64734
R48408 a_71281_n8397.n215 a_71281_n8397.n206 4.64734
R48409 a_71281_n8397.n197 a_71281_n8397.n193 4.64734
R48410 a_71281_n8397.n198 a_71281_n8397.n189 4.64734
R48411 a_71281_n8397.n183 a_71281_n8397.n179 4.64734
R48412 a_71281_n8397.n184 a_71281_n8397.n175 4.64734
R48413 a_71281_n8397.n419 a_71281_n8397.n415 4.64734
R48414 a_71281_n8397.n420 a_71281_n8397.n411 4.64734
R48415 a_71281_n8397.n433 a_71281_n8397.n429 4.64734
R48416 a_71281_n8397.n434 a_71281_n8397.n425 4.64734
R48417 a_71281_n8397.n461 a_71281_n8397.n452 4.64734
R48418 a_71281_n8397.n460 a_71281_n8397.n456 4.64734
R48419 a_71281_n8397.n447 a_71281_n8397.n439 4.64734
R48420 a_71281_n8397.n446 a_71281_n8397.n443 4.64734
R48421 a_71281_n8397.n302 a_71281_n8397.n294 4.64734
R48422 a_71281_n8397.n301 a_71281_n8397.n298 4.64734
R48423 a_71281_n8397.n316 a_71281_n8397.n307 4.64734
R48424 a_71281_n8397.n315 a_71281_n8397.n311 4.64734
R48425 a_71281_n8397.n330 a_71281_n8397.n321 4.64734
R48426 a_71281_n8397.n329 a_71281_n8397.n325 4.64734
R48427 a_71281_n8397.n344 a_71281_n8397.n335 4.64734
R48428 a_71281_n8397.n343 a_71281_n8397.n339 4.64734
R48429 a_71281_n8397.n361 a_71281_n8397.n352 4.64734
R48430 a_71281_n8397.n360 a_71281_n8397.n356 4.64734
R48431 a_71281_n8397.n375 a_71281_n8397.n366 4.64734
R48432 a_71281_n8397.n374 a_71281_n8397.n370 4.64734
R48433 a_71281_n8397.n392 a_71281_n8397.n383 4.64734
R48434 a_71281_n8397.n391 a_71281_n8397.n387 4.64734
R48435 a_71281_n8397.n406 a_71281_n8397.n397 4.64734
R48436 a_71281_n8397.n405 a_71281_n8397.n401 4.64734
R48437 a_71281_n8397.n578 a_71281_n8397.n574 4.64734
R48438 a_71281_n8397.n579 a_71281_n8397.n570 4.64734
R48439 a_71281_n8397.n564 a_71281_n8397.n560 4.64734
R48440 a_71281_n8397.n565 a_71281_n8397.n556 4.64734
R48441 a_71281_n8397.n550 a_71281_n8397.n546 4.64734
R48442 a_71281_n8397.n551 a_71281_n8397.n542 4.64734
R48443 a_71281_n8397.n536 a_71281_n8397.n532 4.64734
R48444 a_71281_n8397.n537 a_71281_n8397.n528 4.64734
R48445 a_71281_n8397.n519 a_71281_n8397.n515 4.64734
R48446 a_71281_n8397.n520 a_71281_n8397.n511 4.64734
R48447 a_71281_n8397.n505 a_71281_n8397.n501 4.64734
R48448 a_71281_n8397.n506 a_71281_n8397.n497 4.64734
R48449 a_71281_n8397.n488 a_71281_n8397.n484 4.64734
R48450 a_71281_n8397.n489 a_71281_n8397.n480 4.64734
R48451 a_71281_n8397.n474 a_71281_n8397.n470 4.64734
R48452 a_71281_n8397.n475 a_71281_n8397.n466 4.64734
R48453 a_71281_n8397.n741 a_71281_n8397.n732 4.64734
R48454 a_71281_n8397.n740 a_71281_n8397.n736 4.64734
R48455 a_71281_n8397.n755 a_71281_n8397.n746 4.64734
R48456 a_71281_n8397.n754 a_71281_n8397.n750 4.64734
R48457 a_71281_n8397.n769 a_71281_n8397.n760 4.64734
R48458 a_71281_n8397.n768 a_71281_n8397.n764 4.64734
R48459 a_71281_n8397.n783 a_71281_n8397.n774 4.64734
R48460 a_71281_n8397.n782 a_71281_n8397.n778 4.64734
R48461 a_71281_n8397.n868 a_71281_n8397.n864 4.64734
R48462 a_71281_n8397.n869 a_71281_n8397.n860 4.64734
R48463 a_71281_n8397.n854 a_71281_n8397.n850 4.64734
R48464 a_71281_n8397.n855 a_71281_n8397.n846 4.64734
R48465 a_71281_n8397.n837 a_71281_n8397.n833 4.64734
R48466 a_71281_n8397.n838 a_71281_n8397.n829 4.64734
R48467 a_71281_n8397.n823 a_71281_n8397.n819 4.64734
R48468 a_71281_n8397.n824 a_71281_n8397.n815 4.64734
R48469 a_71281_n8397.n642 a_71281_n8397.n641 4.01884
R48470 a_71281_n8397.n58 a_71281_n8397.n57 4.01884
R48471 a_71281_n8397.n234 a_71281_n8397.n233 4.01884
R48472 a_71281_n8397.n349 a_71281_n8397.n348 4.01884
R48473 a_71281_n8397.n525 a_71281_n8397.n524 4.01884
R48474 a_71281_n8397.n875 a_71281_n8397.n874 4.01884
R48475 a_71281_n8397.n673 a_71281_n8397.n672 4.00982
R48476 a_71281_n8397.n843 a_71281_n8397.n842 4.00982
R48477 a_71281_n8397.n89 a_71281_n8397.n88 4.00982
R48478 a_71281_n8397.n203 a_71281_n8397.n202 4.00982
R48479 a_71281_n8397.n380 a_71281_n8397.n379 4.00982
R48480 a_71281_n8397.n494 a_71281_n8397.n493 4.00982
R48481 a_71281_n8397.n584 a_71281_n8397.n292 3.61592
R48482 a_71281_n8397.n0 a_71281_n8397.n584 3.61491
R48483 a_71281_n8397.n714 a_71281_n8397.n713 2.25278
R48484 a_71281_n8397.n712 a_71281_n8397.n711 2.25278
R48485 a_71281_n8397.n728 a_71281_n8397.n727 2.25278
R48486 a_71281_n8397.n726 a_71281_n8397.n725 2.25278
R48487 a_71281_n8397.n809 a_71281_n8397.n808 2.25278
R48488 a_71281_n8397.n811 a_71281_n8397.n810 2.25278
R48489 a_71281_n8397.n795 a_71281_n8397.n794 2.25278
R48490 a_71281_n8397.n797 a_71281_n8397.n796 2.25278
R48491 a_71281_n8397.n594 a_71281_n8397.n593 2.25278
R48492 a_71281_n8397.n596 a_71281_n8397.n595 2.25278
R48493 a_71281_n8397.n608 a_71281_n8397.n607 2.25278
R48494 a_71281_n8397.n610 a_71281_n8397.n609 2.25278
R48495 a_71281_n8397.n622 a_71281_n8397.n621 2.25278
R48496 a_71281_n8397.n624 a_71281_n8397.n623 2.25278
R48497 a_71281_n8397.n636 a_71281_n8397.n635 2.25278
R48498 a_71281_n8397.n638 a_71281_n8397.n637 2.25278
R48499 a_71281_n8397.n653 a_71281_n8397.n652 2.25278
R48500 a_71281_n8397.n655 a_71281_n8397.n654 2.25278
R48501 a_71281_n8397.n667 a_71281_n8397.n666 2.25278
R48502 a_71281_n8397.n669 a_71281_n8397.n668 2.25278
R48503 a_71281_n8397.n684 a_71281_n8397.n683 2.25278
R48504 a_71281_n8397.n686 a_71281_n8397.n685 2.25278
R48505 a_71281_n8397.n698 a_71281_n8397.n697 2.25278
R48506 a_71281_n8397.n700 a_71281_n8397.n699 2.25278
R48507 a_71281_n8397.n130 a_71281_n8397.n129 2.25278
R48508 a_71281_n8397.n128 a_71281_n8397.n127 2.25278
R48509 a_71281_n8397.n144 a_71281_n8397.n143 2.25278
R48510 a_71281_n8397.n142 a_71281_n8397.n141 2.25278
R48511 a_71281_n8397.n169 a_71281_n8397.n168 2.25278
R48512 a_71281_n8397.n171 a_71281_n8397.n170 2.25278
R48513 a_71281_n8397.n155 a_71281_n8397.n154 2.25278
R48514 a_71281_n8397.n157 a_71281_n8397.n156 2.25278
R48515 a_71281_n8397.n10 a_71281_n8397.n9 2.25278
R48516 a_71281_n8397.n12 a_71281_n8397.n11 2.25278
R48517 a_71281_n8397.n24 a_71281_n8397.n23 2.25278
R48518 a_71281_n8397.n26 a_71281_n8397.n25 2.25278
R48519 a_71281_n8397.n38 a_71281_n8397.n37 2.25278
R48520 a_71281_n8397.n40 a_71281_n8397.n39 2.25278
R48521 a_71281_n8397.n52 a_71281_n8397.n51 2.25278
R48522 a_71281_n8397.n54 a_71281_n8397.n53 2.25278
R48523 a_71281_n8397.n69 a_71281_n8397.n68 2.25278
R48524 a_71281_n8397.n71 a_71281_n8397.n70 2.25278
R48525 a_71281_n8397.n83 a_71281_n8397.n82 2.25278
R48526 a_71281_n8397.n85 a_71281_n8397.n84 2.25278
R48527 a_71281_n8397.n100 a_71281_n8397.n99 2.25278
R48528 a_71281_n8397.n102 a_71281_n8397.n101 2.25278
R48529 a_71281_n8397.n114 a_71281_n8397.n113 2.25278
R48530 a_71281_n8397.n116 a_71281_n8397.n115 2.25278
R48531 a_71281_n8397.n289 a_71281_n8397.n288 2.25278
R48532 a_71281_n8397.n287 a_71281_n8397.n286 2.25278
R48533 a_71281_n8397.n275 a_71281_n8397.n274 2.25278
R48534 a_71281_n8397.n273 a_71281_n8397.n272 2.25278
R48535 a_71281_n8397.n261 a_71281_n8397.n260 2.25278
R48536 a_71281_n8397.n259 a_71281_n8397.n258 2.25278
R48537 a_71281_n8397.n247 a_71281_n8397.n246 2.25278
R48538 a_71281_n8397.n245 a_71281_n8397.n244 2.25278
R48539 a_71281_n8397.n230 a_71281_n8397.n229 2.25278
R48540 a_71281_n8397.n228 a_71281_n8397.n227 2.25278
R48541 a_71281_n8397.n216 a_71281_n8397.n215 2.25278
R48542 a_71281_n8397.n214 a_71281_n8397.n213 2.25278
R48543 a_71281_n8397.n199 a_71281_n8397.n198 2.25278
R48544 a_71281_n8397.n197 a_71281_n8397.n196 2.25278
R48545 a_71281_n8397.n185 a_71281_n8397.n184 2.25278
R48546 a_71281_n8397.n183 a_71281_n8397.n182 2.25278
R48547 a_71281_n8397.n421 a_71281_n8397.n420 2.25278
R48548 a_71281_n8397.n419 a_71281_n8397.n418 2.25278
R48549 a_71281_n8397.n435 a_71281_n8397.n434 2.25278
R48550 a_71281_n8397.n433 a_71281_n8397.n432 2.25278
R48551 a_71281_n8397.n460 a_71281_n8397.n459 2.25278
R48552 a_71281_n8397.n462 a_71281_n8397.n461 2.25278
R48553 a_71281_n8397.n446 a_71281_n8397.n445 2.25278
R48554 a_71281_n8397.n448 a_71281_n8397.n447 2.25278
R48555 a_71281_n8397.n301 a_71281_n8397.n300 2.25278
R48556 a_71281_n8397.n303 a_71281_n8397.n302 2.25278
R48557 a_71281_n8397.n315 a_71281_n8397.n314 2.25278
R48558 a_71281_n8397.n317 a_71281_n8397.n316 2.25278
R48559 a_71281_n8397.n329 a_71281_n8397.n328 2.25278
R48560 a_71281_n8397.n331 a_71281_n8397.n330 2.25278
R48561 a_71281_n8397.n343 a_71281_n8397.n342 2.25278
R48562 a_71281_n8397.n345 a_71281_n8397.n344 2.25278
R48563 a_71281_n8397.n360 a_71281_n8397.n359 2.25278
R48564 a_71281_n8397.n362 a_71281_n8397.n361 2.25278
R48565 a_71281_n8397.n374 a_71281_n8397.n373 2.25278
R48566 a_71281_n8397.n376 a_71281_n8397.n375 2.25278
R48567 a_71281_n8397.n391 a_71281_n8397.n390 2.25278
R48568 a_71281_n8397.n393 a_71281_n8397.n392 2.25278
R48569 a_71281_n8397.n405 a_71281_n8397.n404 2.25278
R48570 a_71281_n8397.n407 a_71281_n8397.n406 2.25278
R48571 a_71281_n8397.n580 a_71281_n8397.n579 2.25278
R48572 a_71281_n8397.n578 a_71281_n8397.n577 2.25278
R48573 a_71281_n8397.n566 a_71281_n8397.n565 2.25278
R48574 a_71281_n8397.n564 a_71281_n8397.n563 2.25278
R48575 a_71281_n8397.n552 a_71281_n8397.n551 2.25278
R48576 a_71281_n8397.n550 a_71281_n8397.n549 2.25278
R48577 a_71281_n8397.n538 a_71281_n8397.n537 2.25278
R48578 a_71281_n8397.n536 a_71281_n8397.n535 2.25278
R48579 a_71281_n8397.n521 a_71281_n8397.n520 2.25278
R48580 a_71281_n8397.n519 a_71281_n8397.n518 2.25278
R48581 a_71281_n8397.n507 a_71281_n8397.n506 2.25278
R48582 a_71281_n8397.n505 a_71281_n8397.n504 2.25278
R48583 a_71281_n8397.n490 a_71281_n8397.n489 2.25278
R48584 a_71281_n8397.n488 a_71281_n8397.n487 2.25278
R48585 a_71281_n8397.n476 a_71281_n8397.n475 2.25278
R48586 a_71281_n8397.n474 a_71281_n8397.n473 2.25278
R48587 a_71281_n8397.n740 a_71281_n8397.n739 2.25278
R48588 a_71281_n8397.n742 a_71281_n8397.n741 2.25278
R48589 a_71281_n8397.n754 a_71281_n8397.n753 2.25278
R48590 a_71281_n8397.n756 a_71281_n8397.n755 2.25278
R48591 a_71281_n8397.n768 a_71281_n8397.n767 2.25278
R48592 a_71281_n8397.n770 a_71281_n8397.n769 2.25278
R48593 a_71281_n8397.n782 a_71281_n8397.n781 2.25278
R48594 a_71281_n8397.n784 a_71281_n8397.n783 2.25278
R48595 a_71281_n8397.n870 a_71281_n8397.n869 2.25278
R48596 a_71281_n8397.n868 a_71281_n8397.n867 2.25278
R48597 a_71281_n8397.n856 a_71281_n8397.n855 2.25278
R48598 a_71281_n8397.n854 a_71281_n8397.n853 2.25278
R48599 a_71281_n8397.n839 a_71281_n8397.n838 2.25278
R48600 a_71281_n8397.n837 a_71281_n8397.n836 2.25278
R48601 a_71281_n8397.n825 a_71281_n8397.n824 2.25278
R48602 a_71281_n8397.n823 a_71281_n8397.n822 2.25278
R48603 a_71281_n8397.n1 a_71281_n8397.n0 0.0196917
R48604 a_71281_n8397.n14 a_71281_n8397.n2 1.6802
R48605 a_71281_n8397.n159 a_71281_n8397.n147 1.6802
R48606 a_71281_n8397.n305 a_71281_n8397.n293 1.6802
R48607 a_71281_n8397.n450 a_71281_n8397.n438 1.6802
R48608 a_71281_n8397.n598 a_71281_n8397.n586 1.6802
R48609 a_71281_n8397.n799 a_71281_n8397.n787 1.6802
R48610 a_71281_n8397.n180 a_71281_n8397.n174 1.5005
R48611 a_71281_n8397.n194 a_71281_n8397.n188 1.5005
R48612 a_71281_n8397.n211 a_71281_n8397.n205 1.5005
R48613 a_71281_n8397.n225 a_71281_n8397.n219 1.5005
R48614 a_71281_n8397.n235 a_71281_n8397.n234 1.5005
R48615 a_71281_n8397.n242 a_71281_n8397.n236 1.5005
R48616 a_71281_n8397.n256 a_71281_n8397.n250 1.5005
R48617 a_71281_n8397.n270 a_71281_n8397.n264 1.5005
R48618 a_71281_n8397.n284 a_71281_n8397.n278 1.5005
R48619 a_71281_n8397.n118 a_71281_n8397.n117 1.5005
R48620 a_71281_n8397.n104 a_71281_n8397.n103 1.5005
R48621 a_71281_n8397.n87 a_71281_n8397.n86 1.5005
R48622 a_71281_n8397.n73 a_71281_n8397.n72 1.5005
R48623 a_71281_n8397.n59 a_71281_n8397.n58 1.5005
R48624 a_71281_n8397.n56 a_71281_n8397.n55 1.5005
R48625 a_71281_n8397.n42 a_71281_n8397.n41 1.5005
R48626 a_71281_n8397.n28 a_71281_n8397.n27 1.5005
R48627 a_71281_n8397.n14 a_71281_n8397.n13 1.5005
R48628 a_71281_n8397.n204 a_71281_n8397.n203 1.5005
R48629 a_71281_n8397.n90 a_71281_n8397.n89 1.5005
R48630 a_71281_n8397.n159 a_71281_n8397.n158 1.5005
R48631 a_71281_n8397.n173 a_71281_n8397.n172 1.5005
R48632 a_71281_n8397.n167 a_71281_n8397.n160 1.5005
R48633 a_71281_n8397.n187 a_71281_n8397.n186 1.5005
R48634 a_71281_n8397.n201 a_71281_n8397.n200 1.5005
R48635 a_71281_n8397.n218 a_71281_n8397.n217 1.5005
R48636 a_71281_n8397.n232 a_71281_n8397.n231 1.5005
R48637 a_71281_n8397.n249 a_71281_n8397.n248 1.5005
R48638 a_71281_n8397.n263 a_71281_n8397.n262 1.5005
R48639 a_71281_n8397.n277 a_71281_n8397.n276 1.5005
R48640 a_71281_n8397.n291 a_71281_n8397.n290 1.5005
R48641 a_71281_n8397.n139 a_71281_n8397.n133 1.5005
R48642 a_71281_n8397.n146 a_71281_n8397.n145 1.5005
R48643 a_71281_n8397.n125 a_71281_n8397.n119 1.5005
R48644 a_71281_n8397.n132 a_71281_n8397.n131 1.5005
R48645 a_71281_n8397.n112 a_71281_n8397.n105 1.5005
R48646 a_71281_n8397.n98 a_71281_n8397.n91 1.5005
R48647 a_71281_n8397.n81 a_71281_n8397.n74 1.5005
R48648 a_71281_n8397.n67 a_71281_n8397.n60 1.5005
R48649 a_71281_n8397.n50 a_71281_n8397.n43 1.5005
R48650 a_71281_n8397.n36 a_71281_n8397.n29 1.5005
R48651 a_71281_n8397.n22 a_71281_n8397.n15 1.5005
R48652 a_71281_n8397.n471 a_71281_n8397.n465 1.5005
R48653 a_71281_n8397.n485 a_71281_n8397.n479 1.5005
R48654 a_71281_n8397.n502 a_71281_n8397.n496 1.5005
R48655 a_71281_n8397.n516 a_71281_n8397.n510 1.5005
R48656 a_71281_n8397.n526 a_71281_n8397.n525 1.5005
R48657 a_71281_n8397.n533 a_71281_n8397.n527 1.5005
R48658 a_71281_n8397.n547 a_71281_n8397.n541 1.5005
R48659 a_71281_n8397.n561 a_71281_n8397.n555 1.5005
R48660 a_71281_n8397.n575 a_71281_n8397.n569 1.5005
R48661 a_71281_n8397.n409 a_71281_n8397.n408 1.5005
R48662 a_71281_n8397.n395 a_71281_n8397.n394 1.5005
R48663 a_71281_n8397.n378 a_71281_n8397.n377 1.5005
R48664 a_71281_n8397.n364 a_71281_n8397.n363 1.5005
R48665 a_71281_n8397.n350 a_71281_n8397.n349 1.5005
R48666 a_71281_n8397.n347 a_71281_n8397.n346 1.5005
R48667 a_71281_n8397.n333 a_71281_n8397.n332 1.5005
R48668 a_71281_n8397.n319 a_71281_n8397.n318 1.5005
R48669 a_71281_n8397.n305 a_71281_n8397.n304 1.5005
R48670 a_71281_n8397.n495 a_71281_n8397.n494 1.5005
R48671 a_71281_n8397.n381 a_71281_n8397.n380 1.5005
R48672 a_71281_n8397.n450 a_71281_n8397.n449 1.5005
R48673 a_71281_n8397.n464 a_71281_n8397.n463 1.5005
R48674 a_71281_n8397.n458 a_71281_n8397.n451 1.5005
R48675 a_71281_n8397.n478 a_71281_n8397.n477 1.5005
R48676 a_71281_n8397.n492 a_71281_n8397.n491 1.5005
R48677 a_71281_n8397.n509 a_71281_n8397.n508 1.5005
R48678 a_71281_n8397.n523 a_71281_n8397.n522 1.5005
R48679 a_71281_n8397.n540 a_71281_n8397.n539 1.5005
R48680 a_71281_n8397.n554 a_71281_n8397.n553 1.5005
R48681 a_71281_n8397.n568 a_71281_n8397.n567 1.5005
R48682 a_71281_n8397.n582 a_71281_n8397.n581 1.5005
R48683 a_71281_n8397.n430 a_71281_n8397.n424 1.5005
R48684 a_71281_n8397.n437 a_71281_n8397.n436 1.5005
R48685 a_71281_n8397.n416 a_71281_n8397.n410 1.5005
R48686 a_71281_n8397.n423 a_71281_n8397.n422 1.5005
R48687 a_71281_n8397.n403 a_71281_n8397.n396 1.5005
R48688 a_71281_n8397.n389 a_71281_n8397.n382 1.5005
R48689 a_71281_n8397.n372 a_71281_n8397.n365 1.5005
R48690 a_71281_n8397.n358 a_71281_n8397.n351 1.5005
R48691 a_71281_n8397.n341 a_71281_n8397.n334 1.5005
R48692 a_71281_n8397.n327 a_71281_n8397.n320 1.5005
R48693 a_71281_n8397.n313 a_71281_n8397.n306 1.5005
R48694 a_71281_n8397.n820 a_71281_n8397.n814 1.5005
R48695 a_71281_n8397.n834 a_71281_n8397.n828 1.5005
R48696 a_71281_n8397.n851 a_71281_n8397.n845 1.5005
R48697 a_71281_n8397.n865 a_71281_n8397.n859 1.5005
R48698 a_71281_n8397.n786 a_71281_n8397.n785 1.5005
R48699 a_71281_n8397.n772 a_71281_n8397.n771 1.5005
R48700 a_71281_n8397.n758 a_71281_n8397.n757 1.5005
R48701 a_71281_n8397.n744 a_71281_n8397.n743 1.5005
R48702 a_71281_n8397.n702 a_71281_n8397.n701 1.5005
R48703 a_71281_n8397.n688 a_71281_n8397.n687 1.5005
R48704 a_71281_n8397.n671 a_71281_n8397.n670 1.5005
R48705 a_71281_n8397.n657 a_71281_n8397.n656 1.5005
R48706 a_71281_n8397.n643 a_71281_n8397.n642 1.5005
R48707 a_71281_n8397.n640 a_71281_n8397.n639 1.5005
R48708 a_71281_n8397.n626 a_71281_n8397.n625 1.5005
R48709 a_71281_n8397.n612 a_71281_n8397.n611 1.5005
R48710 a_71281_n8397.n598 a_71281_n8397.n597 1.5005
R48711 a_71281_n8397.n844 a_71281_n8397.n843 1.5005
R48712 a_71281_n8397.n674 a_71281_n8397.n673 1.5005
R48713 a_71281_n8397.n799 a_71281_n8397.n798 1.5005
R48714 a_71281_n8397.n813 a_71281_n8397.n812 1.5005
R48715 a_71281_n8397.n807 a_71281_n8397.n800 1.5005
R48716 a_71281_n8397.n827 a_71281_n8397.n826 1.5005
R48717 a_71281_n8397.n841 a_71281_n8397.n840 1.5005
R48718 a_71281_n8397.n858 a_71281_n8397.n857 1.5005
R48719 a_71281_n8397.n872 a_71281_n8397.n871 1.5005
R48720 a_71281_n8397.n780 a_71281_n8397.n773 1.5005
R48721 a_71281_n8397.n766 a_71281_n8397.n759 1.5005
R48722 a_71281_n8397.n752 a_71281_n8397.n745 1.5005
R48723 a_71281_n8397.n738 a_71281_n8397.n731 1.5005
R48724 a_71281_n8397.n723 a_71281_n8397.n717 1.5005
R48725 a_71281_n8397.n730 a_71281_n8397.n729 1.5005
R48726 a_71281_n8397.n709 a_71281_n8397.n703 1.5005
R48727 a_71281_n8397.n716 a_71281_n8397.n715 1.5005
R48728 a_71281_n8397.n696 a_71281_n8397.n689 1.5005
R48729 a_71281_n8397.n682 a_71281_n8397.n675 1.5005
R48730 a_71281_n8397.n665 a_71281_n8397.n658 1.5005
R48731 a_71281_n8397.n651 a_71281_n8397.n644 1.5005
R48732 a_71281_n8397.n634 a_71281_n8397.n627 1.5005
R48733 a_71281_n8397.n620 a_71281_n8397.n613 1.5005
R48734 a_71281_n8397.n606 a_71281_n8397.n599 1.5005
R48735 a_71281_n8397.n874 a_71281_n8397.n873 1.5005
R48736 a_71281_n8397.n672 a_71281_n8397.t31 1.4705
R48737 a_71281_n8397.n672 a_71281_n8397.t27 1.4705
R48738 a_71281_n8397.n842 a_71281_n8397.t21 1.4705
R48739 a_71281_n8397.n842 a_71281_n8397.t51 1.4705
R48740 a_71281_n8397.n641 a_71281_n8397.t55 1.4705
R48741 a_71281_n8397.n641 a_71281_n8397.t33 1.4705
R48742 a_71281_n8397.n88 a_71281_n8397.t45 1.4705
R48743 a_71281_n8397.n88 a_71281_n8397.t19 1.4705
R48744 a_71281_n8397.n202 a_71281_n8397.t63 1.4705
R48745 a_71281_n8397.n202 a_71281_n8397.t11 1.4705
R48746 a_71281_n8397.n57 a_71281_n8397.t41 1.4705
R48747 a_71281_n8397.n57 a_71281_n8397.t9 1.4705
R48748 a_71281_n8397.n233 a_71281_n8397.t29 1.4705
R48749 a_71281_n8397.n233 a_71281_n8397.t37 1.4705
R48750 a_71281_n8397.n379 a_71281_n8397.t57 1.4705
R48751 a_71281_n8397.n379 a_71281_n8397.t25 1.4705
R48752 a_71281_n8397.n493 a_71281_n8397.t35 1.4705
R48753 a_71281_n8397.n493 a_71281_n8397.t47 1.4705
R48754 a_71281_n8397.n348 a_71281_n8397.t53 1.4705
R48755 a_71281_n8397.n348 a_71281_n8397.t23 1.4705
R48756 a_71281_n8397.n524 a_71281_n8397.t67 1.4705
R48757 a_71281_n8397.n524 a_71281_n8397.t69 1.4705
R48758 a_71281_n8397.t71 a_71281_n8397.n875 1.4705
R48759 a_71281_n8397.n875 a_71281_n8397.t39 1.4705
R48760 a_71281_n8397.n584 a_71281_n8397.n583 0.7505
R48761 a_71281_n8397.n714 a_71281_n8397.n705 0.567403
R48762 a_71281_n8397.n711 a_71281_n8397.n710 0.567403
R48763 a_71281_n8397.n728 a_71281_n8397.n719 0.567403
R48764 a_71281_n8397.n725 a_71281_n8397.n724 0.567403
R48765 a_71281_n8397.n808 a_71281_n8397.n806 0.567403
R48766 a_71281_n8397.n811 a_71281_n8397.n802 0.567403
R48767 a_71281_n8397.n794 a_71281_n8397.n793 0.567403
R48768 a_71281_n8397.n797 a_71281_n8397.n789 0.567403
R48769 a_71281_n8397.n593 a_71281_n8397.n592 0.567403
R48770 a_71281_n8397.n596 a_71281_n8397.n588 0.567403
R48771 a_71281_n8397.n607 a_71281_n8397.n605 0.567403
R48772 a_71281_n8397.n610 a_71281_n8397.n601 0.567403
R48773 a_71281_n8397.n621 a_71281_n8397.n619 0.567403
R48774 a_71281_n8397.n624 a_71281_n8397.n615 0.567403
R48775 a_71281_n8397.n635 a_71281_n8397.n633 0.567403
R48776 a_71281_n8397.n638 a_71281_n8397.n629 0.567403
R48777 a_71281_n8397.n652 a_71281_n8397.n650 0.567403
R48778 a_71281_n8397.n655 a_71281_n8397.n646 0.567403
R48779 a_71281_n8397.n666 a_71281_n8397.n664 0.567403
R48780 a_71281_n8397.n669 a_71281_n8397.n660 0.567403
R48781 a_71281_n8397.n683 a_71281_n8397.n681 0.567403
R48782 a_71281_n8397.n686 a_71281_n8397.n677 0.567403
R48783 a_71281_n8397.n697 a_71281_n8397.n695 0.567403
R48784 a_71281_n8397.n700 a_71281_n8397.n691 0.567403
R48785 a_71281_n8397.n130 a_71281_n8397.n121 0.567403
R48786 a_71281_n8397.n127 a_71281_n8397.n126 0.567403
R48787 a_71281_n8397.n144 a_71281_n8397.n135 0.567403
R48788 a_71281_n8397.n141 a_71281_n8397.n140 0.567403
R48789 a_71281_n8397.n168 a_71281_n8397.n166 0.567403
R48790 a_71281_n8397.n171 a_71281_n8397.n162 0.567403
R48791 a_71281_n8397.n154 a_71281_n8397.n153 0.567403
R48792 a_71281_n8397.n157 a_71281_n8397.n149 0.567403
R48793 a_71281_n8397.n9 a_71281_n8397.n8 0.567403
R48794 a_71281_n8397.n12 a_71281_n8397.n4 0.567403
R48795 a_71281_n8397.n23 a_71281_n8397.n21 0.567403
R48796 a_71281_n8397.n26 a_71281_n8397.n17 0.567403
R48797 a_71281_n8397.n37 a_71281_n8397.n35 0.567403
R48798 a_71281_n8397.n40 a_71281_n8397.n31 0.567403
R48799 a_71281_n8397.n51 a_71281_n8397.n49 0.567403
R48800 a_71281_n8397.n54 a_71281_n8397.n45 0.567403
R48801 a_71281_n8397.n68 a_71281_n8397.n66 0.567403
R48802 a_71281_n8397.n71 a_71281_n8397.n62 0.567403
R48803 a_71281_n8397.n82 a_71281_n8397.n80 0.567403
R48804 a_71281_n8397.n85 a_71281_n8397.n76 0.567403
R48805 a_71281_n8397.n99 a_71281_n8397.n97 0.567403
R48806 a_71281_n8397.n102 a_71281_n8397.n93 0.567403
R48807 a_71281_n8397.n113 a_71281_n8397.n111 0.567403
R48808 a_71281_n8397.n116 a_71281_n8397.n107 0.567403
R48809 a_71281_n8397.n289 a_71281_n8397.n280 0.567403
R48810 a_71281_n8397.n286 a_71281_n8397.n285 0.567403
R48811 a_71281_n8397.n275 a_71281_n8397.n266 0.567403
R48812 a_71281_n8397.n272 a_71281_n8397.n271 0.567403
R48813 a_71281_n8397.n261 a_71281_n8397.n252 0.567403
R48814 a_71281_n8397.n258 a_71281_n8397.n257 0.567403
R48815 a_71281_n8397.n247 a_71281_n8397.n238 0.567403
R48816 a_71281_n8397.n244 a_71281_n8397.n243 0.567403
R48817 a_71281_n8397.n230 a_71281_n8397.n221 0.567403
R48818 a_71281_n8397.n227 a_71281_n8397.n226 0.567403
R48819 a_71281_n8397.n216 a_71281_n8397.n207 0.567403
R48820 a_71281_n8397.n213 a_71281_n8397.n212 0.567403
R48821 a_71281_n8397.n199 a_71281_n8397.n190 0.567403
R48822 a_71281_n8397.n196 a_71281_n8397.n195 0.567403
R48823 a_71281_n8397.n185 a_71281_n8397.n176 0.567403
R48824 a_71281_n8397.n182 a_71281_n8397.n181 0.567403
R48825 a_71281_n8397.n421 a_71281_n8397.n412 0.567403
R48826 a_71281_n8397.n418 a_71281_n8397.n417 0.567403
R48827 a_71281_n8397.n435 a_71281_n8397.n426 0.567403
R48828 a_71281_n8397.n432 a_71281_n8397.n431 0.567403
R48829 a_71281_n8397.n459 a_71281_n8397.n457 0.567403
R48830 a_71281_n8397.n462 a_71281_n8397.n453 0.567403
R48831 a_71281_n8397.n445 a_71281_n8397.n444 0.567403
R48832 a_71281_n8397.n448 a_71281_n8397.n440 0.567403
R48833 a_71281_n8397.n300 a_71281_n8397.n299 0.567403
R48834 a_71281_n8397.n303 a_71281_n8397.n295 0.567403
R48835 a_71281_n8397.n314 a_71281_n8397.n312 0.567403
R48836 a_71281_n8397.n317 a_71281_n8397.n308 0.567403
R48837 a_71281_n8397.n328 a_71281_n8397.n326 0.567403
R48838 a_71281_n8397.n331 a_71281_n8397.n322 0.567403
R48839 a_71281_n8397.n342 a_71281_n8397.n340 0.567403
R48840 a_71281_n8397.n345 a_71281_n8397.n336 0.567403
R48841 a_71281_n8397.n359 a_71281_n8397.n357 0.567403
R48842 a_71281_n8397.n362 a_71281_n8397.n353 0.567403
R48843 a_71281_n8397.n373 a_71281_n8397.n371 0.567403
R48844 a_71281_n8397.n376 a_71281_n8397.n367 0.567403
R48845 a_71281_n8397.n390 a_71281_n8397.n388 0.567403
R48846 a_71281_n8397.n393 a_71281_n8397.n384 0.567403
R48847 a_71281_n8397.n404 a_71281_n8397.n402 0.567403
R48848 a_71281_n8397.n407 a_71281_n8397.n398 0.567403
R48849 a_71281_n8397.n580 a_71281_n8397.n571 0.567403
R48850 a_71281_n8397.n577 a_71281_n8397.n576 0.567403
R48851 a_71281_n8397.n566 a_71281_n8397.n557 0.567403
R48852 a_71281_n8397.n563 a_71281_n8397.n562 0.567403
R48853 a_71281_n8397.n552 a_71281_n8397.n543 0.567403
R48854 a_71281_n8397.n549 a_71281_n8397.n548 0.567403
R48855 a_71281_n8397.n538 a_71281_n8397.n529 0.567403
R48856 a_71281_n8397.n535 a_71281_n8397.n534 0.567403
R48857 a_71281_n8397.n521 a_71281_n8397.n512 0.567403
R48858 a_71281_n8397.n518 a_71281_n8397.n517 0.567403
R48859 a_71281_n8397.n507 a_71281_n8397.n498 0.567403
R48860 a_71281_n8397.n504 a_71281_n8397.n503 0.567403
R48861 a_71281_n8397.n490 a_71281_n8397.n481 0.567403
R48862 a_71281_n8397.n487 a_71281_n8397.n486 0.567403
R48863 a_71281_n8397.n476 a_71281_n8397.n467 0.567403
R48864 a_71281_n8397.n473 a_71281_n8397.n472 0.567403
R48865 a_71281_n8397.n739 a_71281_n8397.n737 0.567403
R48866 a_71281_n8397.n742 a_71281_n8397.n733 0.567403
R48867 a_71281_n8397.n753 a_71281_n8397.n751 0.567403
R48868 a_71281_n8397.n756 a_71281_n8397.n747 0.567403
R48869 a_71281_n8397.n767 a_71281_n8397.n765 0.567403
R48870 a_71281_n8397.n770 a_71281_n8397.n761 0.567403
R48871 a_71281_n8397.n781 a_71281_n8397.n779 0.567403
R48872 a_71281_n8397.n784 a_71281_n8397.n775 0.567403
R48873 a_71281_n8397.n870 a_71281_n8397.n861 0.567403
R48874 a_71281_n8397.n867 a_71281_n8397.n866 0.567403
R48875 a_71281_n8397.n856 a_71281_n8397.n847 0.567403
R48876 a_71281_n8397.n853 a_71281_n8397.n852 0.567403
R48877 a_71281_n8397.n839 a_71281_n8397.n830 0.567403
R48878 a_71281_n8397.n836 a_71281_n8397.n835 0.567403
R48879 a_71281_n8397.n825 a_71281_n8397.n816 0.567403
R48880 a_71281_n8397.n822 a_71281_n8397.n821 0.567403
R48881 a_71281_n8397.n706 a_71281_n8397.n704 0.496742
R48882 a_71281_n8397.n708 a_71281_n8397.n707 0.496742
R48883 a_71281_n8397.n720 a_71281_n8397.n718 0.496742
R48884 a_71281_n8397.n722 a_71281_n8397.n721 0.496742
R48885 a_71281_n8397.n805 a_71281_n8397.n804 0.496742
R48886 a_71281_n8397.n803 a_71281_n8397.n801 0.496742
R48887 a_71281_n8397.n792 a_71281_n8397.n791 0.496742
R48888 a_71281_n8397.n790 a_71281_n8397.n788 0.496742
R48889 a_71281_n8397.n591 a_71281_n8397.n590 0.496742
R48890 a_71281_n8397.n589 a_71281_n8397.n587 0.496742
R48891 a_71281_n8397.n604 a_71281_n8397.n603 0.496742
R48892 a_71281_n8397.n602 a_71281_n8397.n600 0.496742
R48893 a_71281_n8397.n618 a_71281_n8397.n617 0.496742
R48894 a_71281_n8397.n616 a_71281_n8397.n614 0.496742
R48895 a_71281_n8397.n632 a_71281_n8397.n631 0.496742
R48896 a_71281_n8397.n630 a_71281_n8397.n628 0.496742
R48897 a_71281_n8397.n649 a_71281_n8397.n648 0.496742
R48898 a_71281_n8397.n647 a_71281_n8397.n645 0.496742
R48899 a_71281_n8397.n663 a_71281_n8397.n662 0.496742
R48900 a_71281_n8397.n661 a_71281_n8397.n659 0.496742
R48901 a_71281_n8397.n680 a_71281_n8397.n679 0.496742
R48902 a_71281_n8397.n678 a_71281_n8397.n676 0.496742
R48903 a_71281_n8397.n694 a_71281_n8397.n693 0.496742
R48904 a_71281_n8397.n692 a_71281_n8397.n690 0.496742
R48905 a_71281_n8397.n122 a_71281_n8397.n120 0.496742
R48906 a_71281_n8397.n124 a_71281_n8397.n123 0.496742
R48907 a_71281_n8397.n136 a_71281_n8397.n134 0.496742
R48908 a_71281_n8397.n138 a_71281_n8397.n137 0.496742
R48909 a_71281_n8397.n165 a_71281_n8397.n164 0.496742
R48910 a_71281_n8397.n163 a_71281_n8397.n161 0.496742
R48911 a_71281_n8397.n152 a_71281_n8397.n151 0.496742
R48912 a_71281_n8397.n150 a_71281_n8397.n148 0.496742
R48913 a_71281_n8397.n7 a_71281_n8397.n6 0.496742
R48914 a_71281_n8397.n5 a_71281_n8397.n3 0.496742
R48915 a_71281_n8397.n20 a_71281_n8397.n19 0.496742
R48916 a_71281_n8397.n18 a_71281_n8397.n16 0.496742
R48917 a_71281_n8397.n34 a_71281_n8397.n33 0.496742
R48918 a_71281_n8397.n32 a_71281_n8397.n30 0.496742
R48919 a_71281_n8397.n48 a_71281_n8397.n47 0.496742
R48920 a_71281_n8397.n46 a_71281_n8397.n44 0.496742
R48921 a_71281_n8397.n65 a_71281_n8397.n64 0.496742
R48922 a_71281_n8397.n63 a_71281_n8397.n61 0.496742
R48923 a_71281_n8397.n79 a_71281_n8397.n78 0.496742
R48924 a_71281_n8397.n77 a_71281_n8397.n75 0.496742
R48925 a_71281_n8397.n96 a_71281_n8397.n95 0.496742
R48926 a_71281_n8397.n94 a_71281_n8397.n92 0.496742
R48927 a_71281_n8397.n110 a_71281_n8397.n109 0.496742
R48928 a_71281_n8397.n108 a_71281_n8397.n106 0.496742
R48929 a_71281_n8397.n281 a_71281_n8397.n279 0.496742
R48930 a_71281_n8397.n283 a_71281_n8397.n282 0.496742
R48931 a_71281_n8397.n267 a_71281_n8397.n265 0.496742
R48932 a_71281_n8397.n269 a_71281_n8397.n268 0.496742
R48933 a_71281_n8397.n253 a_71281_n8397.n251 0.496742
R48934 a_71281_n8397.n255 a_71281_n8397.n254 0.496742
R48935 a_71281_n8397.n239 a_71281_n8397.n237 0.496742
R48936 a_71281_n8397.n241 a_71281_n8397.n240 0.496742
R48937 a_71281_n8397.n222 a_71281_n8397.n220 0.496742
R48938 a_71281_n8397.n224 a_71281_n8397.n223 0.496742
R48939 a_71281_n8397.n208 a_71281_n8397.n206 0.496742
R48940 a_71281_n8397.n210 a_71281_n8397.n209 0.496742
R48941 a_71281_n8397.n191 a_71281_n8397.n189 0.496742
R48942 a_71281_n8397.n193 a_71281_n8397.n192 0.496742
R48943 a_71281_n8397.n177 a_71281_n8397.n175 0.496742
R48944 a_71281_n8397.n179 a_71281_n8397.n178 0.496742
R48945 a_71281_n8397.n413 a_71281_n8397.n411 0.496742
R48946 a_71281_n8397.n415 a_71281_n8397.n414 0.496742
R48947 a_71281_n8397.n427 a_71281_n8397.n425 0.496742
R48948 a_71281_n8397.n429 a_71281_n8397.n428 0.496742
R48949 a_71281_n8397.n456 a_71281_n8397.n455 0.496742
R48950 a_71281_n8397.n454 a_71281_n8397.n452 0.496742
R48951 a_71281_n8397.n443 a_71281_n8397.n442 0.496742
R48952 a_71281_n8397.n441 a_71281_n8397.n439 0.496742
R48953 a_71281_n8397.n298 a_71281_n8397.n297 0.496742
R48954 a_71281_n8397.n296 a_71281_n8397.n294 0.496742
R48955 a_71281_n8397.n311 a_71281_n8397.n310 0.496742
R48956 a_71281_n8397.n309 a_71281_n8397.n307 0.496742
R48957 a_71281_n8397.n325 a_71281_n8397.n324 0.496742
R48958 a_71281_n8397.n323 a_71281_n8397.n321 0.496742
R48959 a_71281_n8397.n339 a_71281_n8397.n338 0.496742
R48960 a_71281_n8397.n337 a_71281_n8397.n335 0.496742
R48961 a_71281_n8397.n356 a_71281_n8397.n355 0.496742
R48962 a_71281_n8397.n354 a_71281_n8397.n352 0.496742
R48963 a_71281_n8397.n370 a_71281_n8397.n369 0.496742
R48964 a_71281_n8397.n368 a_71281_n8397.n366 0.496742
R48965 a_71281_n8397.n387 a_71281_n8397.n386 0.496742
R48966 a_71281_n8397.n385 a_71281_n8397.n383 0.496742
R48967 a_71281_n8397.n401 a_71281_n8397.n400 0.496742
R48968 a_71281_n8397.n399 a_71281_n8397.n397 0.496742
R48969 a_71281_n8397.n572 a_71281_n8397.n570 0.496742
R48970 a_71281_n8397.n574 a_71281_n8397.n573 0.496742
R48971 a_71281_n8397.n558 a_71281_n8397.n556 0.496742
R48972 a_71281_n8397.n560 a_71281_n8397.n559 0.496742
R48973 a_71281_n8397.n544 a_71281_n8397.n542 0.496742
R48974 a_71281_n8397.n546 a_71281_n8397.n545 0.496742
R48975 a_71281_n8397.n530 a_71281_n8397.n528 0.496742
R48976 a_71281_n8397.n532 a_71281_n8397.n531 0.496742
R48977 a_71281_n8397.n513 a_71281_n8397.n511 0.496742
R48978 a_71281_n8397.n515 a_71281_n8397.n514 0.496742
R48979 a_71281_n8397.n499 a_71281_n8397.n497 0.496742
R48980 a_71281_n8397.n501 a_71281_n8397.n500 0.496742
R48981 a_71281_n8397.n482 a_71281_n8397.n480 0.496742
R48982 a_71281_n8397.n484 a_71281_n8397.n483 0.496742
R48983 a_71281_n8397.n468 a_71281_n8397.n466 0.496742
R48984 a_71281_n8397.n470 a_71281_n8397.n469 0.496742
R48985 a_71281_n8397.n736 a_71281_n8397.n735 0.496742
R48986 a_71281_n8397.n734 a_71281_n8397.n732 0.496742
R48987 a_71281_n8397.n750 a_71281_n8397.n749 0.496742
R48988 a_71281_n8397.n748 a_71281_n8397.n746 0.496742
R48989 a_71281_n8397.n764 a_71281_n8397.n763 0.496742
R48990 a_71281_n8397.n762 a_71281_n8397.n760 0.496742
R48991 a_71281_n8397.n778 a_71281_n8397.n777 0.496742
R48992 a_71281_n8397.n776 a_71281_n8397.n774 0.496742
R48993 a_71281_n8397.n862 a_71281_n8397.n860 0.496742
R48994 a_71281_n8397.n864 a_71281_n8397.n863 0.496742
R48995 a_71281_n8397.n848 a_71281_n8397.n846 0.496742
R48996 a_71281_n8397.n850 a_71281_n8397.n849 0.496742
R48997 a_71281_n8397.n831 a_71281_n8397.n829 0.496742
R48998 a_71281_n8397.n833 a_71281_n8397.n832 0.496742
R48999 a_71281_n8397.n817 a_71281_n8397.n815 0.496742
R49000 a_71281_n8397.n819 a_71281_n8397.n818 0.496742
R49001 a_71281_n8397.n292 a_71281_n8397.n291 0.445939
R49002 a_71281_n8397.n583 a_71281_n8397.n582 0.445939
R49003 a_71281_n8397.n292 a_71281_n8397.n146 0.443507
R49004 a_71281_n8397.n583 a_71281_n8397.n437 0.443507
R49005 a_71281_n8397.n0 a_71281_n8397.n730 0.427392
R49006 a_71281_n8397.n56 a_71281_n8397.n43 0.180804
R49007 a_71281_n8397.n132 a_71281_n8397.n119 0.180804
R49008 a_71281_n8397.n249 a_71281_n8397.n236 0.180804
R49009 a_71281_n8397.n173 a_71281_n8397.n160 0.180804
R49010 a_71281_n8397.n347 a_71281_n8397.n334 0.180804
R49011 a_71281_n8397.n423 a_71281_n8397.n410 0.180804
R49012 a_71281_n8397.n540 a_71281_n8397.n527 0.180804
R49013 a_71281_n8397.n464 a_71281_n8397.n451 0.180804
R49014 a_71281_n8397.n640 a_71281_n8397.n627 0.180804
R49015 a_71281_n8397.n716 a_71281_n8397.n703 0.180804
R49016 a_71281_n8397.n786 a_71281_n8397.n773 0.180804
R49017 a_71281_n8397.n813 a_71281_n8397.n800 0.180804
R49018 a_71281_n8397.n42 a_71281_n8397.n29 0.180196
R49019 a_71281_n8397.n73 a_71281_n8397.n60 0.180196
R49020 a_71281_n8397.n87 a_71281_n8397.n74 0.180196
R49021 a_71281_n8397.n118 a_71281_n8397.n105 0.180196
R49022 a_71281_n8397.n146 a_71281_n8397.n133 0.180196
R49023 a_71281_n8397.n291 a_71281_n8397.n278 0.180196
R49024 a_71281_n8397.n263 a_71281_n8397.n250 0.180196
R49025 a_71281_n8397.n232 a_71281_n8397.n219 0.180196
R49026 a_71281_n8397.n218 a_71281_n8397.n205 0.180196
R49027 a_71281_n8397.n187 a_71281_n8397.n174 0.180196
R49028 a_71281_n8397.n333 a_71281_n8397.n320 0.180196
R49029 a_71281_n8397.n364 a_71281_n8397.n351 0.180196
R49030 a_71281_n8397.n378 a_71281_n8397.n365 0.180196
R49031 a_71281_n8397.n409 a_71281_n8397.n396 0.180196
R49032 a_71281_n8397.n437 a_71281_n8397.n424 0.180196
R49033 a_71281_n8397.n582 a_71281_n8397.n569 0.180196
R49034 a_71281_n8397.n554 a_71281_n8397.n541 0.180196
R49035 a_71281_n8397.n523 a_71281_n8397.n510 0.180196
R49036 a_71281_n8397.n509 a_71281_n8397.n496 0.180196
R49037 a_71281_n8397.n478 a_71281_n8397.n465 0.180196
R49038 a_71281_n8397.n626 a_71281_n8397.n613 0.180196
R49039 a_71281_n8397.n657 a_71281_n8397.n644 0.180196
R49040 a_71281_n8397.n671 a_71281_n8397.n658 0.180196
R49041 a_71281_n8397.n702 a_71281_n8397.n689 0.180196
R49042 a_71281_n8397.n730 a_71281_n8397.n717 0.180196
R49043 a_71281_n8397.n744 a_71281_n8397.n731 0.180196
R49044 a_71281_n8397.n772 a_71281_n8397.n759 0.180196
R49045 a_71281_n8397.n872 a_71281_n8397.n859 0.180196
R49046 a_71281_n8397.n858 a_71281_n8397.n845 0.180196
R49047 a_71281_n8397.n827 a_71281_n8397.n814 0.180196
R49048 a_71281_n8397.n28 a_71281_n8397.n15 0.179892
R49049 a_71281_n8397.n104 a_71281_n8397.n91 0.179892
R49050 a_71281_n8397.n277 a_71281_n8397.n264 0.179892
R49051 a_71281_n8397.n201 a_71281_n8397.n188 0.179892
R49052 a_71281_n8397.n319 a_71281_n8397.n306 0.179892
R49053 a_71281_n8397.n395 a_71281_n8397.n382 0.179892
R49054 a_71281_n8397.n568 a_71281_n8397.n555 0.179892
R49055 a_71281_n8397.n492 a_71281_n8397.n479 0.179892
R49056 a_71281_n8397.n612 a_71281_n8397.n599 0.179892
R49057 a_71281_n8397.n688 a_71281_n8397.n675 0.179892
R49058 a_71281_n8397.n758 a_71281_n8397.n745 0.179892
R49059 a_71281_n8397.n841 a_71281_n8397.n828 0.179892
R49060 a_71281_n8397.n715 a_71281_n8397.n704 0.136625
R49061 a_71281_n8397.n709 a_71281_n8397.n708 0.136625
R49062 a_71281_n8397.n729 a_71281_n8397.n718 0.136625
R49063 a_71281_n8397.n723 a_71281_n8397.n722 0.136625
R49064 a_71281_n8397.n807 a_71281_n8397.n805 0.136625
R49065 a_71281_n8397.n812 a_71281_n8397.n801 0.136625
R49066 a_71281_n8397.n792 a_71281_n8397.n787 0.136625
R49067 a_71281_n8397.n798 a_71281_n8397.n788 0.136625
R49068 a_71281_n8397.n591 a_71281_n8397.n586 0.136625
R49069 a_71281_n8397.n597 a_71281_n8397.n587 0.136625
R49070 a_71281_n8397.n606 a_71281_n8397.n604 0.136625
R49071 a_71281_n8397.n611 a_71281_n8397.n600 0.136625
R49072 a_71281_n8397.n620 a_71281_n8397.n618 0.136625
R49073 a_71281_n8397.n625 a_71281_n8397.n614 0.136625
R49074 a_71281_n8397.n634 a_71281_n8397.n632 0.136625
R49075 a_71281_n8397.n639 a_71281_n8397.n628 0.136625
R49076 a_71281_n8397.n651 a_71281_n8397.n649 0.136625
R49077 a_71281_n8397.n656 a_71281_n8397.n645 0.136625
R49078 a_71281_n8397.n665 a_71281_n8397.n663 0.136625
R49079 a_71281_n8397.n670 a_71281_n8397.n659 0.136625
R49080 a_71281_n8397.n682 a_71281_n8397.n680 0.136625
R49081 a_71281_n8397.n687 a_71281_n8397.n676 0.136625
R49082 a_71281_n8397.n696 a_71281_n8397.n694 0.136625
R49083 a_71281_n8397.n701 a_71281_n8397.n690 0.136625
R49084 a_71281_n8397.n131 a_71281_n8397.n120 0.136625
R49085 a_71281_n8397.n125 a_71281_n8397.n124 0.136625
R49086 a_71281_n8397.n145 a_71281_n8397.n134 0.136625
R49087 a_71281_n8397.n139 a_71281_n8397.n138 0.136625
R49088 a_71281_n8397.n167 a_71281_n8397.n165 0.136625
R49089 a_71281_n8397.n172 a_71281_n8397.n161 0.136625
R49090 a_71281_n8397.n152 a_71281_n8397.n147 0.136625
R49091 a_71281_n8397.n158 a_71281_n8397.n148 0.136625
R49092 a_71281_n8397.n7 a_71281_n8397.n2 0.136625
R49093 a_71281_n8397.n13 a_71281_n8397.n3 0.136625
R49094 a_71281_n8397.n22 a_71281_n8397.n20 0.136625
R49095 a_71281_n8397.n27 a_71281_n8397.n16 0.136625
R49096 a_71281_n8397.n36 a_71281_n8397.n34 0.136625
R49097 a_71281_n8397.n41 a_71281_n8397.n30 0.136625
R49098 a_71281_n8397.n50 a_71281_n8397.n48 0.136625
R49099 a_71281_n8397.n55 a_71281_n8397.n44 0.136625
R49100 a_71281_n8397.n67 a_71281_n8397.n65 0.136625
R49101 a_71281_n8397.n72 a_71281_n8397.n61 0.136625
R49102 a_71281_n8397.n81 a_71281_n8397.n79 0.136625
R49103 a_71281_n8397.n86 a_71281_n8397.n75 0.136625
R49104 a_71281_n8397.n98 a_71281_n8397.n96 0.136625
R49105 a_71281_n8397.n103 a_71281_n8397.n92 0.136625
R49106 a_71281_n8397.n112 a_71281_n8397.n110 0.136625
R49107 a_71281_n8397.n117 a_71281_n8397.n106 0.136625
R49108 a_71281_n8397.n290 a_71281_n8397.n279 0.136625
R49109 a_71281_n8397.n284 a_71281_n8397.n283 0.136625
R49110 a_71281_n8397.n276 a_71281_n8397.n265 0.136625
R49111 a_71281_n8397.n270 a_71281_n8397.n269 0.136625
R49112 a_71281_n8397.n262 a_71281_n8397.n251 0.136625
R49113 a_71281_n8397.n256 a_71281_n8397.n255 0.136625
R49114 a_71281_n8397.n248 a_71281_n8397.n237 0.136625
R49115 a_71281_n8397.n242 a_71281_n8397.n241 0.136625
R49116 a_71281_n8397.n231 a_71281_n8397.n220 0.136625
R49117 a_71281_n8397.n225 a_71281_n8397.n224 0.136625
R49118 a_71281_n8397.n217 a_71281_n8397.n206 0.136625
R49119 a_71281_n8397.n211 a_71281_n8397.n210 0.136625
R49120 a_71281_n8397.n200 a_71281_n8397.n189 0.136625
R49121 a_71281_n8397.n194 a_71281_n8397.n193 0.136625
R49122 a_71281_n8397.n186 a_71281_n8397.n175 0.136625
R49123 a_71281_n8397.n180 a_71281_n8397.n179 0.136625
R49124 a_71281_n8397.n422 a_71281_n8397.n411 0.136625
R49125 a_71281_n8397.n416 a_71281_n8397.n415 0.136625
R49126 a_71281_n8397.n436 a_71281_n8397.n425 0.136625
R49127 a_71281_n8397.n430 a_71281_n8397.n429 0.136625
R49128 a_71281_n8397.n458 a_71281_n8397.n456 0.136625
R49129 a_71281_n8397.n463 a_71281_n8397.n452 0.136625
R49130 a_71281_n8397.n443 a_71281_n8397.n438 0.136625
R49131 a_71281_n8397.n449 a_71281_n8397.n439 0.136625
R49132 a_71281_n8397.n298 a_71281_n8397.n293 0.136625
R49133 a_71281_n8397.n304 a_71281_n8397.n294 0.136625
R49134 a_71281_n8397.n313 a_71281_n8397.n311 0.136625
R49135 a_71281_n8397.n318 a_71281_n8397.n307 0.136625
R49136 a_71281_n8397.n327 a_71281_n8397.n325 0.136625
R49137 a_71281_n8397.n332 a_71281_n8397.n321 0.136625
R49138 a_71281_n8397.n341 a_71281_n8397.n339 0.136625
R49139 a_71281_n8397.n346 a_71281_n8397.n335 0.136625
R49140 a_71281_n8397.n358 a_71281_n8397.n356 0.136625
R49141 a_71281_n8397.n363 a_71281_n8397.n352 0.136625
R49142 a_71281_n8397.n372 a_71281_n8397.n370 0.136625
R49143 a_71281_n8397.n377 a_71281_n8397.n366 0.136625
R49144 a_71281_n8397.n389 a_71281_n8397.n387 0.136625
R49145 a_71281_n8397.n394 a_71281_n8397.n383 0.136625
R49146 a_71281_n8397.n403 a_71281_n8397.n401 0.136625
R49147 a_71281_n8397.n408 a_71281_n8397.n397 0.136625
R49148 a_71281_n8397.n581 a_71281_n8397.n570 0.136625
R49149 a_71281_n8397.n575 a_71281_n8397.n574 0.136625
R49150 a_71281_n8397.n567 a_71281_n8397.n556 0.136625
R49151 a_71281_n8397.n561 a_71281_n8397.n560 0.136625
R49152 a_71281_n8397.n553 a_71281_n8397.n542 0.136625
R49153 a_71281_n8397.n547 a_71281_n8397.n546 0.136625
R49154 a_71281_n8397.n539 a_71281_n8397.n528 0.136625
R49155 a_71281_n8397.n533 a_71281_n8397.n532 0.136625
R49156 a_71281_n8397.n522 a_71281_n8397.n511 0.136625
R49157 a_71281_n8397.n516 a_71281_n8397.n515 0.136625
R49158 a_71281_n8397.n508 a_71281_n8397.n497 0.136625
R49159 a_71281_n8397.n502 a_71281_n8397.n501 0.136625
R49160 a_71281_n8397.n491 a_71281_n8397.n480 0.136625
R49161 a_71281_n8397.n485 a_71281_n8397.n484 0.136625
R49162 a_71281_n8397.n477 a_71281_n8397.n466 0.136625
R49163 a_71281_n8397.n471 a_71281_n8397.n470 0.136625
R49164 a_71281_n8397.n738 a_71281_n8397.n736 0.136625
R49165 a_71281_n8397.n743 a_71281_n8397.n732 0.136625
R49166 a_71281_n8397.n752 a_71281_n8397.n750 0.136625
R49167 a_71281_n8397.n757 a_71281_n8397.n746 0.136625
R49168 a_71281_n8397.n766 a_71281_n8397.n764 0.136625
R49169 a_71281_n8397.n771 a_71281_n8397.n760 0.136625
R49170 a_71281_n8397.n780 a_71281_n8397.n778 0.136625
R49171 a_71281_n8397.n785 a_71281_n8397.n774 0.136625
R49172 a_71281_n8397.n871 a_71281_n8397.n860 0.136625
R49173 a_71281_n8397.n865 a_71281_n8397.n864 0.136625
R49174 a_71281_n8397.n857 a_71281_n8397.n846 0.136625
R49175 a_71281_n8397.n851 a_71281_n8397.n850 0.136625
R49176 a_71281_n8397.n840 a_71281_n8397.n829 0.136625
R49177 a_71281_n8397.n834 a_71281_n8397.n833 0.136625
R49178 a_71281_n8397.n826 a_71281_n8397.n815 0.136625
R49179 a_71281_n8397.n820 a_71281_n8397.n819 0.136625
R49180 a_71281_n8397.n15 a_71281_n8397.n14 0.095973
R49181 a_71281_n8397.n29 a_71281_n8397.n28 0.095973
R49182 a_71281_n8397.n43 a_71281_n8397.n42 0.095973
R49183 a_71281_n8397.n74 a_71281_n8397.n73 0.095973
R49184 a_71281_n8397.n105 a_71281_n8397.n104 0.095973
R49185 a_71281_n8397.n119 a_71281_n8397.n118 0.095973
R49186 a_71281_n8397.n133 a_71281_n8397.n132 0.095973
R49187 a_71281_n8397.n278 a_71281_n8397.n277 0.095973
R49188 a_71281_n8397.n264 a_71281_n8397.n263 0.095973
R49189 a_71281_n8397.n250 a_71281_n8397.n249 0.095973
R49190 a_71281_n8397.n219 a_71281_n8397.n218 0.095973
R49191 a_71281_n8397.n188 a_71281_n8397.n187 0.095973
R49192 a_71281_n8397.n174 a_71281_n8397.n173 0.095973
R49193 a_71281_n8397.n160 a_71281_n8397.n159 0.095973
R49194 a_71281_n8397.n306 a_71281_n8397.n305 0.095973
R49195 a_71281_n8397.n320 a_71281_n8397.n319 0.095973
R49196 a_71281_n8397.n334 a_71281_n8397.n333 0.095973
R49197 a_71281_n8397.n365 a_71281_n8397.n364 0.095973
R49198 a_71281_n8397.n396 a_71281_n8397.n395 0.095973
R49199 a_71281_n8397.n410 a_71281_n8397.n409 0.095973
R49200 a_71281_n8397.n424 a_71281_n8397.n423 0.095973
R49201 a_71281_n8397.n569 a_71281_n8397.n568 0.095973
R49202 a_71281_n8397.n555 a_71281_n8397.n554 0.095973
R49203 a_71281_n8397.n541 a_71281_n8397.n540 0.095973
R49204 a_71281_n8397.n510 a_71281_n8397.n509 0.095973
R49205 a_71281_n8397.n479 a_71281_n8397.n478 0.095973
R49206 a_71281_n8397.n465 a_71281_n8397.n464 0.095973
R49207 a_71281_n8397.n451 a_71281_n8397.n450 0.095973
R49208 a_71281_n8397.n599 a_71281_n8397.n598 0.095973
R49209 a_71281_n8397.n613 a_71281_n8397.n612 0.095973
R49210 a_71281_n8397.n627 a_71281_n8397.n626 0.095973
R49211 a_71281_n8397.n658 a_71281_n8397.n657 0.095973
R49212 a_71281_n8397.n689 a_71281_n8397.n688 0.095973
R49213 a_71281_n8397.n703 a_71281_n8397.n702 0.095973
R49214 a_71281_n8397.n717 a_71281_n8397.n716 0.095973
R49215 a_71281_n8397.n745 a_71281_n8397.n744 0.095973
R49216 a_71281_n8397.n759 a_71281_n8397.n758 0.095973
R49217 a_71281_n8397.n773 a_71281_n8397.n772 0.095973
R49218 a_71281_n8397.n859 a_71281_n8397.n858 0.095973
R49219 a_71281_n8397.n828 a_71281_n8397.n827 0.095973
R49220 a_71281_n8397.n814 a_71281_n8397.n813 0.095973
R49221 a_71281_n8397.n800 a_71281_n8397.n799 0.095973
R49222 a_71281_n8397.n715 a_71281_n8397.n714 0.0719743
R49223 a_71281_n8397.n711 a_71281_n8397.n709 0.0719743
R49224 a_71281_n8397.n729 a_71281_n8397.n728 0.0719743
R49225 a_71281_n8397.n725 a_71281_n8397.n723 0.0719743
R49226 a_71281_n8397.n808 a_71281_n8397.n807 0.0719743
R49227 a_71281_n8397.n812 a_71281_n8397.n811 0.0719743
R49228 a_71281_n8397.n794 a_71281_n8397.n787 0.0719743
R49229 a_71281_n8397.n798 a_71281_n8397.n797 0.0719743
R49230 a_71281_n8397.n593 a_71281_n8397.n586 0.0719743
R49231 a_71281_n8397.n597 a_71281_n8397.n596 0.0719743
R49232 a_71281_n8397.n607 a_71281_n8397.n606 0.0719743
R49233 a_71281_n8397.n611 a_71281_n8397.n610 0.0719743
R49234 a_71281_n8397.n621 a_71281_n8397.n620 0.0719743
R49235 a_71281_n8397.n625 a_71281_n8397.n624 0.0719743
R49236 a_71281_n8397.n635 a_71281_n8397.n634 0.0719743
R49237 a_71281_n8397.n639 a_71281_n8397.n638 0.0719743
R49238 a_71281_n8397.n652 a_71281_n8397.n651 0.0719743
R49239 a_71281_n8397.n656 a_71281_n8397.n655 0.0719743
R49240 a_71281_n8397.n666 a_71281_n8397.n665 0.0719743
R49241 a_71281_n8397.n670 a_71281_n8397.n669 0.0719743
R49242 a_71281_n8397.n683 a_71281_n8397.n682 0.0719743
R49243 a_71281_n8397.n687 a_71281_n8397.n686 0.0719743
R49244 a_71281_n8397.n697 a_71281_n8397.n696 0.0719743
R49245 a_71281_n8397.n701 a_71281_n8397.n700 0.0719743
R49246 a_71281_n8397.n131 a_71281_n8397.n130 0.0719743
R49247 a_71281_n8397.n127 a_71281_n8397.n125 0.0719743
R49248 a_71281_n8397.n145 a_71281_n8397.n144 0.0719743
R49249 a_71281_n8397.n141 a_71281_n8397.n139 0.0719743
R49250 a_71281_n8397.n168 a_71281_n8397.n167 0.0719743
R49251 a_71281_n8397.n172 a_71281_n8397.n171 0.0719743
R49252 a_71281_n8397.n154 a_71281_n8397.n147 0.0719743
R49253 a_71281_n8397.n158 a_71281_n8397.n157 0.0719743
R49254 a_71281_n8397.n9 a_71281_n8397.n2 0.0719743
R49255 a_71281_n8397.n13 a_71281_n8397.n12 0.0719743
R49256 a_71281_n8397.n23 a_71281_n8397.n22 0.0719743
R49257 a_71281_n8397.n27 a_71281_n8397.n26 0.0719743
R49258 a_71281_n8397.n37 a_71281_n8397.n36 0.0719743
R49259 a_71281_n8397.n41 a_71281_n8397.n40 0.0719743
R49260 a_71281_n8397.n51 a_71281_n8397.n50 0.0719743
R49261 a_71281_n8397.n55 a_71281_n8397.n54 0.0719743
R49262 a_71281_n8397.n68 a_71281_n8397.n67 0.0719743
R49263 a_71281_n8397.n72 a_71281_n8397.n71 0.0719743
R49264 a_71281_n8397.n82 a_71281_n8397.n81 0.0719743
R49265 a_71281_n8397.n86 a_71281_n8397.n85 0.0719743
R49266 a_71281_n8397.n99 a_71281_n8397.n98 0.0719743
R49267 a_71281_n8397.n103 a_71281_n8397.n102 0.0719743
R49268 a_71281_n8397.n113 a_71281_n8397.n112 0.0719743
R49269 a_71281_n8397.n117 a_71281_n8397.n116 0.0719743
R49270 a_71281_n8397.n290 a_71281_n8397.n289 0.0719743
R49271 a_71281_n8397.n286 a_71281_n8397.n284 0.0719743
R49272 a_71281_n8397.n276 a_71281_n8397.n275 0.0719743
R49273 a_71281_n8397.n272 a_71281_n8397.n270 0.0719743
R49274 a_71281_n8397.n262 a_71281_n8397.n261 0.0719743
R49275 a_71281_n8397.n258 a_71281_n8397.n256 0.0719743
R49276 a_71281_n8397.n248 a_71281_n8397.n247 0.0719743
R49277 a_71281_n8397.n244 a_71281_n8397.n242 0.0719743
R49278 a_71281_n8397.n231 a_71281_n8397.n230 0.0719743
R49279 a_71281_n8397.n227 a_71281_n8397.n225 0.0719743
R49280 a_71281_n8397.n217 a_71281_n8397.n216 0.0719743
R49281 a_71281_n8397.n213 a_71281_n8397.n211 0.0719743
R49282 a_71281_n8397.n200 a_71281_n8397.n199 0.0719743
R49283 a_71281_n8397.n196 a_71281_n8397.n194 0.0719743
R49284 a_71281_n8397.n186 a_71281_n8397.n185 0.0719743
R49285 a_71281_n8397.n182 a_71281_n8397.n180 0.0719743
R49286 a_71281_n8397.n422 a_71281_n8397.n421 0.0719743
R49287 a_71281_n8397.n418 a_71281_n8397.n416 0.0719743
R49288 a_71281_n8397.n436 a_71281_n8397.n435 0.0719743
R49289 a_71281_n8397.n432 a_71281_n8397.n430 0.0719743
R49290 a_71281_n8397.n459 a_71281_n8397.n458 0.0719743
R49291 a_71281_n8397.n463 a_71281_n8397.n462 0.0719743
R49292 a_71281_n8397.n445 a_71281_n8397.n438 0.0719743
R49293 a_71281_n8397.n449 a_71281_n8397.n448 0.0719743
R49294 a_71281_n8397.n300 a_71281_n8397.n293 0.0719743
R49295 a_71281_n8397.n304 a_71281_n8397.n303 0.0719743
R49296 a_71281_n8397.n314 a_71281_n8397.n313 0.0719743
R49297 a_71281_n8397.n318 a_71281_n8397.n317 0.0719743
R49298 a_71281_n8397.n328 a_71281_n8397.n327 0.0719743
R49299 a_71281_n8397.n332 a_71281_n8397.n331 0.0719743
R49300 a_71281_n8397.n342 a_71281_n8397.n341 0.0719743
R49301 a_71281_n8397.n346 a_71281_n8397.n345 0.0719743
R49302 a_71281_n8397.n359 a_71281_n8397.n358 0.0719743
R49303 a_71281_n8397.n363 a_71281_n8397.n362 0.0719743
R49304 a_71281_n8397.n373 a_71281_n8397.n372 0.0719743
R49305 a_71281_n8397.n377 a_71281_n8397.n376 0.0719743
R49306 a_71281_n8397.n390 a_71281_n8397.n389 0.0719743
R49307 a_71281_n8397.n394 a_71281_n8397.n393 0.0719743
R49308 a_71281_n8397.n404 a_71281_n8397.n403 0.0719743
R49309 a_71281_n8397.n408 a_71281_n8397.n407 0.0719743
R49310 a_71281_n8397.n581 a_71281_n8397.n580 0.0719743
R49311 a_71281_n8397.n577 a_71281_n8397.n575 0.0719743
R49312 a_71281_n8397.n567 a_71281_n8397.n566 0.0719743
R49313 a_71281_n8397.n563 a_71281_n8397.n561 0.0719743
R49314 a_71281_n8397.n553 a_71281_n8397.n552 0.0719743
R49315 a_71281_n8397.n549 a_71281_n8397.n547 0.0719743
R49316 a_71281_n8397.n539 a_71281_n8397.n538 0.0719743
R49317 a_71281_n8397.n535 a_71281_n8397.n533 0.0719743
R49318 a_71281_n8397.n522 a_71281_n8397.n521 0.0719743
R49319 a_71281_n8397.n518 a_71281_n8397.n516 0.0719743
R49320 a_71281_n8397.n508 a_71281_n8397.n507 0.0719743
R49321 a_71281_n8397.n504 a_71281_n8397.n502 0.0719743
R49322 a_71281_n8397.n491 a_71281_n8397.n490 0.0719743
R49323 a_71281_n8397.n487 a_71281_n8397.n485 0.0719743
R49324 a_71281_n8397.n477 a_71281_n8397.n476 0.0719743
R49325 a_71281_n8397.n473 a_71281_n8397.n471 0.0719743
R49326 a_71281_n8397.n739 a_71281_n8397.n738 0.0719743
R49327 a_71281_n8397.n743 a_71281_n8397.n742 0.0719743
R49328 a_71281_n8397.n753 a_71281_n8397.n752 0.0719743
R49329 a_71281_n8397.n757 a_71281_n8397.n756 0.0719743
R49330 a_71281_n8397.n767 a_71281_n8397.n766 0.0719743
R49331 a_71281_n8397.n771 a_71281_n8397.n770 0.0719743
R49332 a_71281_n8397.n781 a_71281_n8397.n780 0.0719743
R49333 a_71281_n8397.n785 a_71281_n8397.n784 0.0719743
R49334 a_71281_n8397.n871 a_71281_n8397.n870 0.0719743
R49335 a_71281_n8397.n867 a_71281_n8397.n865 0.0719743
R49336 a_71281_n8397.n857 a_71281_n8397.n856 0.0719743
R49337 a_71281_n8397.n853 a_71281_n8397.n851 0.0719743
R49338 a_71281_n8397.n840 a_71281_n8397.n839 0.0719743
R49339 a_71281_n8397.n836 a_71281_n8397.n834 0.0719743
R49340 a_71281_n8397.n826 a_71281_n8397.n825 0.0719743
R49341 a_71281_n8397.n822 a_71281_n8397.n820 0.0719743
R49342 a_71281_n8397.n60 a_71281_n8397.n59 0.0485405
R49343 a_71281_n8397.n235 a_71281_n8397.n232 0.0485405
R49344 a_71281_n8397.n351 a_71281_n8397.n350 0.0485405
R49345 a_71281_n8397.n526 a_71281_n8397.n523 0.0485405
R49346 a_71281_n8397.n644 a_71281_n8397.n643 0.0485405
R49347 a_71281_n8397.n873 a_71281_n8397.n872 0.0485405
R49348 a_71281_n8397.n90 a_71281_n8397.n87 0.0482365
R49349 a_71281_n8397.n91 a_71281_n8397.n90 0.0482365
R49350 a_71281_n8397.n205 a_71281_n8397.n204 0.0482365
R49351 a_71281_n8397.n204 a_71281_n8397.n201 0.0482365
R49352 a_71281_n8397.n381 a_71281_n8397.n378 0.0482365
R49353 a_71281_n8397.n382 a_71281_n8397.n381 0.0482365
R49354 a_71281_n8397.n496 a_71281_n8397.n495 0.0482365
R49355 a_71281_n8397.n495 a_71281_n8397.n492 0.0482365
R49356 a_71281_n8397.n674 a_71281_n8397.n671 0.0482365
R49357 a_71281_n8397.n675 a_71281_n8397.n674 0.0482365
R49358 a_71281_n8397.n845 a_71281_n8397.n844 0.0482365
R49359 a_71281_n8397.n844 a_71281_n8397.n841 0.0482365
R49360 a_71281_n8397.n59 a_71281_n8397.n56 0.0479324
R49361 a_71281_n8397.n236 a_71281_n8397.n235 0.0479324
R49362 a_71281_n8397.n350 a_71281_n8397.n347 0.0479324
R49363 a_71281_n8397.n527 a_71281_n8397.n526 0.0479324
R49364 a_71281_n8397.n643 a_71281_n8397.n640 0.0479324
R49365 a_71281_n8397.n873 a_71281_n8397.n786 0.0479324
R49366 a_71281_n8397.n731 a_71281_n8397.n1 0.443549
R49367 a_35922_19591.n237 a_35922_19591.n230 10.6966
R49368 a_35922_19591.n234 a_35922_19591.t104 8.75329
R49369 a_35922_19591.n236 a_35922_19591.t86 8.75329
R49370 a_35922_19591.n233 a_35922_19591.t99 8.75329
R49371 a_35922_19591.n235 a_35922_19591.t51 8.75329
R49372 a_35922_19591.n143 a_35922_19591.t38 8.38704
R49373 a_35922_19591.n132 a_35922_19591.t64 8.38704
R49374 a_35922_19591.n100 a_35922_19591.t150 8.46135
R49375 a_35922_19591.n101 a_35922_19591.t155 8.46135
R49376 a_35922_19591.n0 a_35922_19591.t14 8.39293
R49377 a_35922_19591.n109 a_35922_19591.t168 8.39293
R49378 a_35922_19591.n59 a_35922_19591.t132 8.26625
R49379 a_35922_19591.n61 a_35922_19591.t102 8.26625
R49380 a_35922_19591.n62 a_35922_19591.t71 8.26625
R49381 a_35922_19591.n234 a_35922_19591.t61 8.12045
R49382 a_35922_19591.n236 a_35922_19591.t29 8.12045
R49383 a_35922_19591.n233 a_35922_19591.t58 8.12045
R49384 a_35922_19591.n232 a_35922_19591.t124 8.12045
R49385 a_35922_19591.n235 a_35922_19591.t149 8.12045
R49386 a_35922_19591.n90 a_35922_19591.t80 8.10567
R49387 a_35922_19591.n72 a_35922_19591.t173 8.10567
R49388 a_35922_19591.n72 a_35922_19591.t122 8.10567
R49389 a_35922_19591.n72 a_35922_19591.t84 8.10567
R49390 a_35922_19591.n72 a_35922_19591.t183 8.10567
R49391 a_35922_19591.n31 a_35922_19591.t191 8.10567
R49392 a_35922_19591.n31 a_35922_19591.t13 8.10567
R49393 a_35922_19591.n31 a_35922_19591.t138 8.10567
R49394 a_35922_19591.n31 a_35922_19591.t52 8.10567
R49395 a_35922_19591.n34 a_35922_19591.t15 8.10567
R49396 a_35922_19591.n34 a_35922_19591.t174 8.10567
R49397 a_35922_19591.n34 a_35922_19591.t125 8.10567
R49398 a_35922_19591.n34 a_35922_19591.t26 8.10567
R49399 a_35922_19591.n70 a_35922_19591.t59 8.10567
R49400 a_35922_19591.n70 a_35922_19591.t128 8.10567
R49401 a_35922_19591.n70 a_35922_19591.t76 8.10567
R49402 a_35922_19591.n68 a_35922_19591.t74 8.10567
R49403 a_35922_19591.n68 a_35922_19591.t143 8.10567
R49404 a_35922_19591.n68 a_35922_19591.t131 8.10567
R49405 a_35922_19591.n90 a_35922_19591.t45 8.10567
R49406 a_35922_19591.n90 a_35922_19591.t147 8.10567
R49407 a_35922_19591.n90 a_35922_19591.t44 8.10567
R49408 a_35922_19591.n99 a_35922_19591.t77 8.10567
R49409 a_35922_19591.n86 a_35922_19591.t163 8.10567
R49410 a_35922_19591.n86 a_35922_19591.t116 8.10567
R49411 a_35922_19591.n86 a_35922_19591.t82 8.10567
R49412 a_35922_19591.n86 a_35922_19591.t170 8.10567
R49413 a_35922_19591.n48 a_35922_19591.t178 8.10567
R49414 a_35922_19591.n48 a_35922_19591.t187 8.10567
R49415 a_35922_19591.n48 a_35922_19591.t134 8.10567
R49416 a_35922_19591.n48 a_35922_19591.t37 8.10567
R49417 a_35922_19591.n50 a_35922_19591.t190 8.10567
R49418 a_35922_19591.n50 a_35922_19591.t165 8.10567
R49419 a_35922_19591.n50 a_35922_19591.t117 8.10567
R49420 a_35922_19591.n50 a_35922_19591.t12 8.10567
R49421 a_35922_19591.n82 a_35922_19591.t182 8.10567
R49422 a_35922_19591.n82 a_35922_19591.t87 8.10567
R49423 a_35922_19591.n82 a_35922_19591.t33 8.10567
R49424 a_35922_19591.n80 a_35922_19591.t25 8.10567
R49425 a_35922_19591.n80 a_35922_19591.t98 8.10567
R49426 a_35922_19591.n80 a_35922_19591.t89 8.10567
R49427 a_35922_19591.n99 a_35922_19591.t31 8.10567
R49428 a_35922_19591.n99 a_35922_19591.t144 8.10567
R49429 a_35922_19591.n99 a_35922_19591.t30 8.10567
R49430 a_35922_19591.n91 a_35922_19591.t70 8.10567
R49431 a_35922_19591.n74 a_35922_19591.t152 8.10567
R49432 a_35922_19591.n74 a_35922_19591.t101 8.10567
R49433 a_35922_19591.n74 a_35922_19591.t75 8.10567
R49434 a_35922_19591.n74 a_35922_19591.t158 8.10567
R49435 a_35922_19591.n39 a_35922_19591.t160 8.10567
R49436 a_35922_19591.n39 a_35922_19591.t167 8.10567
R49437 a_35922_19591.n39 a_35922_19591.t119 8.10567
R49438 a_35922_19591.n39 a_35922_19591.t19 8.10567
R49439 a_35922_19591.n43 a_35922_19591.t169 8.10567
R49440 a_35922_19591.n43 a_35922_19591.t154 8.10567
R49441 a_35922_19591.n43 a_35922_19591.t103 8.10567
R49442 a_35922_19591.n43 a_35922_19591.t181 8.10567
R49443 a_35922_19591.n66 a_35922_19591.t34 8.10567
R49444 a_35922_19591.n66 a_35922_19591.t105 8.10567
R49445 a_35922_19591.n66 a_35922_19591.t62 8.10567
R49446 a_35922_19591.n64 a_35922_19591.t57 8.10567
R49447 a_35922_19591.n64 a_35922_19591.t123 8.10567
R49448 a_35922_19591.n64 a_35922_19591.t108 8.10567
R49449 a_35922_19591.n91 a_35922_19591.t9 8.10567
R49450 a_35922_19591.n91 a_35922_19591.t137 8.10567
R49451 a_35922_19591.n91 a_35922_19591.t8 8.10567
R49452 a_35922_19591.n94 a_35922_19591.t81 8.10567
R49453 a_35922_19591.n84 a_35922_19591.t176 8.10567
R49454 a_35922_19591.n84 a_35922_19591.t127 8.10567
R49455 a_35922_19591.n84 a_35922_19591.t85 8.10567
R49456 a_35922_19591.n84 a_35922_19591.t185 8.10567
R49457 a_35922_19591.n54 a_35922_19591.t193 8.10567
R49458 a_35922_19591.n54 a_35922_19591.t17 8.10567
R49459 a_35922_19591.n54 a_35922_19591.t141 8.10567
R49460 a_35922_19591.n54 a_35922_19591.t55 8.10567
R49461 a_35922_19591.n56 a_35922_19591.t21 8.10567
R49462 a_35922_19591.n56 a_35922_19591.t180 8.10567
R49463 a_35922_19591.n56 a_35922_19591.t130 8.10567
R49464 a_35922_19591.n56 a_35922_19591.t28 8.10567
R49465 a_35922_19591.n78 a_35922_19591.t11 8.10567
R49466 a_35922_19591.n78 a_35922_19591.t92 8.10567
R49467 a_35922_19591.n78 a_35922_19591.t50 8.10567
R49468 a_35922_19591.n76 a_35922_19591.t42 8.10567
R49469 a_35922_19591.n76 a_35922_19591.t113 8.10567
R49470 a_35922_19591.n76 a_35922_19591.t93 8.10567
R49471 a_35922_19591.n94 a_35922_19591.t49 8.10567
R49472 a_35922_19591.n94 a_35922_19591.t148 8.10567
R49473 a_35922_19591.n94 a_35922_19591.t47 8.10567
R49474 a_35922_19591.n0 a_35922_19591.t32 8.10567
R49475 a_35922_19591.n0 a_35922_19591.t43 8.10567
R49476 a_35922_19591.n0 a_35922_19591.t146 8.10567
R49477 a_35922_19591.n0 a_35922_19591.t69 8.10567
R49478 a_35922_19591.n0 a_35922_19591.t36 8.10567
R49479 a_35922_19591.n0 a_35922_19591.t109 8.10567
R49480 a_35922_19591.n0 a_35922_19591.t66 8.10567
R49481 a_35922_19591.n0 a_35922_19591.t94 8.10567
R49482 a_35922_19591.n0 a_35922_19591.t24 8.10567
R49483 a_35922_19591.n105 a_35922_19591.t88 8.10567
R49484 a_35922_19591.n103 a_35922_19591.t65 8.10567
R49485 a_35922_19591.n131 a_35922_19591.t157 8.10567
R49486 a_35922_19591.n2 a_35922_19591.t60 8.10567
R49487 a_35922_19591.n228 a_35922_19591.t129 8.10567
R49488 a_35922_19591.n227 a_35922_19591.t111 8.10567
R49489 a_35922_19591.n3 a_35922_19591.t46 8.10567
R49490 a_35922_19591.n3 a_35922_19591.t16 8.10567
R49491 a_35922_19591.n3 a_35922_19591.t140 8.10567
R49492 a_35922_19591.n3 a_35922_19591.t54 8.10567
R49493 a_35922_19591.n12 a_35922_19591.t156 8.10567
R49494 a_35922_19591.n12 a_35922_19591.t162 8.10567
R49495 a_35922_19591.n12 a_35922_19591.t115 8.10567
R49496 a_35922_19591.n12 a_35922_19591.t6 8.10567
R49497 a_35922_19591.n27 a_35922_19591.t23 8.10567
R49498 a_35922_19591.n162 a_35922_19591.t97 8.10567
R49499 a_35922_19591.n161 a_35922_19591.t56 8.10567
R49500 a_35922_19591.n28 a_35922_19591.t95 8.10567
R49501 a_35922_19591.n29 a_35922_19591.t73 8.10567
R49502 a_35922_19591.n29 a_35922_19591.t153 8.10567
R49503 a_35922_19591.n4 a_35922_19591.t67 8.10567
R49504 a_35922_19591.n4 a_35922_19591.t189 8.10567
R49505 a_35922_19591.n4 a_35922_19591.t135 8.10567
R49506 a_35922_19591.n25 a_35922_19591.t53 8.10567
R49507 a_35922_19591.n160 a_35922_19591.t118 8.10567
R49508 a_35922_19591.n159 a_35922_19591.t100 8.10567
R49509 a_35922_19591.n17 a_35922_19591.t164 8.10567
R49510 a_35922_19591.n17 a_35922_19591.t151 8.10567
R49511 a_35922_19591.n16 a_35922_19591.t96 8.10567
R49512 a_35922_19591.n16 a_35922_19591.t171 8.10567
R49513 a_35922_19591.n112 a_35922_19591.t184 8.10567
R49514 a_35922_19591.n111 a_35922_19591.t7 8.10567
R49515 a_35922_19591.n110 a_35922_19591.t136 8.10567
R49516 a_35922_19591.n194 a_35922_19591.t48 8.10567
R49517 a_35922_19591.n177 a_35922_19591.t192 8.10567
R49518 a_35922_19591.n178 a_35922_19591.t90 8.10567
R49519 a_35922_19591.n179 a_35922_19591.t41 8.10567
R49520 a_35922_19591.n108 a_35922_19591.t120 8.10567
R49521 a_35922_19591.n107 a_35922_19591.t83 8.10567
R49522 a_35922_19591.n106 a_35922_19591.t179 8.10567
R49523 a_35922_19591.n126 a_35922_19591.t79 8.10567
R49524 a_35922_19591.n124 a_35922_19591.t39 8.10567
R49525 a_35922_19591.n142 a_35922_19591.t145 8.10567
R49526 a_35922_19591.n153 a_35922_19591.t35 8.10567
R49527 a_35922_19591.n152 a_35922_19591.t106 8.10567
R49528 a_35922_19591.n151 a_35922_19591.t91 8.10567
R49529 a_35922_19591.n120 a_35922_19591.t10 8.10567
R49530 a_35922_19591.n119 a_35922_19591.t172 8.10567
R49531 a_35922_19591.n118 a_35922_19591.t121 8.10567
R49532 a_35922_19591.n115 a_35922_19591.t22 8.10567
R49533 a_35922_19591.n10 a_35922_19591.t166 8.10567
R49534 a_35922_19591.n10 a_35922_19591.t175 8.10567
R49535 a_35922_19591.n10 a_35922_19591.t126 8.10567
R49536 a_35922_19591.n10 a_35922_19591.t27 8.10567
R49537 a_35922_19591.n212 a_35922_19591.t40 8.10567
R49538 a_35922_19591.n213 a_35922_19591.t112 8.10567
R49539 a_35922_19591.n9 a_35922_19591.t68 8.10567
R49540 a_35922_19591.n22 a_35922_19591.t107 8.10567
R49541 a_35922_19591.n23 a_35922_19591.t78 8.10567
R49542 a_35922_19591.n23 a_35922_19591.t161 8.10567
R49543 a_35922_19591.n8 a_35922_19591.t72 8.10567
R49544 a_35922_19591.n8 a_35922_19591.t20 8.10567
R49545 a_35922_19591.n8 a_35922_19591.t142 8.10567
R49546 a_35922_19591.n19 a_35922_19591.t63 8.10567
R49547 a_35922_19591.n210 a_35922_19591.t133 8.10567
R49548 a_35922_19591.n209 a_35922_19591.t114 8.10567
R49549 a_35922_19591.n14 a_35922_19591.t177 8.10567
R49550 a_35922_19591.n14 a_35922_19591.t159 8.10567
R49551 a_35922_19591.n20 a_35922_19591.t110 8.10567
R49552 a_35922_19591.n20 a_35922_19591.t186 8.10567
R49553 a_35922_19591.n231 a_35922_19591.t0 6.69607
R49554 a_35922_19591.n240 a_35922_19591.t2 6.0467
R49555 a_35922_19591.n231 a_35922_19591.t1 5.54843
R49556 a_35922_19591.n238 a_35922_19591.t3 5.44096
R49557 a_35922_19591.n238 a_35922_19591.t4 5.41626
R49558 a_35922_19591.n239 a_35922_19591.n237 4.8989
R49559 a_35922_19591.t5 a_35922_19591.n240 4.79524
R49560 a_35922_19591.n1 a_35922_19591.n3 0.426349
R49561 a_35922_19591.n121 a_35922_19591.n120 2.25163
R49562 a_35922_19591.n18 a_35922_19591.n17 0.607617
R49563 a_35922_19591.n15 a_35922_19591.n14 0.607617
R49564 a_35922_19591.n86 a_35922_19591.n87 0.020246
R49565 a_35922_19591.n85 a_35922_19591.n84 0.020246
R49566 a_35922_19591.n48 a_35922_19591.n47 0.150783
R49567 a_35922_19591.n50 a_35922_19591.n46 0.150803
R49568 a_35922_19591.n99 a_35922_19591.n98 0.0676355
R49569 a_35922_19591.n54 a_35922_19591.n53 0.150803
R49570 a_35922_19591.n58 a_35922_19591.n56 0.150806
R49571 a_35922_19591.n95 a_35922_19591.n94 0.0676255
R49572 a_35922_19591.n34 a_35922_19591.n35 0.153625
R49573 a_35922_19591.n31 a_35922_19591.n32 0.153625
R49574 a_35922_19591.n73 a_35922_19591.n72 0.020088
R49575 a_35922_19591.n51 a_35922_19591.n50 0.246907
R49576 a_35922_19591.n48 a_35922_19591.n49 0.246877
R49577 a_35922_19591.n44 a_35922_19591.n43 0.153625
R49578 a_35922_19591.n40 a_35922_19591.n39 0.153625
R49579 a_35922_19591.n74 a_35922_19591.n75 0.020088
R49580 a_35922_19591.n91 a_35922_19591.n92 0.0201939
R49581 a_35922_19591.n43 a_35922_19591.n42 0.246907
R49582 a_35922_19591.n39 a_35922_19591.n38 0.246907
R49583 a_35922_19591.n56 a_35922_19591.n57 0.246907
R49584 a_35922_19591.n55 a_35922_19591.n54 0.246907
R49585 a_35922_19591.n90 a_35922_19591.n89 0.0201939
R49586 a_35922_19591.n36 a_35922_19591.n34 0.246907
R49587 a_35922_19591.n33 a_35922_19591.n31 0.246907
R49588 a_35922_19591.n4 a_35922_19591.n5 0.260442
R49589 a_35922_19591.n26 a_35922_19591.n16 0.591264
R49590 a_35922_19591.n12 a_35922_19591.n13 0.310971
R49591 a_35922_19591.n30 a_35922_19591.n29 0.591264
R49592 a_35922_19591.n28 a_35922_19591.n100 0.332154
R49593 a_35922_19591.n150 a_35922_19591.n140 4.5005
R49594 a_35922_19591.n126 a_35922_19591.n149 4.5005
R49595 a_35922_19591.n148 a_35922_19591.n125 4.5005
R49596 a_35922_19591.n147 a_35922_19591.n146 4.5005
R49597 a_35922_19591.n124 a_35922_19591.n122 4.5005
R49598 a_35922_19591.n123 a_35922_19591.n145 4.5005
R49599 a_35922_19591.n144 a_35922_19591.n141 4.5005
R49600 a_35922_19591.n206 a_35922_19591.n205 4.5005
R49601 a_35922_19591.n115 a_35922_19591.n113 4.5005
R49602 a_35922_19591.n114 a_35922_19591.n204 4.5005
R49603 a_35922_19591.n203 a_35922_19591.n116 4.5005
R49604 a_35922_19591.n202 a_35922_19591.n118 4.5005
R49605 a_35922_19591.n117 a_35922_19591.n154 4.5005
R49606 a_35922_19591.n201 a_35922_19591.n200 4.5005
R49607 a_35922_19591.n199 a_35922_19591.n119 4.5005
R49608 a_35922_19591.n198 a_35922_19591.n197 4.5005
R49609 a_35922_19591.n196 a_35922_19591.n155 4.5005
R49610 a_35922_19591.n181 a_35922_19591.n180 4.5005
R49611 a_35922_19591.n112 a_35922_19591.n182 4.5005
R49612 a_35922_19591.n183 a_35922_19591.n158 4.5005
R49613 a_35922_19591.n185 a_35922_19591.n184 4.5005
R49614 a_35922_19591.n111 a_35922_19591.n186 4.5005
R49615 a_35922_19591.n187 a_35922_19591.n157 4.5005
R49616 a_35922_19591.n189 a_35922_19591.n188 4.5005
R49617 a_35922_19591.n190 a_35922_19591.n110 4.5005
R49618 a_35922_19591.n192 a_35922_19591.n191 4.5005
R49619 a_35922_19591.n193 a_35922_19591.n156 4.5005
R49620 a_35922_19591.n176 a_35922_19591.n175 4.5005
R49621 a_35922_19591.n174 a_35922_19591.n106 4.5005
R49622 a_35922_19591.n173 a_35922_19591.n172 4.5005
R49623 a_35922_19591.n171 a_35922_19591.n165 4.5005
R49624 a_35922_19591.n107 a_35922_19591.n170 4.5005
R49625 a_35922_19591.n169 a_35922_19591.n168 4.5005
R49626 a_35922_19591.n167 a_35922_19591.n166 4.5005
R49627 a_35922_19591.n8 a_35922_19591.n7 0.260442
R49628 a_35922_19591.n21 a_35922_19591.n20 0.591264
R49629 a_35922_19591.n10 a_35922_19591.n11 0.310971
R49630 a_35922_19591.n23 a_35922_19591.n24 0.591264
R49631 a_35922_19591.n22 a_35922_19591.n101 0.332154
R49632 a_35922_19591.n226 a_35922_19591.n225 4.5005
R49633 a_35922_19591.n138 a_35922_19591.n105 4.5005
R49634 a_35922_19591.n104 a_35922_19591.n129 4.5005
R49635 a_35922_19591.n137 a_35922_19591.n136 4.5005
R49636 a_35922_19591.n135 a_35922_19591.n103 4.5005
R49637 a_35922_19591.n102 a_35922_19591.n130 4.5005
R49638 a_35922_19591.n134 a_35922_19591.n133 4.5005
R49639 a_35922_19591.n222 a_35922_19591.n127 3.97759
R49640 a_35922_19591.n240 a_35922_19591.n239 3.0252
R49641 a_35922_19591.n232 a_35922_19591.n231 2.35922
R49642 a_35922_19591.n237 a_35922_19591.n63 2.34557
R49643 a_35922_19591.n208 a_35922_19591.n139 2.30989
R49644 a_35922_19591.n163 a_35922_19591.n93 2.30989
R49645 a_35922_19591.n195 a_35922_19591.n194 2.25752
R49646 a_35922_19591.n71 a_35922_19591.n70 0.427602
R49647 a_35922_19591.n69 a_35922_19591.n68 0.427602
R49648 a_35922_19591.n67 a_35922_19591.n66 0.427602
R49649 a_35922_19591.n65 a_35922_19591.n64 0.427602
R49650 a_35922_19591.n83 a_35922_19591.n82 0.420727
R49651 a_35922_19591.n81 a_35922_19591.n80 0.420727
R49652 a_35922_19591.n79 a_35922_19591.n78 0.420727
R49653 a_35922_19591.n77 a_35922_19591.n76 0.420727
R49654 a_35922_19591.n207 a_35922_19591.n140 2.16725
R49655 a_35922_19591.n181 a_35922_19591.n164 2.16725
R49656 a_35922_19591.n225 a_35922_19591.n224 2.16725
R49657 a_35922_19591.n42 a_35922_19591.n41 2.96488
R49658 a_35922_19591.n37 a_35922_19591.n75 2.94096
R49659 a_35922_19591.n88 a_35922_19591.n36 2.96488
R49660 a_35922_19591.n73 a_35922_19591.n220 2.94096
R49661 a_35922_19591.n222 a_35922_19591.n221 2.09357
R49662 a_35922_19591.n216 a_35922_19591.n97 2.07182
R49663 a_35922_19591.n217 a_35922_19591.n45 2.07182
R49664 a_35922_19591.n97 a_35922_19591.n46 2.75706
R49665 a_35922_19591.n87 a_35922_19591.n45 2.90773
R49666 a_35922_19591.n58 a_35922_19591.n96 2.75704
R49667 a_35922_19591.n52 a_35922_19591.n85 2.90773
R49668 a_35922_19591.n63 a_35922_19591.n60 1.58959
R49669 a_35922_19591.n96 a_35922_19591.n215 1.5005
R49670 a_35922_19591.n41 a_35922_19591.n216 1.5005
R49671 a_35922_19591.n221 a_35922_19591.n88 1.5005
R49672 a_35922_19591.n220 a_35922_19591.n219 1.5005
R49673 a_35922_19591.n218 a_35922_19591.n52 1.5005
R49674 a_35922_19591.n217 a_35922_19591.n37 1.5005
R49675 a_35922_19591.n214 a_35922_19591.n6 1.5005
R49676 a_35922_19591.n208 a_35922_19591.n207 1.5005
R49677 a_35922_19591.n224 a_35922_19591.n223 1.5005
R49678 a_35922_19591.n211 a_35922_19591.n128 1.5005
R49679 a_35922_19591.n164 a_35922_19591.n163 1.5005
R49680 a_35922_19591.n63 a_35922_19591.n62 1.5005
R49681 a_35922_19591.n63 a_35922_19591.n59 1.5005
R49682 a_35922_19591.n239 a_35922_19591.n238 1.5005
R49683 a_35922_19591.n219 a_35922_19591.n127 1.49172
R49684 a_35922_19591.n216 a_35922_19591.n215 1.47516
R49685 a_35922_19591.n218 a_35922_19591.n217 1.47516
R49686 a_35922_19591.n5 a_35922_19591.t188 9.17619
R49687 a_35922_19591.n7 a_35922_19591.t18 9.17619
R49688 a_35922_19591.n223 a_35922_19591.n222 1.37253
R49689 a_35922_19591.n230 a_35922_19591.n229 1.37253
R49690 a_35922_19591.n29 a_35922_19591.n27 1.24866
R49691 a_35922_19591.n16 a_35922_19591.n25 1.24866
R49692 a_35922_19591.n212 a_35922_19591.n23 1.24866
R49693 a_35922_19591.n20 a_35922_19591.n19 1.24866
R49694 a_35922_19591.n159 a_35922_19591.n4 1.24629
R49695 a_35922_19591.n209 a_35922_19591.n8 1.24629
R49696 a_35922_19591.n214 a_35922_19591.n208 1.23709
R49697 a_35922_19591.n163 a_35922_19591.n128 1.23709
R49698 a_35922_19591.n227 a_35922_19591.n226 1.22261
R49699 a_35922_19591.n180 a_35922_19591.n179 1.22261
R49700 a_35922_19591.n151 a_35922_19591.n150 1.22261
R49701 a_35922_19591.n3 a_35922_19591.n2 1.21313
R49702 a_35922_19591.n177 a_35922_19591.n176 1.21313
R49703 a_35922_19591.n205 a_35922_19591.n153 1.21313
R49704 a_35922_19591.n144 a_35922_19591.n143 1.12904
R49705 a_35922_19591.n133 a_35922_19591.n132 1.12904
R49706 a_35922_19591.n223 a_35922_19591.n214 0.809892
R49707 a_35922_19591.n229 a_35922_19591.n128 0.809892
R49708 a_35922_19591.n26 a_35922_19591.n139 1.14908
R49709 a_35922_19591.n93 a_35922_19591.n30 1.14908
R49710 a_35922_19591.n6 a_35922_19591.n21 1.14908
R49711 a_35922_19591.n24 a_35922_19591.n211 1.14908
R49712 a_35922_19591.n207 a_35922_19591.n206 0.71825
R49713 a_35922_19591.n175 a_35922_19591.n164 0.71825
R49714 a_35922_19591.n224 a_35922_19591.n1 1.69988
R49715 a_35922_19591.n228 a_35922_19591.n227 0.673132
R49716 a_35922_19591.n2 a_35922_19591.n228 0.673132
R49717 a_35922_19591.n162 a_35922_19591.n161 0.673132
R49718 a_35922_19591.n27 a_35922_19591.n162 0.673132
R49719 a_35922_19591.n160 a_35922_19591.n159 0.673132
R49720 a_35922_19591.n25 a_35922_19591.n160 0.673132
R49721 a_35922_19591.n179 a_35922_19591.n178 0.673132
R49722 a_35922_19591.n178 a_35922_19591.n177 0.673132
R49723 a_35922_19591.n152 a_35922_19591.n151 0.673132
R49724 a_35922_19591.n153 a_35922_19591.n152 0.673132
R49725 a_35922_19591.n9 a_35922_19591.n213 0.673132
R49726 a_35922_19591.n213 a_35922_19591.n212 0.673132
R49727 a_35922_19591.n210 a_35922_19591.n209 0.673132
R49728 a_35922_19591.n19 a_35922_19591.n210 0.673132
R49729 a_35922_19591.n230 a_35922_19591.n127 0.602344
R49730 a_35922_19591.n221 a_35922_19591.n215 0.571818
R49731 a_35922_19591.n219 a_35922_19591.n218 0.571818
R49732 a_35922_19591.n59 a_35922_19591.n234 0.487111
R49733 a_35922_19591.n61 a_35922_19591.n236 0.487111
R49734 a_35922_19591.n60 a_35922_19591.n233 0.487111
R49735 a_35922_19591.n62 a_35922_19591.n235 0.487111
R49736 a_35922_19591.n109 a_35922_19591.n108 0.321834
R49737 a_35922_19591.n102 a_35922_19591.n134 0.379447
R49738 a_35922_19591.n104 a_35922_19591.n137 0.379447
R49739 a_35922_19591.n172 a_35922_19591.n171 0.379447
R49740 a_35922_19591.n168 a_35922_19591.n167 0.379447
R49741 a_35922_19591.n193 a_35922_19591.n192 0.379447
R49742 a_35922_19591.n188 a_35922_19591.n187 0.379447
R49743 a_35922_19591.n184 a_35922_19591.n183 0.379447
R49744 a_35922_19591.n114 a_35922_19591.n116 0.379447
R49745 a_35922_19591.n117 a_35922_19591.n201 0.379447
R49746 a_35922_19591.n197 a_35922_19591.n196 0.379447
R49747 a_35922_19591.n123 a_35922_19591.n141 0.379447
R49748 a_35922_19591.n146 a_35922_19591.n125 0.379447
R49749 a_35922_19591.n26 a_35922_19591.n18 1.14166
R49750 a_35922_19591.n93 a_35922_19591.n13 2.75347
R49751 a_35922_19591.n100 a_35922_19591.n30 1.60203
R49752 a_35922_19591.n15 a_35922_19591.n21 1.14166
R49753 a_35922_19591.n211 a_35922_19591.n11 2.75347
R49754 a_35922_19591.n101 a_35922_19591.n24 1.60203
R49755 a_35922_19591.n145 a_35922_19591.n144 0.3605
R49756 a_35922_19591.n148 a_35922_19591.n147 0.3605
R49757 a_35922_19591.n204 a_35922_19591.n203 0.3605
R49758 a_35922_19591.n200 a_35922_19591.n154 0.3605
R49759 a_35922_19591.n198 a_35922_19591.n155 0.3605
R49760 a_35922_19591.n191 a_35922_19591.n156 0.3605
R49761 a_35922_19591.n189 a_35922_19591.n157 0.3605
R49762 a_35922_19591.n185 a_35922_19591.n158 0.3605
R49763 a_35922_19591.n173 a_35922_19591.n165 0.3605
R49764 a_35922_19591.n169 a_35922_19591.n166 0.3605
R49765 a_35922_19591.n133 a_35922_19591.n130 0.3605
R49766 a_35922_19591.n136 a_35922_19591.n129 0.3605
R49767 a_35922_19591.n132 a_35922_19591.n131 0.327481
R49768 a_35922_19591.n143 a_35922_19591.n142 0.327481
R49769 a_35922_19591.n195 a_35922_19591.n156 0.208099
R49770 a_35922_19591.n103 a_35922_19591.n102 0.147342
R49771 a_35922_19591.n105 a_35922_19591.n104 0.147342
R49772 a_35922_19591.n176 a_35922_19591.n106 0.147342
R49773 a_35922_19591.n171 a_35922_19591.n107 0.147342
R49774 a_35922_19591.n192 a_35922_19591.n110 0.147342
R49775 a_35922_19591.n187 a_35922_19591.n111 0.147342
R49776 a_35922_19591.n183 a_35922_19591.n112 0.147342
R49777 a_35922_19591.n205 a_35922_19591.n115 0.147342
R49778 a_35922_19591.n118 a_35922_19591.n116 0.147342
R49779 a_35922_19591.n201 a_35922_19591.n119 0.147342
R49780 a_35922_19591.n124 a_35922_19591.n123 0.147342
R49781 a_35922_19591.n126 a_35922_19591.n125 0.147342
R49782 a_35922_19591.n60 a_35922_19591.n232 0.146729
R49783 a_35922_19591.n134 a_35922_19591.n131 0.142605
R49784 a_35922_19591.n194 a_35922_19591.n193 0.142605
R49785 a_35922_19591.n142 a_35922_19591.n141 0.142605
R49786 a_35922_19591.n69 a_35922_19591.n89 2.03311
R49787 a_35922_19591.n35 a_35922_19591.n69 2.04491
R49788 a_35922_19591.n32 a_35922_19591.n35 4.37762
R49789 a_35922_19591.n71 a_35922_19591.n32 1.87961
R49790 a_35922_19591.n71 a_35922_19591.n73 2.19836
R49791 a_35922_19591.n81 a_35922_19591.n98 2.03667
R49792 a_35922_19591.n51 a_35922_19591.n81 2.2172
R49793 a_35922_19591.n51 a_35922_19591.n49 4.49278
R49794 a_35922_19591.n83 a_35922_19591.n49 1.82125
R49795 a_35922_19591.n83 a_35922_19591.n87 2.19319
R49796 a_35922_19591.n98 a_35922_19591.n97 1.65342
R49797 a_35922_19591.n47 a_35922_19591.n46 4.34534
R49798 a_35922_19591.n47 a_35922_19591.n45 1.50598
R49799 a_35922_19591.n65 a_35922_19591.n92 2.03311
R49800 a_35922_19591.n44 a_35922_19591.n65 2.04491
R49801 a_35922_19591.n40 a_35922_19591.n44 4.37762
R49802 a_35922_19591.n67 a_35922_19591.n40 1.87961
R49803 a_35922_19591.n75 a_35922_19591.n67 2.19836
R49804 a_35922_19591.n41 a_35922_19591.n92 1.65903
R49805 a_35922_19591.n42 a_35922_19591.n38 4.49309
R49806 a_35922_19591.n38 a_35922_19591.n37 1.44546
R49807 a_35922_19591.n77 a_35922_19591.n95 2.03657
R49808 a_35922_19591.n77 a_35922_19591.n57 2.21715
R49809 a_35922_19591.n55 a_35922_19591.n57 4.49317
R49810 a_35922_19591.n79 a_35922_19591.n55 1.82113
R49811 a_35922_19591.n85 a_35922_19591.n79 2.19319
R49812 a_35922_19591.n96 a_35922_19591.n95 1.65366
R49813 a_35922_19591.n53 a_35922_19591.n58 4.34574
R49814 a_35922_19591.n53 a_35922_19591.n52 1.50586
R49815 a_35922_19591.n196 a_35922_19591.n120 0.152079
R49816 a_35922_19591.n150 a_35922_19591.n126 0.147342
R49817 a_35922_19591.n146 a_35922_19591.n124 0.147342
R49818 a_35922_19591.n89 a_35922_19591.n88 1.65903
R49819 a_35922_19591.n36 a_35922_19591.n33 4.49309
R49820 a_35922_19591.n33 a_35922_19591.n220 1.44546
R49821 a_35922_19591.n139 a_35922_19591.n5 2.8103
R49822 a_35922_19591.n13 a_35922_19591.n18 4.38327
R49823 a_35922_19591.n145 a_35922_19591.n122 0.14
R49824 a_35922_19591.n147 a_35922_19591.n122 0.14
R49825 a_35922_19591.n149 a_35922_19591.n148 0.14
R49826 a_35922_19591.n149 a_35922_19591.n140 0.14
R49827 a_35922_19591.n206 a_35922_19591.n113 0.14
R49828 a_35922_19591.n204 a_35922_19591.n113 0.14
R49829 a_35922_19591.n203 a_35922_19591.n202 0.14
R49830 a_35922_19591.n202 a_35922_19591.n154 0.14
R49831 a_35922_19591.n200 a_35922_19591.n199 0.14
R49832 a_35922_19591.n199 a_35922_19591.n198 0.14
R49833 a_35922_19591.n121 a_35922_19591.n155 0.208134
R49834 a_35922_19591.n121 a_35922_19591.n195 3.10882
R49835 a_35922_19591.n167 a_35922_19591.n108 0.152079
R49836 a_35922_19591.n197 a_35922_19591.n119 0.147342
R49837 a_35922_19591.n118 a_35922_19591.n117 0.147342
R49838 a_35922_19591.n115 a_35922_19591.n114 0.147342
R49839 a_35922_19591.n180 a_35922_19591.n112 0.147342
R49840 a_35922_19591.n184 a_35922_19591.n111 0.147342
R49841 a_35922_19591.n188 a_35922_19591.n110 0.147342
R49842 a_35922_19591.n191 a_35922_19591.n190 0.14
R49843 a_35922_19591.n190 a_35922_19591.n189 0.14
R49844 a_35922_19591.n186 a_35922_19591.n157 0.14
R49845 a_35922_19591.n186 a_35922_19591.n185 0.14
R49846 a_35922_19591.n182 a_35922_19591.n158 0.14
R49847 a_35922_19591.n182 a_35922_19591.n181 0.14
R49848 a_35922_19591.n175 a_35922_19591.n174 0.14
R49849 a_35922_19591.n174 a_35922_19591.n173 0.14
R49850 a_35922_19591.n170 a_35922_19591.n165 0.14
R49851 a_35922_19591.n170 a_35922_19591.n169 0.14
R49852 a_35922_19591.n109 a_35922_19591.n166 1.12757
R49853 a_35922_19591.n168 a_35922_19591.n107 0.147342
R49854 a_35922_19591.n172 a_35922_19591.n106 0.147342
R49855 a_35922_19591.n226 a_35922_19591.n105 0.147342
R49856 a_35922_19591.n137 a_35922_19591.n103 0.147342
R49857 a_35922_19591.n7 a_35922_19591.n6 2.8103
R49858 a_35922_19591.n15 a_35922_19591.n11 4.38327
R49859 a_35922_19591.n135 a_35922_19591.n130 0.14
R49860 a_35922_19591.n136 a_35922_19591.n135 0.14
R49861 a_35922_19591.n138 a_35922_19591.n129 0.14
R49862 a_35922_19591.n225 a_35922_19591.n138 0.14
R49863 a_35922_19591.n0 a_35922_19591.n1 5.18575
R49864 a_35922_19591.n161 a_35922_19591.n12 2.13563
R49865 a_35922_19591.n10 a_35922_19591.n9 2.13563
R49866 a_35922_19591.n17 a_35922_19591.n16 2.13445
R49867 a_35922_19591.n20 a_35922_19591.n14 2.13445
R49868 a_35922_19591.n63 a_35922_19591.n61 1.89911
R49869 a_35922_19591.n29 a_35922_19591.n28 1.36353
R49870 a_35922_19591.n23 a_35922_19591.n22 1.36353
R49871 a_35922_19591.n0 a_35922_19591.t139 8.54486
R49872 a_35922_19591.n229 a_35922_19591.n0 3.64386
R49873 a_52635_48695.n83 a_52635_48695.n81 7.22198
R49874 a_52635_48695.n119 a_52635_48695.n118 7.22198
R49875 a_52635_48695.n68 a_52635_48695.t125 6.77653
R49876 a_52635_48695.n54 a_52635_48695.t161 6.77653
R49877 a_52635_48695.n60 a_52635_48695.t142 6.7761
R49878 a_52635_48695.n58 a_52635_48695.t92 6.7761
R49879 a_52635_48695.n23 a_52635_48695.t102 6.77231
R49880 a_52635_48695.n33 a_52635_48695.t130 6.77231
R49881 a_52635_48695.n192 a_52635_48695.n191 6.50088
R49882 a_52635_48695.n162 a_52635_48695.n161 6.50088
R49883 a_52635_48695.n72 a_52635_48695.t135 5.50607
R49884 a_52635_48695.n69 a_52635_48695.t99 5.50607
R49885 a_52635_48695.n99 a_52635_48695.t174 5.50607
R49886 a_52635_48695.n55 a_52635_48695.t144 5.50607
R49887 a_52635_48695.n71 a_52635_48695.t138 5.50475
R49888 a_52635_48695.n75 a_52635_48695.t123 5.50475
R49889 a_52635_48695.n76 a_52635_48695.t131 5.50475
R49890 a_52635_48695.n70 a_52635_48695.t127 5.50475
R49891 a_52635_48695.n98 a_52635_48695.t175 5.50475
R49892 a_52635_48695.n102 a_52635_48695.t157 5.50475
R49893 a_52635_48695.n103 a_52635_48695.t170 5.50475
R49894 a_52635_48695.n56 a_52635_48695.t165 5.50475
R49895 a_52635_48695.n137 a_52635_48695.n135 4.92758
R49896 a_52635_48695.n38 a_52635_48695.n36 4.92758
R49897 a_52635_48695.n6 a_52635_48695.n175 4.92217
R49898 a_52635_48695.n13 a_52635_48695.n142 4.92217
R49899 a_52635_48695.n183 a_52635_48695.n0 3.65107
R49900 a_52635_48695.n182 a_52635_48695.n1 3.65107
R49901 a_52635_48695.n181 a_52635_48695.n2 3.65107
R49902 a_52635_48695.n180 a_52635_48695.n3 3.65107
R49903 a_52635_48695.n178 a_52635_48695.n4 3.65107
R49904 a_52635_48695.n177 a_52635_48695.n5 3.65107
R49905 a_52635_48695.n176 a_52635_48695.n6 3.65107
R49906 a_52635_48695.n7 a_52635_48695.n149 3.65107
R49907 a_52635_48695.n8 a_52635_48695.n148 3.65107
R49908 a_52635_48695.n9 a_52635_48695.n147 3.65107
R49909 a_52635_48695.n10 a_52635_48695.n146 3.65107
R49910 a_52635_48695.n145 a_52635_48695.n11 3.65107
R49911 a_52635_48695.n144 a_52635_48695.n12 3.65107
R49912 a_52635_48695.n143 a_52635_48695.n13 3.65107
R49913 a_52635_48695.n14 a_52635_48695.n125 4.0312
R49914 a_52635_48695.t119 a_52635_48695.n15 5.5012
R49915 a_52635_48695.t116 a_52635_48695.n16 5.5012
R49916 a_52635_48695.n124 a_52635_48695.n17 4.0312
R49917 a_52635_48695.t98 a_52635_48695.n18 5.5012
R49918 a_52635_48695.t111 a_52635_48695.n19 5.5012
R49919 a_52635_48695.n123 a_52635_48695.n20 4.0312
R49920 a_52635_48695.t108 a_52635_48695.n21 5.5012
R49921 a_52635_48695.t88 a_52635_48695.n22 5.5012
R49922 a_52635_48695.n51 a_52635_48695.n23 4.0312
R49923 a_52635_48695.n24 a_52635_48695.n93 4.0312
R49924 a_52635_48695.t147 a_52635_48695.n25 5.5012
R49925 a_52635_48695.t145 a_52635_48695.n26 5.5012
R49926 a_52635_48695.n92 a_52635_48695.n27 4.0312
R49927 a_52635_48695.t126 a_52635_48695.n28 5.5012
R49928 a_52635_48695.t139 a_52635_48695.n29 5.5012
R49929 a_52635_48695.n91 a_52635_48695.n30 4.0312
R49930 a_52635_48695.t136 a_52635_48695.n31 5.5012
R49931 a_52635_48695.t110 a_52635_48695.n32 5.5012
R49932 a_52635_48695.n89 a_52635_48695.n33 4.0312
R49933 a_52635_48695.n82 a_52635_48695.t128 4.24002
R49934 a_52635_48695.n62 a_52635_48695.t95 4.24002
R49935 a_52635_48695.n117 a_52635_48695.t100 4.24002
R49936 a_52635_48695.n108 a_52635_48695.t163 4.24002
R49937 a_52635_48695.n156 a_52635_48695.t71 4.06712
R49938 a_52635_48695.n154 a_52635_48695.t62 4.06712
R49939 a_52635_48695.n186 a_52635_48695.t79 4.06712
R49940 a_52635_48695.n48 a_52635_48695.t66 4.06712
R49941 a_52635_48695.n60 a_52635_48695.n59 4.03475
R49942 a_52635_48695.n74 a_52635_48695.n73 4.03475
R49943 a_52635_48695.n78 a_52635_48695.n77 4.03475
R49944 a_52635_48695.n68 a_52635_48695.n67 4.03475
R49945 a_52635_48695.n58 a_52635_48695.n57 4.03475
R49946 a_52635_48695.n101 a_52635_48695.n100 4.03475
R49947 a_52635_48695.n105 a_52635_48695.n104 4.03475
R49948 a_52635_48695.n54 a_52635_48695.n53 4.03475
R49949 a_52635_48695.n128 a_52635_48695.n43 3.97307
R49950 a_52635_48695.n187 a_52635_48695.n185 3.96014
R49951 a_52635_48695.n157 a_52635_48695.n134 3.96014
R49952 a_52635_48695.n156 a_52635_48695.t74 3.86107
R49953 a_52635_48695.n154 a_52635_48695.t63 3.86107
R49954 a_52635_48695.n186 a_52635_48695.t0 3.86107
R49955 a_52635_48695.n48 a_52635_48695.t75 3.86107
R49956 a_52635_48695.n139 a_52635_48695.n137 3.79678
R49957 a_52635_48695.n171 a_52635_48695.n169 3.79678
R49958 a_52635_48695.n40 a_52635_48695.n38 3.79678
R49959 a_52635_48695.n130 a_52635_48695.n35 3.79678
R49960 a_52635_48695.n82 a_52635_48695.t106 3.68818
R49961 a_52635_48695.n62 a_52635_48695.t166 3.68818
R49962 a_52635_48695.n117 a_52635_48695.t148 3.68818
R49963 a_52635_48695.n108 a_52635_48695.t114 3.68818
R49964 a_52635_48695.n132 a_52635_48695.n131 3.65581
R49965 a_52635_48695.n173 a_52635_48695.n172 3.65581
R49966 a_52635_48695.n171 a_52635_48695.n170 3.65581
R49967 a_52635_48695.n169 a_52635_48695.n168 3.65581
R49968 a_52635_48695.n167 a_52635_48695.n166 3.65581
R49969 a_52635_48695.n141 a_52635_48695.n140 3.65581
R49970 a_52635_48695.n139 a_52635_48695.n138 3.65581
R49971 a_52635_48695.n137 a_52635_48695.n136 3.65581
R49972 a_52635_48695.n130 a_52635_48695.n129 3.65581
R49973 a_52635_48695.n35 a_52635_48695.n34 3.65581
R49974 a_52635_48695.n197 a_52635_48695.n196 3.65581
R49975 a_52635_48695.n42 a_52635_48695.n41 3.65581
R49976 a_52635_48695.n40 a_52635_48695.n39 3.65581
R49977 a_52635_48695.n38 a_52635_48695.n37 3.65581
R49978 a_52635_48695.n167 a_52635_48695.n165 3.64443
R49979 a_52635_48695.n196 a_52635_48695.n195 3.64443
R49980 a_52635_48695.n3 a_52635_48695.n179 3.64223
R49981 a_52635_48695.n150 a_52635_48695.n10 3.64223
R49982 a_52635_48695.n88 a_52635_48695.n87 3.23904
R49983 a_52635_48695.n116 a_52635_48695.n50 3.23904
R49984 a_52635_48695.n86 a_52635_48695.n85 2.77002
R49985 a_52635_48695.n65 a_52635_48695.n64 2.77002
R49986 a_52635_48695.n115 a_52635_48695.n114 2.77002
R49987 a_52635_48695.n111 a_52635_48695.n110 2.77002
R49988 a_52635_48695.n66 a_52635_48695.n62 2.73714
R49989 a_52635_48695.n112 a_52635_48695.n108 2.73714
R49990 a_52635_48695.n49 a_52635_48695.n47 2.73714
R49991 a_52635_48695.n155 a_52635_48695.n153 2.73714
R49992 a_52635_48695.n76 a_52635_48695.n75 2.60203
R49993 a_52635_48695.n103 a_52635_48695.n102 2.60203
R49994 a_52635_48695.n160 a_52635_48695.n158 2.59712
R49995 a_52635_48695.n153 a_52635_48695.n151 2.59712
R49996 a_52635_48695.n190 a_52635_48695.n188 2.59712
R49997 a_52635_48695.n47 a_52635_48695.n45 2.59712
R49998 a_52635_48695.n70 a_52635_48695.n69 2.52436
R49999 a_52635_48695.n72 a_52635_48695.n71 2.52436
R50000 a_52635_48695.n56 a_52635_48695.n55 2.52436
R50001 a_52635_48695.n99 a_52635_48695.n98 2.52436
R50002 a_52635_48695.n192 a_52635_48695.n49 2.46014
R50003 a_52635_48695.n162 a_52635_48695.n155 2.46014
R50004 a_52635_48695.n160 a_52635_48695.n159 2.39107
R50005 a_52635_48695.n153 a_52635_48695.n152 2.39107
R50006 a_52635_48695.n190 a_52635_48695.n189 2.39107
R50007 a_52635_48695.n47 a_52635_48695.n46 2.39107
R50008 a_52635_48695.n86 a_52635_48695.n84 2.21818
R50009 a_52635_48695.n65 a_52635_48695.n63 2.21818
R50010 a_52635_48695.n115 a_52635_48695.n113 2.21818
R50011 a_52635_48695.n111 a_52635_48695.n109 2.21818
R50012 a_52635_48695.n80 a_52635_48695.n79 2.13841
R50013 a_52635_48695.n88 a_52635_48695.n61 2.13841
R50014 a_52635_48695.n163 a_52635_48695.n150 2.0852
R50015 a_52635_48695.n133 a_52635_48695.n128 2.02864
R50016 a_52635_48695.n121 a_52635_48695.n43 1.76168
R50017 a_52635_48695.n81 a_52635_48695.n66 1.73904
R50018 a_52635_48695.n119 a_52635_48695.n112 1.73904
R50019 a_52635_48695.n174 a_52635_48695.n173 1.73609
R50020 a_52635_48695.n133 a_52635_48695.n132 1.73609
R50021 a_52635_48695.n120 a_52635_48695.n119 1.5005
R50022 a_52635_48695.n107 a_52635_48695.n106 1.5005
R50023 a_52635_48695.n90 a_52635_48695.n52 1.5005
R50024 a_52635_48695.n81 a_52635_48695.n80 1.5005
R50025 a_52635_48695.n122 a_52635_48695.n121 1.5005
R50026 a_52635_48695.n127 a_52635_48695.n126 1.5005
R50027 a_52635_48695.n97 a_52635_48695.n96 1.5005
R50028 a_52635_48695.n95 a_52635_48695.n94 1.5005
R50029 a_52635_48695.n163 a_52635_48695.n162 1.5005
R50030 a_52635_48695.n193 a_52635_48695.n192 1.5005
R50031 a_52635_48695.n165 a_52635_48695.n164 1.5005
R50032 a_52635_48695.n179 a_52635_48695.n44 1.5005
R50033 a_52635_48695.n195 a_52635_48695.n194 1.5005
R50034 a_52635_48695.n131 a_52635_48695.t46 1.4705
R50035 a_52635_48695.n131 a_52635_48695.t21 1.4705
R50036 a_52635_48695.n158 a_52635_48695.t57 1.4705
R50037 a_52635_48695.n158 a_52635_48695.t37 1.4705
R50038 a_52635_48695.n159 a_52635_48695.t59 1.4705
R50039 a_52635_48695.n159 a_52635_48695.t40 1.4705
R50040 a_52635_48695.n151 a_52635_48695.t36 1.4705
R50041 a_52635_48695.n151 a_52635_48695.t29 1.4705
R50042 a_52635_48695.n152 a_52635_48695.t38 1.4705
R50043 a_52635_48695.n152 a_52635_48695.t30 1.4705
R50044 a_52635_48695.n183 a_52635_48695.t33 1.4705
R50045 a_52635_48695.n183 a_52635_48695.t10 1.4705
R50046 a_52635_48695.n182 a_52635_48695.t5 1.4705
R50047 a_52635_48695.n182 a_52635_48695.t51 1.4705
R50048 a_52635_48695.n181 a_52635_48695.t86 1.4705
R50049 a_52635_48695.n181 a_52635_48695.t4 1.4705
R50050 a_52635_48695.n180 a_52635_48695.t67 1.4705
R50051 a_52635_48695.n180 a_52635_48695.t27 1.4705
R50052 a_52635_48695.n178 a_52635_48695.t8 1.4705
R50053 a_52635_48695.n178 a_52635_48695.t85 1.4705
R50054 a_52635_48695.n177 a_52635_48695.t80 1.4705
R50055 a_52635_48695.n177 a_52635_48695.t32 1.4705
R50056 a_52635_48695.n176 a_52635_48695.t72 1.4705
R50057 a_52635_48695.n176 a_52635_48695.t52 1.4705
R50058 a_52635_48695.n175 a_52635_48695.t73 1.4705
R50059 a_52635_48695.n175 a_52635_48695.t23 1.4705
R50060 a_52635_48695.n172 a_52635_48695.t41 1.4705
R50061 a_52635_48695.n172 a_52635_48695.t18 1.4705
R50062 a_52635_48695.n170 a_52635_48695.t14 1.4705
R50063 a_52635_48695.n170 a_52635_48695.t53 1.4705
R50064 a_52635_48695.n168 a_52635_48695.t7 1.4705
R50065 a_52635_48695.n168 a_52635_48695.t11 1.4705
R50066 a_52635_48695.n166 a_52635_48695.t77 1.4705
R50067 a_52635_48695.n166 a_52635_48695.t31 1.4705
R50068 a_52635_48695.n140 a_52635_48695.t15 1.4705
R50069 a_52635_48695.n140 a_52635_48695.t6 1.4705
R50070 a_52635_48695.n138 a_52635_48695.t3 1.4705
R50071 a_52635_48695.n138 a_52635_48695.t39 1.4705
R50072 a_52635_48695.n136 a_52635_48695.t81 1.4705
R50073 a_52635_48695.n136 a_52635_48695.t55 1.4705
R50074 a_52635_48695.n135 a_52635_48695.t82 1.4705
R50075 a_52635_48695.n135 a_52635_48695.t24 1.4705
R50076 a_52635_48695.n149 a_52635_48695.t26 1.4705
R50077 a_52635_48695.n149 a_52635_48695.t84 1.4705
R50078 a_52635_48695.n148 a_52635_48695.t78 1.4705
R50079 a_52635_48695.n148 a_52635_48695.t47 1.4705
R50080 a_52635_48695.n147 a_52635_48695.t69 1.4705
R50081 a_52635_48695.n147 a_52635_48695.t76 1.4705
R50082 a_52635_48695.n146 a_52635_48695.t56 1.4705
R50083 a_52635_48695.n146 a_52635_48695.t22 1.4705
R50084 a_52635_48695.n145 a_52635_48695.t83 1.4705
R50085 a_52635_48695.n145 a_52635_48695.t68 1.4705
R50086 a_52635_48695.n144 a_52635_48695.t65 1.4705
R50087 a_52635_48695.n144 a_52635_48695.t25 1.4705
R50088 a_52635_48695.n143 a_52635_48695.t60 1.4705
R50089 a_52635_48695.n143 a_52635_48695.t50 1.4705
R50090 a_52635_48695.n142 a_52635_48695.t61 1.4705
R50091 a_52635_48695.n142 a_52635_48695.t16 1.4705
R50092 a_52635_48695.n125 a_52635_48695.t173 1.4705
R50093 a_52635_48695.n125 a_52635_48695.t153 1.4705
R50094 a_52635_48695.n124 a_52635_48695.t146 1.4705
R50095 a_52635_48695.n124 a_52635_48695.t112 1.4705
R50096 a_52635_48695.n123 a_52635_48695.t152 1.4705
R50097 a_52635_48695.n123 a_52635_48695.t121 1.4705
R50098 a_52635_48695.n51 a_52635_48695.t134 1.4705
R50099 a_52635_48695.n51 a_52635_48695.t101 1.4705
R50100 a_52635_48695.n59 a_52635_48695.t94 1.4705
R50101 a_52635_48695.n59 a_52635_48695.t172 1.4705
R50102 a_52635_48695.n73 a_52635_48695.t162 1.4705
R50103 a_52635_48695.n73 a_52635_48695.t132 1.4705
R50104 a_52635_48695.n77 a_52635_48695.t169 1.4705
R50105 a_52635_48695.n77 a_52635_48695.t141 1.4705
R50106 a_52635_48695.n67 a_52635_48695.t154 1.4705
R50107 a_52635_48695.n67 a_52635_48695.t124 1.4705
R50108 a_52635_48695.n84 a_52635_48695.t167 1.4705
R50109 a_52635_48695.n84 a_52635_48695.t120 1.4705
R50110 a_52635_48695.n85 a_52635_48695.t96 1.4705
R50111 a_52635_48695.n85 a_52635_48695.t143 1.4705
R50112 a_52635_48695.n63 a_52635_48695.t158 1.4705
R50113 a_52635_48695.n63 a_52635_48695.t109 1.4705
R50114 a_52635_48695.n64 a_52635_48695.t93 1.4705
R50115 a_52635_48695.n64 a_52635_48695.t133 1.4705
R50116 a_52635_48695.n93 a_52635_48695.t103 1.4705
R50117 a_52635_48695.n93 a_52635_48695.t91 1.4705
R50118 a_52635_48695.n92 a_52635_48695.t168 1.4705
R50119 a_52635_48695.n92 a_52635_48695.t140 1.4705
R50120 a_52635_48695.n91 a_52635_48695.t89 1.4705
R50121 a_52635_48695.n91 a_52635_48695.t149 1.4705
R50122 a_52635_48695.n89 a_52635_48695.t159 1.4705
R50123 a_52635_48695.n89 a_52635_48695.t129 1.4705
R50124 a_52635_48695.n57 a_52635_48695.t137 1.4705
R50125 a_52635_48695.n57 a_52635_48695.t118 1.4705
R50126 a_52635_48695.n100 a_52635_48695.t107 1.4705
R50127 a_52635_48695.n100 a_52635_48695.t171 1.4705
R50128 a_52635_48695.n104 a_52635_48695.t117 1.4705
R50129 a_52635_48695.n104 a_52635_48695.t90 1.4705
R50130 a_52635_48695.n53 a_52635_48695.t97 1.4705
R50131 a_52635_48695.n53 a_52635_48695.t160 1.4705
R50132 a_52635_48695.n113 a_52635_48695.t115 1.4705
R50133 a_52635_48695.n113 a_52635_48695.t155 1.4705
R50134 a_52635_48695.n114 a_52635_48695.t164 1.4705
R50135 a_52635_48695.n114 a_52635_48695.t113 1.4705
R50136 a_52635_48695.n109 a_52635_48695.t105 1.4705
R50137 a_52635_48695.n109 a_52635_48695.t151 1.4705
R50138 a_52635_48695.n110 a_52635_48695.t156 1.4705
R50139 a_52635_48695.n110 a_52635_48695.t104 1.4705
R50140 a_52635_48695.n188 a_52635_48695.t64 1.4705
R50141 a_52635_48695.n188 a_52635_48695.t44 1.4705
R50142 a_52635_48695.n189 a_52635_48695.t70 1.4705
R50143 a_52635_48695.n189 a_52635_48695.t49 1.4705
R50144 a_52635_48695.n45 a_52635_48695.t43 1.4705
R50145 a_52635_48695.n45 a_52635_48695.t34 1.4705
R50146 a_52635_48695.n46 a_52635_48695.t48 1.4705
R50147 a_52635_48695.n46 a_52635_48695.t42 1.4705
R50148 a_52635_48695.n129 a_52635_48695.t19 1.4705
R50149 a_52635_48695.n129 a_52635_48695.t54 1.4705
R50150 a_52635_48695.n34 a_52635_48695.t13 1.4705
R50151 a_52635_48695.n34 a_52635_48695.t17 1.4705
R50152 a_52635_48695.n41 a_52635_48695.t20 1.4705
R50153 a_52635_48695.n41 a_52635_48695.t12 1.4705
R50154 a_52635_48695.n39 a_52635_48695.t9 1.4705
R50155 a_52635_48695.n39 a_52635_48695.t45 1.4705
R50156 a_52635_48695.n37 a_52635_48695.t1 1.4705
R50157 a_52635_48695.n37 a_52635_48695.t58 1.4705
R50158 a_52635_48695.n36 a_52635_48695.t2 1.4705
R50159 a_52635_48695.n36 a_52635_48695.t28 1.4705
R50160 a_52635_48695.t87 a_52635_48695.n197 1.4705
R50161 a_52635_48695.n197 a_52635_48695.t35 1.4705
R50162 a_52635_48695.n87 a_52635_48695.n86 1.46537
R50163 a_52635_48695.n83 a_52635_48695.n82 1.46537
R50164 a_52635_48695.n66 a_52635_48695.n65 1.46537
R50165 a_52635_48695.n116 a_52635_48695.n115 1.46537
R50166 a_52635_48695.n118 a_52635_48695.n117 1.46537
R50167 a_52635_48695.n112 a_52635_48695.n111 1.46537
R50168 a_52635_48695.n157 a_52635_48695.n156 1.46537
R50169 a_52635_48695.n161 a_52635_48695.n160 1.46537
R50170 a_52635_48695.n155 a_52635_48695.n154 1.46537
R50171 a_52635_48695.n187 a_52635_48695.n186 1.46537
R50172 a_52635_48695.n191 a_52635_48695.n190 1.46537
R50173 a_52635_48695.n49 a_52635_48695.n48 1.46537
R50174 a_52635_48695.n194 a_52635_48695.n43 1.42428
R50175 a_52635_48695.n78 a_52635_48695.n76 1.27228
R50176 a_52635_48695.n75 a_52635_48695.n74 1.27228
R50177 a_52635_48695.n87 a_52635_48695.n83 1.27228
R50178 a_52635_48695.n105 a_52635_48695.n103 1.27228
R50179 a_52635_48695.n102 a_52635_48695.n101 1.27228
R50180 a_52635_48695.n118 a_52635_48695.n116 1.27228
R50181 a_52635_48695.n141 a_52635_48695.n139 1.27228
R50182 a_52635_48695.n169 a_52635_48695.n167 1.27228
R50183 a_52635_48695.n173 a_52635_48695.n171 1.27228
R50184 a_52635_48695.n191 a_52635_48695.n187 1.27228
R50185 a_52635_48695.n161 a_52635_48695.n157 1.27228
R50186 a_52635_48695.n196 a_52635_48695.n35 1.27228
R50187 a_52635_48695.n42 a_52635_48695.n40 1.27228
R50188 a_52635_48695.n132 a_52635_48695.n130 1.27228
R50189 a_52635_48695.n69 a_52635_48695.n68 1.26756
R50190 a_52635_48695.n74 a_52635_48695.n72 1.26756
R50191 a_52635_48695.n55 a_52635_48695.n54 1.26756
R50192 a_52635_48695.n101 a_52635_48695.n99 1.26756
R50193 a_52635_48695.n128 a_52635_48695.n127 1.15732
R50194 a_52635_48695.n184 a_52635_48695.n174 0.822966
R50195 a_52635_48695.n164 a_52635_48695.n44 0.822966
R50196 a_52635_48695.n79 a_52635_48695.n70 0.796291
R50197 a_52635_48695.n71 a_52635_48695.n61 0.796291
R50198 a_52635_48695.n106 a_52635_48695.n56 0.796291
R50199 a_52635_48695.n98 a_52635_48695.n97 0.796291
R50200 a_52635_48695.n80 a_52635_48695.n52 0.780703
R50201 a_52635_48695.n121 a_52635_48695.n120 0.780703
R50202 a_52635_48695.n95 a_52635_48695.n88 0.780703
R50203 a_52635_48695.n127 a_52635_48695.n50 0.780703
R50204 a_52635_48695.n185 a_52635_48695.n133 0.639318
R50205 a_52635_48695.n174 a_52635_48695.n134 0.639318
R50206 a_52635_48695.n194 a_52635_48695.n193 0.639318
R50207 a_52635_48695.n164 a_52635_48695.n163 0.639318
R50208 a_52635_48695.n120 a_52635_48695.n107 0.638405
R50209 a_52635_48695.n96 a_52635_48695.n50 0.638405
R50210 a_52635_48695.n107 a_52635_48695.n52 0.628372
R50211 a_52635_48695.n96 a_52635_48695.n95 0.628372
R50212 a_52635_48695.n185 a_52635_48695.n184 0.585196
R50213 a_52635_48695.n193 a_52635_48695.n44 0.585196
R50214 a_52635_48695.n79 a_52635_48695.n78 0.476484
R50215 a_52635_48695.n61 a_52635_48695.n60 0.476484
R50216 a_52635_48695.n106 a_52635_48695.n105 0.476484
R50217 a_52635_48695.n97 a_52635_48695.n58 0.476484
R50218 a_52635_48695.n30 a_52635_48695.n90 0.478684
R50219 a_52635_48695.n94 a_52635_48695.n24 0.478684
R50220 a_52635_48695.n20 a_52635_48695.n122 0.478684
R50221 a_52635_48695.n126 a_52635_48695.n14 0.478684
R50222 a_52635_48695.n165 a_52635_48695.n141 0.236091
R50223 a_52635_48695.n195 a_52635_48695.n42 0.236091
R50224 a_52635_48695.n5 a_52635_48695.n6 3.79678
R50225 a_52635_48695.n4 a_52635_48695.n5 1.27228
R50226 a_52635_48695.n179 a_52635_48695.n4 0.238291
R50227 a_52635_48695.n2 a_52635_48695.n3 1.27228
R50228 a_52635_48695.n1 a_52635_48695.n2 3.79678
R50229 a_52635_48695.n0 a_52635_48695.n1 1.27228
R50230 a_52635_48695.n184 a_52635_48695.n0 1.73829
R50231 a_52635_48695.n12 a_52635_48695.n13 3.79678
R50232 a_52635_48695.n11 a_52635_48695.n12 1.27228
R50233 a_52635_48695.n150 a_52635_48695.n11 0.238291
R50234 a_52635_48695.n9 a_52635_48695.n10 1.27228
R50235 a_52635_48695.n8 a_52635_48695.n9 3.79678
R50236 a_52635_48695.n7 a_52635_48695.n8 1.27228
R50237 a_52635_48695.n134 a_52635_48695.n7 2.32299
R50238 a_52635_48695.n32 a_52635_48695.n33 1.27228
R50239 a_52635_48695.n31 a_52635_48695.n32 2.51878
R50240 a_52635_48695.n90 a_52635_48695.n31 0.794091
R50241 a_52635_48695.n29 a_52635_48695.n30 1.27228
R50242 a_52635_48695.n28 a_52635_48695.n29 2.60203
R50243 a_52635_48695.n27 a_52635_48695.n28 1.27228
R50244 a_52635_48695.n26 a_52635_48695.n27 1.27228
R50245 a_52635_48695.n25 a_52635_48695.n26 2.51878
R50246 a_52635_48695.n94 a_52635_48695.n25 0.794091
R50247 a_52635_48695.t150 a_52635_48695.n24 6.77266
R50248 a_52635_48695.n22 a_52635_48695.n23 1.27228
R50249 a_52635_48695.n21 a_52635_48695.n22 2.51878
R50250 a_52635_48695.n122 a_52635_48695.n21 0.794091
R50251 a_52635_48695.n19 a_52635_48695.n20 1.27228
R50252 a_52635_48695.n18 a_52635_48695.n19 2.60203
R50253 a_52635_48695.n17 a_52635_48695.n18 1.27228
R50254 a_52635_48695.n16 a_52635_48695.n17 1.27228
R50255 a_52635_48695.n15 a_52635_48695.n16 2.51878
R50256 a_52635_48695.n126 a_52635_48695.n15 0.794091
R50257 a_52635_48695.t122 a_52635_48695.n14 6.77266
R50258 a_50751_n19729.n300 a_50751_n19729.t72 12.6064
R50259 a_50751_n19729.t357 a_50751_n19729.n232 10.1674
R50260 a_50751_n19729.n233 a_50751_n19729.t357 10.1674
R50261 a_50751_n19729.t137 a_50751_n19729.n234 10.1674
R50262 a_50751_n19729.n235 a_50751_n19729.t137 10.1674
R50263 a_50751_n19729.t122 a_50751_n19729.n238 10.1674
R50264 a_50751_n19729.n239 a_50751_n19729.t122 10.1674
R50265 a_50751_n19729.t194 a_50751_n19729.n242 10.1674
R50266 a_50751_n19729.n243 a_50751_n19729.t194 10.1674
R50267 a_50751_n19729.t346 a_50751_n19729.n250 10.1674
R50268 a_50751_n19729.n251 a_50751_n19729.t346 10.1674
R50269 a_50751_n19729.n499 a_50751_n19729.t111 10.1674
R50270 a_50751_n19729.t111 a_50751_n19729.n498 10.1674
R50271 a_50751_n19729.n493 a_50751_n19729.t170 10.1674
R50272 a_50751_n19729.n297 a_50751_n19729.t106 10.1674
R50273 a_50751_n19729.t106 a_50751_n19729.n296 10.1674
R50274 a_50751_n19729.n293 a_50751_n19729.t100 10.1674
R50275 a_50751_n19729.t100 a_50751_n19729.n292 10.1674
R50276 a_50751_n19729.n289 a_50751_n19729.t167 10.1674
R50277 a_50751_n19729.t167 a_50751_n19729.n288 10.1674
R50278 a_50751_n19729.t250 a_50751_n19729.n257 10.1674
R50279 a_50751_n19729.n258 a_50751_n19729.t250 10.1674
R50280 a_50751_n19729.t297 a_50751_n19729.n265 10.1674
R50281 a_50751_n19729.n266 a_50751_n19729.t297 10.1674
R50282 a_50751_n19729.n276 a_50751_n19729.t132 10.1674
R50283 a_50751_n19729.t132 a_50751_n19729.n275 10.1674
R50284 a_50751_n19729.n270 a_50751_n19729.t204 10.1674
R50285 a_50751_n19729.n247 a_50751_n19729.t274 10.1674
R50286 a_50751_n19729.t274 a_50751_n19729.n246 10.1674
R50287 a_50751_n19729.t331 a_50751_n19729.n502 10.1674
R50288 a_50751_n19729.n503 a_50751_n19729.t331 10.1674
R50289 a_50751_n19729.t140 a_50751_n19729.n307 10.1674
R50290 a_50751_n19729.n308 a_50751_n19729.t140 10.1674
R50291 a_50751_n19729.t212 a_50751_n19729.n309 10.1674
R50292 a_50751_n19729.n310 a_50751_n19729.t212 10.1674
R50293 a_50751_n19729.t196 a_50751_n19729.n313 10.1674
R50294 a_50751_n19729.n314 a_50751_n19729.t196 10.1674
R50295 a_50751_n19729.n326 a_50751_n19729.t276 10.1674
R50296 a_50751_n19729.t276 a_50751_n19729.n325 10.1674
R50297 a_50751_n19729.n318 a_50751_n19729.t129 10.1674
R50298 a_50751_n19729.t129 a_50751_n19729.n317 10.1674
R50299 a_50751_n19729.t184 a_50751_n19729.n338 10.1674
R50300 a_50751_n19729.n339 a_50751_n19729.t184 10.1674
R50301 a_50751_n19729.n343 a_50751_n19729.t254 10.1674
R50302 a_50751_n19729.n391 a_50751_n19729.t286 10.1674
R50303 a_50751_n19729.t286 a_50751_n19729.n390 10.1674
R50304 a_50751_n19729.n387 a_50751_n19729.t272 10.1674
R50305 a_50751_n19729.t272 a_50751_n19729.n386 10.1674
R50306 a_50751_n19729.n383 a_50751_n19729.t345 10.1674
R50307 a_50751_n19729.t345 a_50751_n19729.n382 10.1674
R50308 a_50751_n19729.t127 a_50751_n19729.n351 10.1674
R50309 a_50751_n19729.n352 a_50751_n19729.t127 10.1674
R50310 a_50751_n19729.t169 a_50751_n19729.n359 10.1674
R50311 a_50751_n19729.n360 a_50751_n19729.t169 10.1674
R50312 a_50751_n19729.n370 a_50751_n19729.t309 10.1674
R50313 a_50751_n19729.t309 a_50751_n19729.n369 10.1674
R50314 a_50751_n19729.n364 a_50751_n19729.t94 10.1674
R50315 a_50751_n19729.t348 a_50751_n19729.n321 10.1674
R50316 a_50751_n19729.n322 a_50751_n19729.t348 10.1674
R50317 a_50751_n19729.n335 a_50751_n19729.t115 10.1674
R50318 a_50751_n19729.t115 a_50751_n19729.n334 10.1674
R50319 a_50751_n19729.n356 a_50751_n19729.t110 10.1674
R50320 a_50751_n19729.t110 a_50751_n19729.n355 10.1674
R50321 a_50751_n19729.t252 a_50751_n19729.n373 10.1674
R50322 a_50751_n19729.n374 a_50751_n19729.t252 10.1674
R50323 a_50751_n19729.t257 a_50751_n19729.n402 10.1674
R50324 a_50751_n19729.n403 a_50751_n19729.t257 10.1674
R50325 a_50751_n19729.t328 a_50751_n19729.n404 10.1674
R50326 a_50751_n19729.n405 a_50751_n19729.t328 10.1674
R50327 a_50751_n19729.t319 a_50751_n19729.n408 10.1674
R50328 a_50751_n19729.n409 a_50751_n19729.t319 10.1674
R50329 a_50751_n19729.n421 a_50751_n19729.t99 10.1674
R50330 a_50751_n19729.t99 a_50751_n19729.n420 10.1674
R50331 a_50751_n19729.n413 a_50751_n19729.t249 10.1674
R50332 a_50751_n19729.t249 a_50751_n19729.n412 10.1674
R50333 a_50751_n19729.t310 a_50751_n19729.n433 10.1674
R50334 a_50751_n19729.n434 a_50751_n19729.t310 10.1674
R50335 a_50751_n19729.n438 a_50751_n19729.t82 10.1674
R50336 a_50751_n19729.n486 a_50751_n19729.t255 10.1674
R50337 a_50751_n19729.t255 a_50751_n19729.n485 10.1674
R50338 a_50751_n19729.n482 a_50751_n19729.t239 10.1674
R50339 a_50751_n19729.t239 a_50751_n19729.n481 10.1674
R50340 a_50751_n19729.n478 a_50751_n19729.t318 10.1674
R50341 a_50751_n19729.t318 a_50751_n19729.n477 10.1674
R50342 a_50751_n19729.t98 a_50751_n19729.n446 10.1674
R50343 a_50751_n19729.n447 a_50751_n19729.t98 10.1674
R50344 a_50751_n19729.t143 a_50751_n19729.n454 10.1674
R50345 a_50751_n19729.n455 a_50751_n19729.t143 10.1674
R50346 a_50751_n19729.n465 a_50751_n19729.t279 10.1674
R50347 a_50751_n19729.t279 a_50751_n19729.n464 10.1674
R50348 a_50751_n19729.n459 a_50751_n19729.t349 10.1674
R50349 a_50751_n19729.t166 a_50751_n19729.n416 10.1674
R50350 a_50751_n19729.n417 a_50751_n19729.t166 10.1674
R50351 a_50751_n19729.n430 a_50751_n19729.t230 10.1674
R50352 a_50751_n19729.t230 a_50751_n19729.n429 10.1674
R50353 a_50751_n19729.n451 a_50751_n19729.t91 10.1674
R50354 a_50751_n19729.t91 a_50751_n19729.n450 10.1674
R50355 a_50751_n19729.t218 a_50751_n19729.n468 10.1674
R50356 a_50751_n19729.n469 a_50751_n19729.t218 10.1674
R50357 a_50751_n19729.n262 a_50751_n19729.t231 10.1674
R50358 a_50751_n19729.t231 a_50751_n19729.n261 10.1674
R50359 a_50751_n19729.t83 a_50751_n19729.n279 10.1674
R50360 a_50751_n19729.n280 a_50751_n19729.t83 10.1674
R50361 a_50751_n19729.n231 a_50751_n19729.t229 10.1674
R50362 a_50751_n19729.t229 a_50751_n19729.n230 10.1674
R50363 a_50751_n19729.t308 a_50751_n19729.n236 10.1674
R50364 a_50751_n19729.n237 a_50751_n19729.t308 10.1674
R50365 a_50751_n19729.t296 a_50751_n19729.n240 10.1674
R50366 a_50751_n19729.n241 a_50751_n19729.t296 10.1674
R50367 a_50751_n19729.t81 a_50751_n19729.n244 10.1674
R50368 a_50751_n19729.n245 a_50751_n19729.t81 10.1674
R50369 a_50751_n19729.t222 a_50751_n19729.n252 10.1674
R50370 a_50751_n19729.n253 a_50751_n19729.t222 10.1674
R50371 a_50751_n19729.n501 a_50751_n19729.t287 10.1674
R50372 a_50751_n19729.t287 a_50751_n19729.n500 10.1674
R50373 a_50751_n19729.n495 a_50751_n19729.t342 10.1674
R50374 a_50751_n19729.n299 a_50751_n19729.t351 10.1674
R50375 a_50751_n19729.t351 a_50751_n19729.n298 10.1674
R50376 a_50751_n19729.n295 a_50751_n19729.t337 10.1674
R50377 a_50751_n19729.t337 a_50751_n19729.n294 10.1674
R50378 a_50751_n19729.n291 a_50751_n19729.t118 10.1674
R50379 a_50751_n19729.t118 a_50751_n19729.n290 10.1674
R50380 a_50751_n19729.t188 a_50751_n19729.n259 10.1674
R50381 a_50751_n19729.n260 a_50751_n19729.t188 10.1674
R50382 a_50751_n19729.t242 a_50751_n19729.n267 10.1674
R50383 a_50751_n19729.n268 a_50751_n19729.t242 10.1674
R50384 a_50751_n19729.n278 a_50751_n19729.t86 10.1674
R50385 a_50751_n19729.t86 a_50751_n19729.n277 10.1674
R50386 a_50751_n19729.n272 a_50751_n19729.t154 10.1674
R50387 a_50751_n19729.n249 a_50751_n19729.t149 10.1674
R50388 a_50751_n19729.t149 a_50751_n19729.n248 10.1674
R50389 a_50751_n19729.t210 a_50751_n19729.n504 10.1674
R50390 a_50751_n19729.n505 a_50751_n19729.t210 10.1674
R50391 a_50751_n19729.n306 a_50751_n19729.t80 10.1674
R50392 a_50751_n19729.t80 a_50751_n19729.n305 10.1674
R50393 a_50751_n19729.t148 a_50751_n19729.n311 10.1674
R50394 a_50751_n19729.n312 a_50751_n19729.t148 10.1674
R50395 a_50751_n19729.t136 a_50751_n19729.n315 10.1674
R50396 a_50751_n19729.n316 a_50751_n19729.t136 10.1674
R50397 a_50751_n19729.n328 a_50751_n19729.t209 10.1674
R50398 a_50751_n19729.t209 a_50751_n19729.n327 10.1674
R50399 a_50751_n19729.n320 a_50751_n19729.t361 10.1674
R50400 a_50751_n19729.t361 a_50751_n19729.n319 10.1674
R50401 a_50751_n19729.t126 a_50751_n19729.n340 10.1674
R50402 a_50751_n19729.n341 a_50751_n19729.t126 10.1674
R50403 a_50751_n19729.n345 a_50751_n19729.t181 10.1674
R50404 a_50751_n19729.n393 a_50751_n19729.t168 10.1674
R50405 a_50751_n19729.t168 a_50751_n19729.n392 10.1674
R50406 a_50751_n19729.n389 a_50751_n19729.t160 10.1674
R50407 a_50751_n19729.t160 a_50751_n19729.n388 10.1674
R50408 a_50751_n19729.n385 a_50751_n19729.t234 10.1674
R50409 a_50751_n19729.t234 a_50751_n19729.n384 10.1674
R50410 a_50751_n19729.t312 a_50751_n19729.n353 10.1674
R50411 a_50751_n19729.n354 a_50751_n19729.t312 10.1674
R50412 a_50751_n19729.t360 a_50751_n19729.n361 10.1674
R50413 a_50751_n19729.n362 a_50751_n19729.t360 10.1674
R50414 a_50751_n19729.n372 a_50751_n19729.t190 10.1674
R50415 a_50751_n19729.t190 a_50751_n19729.n371 10.1674
R50416 a_50751_n19729.n366 a_50751_n19729.t271 10.1674
R50417 a_50751_n19729.t285 a_50751_n19729.n323 10.1674
R50418 a_50751_n19729.n324 a_50751_n19729.t285 10.1674
R50419 a_50751_n19729.n337 a_50751_n19729.t344 10.1674
R50420 a_50751_n19729.t344 a_50751_n19729.n336 10.1674
R50421 a_50751_n19729.n358 a_50751_n19729.t301 10.1674
R50422 a_50751_n19729.t301 a_50751_n19729.n357 10.1674
R50423 a_50751_n19729.t139 a_50751_n19729.n375 10.1674
R50424 a_50751_n19729.n376 a_50751_n19729.t139 10.1674
R50425 a_50751_n19729.n401 a_50751_n19729.t215 10.1674
R50426 a_50751_n19729.t215 a_50751_n19729.n400 10.1674
R50427 a_50751_n19729.t289 a_50751_n19729.n406 10.1674
R50428 a_50751_n19729.n407 a_50751_n19729.t289 10.1674
R50429 a_50751_n19729.t280 a_50751_n19729.n410 10.1674
R50430 a_50751_n19729.n411 a_50751_n19729.t280 10.1674
R50431 a_50751_n19729.n423 a_50751_n19729.t350 10.1674
R50432 a_50751_n19729.t350 a_50751_n19729.n422 10.1674
R50433 a_50751_n19729.n415 a_50751_n19729.t202 10.1674
R50434 a_50751_n19729.t202 a_50751_n19729.n414 10.1674
R50435 a_50751_n19729.t269 a_50751_n19729.n435 10.1674
R50436 a_50751_n19729.n436 a_50751_n19729.t269 10.1674
R50437 a_50751_n19729.n440 a_50751_n19729.t329 10.1674
R50438 a_50751_n19729.n488 a_50751_n19729.t347 10.1674
R50439 a_50751_n19729.t347 a_50751_n19729.n487 10.1674
R50440 a_50751_n19729.n484 a_50751_n19729.t334 10.1674
R50441 a_50751_n19729.t334 a_50751_n19729.n483 10.1674
R50442 a_50751_n19729.n480 a_50751_n19729.t114 10.1674
R50443 a_50751_n19729.t114 a_50751_n19729.n479 10.1674
R50444 a_50751_n19729.t183 a_50751_n19729.n448 10.1674
R50445 a_50751_n19729.n449 a_50751_n19729.t183 10.1674
R50446 a_50751_n19729.t238 a_50751_n19729.n456 10.1674
R50447 a_50751_n19729.n457 a_50751_n19729.t238 10.1674
R50448 a_50751_n19729.n467 a_50751_n19729.t84 10.1674
R50449 a_50751_n19729.t84 a_50751_n19729.n466 10.1674
R50450 a_50751_n19729.n461 a_50751_n19729.t153 10.1674
R50451 a_50751_n19729.t130 a_50751_n19729.n418 10.1674
R50452 a_50751_n19729.n419 a_50751_n19729.t130 10.1674
R50453 a_50751_n19729.n432 a_50751_n19729.t187 10.1674
R50454 a_50751_n19729.t187 a_50751_n19729.n431 10.1674
R50455 a_50751_n19729.n453 a_50751_n19729.t174 10.1674
R50456 a_50751_n19729.t174 a_50751_n19729.n452 10.1674
R50457 a_50751_n19729.t317 a_50751_n19729.n470 10.1674
R50458 a_50751_n19729.n471 a_50751_n19729.t317 10.1674
R50459 a_50751_n19729.n264 a_50751_n19729.t177 10.1674
R50460 a_50751_n19729.t177 a_50751_n19729.n263 10.1674
R50461 a_50751_n19729.t321 a_50751_n19729.n281 10.1674
R50462 a_50751_n19729.n282 a_50751_n19729.t321 10.1674
R50463 a_50751_n19729.t170 a_50751_n19729.n492 10.1409
R50464 a_50751_n19729.t204 a_50751_n19729.n269 10.1409
R50465 a_50751_n19729.t254 a_50751_n19729.n342 10.1409
R50466 a_50751_n19729.t94 a_50751_n19729.n363 10.1409
R50467 a_50751_n19729.t82 a_50751_n19729.n437 10.1409
R50468 a_50751_n19729.t349 a_50751_n19729.n458 10.1409
R50469 a_50751_n19729.t342 a_50751_n19729.n494 10.1409
R50470 a_50751_n19729.t154 a_50751_n19729.n271 10.1409
R50471 a_50751_n19729.t181 a_50751_n19729.n344 10.1409
R50472 a_50751_n19729.t271 a_50751_n19729.n365 10.1409
R50473 a_50751_n19729.t329 a_50751_n19729.n439 10.1409
R50474 a_50751_n19729.t153 a_50751_n19729.n460 10.1409
R50475 a_50751_n19729.t267 a_50751_n19729.n492 9.54631
R50476 a_50751_n19729.n213 a_50751_n19729.t341 9.54631
R50477 a_50751_n19729.t171 a_50751_n19729.n212 9.54631
R50478 a_50751_n19729.n494 a_50751_n19729.t353 9.54631
R50479 a_50751_n19729.t105 a_50751_n19729.n269 9.54631
R50480 a_50751_n19729.n215 a_50751_n19729.t298 9.54631
R50481 a_50751_n19729.t75 a_50751_n19729.n214 9.54631
R50482 a_50751_n19729.n271 a_50751_n19729.t223 9.54631
R50483 a_50751_n19729.t92 a_50751_n19729.n342 9.54631
R50484 a_50751_n19729.n217 a_50751_n19729.t262 9.54631
R50485 a_50751_n19729.t256 a_50751_n19729.n216 9.54631
R50486 a_50751_n19729.n344 a_50751_n19729.t359 9.54631
R50487 a_50751_n19729.t156 a_50751_n19729.n363 9.54631
R50488 a_50751_n19729.n219 a_50751_n19729.t313 9.54631
R50489 a_50751_n19729.t246 a_50751_n19729.n218 9.54631
R50490 a_50751_n19729.n365 a_50751_n19729.t201 9.54631
R50491 a_50751_n19729.t101 a_50751_n19729.n437 9.54631
R50492 a_50751_n19729.n221 a_50751_n19729.t200 9.54631
R50493 a_50751_n19729.t299 a_50751_n19729.n220 9.54631
R50494 a_50751_n19729.n439 a_50751_n19729.t108 9.54631
R50495 a_50751_n19729.t157 a_50751_n19729.n458 9.54631
R50496 a_50751_n19729.n223 a_50751_n19729.t113 9.54631
R50497 a_50751_n19729.t314 a_50751_n19729.n222 9.54631
R50498 a_50751_n19729.n460 a_50751_n19729.t85 9.54631
R50499 a_50751_n19729.n233 a_50751_n19729.t152 9.54355
R50500 a_50751_n19729.t152 a_50751_n19729.n232 9.54355
R50501 a_50751_n19729.t227 a_50751_n19729.n2 9.54355
R50502 a_50751_n19729.n1 a_50751_n19729.t227 9.54355
R50503 a_50751_n19729.n229 a_50751_n19729.t358 9.54355
R50504 a_50751_n19729.n0 a_50751_n19729.t358 9.54355
R50505 a_50751_n19729.n230 a_50751_n19729.t237 9.54355
R50506 a_50751_n19729.n231 a_50751_n19729.t237 9.54355
R50507 a_50751_n19729.n235 a_50751_n19729.t224 9.54355
R50508 a_50751_n19729.t224 a_50751_n19729.n234 9.54355
R50509 a_50751_n19729.t307 a_50751_n19729.n7 9.54355
R50510 a_50751_n19729.n4 a_50751_n19729.t307 9.54355
R50511 a_50751_n19729.n5 a_50751_n19729.t138 9.54355
R50512 a_50751_n19729.t138 a_50751_n19729.n3 9.54355
R50513 a_50751_n19729.n237 a_50751_n19729.t315 9.54355
R50514 a_50751_n19729.n236 a_50751_n19729.t315 9.54355
R50515 a_50751_n19729.n239 a_50751_n19729.t216 9.54355
R50516 a_50751_n19729.t216 a_50751_n19729.n238 9.54355
R50517 a_50751_n19729.t294 a_50751_n19729.n11 9.54355
R50518 a_50751_n19729.n9 a_50751_n19729.t294 9.54355
R50519 a_50751_n19729.n10 a_50751_n19729.t123 9.54355
R50520 a_50751_n19729.t123 a_50751_n19729.n8 9.54355
R50521 a_50751_n19729.n241 a_50751_n19729.t303 9.54355
R50522 a_50751_n19729.n240 a_50751_n19729.t303 9.54355
R50523 a_50751_n19729.n243 a_50751_n19729.t290 9.54355
R50524 a_50751_n19729.t290 a_50751_n19729.n242 9.54355
R50525 a_50751_n19729.t70 a_50751_n19729.n15 9.54355
R50526 a_50751_n19729.n13 a_50751_n19729.t70 9.54355
R50527 a_50751_n19729.n14 a_50751_n19729.t40 9.54355
R50528 a_50751_n19729.t40 a_50751_n19729.n12 9.54355
R50529 a_50751_n19729.n245 a_50751_n19729.t88 9.54355
R50530 a_50751_n19729.n244 a_50751_n19729.t88 9.54355
R50531 a_50751_n19729.n251 a_50751_n19729.t145 9.54355
R50532 a_50751_n19729.t145 a_50751_n19729.n250 9.54355
R50533 a_50751_n19729.t36 a_50751_n19729.n20 9.54355
R50534 a_50751_n19729.n17 a_50751_n19729.t36 9.54355
R50535 a_50751_n19729.n18 a_50751_n19729.t8 9.54355
R50536 a_50751_n19729.t8 a_50751_n19729.n16 9.54355
R50537 a_50751_n19729.n253 a_50751_n19729.t228 9.54355
R50538 a_50751_n19729.n252 a_50751_n19729.t228 9.54355
R50539 a_50751_n19729.t205 a_50751_n19729.n498 9.54355
R50540 a_50751_n19729.n499 a_50751_n19729.t205 9.54355
R50541 a_50751_n19729.n25 a_50751_n19729.t284 9.54355
R50542 a_50751_n19729.t284 a_50751_n19729.n23 9.54355
R50543 a_50751_n19729.t112 a_50751_n19729.n24 9.54355
R50544 a_50751_n19729.n21 a_50751_n19729.t112 9.54355
R50545 a_50751_n19729.n500 a_50751_n19729.t295 9.54355
R50546 a_50751_n19729.n501 a_50751_n19729.t295 9.54355
R50547 a_50751_n19729.n493 a_50751_n19729.t267 9.54355
R50548 a_50751_n19729.t341 a_50751_n19729.n497 9.54355
R50549 a_50751_n19729.n496 a_50751_n19729.t171 9.54355
R50550 a_50751_n19729.n495 a_50751_n19729.t353 9.54355
R50551 a_50751_n19729.t305 a_50751_n19729.n296 9.54355
R50552 a_50751_n19729.n297 a_50751_n19729.t305 9.54355
R50553 a_50751_n19729.n30 a_50751_n19729.t192 9.54355
R50554 a_50751_n19729.t192 a_50751_n19729.n28 9.54355
R50555 a_50751_n19729.t266 a_50751_n19729.n29 9.54355
R50556 a_50751_n19729.n26 a_50751_n19729.t266 9.54355
R50557 a_50751_n19729.n298 a_50751_n19729.t124 9.54355
R50558 a_50751_n19729.n299 a_50751_n19729.t124 9.54355
R50559 a_50751_n19729.t292 a_50751_n19729.n292 9.54355
R50560 a_50751_n19729.n293 a_50751_n19729.t292 9.54355
R50561 a_50751_n19729.n34 a_50751_n19729.t180 9.54355
R50562 a_50751_n19729.t180 a_50751_n19729.n32 9.54355
R50563 a_50751_n19729.t253 a_50751_n19729.n33 9.54355
R50564 a_50751_n19729.n31 a_50751_n19729.t253 9.54355
R50565 a_50751_n19729.n294 a_50751_n19729.t109 9.54355
R50566 a_50751_n19729.n295 a_50751_n19729.t109 9.54355
R50567 a_50751_n19729.t78 a_50751_n19729.n288 9.54355
R50568 a_50751_n19729.n289 a_50751_n19729.t78 9.54355
R50569 a_50751_n19729.n39 a_50751_n19729.t260 9.54355
R50570 a_50751_n19729.t260 a_50751_n19729.n37 9.54355
R50571 a_50751_n19729.t327 a_50751_n19729.n38 9.54355
R50572 a_50751_n19729.n35 a_50751_n19729.t327 9.54355
R50573 a_50751_n19729.n290 a_50751_n19729.t182 9.54355
R50574 a_50751_n19729.n291 a_50751_n19729.t182 9.54355
R50575 a_50751_n19729.n258 a_50751_n19729.t146 9.54355
R50576 a_50751_n19729.t146 a_50751_n19729.n257 9.54355
R50577 a_50751_n19729.t14 a_50751_n19729.n43 9.54355
R50578 a_50751_n19729.n41 a_50751_n19729.t14 9.54355
R50579 a_50751_n19729.n42 a_50751_n19729.t56 9.54355
R50580 a_50751_n19729.t56 a_50751_n19729.n40 9.54355
R50581 a_50751_n19729.n260 a_50751_n19729.t263 9.54355
R50582 a_50751_n19729.n259 a_50751_n19729.t263 9.54355
R50583 a_50751_n19729.n266 a_50751_n19729.t185 9.54355
R50584 a_50751_n19729.t185 a_50751_n19729.n265 9.54355
R50585 a_50751_n19729.t66 a_50751_n19729.n48 9.54355
R50586 a_50751_n19729.n45 a_50751_n19729.t66 9.54355
R50587 a_50751_n19729.n46 a_50751_n19729.t46 9.54355
R50588 a_50751_n19729.t46 a_50751_n19729.n44 9.54355
R50589 a_50751_n19729.n268 a_50751_n19729.t311 9.54355
R50590 a_50751_n19729.n267 a_50751_n19729.t311 9.54355
R50591 a_50751_n19729.t326 a_50751_n19729.n275 9.54355
R50592 a_50751_n19729.n276 a_50751_n19729.t326 9.54355
R50593 a_50751_n19729.n53 a_50751_n19729.t219 9.54355
R50594 a_50751_n19729.t219 a_50751_n19729.n51 9.54355
R50595 a_50751_n19729.t288 a_50751_n19729.n52 9.54355
R50596 a_50751_n19729.n49 a_50751_n19729.t288 9.54355
R50597 a_50751_n19729.n277 a_50751_n19729.t150 9.54355
R50598 a_50751_n19729.n278 a_50751_n19729.t150 9.54355
R50599 a_50751_n19729.n270 a_50751_n19729.t105 9.54355
R50600 a_50751_n19729.t298 a_50751_n19729.n274 9.54355
R50601 a_50751_n19729.n273 a_50751_n19729.t75 9.54355
R50602 a_50751_n19729.n272 a_50751_n19729.t223 9.54355
R50603 a_50751_n19729.t76 a_50751_n19729.n246 9.54355
R50604 a_50751_n19729.n247 a_50751_n19729.t76 9.54355
R50605 a_50751_n19729.n57 a_50751_n19729.t48 9.54355
R50606 a_50751_n19729.t48 a_50751_n19729.n55 9.54355
R50607 a_50751_n19729.t30 a_50751_n19729.n56 9.54355
R50608 a_50751_n19729.n54 a_50751_n19729.t30 9.54355
R50609 a_50751_n19729.n248 a_50751_n19729.t155 9.54355
R50610 a_50751_n19729.n249 a_50751_n19729.t155 9.54355
R50611 a_50751_n19729.n503 a_50751_n19729.t133 9.54355
R50612 a_50751_n19729.t133 a_50751_n19729.n502 9.54355
R50613 a_50751_n19729.t208 a_50751_n19729.n61 9.54355
R50614 a_50751_n19729.n59 a_50751_n19729.t208 9.54355
R50615 a_50751_n19729.n60 a_50751_n19729.t332 9.54355
R50616 a_50751_n19729.t332 a_50751_n19729.n58 9.54355
R50617 a_50751_n19729.n505 a_50751_n19729.t217 9.54355
R50618 a_50751_n19729.n504 a_50751_n19729.t217 9.54355
R50619 a_50751_n19729.n308 a_50751_n19729.t265 9.54355
R50620 a_50751_n19729.t265 a_50751_n19729.n307 9.54355
R50621 a_50751_n19729.t147 a_50751_n19729.n64 9.54355
R50622 a_50751_n19729.n63 a_50751_n19729.t147 9.54355
R50623 a_50751_n19729.n304 a_50751_n19729.t141 9.54355
R50624 a_50751_n19729.n62 a_50751_n19729.t141 9.54355
R50625 a_50751_n19729.n305 a_50751_n19729.t241 9.54355
R50626 a_50751_n19729.n306 a_50751_n19729.t241 9.54355
R50627 a_50751_n19729.n310 a_50751_n19729.t336 9.54355
R50628 a_50751_n19729.t336 a_50751_n19729.n309 9.54355
R50629 a_50751_n19729.t220 a_50751_n19729.n69 9.54355
R50630 a_50751_n19729.n66 a_50751_n19729.t220 9.54355
R50631 a_50751_n19729.n67 a_50751_n19729.t214 9.54355
R50632 a_50751_n19729.t214 a_50751_n19729.n65 9.54355
R50633 a_50751_n19729.n312 a_50751_n19729.t320 9.54355
R50634 a_50751_n19729.n311 a_50751_n19729.t320 9.54355
R50635 a_50751_n19729.n314 a_50751_n19729.t325 9.54355
R50636 a_50751_n19729.t325 a_50751_n19729.n313 9.54355
R50637 a_50751_n19729.t207 a_50751_n19729.n73 9.54355
R50638 a_50751_n19729.n71 a_50751_n19729.t207 9.54355
R50639 a_50751_n19729.n72 a_50751_n19729.t199 9.54355
R50640 a_50751_n19729.t199 a_50751_n19729.n70 9.54355
R50641 a_50751_n19729.n316 a_50751_n19729.t306 9.54355
R50642 a_50751_n19729.n315 a_50751_n19729.t306 9.54355
R50643 a_50751_n19729.t104 a_50751_n19729.n325 9.54355
R50644 a_50751_n19729.n326 a_50751_n19729.t104 9.54355
R50645 a_50751_n19729.n78 a_50751_n19729.t24 9.54355
R50646 a_50751_n19729.t24 a_50751_n19729.n76 9.54355
R50647 a_50751_n19729.t28 a_50751_n19729.n77 9.54355
R50648 a_50751_n19729.n74 a_50751_n19729.t28 9.54355
R50649 a_50751_n19729.n327 a_50751_n19729.t93 9.54355
R50650 a_50751_n19729.n328 a_50751_n19729.t93 9.54355
R50651 a_50751_n19729.t259 a_50751_n19729.n317 9.54355
R50652 a_50751_n19729.n318 a_50751_n19729.t259 9.54355
R50653 a_50751_n19729.n83 a_50751_n19729.t52 9.54355
R50654 a_50751_n19729.t52 a_50751_n19729.n81 9.54355
R50655 a_50751_n19729.t54 a_50751_n19729.n82 9.54355
R50656 a_50751_n19729.n79 a_50751_n19729.t54 9.54355
R50657 a_50751_n19729.n319 a_50751_n19729.t232 9.54355
R50658 a_50751_n19729.n320 a_50751_n19729.t232 9.54355
R50659 a_50751_n19729.n339 a_50751_n19729.t323 9.54355
R50660 a_50751_n19729.t323 a_50751_n19729.n338 9.54355
R50661 a_50751_n19729.t198 a_50751_n19729.n88 9.54355
R50662 a_50751_n19729.n85 a_50751_n19729.t198 9.54355
R50663 a_50751_n19729.n86 a_50751_n19729.t186 9.54355
R50664 a_50751_n19729.t186 a_50751_n19729.n84 9.54355
R50665 a_50751_n19729.n341 a_50751_n19729.t300 9.54355
R50666 a_50751_n19729.n340 a_50751_n19729.t300 9.54355
R50667 a_50751_n19729.n343 a_50751_n19729.t92 9.54355
R50668 a_50751_n19729.t262 a_50751_n19729.n347 9.54355
R50669 a_50751_n19729.n346 a_50751_n19729.t256 9.54355
R50670 a_50751_n19729.n345 a_50751_n19729.t359 9.54355
R50671 a_50751_n19729.t352 a_50751_n19729.n390 9.54355
R50672 a_50751_n19729.n391 a_50751_n19729.t352 9.54355
R50673 a_50751_n19729.n93 a_50751_n19729.t211 9.54355
R50674 a_50751_n19729.t211 a_50751_n19729.n91 9.54355
R50675 a_50751_n19729.t144 a_50751_n19729.n92 9.54355
R50676 a_50751_n19729.n89 a_50751_n19729.t144 9.54355
R50677 a_50751_n19729.n392 a_50751_n19729.t102 9.54355
R50678 a_50751_n19729.n393 a_50751_n19729.t102 9.54355
R50679 a_50751_n19729.t338 a_50751_n19729.n386 9.54355
R50680 a_50751_n19729.n387 a_50751_n19729.t338 9.54355
R50681 a_50751_n19729.n97 a_50751_n19729.t195 9.54355
R50682 a_50751_n19729.t195 a_50751_n19729.n95 9.54355
R50683 a_50751_n19729.t131 a_50751_n19729.n96 9.54355
R50684 a_50751_n19729.n94 a_50751_n19729.t131 9.54355
R50685 a_50751_n19729.n388 a_50751_n19729.t97 9.54355
R50686 a_50751_n19729.n389 a_50751_n19729.t97 9.54355
R50687 a_50751_n19729.t119 a_50751_n19729.n382 9.54355
R50688 a_50751_n19729.n383 a_50751_n19729.t119 9.54355
R50689 a_50751_n19729.n102 a_50751_n19729.t275 9.54355
R50690 a_50751_n19729.t275 a_50751_n19729.n100 9.54355
R50691 a_50751_n19729.t203 a_50751_n19729.n101 9.54355
R50692 a_50751_n19729.n98 a_50751_n19729.t203 9.54355
R50693 a_50751_n19729.n384 a_50751_n19729.t164 9.54355
R50694 a_50751_n19729.n385 a_50751_n19729.t164 9.54355
R50695 a_50751_n19729.n352 a_50751_n19729.t189 9.54355
R50696 a_50751_n19729.t189 a_50751_n19729.n351 9.54355
R50697 a_50751_n19729.t6 a_50751_n19729.n106 9.54355
R50698 a_50751_n19729.n104 a_50751_n19729.t6 9.54355
R50699 a_50751_n19729.n105 a_50751_n19729.t26 9.54355
R50700 a_50751_n19729.t26 a_50751_n19729.n103 9.54355
R50701 a_50751_n19729.n354 a_50751_n19729.t244 9.54355
R50702 a_50751_n19729.n353 a_50751_n19729.t244 9.54355
R50703 a_50751_n19729.n360 a_50751_n19729.t243 9.54355
R50704 a_50751_n19729.t243 a_50751_n19729.n359 9.54355
R50705 a_50751_n19729.t60 a_50751_n19729.n111 9.54355
R50706 a_50751_n19729.n108 a_50751_n19729.t60 9.54355
R50707 a_50751_n19729.n109 a_50751_n19729.t16 9.54355
R50708 a_50751_n19729.t16 a_50751_n19729.n107 9.54355
R50709 a_50751_n19729.n362 a_50751_n19729.t291 9.54355
R50710 a_50751_n19729.n361 a_50751_n19729.t291 9.54355
R50711 a_50751_n19729.t87 a_50751_n19729.n369 9.54355
R50712 a_50751_n19729.n370 a_50751_n19729.t87 9.54355
R50713 a_50751_n19729.n116 a_50751_n19729.t235 9.54355
R50714 a_50751_n19729.t235 a_50751_n19729.n114 9.54355
R50715 a_50751_n19729.t165 a_50751_n19729.n115 9.54355
R50716 a_50751_n19729.n112 a_50751_n19729.t165 9.54355
R50717 a_50751_n19729.n371 a_50751_n19729.t128 9.54355
R50718 a_50751_n19729.n372 a_50751_n19729.t128 9.54355
R50719 a_50751_n19729.n364 a_50751_n19729.t156 9.54355
R50720 a_50751_n19729.t313 a_50751_n19729.n368 9.54355
R50721 a_50751_n19729.n367 a_50751_n19729.t246 9.54355
R50722 a_50751_n19729.n366 a_50751_n19729.t201 9.54355
R50723 a_50751_n19729.n322 a_50751_n19729.t176 9.54355
R50724 a_50751_n19729.t176 a_50751_n19729.n321 9.54355
R50725 a_50751_n19729.t0 a_50751_n19729.n120 9.54355
R50726 a_50751_n19729.n118 a_50751_n19729.t0 9.54355
R50727 a_50751_n19729.n119 a_50751_n19729.t2 9.54355
R50728 a_50751_n19729.t2 a_50751_n19729.n117 9.54355
R50729 a_50751_n19729.n324 a_50751_n19729.t158 9.54355
R50730 a_50751_n19729.n323 a_50751_n19729.t158 9.54355
R50731 a_50751_n19729.t247 a_50751_n19729.n334 9.54355
R50732 a_50751_n19729.n335 a_50751_n19729.t247 9.54355
R50733 a_50751_n19729.n124 a_50751_n19729.t125 9.54355
R50734 a_50751_n19729.t125 a_50751_n19729.n122 9.54355
R50735 a_50751_n19729.t116 a_50751_n19729.n123 9.54355
R50736 a_50751_n19729.n121 a_50751_n19729.t116 9.54355
R50737 a_50751_n19729.n336 a_50751_n19729.t221 9.54355
R50738 a_50751_n19729.n337 a_50751_n19729.t221 9.54355
R50739 a_50751_n19729.t178 a_50751_n19729.n355 9.54355
R50740 a_50751_n19729.n356 a_50751_n19729.t178 9.54355
R50741 a_50751_n19729.n128 a_50751_n19729.t12 9.54355
R50742 a_50751_n19729.t12 a_50751_n19729.n126 9.54355
R50743 a_50751_n19729.t32 a_50751_n19729.n127 9.54355
R50744 a_50751_n19729.n125 a_50751_n19729.t32 9.54355
R50745 a_50751_n19729.n357 a_50751_n19729.t226 9.54355
R50746 a_50751_n19729.n358 a_50751_n19729.t226 9.54355
R50747 a_50751_n19729.n374 a_50751_n19729.t322 9.54355
R50748 a_50751_n19729.t322 a_50751_n19729.n373 9.54355
R50749 a_50751_n19729.t172 a_50751_n19729.n132 9.54355
R50750 a_50751_n19729.n130 a_50751_n19729.t172 9.54355
R50751 a_50751_n19729.n131 a_50751_n19729.t107 9.54355
R50752 a_50751_n19729.t107 a_50751_n19729.n129 9.54355
R50753 a_50751_n19729.n376 a_50751_n19729.t77 9.54355
R50754 a_50751_n19729.n375 a_50751_n19729.t77 9.54355
R50755 a_50751_n19729.n403 a_50751_n19729.t282 9.54355
R50756 a_50751_n19729.t282 a_50751_n19729.n402 9.54355
R50757 a_50751_n19729.t95 a_50751_n19729.n135 9.54355
R50758 a_50751_n19729.n134 a_50751_n19729.t95 9.54355
R50759 a_50751_n19729.n399 a_50751_n19729.t175 9.54355
R50760 a_50751_n19729.n133 a_50751_n19729.t175 9.54355
R50761 a_50751_n19729.n400 a_50751_n19729.t293 9.54355
R50762 a_50751_n19729.n401 a_50751_n19729.t293 9.54355
R50763 a_50751_n19729.n405 a_50751_n19729.t356 9.54355
R50764 a_50751_n19729.t356 a_50751_n19729.n404 9.54355
R50765 a_50751_n19729.t162 a_50751_n19729.n140 9.54355
R50766 a_50751_n19729.n137 a_50751_n19729.t162 9.54355
R50767 a_50751_n19729.n138 a_50751_n19729.t258 9.54355
R50768 a_50751_n19729.t258 a_50751_n19729.n136 9.54355
R50769 a_50751_n19729.n407 a_50751_n19729.t79 9.54355
R50770 a_50751_n19729.n406 a_50751_n19729.t79 9.54355
R50771 a_50751_n19729.n409 a_50751_n19729.t340 9.54355
R50772 a_50751_n19729.t340 a_50751_n19729.n408 9.54355
R50773 a_50751_n19729.t151 a_50751_n19729.n144 9.54355
R50774 a_50751_n19729.n142 a_50751_n19729.t151 9.54355
R50775 a_50751_n19729.n143 a_50751_n19729.t245 9.54355
R50776 a_50751_n19729.t245 a_50751_n19729.n141 9.54355
R50777 a_50751_n19729.n411 a_50751_n19729.t354 9.54355
R50778 a_50751_n19729.n410 a_50751_n19729.t354 9.54355
R50779 a_50751_n19729.t121 a_50751_n19729.n420 9.54355
R50780 a_50751_n19729.n421 a_50751_n19729.t121 9.54355
R50781 a_50751_n19729.n149 a_50751_n19729.t34 9.54355
R50782 a_50751_n19729.t34 a_50751_n19729.n147 9.54355
R50783 a_50751_n19729.t20 a_50751_n19729.n148 9.54355
R50784 a_50751_n19729.n145 a_50751_n19729.t20 9.54355
R50785 a_50751_n19729.n422 a_50751_n19729.t135 9.54355
R50786 a_50751_n19729.n423 a_50751_n19729.t135 9.54355
R50787 a_50751_n19729.t273 a_50751_n19729.n412 9.54355
R50788 a_50751_n19729.n413 a_50751_n19729.t273 9.54355
R50789 a_50751_n19729.n154 a_50751_n19729.t68 9.54355
R50790 a_50751_n19729.t68 a_50751_n19729.n152 9.54355
R50791 a_50751_n19729.t42 a_50751_n19729.n153 9.54355
R50792 a_50751_n19729.n150 a_50751_n19729.t42 9.54355
R50793 a_50751_n19729.n414 a_50751_n19729.t283 9.54355
R50794 a_50751_n19729.n415 a_50751_n19729.t283 9.54355
R50795 a_50751_n19729.n434 a_50751_n19729.t330 9.54355
R50796 a_50751_n19729.t330 a_50751_n19729.n433 9.54355
R50797 a_50751_n19729.t142 a_50751_n19729.n159 9.54355
R50798 a_50751_n19729.n156 a_50751_n19729.t142 9.54355
R50799 a_50751_n19729.n157 a_50751_n19729.t233 9.54355
R50800 a_50751_n19729.t233 a_50751_n19729.n155 9.54355
R50801 a_50751_n19729.n436 a_50751_n19729.t343 9.54355
R50802 a_50751_n19729.n435 a_50751_n19729.t343 9.54355
R50803 a_50751_n19729.n438 a_50751_n19729.t101 9.54355
R50804 a_50751_n19729.t200 a_50751_n19729.n442 9.54355
R50805 a_50751_n19729.n441 a_50751_n19729.t299 9.54355
R50806 a_50751_n19729.n440 a_50751_n19729.t108 9.54355
R50807 a_50751_n19729.t355 a_50751_n19729.n485 9.54355
R50808 a_50751_n19729.n486 a_50751_n19729.t355 9.54355
R50809 a_50751_n19729.n164 a_50751_n19729.t316 9.54355
R50810 a_50751_n19729.t316 a_50751_n19729.n162 9.54355
R50811 a_50751_n19729.t213 a_50751_n19729.n163 9.54355
R50812 a_50751_n19729.n160 a_50751_n19729.t213 9.54355
R50813 a_50751_n19729.n487 a_50751_n19729.t278 9.54355
R50814 a_50751_n19729.n488 a_50751_n19729.t278 9.54355
R50815 a_50751_n19729.t339 a_50751_n19729.n481 9.54355
R50816 a_50751_n19729.n482 a_50751_n19729.t339 9.54355
R50817 a_50751_n19729.n168 a_50751_n19729.t304 9.54355
R50818 a_50751_n19729.t304 a_50751_n19729.n166 9.54355
R50819 a_50751_n19729.t197 a_50751_n19729.n167 9.54355
R50820 a_50751_n19729.n165 a_50751_n19729.t197 9.54355
R50821 a_50751_n19729.n483 a_50751_n19729.t264 9.54355
R50822 a_50751_n19729.n484 a_50751_n19729.t264 9.54355
R50823 a_50751_n19729.t120 a_50751_n19729.n477 9.54355
R50824 a_50751_n19729.n478 a_50751_n19729.t120 9.54355
R50825 a_50751_n19729.n173 a_50751_n19729.t89 9.54355
R50826 a_50751_n19729.t89 a_50751_n19729.n171 9.54355
R50827 a_50751_n19729.t277 a_50751_n19729.n172 9.54355
R50828 a_50751_n19729.n169 a_50751_n19729.t277 9.54355
R50829 a_50751_n19729.n479 a_50751_n19729.t335 9.54355
R50830 a_50751_n19729.n480 a_50751_n19729.t335 9.54355
R50831 a_50751_n19729.n447 a_50751_n19729.t191 9.54355
R50832 a_50751_n19729.t191 a_50751_n19729.n446 9.54355
R50833 a_50751_n19729.t44 a_50751_n19729.n177 9.54355
R50834 a_50751_n19729.n175 a_50751_n19729.t44 9.54355
R50835 a_50751_n19729.n176 a_50751_n19729.t4 9.54355
R50836 a_50751_n19729.t4 a_50751_n19729.n174 9.54355
R50837 a_50751_n19729.n449 a_50751_n19729.t117 9.54355
R50838 a_50751_n19729.n448 a_50751_n19729.t117 9.54355
R50839 a_50751_n19729.n455 a_50751_n19729.t248 9.54355
R50840 a_50751_n19729.t248 a_50751_n19729.n454 9.54355
R50841 a_50751_n19729.t38 a_50751_n19729.n182 9.54355
R50842 a_50751_n19729.n179 a_50751_n19729.t38 9.54355
R50843 a_50751_n19729.n180 a_50751_n19729.t58 9.54355
R50844 a_50751_n19729.t58 a_50751_n19729.n178 9.54355
R50845 a_50751_n19729.n457 a_50751_n19729.t163 9.54355
R50846 a_50751_n19729.n456 a_50751_n19729.t163 9.54355
R50847 a_50751_n19729.t90 a_50751_n19729.n464 9.54355
R50848 a_50751_n19729.n465 a_50751_n19729.t90 9.54355
R50849 a_50751_n19729.n187 a_50751_n19729.t333 9.54355
R50850 a_50751_n19729.t333 a_50751_n19729.n185 9.54355
R50851 a_50751_n19729.t236 a_50751_n19729.n186 9.54355
R50852 a_50751_n19729.n183 a_50751_n19729.t236 9.54355
R50853 a_50751_n19729.n466 a_50751_n19729.t302 9.54355
R50854 a_50751_n19729.n467 a_50751_n19729.t302 9.54355
R50855 a_50751_n19729.n459 a_50751_n19729.t157 9.54355
R50856 a_50751_n19729.t113 a_50751_n19729.n463 9.54355
R50857 a_50751_n19729.n462 a_50751_n19729.t314 9.54355
R50858 a_50751_n19729.n461 a_50751_n19729.t85 9.54355
R50859 a_50751_n19729.n417 a_50751_n19729.t193 9.54355
R50860 a_50751_n19729.t193 a_50751_n19729.n416 9.54355
R50861 a_50751_n19729.t22 a_50751_n19729.n191 9.54355
R50862 a_50751_n19729.n189 a_50751_n19729.t22 9.54355
R50863 a_50751_n19729.n190 a_50751_n19729.t62 9.54355
R50864 a_50751_n19729.t62 a_50751_n19729.n188 9.54355
R50865 a_50751_n19729.n419 a_50751_n19729.t206 9.54355
R50866 a_50751_n19729.n418 a_50751_n19729.t206 9.54355
R50867 a_50751_n19729.t261 a_50751_n19729.n429 9.54355
R50868 a_50751_n19729.n430 a_50751_n19729.t261 9.54355
R50869 a_50751_n19729.n195 a_50751_n19729.t74 9.54355
R50870 a_50751_n19729.t74 a_50751_n19729.n193 9.54355
R50871 a_50751_n19729.t159 a_50751_n19729.n194 9.54355
R50872 a_50751_n19729.n192 a_50751_n19729.t159 9.54355
R50873 a_50751_n19729.n431 a_50751_n19729.t270 9.54355
R50874 a_50751_n19729.n432 a_50751_n19729.t270 9.54355
R50875 a_50751_n19729.t179 a_50751_n19729.n450 9.54355
R50876 a_50751_n19729.n451 a_50751_n19729.t179 9.54355
R50877 a_50751_n19729.n199 a_50751_n19729.t50 9.54355
R50878 a_50751_n19729.t50 a_50751_n19729.n197 9.54355
R50879 a_50751_n19729.t10 a_50751_n19729.n198 9.54355
R50880 a_50751_n19729.n196 a_50751_n19729.t10 9.54355
R50881 a_50751_n19729.n452 a_50751_n19729.t103 9.54355
R50882 a_50751_n19729.n453 a_50751_n19729.t103 9.54355
R50883 a_50751_n19729.n469 a_50751_n19729.t324 9.54355
R50884 a_50751_n19729.t324 a_50751_n19729.n468 9.54355
R50885 a_50751_n19729.t281 a_50751_n19729.n203 9.54355
R50886 a_50751_n19729.n201 a_50751_n19729.t281 9.54355
R50887 a_50751_n19729.n202 a_50751_n19729.t173 9.54355
R50888 a_50751_n19729.t173 a_50751_n19729.n200 9.54355
R50889 a_50751_n19729.n471 a_50751_n19729.t240 9.54355
R50890 a_50751_n19729.n470 a_50751_n19729.t240 9.54355
R50891 a_50751_n19729.t134 a_50751_n19729.n261 9.54355
R50892 a_50751_n19729.n262 a_50751_n19729.t134 9.54355
R50893 a_50751_n19729.n207 a_50751_n19729.t18 9.54355
R50894 a_50751_n19729.t18 a_50751_n19729.n205 9.54355
R50895 a_50751_n19729.t64 a_50751_n19729.n206 9.54355
R50896 a_50751_n19729.n204 a_50751_n19729.t64 9.54355
R50897 a_50751_n19729.n263 a_50751_n19729.t251 9.54355
R50898 a_50751_n19729.n264 a_50751_n19729.t251 9.54355
R50899 a_50751_n19729.n280 a_50751_n19729.t268 9.54355
R50900 a_50751_n19729.t268 a_50751_n19729.n279 9.54355
R50901 a_50751_n19729.t161 a_50751_n19729.n211 9.54355
R50902 a_50751_n19729.n209 a_50751_n19729.t161 9.54355
R50903 a_50751_n19729.n210 a_50751_n19729.t225 9.54355
R50904 a_50751_n19729.t225 a_50751_n19729.n208 9.54355
R50905 a_50751_n19729.n282 a_50751_n19729.t96 9.54355
R50906 a_50751_n19729.n281 a_50751_n19729.t96 9.54355
R50907 a_50751_n19729.n300 a_50751_n19729.t73 7.11376
R50908 a_50751_n19729.n395 a_50751_n19729.n300 6.02769
R50909 a_50751_n19729.n491 a_50751_n19729.n490 3.90251
R50910 a_50751_n19729.n508 a_50751_n19729.t49 3.3605
R50911 a_50751_n19729.n507 a_50751_n19729.t37 3.3605
R50912 a_50751_n19729.n226 a_50751_n19729.t41 3.3605
R50913 a_50751_n19729.n227 a_50751_n19729.t31 3.3605
R50914 a_50751_n19729.n228 a_50751_n19729.t9 3.3605
R50915 a_50751_n19729.n303 a_50751_n19729.t29 3.3605
R50916 a_50751_n19729.n302 a_50751_n19729.t3 3.3605
R50917 a_50751_n19729.n301 a_50751_n19729.t55 3.3605
R50918 a_50751_n19729.n330 a_50751_n19729.t25 3.3605
R50919 a_50751_n19729.n331 a_50751_n19729.t1 3.3605
R50920 a_50751_n19729.n332 a_50751_n19729.t53 3.3605
R50921 a_50751_n19729.n348 a_50751_n19729.t27 3.3605
R50922 a_50751_n19729.n349 a_50751_n19729.t33 3.3605
R50923 a_50751_n19729.n350 a_50751_n19729.t17 3.3605
R50924 a_50751_n19729.n380 a_50751_n19729.t7 3.3605
R50925 a_50751_n19729.n379 a_50751_n19729.t13 3.3605
R50926 a_50751_n19729.n378 a_50751_n19729.t61 3.3605
R50927 a_50751_n19729.n398 a_50751_n19729.t21 3.3605
R50928 a_50751_n19729.n397 a_50751_n19729.t63 3.3605
R50929 a_50751_n19729.n396 a_50751_n19729.t43 3.3605
R50930 a_50751_n19729.n425 a_50751_n19729.t35 3.3605
R50931 a_50751_n19729.n426 a_50751_n19729.t23 3.3605
R50932 a_50751_n19729.n427 a_50751_n19729.t69 3.3605
R50933 a_50751_n19729.n443 a_50751_n19729.t5 3.3605
R50934 a_50751_n19729.n444 a_50751_n19729.t11 3.3605
R50935 a_50751_n19729.n445 a_50751_n19729.t59 3.3605
R50936 a_50751_n19729.n475 a_50751_n19729.t45 3.3605
R50937 a_50751_n19729.n474 a_50751_n19729.t51 3.3605
R50938 a_50751_n19729.n473 a_50751_n19729.t39 3.3605
R50939 a_50751_n19729.n254 a_50751_n19729.t57 3.3605
R50940 a_50751_n19729.n255 a_50751_n19729.t65 3.3605
R50941 a_50751_n19729.n256 a_50751_n19729.t47 3.3605
R50942 a_50751_n19729.n286 a_50751_n19729.t15 3.3605
R50943 a_50751_n19729.n285 a_50751_n19729.t19 3.3605
R50944 a_50751_n19729.n284 a_50751_n19729.t67 3.3605
R50945 a_50751_n19729.t71 a_50751_n19729.n509 3.3605
R50946 a_50751_n19729.n490 a_50751_n19729.n395 3.14899
R50947 a_50751_n19729.n333 a_50751_n19729.n301 2.59662
R50948 a_50751_n19729.n377 a_50751_n19729.n350 2.59662
R50949 a_50751_n19729.n428 a_50751_n19729.n396 2.59662
R50950 a_50751_n19729.n472 a_50751_n19729.n445 2.59662
R50951 a_50751_n19729.n283 a_50751_n19729.n256 2.59662
R50952 a_50751_n19729.n506 a_50751_n19729.n228 2.59662
R50953 a_50751_n19729.n226 a_50751_n19729.n225 2.59544
R50954 a_50751_n19729.n329 a_50751_n19729.n303 2.59544
R50955 a_50751_n19729.n381 a_50751_n19729.n348 2.59544
R50956 a_50751_n19729.n424 a_50751_n19729.n398 2.59544
R50957 a_50751_n19729.n476 a_50751_n19729.n443 2.59544
R50958 a_50751_n19729.n287 a_50751_n19729.n254 2.59544
R50959 a_50751_n19729.n333 a_50751_n19729.n332 2.58354
R50960 a_50751_n19729.n378 a_50751_n19729.n377 2.58354
R50961 a_50751_n19729.n428 a_50751_n19729.n427 2.58354
R50962 a_50751_n19729.n473 a_50751_n19729.n472 2.58354
R50963 a_50751_n19729.n284 a_50751_n19729.n283 2.58354
R50964 a_50751_n19729.n507 a_50751_n19729.n506 2.58354
R50965 a_50751_n19729.n509 a_50751_n19729.n225 2.58235
R50966 a_50751_n19729.n330 a_50751_n19729.n329 2.58235
R50967 a_50751_n19729.n381 a_50751_n19729.n380 2.58235
R50968 a_50751_n19729.n425 a_50751_n19729.n424 2.58235
R50969 a_50751_n19729.n476 a_50751_n19729.n475 2.58235
R50970 a_50751_n19729.n287 a_50751_n19729.n286 2.58235
R50971 a_50751_n19729.n68 a_50751_n19729.n64 1.6805
R50972 a_50751_n19729.n139 a_50751_n19729.n135 1.6805
R50973 a_50751_n19729.n6 a_50751_n19729.n2 1.6805
R50974 a_50751_n19729.n113 a_50751_n19729.n219 1.59324
R50975 a_50751_n19729.n184 a_50751_n19729.n223 1.59324
R50976 a_50751_n19729.n50 a_50751_n19729.n215 1.59324
R50977 a_50751_n19729.n132 a_50751_n19729.n113 1.5005
R50978 a_50751_n19729.n377 a_50751_n19729.n113 1.5005
R50979 a_50751_n19729.n110 a_50751_n19729.n128 1.5005
R50980 a_50751_n19729.n99 a_50751_n19729.n381 1.5005
R50981 a_50751_n19729.n87 a_50751_n19729.n124 1.5005
R50982 a_50751_n19729.n80 a_50751_n19729.n333 1.5005
R50983 a_50751_n19729.n120 a_50751_n19729.n75 1.5005
R50984 a_50751_n19729.n329 a_50751_n19729.n68 1.5005
R50985 a_50751_n19729.n113 a_50751_n19729.n116 1.5005
R50986 a_50751_n19729.n114 a_50751_n19729.n113 1.5005
R50987 a_50751_n19729.n113 a_50751_n19729.n130 1.5005
R50988 a_50751_n19729.n111 a_50751_n19729.n110 1.5005
R50989 a_50751_n19729.n113 a_50751_n19729.n108 1.5005
R50990 a_50751_n19729.n126 a_50751_n19729.n110 1.5005
R50991 a_50751_n19729.n106 a_50751_n19729.n99 1.5005
R50992 a_50751_n19729.n110 a_50751_n19729.n104 1.5005
R50993 a_50751_n19729.n90 a_50751_n19729.n102 1.5005
R50994 a_50751_n19729.n100 a_50751_n19729.n99 1.5005
R50995 a_50751_n19729.n90 a_50751_n19729.n97 1.5005
R50996 a_50751_n19729.n95 a_50751_n19729.n90 1.5005
R50997 a_50751_n19729.n90 a_50751_n19729.n93 1.5005
R50998 a_50751_n19729.n91 a_50751_n19729.n90 1.5005
R50999 a_50751_n19729.n87 a_50751_n19729.n217 1.5005
R51000 a_50751_n19729.n88 a_50751_n19729.n87 1.5005
R51001 a_50751_n19729.n87 a_50751_n19729.n85 1.5005
R51002 a_50751_n19729.n122 a_50751_n19729.n80 1.5005
R51003 a_50751_n19729.n75 a_50751_n19729.n83 1.5005
R51004 a_50751_n19729.n81 a_50751_n19729.n80 1.5005
R51005 a_50751_n19729.n75 a_50751_n19729.n118 1.5005
R51006 a_50751_n19729.n68 a_50751_n19729.n78 1.5005
R51007 a_50751_n19729.n76 a_50751_n19729.n75 1.5005
R51008 a_50751_n19729.n73 a_50751_n19729.n68 1.5005
R51009 a_50751_n19729.n68 a_50751_n19729.n71 1.5005
R51010 a_50751_n19729.n69 a_50751_n19729.n68 1.5005
R51011 a_50751_n19729.n68 a_50751_n19729.n66 1.5005
R51012 a_50751_n19729.n68 a_50751_n19729.n63 1.5005
R51013 a_50751_n19729.n203 a_50751_n19729.n184 1.5005
R51014 a_50751_n19729.n472 a_50751_n19729.n184 1.5005
R51015 a_50751_n19729.n181 a_50751_n19729.n199 1.5005
R51016 a_50751_n19729.n170 a_50751_n19729.n476 1.5005
R51017 a_50751_n19729.n158 a_50751_n19729.n195 1.5005
R51018 a_50751_n19729.n151 a_50751_n19729.n428 1.5005
R51019 a_50751_n19729.n191 a_50751_n19729.n146 1.5005
R51020 a_50751_n19729.n424 a_50751_n19729.n139 1.5005
R51021 a_50751_n19729.n184 a_50751_n19729.n187 1.5005
R51022 a_50751_n19729.n185 a_50751_n19729.n184 1.5005
R51023 a_50751_n19729.n184 a_50751_n19729.n201 1.5005
R51024 a_50751_n19729.n182 a_50751_n19729.n181 1.5005
R51025 a_50751_n19729.n184 a_50751_n19729.n179 1.5005
R51026 a_50751_n19729.n197 a_50751_n19729.n181 1.5005
R51027 a_50751_n19729.n177 a_50751_n19729.n170 1.5005
R51028 a_50751_n19729.n181 a_50751_n19729.n175 1.5005
R51029 a_50751_n19729.n161 a_50751_n19729.n173 1.5005
R51030 a_50751_n19729.n171 a_50751_n19729.n170 1.5005
R51031 a_50751_n19729.n161 a_50751_n19729.n168 1.5005
R51032 a_50751_n19729.n166 a_50751_n19729.n161 1.5005
R51033 a_50751_n19729.n161 a_50751_n19729.n164 1.5005
R51034 a_50751_n19729.n162 a_50751_n19729.n161 1.5005
R51035 a_50751_n19729.n158 a_50751_n19729.n221 1.5005
R51036 a_50751_n19729.n159 a_50751_n19729.n158 1.5005
R51037 a_50751_n19729.n158 a_50751_n19729.n156 1.5005
R51038 a_50751_n19729.n193 a_50751_n19729.n151 1.5005
R51039 a_50751_n19729.n146 a_50751_n19729.n154 1.5005
R51040 a_50751_n19729.n152 a_50751_n19729.n151 1.5005
R51041 a_50751_n19729.n146 a_50751_n19729.n189 1.5005
R51042 a_50751_n19729.n139 a_50751_n19729.n149 1.5005
R51043 a_50751_n19729.n147 a_50751_n19729.n146 1.5005
R51044 a_50751_n19729.n144 a_50751_n19729.n139 1.5005
R51045 a_50751_n19729.n139 a_50751_n19729.n142 1.5005
R51046 a_50751_n19729.n140 a_50751_n19729.n139 1.5005
R51047 a_50751_n19729.n139 a_50751_n19729.n137 1.5005
R51048 a_50751_n19729.n139 a_50751_n19729.n134 1.5005
R51049 a_50751_n19729.n211 a_50751_n19729.n50 1.5005
R51050 a_50751_n19729.n283 a_50751_n19729.n50 1.5005
R51051 a_50751_n19729.n47 a_50751_n19729.n207 1.5005
R51052 a_50751_n19729.n36 a_50751_n19729.n287 1.5005
R51053 a_50751_n19729.n61 a_50751_n19729.n22 1.5005
R51054 a_50751_n19729.n19 a_50751_n19729.n57 1.5005
R51055 a_50751_n19729.n6 a_50751_n19729.n225 1.5005
R51056 a_50751_n19729.n50 a_50751_n19729.n53 1.5005
R51057 a_50751_n19729.n51 a_50751_n19729.n50 1.5005
R51058 a_50751_n19729.n50 a_50751_n19729.n209 1.5005
R51059 a_50751_n19729.n48 a_50751_n19729.n47 1.5005
R51060 a_50751_n19729.n50 a_50751_n19729.n45 1.5005
R51061 a_50751_n19729.n205 a_50751_n19729.n47 1.5005
R51062 a_50751_n19729.n43 a_50751_n19729.n36 1.5005
R51063 a_50751_n19729.n47 a_50751_n19729.n41 1.5005
R51064 a_50751_n19729.n27 a_50751_n19729.n39 1.5005
R51065 a_50751_n19729.n37 a_50751_n19729.n36 1.5005
R51066 a_50751_n19729.n27 a_50751_n19729.n34 1.5005
R51067 a_50751_n19729.n32 a_50751_n19729.n27 1.5005
R51068 a_50751_n19729.n27 a_50751_n19729.n30 1.5005
R51069 a_50751_n19729.n28 a_50751_n19729.n27 1.5005
R51070 a_50751_n19729.n22 a_50751_n19729.n213 1.5005
R51071 a_50751_n19729.n22 a_50751_n19729.n25 1.5005
R51072 a_50751_n19729.n23 a_50751_n19729.n22 1.5005
R51073 a_50751_n19729.n224 a_50751_n19729.n59 1.5005
R51074 a_50751_n19729.n20 a_50751_n19729.n19 1.5005
R51075 a_50751_n19729.n224 a_50751_n19729.n17 1.5005
R51076 a_50751_n19729.n55 a_50751_n19729.n19 1.5005
R51077 a_50751_n19729.n15 a_50751_n19729.n6 1.5005
R51078 a_50751_n19729.n19 a_50751_n19729.n13 1.5005
R51079 a_50751_n19729.n11 a_50751_n19729.n6 1.5005
R51080 a_50751_n19729.n6 a_50751_n19729.n9 1.5005
R51081 a_50751_n19729.n7 a_50751_n19729.n6 1.5005
R51082 a_50751_n19729.n6 a_50751_n19729.n4 1.5005
R51083 a_50751_n19729.n6 a_50751_n19729.n1 1.5005
R51084 a_50751_n19729.n506 a_50751_n19729.n224 1.5005
R51085 a_50751_n19729.n227 a_50751_n19729.n226 1.06274
R51086 a_50751_n19729.n228 a_50751_n19729.n227 1.06274
R51087 a_50751_n19729.n331 a_50751_n19729.n330 1.06274
R51088 a_50751_n19729.n332 a_50751_n19729.n331 1.06274
R51089 a_50751_n19729.n303 a_50751_n19729.n302 1.06274
R51090 a_50751_n19729.n302 a_50751_n19729.n301 1.06274
R51091 a_50751_n19729.n380 a_50751_n19729.n379 1.06274
R51092 a_50751_n19729.n379 a_50751_n19729.n378 1.06274
R51093 a_50751_n19729.n349 a_50751_n19729.n348 1.06274
R51094 a_50751_n19729.n350 a_50751_n19729.n349 1.06274
R51095 a_50751_n19729.n426 a_50751_n19729.n425 1.06274
R51096 a_50751_n19729.n427 a_50751_n19729.n426 1.06274
R51097 a_50751_n19729.n398 a_50751_n19729.n397 1.06274
R51098 a_50751_n19729.n397 a_50751_n19729.n396 1.06274
R51099 a_50751_n19729.n475 a_50751_n19729.n474 1.06274
R51100 a_50751_n19729.n474 a_50751_n19729.n473 1.06274
R51101 a_50751_n19729.n444 a_50751_n19729.n443 1.06274
R51102 a_50751_n19729.n445 a_50751_n19729.n444 1.06274
R51103 a_50751_n19729.n286 a_50751_n19729.n285 1.06274
R51104 a_50751_n19729.n285 a_50751_n19729.n284 1.06274
R51105 a_50751_n19729.n255 a_50751_n19729.n254 1.06274
R51106 a_50751_n19729.n256 a_50751_n19729.n255 1.06274
R51107 a_50751_n19729.n509 a_50751_n19729.n508 1.06274
R51108 a_50751_n19729.n508 a_50751_n19729.n507 1.06274
R51109 a_50751_n19729.n0 a_50751_n19729.n231 0.97759
R51110 a_50751_n19729.n1 a_50751_n19729.n232 0.97759
R51111 a_50751_n19729.n230 a_50751_n19729.n229 0.97759
R51112 a_50751_n19729.n2 a_50751_n19729.n233 0.97759
R51113 a_50751_n19729.n236 a_50751_n19729.n3 0.97759
R51114 a_50751_n19729.n4 a_50751_n19729.n234 0.97759
R51115 a_50751_n19729.n5 a_50751_n19729.n237 0.97759
R51116 a_50751_n19729.n7 a_50751_n19729.n235 0.97759
R51117 a_50751_n19729.n240 a_50751_n19729.n8 0.97759
R51118 a_50751_n19729.n9 a_50751_n19729.n238 0.97759
R51119 a_50751_n19729.n10 a_50751_n19729.n241 0.97759
R51120 a_50751_n19729.n11 a_50751_n19729.n239 0.97759
R51121 a_50751_n19729.n244 a_50751_n19729.n12 0.97759
R51122 a_50751_n19729.n13 a_50751_n19729.n242 0.97759
R51123 a_50751_n19729.n14 a_50751_n19729.n245 0.97759
R51124 a_50751_n19729.n15 a_50751_n19729.n243 0.97759
R51125 a_50751_n19729.n252 a_50751_n19729.n16 0.97759
R51126 a_50751_n19729.n17 a_50751_n19729.n250 0.97759
R51127 a_50751_n19729.n18 a_50751_n19729.n253 0.97759
R51128 a_50751_n19729.n20 a_50751_n19729.n251 0.97759
R51129 a_50751_n19729.n21 a_50751_n19729.n501 0.97759
R51130 a_50751_n19729.n23 a_50751_n19729.n499 0.97759
R51131 a_50751_n19729.n500 a_50751_n19729.n24 0.97759
R51132 a_50751_n19729.n25 a_50751_n19729.n498 0.97759
R51133 a_50751_n19729.n496 a_50751_n19729.n495 0.97759
R51134 a_50751_n19729.n497 a_50751_n19729.n493 0.97759
R51135 a_50751_n19729.n26 a_50751_n19729.n299 0.97759
R51136 a_50751_n19729.n28 a_50751_n19729.n297 0.97759
R51137 a_50751_n19729.n298 a_50751_n19729.n29 0.97759
R51138 a_50751_n19729.n30 a_50751_n19729.n296 0.97759
R51139 a_50751_n19729.n31 a_50751_n19729.n295 0.97759
R51140 a_50751_n19729.n32 a_50751_n19729.n293 0.97759
R51141 a_50751_n19729.n294 a_50751_n19729.n33 0.97759
R51142 a_50751_n19729.n34 a_50751_n19729.n292 0.97759
R51143 a_50751_n19729.n35 a_50751_n19729.n291 0.97759
R51144 a_50751_n19729.n37 a_50751_n19729.n289 0.97759
R51145 a_50751_n19729.n290 a_50751_n19729.n38 0.97759
R51146 a_50751_n19729.n39 a_50751_n19729.n288 0.97759
R51147 a_50751_n19729.n259 a_50751_n19729.n40 0.97759
R51148 a_50751_n19729.n41 a_50751_n19729.n257 0.97759
R51149 a_50751_n19729.n42 a_50751_n19729.n260 0.97759
R51150 a_50751_n19729.n43 a_50751_n19729.n258 0.97759
R51151 a_50751_n19729.n267 a_50751_n19729.n44 0.97759
R51152 a_50751_n19729.n45 a_50751_n19729.n265 0.97759
R51153 a_50751_n19729.n46 a_50751_n19729.n268 0.97759
R51154 a_50751_n19729.n48 a_50751_n19729.n266 0.97759
R51155 a_50751_n19729.n49 a_50751_n19729.n278 0.97759
R51156 a_50751_n19729.n51 a_50751_n19729.n276 0.97759
R51157 a_50751_n19729.n277 a_50751_n19729.n52 0.97759
R51158 a_50751_n19729.n53 a_50751_n19729.n275 0.97759
R51159 a_50751_n19729.n273 a_50751_n19729.n272 0.97759
R51160 a_50751_n19729.n274 a_50751_n19729.n270 0.97759
R51161 a_50751_n19729.n54 a_50751_n19729.n249 0.97759
R51162 a_50751_n19729.n55 a_50751_n19729.n247 0.97759
R51163 a_50751_n19729.n248 a_50751_n19729.n56 0.97759
R51164 a_50751_n19729.n57 a_50751_n19729.n246 0.97759
R51165 a_50751_n19729.n504 a_50751_n19729.n58 0.97759
R51166 a_50751_n19729.n59 a_50751_n19729.n502 0.97759
R51167 a_50751_n19729.n60 a_50751_n19729.n505 0.97759
R51168 a_50751_n19729.n61 a_50751_n19729.n503 0.97759
R51169 a_50751_n19729.n62 a_50751_n19729.n306 0.97759
R51170 a_50751_n19729.n63 a_50751_n19729.n307 0.97759
R51171 a_50751_n19729.n305 a_50751_n19729.n304 0.97759
R51172 a_50751_n19729.n64 a_50751_n19729.n308 0.97759
R51173 a_50751_n19729.n311 a_50751_n19729.n65 0.97759
R51174 a_50751_n19729.n66 a_50751_n19729.n309 0.97759
R51175 a_50751_n19729.n67 a_50751_n19729.n312 0.97759
R51176 a_50751_n19729.n69 a_50751_n19729.n310 0.97759
R51177 a_50751_n19729.n315 a_50751_n19729.n70 0.97759
R51178 a_50751_n19729.n71 a_50751_n19729.n313 0.97759
R51179 a_50751_n19729.n72 a_50751_n19729.n316 0.97759
R51180 a_50751_n19729.n73 a_50751_n19729.n314 0.97759
R51181 a_50751_n19729.n74 a_50751_n19729.n328 0.97759
R51182 a_50751_n19729.n76 a_50751_n19729.n326 0.97759
R51183 a_50751_n19729.n327 a_50751_n19729.n77 0.97759
R51184 a_50751_n19729.n78 a_50751_n19729.n325 0.97759
R51185 a_50751_n19729.n79 a_50751_n19729.n320 0.97759
R51186 a_50751_n19729.n81 a_50751_n19729.n318 0.97759
R51187 a_50751_n19729.n319 a_50751_n19729.n82 0.97759
R51188 a_50751_n19729.n83 a_50751_n19729.n317 0.97759
R51189 a_50751_n19729.n340 a_50751_n19729.n84 0.97759
R51190 a_50751_n19729.n85 a_50751_n19729.n338 0.97759
R51191 a_50751_n19729.n86 a_50751_n19729.n341 0.97759
R51192 a_50751_n19729.n88 a_50751_n19729.n339 0.97759
R51193 a_50751_n19729.n346 a_50751_n19729.n345 0.97759
R51194 a_50751_n19729.n347 a_50751_n19729.n343 0.97759
R51195 a_50751_n19729.n89 a_50751_n19729.n393 0.97759
R51196 a_50751_n19729.n91 a_50751_n19729.n391 0.97759
R51197 a_50751_n19729.n392 a_50751_n19729.n92 0.97759
R51198 a_50751_n19729.n93 a_50751_n19729.n390 0.97759
R51199 a_50751_n19729.n94 a_50751_n19729.n389 0.97759
R51200 a_50751_n19729.n95 a_50751_n19729.n387 0.97759
R51201 a_50751_n19729.n388 a_50751_n19729.n96 0.97759
R51202 a_50751_n19729.n97 a_50751_n19729.n386 0.97759
R51203 a_50751_n19729.n98 a_50751_n19729.n385 0.97759
R51204 a_50751_n19729.n100 a_50751_n19729.n383 0.97759
R51205 a_50751_n19729.n384 a_50751_n19729.n101 0.97759
R51206 a_50751_n19729.n102 a_50751_n19729.n382 0.97759
R51207 a_50751_n19729.n353 a_50751_n19729.n103 0.97759
R51208 a_50751_n19729.n104 a_50751_n19729.n351 0.97759
R51209 a_50751_n19729.n105 a_50751_n19729.n354 0.97759
R51210 a_50751_n19729.n106 a_50751_n19729.n352 0.97759
R51211 a_50751_n19729.n361 a_50751_n19729.n107 0.97759
R51212 a_50751_n19729.n108 a_50751_n19729.n359 0.97759
R51213 a_50751_n19729.n109 a_50751_n19729.n362 0.97759
R51214 a_50751_n19729.n111 a_50751_n19729.n360 0.97759
R51215 a_50751_n19729.n112 a_50751_n19729.n372 0.97759
R51216 a_50751_n19729.n114 a_50751_n19729.n370 0.97759
R51217 a_50751_n19729.n371 a_50751_n19729.n115 0.97759
R51218 a_50751_n19729.n116 a_50751_n19729.n369 0.97759
R51219 a_50751_n19729.n367 a_50751_n19729.n366 0.97759
R51220 a_50751_n19729.n368 a_50751_n19729.n364 0.97759
R51221 a_50751_n19729.n323 a_50751_n19729.n117 0.97759
R51222 a_50751_n19729.n118 a_50751_n19729.n321 0.97759
R51223 a_50751_n19729.n119 a_50751_n19729.n324 0.97759
R51224 a_50751_n19729.n120 a_50751_n19729.n322 0.97759
R51225 a_50751_n19729.n121 a_50751_n19729.n337 0.97759
R51226 a_50751_n19729.n122 a_50751_n19729.n335 0.97759
R51227 a_50751_n19729.n336 a_50751_n19729.n123 0.97759
R51228 a_50751_n19729.n124 a_50751_n19729.n334 0.97759
R51229 a_50751_n19729.n125 a_50751_n19729.n358 0.97759
R51230 a_50751_n19729.n126 a_50751_n19729.n356 0.97759
R51231 a_50751_n19729.n357 a_50751_n19729.n127 0.97759
R51232 a_50751_n19729.n128 a_50751_n19729.n355 0.97759
R51233 a_50751_n19729.n375 a_50751_n19729.n129 0.97759
R51234 a_50751_n19729.n130 a_50751_n19729.n373 0.97759
R51235 a_50751_n19729.n131 a_50751_n19729.n376 0.97759
R51236 a_50751_n19729.n132 a_50751_n19729.n374 0.97759
R51237 a_50751_n19729.n133 a_50751_n19729.n401 0.97759
R51238 a_50751_n19729.n134 a_50751_n19729.n402 0.97759
R51239 a_50751_n19729.n400 a_50751_n19729.n399 0.97759
R51240 a_50751_n19729.n135 a_50751_n19729.n403 0.97759
R51241 a_50751_n19729.n406 a_50751_n19729.n136 0.97759
R51242 a_50751_n19729.n137 a_50751_n19729.n404 0.97759
R51243 a_50751_n19729.n138 a_50751_n19729.n407 0.97759
R51244 a_50751_n19729.n140 a_50751_n19729.n405 0.97759
R51245 a_50751_n19729.n410 a_50751_n19729.n141 0.97759
R51246 a_50751_n19729.n142 a_50751_n19729.n408 0.97759
R51247 a_50751_n19729.n143 a_50751_n19729.n411 0.97759
R51248 a_50751_n19729.n144 a_50751_n19729.n409 0.97759
R51249 a_50751_n19729.n145 a_50751_n19729.n423 0.97759
R51250 a_50751_n19729.n147 a_50751_n19729.n421 0.97759
R51251 a_50751_n19729.n422 a_50751_n19729.n148 0.97759
R51252 a_50751_n19729.n149 a_50751_n19729.n420 0.97759
R51253 a_50751_n19729.n150 a_50751_n19729.n415 0.97759
R51254 a_50751_n19729.n152 a_50751_n19729.n413 0.97759
R51255 a_50751_n19729.n414 a_50751_n19729.n153 0.97759
R51256 a_50751_n19729.n154 a_50751_n19729.n412 0.97759
R51257 a_50751_n19729.n435 a_50751_n19729.n155 0.97759
R51258 a_50751_n19729.n156 a_50751_n19729.n433 0.97759
R51259 a_50751_n19729.n157 a_50751_n19729.n436 0.97759
R51260 a_50751_n19729.n159 a_50751_n19729.n434 0.97759
R51261 a_50751_n19729.n441 a_50751_n19729.n440 0.97759
R51262 a_50751_n19729.n442 a_50751_n19729.n438 0.97759
R51263 a_50751_n19729.n160 a_50751_n19729.n488 0.97759
R51264 a_50751_n19729.n162 a_50751_n19729.n486 0.97759
R51265 a_50751_n19729.n487 a_50751_n19729.n163 0.97759
R51266 a_50751_n19729.n164 a_50751_n19729.n485 0.97759
R51267 a_50751_n19729.n165 a_50751_n19729.n484 0.97759
R51268 a_50751_n19729.n166 a_50751_n19729.n482 0.97759
R51269 a_50751_n19729.n483 a_50751_n19729.n167 0.97759
R51270 a_50751_n19729.n168 a_50751_n19729.n481 0.97759
R51271 a_50751_n19729.n169 a_50751_n19729.n480 0.97759
R51272 a_50751_n19729.n171 a_50751_n19729.n478 0.97759
R51273 a_50751_n19729.n479 a_50751_n19729.n172 0.97759
R51274 a_50751_n19729.n173 a_50751_n19729.n477 0.97759
R51275 a_50751_n19729.n448 a_50751_n19729.n174 0.97759
R51276 a_50751_n19729.n175 a_50751_n19729.n446 0.97759
R51277 a_50751_n19729.n176 a_50751_n19729.n449 0.97759
R51278 a_50751_n19729.n177 a_50751_n19729.n447 0.97759
R51279 a_50751_n19729.n456 a_50751_n19729.n178 0.97759
R51280 a_50751_n19729.n179 a_50751_n19729.n454 0.97759
R51281 a_50751_n19729.n180 a_50751_n19729.n457 0.97759
R51282 a_50751_n19729.n182 a_50751_n19729.n455 0.97759
R51283 a_50751_n19729.n183 a_50751_n19729.n467 0.97759
R51284 a_50751_n19729.n185 a_50751_n19729.n465 0.97759
R51285 a_50751_n19729.n466 a_50751_n19729.n186 0.97759
R51286 a_50751_n19729.n187 a_50751_n19729.n464 0.97759
R51287 a_50751_n19729.n462 a_50751_n19729.n461 0.97759
R51288 a_50751_n19729.n463 a_50751_n19729.n459 0.97759
R51289 a_50751_n19729.n418 a_50751_n19729.n188 0.97759
R51290 a_50751_n19729.n189 a_50751_n19729.n416 0.97759
R51291 a_50751_n19729.n190 a_50751_n19729.n419 0.97759
R51292 a_50751_n19729.n191 a_50751_n19729.n417 0.97759
R51293 a_50751_n19729.n192 a_50751_n19729.n432 0.97759
R51294 a_50751_n19729.n193 a_50751_n19729.n430 0.97759
R51295 a_50751_n19729.n431 a_50751_n19729.n194 0.97759
R51296 a_50751_n19729.n195 a_50751_n19729.n429 0.97759
R51297 a_50751_n19729.n196 a_50751_n19729.n453 0.97759
R51298 a_50751_n19729.n197 a_50751_n19729.n451 0.97759
R51299 a_50751_n19729.n452 a_50751_n19729.n198 0.97759
R51300 a_50751_n19729.n199 a_50751_n19729.n450 0.97759
R51301 a_50751_n19729.n470 a_50751_n19729.n200 0.97759
R51302 a_50751_n19729.n201 a_50751_n19729.n468 0.97759
R51303 a_50751_n19729.n202 a_50751_n19729.n471 0.97759
R51304 a_50751_n19729.n203 a_50751_n19729.n469 0.97759
R51305 a_50751_n19729.n204 a_50751_n19729.n264 0.97759
R51306 a_50751_n19729.n205 a_50751_n19729.n262 0.97759
R51307 a_50751_n19729.n263 a_50751_n19729.n206 0.97759
R51308 a_50751_n19729.n207 a_50751_n19729.n261 0.97759
R51309 a_50751_n19729.n281 a_50751_n19729.n208 0.97759
R51310 a_50751_n19729.n209 a_50751_n19729.n279 0.97759
R51311 a_50751_n19729.n210 a_50751_n19729.n282 0.97759
R51312 a_50751_n19729.n211 a_50751_n19729.n280 0.97759
R51313 a_50751_n19729.n494 a_50751_n19729.n212 0.931516
R51314 a_50751_n19729.n213 a_50751_n19729.n492 0.931516
R51315 a_50751_n19729.n271 a_50751_n19729.n214 0.931516
R51316 a_50751_n19729.n215 a_50751_n19729.n269 0.931516
R51317 a_50751_n19729.n344 a_50751_n19729.n216 0.931516
R51318 a_50751_n19729.n217 a_50751_n19729.n342 0.931516
R51319 a_50751_n19729.n365 a_50751_n19729.n218 0.931516
R51320 a_50751_n19729.n219 a_50751_n19729.n363 0.931516
R51321 a_50751_n19729.n439 a_50751_n19729.n220 0.931516
R51322 a_50751_n19729.n221 a_50751_n19729.n437 0.931516
R51323 a_50751_n19729.n460 a_50751_n19729.n222 0.931516
R51324 a_50751_n19729.n223 a_50751_n19729.n458 0.931516
R51325 a_50751_n19729.n113 a_50751_n19729.n110 0.82023
R51326 a_50751_n19729.n184 a_50751_n19729.n181 0.82023
R51327 a_50751_n19729.n50 a_50751_n19729.n47 0.82023
R51328 a_50751_n19729.n68 a_50751_n19729.n75 0.818405
R51329 a_50751_n19729.n139 a_50751_n19729.n146 0.818405
R51330 a_50751_n19729.n19 a_50751_n19729.n6 0.818405
R51331 a_50751_n19729.n490 a_50751_n19729.n489 0.7505
R51332 a_50751_n19729.n395 a_50751_n19729.n394 0.7505
R51333 a_50751_n19729.n394 a_50751_n19729.n90 0.717155
R51334 a_50751_n19729.n489 a_50751_n19729.n161 0.717155
R51335 a_50751_n19729.n491 a_50751_n19729.n27 0.717155
R51336 a_50751_n19729.n87 a_50751_n19729.n80 0.639622
R51337 a_50751_n19729.n158 a_50751_n19729.n151 0.639622
R51338 a_50751_n19729.n224 a_50751_n19729.n22 0.639622
R51339 a_50751_n19729.n497 a_50751_n19729.n496 0.62434
R51340 a_50751_n19729.n274 a_50751_n19729.n273 0.62434
R51341 a_50751_n19729.n347 a_50751_n19729.n346 0.62434
R51342 a_50751_n19729.n368 a_50751_n19729.n367 0.62434
R51343 a_50751_n19729.n442 a_50751_n19729.n441 0.62434
R51344 a_50751_n19729.n463 a_50751_n19729.n462 0.62434
R51345 a_50751_n19729.n211 a_50751_n19729.n210 0.62434
R51346 a_50751_n19729.n209 a_50751_n19729.n208 0.62434
R51347 a_50751_n19729.n207 a_50751_n19729.n206 0.62434
R51348 a_50751_n19729.n205 a_50751_n19729.n204 0.62434
R51349 a_50751_n19729.n203 a_50751_n19729.n202 0.62434
R51350 a_50751_n19729.n201 a_50751_n19729.n200 0.62434
R51351 a_50751_n19729.n199 a_50751_n19729.n198 0.62434
R51352 a_50751_n19729.n197 a_50751_n19729.n196 0.62434
R51353 a_50751_n19729.n195 a_50751_n19729.n194 0.62434
R51354 a_50751_n19729.n193 a_50751_n19729.n192 0.62434
R51355 a_50751_n19729.n191 a_50751_n19729.n190 0.62434
R51356 a_50751_n19729.n189 a_50751_n19729.n188 0.62434
R51357 a_50751_n19729.n187 a_50751_n19729.n186 0.62434
R51358 a_50751_n19729.n185 a_50751_n19729.n183 0.62434
R51359 a_50751_n19729.n182 a_50751_n19729.n180 0.62434
R51360 a_50751_n19729.n179 a_50751_n19729.n178 0.62434
R51361 a_50751_n19729.n177 a_50751_n19729.n176 0.62434
R51362 a_50751_n19729.n175 a_50751_n19729.n174 0.62434
R51363 a_50751_n19729.n173 a_50751_n19729.n172 0.62434
R51364 a_50751_n19729.n171 a_50751_n19729.n169 0.62434
R51365 a_50751_n19729.n168 a_50751_n19729.n167 0.62434
R51366 a_50751_n19729.n166 a_50751_n19729.n165 0.62434
R51367 a_50751_n19729.n164 a_50751_n19729.n163 0.62434
R51368 a_50751_n19729.n162 a_50751_n19729.n160 0.62434
R51369 a_50751_n19729.n159 a_50751_n19729.n157 0.62434
R51370 a_50751_n19729.n156 a_50751_n19729.n155 0.62434
R51371 a_50751_n19729.n154 a_50751_n19729.n153 0.62434
R51372 a_50751_n19729.n152 a_50751_n19729.n150 0.62434
R51373 a_50751_n19729.n149 a_50751_n19729.n148 0.62434
R51374 a_50751_n19729.n147 a_50751_n19729.n145 0.62434
R51375 a_50751_n19729.n144 a_50751_n19729.n143 0.62434
R51376 a_50751_n19729.n142 a_50751_n19729.n141 0.62434
R51377 a_50751_n19729.n140 a_50751_n19729.n138 0.62434
R51378 a_50751_n19729.n137 a_50751_n19729.n136 0.62434
R51379 a_50751_n19729.n399 a_50751_n19729.n135 0.62434
R51380 a_50751_n19729.n134 a_50751_n19729.n133 0.62434
R51381 a_50751_n19729.n132 a_50751_n19729.n131 0.62434
R51382 a_50751_n19729.n130 a_50751_n19729.n129 0.62434
R51383 a_50751_n19729.n128 a_50751_n19729.n127 0.62434
R51384 a_50751_n19729.n126 a_50751_n19729.n125 0.62434
R51385 a_50751_n19729.n124 a_50751_n19729.n123 0.62434
R51386 a_50751_n19729.n122 a_50751_n19729.n121 0.62434
R51387 a_50751_n19729.n120 a_50751_n19729.n119 0.62434
R51388 a_50751_n19729.n118 a_50751_n19729.n117 0.62434
R51389 a_50751_n19729.n116 a_50751_n19729.n115 0.62434
R51390 a_50751_n19729.n114 a_50751_n19729.n112 0.62434
R51391 a_50751_n19729.n111 a_50751_n19729.n109 0.62434
R51392 a_50751_n19729.n108 a_50751_n19729.n107 0.62434
R51393 a_50751_n19729.n106 a_50751_n19729.n105 0.62434
R51394 a_50751_n19729.n104 a_50751_n19729.n103 0.62434
R51395 a_50751_n19729.n102 a_50751_n19729.n101 0.62434
R51396 a_50751_n19729.n100 a_50751_n19729.n98 0.62434
R51397 a_50751_n19729.n97 a_50751_n19729.n96 0.62434
R51398 a_50751_n19729.n95 a_50751_n19729.n94 0.62434
R51399 a_50751_n19729.n93 a_50751_n19729.n92 0.62434
R51400 a_50751_n19729.n91 a_50751_n19729.n89 0.62434
R51401 a_50751_n19729.n88 a_50751_n19729.n86 0.62434
R51402 a_50751_n19729.n85 a_50751_n19729.n84 0.62434
R51403 a_50751_n19729.n83 a_50751_n19729.n82 0.62434
R51404 a_50751_n19729.n81 a_50751_n19729.n79 0.62434
R51405 a_50751_n19729.n78 a_50751_n19729.n77 0.62434
R51406 a_50751_n19729.n76 a_50751_n19729.n74 0.62434
R51407 a_50751_n19729.n73 a_50751_n19729.n72 0.62434
R51408 a_50751_n19729.n71 a_50751_n19729.n70 0.62434
R51409 a_50751_n19729.n69 a_50751_n19729.n67 0.62434
R51410 a_50751_n19729.n66 a_50751_n19729.n65 0.62434
R51411 a_50751_n19729.n304 a_50751_n19729.n64 0.62434
R51412 a_50751_n19729.n63 a_50751_n19729.n62 0.62434
R51413 a_50751_n19729.n61 a_50751_n19729.n60 0.62434
R51414 a_50751_n19729.n59 a_50751_n19729.n58 0.62434
R51415 a_50751_n19729.n57 a_50751_n19729.n56 0.62434
R51416 a_50751_n19729.n55 a_50751_n19729.n54 0.62434
R51417 a_50751_n19729.n53 a_50751_n19729.n52 0.62434
R51418 a_50751_n19729.n51 a_50751_n19729.n49 0.62434
R51419 a_50751_n19729.n48 a_50751_n19729.n46 0.62434
R51420 a_50751_n19729.n45 a_50751_n19729.n44 0.62434
R51421 a_50751_n19729.n43 a_50751_n19729.n42 0.62434
R51422 a_50751_n19729.n41 a_50751_n19729.n40 0.62434
R51423 a_50751_n19729.n39 a_50751_n19729.n38 0.62434
R51424 a_50751_n19729.n37 a_50751_n19729.n35 0.62434
R51425 a_50751_n19729.n34 a_50751_n19729.n33 0.62434
R51426 a_50751_n19729.n32 a_50751_n19729.n31 0.62434
R51427 a_50751_n19729.n30 a_50751_n19729.n29 0.62434
R51428 a_50751_n19729.n28 a_50751_n19729.n26 0.62434
R51429 a_50751_n19729.n25 a_50751_n19729.n24 0.62434
R51430 a_50751_n19729.n23 a_50751_n19729.n21 0.62434
R51431 a_50751_n19729.n20 a_50751_n19729.n18 0.62434
R51432 a_50751_n19729.n17 a_50751_n19729.n16 0.62434
R51433 a_50751_n19729.n15 a_50751_n19729.n14 0.62434
R51434 a_50751_n19729.n13 a_50751_n19729.n12 0.62434
R51435 a_50751_n19729.n11 a_50751_n19729.n10 0.62434
R51436 a_50751_n19729.n9 a_50751_n19729.n8 0.62434
R51437 a_50751_n19729.n7 a_50751_n19729.n5 0.62434
R51438 a_50751_n19729.n4 a_50751_n19729.n3 0.62434
R51439 a_50751_n19729.n229 a_50751_n19729.n2 0.62434
R51440 a_50751_n19729.n1 a_50751_n19729.n0 0.62434
R51441 a_50751_n19729.n394 a_50751_n19729.n87 0.617426
R51442 a_50751_n19729.n489 a_50751_n19729.n158 0.617426
R51443 a_50751_n19729.n22 a_50751_n19729.n491 0.617426
R51444 a_50751_n19729.n223 a_50751_n19729.n222 0.595087
R51445 a_50751_n19729.n221 a_50751_n19729.n220 0.595087
R51446 a_50751_n19729.n219 a_50751_n19729.n218 0.595087
R51447 a_50751_n19729.n217 a_50751_n19729.n216 0.595087
R51448 a_50751_n19729.n215 a_50751_n19729.n214 0.595087
R51449 a_50751_n19729.n213 a_50751_n19729.n212 0.595087
R51450 a_50751_n19729.n75 a_50751_n19729.n80 0.545973
R51451 a_50751_n19729.n146 a_50751_n19729.n151 0.545973
R51452 a_50751_n19729.n224 a_50751_n19729.n19 0.545973
R51453 a_50751_n19729.n110 a_50751_n19729.n99 0.545365
R51454 a_50751_n19729.n181 a_50751_n19729.n170 0.545365
R51455 a_50751_n19729.n47 a_50751_n19729.n36 0.545365
R51456 a_50751_n19729.n27 a_50751_n19729.n36 0.452324
R51457 a_50751_n19729.n161 a_50751_n19729.n170 0.452324
R51458 a_50751_n19729.n90 a_50751_n19729.n99 0.452324
R51459 a_65486_n36322.n0 a_65486_n36322.t18 13.7934
R51460 a_65486_n36322.n2 a_65486_n36322.t3 10.7024
R51461 a_65486_n36322.n2 a_65486_n36322.t5 10.1668
R51462 a_65486_n36322.n2 a_65486_n36322.t4 9.64458
R51463 a_65486_n36322.n2 a_65486_n36322.t1 9.27635
R51464 a_65486_n36322.n2 a_65486_n36322.n0 8.75198
R51465 a_65486_n36322.n0 a_65486_n36322.t17 8.14051
R51466 a_65486_n36322.n0 a_65486_n36322.t15 8.14051
R51467 a_65486_n36322.n0 a_65486_n36322.t23 8.14051
R51468 a_65486_n36322.n0 a_65486_n36322.t8 8.14051
R51469 a_65486_n36322.n0 a_65486_n36322.t21 8.06917
R51470 a_65486_n36322.n0 a_65486_n36322.t12 8.06917
R51471 a_65486_n36322.n0 a_65486_n36322.t10 8.06917
R51472 a_65486_n36322.n0 a_65486_n36322.t11 8.06917
R51473 a_65486_n36322.n0 a_65486_n36322.t9 8.06917
R51474 a_65486_n36322.n0 a_65486_n36322.t16 8.06917
R51475 a_65486_n36322.n0 a_65486_n36322.t19 8.06917
R51476 a_65486_n36322.n1 a_65486_n36322.t7 7.94157
R51477 a_65486_n36322.n2 a_65486_n36322.t2 7.72643
R51478 a_65486_n36322.n1 a_65486_n36322.t6 7.22925
R51479 a_65486_n36322.t0 a_65486_n36322.n2 7.17912
R51480 a_65486_n36322.n0 a_65486_n36322.t14 8.33554
R51481 a_65486_n36322.t13 a_65486_n36322.n0 8.33554
R51482 a_65486_n36322.n0 a_65486_n36322.t20 8.33647
R51483 a_65486_n36322.t22 a_65486_n36322.n0 8.33647
R51484 a_65486_n36322.n2 a_65486_n36322.n1 7.46075
R51485 a_71342_n30339.n0 a_71342_n30339.t1 10.3838
R51486 a_71342_n30339.n0 a_71342_n30339.t2 10.3566
R51487 a_71342_n30339.n0 a_71342_n30339.t3 10.0407
R51488 a_71342_n30339.t0 a_71342_n30339.n0 9.57605
R51489 a_106809_n17715.t0 a_106809_n17715.t1 12.8122
R51490 a_33249_48695.n109 a_33249_48695.n106 7.94229
R51491 a_33249_48695.n140 a_33249_48695.n137 7.94229
R51492 a_33249_48695.n394 a_33249_48695.n393 7.22198
R51493 a_33249_48695.n364 a_33249_48695.n363 7.22198
R51494 a_33249_48695.n68 a_33249_48695.t317 6.77653
R51495 a_33249_48695.n47 a_33249_48695.t244 6.77653
R51496 a_33249_48695.n64 a_33249_48695.t178 6.7761
R51497 a_33249_48695.n377 a_33249_48695.t253 6.7761
R51498 a_33249_48695.n9 a_33249_48695.t257 6.77231
R51499 a_33249_48695.n19 a_33249_48695.t205 6.77231
R51500 a_33249_48695.n267 a_33249_48695.t42 6.58663
R51501 a_33249_48695.n223 a_33249_48695.t44 6.58663
R51502 a_33249_48695.n335 a_33249_48695.n334 6.50088
R51503 a_33249_48695.n300 a_33249_48695.n296 6.50088
R51504 a_33249_48695.n268 a_33249_48695.n265 5.95439
R51505 a_33249_48695.n224 a_33249_48695.n221 5.95439
R51506 a_33249_48695.n108 a_33249_48695.t308 5.69423
R51507 a_33249_48695.n90 a_33249_48695.t291 5.69423
R51508 a_33249_48695.n139 a_33249_48695.t201 5.69423
R51509 a_33249_48695.n135 a_33249_48695.t186 5.69423
R51510 a_33249_48695.n61 a_33249_48695.t327 5.50607
R51511 a_33249_48695.n48 a_33249_48695.t266 5.50607
R51512 a_33249_48695.n374 a_33249_48695.t224 5.50607
R51513 a_33249_48695.n69 a_33249_48695.t167 5.50607
R51514 a_33249_48695.n62 a_33249_48695.t215 5.50475
R51515 a_33249_48695.n58 a_33249_48695.t319 5.50475
R51516 a_33249_48695.n57 a_33249_48695.t163 5.50475
R51517 a_33249_48695.n375 a_33249_48695.t289 5.50475
R51518 a_33249_48695.n371 a_33249_48695.t214 5.50475
R51519 a_33249_48695.n370 a_33249_48695.t237 5.50475
R51520 a_33249_48695.n70 a_33249_48695.t229 5.50475
R51521 a_33249_48695.t334 a_33249_48695.n397 5.50475
R51522 a_33249_48695.n108 a_33249_48695.n107 5.49558
R51523 a_33249_48695.n139 a_33249_48695.n138 5.49558
R51524 a_33249_48695.n265 a_33249_48695.t59 5.31528
R51525 a_33249_48695.n221 a_33249_48695.t67 5.31528
R51526 a_33249_48695.n80 a_33249_48695.n78 4.92758
R51527 a_33249_48695.n306 a_33249_48695.n304 4.92758
R51528 a_33249_48695.n38 a_33249_48695.n273 4.92217
R51529 a_33249_48695.n45 a_33249_48695.n286 4.92217
R51530 a_33249_48695.n26 a_33249_48695.n88 4.22068
R51531 a_33249_48695.n27 a_33249_48695.t270 5.69068
R51532 a_33249_48695.n28 a_33249_48695.n87 4.22068
R51533 a_33249_48695.n29 a_33249_48695.n131 4.22068
R51534 a_33249_48695.n30 a_33249_48695.t326 5.69068
R51535 a_33249_48695.n31 a_33249_48695.n130 4.22068
R51536 a_33249_48695.n21 a_33249_48695.n184 3.84173
R51537 a_33249_48695.n24 a_33249_48695.n180 3.84173
R51538 a_33249_48695.n32 a_33249_48695.n280 3.65107
R51539 a_33249_48695.n33 a_33249_48695.n279 3.65107
R51540 a_33249_48695.n34 a_33249_48695.n278 3.65107
R51541 a_33249_48695.n35 a_33249_48695.n277 3.65107
R51542 a_33249_48695.n276 a_33249_48695.n36 3.65107
R51543 a_33249_48695.n275 a_33249_48695.n37 3.65107
R51544 a_33249_48695.n274 a_33249_48695.n38 3.65107
R51545 a_33249_48695.n39 a_33249_48695.n293 3.65107
R51546 a_33249_48695.n40 a_33249_48695.n292 3.65107
R51547 a_33249_48695.n41 a_33249_48695.n291 3.65107
R51548 a_33249_48695.n42 a_33249_48695.n290 3.65107
R51549 a_33249_48695.n289 a_33249_48695.n43 3.65107
R51550 a_33249_48695.n288 a_33249_48695.n44 3.65107
R51551 a_33249_48695.n287 a_33249_48695.n45 3.65107
R51552 a_33249_48695.n0 a_33249_48695.n384 4.0312
R51553 a_33249_48695.t230 a_33249_48695.n1 5.5012
R51554 a_33249_48695.t162 a_33249_48695.n2 5.5012
R51555 a_33249_48695.n383 a_33249_48695.n3 4.0312
R51556 a_33249_48695.t333 a_33249_48695.n4 5.5012
R51557 a_33249_48695.t175 a_33249_48695.n5 5.5012
R51558 a_33249_48695.n382 a_33249_48695.n6 4.0312
R51559 a_33249_48695.t170 a_33249_48695.n7 5.5012
R51560 a_33249_48695.t281 a_33249_48695.n8 5.5012
R51561 a_33249_48695.n380 a_33249_48695.n9 4.0312
R51562 a_33249_48695.n10 a_33249_48695.n75 4.0312
R51563 a_33249_48695.n11 a_33249_48695.t180 5.5012
R51564 a_33249_48695.n12 a_33249_48695.t284 5.5012
R51565 a_33249_48695.n13 a_33249_48695.n74 4.0312
R51566 a_33249_48695.n14 a_33249_48695.t280 5.5012
R51567 a_33249_48695.n15 a_33249_48695.t299 5.5012
R51568 a_33249_48695.n16 a_33249_48695.n73 4.0312
R51569 a_33249_48695.t295 a_33249_48695.n17 5.5012
R51570 a_33249_48695.t231 a_33249_48695.n18 5.5012
R51571 a_33249_48695.n72 a_33249_48695.n19 4.0312
R51572 a_33249_48695.n20 a_33249_48695.t81 5.31173
R51573 a_33249_48695.n22 a_33249_48695.t87 5.31173
R51574 a_33249_48695.n23 a_33249_48695.t76 5.31173
R51575 a_33249_48695.n25 a_33249_48695.t79 5.31173
R51576 a_33249_48695.n264 a_33249_48695.n262 4.50663
R51577 a_33249_48695.n220 a_33249_48695.n179 4.50663
R51578 a_33249_48695.n185 a_33249_48695.n22 4.46113
R51579 a_33249_48695.n392 a_33249_48695.t160 4.24002
R51580 a_33249_48695.n52 a_33249_48695.t320 4.24002
R51581 a_33249_48695.n362 a_33249_48695.t282 4.24002
R51582 a_33249_48695.n353 a_33249_48695.t265 4.24002
R51583 a_33249_48695.n106 a_33249_48695.n105 4.22423
R51584 a_33249_48695.n137 a_33249_48695.n136 4.22423
R51585 a_33249_48695.n301 a_33249_48695.t340 4.06712
R51586 a_33249_48695.n284 a_33249_48695.t130 4.06712
R51587 a_33249_48695.n329 a_33249_48695.t335 4.06712
R51588 a_33249_48695.n327 a_33249_48695.t125 4.06712
R51589 a_33249_48695.n96 a_33249_48695.t207 4.05054
R51590 a_33249_48695.n101 a_33249_48695.t246 4.05054
R51591 a_33249_48695.n103 a_33249_48695.t177 4.05054
R51592 a_33249_48695.n116 a_33249_48695.t172 4.05054
R51593 a_33249_48695.n118 a_33249_48695.t189 4.05054
R51594 a_33249_48695.n124 a_33249_48695.t184 4.05054
R51595 a_33249_48695.n126 a_33249_48695.t298 4.05054
R51596 a_33249_48695.n91 a_33249_48695.t269 4.05054
R51597 a_33249_48695.n164 a_33249_48695.t330 4.05054
R51598 a_33249_48695.n169 a_33249_48695.t194 4.05054
R51599 a_33249_48695.n171 a_33249_48695.t302 4.05054
R51600 a_33249_48695.n158 a_33249_48695.t297 4.05054
R51601 a_33249_48695.n156 a_33249_48695.t314 4.05054
R51602 a_33249_48695.n150 a_33249_48695.t311 4.05054
R51603 a_33249_48695.n148 a_33249_48695.t248 4.05054
R51604 a_33249_48695.n142 a_33249_48695.t223 4.05054
R51605 a_33249_48695.n64 a_33249_48695.n63 4.03475
R51606 a_33249_48695.n60 a_33249_48695.n59 4.03475
R51607 a_33249_48695.n50 a_33249_48695.n49 4.03475
R51608 a_33249_48695.n47 a_33249_48695.n46 4.03475
R51609 a_33249_48695.n377 a_33249_48695.n376 4.03475
R51610 a_33249_48695.n373 a_33249_48695.n372 4.03475
R51611 a_33249_48695.n369 a_33249_48695.n368 4.03475
R51612 a_33249_48695.n68 a_33249_48695.n67 4.03475
R51613 a_33249_48695.n330 a_33249_48695.n77 3.96014
R51614 a_33249_48695.n303 a_33249_48695.n302 3.96014
R51615 a_33249_48695.n96 a_33249_48695.t165 3.87765
R51616 a_33249_48695.n101 a_33249_48695.t199 3.87765
R51617 a_33249_48695.n103 a_33249_48695.t310 3.87765
R51618 a_33249_48695.n116 a_33249_48695.t304 3.87765
R51619 a_33249_48695.n118 a_33249_48695.t323 3.87765
R51620 a_33249_48695.n124 a_33249_48695.t318 3.87765
R51621 a_33249_48695.n126 a_33249_48695.t256 3.87765
R51622 a_33249_48695.n91 a_33249_48695.t227 3.87765
R51623 a_33249_48695.n164 a_33249_48695.t239 3.87765
R51624 a_33249_48695.n169 a_33249_48695.t272 3.87765
R51625 a_33249_48695.n171 a_33249_48695.t206 3.87765
R51626 a_33249_48695.n158 a_33249_48695.t198 3.87765
R51627 a_33249_48695.n156 a_33249_48695.t218 3.87765
R51628 a_33249_48695.n150 a_33249_48695.t212 3.87765
R51629 a_33249_48695.n148 a_33249_48695.t328 3.87765
R51630 a_33249_48695.n142 a_33249_48695.t301 3.87765
R51631 a_33249_48695.n301 a_33249_48695.t339 3.86107
R51632 a_33249_48695.n284 a_33249_48695.t128 3.86107
R51633 a_33249_48695.n329 a_33249_48695.t105 3.86107
R51634 a_33249_48695.n327 a_33249_48695.t119 3.86107
R51635 a_33249_48695.n267 a_33249_48695.n266 3.84528
R51636 a_33249_48695.n264 a_33249_48695.n263 3.84528
R51637 a_33249_48695.n223 a_33249_48695.n222 3.84528
R51638 a_33249_48695.n220 a_33249_48695.n219 3.84528
R51639 a_33249_48695.n256 a_33249_48695.n252 3.79678
R51640 a_33249_48695.n239 a_33249_48695.n235 3.79678
R51641 a_33249_48695.n197 a_33249_48695.n193 3.79678
R51642 a_33249_48695.n212 a_33249_48695.n208 3.79678
R51643 a_33249_48695.n82 a_33249_48695.n80 3.79678
R51644 a_33249_48695.n344 a_33249_48695.n342 3.79678
R51645 a_33249_48695.n308 a_33249_48695.n306 3.79678
R51646 a_33249_48695.n317 a_33249_48695.n315 3.79678
R51647 a_33249_48695.n228 a_33249_48695.n25 3.87644
R51648 a_33249_48695.n248 a_33249_48695.n244 3.73034
R51649 a_33249_48695.n217 a_33249_48695.n201 3.73034
R51650 a_33249_48695.n392 a_33249_48695.t292 3.68818
R51651 a_33249_48695.n52 a_33249_48695.t274 3.68818
R51652 a_33249_48695.n362 a_33249_48695.t187 3.68818
R51653 a_33249_48695.n353 a_33249_48695.t173 3.68818
R51654 a_33249_48695.n346 a_33249_48695.n345 3.65581
R51655 a_33249_48695.n344 a_33249_48695.n343 3.65581
R51656 a_33249_48695.n342 a_33249_48695.n341 3.65581
R51657 a_33249_48695.n340 a_33249_48695.n339 3.65581
R51658 a_33249_48695.n84 a_33249_48695.n83 3.65581
R51659 a_33249_48695.n82 a_33249_48695.n81 3.65581
R51660 a_33249_48695.n80 a_33249_48695.n79 3.65581
R51661 a_33249_48695.n319 a_33249_48695.n318 3.65581
R51662 a_33249_48695.n317 a_33249_48695.n316 3.65581
R51663 a_33249_48695.n315 a_33249_48695.n314 3.65581
R51664 a_33249_48695.n313 a_33249_48695.n312 3.65581
R51665 a_33249_48695.n310 a_33249_48695.n309 3.65581
R51666 a_33249_48695.n308 a_33249_48695.n307 3.65581
R51667 a_33249_48695.n306 a_33249_48695.n305 3.65581
R51668 a_33249_48695.n340 a_33249_48695.n338 3.64443
R51669 a_33249_48695.n313 a_33249_48695.n311 3.64443
R51670 a_33249_48695.n322 a_33249_48695.n35 3.64223
R51671 a_33249_48695.n294 a_33249_48695.n42 3.64223
R51672 a_33249_48695.n129 a_33249_48695.n90 3.25667
R51673 a_33249_48695.n391 a_33249_48695.n387 3.23904
R51674 a_33249_48695.n361 a_33249_48695.n66 3.23904
R51675 a_33249_48695.n133 a_33249_48695.n31 3.15553
R51676 a_33249_48695.n177 a_33249_48695.n28 3.15553
R51677 a_33249_48695.n268 a_33249_48695.n267 3.00663
R51678 a_33249_48695.n224 a_33249_48695.n223 3.00663
R51679 a_33249_48695.n231 a_33249_48695.n229 2.7866
R51680 a_33249_48695.n234 a_33249_48695.n232 2.7866
R51681 a_33249_48695.n238 a_33249_48695.n236 2.7866
R51682 a_33249_48695.n242 a_33249_48695.n240 2.7866
R51683 a_33249_48695.n247 a_33249_48695.n245 2.7866
R51684 a_33249_48695.n251 a_33249_48695.n249 2.7866
R51685 a_33249_48695.n255 a_33249_48695.n253 2.7866
R51686 a_33249_48695.n259 a_33249_48695.n257 2.7866
R51687 a_33249_48695.n204 a_33249_48695.n202 2.7866
R51688 a_33249_48695.n207 a_33249_48695.n205 2.7866
R51689 a_33249_48695.n211 a_33249_48695.n209 2.7866
R51690 a_33249_48695.n215 a_33249_48695.n213 2.7866
R51691 a_33249_48695.n200 a_33249_48695.n198 2.7866
R51692 a_33249_48695.n196 a_33249_48695.n194 2.7866
R51693 a_33249_48695.n192 a_33249_48695.n190 2.7866
R51694 a_33249_48695.n188 a_33249_48695.n186 2.7866
R51695 a_33249_48695.n390 a_33249_48695.n389 2.77002
R51696 a_33249_48695.n55 a_33249_48695.n54 2.77002
R51697 a_33249_48695.n360 a_33249_48695.n359 2.77002
R51698 a_33249_48695.n356 a_33249_48695.n355 2.77002
R51699 a_33249_48695.n56 a_33249_48695.n52 2.73714
R51700 a_33249_48695.n357 a_33249_48695.n353 2.73714
R51701 a_33249_48695.n95 a_33249_48695.n91 2.73714
R51702 a_33249_48695.n146 a_33249_48695.n142 2.73714
R51703 a_33249_48695.n328 a_33249_48695.n326 2.73714
R51704 a_33249_48695.n285 a_33249_48695.n283 2.73714
R51705 a_33249_48695.n235 a_33249_48695.n231 2.73672
R51706 a_33249_48695.n208 a_33249_48695.n204 2.73672
R51707 a_33249_48695.n100 a_33249_48695.n96 2.73672
R51708 a_33249_48695.n168 a_33249_48695.n164 2.73672
R51709 a_33249_48695.n371 a_33249_48695.n370 2.60203
R51710 a_33249_48695.n119 a_33249_48695.n117 2.60203
R51711 a_33249_48695.n159 a_33249_48695.n157 2.60203
R51712 a_33249_48695.n58 a_33249_48695.n57 2.60203
R51713 a_33249_48695.n299 a_33249_48695.n297 2.59712
R51714 a_33249_48695.n283 a_33249_48695.n281 2.59712
R51715 a_33249_48695.n333 a_33249_48695.n331 2.59712
R51716 a_33249_48695.n326 a_33249_48695.n324 2.59712
R51717 a_33249_48695.n99 a_33249_48695.n98 2.58054
R51718 a_33249_48695.n114 a_33249_48695.n113 2.58054
R51719 a_33249_48695.n122 a_33249_48695.n121 2.58054
R51720 a_33249_48695.n94 a_33249_48695.n93 2.58054
R51721 a_33249_48695.n167 a_33249_48695.n166 2.58054
R51722 a_33249_48695.n162 a_33249_48695.n161 2.58054
R51723 a_33249_48695.n154 a_33249_48695.n153 2.58054
R51724 a_33249_48695.n145 a_33249_48695.n144 2.58054
R51725 a_33249_48695.n127 a_33249_48695.n125 2.53418
R51726 a_33249_48695.n104 a_33249_48695.n102 2.53418
R51727 a_33249_48695.n151 a_33249_48695.n149 2.53418
R51728 a_33249_48695.n172 a_33249_48695.n170 2.53418
R51729 a_33249_48695.n397 a_33249_48695.n48 2.52471
R51730 a_33249_48695.n70 a_33249_48695.n69 2.52436
R51731 a_33249_48695.n375 a_33249_48695.n374 2.52436
R51732 a_33249_48695.n62 a_33249_48695.n61 2.52436
R51733 a_33249_48695.n135 a_33249_48695.n134 2.51873
R51734 a_33249_48695.n335 a_33249_48695.n328 2.46014
R51735 a_33249_48695.n296 a_33249_48695.n285 2.46014
R51736 a_33249_48695.n99 a_33249_48695.n97 2.40765
R51737 a_33249_48695.n114 a_33249_48695.n112 2.40765
R51738 a_33249_48695.n122 a_33249_48695.n120 2.40765
R51739 a_33249_48695.n94 a_33249_48695.n92 2.40765
R51740 a_33249_48695.n167 a_33249_48695.n165 2.40765
R51741 a_33249_48695.n162 a_33249_48695.n160 2.40765
R51742 a_33249_48695.n154 a_33249_48695.n152 2.40765
R51743 a_33249_48695.n145 a_33249_48695.n143 2.40765
R51744 a_33249_48695.n299 a_33249_48695.n298 2.39107
R51745 a_33249_48695.n283 a_33249_48695.n282 2.39107
R51746 a_33249_48695.n333 a_33249_48695.n332 2.39107
R51747 a_33249_48695.n326 a_33249_48695.n325 2.39107
R51748 a_33249_48695.n227 a_33249_48695.n23 2.37644
R51749 a_33249_48695.n183 a_33249_48695.n20 2.37644
R51750 a_33249_48695.n110 a_33249_48695.n109 2.23844
R51751 a_33249_48695.n390 a_33249_48695.n388 2.21818
R51752 a_33249_48695.n55 a_33249_48695.n53 2.21818
R51753 a_33249_48695.n360 a_33249_48695.n358 2.21818
R51754 a_33249_48695.n356 a_33249_48695.n354 2.21818
R51755 a_33249_48695.n231 a_33249_48695.n230 2.2016
R51756 a_33249_48695.n234 a_33249_48695.n233 2.2016
R51757 a_33249_48695.n238 a_33249_48695.n237 2.2016
R51758 a_33249_48695.n242 a_33249_48695.n241 2.2016
R51759 a_33249_48695.n247 a_33249_48695.n246 2.2016
R51760 a_33249_48695.n251 a_33249_48695.n250 2.2016
R51761 a_33249_48695.n255 a_33249_48695.n254 2.2016
R51762 a_33249_48695.n259 a_33249_48695.n258 2.2016
R51763 a_33249_48695.n204 a_33249_48695.n203 2.2016
R51764 a_33249_48695.n207 a_33249_48695.n206 2.2016
R51765 a_33249_48695.n211 a_33249_48695.n210 2.2016
R51766 a_33249_48695.n215 a_33249_48695.n214 2.2016
R51767 a_33249_48695.n200 a_33249_48695.n199 2.2016
R51768 a_33249_48695.n196 a_33249_48695.n195 2.2016
R51769 a_33249_48695.n192 a_33249_48695.n191 2.2016
R51770 a_33249_48695.n188 a_33249_48695.n187 2.2016
R51771 a_33249_48695.n396 a_33249_48695.n395 2.13841
R51772 a_33249_48695.n387 a_33249_48695.n65 2.13841
R51773 a_33249_48695.n218 a_33249_48695.n183 2.0852
R51774 a_33249_48695.n295 a_33249_48695.n294 2.0852
R51775 a_33249_48695.n348 a_33249_48695.n347 1.95191
R51776 a_33249_48695.n262 a_33249_48695.n178 1.90397
R51777 a_33249_48695.n348 a_33249_48695.n76 1.80854
R51778 a_33249_48695.n178 a_33249_48695.n71 1.80603
R51779 a_33249_48695.n394 a_33249_48695.n56 1.73904
R51780 a_33249_48695.n364 a_33249_48695.n357 1.73904
R51781 a_33249_48695.n347 a_33249_48695.n346 1.73609
R51782 a_33249_48695.n320 a_33249_48695.n319 1.73609
R51783 a_33249_48695.n261 a_33249_48695.n260 1.65018
R51784 a_33249_48695.n189 a_33249_48695.n185 1.65018
R51785 a_33249_48695.n271 a_33249_48695.n270 1.56167
R51786 a_33249_48695.n132 a_33249_48695.n29 1.65553
R51787 a_33249_48695.n176 a_33249_48695.n26 1.65553
R51788 a_33249_48695.n352 a_33249_48695.n351 1.5005
R51789 a_33249_48695.n365 a_33249_48695.n364 1.5005
R51790 a_33249_48695.n367 a_33249_48695.n366 1.5005
R51791 a_33249_48695.n381 a_33249_48695.n51 1.5005
R51792 a_33249_48695.n395 a_33249_48695.n394 1.5005
R51793 a_33249_48695.n225 a_33249_48695.n224 1.5005
R51794 a_33249_48695.n227 a_33249_48695.n226 1.5005
R51795 a_33249_48695.n269 a_33249_48695.n268 1.5005
R51796 a_33249_48695.n218 a_33249_48695.n217 1.5005
R51797 a_33249_48695.n244 a_33249_48695.n85 1.5005
R51798 a_33249_48695.n147 a_33249_48695.n86 1.5005
R51799 a_33249_48695.n129 a_33249_48695.n128 1.5005
R51800 a_33249_48695.n176 a_33249_48695.n175 1.5005
R51801 a_33249_48695.n174 a_33249_48695.n173 1.5005
R51802 a_33249_48695.n141 a_33249_48695.n140 1.5005
R51803 a_33249_48695.n132 a_33249_48695.n89 1.5005
R51804 a_33249_48695.n111 a_33249_48695.n110 1.5005
R51805 a_33249_48695.n336 a_33249_48695.n335 1.5005
R51806 a_33249_48695.n311 a_33249_48695.n272 1.5005
R51807 a_33249_48695.n323 a_33249_48695.n322 1.5005
R51808 a_33249_48695.n338 a_33249_48695.n337 1.5005
R51809 a_33249_48695.n296 a_33249_48695.n295 1.5005
R51810 a_33249_48695.n350 a_33249_48695.n349 1.5005
R51811 a_33249_48695.n379 a_33249_48695.n378 1.5005
R51812 a_33249_48695.n386 a_33249_48695.n385 1.5005
R51813 a_33249_48695.n63 a_33249_48695.t273 1.4705
R51814 a_33249_48695.n63 a_33249_48695.t213 1.4705
R51815 a_33249_48695.n59 a_33249_48695.t264 1.4705
R51816 a_33249_48695.n59 a_33249_48695.t208 1.4705
R51817 a_33249_48695.n49 a_33249_48695.t258 1.4705
R51818 a_33249_48695.n49 a_33249_48695.t221 1.4705
R51819 a_33249_48695.n46 a_33249_48695.t204 1.4705
R51820 a_33249_48695.n46 a_33249_48695.t324 1.4705
R51821 a_33249_48695.n388 a_33249_48695.t234 1.4705
R51822 a_33249_48695.n388 a_33249_48695.t159 1.4705
R51823 a_33249_48695.n389 a_33249_48695.t275 1.4705
R51824 a_33249_48695.n389 a_33249_48695.t200 1.4705
R51825 a_33249_48695.n53 a_33249_48695.t216 1.4705
R51826 a_33249_48695.n53 a_33249_48695.t296 1.4705
R51827 a_33249_48695.n54 a_33249_48695.t260 1.4705
R51828 a_33249_48695.n54 a_33249_48695.t166 1.4705
R51829 a_33249_48695.n384 a_33249_48695.t286 1.4705
R51830 a_33249_48695.n384 a_33249_48695.t228 1.4705
R51831 a_33249_48695.n383 a_33249_48695.t278 1.4705
R51832 a_33249_48695.n383 a_33249_48695.t220 1.4705
R51833 a_33249_48695.n382 a_33249_48695.t268 1.4705
R51834 a_33249_48695.n382 a_33249_48695.t235 1.4705
R51835 a_33249_48695.n380 a_33249_48695.t217 1.4705
R51836 a_33249_48695.n380 a_33249_48695.t161 1.4705
R51837 a_33249_48695.n376 a_33249_48695.t171 1.4705
R51838 a_33249_48695.n376 a_33249_48695.t288 1.4705
R51839 a_33249_48695.n372 a_33249_48695.t164 1.4705
R51840 a_33249_48695.n372 a_33249_48695.t279 1.4705
R51841 a_33249_48695.n368 a_33249_48695.t331 1.4705
R51842 a_33249_48695.n368 a_33249_48695.t293 1.4705
R51843 a_33249_48695.n67 a_33249_48695.t277 1.4705
R51844 a_33249_48695.n67 a_33249_48695.t219 1.4705
R51845 a_33249_48695.n358 a_33249_48695.t307 1.4705
R51846 a_33249_48695.n358 a_33249_48695.t232 1.4705
R51847 a_33249_48695.n359 a_33249_48695.t225 1.4705
R51848 a_33249_48695.n359 a_33249_48695.t329 1.4705
R51849 a_33249_48695.n354 a_33249_48695.t290 1.4705
R51850 a_33249_48695.n354 a_33249_48695.t192 1.4705
R51851 a_33249_48695.n355 a_33249_48695.t210 1.4705
R51852 a_33249_48695.n355 a_33249_48695.t287 1.4705
R51853 a_33249_48695.n75 a_33249_48695.t241 1.4705
R51854 a_33249_48695.n75 a_33249_48695.t179 1.4705
R51855 a_33249_48695.n74 a_33249_48695.t226 1.4705
R51856 a_33249_48695.n74 a_33249_48695.t169 1.4705
R51857 a_33249_48695.n73 a_33249_48695.t222 1.4705
R51858 a_33249_48695.n73 a_33249_48695.t181 1.4705
R51859 a_33249_48695.n72 a_33249_48695.t168 1.4705
R51860 a_33249_48695.n72 a_33249_48695.t283 1.4705
R51861 a_33249_48695.n182 a_33249_48695.t23 1.4705
R51862 a_33249_48695.n182 a_33249_48695.t58 1.4705
R51863 a_33249_48695.n184 a_33249_48695.t31 1.4705
R51864 a_33249_48695.n184 a_33249_48695.t78 1.4705
R51865 a_33249_48695.n229 a_33249_48695.t27 1.4705
R51866 a_33249_48695.n229 a_33249_48695.t45 1.4705
R51867 a_33249_48695.n230 a_33249_48695.t22 1.4705
R51868 a_33249_48695.n230 a_33249_48695.t43 1.4705
R51869 a_33249_48695.n232 a_33249_48695.t26 1.4705
R51870 a_33249_48695.n232 a_33249_48695.t84 1.4705
R51871 a_33249_48695.n233 a_33249_48695.t21 1.4705
R51872 a_33249_48695.n233 a_33249_48695.t80 1.4705
R51873 a_33249_48695.n236 a_33249_48695.t36 1.4705
R51874 a_33249_48695.n236 a_33249_48695.t61 1.4705
R51875 a_33249_48695.n237 a_33249_48695.t25 1.4705
R51876 a_33249_48695.n237 a_33249_48695.t52 1.4705
R51877 a_33249_48695.n240 a_33249_48695.t65 1.4705
R51878 a_33249_48695.n240 a_33249_48695.t90 1.4705
R51879 a_33249_48695.n241 a_33249_48695.t56 1.4705
R51880 a_33249_48695.n241 a_33249_48695.t83 1.4705
R51881 a_33249_48695.n245 a_33249_48695.t24 1.4705
R51882 a_33249_48695.n245 a_33249_48695.t51 1.4705
R51883 a_33249_48695.n246 a_33249_48695.t19 1.4705
R51884 a_33249_48695.n246 a_33249_48695.t46 1.4705
R51885 a_33249_48695.n249 a_33249_48695.t54 1.4705
R51886 a_33249_48695.n249 a_33249_48695.t94 1.4705
R51887 a_33249_48695.n250 a_33249_48695.t50 1.4705
R51888 a_33249_48695.n250 a_33249_48695.t85 1.4705
R51889 a_33249_48695.n253 a_33249_48695.t63 1.4705
R51890 a_33249_48695.n253 a_33249_48695.t86 1.4705
R51891 a_33249_48695.n254 a_33249_48695.t53 1.4705
R51892 a_33249_48695.n254 a_33249_48695.t82 1.4705
R51893 a_33249_48695.n257 a_33249_48695.t15 1.4705
R51894 a_33249_48695.n257 a_33249_48695.t37 1.4705
R51895 a_33249_48695.n258 a_33249_48695.t98 1.4705
R51896 a_33249_48695.n258 a_33249_48695.t28 1.4705
R51897 a_33249_48695.n202 a_33249_48695.t35 1.4705
R51898 a_33249_48695.n202 a_33249_48695.t49 1.4705
R51899 a_33249_48695.n203 a_33249_48695.t33 1.4705
R51900 a_33249_48695.n203 a_33249_48695.t47 1.4705
R51901 a_33249_48695.n205 a_33249_48695.t34 1.4705
R51902 a_33249_48695.n205 a_33249_48695.t89 1.4705
R51903 a_33249_48695.n206 a_33249_48695.t32 1.4705
R51904 a_33249_48695.n206 a_33249_48695.t88 1.4705
R51905 a_33249_48695.n209 a_33249_48695.t40 1.4705
R51906 a_33249_48695.n209 a_33249_48695.t69 1.4705
R51907 a_33249_48695.n210 a_33249_48695.t38 1.4705
R51908 a_33249_48695.n210 a_33249_48695.t66 1.4705
R51909 a_33249_48695.n213 a_33249_48695.t73 1.4705
R51910 a_33249_48695.n213 a_33249_48695.t96 1.4705
R51911 a_33249_48695.n214 a_33249_48695.t72 1.4705
R51912 a_33249_48695.n214 a_33249_48695.t95 1.4705
R51913 a_33249_48695.n198 a_33249_48695.t30 1.4705
R51914 a_33249_48695.n198 a_33249_48695.t57 1.4705
R51915 a_33249_48695.n199 a_33249_48695.t29 1.4705
R51916 a_33249_48695.n199 a_33249_48695.t55 1.4705
R51917 a_33249_48695.n194 a_33249_48695.t62 1.4705
R51918 a_33249_48695.n194 a_33249_48695.t100 1.4705
R51919 a_33249_48695.n195 a_33249_48695.t60 1.4705
R51920 a_33249_48695.n195 a_33249_48695.t99 1.4705
R51921 a_33249_48695.n190 a_33249_48695.t70 1.4705
R51922 a_33249_48695.n190 a_33249_48695.t93 1.4705
R51923 a_33249_48695.n191 a_33249_48695.t68 1.4705
R51924 a_33249_48695.n191 a_33249_48695.t92 1.4705
R51925 a_33249_48695.n186 a_33249_48695.t18 1.4705
R51926 a_33249_48695.n186 a_33249_48695.t41 1.4705
R51927 a_33249_48695.n187 a_33249_48695.t17 1.4705
R51928 a_33249_48695.n187 a_33249_48695.t39 1.4705
R51929 a_33249_48695.n266 a_33249_48695.t64 1.4705
R51930 a_33249_48695.n266 a_33249_48695.t91 1.4705
R51931 a_33249_48695.n263 a_33249_48695.t74 1.4705
R51932 a_33249_48695.n263 a_33249_48695.t101 1.4705
R51933 a_33249_48695.n181 a_33249_48695.t14 1.4705
R51934 a_33249_48695.n181 a_33249_48695.t48 1.4705
R51935 a_33249_48695.n180 a_33249_48695.t20 1.4705
R51936 a_33249_48695.n180 a_33249_48695.t75 1.4705
R51937 a_33249_48695.n222 a_33249_48695.t71 1.4705
R51938 a_33249_48695.n222 a_33249_48695.t97 1.4705
R51939 a_33249_48695.n219 a_33249_48695.t77 1.4705
R51940 a_33249_48695.n219 a_33249_48695.t16 1.4705
R51941 a_33249_48695.n88 a_33249_48695.t267 1.4705
R51942 a_33249_48695.n88 a_33249_48695.t211 1.4705
R51943 a_33249_48695.n87 a_33249_48695.t255 1.4705
R51944 a_33249_48695.n87 a_33249_48695.t195 1.4705
R51945 a_33249_48695.n107 a_33249_48695.t250 1.4705
R51946 a_33249_48695.n107 a_33249_48695.t174 1.4705
R51947 a_33249_48695.n105 a_33249_48695.t233 1.4705
R51948 a_33249_48695.n105 a_33249_48695.t312 1.4705
R51949 a_33249_48695.n97 a_33249_48695.t259 1.4705
R51950 a_33249_48695.n97 a_33249_48695.t197 1.4705
R51951 a_33249_48695.n98 a_33249_48695.t303 1.4705
R51952 a_33249_48695.n98 a_33249_48695.t245 1.4705
R51953 a_33249_48695.n112 a_33249_48695.t252 1.4705
R51954 a_33249_48695.n112 a_33249_48695.t191 1.4705
R51955 a_33249_48695.n113 a_33249_48695.t294 1.4705
R51956 a_33249_48695.n113 a_33249_48695.t238 1.4705
R51957 a_33249_48695.n120 a_33249_48695.t243 1.4705
R51958 a_33249_48695.n120 a_33249_48695.t203 1.4705
R51959 a_33249_48695.n121 a_33249_48695.t285 1.4705
R51960 a_33249_48695.n121 a_33249_48695.t251 1.4705
R51961 a_33249_48695.n92 a_33249_48695.t188 1.4705
R51962 a_33249_48695.n92 a_33249_48695.t309 1.4705
R51963 a_33249_48695.n93 a_33249_48695.t236 1.4705
R51964 a_33249_48695.n93 a_33249_48695.t176 1.4705
R51965 a_33249_48695.n131 a_33249_48695.t321 1.4705
R51966 a_33249_48695.n131 a_33249_48695.t261 1.4705
R51967 a_33249_48695.n130 a_33249_48695.t305 1.4705
R51968 a_33249_48695.n130 a_33249_48695.t247 1.4705
R51969 a_33249_48695.n138 a_33249_48695.t322 1.4705
R51970 a_33249_48695.n138 a_33249_48695.t249 1.4705
R51971 a_33249_48695.n136 a_33249_48695.t306 1.4705
R51972 a_33249_48695.n136 a_33249_48695.t209 1.4705
R51973 a_33249_48695.n165 a_33249_48695.t332 1.4705
R51974 a_33249_48695.n165 a_33249_48695.t271 1.4705
R51975 a_33249_48695.n166 a_33249_48695.t254 1.4705
R51976 a_33249_48695.n166 a_33249_48695.t193 1.4705
R51977 a_33249_48695.n160 a_33249_48695.t325 1.4705
R51978 a_33249_48695.n160 a_33249_48695.t263 1.4705
R51979 a_33249_48695.n161 a_33249_48695.t242 1.4705
R51980 a_33249_48695.n161 a_33249_48695.t183 1.4705
R51981 a_33249_48695.n152 a_33249_48695.t316 1.4705
R51982 a_33249_48695.n152 a_33249_48695.t276 1.4705
R51983 a_33249_48695.n153 a_33249_48695.t240 1.4705
R51984 a_33249_48695.n153 a_33249_48695.t196 1.4705
R51985 a_33249_48695.n143 a_33249_48695.t262 1.4705
R51986 a_33249_48695.n143 a_33249_48695.t202 1.4705
R51987 a_33249_48695.n144 a_33249_48695.t182 1.4705
R51988 a_33249_48695.n144 a_33249_48695.t300 1.4705
R51989 a_33249_48695.n297 a_33249_48695.t134 1.4705
R51990 a_33249_48695.n297 a_33249_48695.t347 1.4705
R51991 a_33249_48695.n298 a_33249_48695.t133 1.4705
R51992 a_33249_48695.n298 a_33249_48695.t346 1.4705
R51993 a_33249_48695.n281 a_33249_48695.t140 1.4705
R51994 a_33249_48695.n281 a_33249_48695.t0 1.4705
R51995 a_33249_48695.n282 a_33249_48695.t139 1.4705
R51996 a_33249_48695.n282 a_33249_48695.t158 1.4705
R51997 a_33249_48695.n345 a_33249_48695.t110 1.4705
R51998 a_33249_48695.n345 a_33249_48695.t104 1.4705
R51999 a_33249_48695.n343 a_33249_48695.t109 1.4705
R52000 a_33249_48695.n343 a_33249_48695.t137 1.4705
R52001 a_33249_48695.n341 a_33249_48695.t6 1.4705
R52002 a_33249_48695.n341 a_33249_48695.t341 1.4705
R52003 a_33249_48695.n339 a_33249_48695.t344 1.4705
R52004 a_33249_48695.n339 a_33249_48695.t142 1.4705
R52005 a_33249_48695.n83 a_33249_48695.t8 1.4705
R52006 a_33249_48695.n83 a_33249_48695.t13 1.4705
R52007 a_33249_48695.n81 a_33249_48695.t337 1.4705
R52008 a_33249_48695.n81 a_33249_48695.t144 1.4705
R52009 a_33249_48695.n79 a_33249_48695.t343 1.4705
R52010 a_33249_48695.n79 a_33249_48695.t138 1.4705
R52011 a_33249_48695.n78 a_33249_48695.t151 1.4705
R52012 a_33249_48695.n78 a_33249_48695.t106 1.4705
R52013 a_33249_48695.n280 a_33249_48695.t4 1.4705
R52014 a_33249_48695.n280 a_33249_48695.t336 1.4705
R52015 a_33249_48695.n279 a_33249_48695.t3 1.4705
R52016 a_33249_48695.n279 a_33249_48695.t146 1.4705
R52017 a_33249_48695.n278 a_33249_48695.t111 1.4705
R52018 a_33249_48695.n278 a_33249_48695.t120 1.4705
R52019 a_33249_48695.n277 a_33249_48695.t124 1.4705
R52020 a_33249_48695.n277 a_33249_48695.t149 1.4705
R52021 a_33249_48695.n276 a_33249_48695.t107 1.4705
R52022 a_33249_48695.n276 a_33249_48695.t345 1.4705
R52023 a_33249_48695.n275 a_33249_48695.t117 1.4705
R52024 a_33249_48695.n275 a_33249_48695.t152 1.4705
R52025 a_33249_48695.n274 a_33249_48695.t121 1.4705
R52026 a_33249_48695.n274 a_33249_48695.t148 1.4705
R52027 a_33249_48695.n273 a_33249_48695.t348 1.4705
R52028 a_33249_48695.n273 a_33249_48695.t112 1.4705
R52029 a_33249_48695.n318 a_33249_48695.t5 1.4705
R52030 a_33249_48695.n318 a_33249_48695.t11 1.4705
R52031 a_33249_48695.n316 a_33249_48695.t1 1.4705
R52032 a_33249_48695.n316 a_33249_48695.t141 1.4705
R52033 a_33249_48695.n314 a_33249_48695.t108 1.4705
R52034 a_33249_48695.n314 a_33249_48695.t115 1.4705
R52035 a_33249_48695.n312 a_33249_48695.t118 1.4705
R52036 a_33249_48695.n312 a_33249_48695.t145 1.4705
R52037 a_33249_48695.n309 a_33249_48695.t157 1.4705
R52038 a_33249_48695.n309 a_33249_48695.t338 1.4705
R52039 a_33249_48695.n307 a_33249_48695.t342 1.4705
R52040 a_33249_48695.n307 a_33249_48695.t147 1.4705
R52041 a_33249_48695.n305 a_33249_48695.t116 1.4705
R52042 a_33249_48695.n305 a_33249_48695.t143 1.4705
R52043 a_33249_48695.n304 a_33249_48695.t154 1.4705
R52044 a_33249_48695.n304 a_33249_48695.t2 1.4705
R52045 a_33249_48695.n293 a_33249_48695.t103 1.4705
R52046 a_33249_48695.n293 a_33249_48695.t114 1.4705
R52047 a_33249_48695.n292 a_33249_48695.t102 1.4705
R52048 a_33249_48695.n292 a_33249_48695.t153 1.4705
R52049 a_33249_48695.n291 a_33249_48695.t10 1.4705
R52050 a_33249_48695.n291 a_33249_48695.t129 1.4705
R52051 a_33249_48695.n290 a_33249_48695.t135 1.4705
R52052 a_33249_48695.n290 a_33249_48695.t351 1.4705
R52053 a_33249_48695.n289 a_33249_48695.t113 1.4705
R52054 a_33249_48695.n289 a_33249_48695.t123 1.4705
R52055 a_33249_48695.n288 a_33249_48695.t126 1.4705
R52056 a_33249_48695.n288 a_33249_48695.t349 1.4705
R52057 a_33249_48695.n287 a_33249_48695.t132 1.4705
R52058 a_33249_48695.n287 a_33249_48695.t156 1.4705
R52059 a_33249_48695.n286 a_33249_48695.t7 1.4705
R52060 a_33249_48695.n286 a_33249_48695.t12 1.4705
R52061 a_33249_48695.n331 a_33249_48695.t127 1.4705
R52062 a_33249_48695.n331 a_33249_48695.t155 1.4705
R52063 a_33249_48695.n332 a_33249_48695.t122 1.4705
R52064 a_33249_48695.n332 a_33249_48695.t150 1.4705
R52065 a_33249_48695.n324 a_33249_48695.t136 1.4705
R52066 a_33249_48695.n324 a_33249_48695.t9 1.4705
R52067 a_33249_48695.n325 a_33249_48695.t131 1.4705
R52068 a_33249_48695.n325 a_33249_48695.t350 1.4705
R52069 a_33249_48695.n391 a_33249_48695.n390 1.46537
R52070 a_33249_48695.n393 a_33249_48695.n392 1.46537
R52071 a_33249_48695.n56 a_33249_48695.n55 1.46537
R52072 a_33249_48695.n361 a_33249_48695.n360 1.46537
R52073 a_33249_48695.n363 a_33249_48695.n362 1.46537
R52074 a_33249_48695.n357 a_33249_48695.n356 1.46537
R52075 a_33249_48695.n100 a_33249_48695.n99 1.46537
R52076 a_33249_48695.n102 a_33249_48695.n101 1.46537
R52077 a_33249_48695.n115 a_33249_48695.n114 1.46537
R52078 a_33249_48695.n117 a_33249_48695.n116 1.46537
R52079 a_33249_48695.n119 a_33249_48695.n118 1.46537
R52080 a_33249_48695.n123 a_33249_48695.n122 1.46537
R52081 a_33249_48695.n125 a_33249_48695.n124 1.46537
R52082 a_33249_48695.n95 a_33249_48695.n94 1.46537
R52083 a_33249_48695.n168 a_33249_48695.n167 1.46537
R52084 a_33249_48695.n170 a_33249_48695.n169 1.46537
R52085 a_33249_48695.n163 a_33249_48695.n162 1.46537
R52086 a_33249_48695.n159 a_33249_48695.n158 1.46537
R52087 a_33249_48695.n157 a_33249_48695.n156 1.46537
R52088 a_33249_48695.n155 a_33249_48695.n154 1.46537
R52089 a_33249_48695.n151 a_33249_48695.n150 1.46537
R52090 a_33249_48695.n146 a_33249_48695.n145 1.46537
R52091 a_33249_48695.n302 a_33249_48695.n301 1.46537
R52092 a_33249_48695.n300 a_33249_48695.n299 1.46537
R52093 a_33249_48695.n285 a_33249_48695.n284 1.46537
R52094 a_33249_48695.n330 a_33249_48695.n329 1.46537
R52095 a_33249_48695.n334 a_33249_48695.n333 1.46537
R52096 a_33249_48695.n328 a_33249_48695.n327 1.46537
R52097 a_33249_48695.n235 a_33249_48695.n234 1.46537
R52098 a_33249_48695.n239 a_33249_48695.n238 1.46537
R52099 a_33249_48695.n243 a_33249_48695.n242 1.46537
R52100 a_33249_48695.n248 a_33249_48695.n247 1.46537
R52101 a_33249_48695.n252 a_33249_48695.n251 1.46537
R52102 a_33249_48695.n256 a_33249_48695.n255 1.46537
R52103 a_33249_48695.n260 a_33249_48695.n259 1.46537
R52104 a_33249_48695.n208 a_33249_48695.n207 1.46537
R52105 a_33249_48695.n212 a_33249_48695.n211 1.46537
R52106 a_33249_48695.n216 a_33249_48695.n215 1.46537
R52107 a_33249_48695.n201 a_33249_48695.n200 1.46537
R52108 a_33249_48695.n197 a_33249_48695.n196 1.46537
R52109 a_33249_48695.n193 a_33249_48695.n192 1.46537
R52110 a_33249_48695.n189 a_33249_48695.n188 1.46537
R52111 a_33249_48695.n104 a_33249_48695.n103 1.46535
R52112 a_33249_48695.n127 a_33249_48695.n126 1.46535
R52113 a_33249_48695.n172 a_33249_48695.n171 1.46535
R52114 a_33249_48695.n149 a_33249_48695.n148 1.46535
R52115 a_33249_48695.n337 a_33249_48695.n271 1.34705
R52116 a_33249_48695.n270 a_33249_48695.n269 1.2981
R52117 a_33249_48695.n175 a_33249_48695.n76 1.27763
R52118 a_33249_48695.n393 a_33249_48695.n391 1.27228
R52119 a_33249_48695.n370 a_33249_48695.n369 1.27228
R52120 a_33249_48695.n373 a_33249_48695.n371 1.27228
R52121 a_33249_48695.n363 a_33249_48695.n361 1.27228
R52122 a_33249_48695.n106 a_33249_48695.n90 1.27228
R52123 a_33249_48695.n125 a_33249_48695.n123 1.27228
R52124 a_33249_48695.n123 a_33249_48695.n119 1.27228
R52125 a_33249_48695.n117 a_33249_48695.n115 1.27228
R52126 a_33249_48695.n102 a_33249_48695.n100 1.27228
R52127 a_33249_48695.n137 a_33249_48695.n135 1.27228
R52128 a_33249_48695.n155 a_33249_48695.n151 1.27228
R52129 a_33249_48695.n157 a_33249_48695.n155 1.27228
R52130 a_33249_48695.n163 a_33249_48695.n159 1.27228
R52131 a_33249_48695.n170 a_33249_48695.n168 1.27228
R52132 a_33249_48695.n57 a_33249_48695.n50 1.27228
R52133 a_33249_48695.n60 a_33249_48695.n58 1.27228
R52134 a_33249_48695.n260 a_33249_48695.n256 1.27228
R52135 a_33249_48695.n252 a_33249_48695.n248 1.27228
R52136 a_33249_48695.n243 a_33249_48695.n239 1.27228
R52137 a_33249_48695.n193 a_33249_48695.n189 1.27228
R52138 a_33249_48695.n201 a_33249_48695.n197 1.27228
R52139 a_33249_48695.n216 a_33249_48695.n212 1.27228
R52140 a_33249_48695.n265 a_33249_48695.n264 1.27228
R52141 a_33249_48695.n221 a_33249_48695.n220 1.27228
R52142 a_33249_48695.n84 a_33249_48695.n82 1.27228
R52143 a_33249_48695.n342 a_33249_48695.n340 1.27228
R52144 a_33249_48695.n346 a_33249_48695.n344 1.27228
R52145 a_33249_48695.n310 a_33249_48695.n308 1.27228
R52146 a_33249_48695.n315 a_33249_48695.n313 1.27228
R52147 a_33249_48695.n319 a_33249_48695.n317 1.27228
R52148 a_33249_48695.n334 a_33249_48695.n330 1.27228
R52149 a_33249_48695.n302 a_33249_48695.n300 1.27228
R52150 a_33249_48695.n69 a_33249_48695.n68 1.26756
R52151 a_33249_48695.n374 a_33249_48695.n373 1.26756
R52152 a_33249_48695.n48 a_33249_48695.n47 1.26756
R52153 a_33249_48695.n61 a_33249_48695.n60 1.26756
R52154 a_33249_48695.n349 a_33249_48695.n348 1.23567
R52155 a_33249_48695.n352 a_33249_48695.n71 1.23455
R52156 a_33249_48695.n178 a_33249_48695.n177 1.18682
R52157 a_33249_48695.n109 a_33249_48695.n108 1.01873
R52158 a_33249_48695.n140 a_33249_48695.n139 1.01873
R52159 a_33249_48695.n323 a_33249_48695.n272 0.822966
R52160 a_33249_48695.n321 a_33249_48695.n320 0.822966
R52161 a_33249_48695.n367 a_33249_48695.n70 0.796291
R52162 a_33249_48695.n378 a_33249_48695.n375 0.796291
R52163 a_33249_48695.n65 a_33249_48695.n62 0.796291
R52164 a_33249_48695.n397 a_33249_48695.n396 0.795934
R52165 a_33249_48695.n395 a_33249_48695.n51 0.780703
R52166 a_33249_48695.n365 a_33249_48695.n352 0.780703
R52167 a_33249_48695.n387 a_33249_48695.n386 0.780703
R52168 a_33249_48695.n349 a_33249_48695.n66 0.780703
R52169 a_33249_48695.n133 a_33249_48695.n129 0.778574
R52170 a_33249_48695.n177 a_33249_48695.n86 0.778574
R52171 a_33249_48695.n110 a_33249_48695.n89 0.778574
R52172 a_33249_48695.n175 a_33249_48695.n174 0.778574
R52173 a_33249_48695.n134 a_33249_48695.n86 0.738439
R52174 a_33249_48695.n174 a_33249_48695.n141 0.738439
R52175 a_33249_48695.n262 a_33249_48695.n261 0.737223
R52176 a_33249_48695.n185 a_33249_48695.n179 0.737223
R52177 a_33249_48695.n269 a_33249_48695.n85 0.737223
R52178 a_33249_48695.n225 a_33249_48695.n218 0.737223
R52179 a_33249_48695.n228 a_33249_48695.n179 0.725061
R52180 a_33249_48695.n226 a_33249_48695.n225 0.725061
R52181 a_33249_48695.n128 a_33249_48695.n127 0.699581
R52182 a_33249_48695.n111 a_33249_48695.n104 0.699581
R52183 a_33249_48695.n149 a_33249_48695.n147 0.699581
R52184 a_33249_48695.n173 a_33249_48695.n172 0.699581
R52185 a_33249_48695.n337 a_33249_48695.n336 0.639318
R52186 a_33249_48695.n295 a_33249_48695.n272 0.639318
R52187 a_33249_48695.n347 a_33249_48695.n77 0.639318
R52188 a_33249_48695.n320 a_33249_48695.n303 0.639318
R52189 a_33249_48695.n366 a_33249_48695.n365 0.638405
R52190 a_33249_48695.n379 a_33249_48695.n66 0.638405
R52191 a_33249_48695.n366 a_33249_48695.n51 0.628372
R52192 a_33249_48695.n386 a_33249_48695.n379 0.628372
R52193 a_33249_48695.n271 a_33249_48695.n71 0.606869
R52194 a_33249_48695.n270 a_33249_48695.n76 0.60536
R52195 a_33249_48695.n261 a_33249_48695.n228 0.585196
R52196 a_33249_48695.n226 a_33249_48695.n85 0.585196
R52197 a_33249_48695.n336 a_33249_48695.n323 0.585196
R52198 a_33249_48695.n321 a_33249_48695.n77 0.585196
R52199 a_33249_48695.n128 a_33249_48695.n95 0.557791
R52200 a_33249_48695.n115 a_33249_48695.n111 0.557791
R52201 a_33249_48695.n147 a_33249_48695.n146 0.557791
R52202 a_33249_48695.n173 a_33249_48695.n163 0.557791
R52203 a_33249_48695.n134 a_33249_48695.n133 0.530466
R52204 a_33249_48695.n141 a_33249_48695.n89 0.530466
R52205 a_33249_48695.n369 a_33249_48695.n367 0.476484
R52206 a_33249_48695.n378 a_33249_48695.n377 0.476484
R52207 a_33249_48695.n396 a_33249_48695.n50 0.476484
R52208 a_33249_48695.n65 a_33249_48695.n64 0.476484
R52209 a_33249_48695.n6 a_33249_48695.n381 0.478684
R52210 a_33249_48695.n385 a_33249_48695.n0 0.478684
R52211 a_33249_48695.n351 a_33249_48695.n16 0.478684
R52212 a_33249_48695.n350 a_33249_48695.n10 0.478684
R52213 a_33249_48695.n338 a_33249_48695.n84 0.236091
R52214 a_33249_48695.n311 a_33249_48695.n310 0.236091
R52215 a_33249_48695.n244 a_33249_48695.n243 0.150184
R52216 a_33249_48695.n217 a_33249_48695.n216 0.150184
R52217 a_33249_48695.n8 a_33249_48695.n9 1.27228
R52218 a_33249_48695.n7 a_33249_48695.n8 2.51878
R52219 a_33249_48695.n381 a_33249_48695.n7 0.794091
R52220 a_33249_48695.n5 a_33249_48695.n6 1.27228
R52221 a_33249_48695.n4 a_33249_48695.n5 2.60203
R52222 a_33249_48695.n3 a_33249_48695.n4 1.27228
R52223 a_33249_48695.n2 a_33249_48695.n3 1.27228
R52224 a_33249_48695.n1 a_33249_48695.n2 2.51878
R52225 a_33249_48695.n385 a_33249_48695.n1 0.794091
R52226 a_33249_48695.t190 a_33249_48695.n0 6.77266
R52227 a_33249_48695.n18 a_33249_48695.n19 1.27228
R52228 a_33249_48695.n17 a_33249_48695.n18 2.51878
R52229 a_33249_48695.n351 a_33249_48695.n17 0.794091
R52230 a_33249_48695.n15 a_33249_48695.n16 1.27228
R52231 a_33249_48695.n14 a_33249_48695.n15 2.60203
R52232 a_33249_48695.n13 a_33249_48695.n14 1.27228
R52233 a_33249_48695.n12 a_33249_48695.n13 1.27228
R52234 a_33249_48695.n11 a_33249_48695.n12 2.51878
R52235 a_33249_48695.n350 a_33249_48695.n11 0.794091
R52236 a_33249_48695.t315 a_33249_48695.n10 6.77266
R52237 a_33249_48695.n24 a_33249_48695.n25 1.26457
R52238 a_33249_48695.n227 a_33249_48695.n24 6.59229
R52239 a_33249_48695.n181 a_33249_48695.n23 5.10549
R52240 a_33249_48695.n21 a_33249_48695.n22 1.26457
R52241 a_33249_48695.n183 a_33249_48695.n21 6.59229
R52242 a_33249_48695.n182 a_33249_48695.n20 5.10549
R52243 a_33249_48695.n30 a_33249_48695.n31 1.27228
R52244 a_33249_48695.n132 a_33249_48695.n30 7.30549
R52245 a_33249_48695.t185 a_33249_48695.n29 6.96214
R52246 a_33249_48695.n27 a_33249_48695.n28 1.27228
R52247 a_33249_48695.n176 a_33249_48695.n27 7.30549
R52248 a_33249_48695.t313 a_33249_48695.n26 6.96214
R52249 a_33249_48695.n37 a_33249_48695.n38 3.79678
R52250 a_33249_48695.n36 a_33249_48695.n37 1.27228
R52251 a_33249_48695.n322 a_33249_48695.n36 0.238291
R52252 a_33249_48695.n34 a_33249_48695.n35 1.27228
R52253 a_33249_48695.n33 a_33249_48695.n34 3.79678
R52254 a_33249_48695.n32 a_33249_48695.n33 1.27228
R52255 a_33249_48695.n321 a_33249_48695.n32 1.73829
R52256 a_33249_48695.n44 a_33249_48695.n45 3.79678
R52257 a_33249_48695.n43 a_33249_48695.n44 1.27228
R52258 a_33249_48695.n294 a_33249_48695.n43 0.238291
R52259 a_33249_48695.n41 a_33249_48695.n42 1.27228
R52260 a_33249_48695.n40 a_33249_48695.n41 3.79678
R52261 a_33249_48695.n39 a_33249_48695.n40 1.27228
R52262 a_33249_48695.n39 a_33249_48695.n303 2.32299
R52263 OUT.n14 OUT.n13 12.1937
R52264 OUT.n13 OUT.t0 11.5094
R52265 OUT.n13 OUT.t1 9.24966
R52266 OUT.n27 OUT.n20 7.94229
R52267 OUT.n80 OUT.n78 7.94229
R52268 OUT.n117 OUT.n14 7.76579
R52269 OUT.n75 OUT.n68 7.169
R52270 OUT.n142 OUT.n141 7.169
R52271 OUT.n121 OUT.t4 6.96668
R52272 OUT.n8 OUT.t81 6.82564
R52273 OUT.n72 OUT.t92 6.82564
R52274 OUT.n14 OUT.n12 6.28314
R52275 OUT.n137 OUT.t18 5.85326
R52276 OUT.n137 OUT.n136 5.84661
R52277 OUT.n19 OUT.t93 5.69423
R52278 OUT.n28 OUT.t68 5.69423
R52279 OUT.n17 OUT.t85 5.69423
R52280 OUT.n81 OUT.t66 5.69423
R52281 OUT.n19 OUT.n18 5.49558
R52282 OUT.n17 OUT.n16 5.49558
R52283 OUT.n10 OUT.n9 4.61332
R52284 OUT.n144 OUT.n143 4.61332
R52285 OUT.n74 OUT.n73 4.61332
R52286 OUT.n67 OUT.n65 4.61332
R52287 OUT.n63 OUT.n60 4.61332
R52288 OUT.n123 OUT.n122 4.61332
R52289 OUT.n2 OUT.n1 4.61332
R52290 OUT.n9 OUT.n8 4.60571
R52291 OUT.n143 OUT.n142 4.60571
R52292 OUT.n73 OUT.n72 4.60571
R52293 OUT.n68 OUT.n67 4.60571
R52294 OUT.n64 OUT.n63 4.60571
R52295 OUT.n122 OUT.n121 4.60571
R52296 OUT.n145 OUT.n1 4.60571
R52297 OUT.n62 OUT.n59 4.5005
R52298 OUT.n66 OUT.n58 4.5005
R52299 OUT.n71 OUT.n69 4.5005
R52300 OUT.n120 OUT.n118 4.5005
R52301 OUT.n4 OUT.n3 4.5005
R52302 OUT.n7 OUT.n5 4.5005
R52303 OUT.n147 OUT.n146 4.5005
R52304 OUT.n4 OUT.t78 4.22462
R52305 OUT.n66 OUT.t82 4.22462
R52306 OUT.n27 OUT.n26 4.22423
R52307 OUT.n80 OUT.n79 4.22423
R52308 OUT.n130 OUT.t17 4.21195
R52309 OUT.n132 OUT.t2 4.21195
R52310 OUT.n47 OUT.t41 4.05054
R52311 OUT.n52 OUT.t39 4.05054
R52312 OUT.n54 OUT.t38 4.05054
R52313 OUT.n41 OUT.t100 4.05054
R52314 OUT.n39 OUT.t34 4.05054
R52315 OUT.n33 OUT.t27 4.05054
R52316 OUT.n31 OUT.t79 4.05054
R52317 OUT.n21 OUT.t107 4.05054
R52318 OUT.n88 OUT.t32 4.05054
R52319 OUT.n93 OUT.t25 4.05054
R52320 OUT.n95 OUT.t21 4.05054
R52321 OUT.n102 OUT.t84 4.05054
R52322 OUT.n104 OUT.t102 4.05054
R52323 OUT.n110 OUT.t97 4.05054
R52324 OUT.n112 OUT.t74 4.05054
R52325 OUT.n83 OUT.t89 4.05054
R52326 OUT.n130 OUT.t9 4.03668
R52327 OUT.n132 OUT.t11 4.03668
R52328 OUT.n47 OUT.t37 3.87765
R52329 OUT.n52 OUT.t33 3.87765
R52330 OUT.n54 OUT.t29 3.87765
R52331 OUT.n41 OUT.t91 3.87765
R52332 OUT.n39 OUT.t22 3.87765
R52333 OUT.n33 OUT.t104 3.87765
R52334 OUT.n31 OUT.t75 3.87765
R52335 OUT.n21 OUT.t95 3.87765
R52336 OUT.n88 OUT.t30 3.87765
R52337 OUT.n93 OUT.t24 3.87765
R52338 OUT.n95 OUT.t20 3.87765
R52339 OUT.n102 OUT.t83 3.87765
R52340 OUT.n104 OUT.t99 3.87765
R52341 OUT.n110 OUT.t96 3.87765
R52342 OUT.n112 OUT.t73 3.87765
R52343 OUT.n83 OUT.t87 3.87765
R52344 OUT.n135 OUT.n123 3.81532
R52345 OUT.n140 OUT.n139 3.544
R52346 OUT.n29 OUT.n28 3.25667
R52347 OUT.n120 OUT.n119 3.12366
R52348 OUT.n60 OUT.n15 3.01925
R52349 OUT.n116 OUT.n2 3.01925
R52350 OUT.n129 OUT.n128 2.95195
R52351 OUT.n126 OUT.n125 2.95195
R52352 OUT.n129 OUT.n127 2.77668
R52353 OUT.n126 OUT.n124 2.77668
R52354 OUT.n7 OUT.n6 2.75462
R52355 OUT.n71 OUT.n70 2.75462
R52356 OUT.n62 OUT.n61 2.75462
R52357 OUT.n25 OUT.n21 2.73714
R52358 OUT.n87 OUT.n83 2.73714
R52359 OUT.n51 OUT.n47 2.73672
R52360 OUT.n92 OUT.n88 2.73672
R52361 OUT.n131 OUT.n129 2.71872
R52362 OUT.n42 OUT.n40 2.60203
R52363 OUT.n105 OUT.n103 2.60203
R52364 OUT.n50 OUT.n49 2.58054
R52365 OUT.n45 OUT.n44 2.58054
R52366 OUT.n37 OUT.n36 2.58054
R52367 OUT.n24 OUT.n23 2.58054
R52368 OUT.n91 OUT.n90 2.58054
R52369 OUT.n100 OUT.n99 2.58054
R52370 OUT.n108 OUT.n107 2.58054
R52371 OUT.n86 OUT.n85 2.58054
R52372 OUT.n133 OUT.n131 2.56118
R52373 OUT.n138 OUT.n137 2.54573
R52374 OUT.n34 OUT.n32 2.53418
R52375 OUT.n55 OUT.n53 2.53418
R52376 OUT.n113 OUT.n111 2.53418
R52377 OUT.n96 OUT.n94 2.53418
R52378 OUT.n82 OUT.n81 2.51873
R52379 OUT.n50 OUT.n48 2.40765
R52380 OUT.n45 OUT.n43 2.40765
R52381 OUT.n37 OUT.n35 2.40765
R52382 OUT.n24 OUT.n22 2.40765
R52383 OUT.n91 OUT.n89 2.40765
R52384 OUT.n100 OUT.n98 2.40765
R52385 OUT.n108 OUT.n106 2.40765
R52386 OUT.n86 OUT.n84 2.40765
R52387 OUT.n139 OUT.n117 2.25854
R52388 OUT.n57 OUT.n20 2.23844
R52389 OUT OUT.n0 2.05949
R52390 OUT.n134 OUT.n126 2.00466
R52391 OUT.n75 OUT.n74 1.51925
R52392 OUT.n141 OUT.n10 1.51925
R52393 OUT.n115 OUT.n114 1.5005
R52394 OUT.n30 OUT.n29 1.5005
R52395 OUT.n135 OUT.n134 1.5005
R52396 OUT.n97 OUT.n11 1.5005
R52397 OUT.n78 OUT.n77 1.5005
R52398 OUT.n76 OUT.n75 1.5005
R52399 OUT.n57 OUT.n56 1.5005
R52400 OUT.n141 OUT.n140 1.5005
R52401 OUT.n0 OUT.t50 1.4705
R52402 OUT.n0 OUT.t45 1.4705
R52403 OUT.n6 OUT.t76 1.4705
R52404 OUT.n6 OUT.t52 1.4705
R52405 OUT.n18 OUT.t69 1.4705
R52406 OUT.n18 OUT.t26 1.4705
R52407 OUT.n26 OUT.t65 1.4705
R52408 OUT.n26 OUT.t98 1.4705
R52409 OUT.n48 OUT.t72 1.4705
R52410 OUT.n48 OUT.t59 1.4705
R52411 OUT.n49 OUT.t77 1.4705
R52412 OUT.n49 OUT.t64 1.4705
R52413 OUT.n43 OUT.t49 1.4705
R52414 OUT.n43 OUT.t23 1.4705
R52415 OUT.n44 OUT.t57 1.4705
R52416 OUT.n44 OUT.t35 1.4705
R52417 OUT.n35 OUT.t58 1.4705
R52418 OUT.n35 OUT.t36 1.4705
R52419 OUT.n36 OUT.t63 1.4705
R52420 OUT.n36 OUT.t40 1.4705
R52421 OUT.n22 OUT.t44 1.4705
R52422 OUT.n22 OUT.t94 1.4705
R52423 OUT.n23 OUT.t48 1.4705
R52424 OUT.n23 OUT.t106 1.4705
R52425 OUT.n70 OUT.t80 1.4705
R52426 OUT.n70 OUT.t62 1.4705
R52427 OUT.n61 OUT.t61 1.4705
R52428 OUT.n61 OUT.t55 1.4705
R52429 OUT.n16 OUT.t67 1.4705
R52430 OUT.n16 OUT.t105 1.4705
R52431 OUT.n79 OUT.t60 1.4705
R52432 OUT.n79 OUT.t90 1.4705
R52433 OUT.n89 OUT.t70 1.4705
R52434 OUT.n89 OUT.t53 1.4705
R52435 OUT.n90 OUT.t71 1.4705
R52436 OUT.n90 OUT.t56 1.4705
R52437 OUT.n98 OUT.t46 1.4705
R52438 OUT.n98 OUT.t101 1.4705
R52439 OUT.n99 OUT.t47 1.4705
R52440 OUT.n99 OUT.t103 1.4705
R52441 OUT.n106 OUT.t51 1.4705
R52442 OUT.n106 OUT.t28 1.4705
R52443 OUT.n107 OUT.t54 1.4705
R52444 OUT.n107 OUT.t31 1.4705
R52445 OUT.n84 OUT.t42 1.4705
R52446 OUT.n84 OUT.t86 1.4705
R52447 OUT.n85 OUT.t43 1.4705
R52448 OUT.n85 OUT.t88 1.4705
R52449 OUT.n51 OUT.n50 1.46537
R52450 OUT.n53 OUT.n52 1.46537
R52451 OUT.n46 OUT.n45 1.46537
R52452 OUT.n42 OUT.n41 1.46537
R52453 OUT.n40 OUT.n39 1.46537
R52454 OUT.n38 OUT.n37 1.46537
R52455 OUT.n34 OUT.n33 1.46537
R52456 OUT.n25 OUT.n24 1.46537
R52457 OUT.n92 OUT.n91 1.46537
R52458 OUT.n94 OUT.n93 1.46537
R52459 OUT.n101 OUT.n100 1.46537
R52460 OUT.n103 OUT.n102 1.46537
R52461 OUT.n105 OUT.n104 1.46537
R52462 OUT.n109 OUT.n108 1.46537
R52463 OUT.n111 OUT.n110 1.46537
R52464 OUT.n87 OUT.n86 1.46537
R52465 OUT.n131 OUT.n130 1.46537
R52466 OUT.n55 OUT.n54 1.46535
R52467 OUT.n32 OUT.n31 1.46535
R52468 OUT.n96 OUT.n95 1.46535
R52469 OUT.n113 OUT.n112 1.46535
R52470 OUT.n133 OUT.n132 1.46535
R52471 OUT.n28 OUT.n27 1.27228
R52472 OUT.n38 OUT.n34 1.27228
R52473 OUT.n40 OUT.n38 1.27228
R52474 OUT.n46 OUT.n42 1.27228
R52475 OUT.n53 OUT.n51 1.27228
R52476 OUT.n81 OUT.n80 1.27228
R52477 OUT.n111 OUT.n109 1.27228
R52478 OUT.n109 OUT.n105 1.27228
R52479 OUT.n103 OUT.n101 1.27228
R52480 OUT.n94 OUT.n92 1.27228
R52481 OUT.n136 OUT.t5 1.2605
R52482 OUT.n136 OUT.t12 1.2605
R52483 OUT.n127 OUT.t7 1.2605
R52484 OUT.n127 OUT.t13 1.2605
R52485 OUT.n128 OUT.t15 1.2605
R52486 OUT.n128 OUT.t3 1.2605
R52487 OUT.n124 OUT.t19 1.2605
R52488 OUT.n124 OUT.t6 1.2605
R52489 OUT.n125 OUT.t8 1.2605
R52490 OUT.n125 OUT.t14 1.2605
R52491 OUT.n119 OUT.t10 1.2605
R52492 OUT.n119 OUT.t16 1.2605
R52493 OUT.n139 OUT.n138 1.25797
R52494 OUT.n117 OUT.n116 1.22361
R52495 OUT.n20 OUT.n19 1.01873
R52496 OUT.n78 OUT.n17 1.01873
R52497 OUT.n65 OUT.n64 0.9995
R52498 OUT.n145 OUT.n144 0.9995
R52499 OUT.n29 OUT.n15 0.778574
R52500 OUT.n116 OUT.n115 0.778574
R52501 OUT.n76 OUT.n57 0.778574
R52502 OUT.n140 OUT.n11 0.778574
R52503 OUT.n115 OUT.n82 0.738439
R52504 OUT.n138 OUT.n135 0.738439
R52505 OUT.n77 OUT.n11 0.738439
R52506 OUT.n32 OUT.n30 0.699581
R52507 OUT.n56 OUT.n55 0.699581
R52508 OUT.n114 OUT.n113 0.699581
R52509 OUT.n97 OUT.n96 0.699581
R52510 OUT.n134 OUT.n133 0.699581
R52511 OUT OUT.n147 0.695632
R52512 OUT.n30 OUT.n25 0.557791
R52513 OUT.n56 OUT.n46 0.557791
R52514 OUT.n114 OUT.n87 0.557791
R52515 OUT.n101 OUT.n97 0.557791
R52516 OUT.n82 OUT.n15 0.530466
R52517 OUT.n77 OUT.n76 0.530466
R52518 OUT.n60 OUT.n59 0.14
R52519 OUT.n64 OUT.n59 0.14
R52520 OUT.n65 OUT.n58 0.14
R52521 OUT.n68 OUT.n58 0.14
R52522 OUT.n74 OUT.n69 0.14
R52523 OUT.n72 OUT.n69 0.14
R52524 OUT.n123 OUT.n118 0.14
R52525 OUT.n121 OUT.n118 0.14
R52526 OUT.n146 OUT.n2 0.14
R52527 OUT.n146 OUT.n145 0.14
R52528 OUT.n144 OUT.n3 0.14
R52529 OUT.n142 OUT.n3 0.14
R52530 OUT.n10 OUT.n5 0.14
R52531 OUT.n8 OUT.n5 0.14
R52532 OUT.n12 OUT.t109 0.134004
R52533 OUT.n12 OUT.t108 0.03175
R52534 OUT.n9 OUT.n7 0.00168421
R52535 OUT.n143 OUT.n4 0.00168421
R52536 OUT.n73 OUT.n71 0.00168421
R52537 OUT.n67 OUT.n66 0.00168421
R52538 OUT.n63 OUT.n62 0.00168421
R52539 OUT.n122 OUT.n120 0.00168421
R52540 OUT.n147 OUT.n1 0.00168421
R52541 a_30324_n30399.t1 a_30324_n30399.t2 24.9025
R52542 a_30324_n30399.t0 a_30324_n30399.t1 19.5272
R52543 a_31284_n30339.t0 a_31284_n30339.t1 26.4056
R52544 a_31284_n30339.t1 a_31284_n30339.t2 18.4133
R52545 a_100992_n29313.t0 a_100992_n29313.t2 23.2303
R52546 a_100992_n29313.t0 a_100992_n29313.t1 21.6695
R52547 a_38097_n5342.t0 a_38097_n5342.t2 123.341
R52548 a_38097_n5342.t2 a_38097_n5342.t1 18.4133
R52549 a_100992_4421.t2 a_100992_4421.t0 21.6693
R52550 a_100992_4421.t1 a_100992_4421.t0 15.3476
R52551 a_71496_10388.n5 a_71496_10388.n1 10.2377
R52552 a_71496_10388.n4 a_71496_10388.t2 10.2108
R52553 a_71496_10388.n4 a_71496_10388.t0 9.99909
R52554 a_71496_10388.n5 a_71496_10388.t5 9.80443
R52555 a_71496_10388.n5 a_71496_10388.t7 9.55135
R52556 a_71496_10388.n0 a_71496_10388.t19 8.17385
R52557 a_71496_10388.n3 a_71496_10388.t12 8.17299
R52558 a_71496_10388.n3 a_71496_10388.t14 8.17134
R52559 a_71496_10388.n0 a_71496_10388.t10 8.16754
R52560 a_71496_10388.n1 a_71496_10388.t11 8.10567
R52561 a_71496_10388.n1 a_71496_10388.t9 8.10567
R52562 a_71496_10388.n3 a_71496_10388.t22 8.10567
R52563 a_71496_10388.n3 a_71496_10388.t23 8.10567
R52564 a_71496_10388.n1 a_71496_10388.t8 8.10567
R52565 a_71496_10388.n1 a_71496_10388.t17 8.10567
R52566 a_71496_10388.n0 a_71496_10388.t13 8.10567
R52567 a_71496_10388.n0 a_71496_10388.t21 8.10567
R52568 a_71496_10388.n6 a_71496_10388.t3 7.74799
R52569 a_71496_10388.n7 a_71496_10388.t6 7.73052
R52570 a_71496_10388.n6 a_71496_10388.t1 7.46478
R52571 a_71496_10388.t4 a_71496_10388.n7 7.1311
R52572 a_71496_10388.n4 a_71496_10388.n6 2.2505
R52573 a_71496_10388.n7 a_71496_10388.n5 2.2505
R52574 a_71496_10388.n1 a_71496_10388.t15 8.35731
R52575 a_71496_10388.n0 a_71496_10388.t20 8.38107
R52576 a_71496_10388.n1 a_71496_10388.t16 8.37583
R52577 a_71496_10388.n1 a_71496_10388.n0 4.35656
R52578 a_71496_10388.n5 a_71496_10388.n4 2.96863
R52579 a_71496_10388.n2 a_71496_10388.n1 1.0882
R52580 a_71496_10388.n2 a_71496_10388.n3 1.08408
R52581 a_71496_10388.n2 a_71496_10388.t18 8.66753
R52582 a_71342_4481.n0 a_71342_4481.t1 10.6581
R52583 a_71342_4481.t2 a_71342_4481.n0 10.2346
R52584 a_71342_4481.n0 a_71342_4481.t3 9.5029
R52585 a_71342_4481.n0 a_71342_4481.t0 9.34796
R52586 a_30152_10448.t3 a_30152_10448.t11 12.7127
R52587 a_30152_10448.t3 a_30152_10448.t6 10.2828
R52588 a_30152_10448.t3 a_30152_10448.t8 10.2828
R52589 a_30152_10448.t3 a_30152_10448.t19 10.2828
R52590 a_30152_10448.t3 a_30152_10448.t14 10.2828
R52591 a_30152_10448.t3 a_30152_10448.t22 10.1333
R52592 a_30152_10448.t3 a_30152_10448.t23 10.1333
R52593 a_30152_10448.t3 a_30152_10448.t10 10.1333
R52594 a_30152_10448.t3 a_30152_10448.t4 10.1333
R52595 a_30152_10448.t3 a_30152_10448.t1 9.72545
R52596 a_30152_10448.t3 a_30152_10448.t21 9.57156
R52597 a_30152_10448.t3 a_30152_10448.t17 9.57156
R52598 a_30152_10448.t3 a_30152_10448.t18 9.57156
R52599 a_30152_10448.t3 a_30152_10448.t13 9.57156
R52600 a_30152_10448.t3 a_30152_10448.t20 9.57156
R52601 a_30152_10448.t3 a_30152_10448.t15 9.57156
R52602 a_30152_10448.t3 a_30152_10448.t16 9.57156
R52603 a_30152_10448.t3 a_30152_10448.t12 9.57156
R52604 a_30152_10448.t1 a_30152_10448.t0 8.02945
R52605 a_30152_10448.t3 a_30152_10448.t2 8.02708
R52606 a_30152_10448.t3 a_30152_10448.t9 7.90829
R52607 a_30152_10448.t3 a_30152_10448.t7 7.90829
R52608 a_30152_10448.t5 a_30152_10448.t3 7.41776
R52609 a_32913_n8930.t0 a_32913_n8930.t1 103.29
R52610 a_32913_n8930.t1 a_32913_n8930.t2 24.9025
R52611 a_31831_n5342.t0 a_31831_n5342.t2 108.376
R52612 a_31831_n5342.t2 a_31831_n5342.t1 18.4133
R52613 a_51711_n5344.t0 a_51711_n5344.t1 13.2434
R52614 a_33379_34917.n1 a_33379_34917.t2 10.937
R52615 a_33379_34917.n1 a_33379_34917.n0 10.9194
R52616 a_33379_34917.n1 a_33379_34917.t1 9.33982
R52617 a_33379_34917.n6 a_33379_34917.n5 1.21431
R52618 a_33379_34917.n9 a_33379_34917.n1 8.36604
R52619 a_33379_34917.n0 a_33379_34917.t82 8.10567
R52620 a_33379_34917.n3 a_33379_34917.t36 8.10567
R52621 a_33379_34917.n3 a_33379_34917.t22 8.10567
R52622 a_33379_34917.n3 a_33379_34917.t78 8.10567
R52623 a_33379_34917.n3 a_33379_34917.t21 8.10567
R52624 a_33379_34917.n0 a_33379_34917.t55 8.10567
R52625 a_33379_34917.n0 a_33379_34917.t27 8.10567
R52626 a_33379_34917.n0 a_33379_34917.t85 8.10567
R52627 a_33379_34917.n0 a_33379_34917.t61 8.10567
R52628 a_33379_34917.n2 a_33379_34917.t44 8.10567
R52629 a_33379_34917.n2 a_33379_34917.t18 8.10567
R52630 a_33379_34917.n2 a_33379_34917.t89 8.10567
R52631 a_33379_34917.n2 a_33379_34917.t49 8.10567
R52632 a_33379_34917.n3 a_33379_34917.t47 8.10567
R52633 a_33379_34917.n3 a_33379_34917.t12 8.10567
R52634 a_33379_34917.n3 a_33379_34917.t71 8.10567
R52635 a_33379_34917.n2 a_33379_34917.t67 8.10567
R52636 a_33379_34917.n2 a_33379_34917.t20 8.10567
R52637 a_33379_34917.n2 a_33379_34917.t77 8.10567
R52638 a_33379_34917.n0 a_33379_34917.t57 8.10567
R52639 a_33379_34917.n0 a_33379_34917.t28 8.10567
R52640 a_33379_34917.n0 a_33379_34917.t6 8.10567
R52641 a_33379_34917.n4 a_33379_34917.t76 8.10567
R52642 a_33379_34917.n0 a_33379_34917.t34 8.10567
R52643 a_33379_34917.n0 a_33379_34917.t16 8.10567
R52644 a_33379_34917.n0 a_33379_34917.t74 8.10567
R52645 a_33379_34917.n0 a_33379_34917.t15 8.10567
R52646 a_33379_34917.n0 a_33379_34917.t50 8.10567
R52647 a_33379_34917.n0 a_33379_34917.t25 8.10567
R52648 a_33379_34917.n0 a_33379_34917.t80 8.10567
R52649 a_33379_34917.n0 a_33379_34917.t54 8.10567
R52650 a_33379_34917.n6 a_33379_34917.t40 8.10567
R52651 a_33379_34917.n6 a_33379_34917.t13 8.10567
R52652 a_33379_34917.n6 a_33379_34917.t84 8.10567
R52653 a_33379_34917.n6 a_33379_34917.t43 8.10567
R52654 a_33379_34917.n0 a_33379_34917.t31 8.10567
R52655 a_33379_34917.n0 a_33379_34917.t81 8.10567
R52656 a_33379_34917.n0 a_33379_34917.t53 8.10567
R52657 a_33379_34917.n4 a_33379_34917.t48 8.10567
R52658 a_33379_34917.n4 a_33379_34917.t91 8.10567
R52659 a_33379_34917.n4 a_33379_34917.t63 8.10567
R52660 a_33379_34917.n4 a_33379_34917.t52 8.10567
R52661 a_33379_34917.n4 a_33379_34917.t26 8.10567
R52662 a_33379_34917.n4 a_33379_34917.t4 8.10567
R52663 a_33379_34917.n0 a_33379_34917.t72 8.10567
R52664 a_33379_34917.n7 a_33379_34917.t32 8.10567
R52665 a_33379_34917.n7 a_33379_34917.t11 8.10567
R52666 a_33379_34917.n7 a_33379_34917.t70 8.10567
R52667 a_33379_34917.n7 a_33379_34917.t10 8.10567
R52668 a_33379_34917.n0 a_33379_34917.t41 8.10567
R52669 a_33379_34917.n0 a_33379_34917.t14 8.10567
R52670 a_33379_34917.n0 a_33379_34917.t73 8.10567
R52671 a_33379_34917.n0 a_33379_34917.t45 8.10567
R52672 a_33379_34917.n0 a_33379_34917.t35 8.10567
R52673 a_33379_34917.n0 a_33379_34917.t8 8.10567
R52674 a_33379_34917.n0 a_33379_34917.t75 8.10567
R52675 a_33379_34917.n0 a_33379_34917.t39 8.10567
R52676 a_33379_34917.n0 a_33379_34917.t37 8.10567
R52677 a_33379_34917.n0 a_33379_34917.t3 8.10567
R52678 a_33379_34917.n0 a_33379_34917.t65 8.10567
R52679 a_33379_34917.n0 a_33379_34917.t64 8.10567
R52680 a_33379_34917.n0 a_33379_34917.t9 8.10567
R52681 a_33379_34917.n0 a_33379_34917.t69 8.10567
R52682 a_33379_34917.n0 a_33379_34917.t42 8.10567
R52683 a_33379_34917.n0 a_33379_34917.t17 8.10567
R52684 a_33379_34917.n0 a_33379_34917.t88 8.10567
R52685 a_33379_34917.n0 a_33379_34917.t83 8.10567
R52686 a_33379_34917.n8 a_33379_34917.t38 8.10567
R52687 a_33379_34917.n8 a_33379_34917.t24 8.10567
R52688 a_33379_34917.n8 a_33379_34917.t79 8.10567
R52689 a_33379_34917.n8 a_33379_34917.t23 8.10567
R52690 a_33379_34917.n0 a_33379_34917.t58 8.10567
R52691 a_33379_34917.n0 a_33379_34917.t29 8.10567
R52692 a_33379_34917.n0 a_33379_34917.t86 8.10567
R52693 a_33379_34917.n0 a_33379_34917.t62 8.10567
R52694 a_33379_34917.n0 a_33379_34917.t46 8.10567
R52695 a_33379_34917.n0 a_33379_34917.t19 8.10567
R52696 a_33379_34917.n0 a_33379_34917.t90 8.10567
R52697 a_33379_34917.n0 a_33379_34917.t51 8.10567
R52698 a_33379_34917.n0 a_33379_34917.t33 8.10567
R52699 a_33379_34917.n0 a_33379_34917.t87 8.10567
R52700 a_33379_34917.n0 a_33379_34917.t60 8.10567
R52701 a_33379_34917.n0 a_33379_34917.t56 8.10567
R52702 a_33379_34917.n0 a_33379_34917.t5 8.10567
R52703 a_33379_34917.n0 a_33379_34917.t66 8.10567
R52704 a_33379_34917.n0 a_33379_34917.t59 8.10567
R52705 a_33379_34917.n0 a_33379_34917.t30 8.10567
R52706 a_33379_34917.n0 a_33379_34917.t7 8.10567
R52707 a_33379_34917.t0 a_33379_34917.n9 6.76216
R52708 a_33379_34917.n9 a_33379_34917.t68 6.15224
R52709 a_33379_34917.n0 a_33379_34917.n2 6.81859
R52710 a_33379_34917.n3 a_33379_34917.n0 6.66138
R52711 a_33379_34917.n5 a_33379_34917.n4 0.358927
R52712 a_33379_34917.n0 a_33379_34917.n5 1.88254
R52713 a_33379_34917.n0 a_33379_34917.n8 5.10926
R52714 a_33379_34917.n7 a_33379_34917.n0 5.07392
R52715 a_45445_n19595.t0 a_45445_n19595.t1 49.4223
R52716 a_45445_n19595.t1 a_45445_n19595.t2 24.9025
R52717 a_71281_n10073.n21 a_71281_n10073.t173 10.5154
R52718 a_71281_n10073.t173 a_71281_n10073.n16 10.5154
R52719 a_71281_n10073.n35 a_71281_n10073.t168 10.5154
R52720 a_71281_n10073.t168 a_71281_n10073.n30 10.5154
R52721 a_71281_n10073.n49 a_71281_n10073.t239 10.5154
R52722 a_71281_n10073.t239 a_71281_n10073.n44 10.5154
R52723 a_71281_n10073.t225 a_71281_n10073.n861 10.5154
R52724 a_71281_n10073.n865 a_71281_n10073.t225 10.5154
R52725 a_71281_n10073.t310 a_71281_n10073.n847 10.5154
R52726 a_71281_n10073.n851 a_71281_n10073.t310 10.5154
R52727 a_71281_n10073.t279 a_71281_n10073.n830 10.5154
R52728 a_71281_n10073.n834 a_71281_n10073.t279 10.5154
R52729 a_71281_n10073.t85 a_71281_n10073.n816 10.5154
R52730 a_71281_n10073.n820 a_71281_n10073.t85 10.5154
R52731 a_71281_n10073.t81 a_71281_n10073.n802 10.5154
R52732 a_71281_n10073.n806 a_71281_n10073.t81 10.5154
R52733 a_71281_n10073.t146 a_71281_n10073.n788 10.5154
R52734 a_71281_n10073.n792 a_71281_n10073.t146 10.5154
R52735 a_71281_n10073.t330 a_71281_n10073.n175 10.5154
R52736 a_71281_n10073.n179 a_71281_n10073.t330 10.5154
R52737 a_71281_n10073.t294 a_71281_n10073.n161 10.5154
R52738 a_71281_n10073.n165 a_71281_n10073.t294 10.5154
R52739 a_71281_n10073.t309 a_71281_n10073.n147 10.5154
R52740 a_71281_n10073.n151 a_71281_n10073.t309 10.5154
R52741 a_71281_n10073.t293 a_71281_n10073.n130 10.5154
R52742 a_71281_n10073.n134 a_71281_n10073.t293 10.5154
R52743 a_71281_n10073.t101 a_71281_n10073.n116 10.5154
R52744 a_71281_n10073.n120 a_71281_n10073.t101 10.5154
R52745 a_71281_n10073.t94 a_71281_n10073.n99 10.5154
R52746 a_71281_n10073.n103 a_71281_n10073.t94 10.5154
R52747 a_71281_n10073.t161 a_71281_n10073.n85 10.5154
R52748 a_71281_n10073.n89 a_71281_n10073.t161 10.5154
R52749 a_71281_n10073.t300 a_71281_n10073.n71 10.5154
R52750 a_71281_n10073.n75 a_71281_n10073.t300 10.5154
R52751 a_71281_n10073.t106 a_71281_n10073.n58 10.5154
R52752 a_71281_n10073.n62 a_71281_n10073.t106 10.5154
R52753 a_71281_n10073.t108 a_71281_n10073.n3 10.5154
R52754 a_71281_n10073.n7 a_71281_n10073.t108 10.5154
R52755 a_71281_n10073.n221 a_71281_n10073.t177 10.5154
R52756 a_71281_n10073.t177 a_71281_n10073.n216 10.5154
R52757 a_71281_n10073.n235 a_71281_n10073.t172 10.5154
R52758 a_71281_n10073.t172 a_71281_n10073.n230 10.5154
R52759 a_71281_n10073.n249 a_71281_n10073.t247 10.5154
R52760 a_71281_n10073.t247 a_71281_n10073.n244 10.5154
R52761 a_71281_n10073.n266 a_71281_n10073.t231 10.5154
R52762 a_71281_n10073.t231 a_71281_n10073.n261 10.5154
R52763 a_71281_n10073.n280 a_71281_n10073.t316 10.5154
R52764 a_71281_n10073.t316 a_71281_n10073.n275 10.5154
R52765 a_71281_n10073.n297 a_71281_n10073.t284 10.5154
R52766 a_71281_n10073.t284 a_71281_n10073.n292 10.5154
R52767 a_71281_n10073.n311 a_71281_n10073.t89 10.5154
R52768 a_71281_n10073.t89 a_71281_n10073.n306 10.5154
R52769 a_71281_n10073.n325 a_71281_n10073.t83 10.5154
R52770 a_71281_n10073.t83 a_71281_n10073.n320 10.5154
R52771 a_71281_n10073.n339 a_71281_n10073.t149 10.5154
R52772 a_71281_n10073.t149 a_71281_n10073.n334 10.5154
R52773 a_71281_n10073.t243 a_71281_n10073.n465 10.5154
R52774 a_71281_n10073.n469 a_71281_n10073.t243 10.5154
R52775 a_71281_n10073.t207 a_71281_n10073.n451 10.5154
R52776 a_71281_n10073.n455 a_71281_n10073.t207 10.5154
R52777 a_71281_n10073.t219 a_71281_n10073.n437 10.5154
R52778 a_71281_n10073.n441 a_71281_n10073.t219 10.5154
R52779 a_71281_n10073.t206 a_71281_n10073.n420 10.5154
R52780 a_71281_n10073.n424 a_71281_n10073.t206 10.5154
R52781 a_71281_n10073.t286 a_71281_n10073.n406 10.5154
R52782 a_71281_n10073.n410 a_71281_n10073.t286 10.5154
R52783 a_71281_n10073.t280 a_71281_n10073.n389 10.5154
R52784 a_71281_n10073.n393 a_71281_n10073.t280 10.5154
R52785 a_71281_n10073.t87 a_71281_n10073.n375 10.5154
R52786 a_71281_n10073.n379 a_71281_n10073.t87 10.5154
R52787 a_71281_n10073.t212 a_71281_n10073.n361 10.5154
R52788 a_71281_n10073.n365 a_71281_n10073.t212 10.5154
R52789 a_71281_n10073.t291 a_71281_n10073.n348 10.5154
R52790 a_71281_n10073.n352 a_71281_n10073.t291 10.5154
R52791 a_71281_n10073.t112 a_71281_n10073.n203 10.5154
R52792 a_71281_n10073.n207 a_71281_n10073.t112 10.5154
R52793 a_71281_n10073.n484 a_71281_n10073.t170 10.5154
R52794 a_71281_n10073.t170 a_71281_n10073.n479 10.5154
R52795 a_71281_n10073.n512 a_71281_n10073.t109 10.5154
R52796 a_71281_n10073.t109 a_71281_n10073.n507 10.5154
R52797 a_71281_n10073.n526 a_71281_n10073.t100 10.5154
R52798 a_71281_n10073.t100 a_71281_n10073.n521 10.5154
R52799 a_71281_n10073.n540 a_71281_n10073.t169 10.5154
R52800 a_71281_n10073.t169 a_71281_n10073.n535 10.5154
R52801 a_71281_n10073.n557 a_71281_n10073.t154 10.5154
R52802 a_71281_n10073.t154 a_71281_n10073.n552 10.5154
R52803 a_71281_n10073.n571 a_71281_n10073.t227 10.5154
R52804 a_71281_n10073.t227 a_71281_n10073.n566 10.5154
R52805 a_71281_n10073.n588 a_71281_n10073.t198 10.5154
R52806 a_71281_n10073.t198 a_71281_n10073.n583 10.5154
R52807 a_71281_n10073.n602 a_71281_n10073.t281 10.5154
R52808 a_71281_n10073.t281 a_71281_n10073.n597 10.5154
R52809 a_71281_n10073.n616 a_71281_n10073.t272 10.5154
R52810 a_71281_n10073.t272 a_71281_n10073.n611 10.5154
R52811 a_71281_n10073.n630 a_71281_n10073.t82 10.5154
R52812 a_71281_n10073.t82 a_71281_n10073.n625 10.5154
R52813 a_71281_n10073.t263 a_71281_n10073.n756 10.5154
R52814 a_71281_n10073.n760 a_71281_n10073.t263 10.5154
R52815 a_71281_n10073.t232 a_71281_n10073.n742 10.5154
R52816 a_71281_n10073.n746 a_71281_n10073.t232 10.5154
R52817 a_71281_n10073.t246 a_71281_n10073.n728 10.5154
R52818 a_71281_n10073.n732 a_71281_n10073.t246 10.5154
R52819 a_71281_n10073.t230 a_71281_n10073.n711 10.5154
R52820 a_71281_n10073.n715 a_71281_n10073.t230 10.5154
R52821 a_71281_n10073.t315 a_71281_n10073.n697 10.5154
R52822 a_71281_n10073.n701 a_71281_n10073.t315 10.5154
R52823 a_71281_n10073.t302 a_71281_n10073.n680 10.5154
R52824 a_71281_n10073.n684 a_71281_n10073.t302 10.5154
R52825 a_71281_n10073.t107 a_71281_n10073.n666 10.5154
R52826 a_71281_n10073.n670 a_71281_n10073.t107 10.5154
R52827 a_71281_n10073.t237 a_71281_n10073.n652 10.5154
R52828 a_71281_n10073.n656 a_71281_n10073.t237 10.5154
R52829 a_71281_n10073.t319 a_71281_n10073.n639 10.5154
R52830 a_71281_n10073.n643 a_71281_n10073.t319 10.5154
R52831 a_71281_n10073.t304 a_71281_n10073.n494 10.5154
R52832 a_71281_n10073.n498 a_71281_n10073.t304 10.5154
R52833 a_71281_n10073.n775 a_71281_n10073.t184 10.5154
R52834 a_71281_n10073.t184 a_71281_n10073.n770 10.5154
R52835 a_71281_n10073.n194 a_71281_n10073.t251 10.5154
R52836 a_71281_n10073.t251 a_71281_n10073.n189 10.5154
R52837 a_71281_n10073.n789 a_71281_n10073.t214 10.515
R52838 a_71281_n10073.n59 a_71281_n10073.t126 10.515
R52839 a_71281_n10073.n336 a_71281_n10073.t218 10.515
R52840 a_71281_n10073.n349 a_71281_n10073.t325 10.515
R52841 a_71281_n10073.n627 a_71281_n10073.t181 10.515
R52842 a_71281_n10073.n640 a_71281_n10073.t202 10.515
R52843 a_71281_n10073.n17 a_71281_n10073.t254 10.515
R52844 a_71281_n10073.n18 a_71281_n10073.t254 10.515
R52845 a_71281_n10073.n31 a_71281_n10073.t241 10.515
R52846 a_71281_n10073.n32 a_71281_n10073.t241 10.515
R52847 a_71281_n10073.n45 a_71281_n10073.t321 10.515
R52848 a_71281_n10073.n46 a_71281_n10073.t321 10.515
R52849 a_71281_n10073.n863 a_71281_n10073.t312 10.515
R52850 a_71281_n10073.n862 a_71281_n10073.t312 10.515
R52851 a_71281_n10073.n849 a_71281_n10073.t114 10.515
R52852 a_71281_n10073.n848 a_71281_n10073.t114 10.515
R52853 a_71281_n10073.n832 a_71281_n10073.t86 10.515
R52854 a_71281_n10073.n831 a_71281_n10073.t86 10.515
R52855 a_71281_n10073.n818 a_71281_n10073.t152 10.515
R52856 a_71281_n10073.n817 a_71281_n10073.t152 10.515
R52857 a_71281_n10073.n804 a_71281_n10073.t148 10.515
R52858 a_71281_n10073.n803 a_71281_n10073.t148 10.515
R52859 a_71281_n10073.n790 a_71281_n10073.t214 10.515
R52860 a_71281_n10073.n177 a_71281_n10073.t76 10.515
R52861 a_71281_n10073.n176 a_71281_n10073.t76 10.515
R52862 a_71281_n10073.n163 a_71281_n10073.t329 10.515
R52863 a_71281_n10073.n162 a_71281_n10073.t329 10.515
R52864 a_71281_n10073.n149 a_71281_n10073.t336 10.515
R52865 a_71281_n10073.n148 a_71281_n10073.t336 10.515
R52866 a_71281_n10073.n132 a_71281_n10073.t328 10.515
R52867 a_71281_n10073.n131 a_71281_n10073.t328 10.515
R52868 a_71281_n10073.n118 a_71281_n10073.t124 10.515
R52869 a_71281_n10073.n117 a_71281_n10073.t124 10.515
R52870 a_71281_n10073.n101 a_71281_n10073.t119 10.515
R52871 a_71281_n10073.n100 a_71281_n10073.t119 10.515
R52872 a_71281_n10073.n87 a_71281_n10073.t183 10.515
R52873 a_71281_n10073.n86 a_71281_n10073.t183 10.515
R52874 a_71281_n10073.n73 a_71281_n10073.t333 10.515
R52875 a_71281_n10073.n72 a_71281_n10073.t333 10.515
R52876 a_71281_n10073.n60 a_71281_n10073.t126 10.515
R52877 a_71281_n10073.n5 a_71281_n10073.t174 10.515
R52878 a_71281_n10073.n4 a_71281_n10073.t174 10.515
R52879 a_71281_n10073.n217 a_71281_n10073.t259 10.515
R52880 a_71281_n10073.n218 a_71281_n10073.t259 10.515
R52881 a_71281_n10073.n231 a_71281_n10073.t250 10.515
R52882 a_71281_n10073.n232 a_71281_n10073.t250 10.515
R52883 a_71281_n10073.n245 a_71281_n10073.t327 10.515
R52884 a_71281_n10073.n246 a_71281_n10073.t327 10.515
R52885 a_71281_n10073.n262 a_71281_n10073.t317 10.515
R52886 a_71281_n10073.n263 a_71281_n10073.t317 10.515
R52887 a_71281_n10073.n276 a_71281_n10073.t118 10.515
R52888 a_71281_n10073.n277 a_71281_n10073.t118 10.515
R52889 a_71281_n10073.n293 a_71281_n10073.t93 10.515
R52890 a_71281_n10073.n294 a_71281_n10073.t93 10.515
R52891 a_71281_n10073.n307 a_71281_n10073.t159 10.515
R52892 a_71281_n10073.n308 a_71281_n10073.t159 10.515
R52893 a_71281_n10073.n321 a_71281_n10073.t150 10.515
R52894 a_71281_n10073.n322 a_71281_n10073.t150 10.515
R52895 a_71281_n10073.n335 a_71281_n10073.t218 10.515
R52896 a_71281_n10073.n467 a_71281_n10073.t264 10.515
R52897 a_71281_n10073.n466 a_71281_n10073.t264 10.515
R52898 a_71281_n10073.n453 a_71281_n10073.t242 10.515
R52899 a_71281_n10073.n452 a_71281_n10073.t242 10.515
R52900 a_71281_n10073.n439 a_71281_n10073.t253 10.515
R52901 a_71281_n10073.n438 a_71281_n10073.t253 10.515
R52902 a_71281_n10073.n422 a_71281_n10073.t240 10.515
R52903 a_71281_n10073.n421 a_71281_n10073.t240 10.515
R52904 a_71281_n10073.n408 a_71281_n10073.t320 10.515
R52905 a_71281_n10073.n407 a_71281_n10073.t320 10.515
R52906 a_71281_n10073.n391 a_71281_n10073.t311 10.515
R52907 a_71281_n10073.n390 a_71281_n10073.t311 10.515
R52908 a_71281_n10073.n377 a_71281_n10073.t113 10.515
R52909 a_71281_n10073.n376 a_71281_n10073.t113 10.515
R52910 a_71281_n10073.n363 a_71281_n10073.t249 10.515
R52911 a_71281_n10073.n362 a_71281_n10073.t249 10.515
R52912 a_71281_n10073.n350 a_71281_n10073.t325 10.515
R52913 a_71281_n10073.n205 a_71281_n10073.t178 10.515
R52914 a_71281_n10073.n204 a_71281_n10073.t178 10.515
R52915 a_71281_n10073.n480 a_71281_n10073.t186 10.515
R52916 a_71281_n10073.n481 a_71281_n10073.t186 10.515
R52917 a_71281_n10073.n508 a_71281_n10073.t195 10.515
R52918 a_71281_n10073.n509 a_71281_n10073.t195 10.515
R52919 a_71281_n10073.n522 a_71281_n10073.t189 10.515
R52920 a_71281_n10073.n523 a_71281_n10073.t189 10.515
R52921 a_71281_n10073.n536 a_71281_n10073.t270 10.515
R52922 a_71281_n10073.n537 a_71281_n10073.t270 10.515
R52923 a_71281_n10073.n553 a_71281_n10073.t267 10.515
R52924 a_71281_n10073.n554 a_71281_n10073.t267 10.515
R52925 a_71281_n10073.n567 a_71281_n10073.t74 10.515
R52926 a_71281_n10073.n568 a_71281_n10073.t74 10.515
R52927 a_71281_n10073.n584 a_71281_n10073.t323 10.515
R52928 a_71281_n10073.n585 a_71281_n10073.t323 10.515
R52929 a_71281_n10073.n598 a_71281_n10073.t122 10.515
R52930 a_71281_n10073.n599 a_71281_n10073.t122 10.515
R52931 a_71281_n10073.n612 a_71281_n10073.t117 10.515
R52932 a_71281_n10073.n613 a_71281_n10073.t117 10.515
R52933 a_71281_n10073.n626 a_71281_n10073.t181 10.515
R52934 a_71281_n10073.n758 a_71281_n10073.t157 10.515
R52935 a_71281_n10073.n757 a_71281_n10073.t157 10.515
R52936 a_71281_n10073.n744 a_71281_n10073.t135 10.515
R52937 a_71281_n10073.n743 a_71281_n10073.t135 10.515
R52938 a_71281_n10073.n730 a_71281_n10073.t145 10.515
R52939 a_71281_n10073.n729 a_71281_n10073.t145 10.515
R52940 a_71281_n10073.n713 a_71281_n10073.t132 10.515
R52941 a_71281_n10073.n712 a_71281_n10073.t132 10.515
R52942 a_71281_n10073.n699 a_71281_n10073.t200 10.515
R52943 a_71281_n10073.n698 a_71281_n10073.t200 10.515
R52944 a_71281_n10073.n682 a_71281_n10073.t192 10.515
R52945 a_71281_n10073.n681 a_71281_n10073.t192 10.515
R52946 a_71281_n10073.n668 a_71281_n10073.t274 10.515
R52947 a_71281_n10073.n667 a_71281_n10073.t274 10.515
R52948 a_71281_n10073.n654 a_71281_n10073.t138 10.515
R52949 a_71281_n10073.n653 a_71281_n10073.t138 10.515
R52950 a_71281_n10073.n641 a_71281_n10073.t202 10.515
R52951 a_71281_n10073.n496 a_71281_n10073.t130 10.515
R52952 a_71281_n10073.n495 a_71281_n10073.t130 10.515
R52953 a_71281_n10073.n771 a_71281_n10073.t92 10.515
R52954 a_71281_n10073.n772 a_71281_n10073.t92 10.515
R52955 a_71281_n10073.n190 a_71281_n10073.t268 10.515
R52956 a_71281_n10073.n191 a_71281_n10073.t268 10.515
R52957 a_71281_n10073.n21 a_71281_n10073.t121 9.57886
R52958 a_71281_n10073.t121 a_71281_n10073.n16 9.57886
R52959 a_71281_n10073.n18 a_71281_n10073.t313 9.57886
R52960 a_71281_n10073.t313 a_71281_n10073.n17 9.57886
R52961 a_71281_n10073.n35 a_71281_n10073.t116 9.57886
R52962 a_71281_n10073.t116 a_71281_n10073.n30 9.57886
R52963 a_71281_n10073.n32 a_71281_n10073.t299 9.57886
R52964 a_71281_n10073.t299 a_71281_n10073.n31 9.57886
R52965 a_71281_n10073.n49 a_71281_n10073.t180 9.57886
R52966 a_71281_n10073.t180 a_71281_n10073.n44 9.57886
R52967 a_71281_n10073.n46 a_71281_n10073.t105 9.57886
R52968 a_71281_n10073.t105 a_71281_n10073.n45 9.57886
R52969 a_71281_n10073.t42 a_71281_n10073.n861 9.57886
R52970 a_71281_n10073.n865 a_71281_n10073.t42 9.57886
R52971 a_71281_n10073.t70 a_71281_n10073.n862 9.57886
R52972 a_71281_n10073.n863 a_71281_n10073.t70 9.57886
R52973 a_71281_n10073.t14 a_71281_n10073.n847 9.57886
R52974 a_71281_n10073.n851 a_71281_n10073.t14 9.57886
R52975 a_71281_n10073.t46 a_71281_n10073.n848 9.57886
R52976 a_71281_n10073.n849 a_71281_n10073.t46 9.57886
R52977 a_71281_n10073.t215 a_71281_n10073.n830 9.57886
R52978 a_71281_n10073.n834 a_71281_n10073.t215 9.57886
R52979 a_71281_n10073.t139 a_71281_n10073.n831 9.57886
R52980 a_71281_n10073.n832 a_71281_n10073.t139 9.57886
R52981 a_71281_n10073.t297 a_71281_n10073.n816 9.57886
R52982 a_71281_n10073.n820 a_71281_n10073.t297 9.57886
R52983 a_71281_n10073.t203 a_71281_n10073.n817 9.57886
R52984 a_71281_n10073.n818 a_71281_n10073.t203 9.57886
R52985 a_71281_n10073.t285 a_71281_n10073.n802 9.57886
R52986 a_71281_n10073.n806 a_71281_n10073.t285 9.57886
R52987 a_71281_n10073.t196 a_71281_n10073.n803 9.57886
R52988 a_71281_n10073.n804 a_71281_n10073.t196 9.57886
R52989 a_71281_n10073.t98 a_71281_n10073.n788 9.57886
R52990 a_71281_n10073.n792 a_71281_n10073.t98 9.57886
R52991 a_71281_n10073.t277 a_71281_n10073.n789 9.57886
R52992 a_71281_n10073.n790 a_71281_n10073.t277 9.57886
R52993 a_71281_n10073.t142 a_71281_n10073.n175 9.57886
R52994 a_71281_n10073.n179 a_71281_n10073.t142 9.57886
R52995 a_71281_n10073.t238 a_71281_n10073.n176 9.57886
R52996 a_71281_n10073.n177 a_71281_n10073.t238 9.57886
R52997 a_71281_n10073.t127 a_71281_n10073.n161 9.57886
R52998 a_71281_n10073.n165 a_71281_n10073.t127 9.57886
R52999 a_71281_n10073.t204 a_71281_n10073.n162 9.57886
R53000 a_71281_n10073.n163 a_71281_n10073.t204 9.57886
R53001 a_71281_n10073.t129 a_71281_n10073.n147 9.57886
R53002 a_71281_n10073.n151 a_71281_n10073.t129 9.57886
R53003 a_71281_n10073.t216 a_71281_n10073.n148 9.57886
R53004 a_71281_n10073.n149 a_71281_n10073.t216 9.57886
R53005 a_71281_n10073.t58 a_71281_n10073.n130 9.57886
R53006 a_71281_n10073.n134 a_71281_n10073.t58 9.57886
R53007 a_71281_n10073.t28 a_71281_n10073.n131 9.57886
R53008 a_71281_n10073.n132 a_71281_n10073.t28 9.57886
R53009 a_71281_n10073.t36 a_71281_n10073.n116 9.57886
R53010 a_71281_n10073.n120 a_71281_n10073.t36 9.57886
R53011 a_71281_n10073.t12 a_71281_n10073.n117 9.57886
R53012 a_71281_n10073.n118 a_71281_n10073.t12 9.57886
R53013 a_71281_n10073.t187 a_71281_n10073.n99 9.57886
R53014 a_71281_n10073.n103 a_71281_n10073.t187 9.57886
R53015 a_71281_n10073.t278 a_71281_n10073.n100 9.57886
R53016 a_71281_n10073.n101 a_71281_n10073.t278 9.57886
R53017 a_71281_n10073.t265 a_71281_n10073.n85 9.57886
R53018 a_71281_n10073.n89 a_71281_n10073.t265 9.57886
R53019 a_71281_n10073.t84 a_71281_n10073.n86 9.57886
R53020 a_71281_n10073.n87 a_71281_n10073.t84 9.57886
R53021 a_71281_n10073.t128 a_71281_n10073.n71 9.57886
R53022 a_71281_n10073.n75 a_71281_n10073.t128 9.57886
R53023 a_71281_n10073.t210 a_71281_n10073.n72 9.57886
R53024 a_71281_n10073.n73 a_71281_n10073.t210 9.57886
R53025 a_71281_n10073.t190 a_71281_n10073.n58 9.57886
R53026 a_71281_n10073.n62 a_71281_n10073.t190 9.57886
R53027 a_71281_n10073.t288 a_71281_n10073.n59 9.57886
R53028 a_71281_n10073.n60 a_71281_n10073.t288 9.57886
R53029 a_71281_n10073.t322 a_71281_n10073.n3 9.57886
R53030 a_71281_n10073.n7 a_71281_n10073.t322 9.57886
R53031 a_71281_n10073.t228 a_71281_n10073.n4 9.57886
R53032 a_71281_n10073.n5 a_71281_n10073.t228 9.57886
R53033 a_71281_n10073.n221 a_71281_n10073.t185 9.57886
R53034 a_71281_n10073.t185 a_71281_n10073.n216 9.57886
R53035 a_71281_n10073.n218 a_71281_n10073.t318 9.57886
R53036 a_71281_n10073.t318 a_71281_n10073.n217 9.57886
R53037 a_71281_n10073.n235 a_71281_n10073.t179 9.57886
R53038 a_71281_n10073.t179 a_71281_n10073.n230 9.57886
R53039 a_71281_n10073.n232 a_71281_n10073.t305 9.57886
R53040 a_71281_n10073.t305 a_71281_n10073.n231 9.57886
R53041 a_71281_n10073.n249 a_71281_n10073.t260 9.57886
R53042 a_71281_n10073.t260 a_71281_n10073.n244 9.57886
R53043 a_71281_n10073.n246 a_71281_n10073.t110 9.57886
R53044 a_71281_n10073.t110 a_71281_n10073.n245 9.57886
R53045 a_71281_n10073.n266 a_71281_n10073.t16 9.57886
R53046 a_71281_n10073.t16 a_71281_n10073.n261 9.57886
R53047 a_71281_n10073.n263 a_71281_n10073.t66 9.57886
R53048 a_71281_n10073.t66 a_71281_n10073.n262 9.57886
R53049 a_71281_n10073.n280 a_71281_n10073.t0 9.57886
R53050 a_71281_n10073.t0 a_71281_n10073.n275 9.57886
R53051 a_71281_n10073.n277 a_71281_n10073.t44 9.57886
R53052 a_71281_n10073.t44 a_71281_n10073.n276 9.57886
R53053 a_71281_n10073.n297 a_71281_n10073.t295 9.57886
R53054 a_71281_n10073.t295 a_71281_n10073.n292 9.57886
R53055 a_71281_n10073.n294 a_71281_n10073.t143 9.57886
R53056 a_71281_n10073.t143 a_71281_n10073.n293 9.57886
R53057 a_71281_n10073.n311 a_71281_n10073.t102 9.57886
R53058 a_71281_n10073.t102 a_71281_n10073.n306 9.57886
R53059 a_71281_n10073.n308 a_71281_n10073.t209 9.57886
R53060 a_71281_n10073.t209 a_71281_n10073.n307 9.57886
R53061 a_71281_n10073.n325 a_71281_n10073.t95 9.57886
R53062 a_71281_n10073.t95 a_71281_n10073.n320 9.57886
R53063 a_71281_n10073.n322 a_71281_n10073.t199 9.57886
R53064 a_71281_n10073.t199 a_71281_n10073.n321 9.57886
R53065 a_71281_n10073.n339 a_71281_n10073.t162 9.57886
R53066 a_71281_n10073.t162 a_71281_n10073.n334 9.57886
R53067 a_71281_n10073.n336 a_71281_n10073.t283 9.57886
R53068 a_71281_n10073.t283 a_71281_n10073.n335 9.57886
R53069 a_71281_n10073.t256 a_71281_n10073.n465 9.57886
R53070 a_71281_n10073.n469 a_71281_n10073.t256 9.57886
R53071 a_71281_n10073.t156 a_71281_n10073.n466 9.57886
R53072 a_71281_n10073.n467 a_71281_n10073.t156 9.57886
R53073 a_71281_n10073.t222 a_71281_n10073.n451 9.57886
R53074 a_71281_n10073.n455 a_71281_n10073.t222 9.57886
R53075 a_71281_n10073.t133 a_71281_n10073.n452 9.57886
R53076 a_71281_n10073.n453 a_71281_n10073.t133 9.57886
R53077 a_71281_n10073.t234 a_71281_n10073.n437 9.57886
R53078 a_71281_n10073.n441 a_71281_n10073.t234 9.57886
R53079 a_71281_n10073.t144 a_71281_n10073.n438 9.57886
R53080 a_71281_n10073.n439 a_71281_n10073.t144 9.57886
R53081 a_71281_n10073.t24 a_71281_n10073.n420 9.57886
R53082 a_71281_n10073.n424 a_71281_n10073.t24 9.57886
R53083 a_71281_n10073.t54 a_71281_n10073.n421 9.57886
R53084 a_71281_n10073.n422 a_71281_n10073.t54 9.57886
R53085 a_71281_n10073.t4 a_71281_n10073.n406 9.57886
R53086 a_71281_n10073.n410 a_71281_n10073.t4 9.57886
R53087 a_71281_n10073.t32 a_71281_n10073.n407 9.57886
R53088 a_71281_n10073.n408 a_71281_n10073.t32 9.57886
R53089 a_71281_n10073.t287 a_71281_n10073.n389 9.57886
R53090 a_71281_n10073.n393 a_71281_n10073.t287 9.57886
R53091 a_71281_n10073.t191 a_71281_n10073.n390 9.57886
R53092 a_71281_n10073.n391 a_71281_n10073.t191 9.57886
R53093 a_71281_n10073.t99 a_71281_n10073.n375 9.57886
R53094 a_71281_n10073.n379 a_71281_n10073.t99 9.57886
R53095 a_71281_n10073.t273 a_71281_n10073.n376 9.57886
R53096 a_71281_n10073.n377 a_71281_n10073.t273 9.57886
R53097 a_71281_n10073.t224 a_71281_n10073.n361 9.57886
R53098 a_71281_n10073.n365 a_71281_n10073.t224 9.57886
R53099 a_71281_n10073.t137 a_71281_n10073.n362 9.57886
R53100 a_71281_n10073.n363 a_71281_n10073.t137 9.57886
R53101 a_71281_n10073.t308 a_71281_n10073.n348 9.57886
R53102 a_71281_n10073.n352 a_71281_n10073.t308 9.57886
R53103 a_71281_n10073.t201 a_71281_n10073.n349 9.57886
R53104 a_71281_n10073.n350 a_71281_n10073.t201 9.57886
R53105 a_71281_n10073.t120 a_71281_n10073.n203 9.57886
R53106 a_71281_n10073.n207 a_71281_n10073.t120 9.57886
R53107 a_71281_n10073.t235 a_71281_n10073.n204 9.57886
R53108 a_71281_n10073.n205 a_71281_n10073.t235 9.57886
R53109 a_71281_n10073.n484 a_71281_n10073.t175 9.57886
R53110 a_71281_n10073.t175 a_71281_n10073.n479 9.57886
R53111 a_71281_n10073.n481 a_71281_n10073.t91 9.57886
R53112 a_71281_n10073.t91 a_71281_n10073.n480 9.57886
R53113 a_71281_n10073.n512 a_71281_n10073.t80 9.57886
R53114 a_71281_n10073.t80 a_71281_n10073.n507 9.57886
R53115 a_71281_n10073.n509 a_71281_n10073.t233 9.57886
R53116 a_71281_n10073.t233 a_71281_n10073.n508 9.57886
R53117 a_71281_n10073.n526 a_71281_n10073.t75 9.57886
R53118 a_71281_n10073.t75 a_71281_n10073.n521 9.57886
R53119 a_71281_n10073.n523 a_71281_n10073.t220 9.57886
R53120 a_71281_n10073.t220 a_71281_n10073.n522 9.57886
R53121 a_71281_n10073.n540 a_71281_n10073.t134 9.57886
R53122 a_71281_n10073.t134 a_71281_n10073.n535 9.57886
R53123 a_71281_n10073.n537 a_71281_n10073.t303 9.57886
R53124 a_71281_n10073.t303 a_71281_n10073.n536 9.57886
R53125 a_71281_n10073.n557 a_71281_n10073.t56 9.57886
R53126 a_71281_n10073.t56 a_71281_n10073.n552 9.57886
R53127 a_71281_n10073.n554 a_71281_n10073.t10 9.57886
R53128 a_71281_n10073.t10 a_71281_n10073.n553 9.57886
R53129 a_71281_n10073.n571 a_71281_n10073.t34 9.57886
R53130 a_71281_n10073.t34 a_71281_n10073.n566 9.57886
R53131 a_71281_n10073.n568 a_71281_n10073.t68 9.57886
R53132 a_71281_n10073.t68 a_71281_n10073.n567 9.57886
R53133 a_71281_n10073.n588 a_71281_n10073.t182 9.57886
R53134 a_71281_n10073.t182 a_71281_n10073.n583 9.57886
R53135 a_71281_n10073.n585 a_71281_n10073.t77 9.57886
R53136 a_71281_n10073.t77 a_71281_n10073.n584 9.57886
R53137 a_71281_n10073.n602 a_71281_n10073.t262 9.57886
R53138 a_71281_n10073.t262 a_71281_n10073.n597 9.57886
R53139 a_71281_n10073.n599 a_71281_n10073.t141 9.57886
R53140 a_71281_n10073.t141 a_71281_n10073.n598 9.57886
R53141 a_71281_n10073.n616 a_71281_n10073.t255 9.57886
R53142 a_71281_n10073.t255 a_71281_n10073.n611 9.57886
R53143 a_71281_n10073.n613 a_71281_n10073.t131 9.57886
R53144 a_71281_n10073.t131 a_71281_n10073.n612 9.57886
R53145 a_71281_n10073.n630 a_71281_n10073.t334 9.57886
R53146 a_71281_n10073.t334 a_71281_n10073.n625 9.57886
R53147 a_71281_n10073.n627 a_71281_n10073.t197 9.57886
R53148 a_71281_n10073.t197 a_71281_n10073.n626 9.57886
R53149 a_71281_n10073.t244 a_71281_n10073.n756 9.57886
R53150 a_71281_n10073.n760 a_71281_n10073.t244 9.57886
R53151 a_71281_n10073.t176 a_71281_n10073.n757 9.57886
R53152 a_71281_n10073.n758 a_71281_n10073.t176 9.57886
R53153 a_71281_n10073.t208 a_71281_n10073.n742 9.57886
R53154 a_71281_n10073.n746 a_71281_n10073.t208 9.57886
R53155 a_71281_n10073.t151 a_71281_n10073.n743 9.57886
R53156 a_71281_n10073.n744 a_71281_n10073.t151 9.57886
R53157 a_71281_n10073.t221 a_71281_n10073.n728 9.57886
R53158 a_71281_n10073.n732 a_71281_n10073.t221 9.57886
R53159 a_71281_n10073.t165 a_71281_n10073.n729 9.57886
R53160 a_71281_n10073.n730 a_71281_n10073.t165 9.57886
R53161 a_71281_n10073.t26 a_71281_n10073.n711 9.57886
R53162 a_71281_n10073.n715 a_71281_n10073.t26 9.57886
R53163 a_71281_n10073.t48 a_71281_n10073.n712 9.57886
R53164 a_71281_n10073.n713 a_71281_n10073.t48 9.57886
R53165 a_71281_n10073.t8 a_71281_n10073.n697 9.57886
R53166 a_71281_n10073.n701 a_71281_n10073.t8 9.57886
R53167 a_71281_n10073.t20 a_71281_n10073.n698 9.57886
R53168 a_71281_n10073.n699 a_71281_n10073.t20 9.57886
R53169 a_71281_n10073.t282 a_71281_n10073.n680 9.57886
R53170 a_71281_n10073.n684 a_71281_n10073.t282 9.57886
R53171 a_71281_n10073.t211 a_71281_n10073.n681 9.57886
R53172 a_71281_n10073.n682 a_71281_n10073.t211 9.57886
R53173 a_71281_n10073.t88 a_71281_n10073.n666 9.57886
R53174 a_71281_n10073.n670 a_71281_n10073.t88 9.57886
R53175 a_71281_n10073.t289 a_71281_n10073.n667 9.57886
R53176 a_71281_n10073.n668 a_71281_n10073.t289 9.57886
R53177 a_71281_n10073.t213 a_71281_n10073.n652 9.57886
R53178 a_71281_n10073.n656 a_71281_n10073.t213 9.57886
R53179 a_71281_n10073.t153 a_71281_n10073.n653 9.57886
R53180 a_71281_n10073.n654 a_71281_n10073.t153 9.57886
R53181 a_71281_n10073.t292 a_71281_n10073.n639 9.57886
R53182 a_71281_n10073.n643 a_71281_n10073.t292 9.57886
R53183 a_71281_n10073.t226 a_71281_n10073.n640 9.57886
R53184 a_71281_n10073.n641 a_71281_n10073.t226 9.57886
R53185 a_71281_n10073.t271 a_71281_n10073.n494 9.57886
R53186 a_71281_n10073.n498 a_71281_n10073.t271 9.57886
R53187 a_71281_n10073.t160 a_71281_n10073.n495 9.57886
R53188 a_71281_n10073.n496 a_71281_n10073.t160 9.57886
R53189 a_71281_n10073.n775 a_71281_n10073.t171 9.57886
R53190 a_71281_n10073.t171 a_71281_n10073.n770 9.57886
R53191 a_71281_n10073.n772 a_71281_n10073.t111 9.57886
R53192 a_71281_n10073.t111 a_71281_n10073.n771 9.57886
R53193 a_71281_n10073.n194 a_71281_n10073.t79 9.57886
R53194 a_71281_n10073.t79 a_71281_n10073.n189 9.57886
R53195 a_71281_n10073.n191 a_71281_n10073.t167 9.57886
R53196 a_71281_n10073.t167 a_71281_n10073.n190 9.57886
R53197 a_71281_n10073.t337 a_71281_n10073.n23 8.10567
R53198 a_71281_n10073.n24 a_71281_n10073.t337 8.10567
R53199 a_71281_n10073.t332 a_71281_n10073.n37 8.10567
R53200 a_71281_n10073.n38 a_71281_n10073.t332 8.10567
R53201 a_71281_n10073.t125 a_71281_n10073.n51 8.10567
R53202 a_71281_n10073.n52 a_71281_n10073.t125 8.10567
R53203 a_71281_n10073.n869 a_71281_n10073.t60 8.10567
R53204 a_71281_n10073.t60 a_71281_n10073.n868 8.10567
R53205 a_71281_n10073.n855 a_71281_n10073.t38 8.10567
R53206 a_71281_n10073.t38 a_71281_n10073.n854 8.10567
R53207 a_71281_n10073.n838 a_71281_n10073.t166 8.10567
R53208 a_71281_n10073.t166 a_71281_n10073.n837 8.10567
R53209 a_71281_n10073.n824 a_71281_n10073.t236 8.10567
R53210 a_71281_n10073.t236 a_71281_n10073.n823 8.10567
R53211 a_71281_n10073.n810 a_71281_n10073.t223 8.10567
R53212 a_71281_n10073.t223 a_71281_n10073.n809 8.10567
R53213 a_71281_n10073.n796 a_71281_n10073.t307 8.10567
R53214 a_71281_n10073.t307 a_71281_n10073.n795 8.10567
R53215 a_71281_n10073.n183 a_71281_n10073.t324 8.10567
R53216 a_71281_n10073.t324 a_71281_n10073.n182 8.10567
R53217 a_71281_n10073.n169 a_71281_n10073.t290 8.10567
R53218 a_71281_n10073.t290 a_71281_n10073.n168 8.10567
R53219 a_71281_n10073.n155 a_71281_n10073.t306 8.10567
R53220 a_71281_n10073.t306 a_71281_n10073.n154 8.10567
R53221 a_71281_n10073.n138 a_71281_n10073.t6 8.10567
R53222 a_71281_n10073.t6 a_71281_n10073.n137 8.10567
R53223 a_71281_n10073.n124 a_71281_n10073.t64 8.10567
R53224 a_71281_n10073.t64 a_71281_n10073.n123 8.10567
R53225 a_71281_n10073.n107 a_71281_n10073.t90 8.10567
R53226 a_71281_n10073.t90 a_71281_n10073.n106 8.10567
R53227 a_71281_n10073.n93 a_71281_n10073.t155 8.10567
R53228 a_71281_n10073.t155 a_71281_n10073.n92 8.10567
R53229 a_71281_n10073.n79 a_71281_n10073.t298 8.10567
R53230 a_71281_n10073.t298 a_71281_n10073.n78 8.10567
R53231 a_71281_n10073.n65 a_71281_n10073.t104 8.10567
R53232 a_71281_n10073.t104 a_71281_n10073.n64 8.10567
R53233 a_71281_n10073.n10 a_71281_n10073.t261 8.10567
R53234 a_71281_n10073.t261 a_71281_n10073.n9 8.10567
R53235 a_71281_n10073.t103 a_71281_n10073.n223 8.10567
R53236 a_71281_n10073.n224 a_71281_n10073.t103 8.10567
R53237 a_71281_n10073.t96 a_71281_n10073.n237 8.10567
R53238 a_71281_n10073.n238 a_71281_n10073.t96 8.10567
R53239 a_71281_n10073.t163 a_71281_n10073.n251 8.10567
R53240 a_71281_n10073.n252 a_71281_n10073.t163 8.10567
R53241 a_71281_n10073.t50 a_71281_n10073.n268 8.10567
R53242 a_71281_n10073.n269 a_71281_n10073.t50 8.10567
R53243 a_71281_n10073.t22 a_71281_n10073.n282 8.10567
R53244 a_71281_n10073.n283 a_71281_n10073.t22 8.10567
R53245 a_71281_n10073.t194 a_71281_n10073.n299 8.10567
R53246 a_71281_n10073.n300 a_71281_n10073.t194 8.10567
R53247 a_71281_n10073.t276 a_71281_n10073.n313 8.10567
R53248 a_71281_n10073.n314 a_71281_n10073.t276 8.10567
R53249 a_71281_n10073.t269 a_71281_n10073.n327 8.10567
R53250 a_71281_n10073.n328 a_71281_n10073.t269 8.10567
R53251 a_71281_n10073.t78 a_71281_n10073.n341 8.10567
R53252 a_71281_n10073.n342 a_71281_n10073.t78 8.10567
R53253 a_71281_n10073.n473 a_71281_n10073.t266 8.10567
R53254 a_71281_n10073.t266 a_71281_n10073.n472 8.10567
R53255 a_71281_n10073.n459 a_71281_n10073.t245 8.10567
R53256 a_71281_n10073.t245 a_71281_n10073.n458 8.10567
R53257 a_71281_n10073.n445 a_71281_n10073.t257 8.10567
R53258 a_71281_n10073.t257 a_71281_n10073.n444 8.10567
R53259 a_71281_n10073.n428 a_71281_n10073.t18 8.10567
R53260 a_71281_n10073.t18 a_71281_n10073.n427 8.10567
R53261 a_71281_n10073.n414 a_71281_n10073.t2 8.10567
R53262 a_71281_n10073.t2 a_71281_n10073.n413 8.10567
R53263 a_71281_n10073.n397 a_71281_n10073.t314 8.10567
R53264 a_71281_n10073.t314 a_71281_n10073.n396 8.10567
R53265 a_71281_n10073.n383 a_71281_n10073.t115 8.10567
R53266 a_71281_n10073.t115 a_71281_n10073.n382 8.10567
R53267 a_71281_n10073.n369 a_71281_n10073.t252 8.10567
R53268 a_71281_n10073.t252 a_71281_n10073.n368 8.10567
R53269 a_71281_n10073.n355 a_71281_n10073.t331 8.10567
R53270 a_71281_n10073.t331 a_71281_n10073.n354 8.10567
R53271 a_71281_n10073.n210 a_71281_n10073.t296 8.10567
R53272 a_71281_n10073.t296 a_71281_n10073.n209 8.10567
R53273 a_71281_n10073.t188 a_71281_n10073.n486 8.10567
R53274 a_71281_n10073.n487 a_71281_n10073.t188 8.10567
R53275 a_71281_n10073.t335 a_71281_n10073.n514 8.10567
R53276 a_71281_n10073.n515 a_71281_n10073.t335 8.10567
R53277 a_71281_n10073.t326 a_71281_n10073.n528 8.10567
R53278 a_71281_n10073.n529 a_71281_n10073.t326 8.10567
R53279 a_71281_n10073.t123 a_71281_n10073.n542 8.10567
R53280 a_71281_n10073.n543 a_71281_n10073.t123 8.10567
R53281 a_71281_n10073.t62 a_71281_n10073.n559 8.10567
R53282 a_71281_n10073.n560 a_71281_n10073.t62 8.10567
R53283 a_71281_n10073.t40 a_71281_n10073.n573 8.10567
R53284 a_71281_n10073.n574 a_71281_n10073.t40 8.10567
R53285 a_71281_n10073.t158 a_71281_n10073.n590 8.10567
R53286 a_71281_n10073.n591 a_71281_n10073.t158 8.10567
R53287 a_71281_n10073.t229 a_71281_n10073.n604 8.10567
R53288 a_71281_n10073.n605 a_71281_n10073.t229 8.10567
R53289 a_71281_n10073.t217 a_71281_n10073.n618 8.10567
R53290 a_71281_n10073.n619 a_71281_n10073.t217 8.10567
R53291 a_71281_n10073.t301 a_71281_n10073.n632 8.10567
R53292 a_71281_n10073.n633 a_71281_n10073.t301 8.10567
R53293 a_71281_n10073.n764 a_71281_n10073.t164 8.10567
R53294 a_71281_n10073.t164 a_71281_n10073.n763 8.10567
R53295 a_71281_n10073.n750 a_71281_n10073.t136 8.10567
R53296 a_71281_n10073.t136 a_71281_n10073.n749 8.10567
R53297 a_71281_n10073.n736 a_71281_n10073.t147 8.10567
R53298 a_71281_n10073.t147 a_71281_n10073.n735 8.10567
R53299 a_71281_n10073.n719 a_71281_n10073.t52 8.10567
R53300 a_71281_n10073.t52 a_71281_n10073.n718 8.10567
R53301 a_71281_n10073.n705 a_71281_n10073.t30 8.10567
R53302 a_71281_n10073.t30 a_71281_n10073.n704 8.10567
R53303 a_71281_n10073.n688 a_71281_n10073.t193 8.10567
R53304 a_71281_n10073.t193 a_71281_n10073.n687 8.10567
R53305 a_71281_n10073.n674 a_71281_n10073.t275 8.10567
R53306 a_71281_n10073.t275 a_71281_n10073.n673 8.10567
R53307 a_71281_n10073.n660 a_71281_n10073.t140 8.10567
R53308 a_71281_n10073.t140 a_71281_n10073.n659 8.10567
R53309 a_71281_n10073.n646 a_71281_n10073.t205 8.10567
R53310 a_71281_n10073.t205 a_71281_n10073.n645 8.10567
R53311 a_71281_n10073.n501 a_71281_n10073.t258 8.10567
R53312 a_71281_n10073.t258 a_71281_n10073.n500 8.10567
R53313 a_71281_n10073.t97 a_71281_n10073.n777 8.10567
R53314 a_71281_n10073.n778 a_71281_n10073.t97 8.10567
R53315 a_71281_n10073.t248 a_71281_n10073.n196 8.10567
R53316 a_71281_n10073.n197 a_71281_n10073.t248 8.10567
R53317 a_71281_n10073.n143 a_71281_n10073.t59 6.12845
R53318 a_71281_n10073.n257 a_71281_n10073.t17 6.12845
R53319 a_71281_n10073.n433 a_71281_n10073.t25 6.12845
R53320 a_71281_n10073.n548 a_71281_n10073.t57 6.12845
R53321 a_71281_n10073.n724 a_71281_n10073.t27 6.12845
R53322 a_71281_n10073.n874 a_71281_n10073.t43 6.12845
R53323 a_71281_n10073.n843 a_71281_n10073.t47 6.12049
R53324 a_71281_n10073.n288 a_71281_n10073.t45 6.12049
R53325 a_71281_n10073.n402 a_71281_n10073.t33 6.12049
R53326 a_71281_n10073.n579 a_71281_n10073.t69 6.12049
R53327 a_71281_n10073.n693 a_71281_n10073.t21 6.12049
R53328 a_71281_n10073.n112 a_71281_n10073.t13 6.12049
R53329 a_71281_n10073.n23 a_71281_n10073.n19 4.64734
R53330 a_71281_n10073.n24 a_71281_n10073.n15 4.64734
R53331 a_71281_n10073.n37 a_71281_n10073.n33 4.64734
R53332 a_71281_n10073.n38 a_71281_n10073.n29 4.64734
R53333 a_71281_n10073.n51 a_71281_n10073.n47 4.64734
R53334 a_71281_n10073.n52 a_71281_n10073.n43 4.64734
R53335 a_71281_n10073.n869 a_71281_n10073.n860 4.64734
R53336 a_71281_n10073.n868 a_71281_n10073.n864 4.64734
R53337 a_71281_n10073.n855 a_71281_n10073.n846 4.64734
R53338 a_71281_n10073.n854 a_71281_n10073.n850 4.64734
R53339 a_71281_n10073.n838 a_71281_n10073.n829 4.64734
R53340 a_71281_n10073.n837 a_71281_n10073.n833 4.64734
R53341 a_71281_n10073.n824 a_71281_n10073.n815 4.64734
R53342 a_71281_n10073.n823 a_71281_n10073.n819 4.64734
R53343 a_71281_n10073.n810 a_71281_n10073.n801 4.64734
R53344 a_71281_n10073.n809 a_71281_n10073.n805 4.64734
R53345 a_71281_n10073.n796 a_71281_n10073.n787 4.64734
R53346 a_71281_n10073.n795 a_71281_n10073.n791 4.64734
R53347 a_71281_n10073.n183 a_71281_n10073.n174 4.64734
R53348 a_71281_n10073.n182 a_71281_n10073.n178 4.64734
R53349 a_71281_n10073.n169 a_71281_n10073.n160 4.64734
R53350 a_71281_n10073.n168 a_71281_n10073.n164 4.64734
R53351 a_71281_n10073.n155 a_71281_n10073.n146 4.64734
R53352 a_71281_n10073.n154 a_71281_n10073.n150 4.64734
R53353 a_71281_n10073.n138 a_71281_n10073.n129 4.64734
R53354 a_71281_n10073.n137 a_71281_n10073.n133 4.64734
R53355 a_71281_n10073.n124 a_71281_n10073.n115 4.64734
R53356 a_71281_n10073.n123 a_71281_n10073.n119 4.64734
R53357 a_71281_n10073.n107 a_71281_n10073.n98 4.64734
R53358 a_71281_n10073.n106 a_71281_n10073.n102 4.64734
R53359 a_71281_n10073.n93 a_71281_n10073.n84 4.64734
R53360 a_71281_n10073.n92 a_71281_n10073.n88 4.64734
R53361 a_71281_n10073.n79 a_71281_n10073.n70 4.64734
R53362 a_71281_n10073.n78 a_71281_n10073.n74 4.64734
R53363 a_71281_n10073.n65 a_71281_n10073.n57 4.64734
R53364 a_71281_n10073.n64 a_71281_n10073.n61 4.64734
R53365 a_71281_n10073.n10 a_71281_n10073.n2 4.64734
R53366 a_71281_n10073.n9 a_71281_n10073.n6 4.64734
R53367 a_71281_n10073.n223 a_71281_n10073.n219 4.64734
R53368 a_71281_n10073.n224 a_71281_n10073.n215 4.64734
R53369 a_71281_n10073.n237 a_71281_n10073.n233 4.64734
R53370 a_71281_n10073.n238 a_71281_n10073.n229 4.64734
R53371 a_71281_n10073.n251 a_71281_n10073.n247 4.64734
R53372 a_71281_n10073.n252 a_71281_n10073.n243 4.64734
R53373 a_71281_n10073.n268 a_71281_n10073.n264 4.64734
R53374 a_71281_n10073.n269 a_71281_n10073.n260 4.64734
R53375 a_71281_n10073.n282 a_71281_n10073.n278 4.64734
R53376 a_71281_n10073.n283 a_71281_n10073.n274 4.64734
R53377 a_71281_n10073.n299 a_71281_n10073.n295 4.64734
R53378 a_71281_n10073.n300 a_71281_n10073.n291 4.64734
R53379 a_71281_n10073.n313 a_71281_n10073.n309 4.64734
R53380 a_71281_n10073.n314 a_71281_n10073.n305 4.64734
R53381 a_71281_n10073.n327 a_71281_n10073.n323 4.64734
R53382 a_71281_n10073.n328 a_71281_n10073.n319 4.64734
R53383 a_71281_n10073.n341 a_71281_n10073.n337 4.64734
R53384 a_71281_n10073.n342 a_71281_n10073.n333 4.64734
R53385 a_71281_n10073.n473 a_71281_n10073.n464 4.64734
R53386 a_71281_n10073.n472 a_71281_n10073.n468 4.64734
R53387 a_71281_n10073.n459 a_71281_n10073.n450 4.64734
R53388 a_71281_n10073.n458 a_71281_n10073.n454 4.64734
R53389 a_71281_n10073.n445 a_71281_n10073.n436 4.64734
R53390 a_71281_n10073.n444 a_71281_n10073.n440 4.64734
R53391 a_71281_n10073.n428 a_71281_n10073.n419 4.64734
R53392 a_71281_n10073.n427 a_71281_n10073.n423 4.64734
R53393 a_71281_n10073.n414 a_71281_n10073.n405 4.64734
R53394 a_71281_n10073.n413 a_71281_n10073.n409 4.64734
R53395 a_71281_n10073.n397 a_71281_n10073.n388 4.64734
R53396 a_71281_n10073.n396 a_71281_n10073.n392 4.64734
R53397 a_71281_n10073.n383 a_71281_n10073.n374 4.64734
R53398 a_71281_n10073.n382 a_71281_n10073.n378 4.64734
R53399 a_71281_n10073.n369 a_71281_n10073.n360 4.64734
R53400 a_71281_n10073.n368 a_71281_n10073.n364 4.64734
R53401 a_71281_n10073.n355 a_71281_n10073.n347 4.64734
R53402 a_71281_n10073.n354 a_71281_n10073.n351 4.64734
R53403 a_71281_n10073.n210 a_71281_n10073.n202 4.64734
R53404 a_71281_n10073.n209 a_71281_n10073.n206 4.64734
R53405 a_71281_n10073.n486 a_71281_n10073.n482 4.64734
R53406 a_71281_n10073.n487 a_71281_n10073.n478 4.64734
R53407 a_71281_n10073.n514 a_71281_n10073.n510 4.64734
R53408 a_71281_n10073.n515 a_71281_n10073.n506 4.64734
R53409 a_71281_n10073.n528 a_71281_n10073.n524 4.64734
R53410 a_71281_n10073.n529 a_71281_n10073.n520 4.64734
R53411 a_71281_n10073.n542 a_71281_n10073.n538 4.64734
R53412 a_71281_n10073.n543 a_71281_n10073.n534 4.64734
R53413 a_71281_n10073.n559 a_71281_n10073.n555 4.64734
R53414 a_71281_n10073.n560 a_71281_n10073.n551 4.64734
R53415 a_71281_n10073.n573 a_71281_n10073.n569 4.64734
R53416 a_71281_n10073.n574 a_71281_n10073.n565 4.64734
R53417 a_71281_n10073.n590 a_71281_n10073.n586 4.64734
R53418 a_71281_n10073.n591 a_71281_n10073.n582 4.64734
R53419 a_71281_n10073.n604 a_71281_n10073.n600 4.64734
R53420 a_71281_n10073.n605 a_71281_n10073.n596 4.64734
R53421 a_71281_n10073.n618 a_71281_n10073.n614 4.64734
R53422 a_71281_n10073.n619 a_71281_n10073.n610 4.64734
R53423 a_71281_n10073.n632 a_71281_n10073.n628 4.64734
R53424 a_71281_n10073.n633 a_71281_n10073.n624 4.64734
R53425 a_71281_n10073.n764 a_71281_n10073.n755 4.64734
R53426 a_71281_n10073.n763 a_71281_n10073.n759 4.64734
R53427 a_71281_n10073.n750 a_71281_n10073.n741 4.64734
R53428 a_71281_n10073.n749 a_71281_n10073.n745 4.64734
R53429 a_71281_n10073.n736 a_71281_n10073.n727 4.64734
R53430 a_71281_n10073.n735 a_71281_n10073.n731 4.64734
R53431 a_71281_n10073.n719 a_71281_n10073.n710 4.64734
R53432 a_71281_n10073.n718 a_71281_n10073.n714 4.64734
R53433 a_71281_n10073.n705 a_71281_n10073.n696 4.64734
R53434 a_71281_n10073.n704 a_71281_n10073.n700 4.64734
R53435 a_71281_n10073.n688 a_71281_n10073.n679 4.64734
R53436 a_71281_n10073.n687 a_71281_n10073.n683 4.64734
R53437 a_71281_n10073.n674 a_71281_n10073.n665 4.64734
R53438 a_71281_n10073.n673 a_71281_n10073.n669 4.64734
R53439 a_71281_n10073.n660 a_71281_n10073.n651 4.64734
R53440 a_71281_n10073.n659 a_71281_n10073.n655 4.64734
R53441 a_71281_n10073.n646 a_71281_n10073.n638 4.64734
R53442 a_71281_n10073.n645 a_71281_n10073.n642 4.64734
R53443 a_71281_n10073.n501 a_71281_n10073.n493 4.64734
R53444 a_71281_n10073.n500 a_71281_n10073.n497 4.64734
R53445 a_71281_n10073.n777 a_71281_n10073.n773 4.64734
R53446 a_71281_n10073.n778 a_71281_n10073.n769 4.64734
R53447 a_71281_n10073.n196 a_71281_n10073.n192 4.64734
R53448 a_71281_n10073.n197 a_71281_n10073.n188 4.64734
R53449 a_71281_n10073.n784 a_71281_n10073.n0 18.9036
R53450 a_71281_n10073.n843 a_71281_n10073.n842 4.01884
R53451 a_71281_n10073.n288 a_71281_n10073.n287 4.01884
R53452 a_71281_n10073.n402 a_71281_n10073.n401 4.01884
R53453 a_71281_n10073.n579 a_71281_n10073.n578 4.01884
R53454 a_71281_n10073.n693 a_71281_n10073.n692 4.01884
R53455 a_71281_n10073.n112 a_71281_n10073.n111 4.01884
R53456 a_71281_n10073.n143 a_71281_n10073.n142 4.00982
R53457 a_71281_n10073.n257 a_71281_n10073.n256 4.00982
R53458 a_71281_n10073.n433 a_71281_n10073.n432 4.00982
R53459 a_71281_n10073.n548 a_71281_n10073.n547 4.00982
R53460 a_71281_n10073.n724 a_71281_n10073.n723 4.00982
R53461 a_71281_n10073.n875 a_71281_n10073.n874 4.00982
R53462 a_71281_n10073.n0 a_71281_n10073.t73 3.7215
R53463 a_71281_n10073.n783 a_71281_n10073.n491 3.61592
R53464 a_71281_n10073.n784 a_71281_n10073.n783 2.86491
R53465 a_71281_n10073.n25 a_71281_n10073.n24 2.25278
R53466 a_71281_n10073.n23 a_71281_n10073.n22 2.25278
R53467 a_71281_n10073.n39 a_71281_n10073.n38 2.25278
R53468 a_71281_n10073.n37 a_71281_n10073.n36 2.25278
R53469 a_71281_n10073.n53 a_71281_n10073.n52 2.25278
R53470 a_71281_n10073.n51 a_71281_n10073.n50 2.25278
R53471 a_71281_n10073.n868 a_71281_n10073.n867 2.25278
R53472 a_71281_n10073.n870 a_71281_n10073.n869 2.25278
R53473 a_71281_n10073.n854 a_71281_n10073.n853 2.25278
R53474 a_71281_n10073.n856 a_71281_n10073.n855 2.25278
R53475 a_71281_n10073.n837 a_71281_n10073.n836 2.25278
R53476 a_71281_n10073.n839 a_71281_n10073.n838 2.25278
R53477 a_71281_n10073.n823 a_71281_n10073.n822 2.25278
R53478 a_71281_n10073.n825 a_71281_n10073.n824 2.25278
R53479 a_71281_n10073.n809 a_71281_n10073.n808 2.25278
R53480 a_71281_n10073.n811 a_71281_n10073.n810 2.25278
R53481 a_71281_n10073.n795 a_71281_n10073.n794 2.25278
R53482 a_71281_n10073.n797 a_71281_n10073.n796 2.25278
R53483 a_71281_n10073.n182 a_71281_n10073.n181 2.25278
R53484 a_71281_n10073.n184 a_71281_n10073.n183 2.25278
R53485 a_71281_n10073.n168 a_71281_n10073.n167 2.25278
R53486 a_71281_n10073.n170 a_71281_n10073.n169 2.25278
R53487 a_71281_n10073.n154 a_71281_n10073.n153 2.25278
R53488 a_71281_n10073.n156 a_71281_n10073.n155 2.25278
R53489 a_71281_n10073.n137 a_71281_n10073.n136 2.25278
R53490 a_71281_n10073.n139 a_71281_n10073.n138 2.25278
R53491 a_71281_n10073.n123 a_71281_n10073.n122 2.25278
R53492 a_71281_n10073.n125 a_71281_n10073.n124 2.25278
R53493 a_71281_n10073.n106 a_71281_n10073.n105 2.25278
R53494 a_71281_n10073.n108 a_71281_n10073.n107 2.25278
R53495 a_71281_n10073.n92 a_71281_n10073.n91 2.25278
R53496 a_71281_n10073.n94 a_71281_n10073.n93 2.25278
R53497 a_71281_n10073.n78 a_71281_n10073.n77 2.25278
R53498 a_71281_n10073.n80 a_71281_n10073.n79 2.25278
R53499 a_71281_n10073.n64 a_71281_n10073.n63 2.25278
R53500 a_71281_n10073.n66 a_71281_n10073.n65 2.25278
R53501 a_71281_n10073.n9 a_71281_n10073.n8 2.25278
R53502 a_71281_n10073.n11 a_71281_n10073.n10 2.25278
R53503 a_71281_n10073.n225 a_71281_n10073.n224 2.25278
R53504 a_71281_n10073.n223 a_71281_n10073.n222 2.25278
R53505 a_71281_n10073.n239 a_71281_n10073.n238 2.25278
R53506 a_71281_n10073.n237 a_71281_n10073.n236 2.25278
R53507 a_71281_n10073.n253 a_71281_n10073.n252 2.25278
R53508 a_71281_n10073.n251 a_71281_n10073.n250 2.25278
R53509 a_71281_n10073.n270 a_71281_n10073.n269 2.25278
R53510 a_71281_n10073.n268 a_71281_n10073.n267 2.25278
R53511 a_71281_n10073.n284 a_71281_n10073.n283 2.25278
R53512 a_71281_n10073.n282 a_71281_n10073.n281 2.25278
R53513 a_71281_n10073.n301 a_71281_n10073.n300 2.25278
R53514 a_71281_n10073.n299 a_71281_n10073.n298 2.25278
R53515 a_71281_n10073.n315 a_71281_n10073.n314 2.25278
R53516 a_71281_n10073.n313 a_71281_n10073.n312 2.25278
R53517 a_71281_n10073.n329 a_71281_n10073.n328 2.25278
R53518 a_71281_n10073.n327 a_71281_n10073.n326 2.25278
R53519 a_71281_n10073.n343 a_71281_n10073.n342 2.25278
R53520 a_71281_n10073.n341 a_71281_n10073.n340 2.25278
R53521 a_71281_n10073.n472 a_71281_n10073.n471 2.25278
R53522 a_71281_n10073.n474 a_71281_n10073.n473 2.25278
R53523 a_71281_n10073.n458 a_71281_n10073.n457 2.25278
R53524 a_71281_n10073.n460 a_71281_n10073.n459 2.25278
R53525 a_71281_n10073.n444 a_71281_n10073.n443 2.25278
R53526 a_71281_n10073.n446 a_71281_n10073.n445 2.25278
R53527 a_71281_n10073.n427 a_71281_n10073.n426 2.25278
R53528 a_71281_n10073.n429 a_71281_n10073.n428 2.25278
R53529 a_71281_n10073.n413 a_71281_n10073.n412 2.25278
R53530 a_71281_n10073.n415 a_71281_n10073.n414 2.25278
R53531 a_71281_n10073.n396 a_71281_n10073.n395 2.25278
R53532 a_71281_n10073.n398 a_71281_n10073.n397 2.25278
R53533 a_71281_n10073.n382 a_71281_n10073.n381 2.25278
R53534 a_71281_n10073.n384 a_71281_n10073.n383 2.25278
R53535 a_71281_n10073.n368 a_71281_n10073.n367 2.25278
R53536 a_71281_n10073.n370 a_71281_n10073.n369 2.25278
R53537 a_71281_n10073.n354 a_71281_n10073.n353 2.25278
R53538 a_71281_n10073.n356 a_71281_n10073.n355 2.25278
R53539 a_71281_n10073.n209 a_71281_n10073.n208 2.25278
R53540 a_71281_n10073.n211 a_71281_n10073.n210 2.25278
R53541 a_71281_n10073.n488 a_71281_n10073.n487 2.25278
R53542 a_71281_n10073.n486 a_71281_n10073.n485 2.25278
R53543 a_71281_n10073.n516 a_71281_n10073.n515 2.25278
R53544 a_71281_n10073.n514 a_71281_n10073.n513 2.25278
R53545 a_71281_n10073.n530 a_71281_n10073.n529 2.25278
R53546 a_71281_n10073.n528 a_71281_n10073.n527 2.25278
R53547 a_71281_n10073.n544 a_71281_n10073.n543 2.25278
R53548 a_71281_n10073.n542 a_71281_n10073.n541 2.25278
R53549 a_71281_n10073.n561 a_71281_n10073.n560 2.25278
R53550 a_71281_n10073.n559 a_71281_n10073.n558 2.25278
R53551 a_71281_n10073.n575 a_71281_n10073.n574 2.25278
R53552 a_71281_n10073.n573 a_71281_n10073.n572 2.25278
R53553 a_71281_n10073.n592 a_71281_n10073.n591 2.25278
R53554 a_71281_n10073.n590 a_71281_n10073.n589 2.25278
R53555 a_71281_n10073.n606 a_71281_n10073.n605 2.25278
R53556 a_71281_n10073.n604 a_71281_n10073.n603 2.25278
R53557 a_71281_n10073.n620 a_71281_n10073.n619 2.25278
R53558 a_71281_n10073.n618 a_71281_n10073.n617 2.25278
R53559 a_71281_n10073.n634 a_71281_n10073.n633 2.25278
R53560 a_71281_n10073.n632 a_71281_n10073.n631 2.25278
R53561 a_71281_n10073.n763 a_71281_n10073.n762 2.25278
R53562 a_71281_n10073.n765 a_71281_n10073.n764 2.25278
R53563 a_71281_n10073.n749 a_71281_n10073.n748 2.25278
R53564 a_71281_n10073.n751 a_71281_n10073.n750 2.25278
R53565 a_71281_n10073.n735 a_71281_n10073.n734 2.25278
R53566 a_71281_n10073.n737 a_71281_n10073.n736 2.25278
R53567 a_71281_n10073.n718 a_71281_n10073.n717 2.25278
R53568 a_71281_n10073.n720 a_71281_n10073.n719 2.25278
R53569 a_71281_n10073.n704 a_71281_n10073.n703 2.25278
R53570 a_71281_n10073.n706 a_71281_n10073.n705 2.25278
R53571 a_71281_n10073.n687 a_71281_n10073.n686 2.25278
R53572 a_71281_n10073.n689 a_71281_n10073.n688 2.25278
R53573 a_71281_n10073.n673 a_71281_n10073.n672 2.25278
R53574 a_71281_n10073.n675 a_71281_n10073.n674 2.25278
R53575 a_71281_n10073.n659 a_71281_n10073.n658 2.25278
R53576 a_71281_n10073.n661 a_71281_n10073.n660 2.25278
R53577 a_71281_n10073.n645 a_71281_n10073.n644 2.25278
R53578 a_71281_n10073.n647 a_71281_n10073.n646 2.25278
R53579 a_71281_n10073.n500 a_71281_n10073.n499 2.25278
R53580 a_71281_n10073.n502 a_71281_n10073.n501 2.25278
R53581 a_71281_n10073.n779 a_71281_n10073.n778 2.25278
R53582 a_71281_n10073.n777 a_71281_n10073.n776 2.25278
R53583 a_71281_n10073.n198 a_71281_n10073.n197 2.25278
R53584 a_71281_n10073.n196 a_71281_n10073.n195 2.25278
R53585 a_71281_n10073.n213 a_71281_n10073.n201 1.6802
R53586 a_71281_n10073.n358 a_71281_n10073.n346 1.6802
R53587 a_71281_n10073.n504 a_71281_n10073.n492 1.6802
R53588 a_71281_n10073.n649 a_71281_n10073.n637 1.6802
R53589 a_71281_n10073.n13 a_71281_n10073.n1 1.6802
R53590 a_71281_n10073.n68 a_71281_n10073.n56 1.6802
R53591 a_71281_n10073.n403 a_71281_n10073.n402 1.5005
R53592 a_71281_n10073.n483 a_71281_n10073.n477 1.5005
R53593 a_71281_n10073.n289 a_71281_n10073.n288 1.5005
R53594 a_71281_n10073.n213 a_71281_n10073.n212 1.5005
R53595 a_71281_n10073.n434 a_71281_n10073.n433 1.5005
R53596 a_71281_n10073.n258 a_71281_n10073.n257 1.5005
R53597 a_71281_n10073.n358 a_71281_n10073.n357 1.5005
R53598 a_71281_n10073.n372 a_71281_n10073.n371 1.5005
R53599 a_71281_n10073.n366 a_71281_n10073.n359 1.5005
R53600 a_71281_n10073.n386 a_71281_n10073.n385 1.5005
R53601 a_71281_n10073.n380 a_71281_n10073.n373 1.5005
R53602 a_71281_n10073.n400 a_71281_n10073.n399 1.5005
R53603 a_71281_n10073.n394 a_71281_n10073.n387 1.5005
R53604 a_71281_n10073.n417 a_71281_n10073.n416 1.5005
R53605 a_71281_n10073.n411 a_71281_n10073.n404 1.5005
R53606 a_71281_n10073.n431 a_71281_n10073.n430 1.5005
R53607 a_71281_n10073.n425 a_71281_n10073.n418 1.5005
R53608 a_71281_n10073.n448 a_71281_n10073.n447 1.5005
R53609 a_71281_n10073.n442 a_71281_n10073.n435 1.5005
R53610 a_71281_n10073.n462 a_71281_n10073.n461 1.5005
R53611 a_71281_n10073.n456 a_71281_n10073.n449 1.5005
R53612 a_71281_n10073.n476 a_71281_n10073.n475 1.5005
R53613 a_71281_n10073.n470 a_71281_n10073.n463 1.5005
R53614 a_71281_n10073.n490 a_71281_n10073.n489 1.5005
R53615 a_71281_n10073.n338 a_71281_n10073.n332 1.5005
R53616 a_71281_n10073.n345 a_71281_n10073.n344 1.5005
R53617 a_71281_n10073.n324 a_71281_n10073.n318 1.5005
R53618 a_71281_n10073.n331 a_71281_n10073.n330 1.5005
R53619 a_71281_n10073.n310 a_71281_n10073.n304 1.5005
R53620 a_71281_n10073.n317 a_71281_n10073.n316 1.5005
R53621 a_71281_n10073.n296 a_71281_n10073.n290 1.5005
R53622 a_71281_n10073.n303 a_71281_n10073.n302 1.5005
R53623 a_71281_n10073.n279 a_71281_n10073.n273 1.5005
R53624 a_71281_n10073.n286 a_71281_n10073.n285 1.5005
R53625 a_71281_n10073.n265 a_71281_n10073.n259 1.5005
R53626 a_71281_n10073.n272 a_71281_n10073.n271 1.5005
R53627 a_71281_n10073.n248 a_71281_n10073.n242 1.5005
R53628 a_71281_n10073.n255 a_71281_n10073.n254 1.5005
R53629 a_71281_n10073.n234 a_71281_n10073.n228 1.5005
R53630 a_71281_n10073.n241 a_71281_n10073.n240 1.5005
R53631 a_71281_n10073.n220 a_71281_n10073.n214 1.5005
R53632 a_71281_n10073.n227 a_71281_n10073.n226 1.5005
R53633 a_71281_n10073.n694 a_71281_n10073.n693 1.5005
R53634 a_71281_n10073.n774 a_71281_n10073.n768 1.5005
R53635 a_71281_n10073.n580 a_71281_n10073.n579 1.5005
R53636 a_71281_n10073.n504 a_71281_n10073.n503 1.5005
R53637 a_71281_n10073.n725 a_71281_n10073.n724 1.5005
R53638 a_71281_n10073.n549 a_71281_n10073.n548 1.5005
R53639 a_71281_n10073.n649 a_71281_n10073.n648 1.5005
R53640 a_71281_n10073.n663 a_71281_n10073.n662 1.5005
R53641 a_71281_n10073.n657 a_71281_n10073.n650 1.5005
R53642 a_71281_n10073.n677 a_71281_n10073.n676 1.5005
R53643 a_71281_n10073.n671 a_71281_n10073.n664 1.5005
R53644 a_71281_n10073.n691 a_71281_n10073.n690 1.5005
R53645 a_71281_n10073.n685 a_71281_n10073.n678 1.5005
R53646 a_71281_n10073.n708 a_71281_n10073.n707 1.5005
R53647 a_71281_n10073.n702 a_71281_n10073.n695 1.5005
R53648 a_71281_n10073.n722 a_71281_n10073.n721 1.5005
R53649 a_71281_n10073.n716 a_71281_n10073.n709 1.5005
R53650 a_71281_n10073.n739 a_71281_n10073.n738 1.5005
R53651 a_71281_n10073.n733 a_71281_n10073.n726 1.5005
R53652 a_71281_n10073.n753 a_71281_n10073.n752 1.5005
R53653 a_71281_n10073.n747 a_71281_n10073.n740 1.5005
R53654 a_71281_n10073.n767 a_71281_n10073.n766 1.5005
R53655 a_71281_n10073.n761 a_71281_n10073.n754 1.5005
R53656 a_71281_n10073.n781 a_71281_n10073.n780 1.5005
R53657 a_71281_n10073.n629 a_71281_n10073.n623 1.5005
R53658 a_71281_n10073.n636 a_71281_n10073.n635 1.5005
R53659 a_71281_n10073.n615 a_71281_n10073.n609 1.5005
R53660 a_71281_n10073.n622 a_71281_n10073.n621 1.5005
R53661 a_71281_n10073.n601 a_71281_n10073.n595 1.5005
R53662 a_71281_n10073.n608 a_71281_n10073.n607 1.5005
R53663 a_71281_n10073.n587 a_71281_n10073.n581 1.5005
R53664 a_71281_n10073.n594 a_71281_n10073.n593 1.5005
R53665 a_71281_n10073.n570 a_71281_n10073.n564 1.5005
R53666 a_71281_n10073.n577 a_71281_n10073.n576 1.5005
R53667 a_71281_n10073.n556 a_71281_n10073.n550 1.5005
R53668 a_71281_n10073.n563 a_71281_n10073.n562 1.5005
R53669 a_71281_n10073.n539 a_71281_n10073.n533 1.5005
R53670 a_71281_n10073.n546 a_71281_n10073.n545 1.5005
R53671 a_71281_n10073.n525 a_71281_n10073.n519 1.5005
R53672 a_71281_n10073.n532 a_71281_n10073.n531 1.5005
R53673 a_71281_n10073.n511 a_71281_n10073.n505 1.5005
R53674 a_71281_n10073.n518 a_71281_n10073.n517 1.5005
R53675 a_71281_n10073.n113 a_71281_n10073.n112 1.5005
R53676 a_71281_n10073.n193 a_71281_n10073.n187 1.5005
R53677 a_71281_n10073.n844 a_71281_n10073.n843 1.5005
R53678 a_71281_n10073.n13 a_71281_n10073.n12 1.5005
R53679 a_71281_n10073.n144 a_71281_n10073.n143 1.5005
R53680 a_71281_n10073.n68 a_71281_n10073.n67 1.5005
R53681 a_71281_n10073.n82 a_71281_n10073.n81 1.5005
R53682 a_71281_n10073.n76 a_71281_n10073.n69 1.5005
R53683 a_71281_n10073.n96 a_71281_n10073.n95 1.5005
R53684 a_71281_n10073.n90 a_71281_n10073.n83 1.5005
R53685 a_71281_n10073.n110 a_71281_n10073.n109 1.5005
R53686 a_71281_n10073.n104 a_71281_n10073.n97 1.5005
R53687 a_71281_n10073.n127 a_71281_n10073.n126 1.5005
R53688 a_71281_n10073.n121 a_71281_n10073.n114 1.5005
R53689 a_71281_n10073.n141 a_71281_n10073.n140 1.5005
R53690 a_71281_n10073.n135 a_71281_n10073.n128 1.5005
R53691 a_71281_n10073.n158 a_71281_n10073.n157 1.5005
R53692 a_71281_n10073.n152 a_71281_n10073.n145 1.5005
R53693 a_71281_n10073.n172 a_71281_n10073.n171 1.5005
R53694 a_71281_n10073.n166 a_71281_n10073.n159 1.5005
R53695 a_71281_n10073.n186 a_71281_n10073.n185 1.5005
R53696 a_71281_n10073.n180 a_71281_n10073.n173 1.5005
R53697 a_71281_n10073.n200 a_71281_n10073.n199 1.5005
R53698 a_71281_n10073.n799 a_71281_n10073.n798 1.5005
R53699 a_71281_n10073.n793 a_71281_n10073.n786 1.5005
R53700 a_71281_n10073.n813 a_71281_n10073.n812 1.5005
R53701 a_71281_n10073.n807 a_71281_n10073.n800 1.5005
R53702 a_71281_n10073.n827 a_71281_n10073.n826 1.5005
R53703 a_71281_n10073.n821 a_71281_n10073.n814 1.5005
R53704 a_71281_n10073.n841 a_71281_n10073.n840 1.5005
R53705 a_71281_n10073.n835 a_71281_n10073.n828 1.5005
R53706 a_71281_n10073.n858 a_71281_n10073.n857 1.5005
R53707 a_71281_n10073.n852 a_71281_n10073.n845 1.5005
R53708 a_71281_n10073.n872 a_71281_n10073.n871 1.5005
R53709 a_71281_n10073.n866 a_71281_n10073.n859 1.5005
R53710 a_71281_n10073.n48 a_71281_n10073.n42 1.5005
R53711 a_71281_n10073.n55 a_71281_n10073.n54 1.5005
R53712 a_71281_n10073.n34 a_71281_n10073.n28 1.5005
R53713 a_71281_n10073.n41 a_71281_n10073.n40 1.5005
R53714 a_71281_n10073.n20 a_71281_n10073.n14 1.5005
R53715 a_71281_n10073.n27 a_71281_n10073.n26 1.5005
R53716 a_71281_n10073.n874 a_71281_n10073.n873 1.5005
R53717 a_71281_n10073.n142 a_71281_n10073.t29 1.4705
R53718 a_71281_n10073.n142 a_71281_n10073.t7 1.4705
R53719 a_71281_n10073.n842 a_71281_n10073.t39 1.4705
R53720 a_71281_n10073.n842 a_71281_n10073.t15 1.4705
R53721 a_71281_n10073.n256 a_71281_n10073.t67 1.4705
R53722 a_71281_n10073.n256 a_71281_n10073.t51 1.4705
R53723 a_71281_n10073.n432 a_71281_n10073.t55 1.4705
R53724 a_71281_n10073.n432 a_71281_n10073.t19 1.4705
R53725 a_71281_n10073.n287 a_71281_n10073.t23 1.4705
R53726 a_71281_n10073.n287 a_71281_n10073.t1 1.4705
R53727 a_71281_n10073.n401 a_71281_n10073.t3 1.4705
R53728 a_71281_n10073.n401 a_71281_n10073.t5 1.4705
R53729 a_71281_n10073.n547 a_71281_n10073.t11 1.4705
R53730 a_71281_n10073.n547 a_71281_n10073.t63 1.4705
R53731 a_71281_n10073.n723 a_71281_n10073.t49 1.4705
R53732 a_71281_n10073.n723 a_71281_n10073.t53 1.4705
R53733 a_71281_n10073.n578 a_71281_n10073.t41 1.4705
R53734 a_71281_n10073.n578 a_71281_n10073.t35 1.4705
R53735 a_71281_n10073.n692 a_71281_n10073.t31 1.4705
R53736 a_71281_n10073.n692 a_71281_n10073.t9 1.4705
R53737 a_71281_n10073.n111 a_71281_n10073.t65 1.4705
R53738 a_71281_n10073.n111 a_71281_n10073.t37 1.4705
R53739 a_71281_n10073.t71 a_71281_n10073.n875 1.4705
R53740 a_71281_n10073.n875 a_71281_n10073.t61 1.4705
R53741 a_71281_n10073.n783 a_71281_n10073.n782 0.7505
R53742 a_71281_n10073.n785 a_71281_n10073.n784 0.7505
R53743 a_71281_n10073.n25 a_71281_n10073.n16 0.567403
R53744 a_71281_n10073.n22 a_71281_n10073.n21 0.567403
R53745 a_71281_n10073.n39 a_71281_n10073.n30 0.567403
R53746 a_71281_n10073.n36 a_71281_n10073.n35 0.567403
R53747 a_71281_n10073.n53 a_71281_n10073.n44 0.567403
R53748 a_71281_n10073.n50 a_71281_n10073.n49 0.567403
R53749 a_71281_n10073.n867 a_71281_n10073.n865 0.567403
R53750 a_71281_n10073.n870 a_71281_n10073.n861 0.567403
R53751 a_71281_n10073.n853 a_71281_n10073.n851 0.567403
R53752 a_71281_n10073.n856 a_71281_n10073.n847 0.567403
R53753 a_71281_n10073.n836 a_71281_n10073.n834 0.567403
R53754 a_71281_n10073.n839 a_71281_n10073.n830 0.567403
R53755 a_71281_n10073.n822 a_71281_n10073.n820 0.567403
R53756 a_71281_n10073.n825 a_71281_n10073.n816 0.567403
R53757 a_71281_n10073.n808 a_71281_n10073.n806 0.567403
R53758 a_71281_n10073.n811 a_71281_n10073.n802 0.567403
R53759 a_71281_n10073.n794 a_71281_n10073.n792 0.567403
R53760 a_71281_n10073.n797 a_71281_n10073.n788 0.567403
R53761 a_71281_n10073.n181 a_71281_n10073.n179 0.567403
R53762 a_71281_n10073.n184 a_71281_n10073.n175 0.567403
R53763 a_71281_n10073.n167 a_71281_n10073.n165 0.567403
R53764 a_71281_n10073.n170 a_71281_n10073.n161 0.567403
R53765 a_71281_n10073.n153 a_71281_n10073.n151 0.567403
R53766 a_71281_n10073.n156 a_71281_n10073.n147 0.567403
R53767 a_71281_n10073.n136 a_71281_n10073.n134 0.567403
R53768 a_71281_n10073.n139 a_71281_n10073.n130 0.567403
R53769 a_71281_n10073.n122 a_71281_n10073.n120 0.567403
R53770 a_71281_n10073.n125 a_71281_n10073.n116 0.567403
R53771 a_71281_n10073.n105 a_71281_n10073.n103 0.567403
R53772 a_71281_n10073.n108 a_71281_n10073.n99 0.567403
R53773 a_71281_n10073.n91 a_71281_n10073.n89 0.567403
R53774 a_71281_n10073.n94 a_71281_n10073.n85 0.567403
R53775 a_71281_n10073.n77 a_71281_n10073.n75 0.567403
R53776 a_71281_n10073.n80 a_71281_n10073.n71 0.567403
R53777 a_71281_n10073.n63 a_71281_n10073.n62 0.567403
R53778 a_71281_n10073.n66 a_71281_n10073.n58 0.567403
R53779 a_71281_n10073.n8 a_71281_n10073.n7 0.567403
R53780 a_71281_n10073.n11 a_71281_n10073.n3 0.567403
R53781 a_71281_n10073.n225 a_71281_n10073.n216 0.567403
R53782 a_71281_n10073.n222 a_71281_n10073.n221 0.567403
R53783 a_71281_n10073.n239 a_71281_n10073.n230 0.567403
R53784 a_71281_n10073.n236 a_71281_n10073.n235 0.567403
R53785 a_71281_n10073.n253 a_71281_n10073.n244 0.567403
R53786 a_71281_n10073.n250 a_71281_n10073.n249 0.567403
R53787 a_71281_n10073.n270 a_71281_n10073.n261 0.567403
R53788 a_71281_n10073.n267 a_71281_n10073.n266 0.567403
R53789 a_71281_n10073.n284 a_71281_n10073.n275 0.567403
R53790 a_71281_n10073.n281 a_71281_n10073.n280 0.567403
R53791 a_71281_n10073.n301 a_71281_n10073.n292 0.567403
R53792 a_71281_n10073.n298 a_71281_n10073.n297 0.567403
R53793 a_71281_n10073.n315 a_71281_n10073.n306 0.567403
R53794 a_71281_n10073.n312 a_71281_n10073.n311 0.567403
R53795 a_71281_n10073.n329 a_71281_n10073.n320 0.567403
R53796 a_71281_n10073.n326 a_71281_n10073.n325 0.567403
R53797 a_71281_n10073.n343 a_71281_n10073.n334 0.567403
R53798 a_71281_n10073.n340 a_71281_n10073.n339 0.567403
R53799 a_71281_n10073.n471 a_71281_n10073.n469 0.567403
R53800 a_71281_n10073.n474 a_71281_n10073.n465 0.567403
R53801 a_71281_n10073.n457 a_71281_n10073.n455 0.567403
R53802 a_71281_n10073.n460 a_71281_n10073.n451 0.567403
R53803 a_71281_n10073.n443 a_71281_n10073.n441 0.567403
R53804 a_71281_n10073.n446 a_71281_n10073.n437 0.567403
R53805 a_71281_n10073.n426 a_71281_n10073.n424 0.567403
R53806 a_71281_n10073.n429 a_71281_n10073.n420 0.567403
R53807 a_71281_n10073.n412 a_71281_n10073.n410 0.567403
R53808 a_71281_n10073.n415 a_71281_n10073.n406 0.567403
R53809 a_71281_n10073.n395 a_71281_n10073.n393 0.567403
R53810 a_71281_n10073.n398 a_71281_n10073.n389 0.567403
R53811 a_71281_n10073.n381 a_71281_n10073.n379 0.567403
R53812 a_71281_n10073.n384 a_71281_n10073.n375 0.567403
R53813 a_71281_n10073.n367 a_71281_n10073.n365 0.567403
R53814 a_71281_n10073.n370 a_71281_n10073.n361 0.567403
R53815 a_71281_n10073.n353 a_71281_n10073.n352 0.567403
R53816 a_71281_n10073.n356 a_71281_n10073.n348 0.567403
R53817 a_71281_n10073.n208 a_71281_n10073.n207 0.567403
R53818 a_71281_n10073.n211 a_71281_n10073.n203 0.567403
R53819 a_71281_n10073.n488 a_71281_n10073.n479 0.567403
R53820 a_71281_n10073.n485 a_71281_n10073.n484 0.567403
R53821 a_71281_n10073.n516 a_71281_n10073.n507 0.567403
R53822 a_71281_n10073.n513 a_71281_n10073.n512 0.567403
R53823 a_71281_n10073.n530 a_71281_n10073.n521 0.567403
R53824 a_71281_n10073.n527 a_71281_n10073.n526 0.567403
R53825 a_71281_n10073.n544 a_71281_n10073.n535 0.567403
R53826 a_71281_n10073.n541 a_71281_n10073.n540 0.567403
R53827 a_71281_n10073.n561 a_71281_n10073.n552 0.567403
R53828 a_71281_n10073.n558 a_71281_n10073.n557 0.567403
R53829 a_71281_n10073.n575 a_71281_n10073.n566 0.567403
R53830 a_71281_n10073.n572 a_71281_n10073.n571 0.567403
R53831 a_71281_n10073.n592 a_71281_n10073.n583 0.567403
R53832 a_71281_n10073.n589 a_71281_n10073.n588 0.567403
R53833 a_71281_n10073.n606 a_71281_n10073.n597 0.567403
R53834 a_71281_n10073.n603 a_71281_n10073.n602 0.567403
R53835 a_71281_n10073.n620 a_71281_n10073.n611 0.567403
R53836 a_71281_n10073.n617 a_71281_n10073.n616 0.567403
R53837 a_71281_n10073.n634 a_71281_n10073.n625 0.567403
R53838 a_71281_n10073.n631 a_71281_n10073.n630 0.567403
R53839 a_71281_n10073.n762 a_71281_n10073.n760 0.567403
R53840 a_71281_n10073.n765 a_71281_n10073.n756 0.567403
R53841 a_71281_n10073.n748 a_71281_n10073.n746 0.567403
R53842 a_71281_n10073.n751 a_71281_n10073.n742 0.567403
R53843 a_71281_n10073.n734 a_71281_n10073.n732 0.567403
R53844 a_71281_n10073.n737 a_71281_n10073.n728 0.567403
R53845 a_71281_n10073.n717 a_71281_n10073.n715 0.567403
R53846 a_71281_n10073.n720 a_71281_n10073.n711 0.567403
R53847 a_71281_n10073.n703 a_71281_n10073.n701 0.567403
R53848 a_71281_n10073.n706 a_71281_n10073.n697 0.567403
R53849 a_71281_n10073.n686 a_71281_n10073.n684 0.567403
R53850 a_71281_n10073.n689 a_71281_n10073.n680 0.567403
R53851 a_71281_n10073.n672 a_71281_n10073.n670 0.567403
R53852 a_71281_n10073.n675 a_71281_n10073.n666 0.567403
R53853 a_71281_n10073.n658 a_71281_n10073.n656 0.567403
R53854 a_71281_n10073.n661 a_71281_n10073.n652 0.567403
R53855 a_71281_n10073.n644 a_71281_n10073.n643 0.567403
R53856 a_71281_n10073.n647 a_71281_n10073.n639 0.567403
R53857 a_71281_n10073.n499 a_71281_n10073.n498 0.567403
R53858 a_71281_n10073.n502 a_71281_n10073.n494 0.567403
R53859 a_71281_n10073.n779 a_71281_n10073.n770 0.567403
R53860 a_71281_n10073.n776 a_71281_n10073.n775 0.567403
R53861 a_71281_n10073.n198 a_71281_n10073.n189 0.567403
R53862 a_71281_n10073.n195 a_71281_n10073.n194 0.567403
R53863 a_71281_n10073.n17 a_71281_n10073.n15 0.496742
R53864 a_71281_n10073.n19 a_71281_n10073.n18 0.496742
R53865 a_71281_n10073.n31 a_71281_n10073.n29 0.496742
R53866 a_71281_n10073.n33 a_71281_n10073.n32 0.496742
R53867 a_71281_n10073.n45 a_71281_n10073.n43 0.496742
R53868 a_71281_n10073.n47 a_71281_n10073.n46 0.496742
R53869 a_71281_n10073.n864 a_71281_n10073.n863 0.496742
R53870 a_71281_n10073.n862 a_71281_n10073.n860 0.496742
R53871 a_71281_n10073.n850 a_71281_n10073.n849 0.496742
R53872 a_71281_n10073.n848 a_71281_n10073.n846 0.496742
R53873 a_71281_n10073.n833 a_71281_n10073.n832 0.496742
R53874 a_71281_n10073.n831 a_71281_n10073.n829 0.496742
R53875 a_71281_n10073.n819 a_71281_n10073.n818 0.496742
R53876 a_71281_n10073.n817 a_71281_n10073.n815 0.496742
R53877 a_71281_n10073.n805 a_71281_n10073.n804 0.496742
R53878 a_71281_n10073.n803 a_71281_n10073.n801 0.496742
R53879 a_71281_n10073.n791 a_71281_n10073.n790 0.496742
R53880 a_71281_n10073.n789 a_71281_n10073.n787 0.496742
R53881 a_71281_n10073.n178 a_71281_n10073.n177 0.496742
R53882 a_71281_n10073.n176 a_71281_n10073.n174 0.496742
R53883 a_71281_n10073.n164 a_71281_n10073.n163 0.496742
R53884 a_71281_n10073.n162 a_71281_n10073.n160 0.496742
R53885 a_71281_n10073.n150 a_71281_n10073.n149 0.496742
R53886 a_71281_n10073.n148 a_71281_n10073.n146 0.496742
R53887 a_71281_n10073.n133 a_71281_n10073.n132 0.496742
R53888 a_71281_n10073.n131 a_71281_n10073.n129 0.496742
R53889 a_71281_n10073.n119 a_71281_n10073.n118 0.496742
R53890 a_71281_n10073.n117 a_71281_n10073.n115 0.496742
R53891 a_71281_n10073.n102 a_71281_n10073.n101 0.496742
R53892 a_71281_n10073.n100 a_71281_n10073.n98 0.496742
R53893 a_71281_n10073.n88 a_71281_n10073.n87 0.496742
R53894 a_71281_n10073.n86 a_71281_n10073.n84 0.496742
R53895 a_71281_n10073.n74 a_71281_n10073.n73 0.496742
R53896 a_71281_n10073.n72 a_71281_n10073.n70 0.496742
R53897 a_71281_n10073.n61 a_71281_n10073.n60 0.496742
R53898 a_71281_n10073.n59 a_71281_n10073.n57 0.496742
R53899 a_71281_n10073.n6 a_71281_n10073.n5 0.496742
R53900 a_71281_n10073.n4 a_71281_n10073.n2 0.496742
R53901 a_71281_n10073.n217 a_71281_n10073.n215 0.496742
R53902 a_71281_n10073.n219 a_71281_n10073.n218 0.496742
R53903 a_71281_n10073.n231 a_71281_n10073.n229 0.496742
R53904 a_71281_n10073.n233 a_71281_n10073.n232 0.496742
R53905 a_71281_n10073.n245 a_71281_n10073.n243 0.496742
R53906 a_71281_n10073.n247 a_71281_n10073.n246 0.496742
R53907 a_71281_n10073.n262 a_71281_n10073.n260 0.496742
R53908 a_71281_n10073.n264 a_71281_n10073.n263 0.496742
R53909 a_71281_n10073.n276 a_71281_n10073.n274 0.496742
R53910 a_71281_n10073.n278 a_71281_n10073.n277 0.496742
R53911 a_71281_n10073.n293 a_71281_n10073.n291 0.496742
R53912 a_71281_n10073.n295 a_71281_n10073.n294 0.496742
R53913 a_71281_n10073.n307 a_71281_n10073.n305 0.496742
R53914 a_71281_n10073.n309 a_71281_n10073.n308 0.496742
R53915 a_71281_n10073.n321 a_71281_n10073.n319 0.496742
R53916 a_71281_n10073.n323 a_71281_n10073.n322 0.496742
R53917 a_71281_n10073.n335 a_71281_n10073.n333 0.496742
R53918 a_71281_n10073.n337 a_71281_n10073.n336 0.496742
R53919 a_71281_n10073.n468 a_71281_n10073.n467 0.496742
R53920 a_71281_n10073.n466 a_71281_n10073.n464 0.496742
R53921 a_71281_n10073.n454 a_71281_n10073.n453 0.496742
R53922 a_71281_n10073.n452 a_71281_n10073.n450 0.496742
R53923 a_71281_n10073.n440 a_71281_n10073.n439 0.496742
R53924 a_71281_n10073.n438 a_71281_n10073.n436 0.496742
R53925 a_71281_n10073.n423 a_71281_n10073.n422 0.496742
R53926 a_71281_n10073.n421 a_71281_n10073.n419 0.496742
R53927 a_71281_n10073.n409 a_71281_n10073.n408 0.496742
R53928 a_71281_n10073.n407 a_71281_n10073.n405 0.496742
R53929 a_71281_n10073.n392 a_71281_n10073.n391 0.496742
R53930 a_71281_n10073.n390 a_71281_n10073.n388 0.496742
R53931 a_71281_n10073.n378 a_71281_n10073.n377 0.496742
R53932 a_71281_n10073.n376 a_71281_n10073.n374 0.496742
R53933 a_71281_n10073.n364 a_71281_n10073.n363 0.496742
R53934 a_71281_n10073.n362 a_71281_n10073.n360 0.496742
R53935 a_71281_n10073.n351 a_71281_n10073.n350 0.496742
R53936 a_71281_n10073.n349 a_71281_n10073.n347 0.496742
R53937 a_71281_n10073.n206 a_71281_n10073.n205 0.496742
R53938 a_71281_n10073.n204 a_71281_n10073.n202 0.496742
R53939 a_71281_n10073.n480 a_71281_n10073.n478 0.496742
R53940 a_71281_n10073.n482 a_71281_n10073.n481 0.496742
R53941 a_71281_n10073.n508 a_71281_n10073.n506 0.496742
R53942 a_71281_n10073.n510 a_71281_n10073.n509 0.496742
R53943 a_71281_n10073.n522 a_71281_n10073.n520 0.496742
R53944 a_71281_n10073.n524 a_71281_n10073.n523 0.496742
R53945 a_71281_n10073.n536 a_71281_n10073.n534 0.496742
R53946 a_71281_n10073.n538 a_71281_n10073.n537 0.496742
R53947 a_71281_n10073.n553 a_71281_n10073.n551 0.496742
R53948 a_71281_n10073.n555 a_71281_n10073.n554 0.496742
R53949 a_71281_n10073.n567 a_71281_n10073.n565 0.496742
R53950 a_71281_n10073.n569 a_71281_n10073.n568 0.496742
R53951 a_71281_n10073.n584 a_71281_n10073.n582 0.496742
R53952 a_71281_n10073.n586 a_71281_n10073.n585 0.496742
R53953 a_71281_n10073.n598 a_71281_n10073.n596 0.496742
R53954 a_71281_n10073.n600 a_71281_n10073.n599 0.496742
R53955 a_71281_n10073.n612 a_71281_n10073.n610 0.496742
R53956 a_71281_n10073.n614 a_71281_n10073.n613 0.496742
R53957 a_71281_n10073.n626 a_71281_n10073.n624 0.496742
R53958 a_71281_n10073.n628 a_71281_n10073.n627 0.496742
R53959 a_71281_n10073.n759 a_71281_n10073.n758 0.496742
R53960 a_71281_n10073.n757 a_71281_n10073.n755 0.496742
R53961 a_71281_n10073.n745 a_71281_n10073.n744 0.496742
R53962 a_71281_n10073.n743 a_71281_n10073.n741 0.496742
R53963 a_71281_n10073.n731 a_71281_n10073.n730 0.496742
R53964 a_71281_n10073.n729 a_71281_n10073.n727 0.496742
R53965 a_71281_n10073.n714 a_71281_n10073.n713 0.496742
R53966 a_71281_n10073.n712 a_71281_n10073.n710 0.496742
R53967 a_71281_n10073.n700 a_71281_n10073.n699 0.496742
R53968 a_71281_n10073.n698 a_71281_n10073.n696 0.496742
R53969 a_71281_n10073.n683 a_71281_n10073.n682 0.496742
R53970 a_71281_n10073.n681 a_71281_n10073.n679 0.496742
R53971 a_71281_n10073.n669 a_71281_n10073.n668 0.496742
R53972 a_71281_n10073.n667 a_71281_n10073.n665 0.496742
R53973 a_71281_n10073.n655 a_71281_n10073.n654 0.496742
R53974 a_71281_n10073.n653 a_71281_n10073.n651 0.496742
R53975 a_71281_n10073.n642 a_71281_n10073.n641 0.496742
R53976 a_71281_n10073.n640 a_71281_n10073.n638 0.496742
R53977 a_71281_n10073.n497 a_71281_n10073.n496 0.496742
R53978 a_71281_n10073.n495 a_71281_n10073.n493 0.496742
R53979 a_71281_n10073.n771 a_71281_n10073.n769 0.496742
R53980 a_71281_n10073.n773 a_71281_n10073.n772 0.496742
R53981 a_71281_n10073.n190 a_71281_n10073.n188 0.496742
R53982 a_71281_n10073.n192 a_71281_n10073.n191 0.496742
R53983 a_71281_n10073.n491 a_71281_n10073.n345 0.445939
R53984 a_71281_n10073.n782 a_71281_n10073.n636 0.445939
R53985 a_71281_n10073.n786 a_71281_n10073.n785 0.445939
R53986 a_71281_n10073.n491 a_71281_n10073.n490 0.443507
R53987 a_71281_n10073.n782 a_71281_n10073.n781 0.443507
R53988 a_71281_n10073.n785 a_71281_n10073.n200 0.443507
R53989 a_71281_n10073.n227 a_71281_n10073.n214 0.180804
R53990 a_71281_n10073.n303 a_71281_n10073.n290 0.180804
R53991 a_71281_n10073.n476 a_71281_n10073.n463 0.180804
R53992 a_71281_n10073.n400 a_71281_n10073.n387 0.180804
R53993 a_71281_n10073.n518 a_71281_n10073.n505 0.180804
R53994 a_71281_n10073.n594 a_71281_n10073.n581 0.180804
R53995 a_71281_n10073.n767 a_71281_n10073.n754 0.180804
R53996 a_71281_n10073.n691 a_71281_n10073.n678 0.180804
R53997 a_71281_n10073.n27 a_71281_n10073.n14 0.180804
R53998 a_71281_n10073.n841 a_71281_n10073.n828 0.180804
R53999 a_71281_n10073.n186 a_71281_n10073.n173 0.180804
R54000 a_71281_n10073.n110 a_71281_n10073.n97 0.180804
R54001 a_71281_n10073.n241 a_71281_n10073.n228 0.180196
R54002 a_71281_n10073.n272 a_71281_n10073.n259 0.180196
R54003 a_71281_n10073.n286 a_71281_n10073.n273 0.180196
R54004 a_71281_n10073.n317 a_71281_n10073.n304 0.180196
R54005 a_71281_n10073.n345 a_71281_n10073.n332 0.180196
R54006 a_71281_n10073.n490 a_71281_n10073.n477 0.180196
R54007 a_71281_n10073.n462 a_71281_n10073.n449 0.180196
R54008 a_71281_n10073.n431 a_71281_n10073.n418 0.180196
R54009 a_71281_n10073.n417 a_71281_n10073.n404 0.180196
R54010 a_71281_n10073.n386 a_71281_n10073.n373 0.180196
R54011 a_71281_n10073.n532 a_71281_n10073.n519 0.180196
R54012 a_71281_n10073.n563 a_71281_n10073.n550 0.180196
R54013 a_71281_n10073.n577 a_71281_n10073.n564 0.180196
R54014 a_71281_n10073.n608 a_71281_n10073.n595 0.180196
R54015 a_71281_n10073.n636 a_71281_n10073.n623 0.180196
R54016 a_71281_n10073.n781 a_71281_n10073.n768 0.180196
R54017 a_71281_n10073.n753 a_71281_n10073.n740 0.180196
R54018 a_71281_n10073.n722 a_71281_n10073.n709 0.180196
R54019 a_71281_n10073.n708 a_71281_n10073.n695 0.180196
R54020 a_71281_n10073.n677 a_71281_n10073.n664 0.180196
R54021 a_71281_n10073.n41 a_71281_n10073.n28 0.180196
R54022 a_71281_n10073.n872 a_71281_n10073.n859 0.180196
R54023 a_71281_n10073.n858 a_71281_n10073.n845 0.180196
R54024 a_71281_n10073.n827 a_71281_n10073.n814 0.180196
R54025 a_71281_n10073.n799 a_71281_n10073.n786 0.180196
R54026 a_71281_n10073.n200 a_71281_n10073.n187 0.180196
R54027 a_71281_n10073.n172 a_71281_n10073.n159 0.180196
R54028 a_71281_n10073.n141 a_71281_n10073.n128 0.180196
R54029 a_71281_n10073.n127 a_71281_n10073.n114 0.180196
R54030 a_71281_n10073.n96 a_71281_n10073.n83 0.180196
R54031 a_71281_n10073.n255 a_71281_n10073.n242 0.179892
R54032 a_71281_n10073.n331 a_71281_n10073.n318 0.179892
R54033 a_71281_n10073.n448 a_71281_n10073.n435 0.179892
R54034 a_71281_n10073.n372 a_71281_n10073.n359 0.179892
R54035 a_71281_n10073.n546 a_71281_n10073.n533 0.179892
R54036 a_71281_n10073.n622 a_71281_n10073.n609 0.179892
R54037 a_71281_n10073.n739 a_71281_n10073.n726 0.179892
R54038 a_71281_n10073.n663 a_71281_n10073.n650 0.179892
R54039 a_71281_n10073.n55 a_71281_n10073.n42 0.179892
R54040 a_71281_n10073.n813 a_71281_n10073.n800 0.179892
R54041 a_71281_n10073.n158 a_71281_n10073.n145 0.179892
R54042 a_71281_n10073.n82 a_71281_n10073.n69 0.179892
R54043 a_71281_n10073.n26 a_71281_n10073.n15 0.136625
R54044 a_71281_n10073.n20 a_71281_n10073.n19 0.136625
R54045 a_71281_n10073.n40 a_71281_n10073.n29 0.136625
R54046 a_71281_n10073.n34 a_71281_n10073.n33 0.136625
R54047 a_71281_n10073.n54 a_71281_n10073.n43 0.136625
R54048 a_71281_n10073.n48 a_71281_n10073.n47 0.136625
R54049 a_71281_n10073.n866 a_71281_n10073.n864 0.136625
R54050 a_71281_n10073.n871 a_71281_n10073.n860 0.136625
R54051 a_71281_n10073.n852 a_71281_n10073.n850 0.136625
R54052 a_71281_n10073.n857 a_71281_n10073.n846 0.136625
R54053 a_71281_n10073.n835 a_71281_n10073.n833 0.136625
R54054 a_71281_n10073.n840 a_71281_n10073.n829 0.136625
R54055 a_71281_n10073.n821 a_71281_n10073.n819 0.136625
R54056 a_71281_n10073.n826 a_71281_n10073.n815 0.136625
R54057 a_71281_n10073.n807 a_71281_n10073.n805 0.136625
R54058 a_71281_n10073.n812 a_71281_n10073.n801 0.136625
R54059 a_71281_n10073.n793 a_71281_n10073.n791 0.136625
R54060 a_71281_n10073.n798 a_71281_n10073.n787 0.136625
R54061 a_71281_n10073.n180 a_71281_n10073.n178 0.136625
R54062 a_71281_n10073.n185 a_71281_n10073.n174 0.136625
R54063 a_71281_n10073.n166 a_71281_n10073.n164 0.136625
R54064 a_71281_n10073.n171 a_71281_n10073.n160 0.136625
R54065 a_71281_n10073.n152 a_71281_n10073.n150 0.136625
R54066 a_71281_n10073.n157 a_71281_n10073.n146 0.136625
R54067 a_71281_n10073.n135 a_71281_n10073.n133 0.136625
R54068 a_71281_n10073.n140 a_71281_n10073.n129 0.136625
R54069 a_71281_n10073.n121 a_71281_n10073.n119 0.136625
R54070 a_71281_n10073.n126 a_71281_n10073.n115 0.136625
R54071 a_71281_n10073.n104 a_71281_n10073.n102 0.136625
R54072 a_71281_n10073.n109 a_71281_n10073.n98 0.136625
R54073 a_71281_n10073.n90 a_71281_n10073.n88 0.136625
R54074 a_71281_n10073.n95 a_71281_n10073.n84 0.136625
R54075 a_71281_n10073.n76 a_71281_n10073.n74 0.136625
R54076 a_71281_n10073.n81 a_71281_n10073.n70 0.136625
R54077 a_71281_n10073.n61 a_71281_n10073.n56 0.136625
R54078 a_71281_n10073.n67 a_71281_n10073.n57 0.136625
R54079 a_71281_n10073.n6 a_71281_n10073.n1 0.136625
R54080 a_71281_n10073.n12 a_71281_n10073.n2 0.136625
R54081 a_71281_n10073.n226 a_71281_n10073.n215 0.136625
R54082 a_71281_n10073.n220 a_71281_n10073.n219 0.136625
R54083 a_71281_n10073.n240 a_71281_n10073.n229 0.136625
R54084 a_71281_n10073.n234 a_71281_n10073.n233 0.136625
R54085 a_71281_n10073.n254 a_71281_n10073.n243 0.136625
R54086 a_71281_n10073.n248 a_71281_n10073.n247 0.136625
R54087 a_71281_n10073.n271 a_71281_n10073.n260 0.136625
R54088 a_71281_n10073.n265 a_71281_n10073.n264 0.136625
R54089 a_71281_n10073.n285 a_71281_n10073.n274 0.136625
R54090 a_71281_n10073.n279 a_71281_n10073.n278 0.136625
R54091 a_71281_n10073.n302 a_71281_n10073.n291 0.136625
R54092 a_71281_n10073.n296 a_71281_n10073.n295 0.136625
R54093 a_71281_n10073.n316 a_71281_n10073.n305 0.136625
R54094 a_71281_n10073.n310 a_71281_n10073.n309 0.136625
R54095 a_71281_n10073.n330 a_71281_n10073.n319 0.136625
R54096 a_71281_n10073.n324 a_71281_n10073.n323 0.136625
R54097 a_71281_n10073.n344 a_71281_n10073.n333 0.136625
R54098 a_71281_n10073.n338 a_71281_n10073.n337 0.136625
R54099 a_71281_n10073.n470 a_71281_n10073.n468 0.136625
R54100 a_71281_n10073.n475 a_71281_n10073.n464 0.136625
R54101 a_71281_n10073.n456 a_71281_n10073.n454 0.136625
R54102 a_71281_n10073.n461 a_71281_n10073.n450 0.136625
R54103 a_71281_n10073.n442 a_71281_n10073.n440 0.136625
R54104 a_71281_n10073.n447 a_71281_n10073.n436 0.136625
R54105 a_71281_n10073.n425 a_71281_n10073.n423 0.136625
R54106 a_71281_n10073.n430 a_71281_n10073.n419 0.136625
R54107 a_71281_n10073.n411 a_71281_n10073.n409 0.136625
R54108 a_71281_n10073.n416 a_71281_n10073.n405 0.136625
R54109 a_71281_n10073.n394 a_71281_n10073.n392 0.136625
R54110 a_71281_n10073.n399 a_71281_n10073.n388 0.136625
R54111 a_71281_n10073.n380 a_71281_n10073.n378 0.136625
R54112 a_71281_n10073.n385 a_71281_n10073.n374 0.136625
R54113 a_71281_n10073.n366 a_71281_n10073.n364 0.136625
R54114 a_71281_n10073.n371 a_71281_n10073.n360 0.136625
R54115 a_71281_n10073.n351 a_71281_n10073.n346 0.136625
R54116 a_71281_n10073.n357 a_71281_n10073.n347 0.136625
R54117 a_71281_n10073.n206 a_71281_n10073.n201 0.136625
R54118 a_71281_n10073.n212 a_71281_n10073.n202 0.136625
R54119 a_71281_n10073.n489 a_71281_n10073.n478 0.136625
R54120 a_71281_n10073.n483 a_71281_n10073.n482 0.136625
R54121 a_71281_n10073.n517 a_71281_n10073.n506 0.136625
R54122 a_71281_n10073.n511 a_71281_n10073.n510 0.136625
R54123 a_71281_n10073.n531 a_71281_n10073.n520 0.136625
R54124 a_71281_n10073.n525 a_71281_n10073.n524 0.136625
R54125 a_71281_n10073.n545 a_71281_n10073.n534 0.136625
R54126 a_71281_n10073.n539 a_71281_n10073.n538 0.136625
R54127 a_71281_n10073.n562 a_71281_n10073.n551 0.136625
R54128 a_71281_n10073.n556 a_71281_n10073.n555 0.136625
R54129 a_71281_n10073.n576 a_71281_n10073.n565 0.136625
R54130 a_71281_n10073.n570 a_71281_n10073.n569 0.136625
R54131 a_71281_n10073.n593 a_71281_n10073.n582 0.136625
R54132 a_71281_n10073.n587 a_71281_n10073.n586 0.136625
R54133 a_71281_n10073.n607 a_71281_n10073.n596 0.136625
R54134 a_71281_n10073.n601 a_71281_n10073.n600 0.136625
R54135 a_71281_n10073.n621 a_71281_n10073.n610 0.136625
R54136 a_71281_n10073.n615 a_71281_n10073.n614 0.136625
R54137 a_71281_n10073.n635 a_71281_n10073.n624 0.136625
R54138 a_71281_n10073.n629 a_71281_n10073.n628 0.136625
R54139 a_71281_n10073.n761 a_71281_n10073.n759 0.136625
R54140 a_71281_n10073.n766 a_71281_n10073.n755 0.136625
R54141 a_71281_n10073.n747 a_71281_n10073.n745 0.136625
R54142 a_71281_n10073.n752 a_71281_n10073.n741 0.136625
R54143 a_71281_n10073.n733 a_71281_n10073.n731 0.136625
R54144 a_71281_n10073.n738 a_71281_n10073.n727 0.136625
R54145 a_71281_n10073.n716 a_71281_n10073.n714 0.136625
R54146 a_71281_n10073.n721 a_71281_n10073.n710 0.136625
R54147 a_71281_n10073.n702 a_71281_n10073.n700 0.136625
R54148 a_71281_n10073.n707 a_71281_n10073.n696 0.136625
R54149 a_71281_n10073.n685 a_71281_n10073.n683 0.136625
R54150 a_71281_n10073.n690 a_71281_n10073.n679 0.136625
R54151 a_71281_n10073.n671 a_71281_n10073.n669 0.136625
R54152 a_71281_n10073.n676 a_71281_n10073.n665 0.136625
R54153 a_71281_n10073.n657 a_71281_n10073.n655 0.136625
R54154 a_71281_n10073.n662 a_71281_n10073.n651 0.136625
R54155 a_71281_n10073.n642 a_71281_n10073.n637 0.136625
R54156 a_71281_n10073.n648 a_71281_n10073.n638 0.136625
R54157 a_71281_n10073.n497 a_71281_n10073.n492 0.136625
R54158 a_71281_n10073.n503 a_71281_n10073.n493 0.136625
R54159 a_71281_n10073.n780 a_71281_n10073.n769 0.136625
R54160 a_71281_n10073.n774 a_71281_n10073.n773 0.136625
R54161 a_71281_n10073.n199 a_71281_n10073.n188 0.136625
R54162 a_71281_n10073.n193 a_71281_n10073.n192 0.136625
R54163 a_71281_n10073.n214 a_71281_n10073.n213 0.095973
R54164 a_71281_n10073.n228 a_71281_n10073.n227 0.095973
R54165 a_71281_n10073.n242 a_71281_n10073.n241 0.095973
R54166 a_71281_n10073.n273 a_71281_n10073.n272 0.095973
R54167 a_71281_n10073.n304 a_71281_n10073.n303 0.095973
R54168 a_71281_n10073.n318 a_71281_n10073.n317 0.095973
R54169 a_71281_n10073.n332 a_71281_n10073.n331 0.095973
R54170 a_71281_n10073.n477 a_71281_n10073.n476 0.095973
R54171 a_71281_n10073.n463 a_71281_n10073.n462 0.095973
R54172 a_71281_n10073.n449 a_71281_n10073.n448 0.095973
R54173 a_71281_n10073.n418 a_71281_n10073.n417 0.095973
R54174 a_71281_n10073.n387 a_71281_n10073.n386 0.095973
R54175 a_71281_n10073.n373 a_71281_n10073.n372 0.095973
R54176 a_71281_n10073.n359 a_71281_n10073.n358 0.095973
R54177 a_71281_n10073.n505 a_71281_n10073.n504 0.095973
R54178 a_71281_n10073.n519 a_71281_n10073.n518 0.095973
R54179 a_71281_n10073.n533 a_71281_n10073.n532 0.095973
R54180 a_71281_n10073.n564 a_71281_n10073.n563 0.095973
R54181 a_71281_n10073.n595 a_71281_n10073.n594 0.095973
R54182 a_71281_n10073.n609 a_71281_n10073.n608 0.095973
R54183 a_71281_n10073.n623 a_71281_n10073.n622 0.095973
R54184 a_71281_n10073.n768 a_71281_n10073.n767 0.095973
R54185 a_71281_n10073.n754 a_71281_n10073.n753 0.095973
R54186 a_71281_n10073.n740 a_71281_n10073.n739 0.095973
R54187 a_71281_n10073.n709 a_71281_n10073.n708 0.095973
R54188 a_71281_n10073.n678 a_71281_n10073.n677 0.095973
R54189 a_71281_n10073.n664 a_71281_n10073.n663 0.095973
R54190 a_71281_n10073.n650 a_71281_n10073.n649 0.095973
R54191 a_71281_n10073.n14 a_71281_n10073.n13 0.095973
R54192 a_71281_n10073.n28 a_71281_n10073.n27 0.095973
R54193 a_71281_n10073.n42 a_71281_n10073.n41 0.095973
R54194 a_71281_n10073.n859 a_71281_n10073.n858 0.095973
R54195 a_71281_n10073.n828 a_71281_n10073.n827 0.095973
R54196 a_71281_n10073.n814 a_71281_n10073.n813 0.095973
R54197 a_71281_n10073.n800 a_71281_n10073.n799 0.095973
R54198 a_71281_n10073.n187 a_71281_n10073.n186 0.095973
R54199 a_71281_n10073.n173 a_71281_n10073.n172 0.095973
R54200 a_71281_n10073.n159 a_71281_n10073.n158 0.095973
R54201 a_71281_n10073.n128 a_71281_n10073.n127 0.095973
R54202 a_71281_n10073.n97 a_71281_n10073.n96 0.095973
R54203 a_71281_n10073.n83 a_71281_n10073.n82 0.095973
R54204 a_71281_n10073.n69 a_71281_n10073.n68 0.095973
R54205 a_71281_n10073.n26 a_71281_n10073.n25 0.0719743
R54206 a_71281_n10073.n22 a_71281_n10073.n20 0.0719743
R54207 a_71281_n10073.n40 a_71281_n10073.n39 0.0719743
R54208 a_71281_n10073.n36 a_71281_n10073.n34 0.0719743
R54209 a_71281_n10073.n54 a_71281_n10073.n53 0.0719743
R54210 a_71281_n10073.n50 a_71281_n10073.n48 0.0719743
R54211 a_71281_n10073.n867 a_71281_n10073.n866 0.0719743
R54212 a_71281_n10073.n871 a_71281_n10073.n870 0.0719743
R54213 a_71281_n10073.n853 a_71281_n10073.n852 0.0719743
R54214 a_71281_n10073.n857 a_71281_n10073.n856 0.0719743
R54215 a_71281_n10073.n836 a_71281_n10073.n835 0.0719743
R54216 a_71281_n10073.n840 a_71281_n10073.n839 0.0719743
R54217 a_71281_n10073.n822 a_71281_n10073.n821 0.0719743
R54218 a_71281_n10073.n826 a_71281_n10073.n825 0.0719743
R54219 a_71281_n10073.n808 a_71281_n10073.n807 0.0719743
R54220 a_71281_n10073.n812 a_71281_n10073.n811 0.0719743
R54221 a_71281_n10073.n794 a_71281_n10073.n793 0.0719743
R54222 a_71281_n10073.n798 a_71281_n10073.n797 0.0719743
R54223 a_71281_n10073.n181 a_71281_n10073.n180 0.0719743
R54224 a_71281_n10073.n185 a_71281_n10073.n184 0.0719743
R54225 a_71281_n10073.n167 a_71281_n10073.n166 0.0719743
R54226 a_71281_n10073.n171 a_71281_n10073.n170 0.0719743
R54227 a_71281_n10073.n153 a_71281_n10073.n152 0.0719743
R54228 a_71281_n10073.n157 a_71281_n10073.n156 0.0719743
R54229 a_71281_n10073.n136 a_71281_n10073.n135 0.0719743
R54230 a_71281_n10073.n140 a_71281_n10073.n139 0.0719743
R54231 a_71281_n10073.n122 a_71281_n10073.n121 0.0719743
R54232 a_71281_n10073.n126 a_71281_n10073.n125 0.0719743
R54233 a_71281_n10073.n105 a_71281_n10073.n104 0.0719743
R54234 a_71281_n10073.n109 a_71281_n10073.n108 0.0719743
R54235 a_71281_n10073.n91 a_71281_n10073.n90 0.0719743
R54236 a_71281_n10073.n95 a_71281_n10073.n94 0.0719743
R54237 a_71281_n10073.n77 a_71281_n10073.n76 0.0719743
R54238 a_71281_n10073.n81 a_71281_n10073.n80 0.0719743
R54239 a_71281_n10073.n63 a_71281_n10073.n56 0.0719743
R54240 a_71281_n10073.n67 a_71281_n10073.n66 0.0719743
R54241 a_71281_n10073.n8 a_71281_n10073.n1 0.0719743
R54242 a_71281_n10073.n12 a_71281_n10073.n11 0.0719743
R54243 a_71281_n10073.n226 a_71281_n10073.n225 0.0719743
R54244 a_71281_n10073.n222 a_71281_n10073.n220 0.0719743
R54245 a_71281_n10073.n240 a_71281_n10073.n239 0.0719743
R54246 a_71281_n10073.n236 a_71281_n10073.n234 0.0719743
R54247 a_71281_n10073.n254 a_71281_n10073.n253 0.0719743
R54248 a_71281_n10073.n250 a_71281_n10073.n248 0.0719743
R54249 a_71281_n10073.n271 a_71281_n10073.n270 0.0719743
R54250 a_71281_n10073.n267 a_71281_n10073.n265 0.0719743
R54251 a_71281_n10073.n285 a_71281_n10073.n284 0.0719743
R54252 a_71281_n10073.n281 a_71281_n10073.n279 0.0719743
R54253 a_71281_n10073.n302 a_71281_n10073.n301 0.0719743
R54254 a_71281_n10073.n298 a_71281_n10073.n296 0.0719743
R54255 a_71281_n10073.n316 a_71281_n10073.n315 0.0719743
R54256 a_71281_n10073.n312 a_71281_n10073.n310 0.0719743
R54257 a_71281_n10073.n330 a_71281_n10073.n329 0.0719743
R54258 a_71281_n10073.n326 a_71281_n10073.n324 0.0719743
R54259 a_71281_n10073.n344 a_71281_n10073.n343 0.0719743
R54260 a_71281_n10073.n340 a_71281_n10073.n338 0.0719743
R54261 a_71281_n10073.n471 a_71281_n10073.n470 0.0719743
R54262 a_71281_n10073.n475 a_71281_n10073.n474 0.0719743
R54263 a_71281_n10073.n457 a_71281_n10073.n456 0.0719743
R54264 a_71281_n10073.n461 a_71281_n10073.n460 0.0719743
R54265 a_71281_n10073.n443 a_71281_n10073.n442 0.0719743
R54266 a_71281_n10073.n447 a_71281_n10073.n446 0.0719743
R54267 a_71281_n10073.n426 a_71281_n10073.n425 0.0719743
R54268 a_71281_n10073.n430 a_71281_n10073.n429 0.0719743
R54269 a_71281_n10073.n412 a_71281_n10073.n411 0.0719743
R54270 a_71281_n10073.n416 a_71281_n10073.n415 0.0719743
R54271 a_71281_n10073.n395 a_71281_n10073.n394 0.0719743
R54272 a_71281_n10073.n399 a_71281_n10073.n398 0.0719743
R54273 a_71281_n10073.n381 a_71281_n10073.n380 0.0719743
R54274 a_71281_n10073.n385 a_71281_n10073.n384 0.0719743
R54275 a_71281_n10073.n367 a_71281_n10073.n366 0.0719743
R54276 a_71281_n10073.n371 a_71281_n10073.n370 0.0719743
R54277 a_71281_n10073.n353 a_71281_n10073.n346 0.0719743
R54278 a_71281_n10073.n357 a_71281_n10073.n356 0.0719743
R54279 a_71281_n10073.n208 a_71281_n10073.n201 0.0719743
R54280 a_71281_n10073.n212 a_71281_n10073.n211 0.0719743
R54281 a_71281_n10073.n489 a_71281_n10073.n488 0.0719743
R54282 a_71281_n10073.n485 a_71281_n10073.n483 0.0719743
R54283 a_71281_n10073.n517 a_71281_n10073.n516 0.0719743
R54284 a_71281_n10073.n513 a_71281_n10073.n511 0.0719743
R54285 a_71281_n10073.n531 a_71281_n10073.n530 0.0719743
R54286 a_71281_n10073.n527 a_71281_n10073.n525 0.0719743
R54287 a_71281_n10073.n545 a_71281_n10073.n544 0.0719743
R54288 a_71281_n10073.n541 a_71281_n10073.n539 0.0719743
R54289 a_71281_n10073.n562 a_71281_n10073.n561 0.0719743
R54290 a_71281_n10073.n558 a_71281_n10073.n556 0.0719743
R54291 a_71281_n10073.n576 a_71281_n10073.n575 0.0719743
R54292 a_71281_n10073.n572 a_71281_n10073.n570 0.0719743
R54293 a_71281_n10073.n593 a_71281_n10073.n592 0.0719743
R54294 a_71281_n10073.n589 a_71281_n10073.n587 0.0719743
R54295 a_71281_n10073.n607 a_71281_n10073.n606 0.0719743
R54296 a_71281_n10073.n603 a_71281_n10073.n601 0.0719743
R54297 a_71281_n10073.n621 a_71281_n10073.n620 0.0719743
R54298 a_71281_n10073.n617 a_71281_n10073.n615 0.0719743
R54299 a_71281_n10073.n635 a_71281_n10073.n634 0.0719743
R54300 a_71281_n10073.n631 a_71281_n10073.n629 0.0719743
R54301 a_71281_n10073.n762 a_71281_n10073.n761 0.0719743
R54302 a_71281_n10073.n766 a_71281_n10073.n765 0.0719743
R54303 a_71281_n10073.n748 a_71281_n10073.n747 0.0719743
R54304 a_71281_n10073.n752 a_71281_n10073.n751 0.0719743
R54305 a_71281_n10073.n734 a_71281_n10073.n733 0.0719743
R54306 a_71281_n10073.n738 a_71281_n10073.n737 0.0719743
R54307 a_71281_n10073.n717 a_71281_n10073.n716 0.0719743
R54308 a_71281_n10073.n721 a_71281_n10073.n720 0.0719743
R54309 a_71281_n10073.n703 a_71281_n10073.n702 0.0719743
R54310 a_71281_n10073.n707 a_71281_n10073.n706 0.0719743
R54311 a_71281_n10073.n686 a_71281_n10073.n685 0.0719743
R54312 a_71281_n10073.n690 a_71281_n10073.n689 0.0719743
R54313 a_71281_n10073.n672 a_71281_n10073.n671 0.0719743
R54314 a_71281_n10073.n676 a_71281_n10073.n675 0.0719743
R54315 a_71281_n10073.n658 a_71281_n10073.n657 0.0719743
R54316 a_71281_n10073.n662 a_71281_n10073.n661 0.0719743
R54317 a_71281_n10073.n644 a_71281_n10073.n637 0.0719743
R54318 a_71281_n10073.n648 a_71281_n10073.n647 0.0719743
R54319 a_71281_n10073.n499 a_71281_n10073.n492 0.0719743
R54320 a_71281_n10073.n503 a_71281_n10073.n502 0.0719743
R54321 a_71281_n10073.n780 a_71281_n10073.n779 0.0719743
R54322 a_71281_n10073.n776 a_71281_n10073.n774 0.0719743
R54323 a_71281_n10073.n199 a_71281_n10073.n198 0.0719743
R54324 a_71281_n10073.n195 a_71281_n10073.n193 0.0719743
R54325 a_71281_n10073.n289 a_71281_n10073.n286 0.0485405
R54326 a_71281_n10073.n404 a_71281_n10073.n403 0.0485405
R54327 a_71281_n10073.n580 a_71281_n10073.n577 0.0485405
R54328 a_71281_n10073.n695 a_71281_n10073.n694 0.0485405
R54329 a_71281_n10073.n845 a_71281_n10073.n844 0.0485405
R54330 a_71281_n10073.n114 a_71281_n10073.n113 0.0485405
R54331 a_71281_n10073.n258 a_71281_n10073.n255 0.0482365
R54332 a_71281_n10073.n259 a_71281_n10073.n258 0.0482365
R54333 a_71281_n10073.n435 a_71281_n10073.n434 0.0482365
R54334 a_71281_n10073.n434 a_71281_n10073.n431 0.0482365
R54335 a_71281_n10073.n549 a_71281_n10073.n546 0.0482365
R54336 a_71281_n10073.n550 a_71281_n10073.n549 0.0482365
R54337 a_71281_n10073.n726 a_71281_n10073.n725 0.0482365
R54338 a_71281_n10073.n725 a_71281_n10073.n722 0.0482365
R54339 a_71281_n10073.n873 a_71281_n10073.n55 0.0482365
R54340 a_71281_n10073.n873 a_71281_n10073.n872 0.0482365
R54341 a_71281_n10073.n145 a_71281_n10073.n144 0.0482365
R54342 a_71281_n10073.n144 a_71281_n10073.n141 0.0482365
R54343 a_71281_n10073.n290 a_71281_n10073.n289 0.0479324
R54344 a_71281_n10073.n403 a_71281_n10073.n400 0.0479324
R54345 a_71281_n10073.n581 a_71281_n10073.n580 0.0479324
R54346 a_71281_n10073.n694 a_71281_n10073.n691 0.0479324
R54347 a_71281_n10073.n844 a_71281_n10073.n841 0.0479324
R54348 a_71281_n10073.n113 a_71281_n10073.n110 0.0479324
R54349 a_71281_n10073.t72 a_71281_n10073.n0 3.76597
R54350 a_60677_10448.t0 a_60677_10448.t2 60.9362
R54351 a_60677_10448.t2 a_60677_10448.t5 12.9273
R54352 a_60677_10448.t2 a_60677_10448.t1 10.1307
R54353 a_60677_10448.t2 a_60677_10448.t4 8.54643
R54354 a_60677_10448.t2 a_60677_10448.t3 7.50895
R54355 a_33379_34007.t2 a_33379_34007.n351 10.937
R54356 a_33379_34007.t27 a_33379_34007.n350 9.74618
R54357 a_33379_34007.n351 a_33379_34007.t3 9.33982
R54358 a_33379_34007.n180 a_33379_34007.t8 8.38704
R54359 a_33379_34007.n305 a_33379_34007.t20 8.38704
R54360 a_33379_34007.n139 a_33379_34007.t33 8.37857
R54361 a_33379_34007.n286 a_33379_34007.t36 8.37857
R54362 a_33379_34007.n55 a_33379_34007.t40 8.39293
R54363 a_33379_34007.n83 a_33379_34007.t50 8.39293
R54364 a_33379_34007.n37 a_33379_34007.t45 8.10567
R54365 a_33379_34007.n133 a_33379_34007.t19 8.10567
R54366 a_33379_34007.n6 a_33379_34007.t78 8.10567
R54367 a_33379_34007.n25 a_33379_34007.t48 8.10567
R54368 a_33379_34007.n148 a_33379_34007.t39 8.10567
R54369 a_33379_34007.n149 a_33379_34007.t91 8.10567
R54370 a_33379_34007.n150 a_33379_34007.t63 8.10567
R54371 a_33379_34007.n138 a_33379_34007.t13 8.10567
R54372 a_33379_34007.n3 a_33379_34007.t73 8.10567
R54373 a_33379_34007.n23 a_33379_34007.t12 8.10567
R54374 a_33379_34007.n42 a_33379_34007.t74 8.10567
R54375 a_33379_34007.n120 a_33379_34007.t47 8.10567
R54376 a_33379_34007.n12 a_33379_34007.t21 8.10567
R54377 a_33379_34007.n128 a_33379_34007.t61 8.10567
R54378 a_33379_34007.n127 a_33379_34007.t11 8.10567
R54379 a_33379_34007.n126 a_33379_34007.t72 8.10567
R54380 a_33379_34007.n38 a_33379_34007.t38 8.10567
R54381 a_33379_34007.n130 a_33379_34007.t10 8.10567
R54382 a_33379_34007.n9 a_33379_34007.t80 8.10567
R54383 a_33379_34007.n29 a_33379_34007.t41 8.10567
R54384 a_33379_34007.n60 a_33379_34007.t56 8.10567
R54385 a_33379_34007.n58 a_33379_34007.t28 8.10567
R54386 a_33379_34007.n56 a_33379_34007.t85 8.10567
R54387 a_33379_34007.n222 a_33379_34007.t60 8.10567
R54388 a_33379_34007.n207 a_33379_34007.t34 8.10567
R54389 a_33379_34007.n208 a_33379_34007.t86 8.10567
R54390 a_33379_34007.n209 a_33379_34007.t58 8.10567
R54391 a_33379_34007.n54 a_33379_34007.t26 8.10567
R54392 a_33379_34007.n53 a_33379_34007.t82 8.10567
R54393 a_33379_34007.n51 a_33379_34007.t25 8.10567
R54394 a_33379_34007.n75 a_33379_34007.t84 8.10567
R54395 a_33379_34007.n72 a_33379_34007.t57 8.10567
R54396 a_33379_34007.n179 a_33379_34007.t29 8.10567
R54397 a_33379_34007.n189 a_33379_34007.t55 8.10567
R54398 a_33379_34007.n188 a_33379_34007.t4 8.10567
R54399 a_33379_34007.n187 a_33379_34007.t67 8.10567
R54400 a_33379_34007.n68 a_33379_34007.t49 8.10567
R54401 a_33379_34007.n67 a_33379_34007.t22 8.10567
R54402 a_33379_34007.n66 a_33379_34007.t88 8.10567
R54403 a_33379_34007.n63 a_33379_34007.t53 8.10567
R54404 a_33379_34007.n45 a_33379_34007.t51 8.10567
R54405 a_33379_34007.n275 a_33379_34007.t23 8.10567
R54406 a_33379_34007.n18 a_33379_34007.t81 8.10567
R54407 a_33379_34007.n33 a_33379_34007.t54 8.10567
R54408 a_33379_34007.n283 a_33379_34007.t44 8.10567
R54409 a_33379_34007.n282 a_33379_34007.t7 8.10567
R54410 a_33379_34007.n281 a_33379_34007.t70 8.10567
R54411 a_33379_34007.n285 a_33379_34007.t18 8.10567
R54412 a_33379_34007.n15 a_33379_34007.t77 8.10567
R54413 a_33379_34007.n32 a_33379_34007.t17 8.10567
R54414 a_33379_34007.n50 a_33379_34007.t79 8.10567
R54415 a_33379_34007.n243 a_33379_34007.t52 8.10567
R54416 a_33379_34007.n20 a_33379_34007.t24 8.10567
R54417 a_33379_34007.n254 a_33379_34007.t66 8.10567
R54418 a_33379_34007.n253 a_33379_34007.t16 8.10567
R54419 a_33379_34007.n252 a_33379_34007.t76 8.10567
R54420 a_33379_34007.n47 a_33379_34007.t42 8.10567
R54421 a_33379_34007.n264 a_33379_34007.t14 8.10567
R54422 a_33379_34007.n19 a_33379_34007.t83 8.10567
R54423 a_33379_34007.n36 a_33379_34007.t46 8.10567
R54424 a_33379_34007.n92 a_33379_34007.t65 8.10567
R54425 a_33379_34007.n89 a_33379_34007.t35 8.10567
R54426 a_33379_34007.n86 a_33379_34007.t5 8.10567
R54427 a_33379_34007.n298 a_33379_34007.t71 8.10567
R54428 a_33379_34007.n339 a_33379_34007.t43 8.10567
R54429 a_33379_34007.n338 a_33379_34007.t6 8.10567
R54430 a_33379_34007.n337 a_33379_34007.t69 8.10567
R54431 a_33379_34007.n82 a_33379_34007.t32 8.10567
R54432 a_33379_34007.n81 a_33379_34007.t89 8.10567
R54433 a_33379_34007.n78 a_33379_34007.t31 8.10567
R54434 a_33379_34007.n106 a_33379_34007.t92 8.10567
R54435 a_33379_34007.n104 a_33379_34007.t68 8.10567
R54436 a_33379_34007.n304 a_33379_34007.t37 8.10567
R54437 a_33379_34007.n317 a_33379_34007.t64 8.10567
R54438 a_33379_34007.n316 a_33379_34007.t15 8.10567
R54439 a_33379_34007.n315 a_33379_34007.t75 8.10567
R54440 a_33379_34007.n101 a_33379_34007.t59 8.10567
R54441 a_33379_34007.n99 a_33379_34007.t30 8.10567
R54442 a_33379_34007.n96 a_33379_34007.t9 8.10567
R54443 a_33379_34007.n94 a_33379_34007.t62 8.10567
R54444 a_33379_34007.n350 a_33379_34007.n349 6.72496
R54445 a_33379_34007.n69 a_33379_34007.n68 2.25163
R54446 a_33379_34007.n102 a_33379_34007.n101 2.25163
R54447 a_33379_34007.n39 a_33379_34007.n38 2.24588
R54448 a_33379_34007.n48 a_33379_34007.n47 2.24588
R54449 a_33379_34007.n26 a_33379_34007.n25 2.2453
R54450 a_33379_34007.n34 a_33379_34007.n33 2.2453
R54451 a_33379_34007.n117 a_33379_34007.n11 4.5005
R54452 a_33379_34007.n119 a_33379_34007.n118 4.5005
R54453 a_33379_34007.n121 a_33379_34007.n116 4.5005
R54454 a_33379_34007.n123 a_33379_34007.n122 4.5005
R54455 a_33379_34007.n124 a_33379_34007.n41 4.5005
R54456 a_33379_34007.n42 a_33379_34007.n40 4.5005
R54457 a_33379_34007.n125 a_33379_34007.n115 4.5005
R54458 a_33379_34007.n175 a_33379_34007.n174 4.5005
R54459 a_33379_34007.n29 a_33379_34007.n27 4.5005
R54460 a_33379_34007.n28 a_33379_34007.n173 4.5005
R54461 a_33379_34007.n172 a_33379_34007.n8 4.5005
R54462 a_33379_34007.n171 a_33379_34007.n9 4.5005
R54463 a_33379_34007.n7 a_33379_34007.n129 4.5005
R54464 a_33379_34007.n170 a_33379_34007.n169 4.5005
R54465 a_33379_34007.n168 a_33379_34007.n167 4.5005
R54466 a_33379_34007.n166 a_33379_34007.n131 4.5005
R54467 a_33379_34007.n165 a_33379_34007.n164 4.5005
R54468 a_33379_34007.n24 a_33379_34007.n163 4.5005
R54469 a_33379_34007.n162 a_33379_34007.n5 4.5005
R54470 a_33379_34007.n161 a_33379_34007.n6 4.5005
R54471 a_33379_34007.n4 a_33379_34007.n132 4.5005
R54472 a_33379_34007.n160 a_33379_34007.n159 4.5005
R54473 a_33379_34007.n158 a_33379_34007.n157 4.5005
R54474 a_33379_34007.n156 a_33379_34007.n134 4.5005
R54475 a_33379_34007.n155 a_33379_34007.n154 4.5005
R54476 a_33379_34007.n153 a_33379_34007.n37 4.5005
R54477 a_33379_34007.n152 a_33379_34007.n151 4.5005
R54478 a_33379_34007.n147 a_33379_34007.n146 4.5005
R54479 a_33379_34007.n145 a_33379_34007.n23 4.5005
R54480 a_33379_34007.n22 a_33379_34007.n136 4.5005
R54481 a_33379_34007.n144 a_33379_34007.n143 4.5005
R54482 a_33379_34007.n142 a_33379_34007.n3 4.5005
R54483 a_33379_34007.n2 a_33379_34007.n137 4.5005
R54484 a_33379_34007.n141 a_33379_34007.n140 4.5005
R54485 a_33379_34007.n186 a_33379_34007.n177 4.5005
R54486 a_33379_34007.n75 a_33379_34007.n73 4.5005
R54487 a_33379_34007.n185 a_33379_34007.n74 4.5005
R54488 a_33379_34007.n184 a_33379_34007.n183 4.5005
R54489 a_33379_34007.n72 a_33379_34007.n70 4.5005
R54490 a_33379_34007.n71 a_33379_34007.n182 4.5005
R54491 a_33379_34007.n181 a_33379_34007.n178 4.5005
R54492 a_33379_34007.n234 a_33379_34007.n233 4.5005
R54493 a_33379_34007.n63 a_33379_34007.n61 4.5005
R54494 a_33379_34007.n62 a_33379_34007.n232 4.5005
R54495 a_33379_34007.n231 a_33379_34007.n64 4.5005
R54496 a_33379_34007.n230 a_33379_34007.n66 4.5005
R54497 a_33379_34007.n65 a_33379_34007.n190 4.5005
R54498 a_33379_34007.n229 a_33379_34007.n228 4.5005
R54499 a_33379_34007.n227 a_33379_34007.n67 4.5005
R54500 a_33379_34007.n226 a_33379_34007.n225 4.5005
R54501 a_33379_34007.n224 a_33379_34007.n191 4.5005
R54502 a_33379_34007.n211 a_33379_34007.n210 4.5005
R54503 a_33379_34007.n60 a_33379_34007.n59 4.5005
R54504 a_33379_34007.n212 a_33379_34007.n194 4.5005
R54505 a_33379_34007.n214 a_33379_34007.n213 4.5005
R54506 a_33379_34007.n58 a_33379_34007.n57 4.5005
R54507 a_33379_34007.n215 a_33379_34007.n193 4.5005
R54508 a_33379_34007.n217 a_33379_34007.n216 4.5005
R54509 a_33379_34007.n218 a_33379_34007.n56 4.5005
R54510 a_33379_34007.n220 a_33379_34007.n219 4.5005
R54511 a_33379_34007.n221 a_33379_34007.n192 4.5005
R54512 a_33379_34007.n206 a_33379_34007.n205 4.5005
R54513 a_33379_34007.n204 a_33379_34007.n51 4.5005
R54514 a_33379_34007.n203 a_33379_34007.n202 4.5005
R54515 a_33379_34007.n201 a_33379_34007.n196 4.5005
R54516 a_33379_34007.n53 a_33379_34007.n52 4.5005
R54517 a_33379_34007.n200 a_33379_34007.n199 4.5005
R54518 a_33379_34007.n198 a_33379_34007.n197 4.5005
R54519 a_33379_34007.n242 a_33379_34007.n241 4.5005
R54520 a_33379_34007.n245 a_33379_34007.n244 4.5005
R54521 a_33379_34007.n246 a_33379_34007.n240 4.5005
R54522 a_33379_34007.n248 a_33379_34007.n247 4.5005
R54523 a_33379_34007.n49 a_33379_34007.n239 4.5005
R54524 a_33379_34007.n249 a_33379_34007.n50 4.5005
R54525 a_33379_34007.n251 a_33379_34007.n250 4.5005
R54526 a_33379_34007.n256 a_33379_34007.n255 4.5005
R54527 a_33379_34007.n36 a_33379_34007.n35 4.5005
R54528 a_33379_34007.n257 a_33379_34007.n114 4.5005
R54529 a_33379_34007.n259 a_33379_34007.n258 4.5005
R54530 a_33379_34007.n260 a_33379_34007.n19 4.5005
R54531 a_33379_34007.n262 a_33379_34007.n261 4.5005
R54532 a_33379_34007.n263 a_33379_34007.n113 4.5005
R54533 a_33379_34007.n266 a_33379_34007.n265 4.5005
R54534 a_33379_34007.n267 a_33379_34007.n112 4.5005
R54535 a_33379_34007.n46 a_33379_34007.n268 4.5005
R54536 a_33379_34007.n270 a_33379_34007.n269 4.5005
R54537 a_33379_34007.n17 a_33379_34007.n111 4.5005
R54538 a_33379_34007.n271 a_33379_34007.n18 4.5005
R54539 a_33379_34007.n272 a_33379_34007.n16 4.5005
R54540 a_33379_34007.n274 a_33379_34007.n273 4.5005
R54541 a_33379_34007.n276 a_33379_34007.n110 4.5005
R54542 a_33379_34007.n278 a_33379_34007.n277 4.5005
R54543 a_33379_34007.n279 a_33379_34007.n44 4.5005
R54544 a_33379_34007.n45 a_33379_34007.n43 4.5005
R54545 a_33379_34007.n280 a_33379_34007.n109 4.5005
R54546 a_33379_34007.n293 a_33379_34007.n292 4.5005
R54547 a_33379_34007.n32 a_33379_34007.n30 4.5005
R54548 a_33379_34007.n31 a_33379_34007.n291 4.5005
R54549 a_33379_34007.n290 a_33379_34007.n14 4.5005
R54550 a_33379_34007.n289 a_33379_34007.n15 4.5005
R54551 a_33379_34007.n13 a_33379_34007.n284 4.5005
R54552 a_33379_34007.n288 a_33379_34007.n287 4.5005
R54553 a_33379_34007.n314 a_33379_34007.n313 4.5005
R54554 a_33379_34007.n311 a_33379_34007.n106 4.5005
R54555 a_33379_34007.n105 a_33379_34007.n302 4.5005
R54556 a_33379_34007.n310 a_33379_34007.n309 4.5005
R54557 a_33379_34007.n308 a_33379_34007.n104 4.5005
R54558 a_33379_34007.n103 a_33379_34007.n303 4.5005
R54559 a_33379_34007.n307 a_33379_34007.n306 4.5005
R54560 a_33379_34007.n93 a_33379_34007.n301 4.5005
R54561 a_33379_34007.n318 a_33379_34007.n94 4.5005
R54562 a_33379_34007.n320 a_33379_34007.n319 4.5005
R54563 a_33379_34007.n95 a_33379_34007.n300 4.5005
R54564 a_33379_34007.n321 a_33379_34007.n96 4.5005
R54565 a_33379_34007.n323 a_33379_34007.n322 4.5005
R54566 a_33379_34007.n97 a_33379_34007.n299 4.5005
R54567 a_33379_34007.n324 a_33379_34007.n99 4.5005
R54568 a_33379_34007.n325 a_33379_34007.n98 4.5005
R54569 a_33379_34007.n100 a_33379_34007.n326 4.5005
R54570 a_33379_34007.n336 a_33379_34007.n296 4.5005
R54571 a_33379_34007.n92 a_33379_34007.n90 4.5005
R54572 a_33379_34007.n335 a_33379_34007.n91 4.5005
R54573 a_33379_34007.n334 a_33379_34007.n333 4.5005
R54574 a_33379_34007.n89 a_33379_34007.n87 4.5005
R54575 a_33379_34007.n88 a_33379_34007.n332 4.5005
R54576 a_33379_34007.n331 a_33379_34007.n85 4.5005
R54577 a_33379_34007.n330 a_33379_34007.n86 4.5005
R54578 a_33379_34007.n84 a_33379_34007.n297 4.5005
R54579 a_33379_34007.n329 a_33379_34007.n328 4.5005
R54580 a_33379_34007.n347 a_33379_34007.n346 4.5005
R54581 a_33379_34007.n78 a_33379_34007.n76 4.5005
R54582 a_33379_34007.n77 a_33379_34007.n345 4.5005
R54583 a_33379_34007.n344 a_33379_34007.n79 4.5005
R54584 a_33379_34007.n343 a_33379_34007.n81 4.5005
R54585 a_33379_34007.n80 a_33379_34007.n340 4.5005
R54586 a_33379_34007.n342 a_33379_34007.n341 4.5005
R54587 a_33379_34007.n1 a_33379_34007.n0 0.49013
R54588 a_33379_34007.t27 a_33379_34007.n1 7.88634
R54589 a_33379_34007.n135 a_33379_34007.n108 2.30989
R54590 a_33379_34007.n236 a_33379_34007.n176 2.30989
R54591 a_33379_34007.n223 a_33379_34007.n222 2.25752
R54592 a_33379_34007.n327 a_33379_34007.n298 2.25752
R54593 a_33379_34007.n176 a_33379_34007.n115 2.18975
R54594 a_33379_34007.n152 a_33379_34007.n135 2.18975
R54595 a_33379_34007.n250 a_33379_34007.n238 2.18975
R54596 a_33379_34007.n294 a_33379_34007.n109 2.18975
R54597 a_33379_34007.n235 a_33379_34007.n177 2.16725
R54598 a_33379_34007.n211 a_33379_34007.n195 2.16725
R54599 a_33379_34007.n313 a_33379_34007.n312 2.16725
R54600 a_33379_34007.n348 a_33379_34007.n296 2.16725
R54601 a_33379_34007.n349 a_33379_34007.n348 1.5005
R54602 a_33379_34007.n295 a_33379_34007.n294 1.5005
R54603 a_33379_34007.n195 a_33379_34007.n108 1.5005
R54604 a_33379_34007.n312 a_33379_34007.n107 1.5005
R54605 a_33379_34007.n238 a_33379_34007.n237 1.5005
R54606 a_33379_34007.n236 a_33379_34007.n235 1.5005
R54607 a_33379_34007.n10 a_33379_34007.t87 8.40801
R54608 a_33379_34007.n21 a_33379_34007.t90 8.40801
R54609 a_33379_34007.n148 a_33379_34007.n147 1.24866
R54610 a_33379_34007.n174 a_33379_34007.n128 1.24866
R54611 a_33379_34007.n292 a_33379_34007.n283 1.24866
R54612 a_33379_34007.n255 a_33379_34007.n254 1.24866
R54613 a_33379_34007.n151 a_33379_34007.n150 1.24629
R54614 a_33379_34007.n126 a_33379_34007.n125 1.24629
R54615 a_33379_34007.n281 a_33379_34007.n280 1.24629
R54616 a_33379_34007.n252 a_33379_34007.n251 1.24629
R54617 a_33379_34007.n295 a_33379_34007.n108 1.23709
R54618 a_33379_34007.n237 a_33379_34007.n236 1.23709
R54619 a_33379_34007.n210 a_33379_34007.n209 1.22261
R54620 a_33379_34007.n187 a_33379_34007.n186 1.22261
R54621 a_33379_34007.n337 a_33379_34007.n336 1.22261
R54622 a_33379_34007.n315 a_33379_34007.n314 1.22261
R54623 a_33379_34007.n207 a_33379_34007.n206 1.21313
R54624 a_33379_34007.n233 a_33379_34007.n189 1.21313
R54625 a_33379_34007.n346 a_33379_34007.n339 1.21313
R54626 a_33379_34007.n93 a_33379_34007.n317 1.21313
R54627 a_33379_34007.n181 a_33379_34007.n180 1.12904
R54628 a_33379_34007.n306 a_33379_34007.n305 1.12904
R54629 a_33379_34007.n140 a_33379_34007.n139 1.11862
R54630 a_33379_34007.n287 a_33379_34007.n286 1.11862
R54631 a_33379_34007.n349 a_33379_34007.n295 0.809892
R54632 a_33379_34007.n237 a_33379_34007.n107 0.809892
R54633 a_33379_34007.t0 a_33379_34007.n1 0.311051
R54634 a_33379_34007.n176 a_33379_34007.n175 0.752
R54635 a_33379_34007.n146 a_33379_34007.n135 0.752
R54636 a_33379_34007.n256 a_33379_34007.n238 0.752
R54637 a_33379_34007.n294 a_33379_34007.n293 0.752
R54638 a_33379_34007.n235 a_33379_34007.n234 0.71825
R54639 a_33379_34007.n205 a_33379_34007.n195 0.71825
R54640 a_33379_34007.n312 a_33379_34007.n301 0.71825
R54641 a_33379_34007.n348 a_33379_34007.n347 0.71825
R54642 a_33379_34007.n150 a_33379_34007.n149 0.673132
R54643 a_33379_34007.n149 a_33379_34007.n148 0.673132
R54644 a_33379_34007.n127 a_33379_34007.n126 0.673132
R54645 a_33379_34007.n128 a_33379_34007.n127 0.673132
R54646 a_33379_34007.n209 a_33379_34007.n208 0.673132
R54647 a_33379_34007.n208 a_33379_34007.n207 0.673132
R54648 a_33379_34007.n188 a_33379_34007.n187 0.673132
R54649 a_33379_34007.n189 a_33379_34007.n188 0.673132
R54650 a_33379_34007.n282 a_33379_34007.n281 0.673132
R54651 a_33379_34007.n283 a_33379_34007.n282 0.673132
R54652 a_33379_34007.n253 a_33379_34007.n252 0.673132
R54653 a_33379_34007.n254 a_33379_34007.n253 0.673132
R54654 a_33379_34007.n338 a_33379_34007.n337 0.673132
R54655 a_33379_34007.n339 a_33379_34007.n338 0.673132
R54656 a_33379_34007.n316 a_33379_34007.n315 0.673132
R54657 a_33379_34007.n317 a_33379_34007.n316 0.673132
R54658 a_33379_34007.n350 a_33379_34007.n107 0.647527
R54659 a_33379_34007.n55 a_33379_34007.n54 0.321834
R54660 a_33379_34007.n83 a_33379_34007.n82 0.321834
R54661 a_33379_34007.n12 a_33379_34007.n10 0.307602
R54662 a_33379_34007.n21 a_33379_34007.n20 0.307602
R54663 a_33379_34007.n2 a_33379_34007.n141 0.394842
R54664 a_33379_34007.n4 a_33379_34007.n160 0.394842
R54665 a_33379_34007.n7 a_33379_34007.n170 0.394842
R54666 a_33379_34007.n119 a_33379_34007.n11 0.394842
R54667 a_33379_34007.n13 a_33379_34007.n288 0.394842
R54668 a_33379_34007.n274 a_33379_34007.n16 0.394842
R54669 a_33379_34007.n263 a_33379_34007.n262 0.394842
R54670 a_33379_34007.n244 a_33379_34007.n242 0.394842
R54671 a_33379_34007.n22 a_33379_34007.n144 0.381816
R54672 a_33379_34007.n24 a_33379_34007.n5 0.381816
R54673 a_33379_34007.n28 a_33379_34007.n8 0.381816
R54674 a_33379_34007.n31 a_33379_34007.n14 0.381816
R54675 a_33379_34007.n17 a_33379_34007.n270 0.381816
R54676 a_33379_34007.n258 a_33379_34007.n257 0.381816
R54677 a_33379_34007.n202 a_33379_34007.n201 0.379447
R54678 a_33379_34007.n199 a_33379_34007.n198 0.379447
R54679 a_33379_34007.n221 a_33379_34007.n220 0.379447
R54680 a_33379_34007.n216 a_33379_34007.n215 0.379447
R54681 a_33379_34007.n213 a_33379_34007.n212 0.379447
R54682 a_33379_34007.n62 a_33379_34007.n64 0.379447
R54683 a_33379_34007.n65 a_33379_34007.n229 0.379447
R54684 a_33379_34007.n225 a_33379_34007.n224 0.379447
R54685 a_33379_34007.n71 a_33379_34007.n178 0.379447
R54686 a_33379_34007.n183 a_33379_34007.n74 0.379447
R54687 a_33379_34007.n77 a_33379_34007.n79 0.379447
R54688 a_33379_34007.n80 a_33379_34007.n342 0.379447
R54689 a_33379_34007.n84 a_33379_34007.n329 0.379447
R54690 a_33379_34007.n88 a_33379_34007.n85 0.379447
R54691 a_33379_34007.n333 a_33379_34007.n91 0.379447
R54692 a_33379_34007.n95 a_33379_34007.n320 0.379447
R54693 a_33379_34007.n97 a_33379_34007.n323 0.379447
R54694 a_33379_34007.n100 a_33379_34007.n98 0.379447
R54695 a_33379_34007.n103 a_33379_34007.n307 0.379447
R54696 a_33379_34007.n105 a_33379_34007.n310 0.379447
R54697 a_33379_34007.n118 a_33379_34007.n117 0.375125
R54698 a_33379_34007.n169 a_33379_34007.n129 0.375125
R54699 a_33379_34007.n159 a_33379_34007.n132 0.375125
R54700 a_33379_34007.n140 a_33379_34007.n137 0.375125
R54701 a_33379_34007.n245 a_33379_34007.n241 0.375125
R54702 a_33379_34007.n261 a_33379_34007.n113 0.375125
R54703 a_33379_34007.n273 a_33379_34007.n272 0.375125
R54704 a_33379_34007.n287 a_33379_34007.n284 0.375125
R54705 a_33379_34007.n173 a_33379_34007.n172 0.36275
R54706 a_33379_34007.n163 a_33379_34007.n162 0.36275
R54707 a_33379_34007.n143 a_33379_34007.n136 0.36275
R54708 a_33379_34007.n259 a_33379_34007.n114 0.36275
R54709 a_33379_34007.n269 a_33379_34007.n111 0.36275
R54710 a_33379_34007.n291 a_33379_34007.n290 0.36275
R54711 a_33379_34007.n182 a_33379_34007.n181 0.3605
R54712 a_33379_34007.n185 a_33379_34007.n184 0.3605
R54713 a_33379_34007.n232 a_33379_34007.n231 0.3605
R54714 a_33379_34007.n228 a_33379_34007.n190 0.3605
R54715 a_33379_34007.n226 a_33379_34007.n191 0.3605
R54716 a_33379_34007.n219 a_33379_34007.n192 0.3605
R54717 a_33379_34007.n217 a_33379_34007.n193 0.3605
R54718 a_33379_34007.n214 a_33379_34007.n194 0.3605
R54719 a_33379_34007.n203 a_33379_34007.n196 0.3605
R54720 a_33379_34007.n200 a_33379_34007.n197 0.3605
R54721 a_33379_34007.n306 a_33379_34007.n303 0.3605
R54722 a_33379_34007.n309 a_33379_34007.n302 0.3605
R54723 a_33379_34007.n319 a_33379_34007.n300 0.3605
R54724 a_33379_34007.n322 a_33379_34007.n299 0.3605
R54725 a_33379_34007.n326 a_33379_34007.n325 0.3605
R54726 a_33379_34007.n328 a_33379_34007.n297 0.3605
R54727 a_33379_34007.n332 a_33379_34007.n331 0.3605
R54728 a_33379_34007.n335 a_33379_34007.n334 0.3605
R54729 a_33379_34007.n345 a_33379_34007.n344 0.3605
R54730 a_33379_34007.n341 a_33379_34007.n340 0.3605
R54731 a_33379_34007.n139 a_33379_34007.n138 0.348488
R54732 a_33379_34007.n286 a_33379_34007.n285 0.348488
R54733 a_33379_34007.n180 a_33379_34007.n179 0.327481
R54734 a_33379_34007.n305 a_33379_34007.n304 0.327481
R54735 a_33379_34007.n156 a_33379_34007.n155 0.302474
R54736 a_33379_34007.n166 a_33379_34007.n165 0.302474
R54737 a_33379_34007.n122 a_33379_34007.n41 0.302474
R54738 a_33379_34007.n277 a_33379_34007.n44 0.302474
R54739 a_33379_34007.n46 a_33379_34007.n112 0.302474
R54740 a_33379_34007.n49 a_33379_34007.n248 0.302474
R54741 a_33379_34007.n124 a_33379_34007.n123 0.287375
R54742 a_33379_34007.n164 a_33379_34007.n131 0.287375
R54743 a_33379_34007.n154 a_33379_34007.n134 0.287375
R54744 a_33379_34007.n247 a_33379_34007.n239 0.287375
R54745 a_33379_34007.n268 a_33379_34007.n267 0.287375
R54746 a_33379_34007.n279 a_33379_34007.n278 0.287375
R54747 a_33379_34007.n223 a_33379_34007.n192 0.208099
R54748 a_33379_34007.n328 a_33379_34007.n327 0.208099
R54749 a_33379_34007.n101 a_33379_34007.n100 0.152079
R54750 a_33379_34007.n314 a_33379_34007.n106 0.147342
R54751 a_33379_34007.n310 a_33379_34007.n104 0.147342
R54752 a_33379_34007.n23 a_33379_34007.n22 0.147342
R54753 a_33379_34007.n3 a_33379_34007.n2 0.147342
R54754 a_33379_34007.n6 a_33379_34007.n4 0.147342
R54755 a_33379_34007.n157 a_33379_34007.n156 0.147342
R54756 a_33379_34007.n155 a_33379_34007.n37 0.147342
R54757 a_33379_34007.n29 a_33379_34007.n28 0.147342
R54758 a_33379_34007.n9 a_33379_34007.n7 0.147342
R54759 a_33379_34007.n167 a_33379_34007.n166 0.147342
R54760 a_33379_34007.n122 a_33379_34007.n121 0.147342
R54761 a_33379_34007.n42 a_33379_34007.n41 0.147342
R54762 a_33379_34007.n206 a_33379_34007.n51 0.147342
R54763 a_33379_34007.n201 a_33379_34007.n53 0.147342
R54764 a_33379_34007.n220 a_33379_34007.n56 0.147342
R54765 a_33379_34007.n215 a_33379_34007.n58 0.147342
R54766 a_33379_34007.n212 a_33379_34007.n60 0.147342
R54767 a_33379_34007.n233 a_33379_34007.n63 0.147342
R54768 a_33379_34007.n66 a_33379_34007.n64 0.147342
R54769 a_33379_34007.n229 a_33379_34007.n67 0.147342
R54770 a_33379_34007.n72 a_33379_34007.n71 0.147342
R54771 a_33379_34007.n75 a_33379_34007.n74 0.147342
R54772 a_33379_34007.n32 a_33379_34007.n31 0.147342
R54773 a_33379_34007.n15 a_33379_34007.n13 0.147342
R54774 a_33379_34007.n18 a_33379_34007.n16 0.147342
R54775 a_33379_34007.n277 a_33379_34007.n276 0.147342
R54776 a_33379_34007.n45 a_33379_34007.n44 0.147342
R54777 a_33379_34007.n257 a_33379_34007.n36 0.147342
R54778 a_33379_34007.n262 a_33379_34007.n19 0.147342
R54779 a_33379_34007.n265 a_33379_34007.n112 0.147342
R54780 a_33379_34007.n248 a_33379_34007.n240 0.147342
R54781 a_33379_34007.n50 a_33379_34007.n49 0.147342
R54782 a_33379_34007.n346 a_33379_34007.n78 0.147342
R54783 a_33379_34007.n81 a_33379_34007.n79 0.147342
R54784 a_33379_34007.n86 a_33379_34007.n84 0.147342
R54785 a_33379_34007.n89 a_33379_34007.n88 0.147342
R54786 a_33379_34007.n92 a_33379_34007.n91 0.147342
R54787 a_33379_34007.n94 a_33379_34007.n93 0.147342
R54788 a_33379_34007.n96 a_33379_34007.n95 0.147342
R54789 a_33379_34007.n99 a_33379_34007.n97 0.147342
R54790 a_33379_34007.n104 a_33379_34007.n103 0.147342
R54791 a_33379_34007.n106 a_33379_34007.n105 0.147342
R54792 a_33379_34007.n222 a_33379_34007.n221 0.142605
R54793 a_33379_34007.n179 a_33379_34007.n178 0.142605
R54794 a_33379_34007.n329 a_33379_34007.n298 0.142605
R54795 a_33379_34007.n307 a_33379_34007.n304 0.142605
R54796 a_33379_34007.n117 a_33379_34007.n10 1.12843
R54797 a_33379_34007.n118 a_33379_34007.n116 0.14
R54798 a_33379_34007.n123 a_33379_34007.n116 0.14
R54799 a_33379_34007.n40 a_33379_34007.n124 0.14
R54800 a_33379_34007.n40 a_33379_34007.n115 0.14
R54801 a_33379_34007.n175 a_33379_34007.n27 0.14
R54802 a_33379_34007.n173 a_33379_34007.n27 0.14
R54803 a_33379_34007.n172 a_33379_34007.n171 0.14
R54804 a_33379_34007.n171 a_33379_34007.n129 0.14
R54805 a_33379_34007.n169 a_33379_34007.n168 0.14
R54806 a_33379_34007.n168 a_33379_34007.n131 0.14
R54807 a_33379_34007.n164 a_33379_34007.n39 0.208307
R54808 a_33379_34007.n39 a_33379_34007.n26 3.16466
R54809 a_33379_34007.n163 a_33379_34007.n26 0.208324
R54810 a_33379_34007.n162 a_33379_34007.n161 0.14
R54811 a_33379_34007.n161 a_33379_34007.n132 0.14
R54812 a_33379_34007.n159 a_33379_34007.n158 0.14
R54813 a_33379_34007.n158 a_33379_34007.n134 0.14
R54814 a_33379_34007.n154 a_33379_34007.n153 0.14
R54815 a_33379_34007.n153 a_33379_34007.n152 0.14
R54816 a_33379_34007.n146 a_33379_34007.n145 0.14
R54817 a_33379_34007.n145 a_33379_34007.n136 0.14
R54818 a_33379_34007.n143 a_33379_34007.n142 0.14
R54819 a_33379_34007.n142 a_33379_34007.n137 0.14
R54820 a_33379_34007.n182 a_33379_34007.n70 0.14
R54821 a_33379_34007.n184 a_33379_34007.n70 0.14
R54822 a_33379_34007.n73 a_33379_34007.n185 0.14
R54823 a_33379_34007.n73 a_33379_34007.n177 0.14
R54824 a_33379_34007.n234 a_33379_34007.n61 0.14
R54825 a_33379_34007.n232 a_33379_34007.n61 0.14
R54826 a_33379_34007.n231 a_33379_34007.n230 0.14
R54827 a_33379_34007.n230 a_33379_34007.n190 0.14
R54828 a_33379_34007.n228 a_33379_34007.n227 0.14
R54829 a_33379_34007.n227 a_33379_34007.n226 0.14
R54830 a_33379_34007.n69 a_33379_34007.n191 0.208134
R54831 a_33379_34007.n69 a_33379_34007.n223 3.10882
R54832 a_33379_34007.n219 a_33379_34007.n218 0.14
R54833 a_33379_34007.n218 a_33379_34007.n217 0.14
R54834 a_33379_34007.n57 a_33379_34007.n193 0.14
R54835 a_33379_34007.n57 a_33379_34007.n214 0.14
R54836 a_33379_34007.n59 a_33379_34007.n194 0.14
R54837 a_33379_34007.n59 a_33379_34007.n211 0.14
R54838 a_33379_34007.n205 a_33379_34007.n204 0.14
R54839 a_33379_34007.n204 a_33379_34007.n203 0.14
R54840 a_33379_34007.n52 a_33379_34007.n196 0.14
R54841 a_33379_34007.n52 a_33379_34007.n200 0.14
R54842 a_33379_34007.n55 a_33379_34007.n197 1.12757
R54843 a_33379_34007.n21 a_33379_34007.n241 1.12843
R54844 a_33379_34007.n246 a_33379_34007.n245 0.14
R54845 a_33379_34007.n247 a_33379_34007.n246 0.14
R54846 a_33379_34007.n249 a_33379_34007.n239 0.14
R54847 a_33379_34007.n250 a_33379_34007.n249 0.14
R54848 a_33379_34007.n35 a_33379_34007.n256 0.14
R54849 a_33379_34007.n35 a_33379_34007.n114 0.14
R54850 a_33379_34007.n260 a_33379_34007.n259 0.14
R54851 a_33379_34007.n261 a_33379_34007.n260 0.14
R54852 a_33379_34007.n266 a_33379_34007.n113 0.14
R54853 a_33379_34007.n267 a_33379_34007.n266 0.14
R54854 a_33379_34007.n268 a_33379_34007.n48 0.208307
R54855 a_33379_34007.n34 a_33379_34007.n48 3.16466
R54856 a_33379_34007.n269 a_33379_34007.n34 0.208324
R54857 a_33379_34007.n271 a_33379_34007.n111 0.14
R54858 a_33379_34007.n272 a_33379_34007.n271 0.14
R54859 a_33379_34007.n273 a_33379_34007.n110 0.14
R54860 a_33379_34007.n278 a_33379_34007.n110 0.14
R54861 a_33379_34007.n43 a_33379_34007.n279 0.14
R54862 a_33379_34007.n43 a_33379_34007.n109 0.14
R54863 a_33379_34007.n293 a_33379_34007.n30 0.14
R54864 a_33379_34007.n291 a_33379_34007.n30 0.14
R54865 a_33379_34007.n290 a_33379_34007.n289 0.14
R54866 a_33379_34007.n289 a_33379_34007.n284 0.14
R54867 a_33379_34007.n308 a_33379_34007.n303 0.14
R54868 a_33379_34007.n309 a_33379_34007.n308 0.14
R54869 a_33379_34007.n311 a_33379_34007.n302 0.14
R54870 a_33379_34007.n313 a_33379_34007.n311 0.14
R54871 a_33379_34007.n318 a_33379_34007.n301 0.14
R54872 a_33379_34007.n319 a_33379_34007.n318 0.14
R54873 a_33379_34007.n321 a_33379_34007.n300 0.14
R54874 a_33379_34007.n322 a_33379_34007.n321 0.14
R54875 a_33379_34007.n324 a_33379_34007.n299 0.14
R54876 a_33379_34007.n325 a_33379_34007.n324 0.14
R54877 a_33379_34007.n326 a_33379_34007.n102 0.208134
R54878 a_33379_34007.n327 a_33379_34007.n102 3.10882
R54879 a_33379_34007.n342 a_33379_34007.n82 0.152079
R54880 a_33379_34007.n99 a_33379_34007.n98 0.147342
R54881 a_33379_34007.n323 a_33379_34007.n96 0.147342
R54882 a_33379_34007.n320 a_33379_34007.n94 0.147342
R54883 a_33379_34007.n336 a_33379_34007.n92 0.147342
R54884 a_33379_34007.n333 a_33379_34007.n89 0.147342
R54885 a_33379_34007.n86 a_33379_34007.n85 0.147342
R54886 a_33379_34007.n330 a_33379_34007.n297 0.14
R54887 a_33379_34007.n331 a_33379_34007.n330 0.14
R54888 a_33379_34007.n332 a_33379_34007.n87 0.14
R54889 a_33379_34007.n334 a_33379_34007.n87 0.14
R54890 a_33379_34007.n90 a_33379_34007.n335 0.14
R54891 a_33379_34007.n90 a_33379_34007.n296 0.14
R54892 a_33379_34007.n347 a_33379_34007.n76 0.14
R54893 a_33379_34007.n345 a_33379_34007.n76 0.14
R54894 a_33379_34007.n344 a_33379_34007.n343 0.14
R54895 a_33379_34007.n343 a_33379_34007.n340 0.14
R54896 a_33379_34007.n341 a_33379_34007.n83 1.12757
R54897 a_33379_34007.n242 a_33379_34007.n20 0.1805
R54898 a_33379_34007.n12 a_33379_34007.n11 0.1805
R54899 a_33379_34007.n270 a_33379_34007.n33 0.178132
R54900 a_33379_34007.n25 a_33379_34007.n24 0.178132
R54901 a_33379_34007.n47 a_33379_34007.n46 0.175763
R54902 a_33379_34007.n165 a_33379_34007.n38 0.175763
R54903 a_33379_34007.n224 a_33379_34007.n68 0.152079
R54904 a_33379_34007.n198 a_33379_34007.n54 0.152079
R54905 a_33379_34007.n81 a_33379_34007.n80 0.147342
R54906 a_33379_34007.n78 a_33379_34007.n77 0.147342
R54907 a_33379_34007.n186 a_33379_34007.n75 0.147342
R54908 a_33379_34007.n183 a_33379_34007.n72 0.147342
R54909 a_33379_34007.n225 a_33379_34007.n67 0.147342
R54910 a_33379_34007.n66 a_33379_34007.n65 0.147342
R54911 a_33379_34007.n63 a_33379_34007.n62 0.147342
R54912 a_33379_34007.n210 a_33379_34007.n60 0.147342
R54913 a_33379_34007.n213 a_33379_34007.n58 0.147342
R54914 a_33379_34007.n216 a_33379_34007.n56 0.147342
R54915 a_33379_34007.n199 a_33379_34007.n53 0.147342
R54916 a_33379_34007.n202 a_33379_34007.n51 0.147342
R54917 a_33379_34007.n251 a_33379_34007.n50 0.147342
R54918 a_33379_34007.n280 a_33379_34007.n45 0.147342
R54919 a_33379_34007.n125 a_33379_34007.n42 0.147342
R54920 a_33379_34007.n151 a_33379_34007.n37 0.147342
R54921 a_33379_34007.n255 a_33379_34007.n36 0.147342
R54922 a_33379_34007.n292 a_33379_34007.n32 0.147342
R54923 a_33379_34007.n174 a_33379_34007.n29 0.147342
R54924 a_33379_34007.n147 a_33379_34007.n23 0.147342
R54925 a_33379_34007.n258 a_33379_34007.n19 0.147342
R54926 a_33379_34007.n18 a_33379_34007.n17 0.147342
R54927 a_33379_34007.n15 a_33379_34007.n14 0.147342
R54928 a_33379_34007.n9 a_33379_34007.n8 0.147342
R54929 a_33379_34007.n6 a_33379_34007.n5 0.147342
R54930 a_33379_34007.n144 a_33379_34007.n3 0.147342
R54931 a_33379_34007.n141 a_33379_34007.n138 0.0987895
R54932 a_33379_34007.n160 a_33379_34007.n133 0.0987895
R54933 a_33379_34007.n170 a_33379_34007.n130 0.0987895
R54934 a_33379_34007.n120 a_33379_34007.n119 0.0987895
R54935 a_33379_34007.n288 a_33379_34007.n285 0.0987895
R54936 a_33379_34007.n275 a_33379_34007.n274 0.0987895
R54937 a_33379_34007.n264 a_33379_34007.n263 0.0987895
R54938 a_33379_34007.n244 a_33379_34007.n243 0.0987895
R54939 a_33379_34007.n157 a_33379_34007.n133 0.0490526
R54940 a_33379_34007.n167 a_33379_34007.n130 0.0490526
R54941 a_33379_34007.n121 a_33379_34007.n120 0.0490526
R54942 a_33379_34007.n276 a_33379_34007.n275 0.0490526
R54943 a_33379_34007.n265 a_33379_34007.n264 0.0490526
R54944 a_33379_34007.n243 a_33379_34007.n240 0.0490526
R54945 a_33379_34007.n0 a_33379_34007.t1 0.295568
R54946 a_33379_34007.n0 a_33379_34007.n351 16.9974
R54947 a_33249_34067.n114 a_33249_34067.n113 8.18538
R54948 a_33249_34067.n125 a_33249_34067.n123 7.22198
R54949 a_33249_34067.n153 a_33249_34067.n28 7.22198
R54950 a_33249_34067.n30 a_33249_34067.t23 6.77653
R54951 a_33249_34067.n132 a_33249_34067.t20 6.77653
R54952 a_33249_34067.n48 a_33249_34067.t77 6.7761
R54953 a_33249_34067.n145 a_33249_34067.t74 6.7761
R54954 a_33249_34067.n25 a_33249_34067.t133 6.86989
R54955 a_33249_34067.n9 a_33249_34067.t101 6.77231
R54956 a_33249_34067.n19 a_33249_34067.t89 6.77231
R54957 a_33249_34067.n109 a_33249_34067.t7 6.53862
R54958 a_33249_34067.n114 a_33249_34067.n55 5.95467
R54959 a_33249_34067.n79 a_33249_34067.n77 5.89898
R54960 a_33249_34067.n93 a_33249_34067.t126 5.66511
R54961 a_33249_34067.n86 a_33249_34067.t111 5.66511
R54962 a_33249_34067.n94 a_33249_34067.t131 5.66379
R54963 a_33249_34067.n87 a_33249_34067.t116 5.66379
R54964 a_33249_34067.n86 a_33249_34067.n85 5.65285
R54965 a_33249_34067.n73 a_33249_34067.t130 5.61877
R54966 a_33249_34067.n74 a_33249_34067.t109 5.61877
R54967 a_33249_34067.n70 a_33249_34067.t114 5.61877
R54968 a_33249_34067.n45 a_33249_34067.t65 5.50607
R54969 a_33249_34067.n31 a_33249_34067.t36 5.50607
R54970 a_33249_34067.n142 a_33249_34067.t59 5.50607
R54971 a_33249_34067.n133 a_33249_34067.t31 5.50607
R54972 a_33249_34067.n46 a_33249_34067.t97 5.50475
R54973 a_33249_34067.n42 a_33249_34067.t62 5.50475
R54974 a_33249_34067.n41 a_33249_34067.t72 5.50475
R54975 a_33249_34067.n32 a_33249_34067.t69 5.50475
R54976 a_33249_34067.n143 a_33249_34067.t92 5.50475
R54977 a_33249_34067.n139 a_33249_34067.t56 5.50475
R54978 a_33249_34067.n138 a_33249_34067.t68 5.50475
R54979 a_33249_34067.n134 a_33249_34067.t64 5.50475
R54980 a_33249_34067.n112 a_33249_34067.t1 5.28484
R54981 a_33249_34067.n22 a_33249_34067.n99 5.29079
R54982 a_33249_34067.n96 a_33249_34067.n95 4.88835
R54983 a_33249_34067.n63 a_33249_34067.n62 4.88517
R54984 a_33249_34067.n100 a_33249_34067.n21 4.02009
R54985 a_33249_34067.t11 a_33249_34067.n20 5.28011
R54986 a_33249_34067.t10 a_33249_34067.n22 5.28011
R54987 a_33249_34067.n0 a_33249_34067.n38 4.0312
R54988 a_33249_34067.n1 a_33249_34067.t84 5.5012
R54989 a_33249_34067.n2 a_33249_34067.t54 5.5012
R54990 a_33249_34067.n3 a_33249_34067.n37 4.0312
R54991 a_33249_34067.n4 a_33249_34067.t50 5.5012
R54992 a_33249_34067.n5 a_33249_34067.t61 5.5012
R54993 a_33249_34067.n6 a_33249_34067.n36 4.0312
R54994 a_33249_34067.t57 a_33249_34067.n7 5.5012
R54995 a_33249_34067.t26 a_33249_34067.n8 5.5012
R54996 a_33249_34067.n35 a_33249_34067.n9 4.0312
R54997 a_33249_34067.n10 a_33249_34067.n118 4.0312
R54998 a_33249_34067.n11 a_33249_34067.t79 5.5012
R54999 a_33249_34067.n12 a_33249_34067.t45 5.5012
R55000 a_33249_34067.n13 a_33249_34067.n117 4.0312
R55001 a_33249_34067.n14 a_33249_34067.t39 5.5012
R55002 a_33249_34067.n15 a_33249_34067.t51 5.5012
R55003 a_33249_34067.n16 a_33249_34067.n116 4.0312
R55004 a_33249_34067.t48 a_33249_34067.n17 5.5012
R55005 a_33249_34067.t18 a_33249_34067.n18 5.5012
R55006 a_33249_34067.n115 a_33249_34067.n19 4.0312
R55007 a_33249_34067.n23 a_33249_34067.n72 4.40099
R55008 a_33249_34067.n24 a_33249_34067.n71 4.40099
R55009 a_33249_34067.n69 a_33249_34067.n25 4.40099
R55010 a_33249_34067.n92 a_33249_34067.n91 4.40379
R55011 a_33249_34067.n90 a_33249_34067.n89 4.40379
R55012 a_33249_34067.n78 a_33249_34067.t136 4.40142
R55013 a_33249_34067.n64 a_33249_34067.t125 4.40142
R55014 a_33249_34067.n27 a_33249_34067.t52 4.24002
R55015 a_33249_34067.n26 a_33249_34067.t43 4.24002
R55016 a_33249_34067.n124 a_33249_34067.t41 4.24002
R55017 a_33249_34067.n56 a_33249_34067.t35 4.24002
R55018 a_33249_34067.n105 a_33249_34067.t3 4.22616
R55019 a_33249_34067.n48 a_33249_34067.n47 4.03475
R55020 a_33249_34067.n44 a_33249_34067.n43 4.03475
R55021 a_33249_34067.n40 a_33249_34067.n39 4.03475
R55022 a_33249_34067.n30 a_33249_34067.n29 4.03475
R55023 a_33249_34067.n145 a_33249_34067.n144 4.03475
R55024 a_33249_34067.n141 a_33249_34067.n140 4.03475
R55025 a_33249_34067.n137 a_33249_34067.n136 4.03475
R55026 a_33249_34067.n132 a_33249_34067.n131 4.03475
R55027 a_33249_34067.n111 a_33249_34067.n110 4.02484
R55028 a_33249_34067.n109 a_33249_34067.n108 4.02484
R55029 a_33249_34067.n105 a_33249_34067.t9 4.02247
R55030 a_33249_34067.n107 a_33249_34067.n106 3.96014
R55031 a_33249_34067.n98 a_33249_34067.n61 3.94195
R55032 a_33249_34067.n78 a_33249_34067.t141 3.84721
R55033 a_33249_34067.n64 a_33249_34067.t129 3.84721
R55034 a_33249_34067.n92 a_33249_34067.n90 3.81703
R55035 a_33249_34067.n111 a_33249_34067.n109 3.80578
R55036 a_33249_34067.n27 a_33249_34067.t47 3.68818
R55037 a_33249_34067.n26 a_33249_34067.t38 3.68818
R55038 a_33249_34067.n124 a_33249_34067.t40 3.68818
R55039 a_33249_34067.n56 a_33249_34067.t34 3.68818
R55040 a_33249_34067.n130 a_33249_34067.n129 3.23904
R55041 a_33249_34067.n54 a_33249_34067.n53 3.23904
R55042 a_33249_34067.n84 a_33249_34067.n83 3.23004
R55043 a_33249_34067.n82 a_33249_34067.n81 3.14142
R55044 a_33249_34067.n67 a_33249_34067.n66 3.14142
R55045 a_33249_34067.n104 a_33249_34067.n102 2.96616
R55046 a_33249_34067.n52 a_33249_34067.n51 2.77002
R55047 a_33249_34067.n128 a_33249_34067.n127 2.77002
R55048 a_33249_34067.n59 a_33249_34067.n58 2.77002
R55049 a_33249_34067.n157 a_33249_34067.n156 2.77002
R55050 a_33249_34067.n104 a_33249_34067.n103 2.76247
R55051 a_33249_34067.n154 a_33249_34067.n26 2.7375
R55052 a_33249_34067.n60 a_33249_34067.n56 2.73714
R55053 a_33249_34067.n106 a_33249_34067.n104 2.71914
R55054 a_33249_34067.n68 a_33249_34067.n64 2.71914
R55055 a_33249_34067.n98 a_33249_34067.n97 2.64424
R55056 a_33249_34067.n42 a_33249_34067.n41 2.60203
R55057 a_33249_34067.n139 a_33249_34067.n138 2.60203
R55058 a_33249_34067.n82 a_33249_34067.n80 2.58721
R55059 a_33249_34067.n67 a_33249_34067.n65 2.58721
R55060 a_33249_34067.n87 a_33249_34067.n86 2.55136
R55061 a_33249_34067.n94 a_33249_34067.n93 2.55136
R55062 a_33249_34067.n32 a_33249_34067.n31 2.52436
R55063 a_33249_34067.n46 a_33249_34067.n45 2.52436
R55064 a_33249_34067.n134 a_33249_34067.n133 2.52436
R55065 a_33249_34067.n143 a_33249_34067.n142 2.52436
R55066 a_33249_34067.n76 a_33249_34067.n75 2.2807
R55067 a_33249_34067.n84 a_33249_34067.n63 2.2807
R55068 a_33249_34067.n52 a_33249_34067.n50 2.21818
R55069 a_33249_34067.n128 a_33249_34067.n126 2.21818
R55070 a_33249_34067.n59 a_33249_34067.n57 2.21818
R55071 a_33249_34067.n156 a_33249_34067.n155 2.21818
R55072 a_33249_34067.n152 a_33249_34067.n33 2.13841
R55073 a_33249_34067.n54 a_33249_34067.n49 2.13841
R55074 a_33249_34067.n123 a_33249_34067.n60 1.73904
R55075 a_33249_34067.n154 a_33249_34067.n153 1.73868
R55076 a_33249_34067.n113 a_33249_34067.n112 1.73609
R55077 a_33249_34067.n77 a_33249_34067.n68 1.73004
R55078 a_33249_34067.n121 a_33249_34067.n120 1.5005
R55079 a_33249_34067.n123 a_33249_34067.n122 1.5005
R55080 a_33249_34067.n135 a_33249_34067.n34 1.5005
R55081 a_33249_34067.n151 a_33249_34067.n150 1.5005
R55082 a_33249_34067.n77 a_33249_34067.n76 1.5005
R55083 a_33249_34067.n88 a_33249_34067.n61 1.5005
R55084 a_33249_34067.n97 a_33249_34067.n96 1.5005
R55085 a_33249_34067.n119 a_33249_34067.n55 1.5005
R55086 a_33249_34067.n147 a_33249_34067.n146 1.5005
R55087 a_33249_34067.n149 a_33249_34067.n148 1.5005
R55088 a_33249_34067.n153 a_33249_34067.n152 1.5005
R55089 a_33249_34067.n155 a_33249_34067.t98 1.4705
R55090 a_33249_34067.n155 a_33249_34067.t49 1.4705
R55091 a_33249_34067.n50 a_33249_34067.t19 1.4705
R55092 a_33249_34067.n50 a_33249_34067.t71 1.4705
R55093 a_33249_34067.n51 a_33249_34067.t24 1.4705
R55094 a_33249_34067.n51 a_33249_34067.t76 1.4705
R55095 a_33249_34067.n47 a_33249_34067.t37 1.4705
R55096 a_33249_34067.n47 a_33249_34067.t96 1.4705
R55097 a_33249_34067.n43 a_33249_34067.t32 1.4705
R55098 a_33249_34067.n43 a_33249_34067.t90 1.4705
R55099 a_33249_34067.n39 a_33249_34067.t30 1.4705
R55100 a_33249_34067.n39 a_33249_34067.t99 1.4705
R55101 a_33249_34067.n29 a_33249_34067.t88 1.4705
R55102 a_33249_34067.n29 a_33249_34067.t63 1.4705
R55103 a_33249_34067.n38 a_33249_34067.t28 1.4705
R55104 a_33249_34067.n38 a_33249_34067.t83 1.4705
R55105 a_33249_34067.n37 a_33249_34067.t25 1.4705
R55106 a_33249_34067.n37 a_33249_34067.t82 1.4705
R55107 a_33249_34067.n36 a_33249_34067.t22 1.4705
R55108 a_33249_34067.n36 a_33249_34067.t87 1.4705
R55109 a_33249_34067.n35 a_33249_34067.t81 1.4705
R55110 a_33249_34067.n35 a_33249_34067.t53 1.4705
R55111 a_33249_34067.n144 a_33249_34067.t33 1.4705
R55112 a_33249_34067.n144 a_33249_34067.t91 1.4705
R55113 a_33249_34067.n140 a_33249_34067.t29 1.4705
R55114 a_33249_34067.n140 a_33249_34067.t86 1.4705
R55115 a_33249_34067.n136 a_33249_34067.t27 1.4705
R55116 a_33249_34067.n136 a_33249_34067.t95 1.4705
R55117 a_33249_34067.n131 a_33249_34067.t85 1.4705
R55118 a_33249_34067.n131 a_33249_34067.t58 1.4705
R55119 a_33249_34067.n126 a_33249_34067.t102 1.4705
R55120 a_33249_34067.n126 a_33249_34067.t66 1.4705
R55121 a_33249_34067.n127 a_33249_34067.t103 1.4705
R55122 a_33249_34067.n127 a_33249_34067.t67 1.4705
R55123 a_33249_34067.n57 a_33249_34067.t93 1.4705
R55124 a_33249_34067.n57 a_33249_34067.t44 1.4705
R55125 a_33249_34067.n58 a_33249_34067.t94 1.4705
R55126 a_33249_34067.n58 a_33249_34067.t46 1.4705
R55127 a_33249_34067.n118 a_33249_34067.t21 1.4705
R55128 a_33249_34067.n118 a_33249_34067.t78 1.4705
R55129 a_33249_34067.n117 a_33249_34067.t104 1.4705
R55130 a_33249_34067.n117 a_33249_34067.t75 1.4705
R55131 a_33249_34067.n116 a_33249_34067.t100 1.4705
R55132 a_33249_34067.n116 a_33249_34067.t80 1.4705
R55133 a_33249_34067.n115 a_33249_34067.t73 1.4705
R55134 a_33249_34067.n115 a_33249_34067.t42 1.4705
R55135 a_33249_34067.t105 a_33249_34067.n157 1.4705
R55136 a_33249_34067.n157 a_33249_34067.t55 1.4705
R55137 a_33249_34067.n53 a_33249_34067.n52 1.46537
R55138 a_33249_34067.n28 a_33249_34067.n27 1.46537
R55139 a_33249_34067.n129 a_33249_34067.n128 1.46537
R55140 a_33249_34067.n125 a_33249_34067.n124 1.46537
R55141 a_33249_34067.n60 a_33249_34067.n59 1.46537
R55142 a_33249_34067.n83 a_33249_34067.n82 1.46537
R55143 a_33249_34067.n79 a_33249_34067.n78 1.46537
R55144 a_33249_34067.n68 a_33249_34067.n67 1.46537
R55145 a_33249_34067.n156 a_33249_34067.n154 1.46537
R55146 a_33249_34067.n106 a_33249_34067.n105 1.46537
R55147 a_33249_34067.n121 a_33249_34067.n114 1.37875
R55148 a_33249_34067.n41 a_33249_34067.n40 1.27228
R55149 a_33249_34067.n44 a_33249_34067.n42 1.27228
R55150 a_33249_34067.n138 a_33249_34067.n137 1.27228
R55151 a_33249_34067.n141 a_33249_34067.n139 1.27228
R55152 a_33249_34067.n129 a_33249_34067.n125 1.27228
R55153 a_33249_34067.n53 a_33249_34067.n28 1.27228
R55154 a_33249_34067.n31 a_33249_34067.n30 1.26756
R55155 a_33249_34067.n45 a_33249_34067.n44 1.26756
R55156 a_33249_34067.n133 a_33249_34067.n132 1.26756
R55157 a_33249_34067.n142 a_33249_34067.n141 1.26756
R55158 a_33249_34067.n101 a_33249_34067.n98 1.26344
R55159 a_33249_34067.n110 a_33249_34067.t15 1.2605
R55160 a_33249_34067.n110 a_33249_34067.t14 1.2605
R55161 a_33249_34067.n108 a_33249_34067.t12 1.2605
R55162 a_33249_34067.n108 a_33249_34067.t0 1.2605
R55163 a_33249_34067.n100 a_33249_34067.t6 1.2605
R55164 a_33249_34067.n100 a_33249_34067.t5 1.2605
R55165 a_33249_34067.n99 a_33249_34067.t17 1.2605
R55166 a_33249_34067.n99 a_33249_34067.t4 1.2605
R55167 a_33249_34067.n102 a_33249_34067.t8 1.2605
R55168 a_33249_34067.n102 a_33249_34067.t13 1.2605
R55169 a_33249_34067.n103 a_33249_34067.t16 1.2605
R55170 a_33249_34067.n103 a_33249_34067.t2 1.2605
R55171 a_33249_34067.n62 a_33249_34067.t106 1.2605
R55172 a_33249_34067.n62 a_33249_34067.t120 1.2605
R55173 a_33249_34067.n72 a_33249_34067.t118 1.2605
R55174 a_33249_34067.n72 a_33249_34067.t122 1.2605
R55175 a_33249_34067.n71 a_33249_34067.t123 1.2605
R55176 a_33249_34067.n71 a_33249_34067.t135 1.2605
R55177 a_33249_34067.n69 a_33249_34067.t110 1.2605
R55178 a_33249_34067.n69 a_33249_34067.t108 1.2605
R55179 a_33249_34067.n95 a_33249_34067.t107 1.2605
R55180 a_33249_34067.n95 a_33249_34067.t124 1.2605
R55181 a_33249_34067.n91 a_33249_34067.t112 1.2605
R55182 a_33249_34067.n91 a_33249_34067.t119 1.2605
R55183 a_33249_34067.n89 a_33249_34067.t127 1.2605
R55184 a_33249_34067.n89 a_33249_34067.t138 1.2605
R55185 a_33249_34067.n85 a_33249_34067.t137 1.2605
R55186 a_33249_34067.n85 a_33249_34067.t113 1.2605
R55187 a_33249_34067.n80 a_33249_34067.t139 1.2605
R55188 a_33249_34067.n80 a_33249_34067.t117 1.2605
R55189 a_33249_34067.n81 a_33249_34067.t132 1.2605
R55190 a_33249_34067.n81 a_33249_34067.t115 1.2605
R55191 a_33249_34067.n65 a_33249_34067.t128 1.2605
R55192 a_33249_34067.n65 a_33249_34067.t140 1.2605
R55193 a_33249_34067.n66 a_33249_34067.t121 1.2605
R55194 a_33249_34067.n66 a_33249_34067.t134 1.2605
R55195 a_33249_34067.n83 a_33249_34067.n79 1.25428
R55196 a_33249_34067.n112 a_33249_34067.n111 1.25428
R55197 a_33249_34067.n93 a_33249_34067.n92 1.24956
R55198 a_33249_34067.n74 a_33249_34067.n23 1.25162
R55199 a_33249_34067.n33 a_33249_34067.n32 0.796291
R55200 a_33249_34067.n49 a_33249_34067.n46 0.796291
R55201 a_33249_34067.n135 a_33249_34067.n134 0.796291
R55202 a_33249_34067.n146 a_33249_34067.n143 0.796291
R55203 a_33249_34067.n152 a_33249_34067.n151 0.780703
R55204 a_33249_34067.n122 a_33249_34067.n121 0.780703
R55205 a_33249_34067.n148 a_33249_34067.n54 0.780703
R55206 a_33249_34067.n130 a_33249_34067.n55 0.780703
R55207 a_33249_34067.n88 a_33249_34067.n87 0.769291
R55208 a_33249_34067.n96 a_33249_34067.n94 0.769291
R55209 a_33249_34067.n75 a_33249_34067.n70 0.767125
R55210 a_33249_34067.n73 a_33249_34067.n63 0.767125
R55211 a_33249_34067.n113 a_33249_34067.n107 0.639318
R55212 a_33249_34067.n122 a_33249_34067.n34 0.638405
R55213 a_33249_34067.n76 a_33249_34067.n61 0.638405
R55214 a_33249_34067.n97 a_33249_34067.n84 0.638405
R55215 a_33249_34067.n147 a_33249_34067.n130 0.638405
R55216 a_33249_34067.n151 a_33249_34067.n34 0.628372
R55217 a_33249_34067.n148 a_33249_34067.n147 0.628372
R55218 a_33249_34067.n107 a_33249_34067.n101 0.585196
R55219 a_33249_34067.n90 a_33249_34067.n88 0.485484
R55220 a_33249_34067.n40 a_33249_34067.n33 0.476484
R55221 a_33249_34067.n49 a_33249_34067.n48 0.476484
R55222 a_33249_34067.n137 a_33249_34067.n135 0.476484
R55223 a_33249_34067.n146 a_33249_34067.n145 0.476484
R55224 a_33249_34067.n75 a_33249_34067.n24 0.484998
R55225 a_33249_34067.n150 a_33249_34067.n6 0.478684
R55226 a_33249_34067.n149 a_33249_34067.n0 0.478684
R55227 a_33249_34067.n120 a_33249_34067.n16 0.478684
R55228 a_33249_34067.n119 a_33249_34067.n10 0.478684
R55229 a_33249_34067.n8 a_33249_34067.n9 1.27228
R55230 a_33249_34067.n7 a_33249_34067.n8 2.51878
R55231 a_33249_34067.n150 a_33249_34067.n7 0.794091
R55232 a_33249_34067.n5 a_33249_34067.n6 1.27228
R55233 a_33249_34067.n4 a_33249_34067.n5 2.60203
R55234 a_33249_34067.n3 a_33249_34067.n4 1.27228
R55235 a_33249_34067.n2 a_33249_34067.n3 1.27228
R55236 a_33249_34067.n1 a_33249_34067.n2 2.51878
R55237 a_33249_34067.n149 a_33249_34067.n1 0.794091
R55238 a_33249_34067.t70 a_33249_34067.n0 6.77266
R55239 a_33249_34067.n18 a_33249_34067.n19 1.27228
R55240 a_33249_34067.n17 a_33249_34067.n18 2.51878
R55241 a_33249_34067.n120 a_33249_34067.n17 0.794091
R55242 a_33249_34067.n15 a_33249_34067.n16 1.27228
R55243 a_33249_34067.n14 a_33249_34067.n15 2.60203
R55244 a_33249_34067.n13 a_33249_34067.n14 1.27228
R55245 a_33249_34067.n12 a_33249_34067.n13 1.27228
R55246 a_33249_34067.n11 a_33249_34067.n12 2.51878
R55247 a_33249_34067.n119 a_33249_34067.n11 0.794091
R55248 a_33249_34067.t60 a_33249_34067.n10 6.77266
R55249 a_33249_34067.n21 a_33249_34067.n22 3.15817
R55250 a_33249_34067.n20 a_33249_34067.n21 1.27188
R55251 a_33249_34067.n101 a_33249_34067.n20 1.73829
R55252 a_33249_34067.n70 a_33249_34067.n25 3.17898
R55253 a_33249_34067.n74 a_33249_34067.n24 3.19023
R55254 a_33249_34067.n73 a_33249_34067.n23 3.17898
R55255 a_65486_n35156.t8 a_65486_n35156.t3 12.7136
R55256 a_65486_n35156.t8 a_65486_n35156.t14 10.2828
R55257 a_65486_n35156.t8 a_65486_n35156.t6 10.2828
R55258 a_65486_n35156.t8 a_65486_n35156.t13 10.2828
R55259 a_65486_n35156.t8 a_65486_n35156.t4 10.2828
R55260 a_65486_n35156.t8 a_65486_n35156.t0 10.1333
R55261 a_65486_n35156.t8 a_65486_n35156.t21 10.1333
R55262 a_65486_n35156.t8 a_65486_n35156.t2 10.1333
R55263 a_65486_n35156.t8 a_65486_n35156.t22 10.1333
R55264 a_65486_n35156.t8 a_65486_n35156.t11 9.72545
R55265 a_65486_n35156.t8 a_65486_n35156.t20 9.57156
R55266 a_65486_n35156.t8 a_65486_n35156.t17 9.57156
R55267 a_65486_n35156.t8 a_65486_n35156.t19 9.57156
R55268 a_65486_n35156.t8 a_65486_n35156.t18 9.57156
R55269 a_65486_n35156.t8 a_65486_n35156.t16 9.57156
R55270 a_65486_n35156.t8 a_65486_n35156.t23 9.57156
R55271 a_65486_n35156.t8 a_65486_n35156.t15 9.57156
R55272 a_65486_n35156.t8 a_65486_n35156.t12 9.57156
R55273 a_65486_n35156.t11 a_65486_n35156.t10 8.02827
R55274 a_65486_n35156.t8 a_65486_n35156.t9 8.0259
R55275 a_65486_n35156.t8 a_65486_n35156.t5 7.90799
R55276 a_65486_n35156.t8 a_65486_n35156.t7 7.90799
R55277 a_65486_n35156.t1 a_65486_n35156.t8 7.41865
R55278 a_100820_n36322.n0 a_100820_n36322.t16 13.7934
R55279 a_100820_n36322.n2 a_100820_n36322.t1 10.7024
R55280 a_100820_n36322.n2 a_100820_n36322.t4 10.1668
R55281 a_100820_n36322.n2 a_100820_n36322.t7 9.64458
R55282 a_100820_n36322.n2 a_100820_n36322.t3 9.27635
R55283 a_100820_n36322.n2 a_100820_n36322.n0 8.75198
R55284 a_100820_n36322.n0 a_100820_n36322.t20 8.14051
R55285 a_100820_n36322.n0 a_100820_n36322.t18 8.14051
R55286 a_100820_n36322.n0 a_100820_n36322.t10 8.14051
R55287 a_100820_n36322.n0 a_100820_n36322.t11 8.14051
R55288 a_100820_n36322.n0 a_100820_n36322.t17 8.06917
R55289 a_100820_n36322.n0 a_100820_n36322.t15 8.06917
R55290 a_100820_n36322.n0 a_100820_n36322.t14 8.06917
R55291 a_100820_n36322.n0 a_100820_n36322.t9 8.06917
R55292 a_100820_n36322.n0 a_100820_n36322.t23 8.06917
R55293 a_100820_n36322.n0 a_100820_n36322.t19 8.06917
R55294 a_100820_n36322.n0 a_100820_n36322.t22 8.06917
R55295 a_100820_n36322.n1 a_100820_n36322.t6 7.94157
R55296 a_100820_n36322.t0 a_100820_n36322.n2 7.72643
R55297 a_100820_n36322.n1 a_100820_n36322.t5 7.22925
R55298 a_100820_n36322.n2 a_100820_n36322.t2 7.17912
R55299 a_100820_n36322.n0 a_100820_n36322.t8 8.33554
R55300 a_100820_n36322.t21 a_100820_n36322.n0 8.33554
R55301 a_100820_n36322.n0 a_100820_n36322.t12 8.33647
R55302 a_100820_n36322.t13 a_100820_n36322.n0 8.33647
R55303 a_100820_n36322.n2 a_100820_n36322.n1 7.46075
R55304 a_106676_n30339.n0 a_106676_n30339.t3 10.3838
R55305 a_106676_n30339.n0 a_106676_n30339.t1 10.3566
R55306 a_106676_n30339.n0 a_106676_n30339.t0 10.0407
R55307 a_106676_n30339.t2 a_106676_n30339.n0 9.57605
R55308 a_83153_11614.n2 a_83153_11614.t15 12.8637
R55309 a_83153_11614.n1 a_83153_11614.t6 10.7018
R55310 a_83153_11614.n1 a_83153_11614.t2 10.1659
R55311 a_83153_11614.n1 a_83153_11614.t1 9.64387
R55312 a_83153_11614.t4 a_83153_11614.n1 9.27665
R55313 a_83153_11614.n1 a_83153_11614.n2 8.75198
R55314 a_83153_11614.n2 a_83153_11614.t14 8.14051
R55315 a_83153_11614.n2 a_83153_11614.t10 8.14051
R55316 a_83153_11614.n2 a_83153_11614.t22 8.14051
R55317 a_83153_11614.n2 a_83153_11614.t16 8.14051
R55318 a_83153_11614.n2 a_83153_11614.t23 8.06917
R55319 a_83153_11614.n2 a_83153_11614.t20 8.06917
R55320 a_83153_11614.n2 a_83153_11614.t9 8.06917
R55321 a_83153_11614.n2 a_83153_11614.t12 8.06917
R55322 a_83153_11614.n2 a_83153_11614.t19 8.06917
R55323 a_83153_11614.n2 a_83153_11614.t11 8.06917
R55324 a_83153_11614.n2 a_83153_11614.t21 8.06917
R55325 a_83153_11614.n0 a_83153_11614.t3 7.94068
R55326 a_83153_11614.n1 a_83153_11614.t7 7.72524
R55327 a_83153_11614.n0 a_83153_11614.t0 7.22855
R55328 a_83153_11614.n1 a_83153_11614.t5 7.17942
R55329 a_83153_11614.t13 a_83153_11614.n2 8.33649
R55330 a_83153_11614.n2 a_83153_11614.t17 8.33649
R55331 a_83153_11614.t18 a_83153_11614.n2 8.33556
R55332 a_83153_11614.n2 a_83153_11614.t8 8.33556
R55333 a_83153_11614.n1 a_83153_11614.n0 7.46075
R55334 a_86903_n14095.t0 a_86903_n14095.t2 61.4377
R55335 a_86903_n14095.t0 a_86903_n14095.n0 13.0169
R55336 a_86903_n14095.n1 a_86903_n14095.n0 10.9309
R55337 a_86903_n14095.t0 a_86903_n14095.t1 8.5021
R55338 a_86903_n14095.n1 a_86903_n14095.t6 8.44198
R55339 a_86903_n14095.n1 a_86903_n14095.t8 8.44198
R55340 a_86903_n14095.n0 a_86903_n14095.t3 8.44198
R55341 a_86903_n14095.n0 a_86903_n14095.t7 8.44198
R55342 a_86903_n14095.n1 a_86903_n14095.t9 8.10567
R55343 a_86903_n14095.n0 a_86903_n14095.t10 9.26955
R55344 a_86903_n14095.n1 a_86903_n14095.t4 8.65823
R55345 a_86903_n14095.n0 a_86903_n14095.t5 8.77493
R55346 a_89715_n17715.t0 a_89715_n17715.t3 64.7456
R55347 a_89715_n17715.t3 a_89715_n17715.t1 12.9273
R55348 a_89715_n17715.t3 a_89715_n17715.t5 10.1307
R55349 a_89715_n17715.t3 a_89715_n17715.t4 8.54643
R55350 a_89715_n17715.t3 a_89715_n17715.t2 7.50895
R55351 a_112559_4481.n1 a_112559_4481.t4 10.2515
R55352 a_112559_4481.n1 a_112559_4481.t0 10.2515
R55353 a_112559_4481.n1 a_112559_4481.t12 10.2515
R55354 a_112559_4481.n1 a_112559_4481.t17 10.2515
R55355 a_112559_4481.n1 a_112559_4481.t2 10.096
R55356 a_112559_4481.n1 a_112559_4481.t22 10.0935
R55357 a_112559_4481.n1 a_112559_4481.t6 10.0859
R55358 a_112559_4481.n1 a_112559_4481.t15 10.0808
R55359 a_112559_4481.n1 a_112559_4481.t19 9.53981
R55360 a_112559_4481.n1 a_112559_4481.t16 9.53981
R55361 a_112559_4481.n1 a_112559_4481.t11 9.53981
R55362 a_112559_4481.n1 a_112559_4481.t13 9.53981
R55363 a_112559_4481.n1 a_112559_4481.t21 9.53744
R55364 a_112559_4481.n1 a_112559_4481.t20 9.53744
R55365 a_112559_4481.n1 a_112559_4481.t14 9.53744
R55366 a_112559_4481.n1 a_112559_4481.t18 9.53744
R55367 a_112559_4481.n1 a_112559_4481.n0 8.41434
R55368 a_112559_4481.n1 a_112559_4481.t5 8.14082
R55369 a_112559_4481.n0 a_112559_4481.t1 8.13828
R55370 a_112559_4481.t8 a_112559_4481.t9 7.96115
R55371 a_112559_4481.t9 a_112559_4481.t10 7.94694
R55372 a_112559_4481.t9 a_112559_4481.n1 7.50666
R55373 a_112559_4481.n0 a_112559_4481.t3 7.48586
R55374 a_112559_4481.n1 a_112559_4481.t7 7.48333
R55375 a_30152_n36322.n0 a_30152_n36322.t14 13.7934
R55376 a_30152_n36322.n2 a_30152_n36322.t7 10.7024
R55377 a_30152_n36322.n2 a_30152_n36322.t0 10.1668
R55378 a_30152_n36322.n2 a_30152_n36322.t2 9.64458
R55379 a_30152_n36322.n2 a_30152_n36322.t5 9.27635
R55380 a_30152_n36322.n2 a_30152_n36322.n0 8.75198
R55381 a_30152_n36322.n0 a_30152_n36322.t13 8.14051
R55382 a_30152_n36322.n0 a_30152_n36322.t11 8.14051
R55383 a_30152_n36322.n0 a_30152_n36322.t18 8.14051
R55384 a_30152_n36322.n0 a_30152_n36322.t21 8.14051
R55385 a_30152_n36322.n0 a_30152_n36322.t15 8.06917
R55386 a_30152_n36322.n0 a_30152_n36322.t20 8.06917
R55387 a_30152_n36322.n0 a_30152_n36322.t17 8.06917
R55388 a_30152_n36322.n0 a_30152_n36322.t23 8.06917
R55389 a_30152_n36322.n0 a_30152_n36322.t22 8.06917
R55390 a_30152_n36322.n0 a_30152_n36322.t8 8.06917
R55391 a_30152_n36322.n0 a_30152_n36322.t9 8.06917
R55392 a_30152_n36322.n1 a_30152_n36322.t3 7.94157
R55393 a_30152_n36322.n2 a_30152_n36322.t6 7.72643
R55394 a_30152_n36322.n1 a_30152_n36322.t1 7.22925
R55395 a_30152_n36322.t4 a_30152_n36322.n2 7.17912
R55396 a_30152_n36322.n0 a_30152_n36322.t12 8.33554
R55397 a_30152_n36322.t10 a_30152_n36322.n0 8.33554
R55398 a_30152_n36322.n0 a_30152_n36322.t16 8.33647
R55399 a_30152_n36322.t19 a_30152_n36322.n0 8.33647
R55400 a_30152_n36322.n2 a_30152_n36322.n1 7.46075
R55401 a_47819_n35156.t2 a_47819_n35156.t8 12.7136
R55402 a_47819_n35156.t2 a_47819_n35156.t13 10.2828
R55403 a_47819_n35156.t2 a_47819_n35156.t9 10.2828
R55404 a_47819_n35156.t2 a_47819_n35156.t12 10.2828
R55405 a_47819_n35156.t2 a_47819_n35156.t5 10.2828
R55406 a_47819_n35156.t2 a_47819_n35156.t3 10.1333
R55407 a_47819_n35156.t2 a_47819_n35156.t20 10.1333
R55408 a_47819_n35156.t2 a_47819_n35156.t7 10.1333
R55409 a_47819_n35156.t2 a_47819_n35156.t22 10.1333
R55410 a_47819_n35156.t2 a_47819_n35156.t11 9.72545
R55411 a_47819_n35156.t2 a_47819_n35156.t19 9.57156
R55412 a_47819_n35156.t2 a_47819_n35156.t16 9.57156
R55413 a_47819_n35156.t2 a_47819_n35156.t18 9.57156
R55414 a_47819_n35156.t2 a_47819_n35156.t17 9.57156
R55415 a_47819_n35156.t2 a_47819_n35156.t15 9.57156
R55416 a_47819_n35156.t2 a_47819_n35156.t21 9.57156
R55417 a_47819_n35156.t2 a_47819_n35156.t14 9.57156
R55418 a_47819_n35156.t2 a_47819_n35156.t23 9.57156
R55419 a_47819_n35156.t11 a_47819_n35156.t0 8.02827
R55420 a_47819_n35156.t2 a_47819_n35156.t1 8.0259
R55421 a_47819_n35156.t2 a_47819_n35156.t6 7.90799
R55422 a_47819_n35156.t2 a_47819_n35156.t10 7.90799
R55423 a_47819_n35156.t4 a_47819_n35156.t2 7.41865
R55424 a_51711_n12421.t0 a_51711_n12421.t1 78.206
R55425 a_51711_n12421.t0 a_51711_n12421.t2 24.9014
R55426 a_100820_n35156.t0 a_100820_n35156.t7 12.7136
R55427 a_100820_n35156.t0 a_100820_n35156.t21 10.2828
R55428 a_100820_n35156.t0 a_100820_n35156.t10 10.2828
R55429 a_100820_n35156.t0 a_100820_n35156.t20 10.2828
R55430 a_100820_n35156.t0 a_100820_n35156.t8 10.2828
R55431 a_100820_n35156.t0 a_100820_n35156.t4 10.1333
R55432 a_100820_n35156.t0 a_100820_n35156.t12 10.1333
R55433 a_100820_n35156.t0 a_100820_n35156.t6 10.1333
R55434 a_100820_n35156.t0 a_100820_n35156.t13 10.1333
R55435 a_100820_n35156.t0 a_100820_n35156.t2 9.72545
R55436 a_100820_n35156.t0 a_100820_n35156.t17 9.57156
R55437 a_100820_n35156.t0 a_100820_n35156.t14 9.57156
R55438 a_100820_n35156.t0 a_100820_n35156.t16 9.57156
R55439 a_100820_n35156.t0 a_100820_n35156.t15 9.57156
R55440 a_100820_n35156.t0 a_100820_n35156.t23 9.57156
R55441 a_100820_n35156.t0 a_100820_n35156.t18 9.57156
R55442 a_100820_n35156.t0 a_100820_n35156.t22 9.57156
R55443 a_100820_n35156.t0 a_100820_n35156.t19 9.57156
R55444 a_100820_n35156.t2 a_100820_n35156.t1 8.02827
R55445 a_100820_n35156.t0 a_100820_n35156.t3 8.0259
R55446 a_100820_n35156.t0 a_100820_n35156.t9 7.90799
R55447 a_100820_n35156.t0 a_100820_n35156.t11 7.90799
R55448 a_100820_n35156.t5 a_100820_n35156.t0 7.41865
R55449 a_77225_4481.n1 a_77225_4481.t4 10.2515
R55450 a_77225_4481.n1 a_77225_4481.t6 10.2515
R55451 a_77225_4481.n1 a_77225_4481.t13 10.2515
R55452 a_77225_4481.n1 a_77225_4481.t16 10.2515
R55453 a_77225_4481.n1 a_77225_4481.t0 10.096
R55454 a_77225_4481.n1 a_77225_4481.t19 10.0935
R55455 a_77225_4481.n1 a_77225_4481.t2 10.0859
R55456 a_77225_4481.n1 a_77225_4481.t11 10.0808
R55457 a_77225_4481.n1 a_77225_4481.t21 9.53981
R55458 a_77225_4481.n1 a_77225_4481.t20 9.53981
R55459 a_77225_4481.n1 a_77225_4481.t17 9.53981
R55460 a_77225_4481.n1 a_77225_4481.t18 9.53981
R55461 a_77225_4481.n1 a_77225_4481.t15 9.53744
R55462 a_77225_4481.n1 a_77225_4481.t14 9.53744
R55463 a_77225_4481.n1 a_77225_4481.t22 9.53744
R55464 a_77225_4481.n1 a_77225_4481.t12 9.53744
R55465 a_77225_4481.n1 a_77225_4481.n0 8.41434
R55466 a_77225_4481.n1 a_77225_4481.t5 8.14082
R55467 a_77225_4481.n0 a_77225_4481.t7 8.13828
R55468 a_77225_4481.t8 a_77225_4481.t10 7.96115
R55469 a_77225_4481.t8 a_77225_4481.t9 7.94694
R55470 a_77225_4481.t8 a_77225_4481.n1 7.50666
R55471 a_77225_4481.n0 a_77225_4481.t1 7.48586
R55472 a_77225_4481.n1 a_77225_4481.t3 7.48333
R55473 a_106830_10388.n6 a_106830_10388.n1 10.2377
R55474 a_106830_10388.n5 a_106830_10388.t1 10.2108
R55475 a_106830_10388.n5 a_106830_10388.t0 9.99909
R55476 a_106830_10388.t4 a_106830_10388.n6 9.80443
R55477 a_106830_10388.n6 a_106830_10388.t6 9.55135
R55478 a_106830_10388.n0 a_106830_10388.t18 8.17385
R55479 a_106830_10388.n3 a_106830_10388.t15 8.17299
R55480 a_106830_10388.n3 a_106830_10388.t17 8.17134
R55481 a_106830_10388.n0 a_106830_10388.t14 8.16754
R55482 a_106830_10388.n1 a_106830_10388.t11 8.10567
R55483 a_106830_10388.n1 a_106830_10388.t10 8.10567
R55484 a_106830_10388.n3 a_106830_10388.t23 8.10567
R55485 a_106830_10388.n3 a_106830_10388.t8 8.10567
R55486 a_106830_10388.n1 a_106830_10388.t9 8.10567
R55487 a_106830_10388.n1 a_106830_10388.t16 8.10567
R55488 a_106830_10388.n0 a_106830_10388.t13 8.10567
R55489 a_106830_10388.n0 a_106830_10388.t21 8.10567
R55490 a_106830_10388.n7 a_106830_10388.t3 7.74799
R55491 a_106830_10388.n4 a_106830_10388.t5 7.73052
R55492 a_106830_10388.n7 a_106830_10388.t2 7.46478
R55493 a_106830_10388.n4 a_106830_10388.t7 7.1311
R55494 a_106830_10388.n5 a_106830_10388.n7 2.2505
R55495 a_106830_10388.n6 a_106830_10388.n4 2.2505
R55496 a_106830_10388.n1 a_106830_10388.t19 8.35731
R55497 a_106830_10388.n0 a_106830_10388.t12 8.38107
R55498 a_106830_10388.n1 a_106830_10388.t20 8.37583
R55499 a_106830_10388.n1 a_106830_10388.n0 4.35656
R55500 a_106830_10388.n6 a_106830_10388.n5 2.96863
R55501 a_106830_10388.n2 a_106830_10388.n1 1.0882
R55502 a_106830_10388.n2 a_106830_10388.n3 1.08408
R55503 a_106830_10388.n2 a_106830_10388.t22 8.66753
R55504 a_106676_4481.n0 a_106676_4481.t3 10.6581
R55505 a_106676_4481.n0 a_106676_4481.t1 10.2356
R55506 a_106676_4481.t0 a_106676_4481.n0 9.5019
R55507 a_106676_4481.n0 a_106676_4481.t2 9.34796
R55508 a_36032_n35156.t0 a_36032_n35156.n3 96.9245
R55509 a_36032_n35156.n1 a_36032_n35156.n0 10.9327
R55510 a_36032_n35156.n0 a_36032_n35156.t8 8.44198
R55511 a_36032_n35156.n0 a_36032_n35156.t10 8.44198
R55512 a_36032_n35156.n1 a_36032_n35156.t7 8.44198
R55513 a_36032_n35156.n1 a_36032_n35156.t9 8.44198
R55514 a_36032_n35156.n0 a_36032_n35156.t5 9.26917
R55515 a_36032_n35156.n1 a_36032_n35156.t6 8.10567
R55516 a_36032_n35156.n3 a_36032_n35156.t1 6.51122
R55517 a_36032_n35156.n3 a_36032_n35156.n0 6.50622
R55518 a_36032_n35156.t1 a_36032_n35156.t2 6.36267
R55519 a_36032_n35156.t1 a_36032_n35156.n2 4.84877
R55520 a_36032_n35156.n2 a_36032_n35156.t4 3.65383
R55521 a_36032_n35156.n1 a_36032_n35156.t12 8.65827
R55522 a_36032_n35156.n2 a_36032_n35156.t3 3.57094
R55523 a_36032_n35156.n0 a_36032_n35156.t11 8.77499
R55524 a_30152_n35156.t0 a_30152_n35156.t11 12.7136
R55525 a_30152_n35156.t0 a_30152_n35156.t18 10.2828
R55526 a_30152_n35156.t0 a_30152_n35156.t4 10.2828
R55527 a_30152_n35156.t0 a_30152_n35156.t17 10.2828
R55528 a_30152_n35156.t0 a_30152_n35156.t6 10.2828
R55529 a_30152_n35156.t0 a_30152_n35156.t8 10.1333
R55530 a_30152_n35156.t0 a_30152_n35156.t19 10.1333
R55531 a_30152_n35156.t0 a_30152_n35156.t10 10.1333
R55532 a_30152_n35156.t0 a_30152_n35156.t20 10.1333
R55533 a_30152_n35156.t0 a_30152_n35156.t3 9.72545
R55534 a_30152_n35156.t0 a_30152_n35156.t16 9.57156
R55535 a_30152_n35156.t0 a_30152_n35156.t22 9.57156
R55536 a_30152_n35156.t0 a_30152_n35156.t15 9.57156
R55537 a_30152_n35156.t0 a_30152_n35156.t12 9.57156
R55538 a_30152_n35156.t0 a_30152_n35156.t14 9.57156
R55539 a_30152_n35156.t0 a_30152_n35156.t21 9.57156
R55540 a_30152_n35156.t0 a_30152_n35156.t13 9.57156
R55541 a_30152_n35156.t0 a_30152_n35156.t23 9.57156
R55542 a_30152_n35156.t3 a_30152_n35156.t1 8.02827
R55543 a_30152_n35156.t0 a_30152_n35156.t2 8.0259
R55544 a_30152_n35156.t0 a_30152_n35156.t7 7.90799
R55545 a_30152_n35156.t5 a_30152_n35156.t0 7.90799
R55546 a_30152_n35156.t0 a_30152_n35156.t9 7.41865
R55547 a_89163_10388.n6 a_89163_10388.n1 10.2377
R55548 a_89163_10388.n5 a_89163_10388.t3 10.2108
R55549 a_89163_10388.n5 a_89163_10388.t2 9.99909
R55550 a_89163_10388.n6 a_89163_10388.t6 9.80443
R55551 a_89163_10388.t4 a_89163_10388.n6 9.55135
R55552 a_89163_10388.n0 a_89163_10388.t17 8.17385
R55553 a_89163_10388.n3 a_89163_10388.t9 8.17299
R55554 a_89163_10388.n3 a_89163_10388.t11 8.17134
R55555 a_89163_10388.n0 a_89163_10388.t8 8.16754
R55556 a_89163_10388.n1 a_89163_10388.t16 8.10567
R55557 a_89163_10388.n1 a_89163_10388.t14 8.10567
R55558 a_89163_10388.n3 a_89163_10388.t20 8.10567
R55559 a_89163_10388.n3 a_89163_10388.t21 8.10567
R55560 a_89163_10388.n1 a_89163_10388.t13 8.10567
R55561 a_89163_10388.n1 a_89163_10388.t18 8.10567
R55562 a_89163_10388.n0 a_89163_10388.t12 8.10567
R55563 a_89163_10388.n0 a_89163_10388.t19 8.10567
R55564 a_89163_10388.n7 a_89163_10388.t0 7.74799
R55565 a_89163_10388.n4 a_89163_10388.t7 7.73052
R55566 a_89163_10388.n7 a_89163_10388.t1 7.46478
R55567 a_89163_10388.n4 a_89163_10388.t5 7.1311
R55568 a_89163_10388.n5 a_89163_10388.n7 2.2505
R55569 a_89163_10388.n6 a_89163_10388.n4 2.2505
R55570 a_89163_10388.n1 a_89163_10388.t22 8.35731
R55571 a_89163_10388.n0 a_89163_10388.t15 8.38107
R55572 a_89163_10388.n1 a_89163_10388.t23 8.37583
R55573 a_89163_10388.n1 a_89163_10388.n0 4.35656
R55574 a_89163_10388.n6 a_89163_10388.n5 2.96863
R55575 a_89163_10388.n2 a_89163_10388.n1 1.0882
R55576 a_89163_10388.n2 a_89163_10388.n3 1.08408
R55577 a_89163_10388.n2 a_89163_10388.t10 8.66753
R55578 a_89033_13546.n1 a_89033_13546.n0 26.5215
R55579 a_89033_13546.n0 a_89033_13546.t3 11.5094
R55580 a_89033_13546.n1 a_89033_13546.t1 10.937
R55581 a_89033_13546.t0 a_89033_13546.n1 9.33982
R55582 a_89033_13546.n0 a_89033_13546.t2 9.24966
R55583 a_65486_10448.n0 a_65486_10448.t4 10.2828
R55584 a_65486_10448.t10 a_65486_10448.t2 10.2828
R55585 a_65486_10448.n0 a_65486_10448.t19 10.2828
R55586 a_65486_10448.n0 a_65486_10448.t16 10.2828
R55587 a_65486_10448.n0 a_65486_10448.t17 10.1333
R55588 a_65486_10448.t10 a_65486_10448.t18 10.1333
R55589 a_65486_10448.n0 a_65486_10448.t0 10.1333
R55590 a_65486_10448.n0 a_65486_10448.t6 10.1333
R55591 a_65486_10448.n0 a_65486_10448.t13 9.57156
R55592 a_65486_10448.n0 a_65486_10448.t11 9.57156
R55593 a_65486_10448.t10 a_65486_10448.t12 9.57156
R55594 a_65486_10448.n0 a_65486_10448.t15 9.57156
R55595 a_65486_10448.n0 a_65486_10448.t22 9.57156
R55596 a_65486_10448.n0 a_65486_10448.t20 9.57156
R55597 a_65486_10448.t10 a_65486_10448.t21 9.57156
R55598 a_65486_10448.n0 a_65486_10448.t14 9.57156
R55599 a_65486_10448.t10 a_65486_10448.n1 8.94763
R55600 a_65486_10448.t10 a_65486_10448.t9 8.02945
R55601 a_65486_10448.t10 a_65486_10448.t8 8.02708
R55602 a_65486_10448.t10 a_65486_10448.t5 7.90829
R55603 a_65486_10448.n1 a_65486_10448.t3 7.90829
R55604 a_65486_10448.n1 a_65486_10448.t7 7.41776
R55605 a_65486_10448.t1 a_65486_10448.t10 7.41776
R55606 a_65486_10448.t10 a_65486_10448.n0 7.31642
R55607 a_36032_11614.t0 a_36032_11614.n2 74.3465
R55608 a_36032_11614.n1 a_36032_11614.n0 10.9309
R55609 a_36032_11614.t1 a_36032_11614.t2 8.5021
R55610 a_36032_11614.n1 a_36032_11614.t9 8.44198
R55611 a_36032_11614.n1 a_36032_11614.t5 8.44198
R55612 a_36032_11614.n0 a_36032_11614.t6 8.44198
R55613 a_36032_11614.n0 a_36032_11614.t10 8.44198
R55614 a_36032_11614.n1 a_36032_11614.t3 8.10567
R55615 a_36032_11614.n0 a_36032_11614.t4 9.26955
R55616 a_36032_11614.n2 a_36032_11614.t1 6.51122
R55617 a_36032_11614.n2 a_36032_11614.n0 6.50622
R55618 a_36032_11614.n1 a_36032_11614.t7 8.65823
R55619 a_36032_11614.n0 a_36032_11614.t8 8.77493
R55620 a_43010_10448.t0 a_43010_10448.t3 76.8811
R55621 a_43010_10448.t0 a_43010_10448.t1 13.8923
R55622 a_43010_10448.t0 a_43010_10448.t4 10.1307
R55623 a_43010_10448.t0 a_43010_10448.t2 8.54643
R55624 a_81205_n14095.t0 a_81205_n14095.n2 45.7073
R55625 a_81205_n14095.n1 a_81205_n14095.n0 10.9309
R55626 a_81205_n14095.t1 a_81205_n14095.t2 8.5021
R55627 a_81205_n14095.n1 a_81205_n14095.t3 8.44198
R55628 a_81205_n14095.n1 a_81205_n14095.t7 8.44198
R55629 a_81205_n14095.n0 a_81205_n14095.t8 8.44198
R55630 a_81205_n14095.n0 a_81205_n14095.t4 8.44198
R55631 a_81205_n14095.n1 a_81205_n14095.t5 8.10567
R55632 a_81205_n14095.n0 a_81205_n14095.t6 9.26955
R55633 a_81205_n14095.n2 a_81205_n14095.t1 6.51122
R55634 a_81205_n14095.n2 a_81205_n14095.n0 6.50622
R55635 a_81205_n14095.n1 a_81205_n14095.t9 8.65823
R55636 a_81205_n14095.n0 a_81205_n14095.t10 8.77493
R55637 a_89163_n36382.n5 a_89163_n36382.n1 10.2377
R55638 a_89163_n36382.n4 a_89163_n36382.t2 10.2105
R55639 a_89163_n36382.n4 a_89163_n36382.t1 9.99998
R55640 a_89163_n36382.n5 a_89163_n36382.t7 9.80532
R55641 a_89163_n36382.n5 a_89163_n36382.t5 9.55206
R55642 a_89163_n36382.n0 a_89163_n36382.t12 8.17385
R55643 a_89163_n36382.n3 a_89163_n36382.t10 8.17299
R55644 a_89163_n36382.n3 a_89163_n36382.t13 8.17134
R55645 a_89163_n36382.n0 a_89163_n36382.t11 8.16754
R55646 a_89163_n36382.n1 a_89163_n36382.t14 8.10567
R55647 a_89163_n36382.n1 a_89163_n36382.t19 8.10567
R55648 a_89163_n36382.n3 a_89163_n36382.t9 8.10567
R55649 a_89163_n36382.n3 a_89163_n36382.t22 8.10567
R55650 a_89163_n36382.n1 a_89163_n36382.t16 8.10567
R55651 a_89163_n36382.n1 a_89163_n36382.t18 8.10567
R55652 a_89163_n36382.n0 a_89163_n36382.t8 8.10567
R55653 a_89163_n36382.n0 a_89163_n36382.t23 8.10567
R55654 a_89163_n36382.n6 a_89163_n36382.t0 7.74888
R55655 a_89163_n36382.n7 a_89163_n36382.t6 7.73141
R55656 a_89163_n36382.n6 a_89163_n36382.t3 7.46359
R55657 a_89163_n36382.t4 a_89163_n36382.n7 7.13081
R55658 a_89163_n36382.n4 a_89163_n36382.n6 2.2505
R55659 a_89163_n36382.n7 a_89163_n36382.n5 2.2505
R55660 a_89163_n36382.t17 a_89163_n36382.n1 8.35729
R55661 a_89163_n36382.n1 a_89163_n36382.t15 8.37586
R55662 a_89163_n36382.n0 a_89163_n36382.t20 8.38104
R55663 a_89163_n36382.n1 a_89163_n36382.n0 4.35658
R55664 a_89163_n36382.n5 a_89163_n36382.n4 2.96863
R55665 a_89163_n36382.n2 a_89163_n36382.n1 1.08819
R55666 a_89163_n36382.n2 a_89163_n36382.n3 1.08408
R55667 a_89163_n36382.n2 a_89163_n36382.t21 8.6675
R55668 a_106809_n5150.t1 a_106809_n5150.t2 42.6546
R55669 a_106809_n5150.t1 a_106809_n5150.t3 9.77323
R55670 a_106809_n5150.t0 a_106809_n5150.t1 8.17727
R55671 a_41891_n29181.n0 a_41891_n29181.t14 10.2515
R55672 a_41891_n29181.n1 a_41891_n29181.t7 10.2515
R55673 a_41891_n29181.n0 a_41891_n29181.t18 10.2515
R55674 a_41891_n29181.n0 a_41891_n29181.t5 10.2515
R55675 a_41891_n29181.n0 a_41891_n29181.t9 10.096
R55676 a_41891_n29181.n1 a_41891_n29181.t19 10.0935
R55677 a_41891_n29181.n0 a_41891_n29181.t3 10.0859
R55678 a_41891_n29181.n0 a_41891_n29181.t12 10.0808
R55679 a_41891_n29181.n0 a_41891_n29181.t11 9.53981
R55680 a_41891_n29181.n1 a_41891_n29181.t22 9.53981
R55681 a_41891_n29181.n0 a_41891_n29181.t16 9.53981
R55682 a_41891_n29181.n0 a_41891_n29181.t17 9.53981
R55683 a_41891_n29181.n0 a_41891_n29181.t21 9.53744
R55684 a_41891_n29181.n1 a_41891_n29181.t20 9.53744
R55685 a_41891_n29181.n0 a_41891_n29181.t13 9.53744
R55686 a_41891_n29181.n0 a_41891_n29181.t15 9.53744
R55687 a_41891_n29181.n1 a_41891_n29181.n0 9.16839
R55688 a_41891_n29181.n1 a_41891_n29181.t6 8.14051
R55689 a_41891_n29181.n1 a_41891_n29181.t8 8.13798
R55690 a_41891_n29181.t0 a_41891_n29181.t1 7.95997
R55691 a_41891_n29181.t0 a_41891_n29181.t2 7.94576
R55692 a_41891_n29181.t0 a_41891_n29181.n1 7.50666
R55693 a_41891_n29181.n1 a_41891_n29181.t10 7.48675
R55694 a_41891_n29181.n1 a_41891_n29181.t4 7.48422
R55695 a_89009_n27257.n0 a_89009_n27257.t1 10.6581
R55696 a_89009_n27257.n0 a_89009_n27257.t3 10.2358
R55697 a_89009_n27257.t2 a_89009_n27257.n0 9.50202
R55698 a_89009_n27257.n0 a_89009_n27257.t0 9.34796
R55699 a_71496_n36382.n5 a_71496_n36382.n1 10.2377
R55700 a_71496_n36382.n4 a_71496_n36382.t3 10.2105
R55701 a_71496_n36382.n4 a_71496_n36382.t4 9.99998
R55702 a_71496_n36382.n5 a_71496_n36382.t7 9.80532
R55703 a_71496_n36382.n5 a_71496_n36382.t1 9.55206
R55704 a_71496_n36382.n0 a_71496_n36382.t10 8.17385
R55705 a_71496_n36382.n3 a_71496_n36382.t18 8.17299
R55706 a_71496_n36382.n3 a_71496_n36382.t11 8.17134
R55707 a_71496_n36382.n0 a_71496_n36382.t23 8.16754
R55708 a_71496_n36382.n1 a_71496_n36382.t16 8.10567
R55709 a_71496_n36382.n1 a_71496_n36382.t20 8.10567
R55710 a_71496_n36382.n3 a_71496_n36382.t15 8.10567
R55711 a_71496_n36382.n3 a_71496_n36382.t22 8.10567
R55712 a_71496_n36382.n1 a_71496_n36382.t17 8.10567
R55713 a_71496_n36382.n1 a_71496_n36382.t19 8.10567
R55714 a_71496_n36382.n0 a_71496_n36382.t14 8.10567
R55715 a_71496_n36382.n0 a_71496_n36382.t9 8.10567
R55716 a_71496_n36382.n6 a_71496_n36382.t2 7.74888
R55717 a_71496_n36382.n7 a_71496_n36382.t6 7.73141
R55718 a_71496_n36382.n6 a_71496_n36382.t5 7.46359
R55719 a_71496_n36382.t0 a_71496_n36382.n7 7.13081
R55720 a_71496_n36382.n4 a_71496_n36382.n6 2.2505
R55721 a_71496_n36382.n7 a_71496_n36382.n5 2.2505
R55722 a_71496_n36382.t8 a_71496_n36382.n1 8.35729
R55723 a_71496_n36382.n1 a_71496_n36382.t21 8.37586
R55724 a_71496_n36382.n0 a_71496_n36382.t12 8.38104
R55725 a_71496_n36382.n1 a_71496_n36382.n0 4.35658
R55726 a_71496_n36382.n5 a_71496_n36382.n4 2.96863
R55727 a_71496_n36382.n2 a_71496_n36382.n1 1.08819
R55728 a_71496_n36382.n2 a_71496_n36382.n3 1.08408
R55729 a_71496_n36382.n2 a_71496_n36382.t13 8.6675
R55730 a_53699_n36322.n1 a_53699_n36322.n0 26.5254
R55731 a_53699_n36322.t0 a_53699_n36322.n1 11.5094
R55732 a_53699_n36322.n0 a_53699_n36322.t3 10.937
R55733 a_53699_n36322.n0 a_53699_n36322.t2 9.33982
R55734 a_53699_n36322.n1 a_53699_n36322.t1 9.24966
R55735 a_44363_n16007.t0 a_44363_n16007.t2 56.3087
R55736 a_44363_n16007.t2 a_44363_n16007.t1 18.4133
R55737 a_71366_n35156.t0 a_71366_n35156.n3 69.4088
R55738 a_71366_n35156.n1 a_71366_n35156.n0 10.9327
R55739 a_71366_n35156.n0 a_71366_n35156.t9 8.44198
R55740 a_71366_n35156.n0 a_71366_n35156.t11 8.44198
R55741 a_71366_n35156.n1 a_71366_n35156.t8 8.44198
R55742 a_71366_n35156.n1 a_71366_n35156.t10 8.44198
R55743 a_71366_n35156.n0 a_71366_n35156.t12 9.26917
R55744 a_71366_n35156.n1 a_71366_n35156.t5 8.10567
R55745 a_71366_n35156.n3 a_71366_n35156.t3 6.51122
R55746 a_71366_n35156.n3 a_71366_n35156.n0 6.50622
R55747 a_71366_n35156.t3 a_71366_n35156.t2 6.36267
R55748 a_71366_n35156.t3 a_71366_n35156.n2 4.84877
R55749 a_71366_n35156.n2 a_71366_n35156.t4 3.65383
R55750 a_71366_n35156.n1 a_71366_n35156.t7 8.65827
R55751 a_71366_n35156.n2 a_71366_n35156.t1 3.57094
R55752 a_71366_n35156.n0 a_71366_n35156.t6 8.77499
R55753 a_78344_n36322.t0 a_78344_n36322.t2 67.5623
R55754 a_78344_n36322.t2 a_78344_n36322.t1 9.77323
R55755 a_78344_n36322.t2 a_78344_n36322.t3 8.17727
R55756 a_39179_n19595.t0 a_39179_n19595.t1 34.4821
R55757 a_39179_n19595.t0 a_39179_n19595.t2 24.9025
R55758 a_59558_4481.n1 a_59558_4481.t4 10.2515
R55759 a_59558_4481.n1 a_59558_4481.t6 10.2515
R55760 a_59558_4481.n1 a_59558_4481.t14 10.2515
R55761 a_59558_4481.n1 a_59558_4481.t19 10.2515
R55762 a_59558_4481.n1 a_59558_4481.t0 10.096
R55763 a_59558_4481.n1 a_59558_4481.t13 10.0935
R55764 a_59558_4481.n1 a_59558_4481.t2 10.0859
R55765 a_59558_4481.n1 a_59558_4481.t18 10.0808
R55766 a_59558_4481.n1 a_59558_4481.t21 9.53981
R55767 a_59558_4481.n1 a_59558_4481.t17 9.53981
R55768 a_59558_4481.n1 a_59558_4481.t12 9.53981
R55769 a_59558_4481.n1 a_59558_4481.t15 9.53981
R55770 a_59558_4481.n1 a_59558_4481.t11 9.53744
R55771 a_59558_4481.n1 a_59558_4481.t22 9.53744
R55772 a_59558_4481.n1 a_59558_4481.t16 9.53744
R55773 a_59558_4481.n1 a_59558_4481.t20 9.53744
R55774 a_59558_4481.n1 a_59558_4481.n0 8.41434
R55775 a_59558_4481.n1 a_59558_4481.t5 8.14082
R55776 a_59558_4481.n0 a_59558_4481.t7 8.13828
R55777 a_59558_4481.t8 a_59558_4481.t10 7.96115
R55778 a_59558_4481.t10 a_59558_4481.t9 7.94694
R55779 a_59558_4481.t10 a_59558_4481.n1 7.50666
R55780 a_59558_4481.n0 a_59558_4481.t1 7.48586
R55781 a_59558_4481.n1 a_59558_4481.t3 7.48333
R55782 a_53699_n35156.n1 a_53699_n35156.t2 80.9771
R55783 a_53699_n35156.n1 a_53699_n35156.t0 11.3595
R55784 a_53699_n35156.n2 a_53699_n35156.n0 10.9327
R55785 a_53699_n35156.n0 a_53699_n35156.t10 8.44198
R55786 a_53699_n35156.n0 a_53699_n35156.t6 8.44198
R55787 a_53699_n35156.n2 a_53699_n35156.t9 8.44198
R55788 a_53699_n35156.n2 a_53699_n35156.t5 8.44198
R55789 a_53699_n35156.n0 a_53699_n35156.t3 9.26917
R55790 a_53699_n35156.n2 a_53699_n35156.t4 8.10567
R55791 a_53699_n35156.n1 a_53699_n35156.n0 6.50622
R55792 a_53699_n35156.t0 a_53699_n35156.t1 3.65383
R55793 a_53699_n35156.n2 a_53699_n35156.t8 8.65827
R55794 a_53699_n35156.n0 a_53699_n35156.t7 8.77499
R55795 a_83325_n29313.t0 a_83325_n29313.t1 23.2303
R55796 a_83325_n29313.t0 a_83325_n29313.t2 21.6695
R55797 a_94892_n29181.n0 a_94892_n29181.t18 10.2515
R55798 a_94892_n29181.n1 a_94892_n29181.t5 10.2515
R55799 a_94892_n29181.n0 a_94892_n29181.t22 10.2515
R55800 a_94892_n29181.n0 a_94892_n29181.t3 10.2515
R55801 a_94892_n29181.n0 a_94892_n29181.t9 10.096
R55802 a_94892_n29181.n1 a_94892_n29181.t11 10.0935
R55803 a_94892_n29181.n0 a_94892_n29181.t7 10.0859
R55804 a_94892_n29181.n0 a_94892_n29181.t16 10.0808
R55805 a_94892_n29181.n0 a_94892_n29181.t15 9.53981
R55806 a_94892_n29181.n1 a_94892_n29181.t14 9.53981
R55807 a_94892_n29181.n0 a_94892_n29181.t20 9.53981
R55808 a_94892_n29181.n0 a_94892_n29181.t21 9.53981
R55809 a_94892_n29181.n0 a_94892_n29181.t13 9.53744
R55810 a_94892_n29181.n1 a_94892_n29181.t12 9.53744
R55811 a_94892_n29181.n0 a_94892_n29181.t17 9.53744
R55812 a_94892_n29181.n0 a_94892_n29181.t19 9.53744
R55813 a_94892_n29181.n1 a_94892_n29181.n0 9.16839
R55814 a_94892_n29181.n1 a_94892_n29181.t4 8.14051
R55815 a_94892_n29181.n1 a_94892_n29181.t6 8.13798
R55816 a_94892_n29181.t1 a_94892_n29181.t2 7.95997
R55817 a_94892_n29181.t0 a_94892_n29181.t1 7.94576
R55818 a_94892_n29181.t1 a_94892_n29181.n1 7.50666
R55819 a_94892_n29181.n1 a_94892_n29181.t10 7.48675
R55820 a_94892_n29181.n1 a_94892_n29181.t8 7.48422
R55821 I1U I1U.t1 3.63879
R55822 I1U.n0 I1U.t5 2.56243
R55823 I1U.n0 I1U.t4 2.32184
R55824 I1U.n1 I1U.t2 2.32184
R55825 I1U.n2 I1U.t3 2.32184
R55826 I1U.n3 I1U.t6 2.32184
R55827 I1U.n4 I1U.t0 1.34815
R55828 I1U.n4 I1U.n3 1.20346
R55829 I1U I1U.n4 1.12236
R55830 I1U.n1 I1U.n0 0.242306
R55831 I1U.n3 I1U.n2 0.241697
R55832 I1U.n2 I1U.n1 0.241089
R55833 a_77225_n29181.n0 a_77225_n29181.t15 10.2515
R55834 a_77225_n29181.n1 a_77225_n29181.t7 10.2515
R55835 a_77225_n29181.n0 a_77225_n29181.t19 10.2515
R55836 a_77225_n29181.n0 a_77225_n29181.t5 10.2515
R55837 a_77225_n29181.n0 a_77225_n29181.t3 10.096
R55838 a_77225_n29181.n1 a_77225_n29181.t13 10.0935
R55839 a_77225_n29181.n0 a_77225_n29181.t9 10.0859
R55840 a_77225_n29181.n0 a_77225_n29181.t18 10.0808
R55841 a_77225_n29181.n0 a_77225_n29181.t16 9.53981
R55842 a_77225_n29181.n1 a_77225_n29181.t14 9.53981
R55843 a_77225_n29181.n0 a_77225_n29181.t21 9.53981
R55844 a_77225_n29181.n0 a_77225_n29181.t22 9.53981
R55845 a_77225_n29181.n0 a_77225_n29181.t20 9.53744
R55846 a_77225_n29181.n1 a_77225_n29181.t17 9.53744
R55847 a_77225_n29181.n0 a_77225_n29181.t11 9.53744
R55848 a_77225_n29181.n0 a_77225_n29181.t12 9.53744
R55849 a_77225_n29181.n1 a_77225_n29181.n0 9.16839
R55850 a_77225_n29181.n1 a_77225_n29181.t6 8.14051
R55851 a_77225_n29181.n1 a_77225_n29181.t8 8.13798
R55852 a_77225_n29181.t2 a_77225_n29181.t1 7.95997
R55853 a_77225_n29181.t0 a_77225_n29181.t2 7.94576
R55854 a_77225_n29181.t2 a_77225_n29181.n1 7.50666
R55855 a_77225_n29181.n1 a_77225_n29181.t4 7.48675
R55856 a_77225_n29181.n1 a_77225_n29181.t10 7.48422
R55857 a_64243_n1756.t1 a_64243_n1756.t2 24.9014
R55858 a_64243_n1756.t0 a_64243_n1756.t1 23.8039
R55859 a_63161_n5344.t0 a_63161_n5344.t1 30.6913
R55860 a_63161_n5344.t1 a_63161_n5344.t2 15.0742
R55861 a_30152_11614.n2 a_30152_11614.t22 12.8637
R55862 a_30152_11614.n1 a_30152_11614.t7 10.7018
R55863 a_30152_11614.n1 a_30152_11614.t3 10.1659
R55864 a_30152_11614.n1 a_30152_11614.t1 9.64387
R55865 a_30152_11614.n1 a_30152_11614.t6 9.27665
R55866 a_30152_11614.n1 a_30152_11614.n2 8.75198
R55867 a_30152_11614.n2 a_30152_11614.t19 8.14051
R55868 a_30152_11614.n2 a_30152_11614.t15 8.14051
R55869 a_30152_11614.n2 a_30152_11614.t12 8.14051
R55870 a_30152_11614.n2 a_30152_11614.t23 8.14051
R55871 a_30152_11614.n2 a_30152_11614.t16 8.06917
R55872 a_30152_11614.n2 a_30152_11614.t13 8.06917
R55873 a_30152_11614.n2 a_30152_11614.t14 8.06917
R55874 a_30152_11614.n2 a_30152_11614.t18 8.06917
R55875 a_30152_11614.n2 a_30152_11614.t10 8.06917
R55876 a_30152_11614.n2 a_30152_11614.t20 8.06917
R55877 a_30152_11614.n2 a_30152_11614.t11 8.06917
R55878 a_30152_11614.n0 a_30152_11614.t2 7.94068
R55879 a_30152_11614.n1 a_30152_11614.t5 7.72524
R55880 a_30152_11614.n0 a_30152_11614.t0 7.22855
R55881 a_30152_11614.t4 a_30152_11614.n1 7.17942
R55882 a_30152_11614.t21 a_30152_11614.n2 8.33649
R55883 a_30152_11614.n2 a_30152_11614.t8 8.33649
R55884 a_30152_11614.t9 a_30152_11614.n2 8.33556
R55885 a_30152_11614.n2 a_30152_11614.t17 8.33556
R55886 a_30152_11614.n1 a_30152_11614.n0 7.46075
R55887 a_36008_4481.n0 a_36008_4481.t1 10.6581
R55888 a_36008_4481.t2 a_36008_4481.n0 10.2346
R55889 a_36008_4481.n0 a_36008_4481.t3 9.5029
R55890 a_36008_4481.n0 a_36008_4481.t0 9.34796
R55891 a_96011_n36322.t1 a_96011_n36322.t3 39.014
R55892 a_96011_n36322.t1 a_96011_n36322.t0 12.0003
R55893 a_96011_n36322.t1 a_96011_n36322.t2 8.17727
R55894 a_89033_n35156.t0 a_89033_n35156.n3 36.8446
R55895 a_89033_n35156.n1 a_89033_n35156.n0 10.9327
R55896 a_89033_n35156.n0 a_89033_n35156.t6 8.44198
R55897 a_89033_n35156.n0 a_89033_n35156.t8 8.44198
R55898 a_89033_n35156.n1 a_89033_n35156.t5 8.44198
R55899 a_89033_n35156.n1 a_89033_n35156.t7 8.44198
R55900 a_89033_n35156.n0 a_89033_n35156.t11 9.26917
R55901 a_89033_n35156.n1 a_89033_n35156.t12 8.10567
R55902 a_89033_n35156.n3 a_89033_n35156.t3 6.51122
R55903 a_89033_n35156.n3 a_89033_n35156.n0 6.50622
R55904 a_89033_n35156.t3 a_89033_n35156.t4 6.36267
R55905 a_89033_n35156.t3 a_89033_n35156.n2 4.84877
R55906 a_89033_n35156.n2 a_89033_n35156.t1 3.65383
R55907 a_89033_n35156.n1 a_89033_n35156.t10 8.65827
R55908 a_89033_n35156.n2 a_89033_n35156.t2 3.57094
R55909 a_89033_n35156.n0 a_89033_n35156.t9 8.77499
R55910 a_83153_n35156.n0 a_83153_n35156.t20 10.2828
R55911 a_83153_n35156.t8 a_83153_n35156.t4 10.2828
R55912 a_83153_n35156.n0 a_83153_n35156.t19 10.2828
R55913 a_83153_n35156.n0 a_83153_n35156.t0 10.2828
R55914 a_83153_n35156.n0 a_83153_n35156.t6 10.1333
R55915 a_83153_n35156.t8 a_83153_n35156.t21 10.1333
R55916 a_83153_n35156.n0 a_83153_n35156.t2 10.1333
R55917 a_83153_n35156.n0 a_83153_n35156.t22 10.1333
R55918 a_83153_n35156.n0 a_83153_n35156.t18 9.57156
R55919 a_83153_n35156.t8 a_83153_n35156.t12 9.57156
R55920 a_83153_n35156.n0 a_83153_n35156.t17 9.57156
R55921 a_83153_n35156.n0 a_83153_n35156.t14 9.57156
R55922 a_83153_n35156.n0 a_83153_n35156.t16 9.57156
R55923 a_83153_n35156.t8 a_83153_n35156.t11 9.57156
R55924 a_83153_n35156.n0 a_83153_n35156.t15 9.57156
R55925 a_83153_n35156.n0 a_83153_n35156.t13 9.57156
R55926 a_83153_n35156.t8 a_83153_n35156.n1 8.94763
R55927 a_83153_n35156.t8 a_83153_n35156.t9 8.02827
R55928 a_83153_n35156.t8 a_83153_n35156.t10 8.0259
R55929 a_83153_n35156.n1 a_83153_n35156.t5 7.90799
R55930 a_83153_n35156.t1 a_83153_n35156.t8 7.90799
R55931 a_83153_n35156.n1 a_83153_n35156.t7 7.41865
R55932 a_83153_n35156.t8 a_83153_n35156.t3 7.41865
R55933 a_83153_n35156.t8 a_83153_n35156.n0 7.31642
R55934 a_56895_n16009.t0 a_56895_n16009.t1 97.9575
R55935 a_56895_n16009.t1 a_56895_n16009.t2 15.0742
R55936 a_30324_n29313.t0 a_30324_n29313.t2 23.2303
R55937 a_30324_n29313.t0 a_30324_n29313.t1 21.6695
R55938 a_112559_n29181.n0 a_112559_n29181.t14 10.2515
R55939 a_112559_n29181.n1 a_112559_n29181.t9 10.2515
R55940 a_112559_n29181.n0 a_112559_n29181.t20 10.2515
R55941 a_112559_n29181.n0 a_112559_n29181.t3 10.2515
R55942 a_112559_n29181.n0 a_112559_n29181.t7 10.096
R55943 a_112559_n29181.n1 a_112559_n29181.t16 10.0935
R55944 a_112559_n29181.n0 a_112559_n29181.t5 10.0859
R55945 a_112559_n29181.n0 a_112559_n29181.t21 10.0808
R55946 a_112559_n29181.n0 a_112559_n29181.t13 9.53981
R55947 a_112559_n29181.n1 a_112559_n29181.t11 9.53981
R55948 a_112559_n29181.n0 a_112559_n29181.t17 9.53981
R55949 a_112559_n29181.n0 a_112559_n29181.t19 9.53981
R55950 a_112559_n29181.n0 a_112559_n29181.t12 9.53744
R55951 a_112559_n29181.n1 a_112559_n29181.t22 9.53744
R55952 a_112559_n29181.n0 a_112559_n29181.t15 9.53744
R55953 a_112559_n29181.n0 a_112559_n29181.t18 9.53744
R55954 a_112559_n29181.n1 a_112559_n29181.n0 9.16839
R55955 a_112559_n29181.n1 a_112559_n29181.t4 8.14051
R55956 a_112559_n29181.n1 a_112559_n29181.t10 8.13798
R55957 a_112559_n29181.t0 a_112559_n29181.t1 7.95997
R55958 a_112559_n29181.t1 a_112559_n29181.t2 7.94576
R55959 a_112559_n29181.t1 a_112559_n29181.n1 7.50666
R55960 a_112559_n29181.n1 a_112559_n29181.t8 7.48675
R55961 a_112559_n29181.n1 a_112559_n29181.t6 7.48422
R55962 a_47819_10448.n0 a_47819_10448.t0 10.2828
R55963 a_47819_10448.t9 a_47819_10448.t2 10.2828
R55964 a_47819_10448.n0 a_47819_10448.t19 10.2828
R55965 a_47819_10448.n0 a_47819_10448.t15 10.2828
R55966 a_47819_10448.n0 a_47819_10448.t12 10.1333
R55967 a_47819_10448.t9 a_47819_10448.t13 10.1333
R55968 a_47819_10448.n0 a_47819_10448.t6 10.1333
R55969 a_47819_10448.n0 a_47819_10448.t4 10.1333
R55970 a_47819_10448.n0 a_47819_10448.t18 9.57156
R55971 a_47819_10448.n0 a_47819_10448.t16 9.57156
R55972 a_47819_10448.t9 a_47819_10448.t17 9.57156
R55973 a_47819_10448.n0 a_47819_10448.t11 9.57156
R55974 a_47819_10448.n0 a_47819_10448.t22 9.57156
R55975 a_47819_10448.n0 a_47819_10448.t20 9.57156
R55976 a_47819_10448.t9 a_47819_10448.t21 9.57156
R55977 a_47819_10448.n0 a_47819_10448.t14 9.57156
R55978 a_47819_10448.t9 a_47819_10448.n1 8.94763
R55979 a_47819_10448.t9 a_47819_10448.t10 8.02945
R55980 a_47819_10448.t9 a_47819_10448.t8 8.02708
R55981 a_47819_10448.n1 a_47819_10448.t3 7.90829
R55982 a_47819_10448.t1 a_47819_10448.t9 7.90829
R55983 a_47819_10448.n1 a_47819_10448.t5 7.41776
R55984 a_47819_10448.t9 a_47819_10448.t7 7.41776
R55985 a_47819_10448.t9 a_47819_10448.n0 7.31642
R55986 a_47819_n36322.n0 a_47819_n36322.t13 13.7934
R55987 a_47819_n36322.n2 a_47819_n36322.t1 10.7024
R55988 a_47819_n36322.n2 a_47819_n36322.t4 10.1668
R55989 a_47819_n36322.n2 a_47819_n36322.t7 9.64458
R55990 a_47819_n36322.n2 a_47819_n36322.t3 9.27635
R55991 a_47819_n36322.n2 a_47819_n36322.n0 8.75198
R55992 a_47819_n36322.n0 a_47819_n36322.t17 8.14051
R55993 a_47819_n36322.n0 a_47819_n36322.t15 8.14051
R55994 a_47819_n36322.n0 a_47819_n36322.t23 8.14051
R55995 a_47819_n36322.n0 a_47819_n36322.t8 8.14051
R55996 a_47819_n36322.n0 a_47819_n36322.t14 8.06917
R55997 a_47819_n36322.n0 a_47819_n36322.t12 8.06917
R55998 a_47819_n36322.n0 a_47819_n36322.t11 8.06917
R55999 a_47819_n36322.n0 a_47819_n36322.t22 8.06917
R56000 a_47819_n36322.n0 a_47819_n36322.t20 8.06917
R56001 a_47819_n36322.n0 a_47819_n36322.t16 8.06917
R56002 a_47819_n36322.n0 a_47819_n36322.t19 8.06917
R56003 a_47819_n36322.n1 a_47819_n36322.t5 7.94157
R56004 a_47819_n36322.n2 a_47819_n36322.t2 7.72643
R56005 a_47819_n36322.n1 a_47819_n36322.t6 7.22925
R56006 a_47819_n36322.t0 a_47819_n36322.n2 7.17912
R56007 a_47819_n36322.n0 a_47819_n36322.t21 8.33554
R56008 a_47819_n36322.t18 a_47819_n36322.n0 8.33554
R56009 a_47819_n36322.n0 a_47819_n36322.t9 8.33647
R56010 a_47819_n36322.t10 a_47819_n36322.n0 8.33647
R56011 a_47819_n36322.n2 a_47819_n36322.n1 7.46075
R56012 a_83325_4421.t2 a_83325_4421.t0 21.6693
R56013 a_83325_4421.t1 a_83325_4421.t0 15.3476
R56014 a_84017_n17715.t0 a_84017_n17715.t2 49.0231
R56015 a_84017_n17715.t2 a_84017_n17715.t3 12.9273
R56016 a_84017_n17715.t2 a_84017_n17715.t5 10.1307
R56017 a_84017_n17715.t2 a_84017_n17715.t4 8.54643
R56018 a_84017_n17715.t2 a_84017_n17715.t1 7.50895
R56019 a_83153_n36322.n0 a_83153_n36322.t16 13.7934
R56020 a_83153_n36322.n2 a_83153_n36322.t6 10.7024
R56021 a_83153_n36322.n2 a_83153_n36322.t3 10.1668
R56022 a_83153_n36322.n2 a_83153_n36322.t1 9.64458
R56023 a_83153_n36322.n2 a_83153_n36322.t7 9.27635
R56024 a_83153_n36322.n2 a_83153_n36322.n0 8.75198
R56025 a_83153_n36322.n0 a_83153_n36322.t22 8.14051
R56026 a_83153_n36322.n0 a_83153_n36322.t20 8.14051
R56027 a_83153_n36322.n0 a_83153_n36322.t10 8.14051
R56028 a_83153_n36322.n0 a_83153_n36322.t13 8.14051
R56029 a_83153_n36322.n0 a_83153_n36322.t17 8.06917
R56030 a_83153_n36322.n0 a_83153_n36322.t11 8.06917
R56031 a_83153_n36322.n0 a_83153_n36322.t9 8.06917
R56032 a_83153_n36322.n0 a_83153_n36322.t8 8.06917
R56033 a_83153_n36322.n0 a_83153_n36322.t23 8.06917
R56034 a_83153_n36322.n0 a_83153_n36322.t15 8.06917
R56035 a_83153_n36322.n0 a_83153_n36322.t18 8.06917
R56036 a_83153_n36322.n1 a_83153_n36322.t0 7.94157
R56037 a_83153_n36322.n2 a_83153_n36322.t5 7.72643
R56038 a_83153_n36322.n1 a_83153_n36322.t2 7.22925
R56039 a_83153_n36322.t4 a_83153_n36322.n2 7.17912
R56040 a_83153_n36322.n0 a_83153_n36322.t14 8.33554
R56041 a_83153_n36322.t12 a_83153_n36322.n0 8.33554
R56042 a_83153_n36322.n0 a_83153_n36322.t19 8.33647
R56043 a_83153_n36322.t21 a_83153_n36322.n0 8.33647
R56044 a_83153_n36322.n2 a_83153_n36322.n1 7.46075
R56045 a_83153_10448.n0 a_83153_10448.t10 10.2828
R56046 a_83153_10448.n1 a_83153_10448.t8 10.2828
R56047 a_83153_10448.n0 a_83153_10448.t17 10.2828
R56048 a_83153_10448.n0 a_83153_10448.t12 10.2828
R56049 a_83153_10448.n0 a_83153_10448.t20 10.1333
R56050 a_83153_10448.n1 a_83153_10448.t21 10.1333
R56051 a_83153_10448.n0 a_83153_10448.t6 10.1333
R56052 a_83153_10448.n0 a_83153_10448.t4 10.1333
R56053 a_83153_10448.n0 a_83153_10448.t19 9.57156
R56054 a_83153_10448.n0 a_83153_10448.t15 9.57156
R56055 a_83153_10448.n1 a_83153_10448.t16 9.57156
R56056 a_83153_10448.n0 a_83153_10448.t23 9.57156
R56057 a_83153_10448.n0 a_83153_10448.t18 9.57156
R56058 a_83153_10448.n0 a_83153_10448.t13 9.57156
R56059 a_83153_10448.n1 a_83153_10448.t14 9.57156
R56060 a_83153_10448.n0 a_83153_10448.t22 9.57156
R56061 a_83153_10448.n1 a_83153_10448.t3 8.02945
R56062 a_83153_10448.n1 a_83153_10448.t2 8.02708
R56063 a_83153_10448.n2 a_83153_10448.t9 7.90829
R56064 a_83153_10448.t11 a_83153_10448.n3 7.90829
R56065 a_83153_10448.n2 a_83153_10448.t5 7.41776
R56066 a_83153_10448.n3 a_83153_10448.t7 7.41776
R56067 a_83153_10448.n1 a_83153_10448.n0 7.31642
R56068 a_83153_10448.n1 a_83153_10448.t0 6.88906
R56069 a_83153_10448.n1 a_83153_10448.t1 6.88669
R56070 a_83153_10448.n1 a_83153_10448.n2 4.5005
R56071 a_83153_10448.n3 a_83153_10448.n1 4.44762
R56072 a_47819_11614.n2 a_47819_11614.t12 12.8637
R56073 a_47819_11614.t0 a_47819_11614.n1 10.7018
R56074 a_47819_11614.n1 a_47819_11614.t4 10.1659
R56075 a_47819_11614.n1 a_47819_11614.t6 9.64387
R56076 a_47819_11614.n1 a_47819_11614.t3 9.27665
R56077 a_47819_11614.n1 a_47819_11614.n2 8.75198
R56078 a_47819_11614.n2 a_47819_11614.t23 8.14051
R56079 a_47819_11614.n2 a_47819_11614.t19 8.14051
R56080 a_47819_11614.n2 a_47819_11614.t17 8.14051
R56081 a_47819_11614.n2 a_47819_11614.t10 8.14051
R56082 a_47819_11614.n2 a_47819_11614.t14 8.06917
R56083 a_47819_11614.n2 a_47819_11614.t11 8.06917
R56084 a_47819_11614.n2 a_47819_11614.t20 8.06917
R56085 a_47819_11614.n2 a_47819_11614.t8 8.06917
R56086 a_47819_11614.n2 a_47819_11614.t22 8.06917
R56087 a_47819_11614.n2 a_47819_11614.t16 8.06917
R56088 a_47819_11614.n2 a_47819_11614.t18 8.06917
R56089 a_47819_11614.n0 a_47819_11614.t7 7.94068
R56090 a_47819_11614.n1 a_47819_11614.t1 7.72524
R56091 a_47819_11614.n0 a_47819_11614.t5 7.22855
R56092 a_47819_11614.n1 a_47819_11614.t2 7.17942
R56093 a_47819_11614.t9 a_47819_11614.n2 8.33649
R56094 a_47819_11614.n2 a_47819_11614.t13 8.33649
R56095 a_47819_11614.t15 a_47819_11614.n2 8.33556
R56096 a_47819_11614.n2 a_47819_11614.t21 8.33556
R56097 a_47819_11614.n1 a_47819_11614.n0 7.46075
R56098 a_47991_4421.t2 a_47991_4421.t0 21.6693
R56099 a_47991_4421.t1 a_47991_4421.t0 15.3476
R56100 a_57977_n5344.t0 a_57977_n5344.t1 13.2434
R56101 a_103997_n8770.t0 a_103997_n8770.n3 39.3605
R56102 a_103997_n8770.n1 a_103997_n8770.n0 10.9327
R56103 a_103997_n8770.n0 a_103997_n8770.t12 8.44198
R56104 a_103997_n8770.n0 a_103997_n8770.t8 8.44198
R56105 a_103997_n8770.n1 a_103997_n8770.t11 8.44198
R56106 a_103997_n8770.n1 a_103997_n8770.t7 8.44198
R56107 a_103997_n8770.n0 a_103997_n8770.t5 9.26917
R56108 a_103997_n8770.n1 a_103997_n8770.t6 8.10567
R56109 a_103997_n8770.n3 a_103997_n8770.t1 6.51122
R56110 a_103997_n8770.n3 a_103997_n8770.n0 6.50622
R56111 a_103997_n8770.t1 a_103997_n8770.t2 6.36267
R56112 a_103997_n8770.t1 a_103997_n8770.n2 4.84877
R56113 a_103997_n8770.n2 a_103997_n8770.t4 3.65383
R56114 a_103997_n8770.n1 a_103997_n8770.t10 8.65827
R56115 a_103997_n8770.n2 a_103997_n8770.t3 3.57094
R56116 a_103997_n8770.n0 a_103997_n8770.t9 8.77499
R56117 a_47991_5507.t1 a_47991_5507.t2 24.9014
R56118 a_47991_5507.t0 a_47991_5507.t1 15.5881
R56119 a_48951_4481.t0 a_48951_4481.t1 26.1287
R56120 a_48951_4481.t1 a_48951_4481.t2 15.0742
R56121 a_47991_n29313.t0 a_47991_n29313.t1 23.2303
R56122 a_47991_n29313.t0 a_47991_n29313.t2 21.6695
R56123 a_59558_n29181.n0 a_59558_n29181.t11 10.2515
R56124 a_59558_n29181.n1 a_59558_n29181.t5 10.2515
R56125 a_59558_n29181.n0 a_59558_n29181.t17 10.2515
R56126 a_59558_n29181.n0 a_59558_n29181.t3 10.2515
R56127 a_59558_n29181.n0 a_59558_n29181.t7 10.096
R56128 a_59558_n29181.n1 a_59558_n29181.t18 10.0935
R56129 a_59558_n29181.n0 a_59558_n29181.t9 10.0859
R56130 a_59558_n29181.n0 a_59558_n29181.t12 10.0808
R56131 a_59558_n29181.n0 a_59558_n29181.t22 9.53981
R56132 a_59558_n29181.n1 a_59558_n29181.t20 9.53981
R56133 a_59558_n29181.n0 a_59558_n29181.t14 9.53981
R56134 a_59558_n29181.n0 a_59558_n29181.t16 9.53981
R56135 a_59558_n29181.n0 a_59558_n29181.t21 9.53744
R56136 a_59558_n29181.n1 a_59558_n29181.t19 9.53744
R56137 a_59558_n29181.n0 a_59558_n29181.t13 9.53744
R56138 a_59558_n29181.n0 a_59558_n29181.t15 9.53744
R56139 a_59558_n29181.n1 a_59558_n29181.n0 9.16839
R56140 a_59558_n29181.n1 a_59558_n29181.t4 8.14051
R56141 a_59558_n29181.n1 a_59558_n29181.t6 8.13798
R56142 a_59558_n29181.t0 a_59558_n29181.t2 7.95997
R56143 a_59558_n29181.t0 a_59558_n29181.t1 7.94576
R56144 a_59558_n29181.t0 a_59558_n29181.n1 7.50666
R56145 a_59558_n29181.n1 a_59558_n29181.t8 7.48675
R56146 a_59558_n29181.n1 a_59558_n29181.t10 7.48422
R56147 a_53675_n30339.n0 a_53675_n30339.t1 10.3838
R56148 a_53675_n30339.n0 a_53675_n30339.t3 10.3566
R56149 a_53675_n30339.n0 a_53675_n30339.t2 10.0407
R56150 a_53675_n30339.t0 a_53675_n30339.n0 9.57605
R56151 a_60677_n36322.t0 a_60677_n36322.t1 83.5159
R56152 a_60677_n36322.t1 a_60677_n36322.t3 9.77323
R56153 a_60677_n36322.t1 a_60677_n36322.t2 8.17727
R56154 a_65486_11614.n2 a_65486_11614.t23 12.8637
R56155 a_65486_11614.n1 a_65486_11614.t3 10.7018
R56156 a_65486_11614.n1 a_65486_11614.t4 10.1659
R56157 a_65486_11614.n1 a_65486_11614.t7 9.64387
R56158 a_65486_11614.n1 a_65486_11614.t1 9.27665
R56159 a_65486_11614.n1 a_65486_11614.n2 8.75198
R56160 a_65486_11614.n2 a_65486_11614.t18 8.14051
R56161 a_65486_11614.n2 a_65486_11614.t14 8.14051
R56162 a_65486_11614.n2 a_65486_11614.t10 8.14051
R56163 a_65486_11614.n2 a_65486_11614.t22 8.14051
R56164 a_65486_11614.n2 a_65486_11614.t15 8.06917
R56165 a_65486_11614.n2 a_65486_11614.t11 8.06917
R56166 a_65486_11614.n2 a_65486_11614.t16 8.06917
R56167 a_65486_11614.n2 a_65486_11614.t20 8.06917
R56168 a_65486_11614.n2 a_65486_11614.t8 8.06917
R56169 a_65486_11614.n2 a_65486_11614.t19 8.06917
R56170 a_65486_11614.n2 a_65486_11614.t12 8.06917
R56171 a_65486_11614.n0 a_65486_11614.t6 7.94068
R56172 a_65486_11614.n1 a_65486_11614.t2 7.72524
R56173 a_65486_11614.n0 a_65486_11614.t5 7.22855
R56174 a_65486_11614.t0 a_65486_11614.n1 7.17942
R56175 a_65486_11614.t13 a_65486_11614.n2 8.33649
R56176 a_65486_11614.n2 a_65486_11614.t17 8.33649
R56177 a_65486_11614.t21 a_65486_11614.n2 8.33556
R56178 a_65486_11614.n2 a_65486_11614.t9 8.33556
R56179 a_65486_11614.n1 a_65486_11614.n0 7.46075
R56180 a_53829_10388.n5 a_53829_10388.n1 10.2377
R56181 a_53829_10388.n4 a_53829_10388.t6 10.2108
R56182 a_53829_10388.n4 a_53829_10388.t5 9.99909
R56183 a_53829_10388.n5 a_53829_10388.t1 9.80443
R56184 a_53829_10388.n5 a_53829_10388.t7 9.55135
R56185 a_53829_10388.n0 a_53829_10388.t16 8.17385
R56186 a_53829_10388.n3 a_53829_10388.t9 8.17299
R56187 a_53829_10388.n3 a_53829_10388.t10 8.17134
R56188 a_53829_10388.n0 a_53829_10388.t8 8.16754
R56189 a_53829_10388.n1 a_53829_10388.t20 8.10567
R56190 a_53829_10388.n1 a_53829_10388.t19 8.10567
R56191 a_53829_10388.n3 a_53829_10388.t15 8.10567
R56192 a_53829_10388.n3 a_53829_10388.t17 8.10567
R56193 a_53829_10388.n1 a_53829_10388.t18 8.10567
R56194 a_53829_10388.n1 a_53829_10388.t23 8.10567
R56195 a_53829_10388.n0 a_53829_10388.t22 8.10567
R56196 a_53829_10388.n0 a_53829_10388.t13 8.10567
R56197 a_53829_10388.n6 a_53829_10388.t4 7.74799
R56198 a_53829_10388.n7 a_53829_10388.t2 7.73052
R56199 a_53829_10388.n6 a_53829_10388.t3 7.46478
R56200 a_53829_10388.t0 a_53829_10388.n7 7.1311
R56201 a_53829_10388.n4 a_53829_10388.n6 2.2505
R56202 a_53829_10388.n7 a_53829_10388.n5 2.2505
R56203 a_53829_10388.n1 a_53829_10388.t11 8.35731
R56204 a_53829_10388.n0 a_53829_10388.t21 8.38107
R56205 a_53829_10388.n1 a_53829_10388.t12 8.37583
R56206 a_53829_10388.n1 a_53829_10388.n0 4.35656
R56207 a_53829_10388.n5 a_53829_10388.n4 2.96863
R56208 a_53829_10388.n2 a_53829_10388.n1 1.0882
R56209 a_53829_10388.n2 a_53829_10388.n3 1.08408
R56210 a_53829_10388.n2 a_53829_10388.t14 8.66753
R56211 a_53699_13546.n1 a_53699_13546.n0 26.5254
R56212 a_53699_13546.n1 a_53699_13546.t1 11.5094
R56213 a_53699_13546.n0 a_53699_13546.t2 10.937
R56214 a_53699_13546.n0 a_53699_13546.t3 9.33982
R56215 a_53699_13546.t0 a_53699_13546.n1 9.24966
R56216 a_53699_11614.t0 a_53699_11614.n2 58.3955
R56217 a_53699_11614.n1 a_53699_11614.n0 10.9309
R56218 a_53699_11614.t1 a_53699_11614.t2 8.5021
R56219 a_53699_11614.n1 a_53699_11614.t9 8.44198
R56220 a_53699_11614.n1 a_53699_11614.t3 8.44198
R56221 a_53699_11614.n0 a_53699_11614.t6 8.44198
R56222 a_53699_11614.n0 a_53699_11614.t10 8.44198
R56223 a_53699_11614.n1 a_53699_11614.t4 8.10567
R56224 a_53699_11614.n0 a_53699_11614.t5 9.26955
R56225 a_53699_11614.n2 a_53699_11614.t1 6.51122
R56226 a_53699_11614.n2 a_53699_11614.n0 6.50622
R56227 a_53699_11614.n1 a_53699_11614.t7 8.65823
R56228 a_53699_11614.n0 a_53699_11614.t8 8.77493
R56229 a_65658_4421.t1 a_65658_4421.t0 21.6693
R56230 a_65658_4421.t2 a_65658_4421.t0 15.3476
R56231 I1N.n8 I1N.t1 10.2879
R56232 I1N.n32 I1N.n31 6.37738
R56233 I1N.t0 I1N.n9 4.39661
R56234 I1N.n7 I1N.t12 4.39661
R56235 I1N.t17 I1N.n1 4.39661
R56236 I1N.t6 I1N.n25 4.39661
R56237 I1N.n10 I1N.t0 4.39661
R56238 I1N.n26 I1N.t6 4.39661
R56239 I1N.n13 I1N.t7 4.39651
R56240 I1N.n12 I1N.t7 4.39651
R56241 I1N.n21 I1N.t4 4.39651
R56242 I1N.n19 I1N.t10 4.39651
R56243 I1N.n29 I1N.t2 4.39651
R56244 I1N.n28 I1N.t2 4.39651
R56245 I1N.n32 I1N.t3 3.9368
R56246 I1N.n13 I1N.t9 2.96638
R56247 I1N.t9 I1N.n12 2.96638
R56248 I1N.t14 I1N.n9 2.96638
R56249 I1N.n10 I1N.t14 2.96638
R56250 I1N.t8 I1N.n1 2.96638
R56251 I1N.n7 I1N.t5 2.96638
R56252 I1N.n21 I1N.t11 2.96638
R56253 I1N.n29 I1N.t16 2.96638
R56254 I1N.t16 I1N.n28 2.96638
R56255 I1N.t13 I1N.n25 2.96638
R56256 I1N.n26 I1N.t13 2.96638
R56257 I1N.t15 I1N.n19 2.96638
R56258 I1N.n6 I1N.t8 2.52844
R56259 I1N.n18 I1N.t4 2.52844
R56260 I1N.t10 I1N.n18 2.52844
R56261 I1N.t5 I1N.n6 2.52844
R56262 I1N.n3 I1N.t12 2.52844
R56263 I1N.n20 I1N.t15 2.52844
R56264 I1N.t11 I1N.n20 2.52844
R56265 I1N.n3 I1N.t17 2.52844
R56266 I1N.n31 I1N.n30 1.5005
R56267 I1N.n27 I1N.n24 1.5005
R56268 I1N.n23 I1N.n22 1.5005
R56269 I1N.n4 I1N.n0 1.5005
R56270 I1N.n17 I1N.n16 1.5005
R56271 I1N.n15 I1N.n14 1.5005
R56272 I1N.n11 I1N.n8 1.5005
R56273 I1N.n5 I1N.n4 1.19221
R56274 I1N.n4 I1N.n2 1.16411
R56275 I1N.n11 I1N.n10 0.88285
R56276 I1N.n14 I1N.n9 0.88285
R56277 I1N.n17 I1N.n7 0.88285
R56278 I1N.n22 I1N.n1 0.88285
R56279 I1N.n27 I1N.n26 0.88285
R56280 I1N.n30 I1N.n25 0.88285
R56281 I1N.n12 I1N.n11 0.858643
R56282 I1N.n14 I1N.n13 0.858643
R56283 I1N.n19 I1N.n17 0.858643
R56284 I1N.n22 I1N.n21 0.858643
R56285 I1N.n28 I1N.n27 0.858643
R56286 I1N.n30 I1N.n29 0.858643
R56287 I1N.n18 I1N.n2 0.367144
R56288 I1N.n5 I1N.n3 0.365787
R56289 I1N.n16 I1N.n0 0.210297
R56290 I1N.n23 I1N.n0 0.207257
R56291 I1N.n31 I1N.n24 0.1805
R56292 I1N.n15 I1N.n8 0.179588
R56293 I1N.n16 I1N.n15 0.0935405
R56294 I1N.n24 I1N.n23 0.0935405
R56295 I1N.n6 I1N.n5 0.0804816
R56296 I1N.n20 I1N.n2 0.0795377
R56297 I1N I1N.n32 0.0159334
R56298 a_89715_n16810.t0 a_89715_n16810.t1 12.8122
R56299 a_71366_13546.n1 a_71366_13546.n0 26.5281
R56300 a_71366_13546.n0 a_71366_13546.t3 11.5094
R56301 a_71366_13546.t0 a_71366_13546.n1 10.937
R56302 a_71366_13546.n1 a_71366_13546.t1 9.33982
R56303 a_71366_13546.n0 a_71366_13546.t2 9.24966
R56304 a_36162_n36382.n5 a_36162_n36382.n1 10.2377
R56305 a_36162_n36382.n4 a_36162_n36382.t3 10.2105
R56306 a_36162_n36382.n4 a_36162_n36382.t2 9.99998
R56307 a_36162_n36382.n5 a_36162_n36382.t5 9.80532
R56308 a_36162_n36382.n5 a_36162_n36382.t6 9.55206
R56309 a_36162_n36382.n0 a_36162_n36382.t22 8.17385
R56310 a_36162_n36382.n3 a_36162_n36382.t20 8.17299
R56311 a_36162_n36382.n3 a_36162_n36382.t23 8.17134
R56312 a_36162_n36382.n0 a_36162_n36382.t21 8.16754
R56313 a_36162_n36382.n1 a_36162_n36382.t9 8.10567
R56314 a_36162_n36382.n1 a_36162_n36382.t17 8.10567
R56315 a_36162_n36382.n3 a_36162_n36382.t15 8.10567
R56316 a_36162_n36382.n3 a_36162_n36382.t8 8.10567
R56317 a_36162_n36382.n1 a_36162_n36382.t12 8.10567
R56318 a_36162_n36382.n1 a_36162_n36382.t16 8.10567
R56319 a_36162_n36382.n0 a_36162_n36382.t14 8.10567
R56320 a_36162_n36382.n0 a_36162_n36382.t10 8.10567
R56321 a_36162_n36382.n6 a_36162_n36382.t1 7.74888
R56322 a_36162_n36382.n7 a_36162_n36382.t7 7.73141
R56323 a_36162_n36382.n6 a_36162_n36382.t0 7.46359
R56324 a_36162_n36382.t4 a_36162_n36382.n7 7.13081
R56325 a_36162_n36382.n4 a_36162_n36382.n6 2.2505
R56326 a_36162_n36382.n7 a_36162_n36382.n5 2.2505
R56327 a_36162_n36382.t13 a_36162_n36382.n1 8.35729
R56328 a_36162_n36382.n1 a_36162_n36382.t11 8.37586
R56329 a_36162_n36382.n0 a_36162_n36382.t18 8.38104
R56330 a_36162_n36382.n1 a_36162_n36382.n0 4.35658
R56331 a_36162_n36382.n5 a_36162_n36382.n4 2.96863
R56332 a_36162_n36382.n2 a_36162_n36382.n1 1.08819
R56333 a_36162_n36382.n2 a_36162_n36382.n3 1.08408
R56334 a_36162_n36382.n2 a_36162_n36382.t19 8.6675
R56335 a_71342_7563.t2 a_71342_7563.n0 10.3829
R56336 a_71342_7563.n0 a_71342_7563.t0 10.3566
R56337 a_71342_7563.n0 a_71342_7563.t1 10.0407
R56338 a_71342_7563.n0 a_71342_7563.t3 9.57605
R56339 a_71366_11614.t0 a_71366_11614.n2 42.1702
R56340 a_71366_11614.n1 a_71366_11614.n0 10.9309
R56341 a_71366_11614.t1 a_71366_11614.t2 8.5021
R56342 a_71366_11614.n1 a_71366_11614.t7 8.44198
R56343 a_71366_11614.n1 a_71366_11614.t3 8.44198
R56344 a_71366_11614.n0 a_71366_11614.t4 8.44198
R56345 a_71366_11614.n0 a_71366_11614.t10 8.44198
R56346 a_71366_11614.n1 a_71366_11614.t5 8.10567
R56347 a_71366_11614.n0 a_71366_11614.t6 9.26955
R56348 a_71366_11614.n2 a_71366_11614.t1 6.51122
R56349 a_71366_11614.n2 a_71366_11614.n0 6.50622
R56350 a_71366_11614.n1 a_71366_11614.t8 8.65823
R56351 a_71366_11614.n0 a_71366_11614.t9 8.77493
R56352 a_78344_10448.t0 a_78344_10448.t1 44.9816
R56353 a_78344_10448.t1 a_78344_10448.t5 12.9273
R56354 a_78344_10448.t1 a_78344_10448.t4 10.1307
R56355 a_78344_10448.t1 a_78344_10448.t2 8.54643
R56356 a_78344_10448.t1 a_78344_10448.t3 7.50895
R56357 a_38097_n16007.t0 a_38097_n16007.t2 41.3378
R56358 a_38097_n16007.t2 a_38097_n16007.t1 18.4133
R56359 a_53675_4481.n0 a_53675_4481.t2 10.6581
R56360 a_53675_4481.n0 a_53675_4481.t1 10.2356
R56361 a_53675_4481.t0 a_53675_4481.n0 9.5019
R56362 a_53675_4481.n0 a_53675_4481.t3 9.34796
R56363 a_36162_10388.n6 a_36162_10388.n1 10.2377
R56364 a_36162_10388.n5 a_36162_10388.t2 10.2108
R56365 a_36162_10388.n5 a_36162_10388.t3 9.99909
R56366 a_36162_10388.n6 a_36162_10388.t6 9.80443
R56367 a_36162_10388.t4 a_36162_10388.n6 9.55135
R56368 a_36162_10388.n0 a_36162_10388.t20 8.17385
R56369 a_36162_10388.n3 a_36162_10388.t16 8.17299
R56370 a_36162_10388.n3 a_36162_10388.t17 8.17134
R56371 a_36162_10388.n0 a_36162_10388.t15 8.16754
R56372 a_36162_10388.n1 a_36162_10388.t14 8.10567
R56373 a_36162_10388.n1 a_36162_10388.t11 8.10567
R56374 a_36162_10388.n3 a_36162_10388.t9 8.10567
R56375 a_36162_10388.n3 a_36162_10388.t13 8.10567
R56376 a_36162_10388.n1 a_36162_10388.t10 8.10567
R56377 a_36162_10388.n1 a_36162_10388.t19 8.10567
R56378 a_36162_10388.n0 a_36162_10388.t18 8.10567
R56379 a_36162_10388.n0 a_36162_10388.t8 8.10567
R56380 a_36162_10388.n7 a_36162_10388.t1 7.74799
R56381 a_36162_10388.n4 a_36162_10388.t7 7.73052
R56382 a_36162_10388.n7 a_36162_10388.t0 7.46478
R56383 a_36162_10388.n4 a_36162_10388.t5 7.1311
R56384 a_36162_10388.n5 a_36162_10388.n7 2.2505
R56385 a_36162_10388.n6 a_36162_10388.n4 2.2505
R56386 a_36162_10388.n1 a_36162_10388.t21 8.35731
R56387 a_36162_10388.n0 a_36162_10388.t12 8.38107
R56388 a_36162_10388.n1 a_36162_10388.t22 8.37583
R56389 a_36162_10388.n1 a_36162_10388.n0 4.35656
R56390 a_36162_10388.n6 a_36162_10388.n5 2.96863
R56391 a_36162_10388.n2 a_36162_10388.n1 1.0882
R56392 a_36162_10388.n2 a_36162_10388.n3 1.08408
R56393 a_36162_10388.n2 a_36162_10388.t23 8.66753
R56394 a_32913_n5342.t0 a_32913_n5342.t1 13.2434
R56395 a_65658_n29313.t0 a_65658_n29313.t1 23.2303
R56396 a_65658_n29313.t0 a_65658_n29313.t2 21.6695
R56397 a_39179_n16007.t0 a_39179_n16007.t1 13.2434
R56398 a_71366_n36322.n1 a_71366_n36322.n0 26.5281
R56399 a_71366_n36322.n1 a_71366_n36322.t1 11.5094
R56400 a_71366_n36322.n0 a_71366_n36322.t3 10.937
R56401 a_71366_n36322.n0 a_71366_n36322.t2 9.33982
R56402 a_71366_n36322.t0 a_71366_n36322.n1 9.24966
R56403 a_30324_5507.t0 a_30324_5507.t1 30.2725
R56404 a_30324_5507.t1 a_30324_5507.t2 24.9014
R56405 a_71342_n27257.n0 a_71342_n27257.t2 10.6581
R56406 a_71342_n27257.n0 a_71342_n27257.t1 10.2358
R56407 a_71342_n27257.t0 a_71342_n27257.n0 9.50202
R56408 a_71342_n27257.n0 a_71342_n27257.t3 9.34796
R56409 a_50629_n16009.t0 a_50629_n16009.t1 82.9933
R56410 a_50629_n16009.t1 a_50629_n16009.t2 15.0742
R56411 a_39179_n8930.t0 a_39179_n8930.t1 118.243
R56412 a_39179_n8930.t1 a_39179_n8930.t2 24.9025
R56413 a_106676_7563.t0 a_106676_7563.n0 10.3829
R56414 a_106676_7563.n0 a_106676_7563.t2 10.3566
R56415 a_106676_7563.n0 a_106676_7563.t3 10.0407
R56416 a_106676_7563.n0 a_106676_7563.t1 9.57605
R56417 a_106830_n36382.n5 a_106830_n36382.n1 10.2377
R56418 a_106830_n36382.n4 a_106830_n36382.t7 10.2105
R56419 a_106830_n36382.n4 a_106830_n36382.t5 9.99998
R56420 a_106830_n36382.n5 a_106830_n36382.t1 9.80532
R56421 a_106830_n36382.n5 a_106830_n36382.t3 9.55206
R56422 a_106830_n36382.n0 a_106830_n36382.t20 8.17385
R56423 a_106830_n36382.n3 a_106830_n36382.t16 8.17299
R56424 a_106830_n36382.n3 a_106830_n36382.t21 8.17134
R56425 a_106830_n36382.n0 a_106830_n36382.t17 8.16754
R56426 a_106830_n36382.n1 a_106830_n36382.t18 8.10567
R56427 a_106830_n36382.n1 a_106830_n36382.t23 8.10567
R56428 a_106830_n36382.n3 a_106830_n36382.t15 8.10567
R56429 a_106830_n36382.n3 a_106830_n36382.t10 8.10567
R56430 a_106830_n36382.n1 a_106830_n36382.t19 8.10567
R56431 a_106830_n36382.n1 a_106830_n36382.t22 8.10567
R56432 a_106830_n36382.n0 a_106830_n36382.t14 8.10567
R56433 a_106830_n36382.n0 a_106830_n36382.t13 8.10567
R56434 a_106830_n36382.n6 a_106830_n36382.t6 7.74888
R56435 a_106830_n36382.n7 a_106830_n36382.t2 7.73141
R56436 a_106830_n36382.n6 a_106830_n36382.t4 7.46359
R56437 a_106830_n36382.t0 a_106830_n36382.n7 7.13081
R56438 a_106830_n36382.n4 a_106830_n36382.n6 2.2505
R56439 a_106830_n36382.n7 a_106830_n36382.n5 2.2505
R56440 a_106830_n36382.t9 a_106830_n36382.n1 8.35729
R56441 a_106830_n36382.n1 a_106830_n36382.t8 8.37586
R56442 a_106830_n36382.n0 a_106830_n36382.t11 8.38104
R56443 a_106830_n36382.n1 a_106830_n36382.n0 4.35658
R56444 a_106830_n36382.n5 a_106830_n36382.n4 2.96863
R56445 a_106830_n36382.n2 a_106830_n36382.n1 1.08819
R56446 a_106830_n36382.n2 a_106830_n36382.n3 1.08408
R56447 a_106830_n36382.n2 a_106830_n36382.t12 8.6675
R56448 a_36008_7563.t0 a_36008_7563.n0 10.3829
R56449 a_36008_7563.n0 a_36008_7563.t3 10.3566
R56450 a_36008_7563.n0 a_36008_7563.t2 10.0407
R56451 a_36008_7563.n0 a_36008_7563.t1 9.57605
R56452 a_89009_7563.t2 a_89009_7563.n0 10.3829
R56453 a_89009_7563.n0 a_89009_7563.t1 10.3566
R56454 a_89009_7563.n0 a_89009_7563.t0 10.0407
R56455 a_89009_7563.n0 a_89009_7563.t3 9.57605
R56456 a_36032_13546.n1 a_36032_13546.n0 26.5241
R56457 a_36032_13546.n0 a_36032_13546.t3 11.5094
R56458 a_36032_13546.n1 a_36032_13546.t1 10.937
R56459 a_36032_13546.t0 a_36032_13546.n1 9.33982
R56460 a_36032_13546.n0 a_36032_13546.t2 9.24966
R56461 a_101111_n6055.t0 a_101111_n6055.t1 12.8122
R56462 IN_POS.n32 IN_POS.n31 17.0316
R56463 IN_POS.n15 IN_POS.n1 3.06497
R56464 IN_POS.n27 IN_POS.n0 2.80204
R56465 IN_POS.n23 IN_POS.n22 2.55189
R56466 IN_POS.n29 IN_POS.n28 2.44888
R56467 IN_POS.n13 IN_POS.n12 2.44888
R56468 IN_POS.n11 IN_POS.n10 2.44888
R56469 IN_POS.n17 IN_POS.n16 2.44888
R56470 IN_POS.n20 IN_POS.n19 2.44888
R56471 IN_POS.n25 IN_POS.n24 2.44888
R56472 IN_POS IN_POS.n32 2.30113
R56473 IN_POS IN_POS.n32 2.27938
R56474 IN_POS.n31 IN_POS.n0 1.75374
R56475 IN_POS.t0 IN_POS.n8 1.1935
R56476 IN_POS.t0 IN_POS.n18 1.19272
R56477 IN_POS.n23 IN_POS.n9 1.18175
R56478 IN_POS.n27 IN_POS.t0 1.0998
R56479 IN_POS.t0 IN_POS.n15 1.08916
R56480 IN_POS.n28 IN_POS.n27 0.958371
R56481 IN_POS.n17 IN_POS.n15 0.907386
R56482 IN_POS.t0 IN_POS.n9 0.752643
R56483 IN_POS.n13 IN_POS.n8 0.706267
R56484 IN_POS.n20 IN_POS.n18 0.672835
R56485 IN_POS.n16 IN_POS.n1 0.66672
R56486 IN_POS.t0 IN_POS.n14 0.629953
R56487 IN_POS.n30 IN_POS.n29 0.622487
R56488 IN_POS.t0 IN_POS.n21 0.604576
R56489 IN_POS.n25 IN_POS.n21 0.585642
R56490 IN_POS.n14 IN_POS.n11 0.583689
R56491 IN_POS.n21 IN_POS.n20 0.559641
R56492 IN_POS.n26 IN_POS.n25 0.549445
R56493 IN_POS.n28 IN_POS.n8 0.540673
R56494 IN_POS.n14 IN_POS.n13 0.529423
R56495 IN_POS.n18 IN_POS.n17 0.519089
R56496 IN_POS.n12 IN_POS.n7 0.514976
R56497 IN_POS.n19 IN_POS.n4 0.499862
R56498 IN_POS.t1 IN_POS.n30 0.47657
R56499 IN_POS.n30 IN_POS.n0 0.424689
R56500 IN_POS.n29 IN_POS.n7 0.383261
R56501 IN_POS.n16 IN_POS.n4 0.36773
R56502 IN_POS.n10 IN_POS.n6 0.365351
R56503 IN_POS.n24 IN_POS.n3 0.362981
R56504 IN_POS.n19 IN_POS.n3 0.348693
R56505 IN_POS.n12 IN_POS.n6 0.337682
R56506 IN_POS.t1 IN_POS.n1 0.323064
R56507 IN_POS.t1 IN_POS.n4 0.304037
R56508 IN_POS.t1 IN_POS.n7 0.300094
R56509 IN_POS.n10 IN_POS.n5 0.256772
R56510 IN_POS.n24 IN_POS.n2 0.246737
R56511 IN_POS.t1 IN_POS.n6 0.136362
R56512 IN_POS.t1 IN_POS.n3 0.128975
R56513 IN_POS.n11 IN_POS.n9 0.104562
R56514 IN_POS.n22 IN_POS.n2 0.0290825
R56515 IN_POS.n22 IN_POS.n5 0.0207691
R56516 IN_POS.n26 IN_POS.n23 0.00666077
R56517 IN_POS.t1 IN_POS.n2 0.00482948
R56518 IN_POS.t0 IN_POS.n26 0.00449532
R56519 IN_POS.t1 IN_POS.n5 0.00410811
R56520 IN_POS.n31 IN_POS.t1 0.00330619
R56521 a_94892_4481.n1 a_94892_4481.t2 10.2515
R56522 a_94892_4481.n1 a_94892_4481.t0 10.2515
R56523 a_94892_4481.n1 a_94892_4481.t14 10.2515
R56524 a_94892_4481.n1 a_94892_4481.t20 10.2515
R56525 a_94892_4481.n1 a_94892_4481.t4 10.096
R56526 a_94892_4481.n1 a_94892_4481.t13 10.0935
R56527 a_94892_4481.n1 a_94892_4481.t6 10.0859
R56528 a_94892_4481.n1 a_94892_4481.t19 10.0808
R56529 a_94892_4481.n1 a_94892_4481.t22 9.53981
R56530 a_94892_4481.n1 a_94892_4481.t18 9.53981
R56531 a_94892_4481.n1 a_94892_4481.t12 9.53981
R56532 a_94892_4481.n1 a_94892_4481.t16 9.53981
R56533 a_94892_4481.n1 a_94892_4481.t21 9.53744
R56534 a_94892_4481.n1 a_94892_4481.t17 9.53744
R56535 a_94892_4481.n1 a_94892_4481.t11 9.53744
R56536 a_94892_4481.n1 a_94892_4481.t15 9.53744
R56537 a_94892_4481.n1 a_94892_4481.n0 8.41434
R56538 a_94892_4481.n1 a_94892_4481.t3 8.14082
R56539 a_94892_4481.n0 a_94892_4481.t1 8.13828
R56540 a_94892_4481.t8 a_94892_4481.t9 7.96115
R56541 a_94892_4481.t8 a_94892_4481.t10 7.94694
R56542 a_94892_4481.t8 a_94892_4481.n1 7.50666
R56543 a_94892_4481.n0 a_94892_4481.t5 7.48586
R56544 a_94892_4481.n1 a_94892_4481.t7 7.48333
R56545 a_89033_n36322.n1 a_89033_n36322.n0 26.5215
R56546 a_89033_n36322.n0 a_89033_n36322.t3 11.5094
R56547 a_89033_n36322.n1 a_89033_n36322.t1 10.937
R56548 a_89033_n36322.t0 a_89033_n36322.n1 9.33982
R56549 a_89033_n36322.n0 a_89033_n36322.t2 9.24966
R56550 a_53675_n27257.n0 a_53675_n27257.t3 10.6581
R56551 a_53675_n27257.t0 a_53675_n27257.n0 10.2348
R56552 a_53675_n27257.n0 a_53675_n27257.t1 9.50202
R56553 a_53675_n27257.n0 a_53675_n27257.t2 9.34796
R56554 a_51711_n16009.t0 a_51711_n16009.t1 13.2434
R56555 a_89715_n5150.t0 a_89715_n5150.t1 12.8122
R56556 a_64243_n5344.t0 a_64243_n5344.t1 13.2434
R56557 a_89009_4481.n0 a_89009_4481.t0 10.6581
R56558 a_89009_4481.t2 a_89009_4481.n0 10.2346
R56559 a_89009_4481.n0 a_89009_4481.t3 9.5029
R56560 a_89009_4481.n0 a_89009_4481.t1 9.34796
R56561 a_39179_n5342.t0 a_39179_n5342.t1 13.2434
R56562 a_106809_n6055.t0 a_106809_n6055.t1 12.8114
R56563 VCM.n1 VCM.t0 11.5094
R56564 VCM.n2 VCM.n1 10.2743
R56565 VCM.n1 VCM.t1 9.24966
R56566 VCM VCM.n2 4.98085
R56567 VCM.n2 VCM.n0 4.18387
R56568 VCM.n0 VCM.t2 0.111029
R56569 VCM.n0 VCM.t3 0.03175
R56570 a_36008_n30339.n0 a_36008_n30339.t3 10.3838
R56571 a_36008_n30339.n0 a_36008_n30339.t1 10.3566
R56572 a_36008_n30339.n0 a_36008_n30339.t0 10.0407
R56573 a_36008_n30339.t2 a_36008_n30339.n0 9.57605
R56574 a_89009_n30339.t2 a_89009_n30339.n0 10.3838
R56575 a_89009_n30339.n0 a_89009_n30339.t0 10.3566
R56576 a_89009_n30339.n0 a_89009_n30339.t1 10.0407
R56577 a_89009_n30339.n0 a_89009_n30339.t3 9.57605
R56578 a_112507_n17715.t0 a_112507_n17715.t1 12.8114
R56579 a_53675_7563.t0 a_53675_7563.n0 10.3829
R56580 a_53675_7563.n0 a_53675_7563.t3 10.3566
R56581 a_53675_7563.n0 a_53675_7563.t2 10.0407
R56582 a_53675_7563.n0 a_53675_7563.t1 9.57605
R56583 a_45445_n5342.t0 a_45445_n5342.t1 13.2434
R56584 a_43010_n36322.t0 a_43010_n36322.t3 99.4592
R56585 a_43010_n36322.t3 a_43010_n36322.t1 9.77323
R56586 a_43010_n36322.t3 a_43010_n36322.t2 8.17727
R56587 a_64243_n16009.t0 a_64243_n16009.t1 13.2434
R56588 a_57977_n16009.t0 a_57977_n16009.t1 13.2434
R56589 a_36008_n27257.n0 a_36008_n27257.t1 10.6581
R56590 a_36008_n27257.n0 a_36008_n27257.t3 10.2358
R56591 a_36008_n27257.t2 a_36008_n27257.n0 9.50202
R56592 a_36008_n27257.n0 a_36008_n27257.t0 9.34796
R56593 a_71266_n4019.t2 a_71266_n4019.t0 11.1705
R56594 a_84017_n5150.t0 a_84017_n5150.t1 12.8114
R56595 a_106676_n27257.n0 a_106676_n27257.t0 10.6581
R56596 a_106676_n27257.n0 a_106676_n27257.t3 10.2358
R56597 a_106676_n27257.t2 a_106676_n27257.n0 9.50202
R56598 a_106676_n27257.n0 a_106676_n27257.t1 9.34796
R56599 a_95413_n5150.t0 a_95413_n5150.t1 12.8114
R56600 a_112507_n6055.t0 a_112507_n6055.t1 12.8114
R56601 a_95413_n16810.t0 a_95413_n16810.t1 12.8114
R56602 a_32913_n16007.t0 a_32913_n16007.t1 13.2434
R56603 a_45445_n16007.t0 a_45445_n16007.t1 13.2434
R56604 IBPOUT IBPOUT.t0 3.31278
R56605 a_84017_n16810.t0 a_84017_n16810.t1 12.8122
R56606 IN_NEG.n30 IN_NEG.t0 24.6019
R56607 IN_NEG.n8 IN_NEG.n0 3.09085
R56608 IN_NEG.n29 IN_NEG.n7 3.06463
R56609 IN_NEG.n19 IN_NEG.n18 2.55189
R56610 IN_NEG.n13 IN_NEG.n12 2.44888
R56611 IN_NEG.n10 IN_NEG.n9 2.44888
R56612 IN_NEG.n22 IN_NEG.n21 2.44888
R56613 IN_NEG.n25 IN_NEG.n24 2.44888
R56614 IN_NEG.n28 IN_NEG.n27 2.44888
R56615 IN_NEG.n16 IN_NEG.n15 2.44888
R56616 IN_NEG IN_NEG.n30 2.29437
R56617 IN_NEG IN_NEG.n30 2.28612
R56618 IN_NEG.t0 IN_NEG.n1 1.1935
R56619 IN_NEG.t0 IN_NEG.n6 1.19272
R56620 IN_NEG.t0 IN_NEG.n0 1.0998
R56621 IN_NEG.t0 IN_NEG.n29 1.08916
R56622 IN_NEG.n9 IN_NEG.n0 0.958371
R56623 IN_NEG.n29 IN_NEG.n28 0.907386
R56624 IN_NEG.n12 IN_NEG.n1 0.706267
R56625 IN_NEG.n10 IN_NEG.n8 0.694516
R56626 IN_NEG.n24 IN_NEG.n6 0.672835
R56627 IN_NEG.n27 IN_NEG.n7 0.66725
R56628 IN_NEG.t0 IN_NEG.n2 0.629953
R56629 IN_NEG.t0 IN_NEG.n5 0.604576
R56630 IN_NEG.n21 IN_NEG.n5 0.585642
R56631 IN_NEG.n15 IN_NEG.n2 0.583689
R56632 IN_NEG.n15 IN_NEG.n3 0.563066
R56633 IN_NEG.n24 IN_NEG.n5 0.559641
R56634 IN_NEG.n9 IN_NEG.n1 0.540673
R56635 IN_NEG.n12 IN_NEG.n2 0.529423
R56636 IN_NEG.n28 IN_NEG.n6 0.519089
R56637 IN_NEG.n13 IN_NEG.n11 0.514976
R56638 IN_NEG.n21 IN_NEG.n4 0.513594
R56639 IN_NEG.n26 IN_NEG.n25 0.500509
R56640 IN_NEG.n11 IN_NEG.n10 0.383261
R56641 IN_NEG.n27 IN_NEG.n26 0.367123
R56642 IN_NEG.n16 IN_NEG.n14 0.365351
R56643 IN_NEG.n23 IN_NEG.n22 0.3637
R56644 IN_NEG.n25 IN_NEG.n23 0.347986
R56645 IN_NEG.n14 IN_NEG.n13 0.337682
R56646 IN_NEG.n8 IN_NEG.t1 0.323963
R56647 IN_NEG.t1 IN_NEG.n7 0.323141
R56648 IN_NEG.n26 IN_NEG.t1 0.304079
R56649 IN_NEG.n11 IN_NEG.t1 0.300094
R56650 IN_NEG.n22 IN_NEG.n20 0.247682
R56651 IN_NEG.n17 IN_NEG.n16 0.229987
R56652 IN_NEG.n19 IN_NEG.n17 0.222212
R56653 IN_NEG.n14 IN_NEG.t1 0.136362
R56654 IN_NEG.n23 IN_NEG.t1 0.129075
R56655 IN_NEG.n18 IN_NEG.n4 0.100573
R56656 IN_NEG.t0 IN_NEG.n4 0.0624826
R56657 IN_NEG.n17 IN_NEG.t1 0.0337966
R56658 IN_NEG.n20 IN_NEG.n19 0.0147343
R56659 IN_NEG.n18 IN_NEG.n3 0.00689777
R56660 IN_NEG.t0 IN_NEG.n3 0.00476406
R56661 IN_NEG.n20 IN_NEG.t1 0.00295152
R56662 IBNOUT IBNOUT.t0 3.42291
R56663 a_101111_n17715.t0 a_101111_n17715.t1 12.8114
C0 a_101641_n18620# VDD 1.15407f
C1 a_81205_n9675# VDD 1.03081f
C2 a_109695_n21335# VDD 1.27413f
C3 a_107339_n18620# VDD 1.18674f
C4 a_81205_n16810# VDD 1.20767f
C5 a_84547_n6960# VDD 1.15365f
C6 a_86903_n9675# VDD 1.03237f
C7 a_113037_n18620# VDD 1.1868f
C8 a_86903_n16810# VDD 1.27745f
C9 a_90245_n6960# VDD 1.18674f
C10 a_92601_n9675# VDD 1.40063f
C11 IN_POS IN_NEG 3.17862f
C12 VDD I1U 1.71173f
C13 a_92601_n16810# VDD 1.28143f
C14 a_95943_n6960# VDD 1.18674f
C15 a_98299_n9675# VDD 1.27279f
C16 VDD I1N 1.34057f
C17 a_98299_n16810# VDD 1.03823f
C18 a_103997_n9675# VDD 1.27279f
C19 VDD VCM 6.7918f
C20 a_101641_n6960# VDD 1.18674f
C21 a_103997_n16810# VDD 1.04258f
C22 VDD IN_NEG 2.89387f
C23 a_107339_n6960# VDD 1.18674f
C24 a_109695_n9675# VDD 1.60209f
C25 a_109695_n16810# VDD 1.40063f
C26 a_113037_n6960# VDD 1.28333f
C27 a_81205_n21335# VDD 1.33016f
C28 a_84547_n18620# VDD 1.18674f
C29 a_86903_n21335# VDD 1.40049f
C30 a_92601_n5150# VDD 1.28138f
C31 VDD OUT 47.331f
C32 a_90245_n18620# VDD 1.18674f
C33 a_92601_n21335# VDD 1.40049f
C34 VDD IBNOUT 1.55863f
C35 a_98299_n5150# VDD 1.40049f
C36 a_95943_n18620# VDD 1.25121f
C37 VDD IBPOUT 3.44382f
C38 a_103997_n5150# VDD 1.40049f
C39 w_27790_n38888# VDD 96.053f
C40 VDD IN_POS 6.65925f
C41 a_109695_n5150# VDD 1.40049f
C42 IN_NEG VSS 50.44224f
C43 IN_POS VSS 38.26637f
C44 VCM VSS 16.767963f
C45 IBPOUT VSS 11.58886f
C46 I1N VSS 53.45688f
C47 IBNOUT VSS 9.23631f
C48 I1U VSS 33.7696f
C49 OUT VSS 44.56392f
C50 VDD VSS 10.164393p
C51 a_64243_n19597# VSS 1.20649f
C52 a_65677_n17803# VSS 1.46283f
C53 a_57977_n19597# VSS 1.20649f
C54 a_59411_n17803# VSS 1.45216f
C55 a_51711_n19597# VSS 1.20649f
C56 a_53145_n17803# VSS 1.45216f
C57 a_46879_n14213# VSS 1.45219f
C58 a_45445_n12419# VSS 1.14257f
C59 a_40613_n14213# VSS 1.45216f
C60 a_39179_n12419# VSS 1.10481f
C61 a_34347_n14213# VSS 1.29606f
C62 a_32913_n12419# VSS 1.14404f
C63 a_64243_n8932# VSS 1.10481f
C64 a_65677_n7138# VSS 1.28647f
C65 a_57977_n8932# VSS 1.10481f
C66 a_59411_n7138# VSS 1.45216f
C67 a_51711_n8932# VSS 1.13141f
C68 a_53145_n7138# VSS 1.28672f
C69 a_46879_n3548# VSS 1.28675f
C70 a_45445_n1754# VSS 1.20649f
C71 a_40613_n3548# VSS 1.45216f
C72 a_39179_n1754# VSS 1.20649f
C73 a_34347_n3548# VSS 1.45216f
C74 a_32913_n1754# VSS 1.20649f
C75 w_27790_n38888# VSS 0.430923p $ **FLOATING
C76 a_101111_n17715.t0 VSS 1.00448f
C77 IN_NEG.n0 VSS 2.14417f
C78 IN_NEG.n7 VSS 3.88312f
C79 IN_NEG.t1 VSS -11.2283f
C80 IN_NEG.n8 VSS 3.9473f
C81 IN_NEG.n9 VSS 1.12359f
C82 IN_NEG.n10 VSS 2.68065f
C83 IN_NEG.n13 VSS 1.8676f
C84 IN_NEG.n16 VSS 1.08259f
C85 IN_NEG.n22 VSS 1.06551f
C86 IN_NEG.n25 VSS 1.87274f
C87 IN_NEG.n27 VSS 2.63138f
C88 IN_NEG.n28 VSS 1.09392f
C89 IN_NEG.n29 VSS 2.1073f
C90 IN_NEG.t0 VSS 12.679f
C91 IN_NEG.n30 VSS 7.87284f
C92 a_84017_n16810.t1 VSS 1.00453f
C93 a_45445_n16007.t1 VSS 1.26793f
C94 a_45445_n16007.t0 VSS 1.23207f
C95 a_32913_n16007.t1 VSS 1.23207f
C96 a_32913_n16007.t0 VSS 1.26793f
C97 a_95413_n16810.t0 VSS 1.00448f
C98 a_112507_n6055.t0 VSS 1.00448f
C99 a_95413_n5150.t0 VSS 1.00448f
C100 a_106676_n27257.n0 VSS 9.95669f
C101 a_84017_n5150.t0 VSS 1.00448f
C102 a_71266_n4019.t0 VSS 21.298f
C103 a_71266_n4019.t2 VSS 14.601999f
C104 a_36008_n27257.n0 VSS 9.95669f
C105 a_57977_n16009.t1 VSS 1.26787f
C106 a_57977_n16009.t0 VSS 1.23213f
C107 a_64243_n16009.t1 VSS 1.26787f
C108 a_64243_n16009.t0 VSS 1.23213f
C109 a_43010_n36322.t2 VSS 3.08334f
C110 a_43010_n36322.t3 VSS 51.9824f
C111 a_43010_n36322.t1 VSS 1.84861f
C112 a_43010_n36322.t0 VSS 33.8856f
C113 a_45445_n5342.t1 VSS 1.26793f
C114 a_45445_n5342.t0 VSS 1.23207f
C115 a_53675_7563.n0 VSS 10.6245f
C116 a_112507_n17715.t0 VSS 1.00448f
C117 a_89009_n30339.n0 VSS 10.6245f
C118 a_36008_n30339.n0 VSS 10.6245f
C119 VCM.t2 VSS 3.82305f
C120 VCM.t3 VSS 2.11966f
C121 VCM.n0 VSS 4.64613f
C122 VCM.n1 VSS 3.62553f
C123 VCM.n2 VSS 5.40563f
C124 a_106809_n6055.t0 VSS 1.00448f
C125 a_39179_n5342.t1 VSS 1.26793f
C126 a_39179_n5342.t0 VSS 1.23207f
C127 a_89009_4481.n0 VSS 9.956611f
C128 a_64243_n5344.t1 VSS 1.26787f
C129 a_64243_n5344.t0 VSS 1.23213f
C130 a_89715_n5150.t1 VSS 1.00453f
C131 a_51711_n16009.t1 VSS 1.26787f
C132 a_51711_n16009.t0 VSS 1.23213f
C133 a_53675_n27257.n0 VSS 9.956639f
C134 a_89033_n36322.n0 VSS 8.139339f
C135 a_89033_n36322.n1 VSS 8.25763f
C136 a_94892_4481.t8 VSS 3.64456f
C137 a_94892_4481.n1 VSS 7.74464f
C138 IN_POS.n0 VSS 4.48494f
C139 IN_POS.n1 VSS 4.29823f
C140 IN_POS.n10 VSS 1.21126f
C141 IN_POS.n12 VSS 2.06759f
C142 IN_POS.n15 VSS 2.3333f
C143 IN_POS.n16 VSS 2.91269f
C144 IN_POS.n17 VSS 1.21105f
C145 IN_POS.n19 VSS 2.07287f
C146 IN_POS.n24 VSS 1.17853f
C147 IN_POS.n27 VSS 1.94474f
C148 IN_POS.n28 VSS 1.2439f
C149 IN_POS.n29 VSS 2.94329f
C150 IN_POS.t1 VSS -14.683901f
C151 IN_POS.n31 VSS 12.7299f
C152 IN_POS.n32 VSS 5.28104f
C153 a_101111_n6055.t1 VSS 1.00453f
C154 a_36032_13546.n0 VSS 7.9691f
C155 a_36032_13546.n1 VSS 8.089789f
C156 a_89009_7563.n0 VSS 10.6245f
C157 a_36008_7563.n0 VSS 10.6245f
C158 a_106830_n36382.n0 VSS 2.51436f
C159 a_106830_n36382.n1 VSS 9.83545f
C160 a_106830_n36382.n3 VSS 1.58916f
C161 a_106830_n36382.n4 VSS 5.82997f
C162 a_106830_n36382.n5 VSS 7.8766f
C163 a_106676_7563.n0 VSS 10.6245f
C164 a_39179_n8930.t1 VSS 59.5026f
C165 a_39179_n8930.t2 VSS 2.36783f
C166 a_39179_n8930.t0 VSS 30.229502f
C167 a_50629_n16009.t2 VSS 4.46728f
C168 a_50629_n16009.t1 VSS 50.2255f
C169 a_50629_n16009.t0 VSS 33.0072f
C170 a_71342_n27257.n0 VSS 9.95669f
C171 a_30324_5507.t1 VSS 34.531998f
C172 a_30324_5507.t2 VSS 1.63453f
C173 a_30324_5507.t0 VSS 16.5335f
C174 a_71366_n36322.n0 VSS 8.385951f
C175 a_71366_n36322.n1 VSS 8.26458f
C176 a_39179_n16007.t1 VSS 1.26793f
C177 a_39179_n16007.t0 VSS 1.23207f
C178 a_65658_n29313.t0 VSS 23.122198f
C179 a_65658_n29313.t1 VSS 8.80583f
C180 a_65658_n29313.t2 VSS 7.57194f
C181 a_32913_n5342.t1 VSS 1.23207f
C182 a_32913_n5342.t0 VSS 1.26793f
C183 a_36162_10388.n0 VSS 2.54961f
C184 a_36162_10388.n1 VSS 9.97333f
C185 a_36162_10388.n3 VSS 1.61144f
C186 a_36162_10388.n5 VSS 5.9117f
C187 a_36162_10388.n6 VSS 7.98701f
C188 a_53675_4481.n0 VSS 9.95668f
C189 a_38097_n16007.t1 VSS 6.98815f
C190 a_38097_n16007.t2 VSS 51.744198f
C191 a_38097_n16007.t0 VSS 24.7676f
C192 a_78344_10448.t1 VSS 60.4635f
C193 a_78344_10448.t0 VSS 27.6967f
C194 a_71366_11614.n0 VSS 11.663199f
C195 a_71366_11614.n1 VSS 4.27801f
C196 a_71366_11614.t1 VSS 5.09994f
C197 a_71366_11614.n2 VSS 53.2523f
C198 a_71366_11614.t0 VSS 19.8417f
C199 a_71342_7563.n0 VSS 10.6245f
C200 a_36162_n36382.n0 VSS 2.54373f
C201 a_36162_n36382.n1 VSS 9.950349f
C202 a_36162_n36382.n3 VSS 1.60773f
C203 a_36162_n36382.n4 VSS 5.89808f
C204 a_36162_n36382.n5 VSS 7.96862f
C205 a_71366_13546.n0 VSS 7.84506f
C206 a_71366_13546.n1 VSS 7.96027f
C207 a_89715_n16810.t1 VSS 1.00453f
C208 I1N.n31 VSS -6.14373f
C209 a_65658_4421.t0 VSS 25.151001f
C210 a_65658_4421.t2 VSS 13.2043f
C211 a_65658_4421.t1 VSS 1.14464f
C212 a_53699_11614.n0 VSS 11.7253f
C213 a_53699_11614.n1 VSS 4.30079f
C214 a_53699_11614.t1 VSS 5.1271f
C215 a_53699_11614.n2 VSS 49.478897f
C216 a_53699_11614.t0 VSS 23.3596f
C217 a_53699_13546.n0 VSS 8.0887f
C218 a_53699_13546.n1 VSS 7.97019f
C219 a_53829_10388.n0 VSS 2.53786f
C220 a_53829_10388.n1 VSS 9.92737f
C221 a_53829_10388.n3 VSS 1.60401f
C222 a_53829_10388.n4 VSS 5.88445f
C223 a_53829_10388.n5 VSS 7.950201f
C224 a_65486_11614.n1 VSS 11.477901f
C225 a_65486_11614.n2 VSS 11.550099f
C226 a_60677_n36322.t2 VSS 3.06439f
C227 a_60677_n36322.t1 VSS 57.1458f
C228 a_60677_n36322.t3 VSS 1.83725f
C229 a_60677_n36322.t0 VSS 28.752499f
C230 a_53675_n30339.n0 VSS 10.6245f
C231 a_59558_n29181.t0 VSS 3.64456f
C232 a_59558_n29181.n0 VSS 4.17871f
C233 a_59558_n29181.n1 VSS 4.01532f
C234 a_47991_n29313.t0 VSS 23.122198f
C235 a_47991_n29313.t1 VSS 8.80583f
C236 a_47991_n29313.t2 VSS 7.57194f
C237 a_48951_4481.t2 VSS 5.00668f
C238 a_48951_4481.t1 VSS 46.7297f
C239 a_48951_4481.t0 VSS 31.663698f
C240 a_47991_5507.t1 VSS 71.2991f
C241 a_47991_5507.t2 VSS 2.73325f
C242 a_47991_5507.t0 VSS 14.967599f
C243 a_103997_n8770.n0 VSS 11.0025f
C244 a_103997_n8770.n1 VSS 4.03565f
C245 a_103997_n8770.t1 VSS 3.70434f
C246 a_103997_n8770.n3 VSS 57.1449f
C247 a_103997_n8770.t0 VSS 25.2037f
C248 a_57977_n5344.t1 VSS 1.26787f
C249 a_57977_n5344.t0 VSS 1.23213f
C250 a_47991_4421.t0 VSS 25.151001f
C251 a_47991_4421.t1 VSS 13.2043f
C252 a_47991_4421.t2 VSS 1.14464f
C253 a_47819_11614.n1 VSS 11.477901f
C254 a_47819_11614.n2 VSS 11.550099f
C255 a_83153_10448.n0 VSS 7.87162f
C256 a_83153_10448.n1 VSS 12.123099f
C257 a_83153_n36322.n0 VSS 11.550099f
C258 a_83153_n36322.n2 VSS 11.477901f
C259 a_84017_n17715.t2 VSS 61.9764f
C260 a_84017_n17715.t0 VSS 34.5288f
C261 a_83325_4421.t0 VSS 25.151001f
C262 a_83325_4421.t1 VSS 13.2043f
C263 a_83325_4421.t2 VSS 1.14464f
C264 a_47819_n36322.n0 VSS 11.550099f
C265 a_47819_n36322.n2 VSS 11.477901f
C266 a_47819_10448.n0 VSS 7.87162f
C267 a_47819_10448.t9 VSS 13.622499f
C268 a_112559_n29181.n0 VSS 4.20259f
C269 a_112559_n29181.n1 VSS 4.03827f
C270 a_112559_n29181.t1 VSS 3.66539f
C271 a_30324_n29313.t0 VSS 23.414902f
C272 a_30324_n29313.t2 VSS 8.917299f
C273 a_30324_n29313.t1 VSS 7.66778f
C274 a_56895_n16009.t2 VSS 4.41403f
C275 a_56895_n16009.t1 VSS 46.3764f
C276 a_56895_n16009.t0 VSS 36.409603f
C277 a_83153_n35156.n0 VSS 7.87162f
C278 a_83153_n35156.t8 VSS 13.622499f
C279 a_89033_n35156.n0 VSS 11.033299f
C280 a_89033_n35156.n1 VSS 4.04697f
C281 a_89033_n35156.t3 VSS 3.71473f
C282 a_89033_n35156.n3 VSS 62.454002f
C283 a_89033_n35156.t0 VSS 19.6173f
C284 a_96011_n36322.t2 VSS 2.81139f
C285 a_96011_n36322.t0 VSS 2.07143f
C286 a_96011_n36322.t1 VSS 67.07571f
C287 a_96011_n36322.t3 VSS 27.041399f
C288 a_36008_4481.n0 VSS 9.956611f
C289 a_30152_11614.n1 VSS 11.5118f
C290 a_30152_11614.n2 VSS 11.584201f
C291 a_63161_n5344.t2 VSS 4.9628f
C292 a_63161_n5344.t1 VSS 49.1395f
C293 a_63161_n5344.t0 VSS 29.1977f
C294 a_64243_n1756.t1 VSS 69.347206f
C295 a_64243_n1756.t2 VSS 2.72276f
C296 a_64243_n1756.t0 VSS 16.93f
C297 a_77225_n29181.n0 VSS 4.17871f
C298 a_77225_n29181.n1 VSS 4.01532f
C299 a_77225_n29181.t2 VSS 3.64456f
C300 a_94892_n29181.n0 VSS 4.17871f
C301 a_94892_n29181.n1 VSS 4.01532f
C302 a_94892_n29181.t1 VSS 3.64456f
C303 a_83325_n29313.t0 VSS 23.122198f
C304 a_83325_n29313.t1 VSS 8.80583f
C305 a_83325_n29313.t2 VSS 7.57194f
C306 a_53699_n35156.t0 VSS 3.84924f
C307 a_53699_n35156.n0 VSS 11.7377f
C308 a_53699_n35156.n1 VSS 53.8229f
C309 a_53699_n35156.n2 VSS 4.30534f
C310 a_53699_n35156.t2 VSS 20.954401f
C311 a_59558_4481.n1 VSS 7.74464f
C312 a_59558_4481.t10 VSS 3.64456f
C313 a_39179_n19595.t0 VSS 72.542206f
C314 a_39179_n19595.t2 VSS 2.69368f
C315 a_39179_n19595.t1 VSS 13.8641f
C316 a_78344_n36322.t3 VSS 3.04902f
C317 a_78344_n36322.t2 VSS 61.7295f
C318 a_78344_n36322.t1 VSS 1.82803f
C319 a_78344_n36322.t0 VSS 24.293499f
C320 a_71366_n35156.n0 VSS 11.6917f
C321 a_71366_n35156.n1 VSS 4.28844f
C322 a_71366_n35156.t3 VSS 3.93638f
C323 a_71366_n35156.n3 VSS 57.0977f
C324 a_71366_n35156.t0 VSS 16.425098f
C325 a_44363_n16007.t1 VSS 6.93736f
C326 a_44363_n16007.t2 VSS 50.117397f
C327 a_44363_n16007.t0 VSS 26.445198f
C328 a_53699_n36322.n0 VSS 8.25899f
C329 a_53699_n36322.n1 VSS 8.13798f
C330 a_71496_n36382.n0 VSS 2.53786f
C331 a_71496_n36382.n1 VSS 9.92737f
C332 a_71496_n36382.n3 VSS 1.60401f
C333 a_71496_n36382.n4 VSS 5.88446f
C334 a_71496_n36382.n5 VSS 7.95021f
C335 a_89009_n27257.n0 VSS 9.95669f
C336 a_41891_n29181.t0 VSS 3.64456f
C337 a_41891_n29181.n0 VSS 4.17871f
C338 a_41891_n29181.n1 VSS 4.01532f
C339 a_106809_n5150.t0 VSS 1.82106f
C340 a_106809_n5150.t1 VSS 39.92f
C341 a_106809_n5150.t3 VSS 1.09181f
C342 a_106809_n5150.t2 VSS 21.6672f
C343 a_89163_n36382.n0 VSS 2.53786f
C344 a_89163_n36382.n1 VSS 9.92737f
C345 a_89163_n36382.n3 VSS 1.60401f
C346 a_89163_n36382.n4 VSS 5.88446f
C347 a_89163_n36382.n5 VSS 7.95021f
C348 a_81205_n14095.n0 VSS 10.8627f
C349 a_81205_n14095.n1 VSS 3.98441f
C350 a_81205_n14095.t1 VSS 4.74993f
C351 a_81205_n14095.n2 VSS 55.6066f
C352 a_81205_n14095.t0 VSS 26.1919f
C353 a_43010_10448.t0 VSS 51.9369f
C354 a_43010_10448.t3 VSS 36.6491f
C355 a_36032_11614.n0 VSS 11.817201f
C356 a_36032_11614.n1 VSS 4.3345f
C357 a_36032_11614.t1 VSS 5.16728f
C358 a_36032_11614.n2 VSS 44.9672f
C359 a_36032_11614.t0 VSS 27.941301f
C360 a_65486_10448.n0 VSS 7.87162f
C361 a_65486_10448.t10 VSS 13.622499f
C362 a_89033_13546.n0 VSS 7.84565f
C363 a_89033_13546.n1 VSS 7.959681f
C364 a_89163_10388.n0 VSS 2.53786f
C365 a_89163_10388.n1 VSS 9.92737f
C366 a_89163_10388.n3 VSS 1.60401f
C367 a_89163_10388.n5 VSS 5.88445f
C368 a_89163_10388.n6 VSS 7.950201f
C369 a_30152_n35156.t0 VSS 20.5853f
C370 a_30152_n35156.t3 VSS 1.77452f
C371 a_36032_n35156.n0 VSS 11.7943f
C372 a_36032_n35156.n1 VSS 4.32611f
C373 a_36032_n35156.t1 VSS 3.97095f
C374 a_36032_n35156.n3 VSS 47.1512f
C375 a_36032_n35156.t0 VSS 25.5144f
C376 a_106676_4481.n0 VSS 9.95668f
C377 a_106830_10388.n0 VSS 2.51436f
C378 a_106830_10388.n1 VSS 9.83545f
C379 a_106830_10388.n3 VSS 1.58916f
C380 a_106830_10388.n5 VSS 5.82997f
C381 a_106830_10388.n6 VSS 7.87659f
C382 a_77225_4481.t8 VSS 3.64456f
C383 a_77225_4481.n1 VSS 7.74464f
C384 a_100820_n35156.t0 VSS 20.5853f
C385 a_100820_n35156.t2 VSS 1.77452f
C386 a_51711_n12421.t0 VSS 63.9549f
C387 a_51711_n12421.t2 VSS 2.46089f
C388 a_51711_n12421.t1 VSS 26.9842f
C389 a_47819_n35156.t2 VSS 20.5853f
C390 a_47819_n35156.t11 VSS 1.77452f
C391 a_30152_n36322.n0 VSS 11.584201f
C392 a_30152_n36322.n2 VSS 11.5119f
C393 a_112559_4481.n1 VSS 7.78889f
C394 a_112559_4481.t9 VSS 3.66538f
C395 a_89715_n17715.t3 VSS 36.1964f
C396 a_89715_n17715.t0 VSS 26.2966f
C397 a_86903_n14095.n0 VSS 10.9263f
C398 a_86903_n14095.t0 VSS 55.2877f
C399 a_86903_n14095.n1 VSS 4.00774f
C400 a_86903_n14095.t2 VSS 32.2293f
C401 a_83153_11614.n1 VSS 11.477901f
C402 a_83153_11614.n2 VSS 11.550099f
C403 a_106676_n30339.n0 VSS 10.6245f
C404 a_100820_n36322.n0 VSS 11.550099f
C405 a_100820_n36322.n2 VSS 11.477901f
C406 a_65486_n35156.t8 VSS 20.5853f
C407 a_65486_n35156.t11 VSS 1.77452f
C408 a_33249_34067.n9 VSS 1.10607f
C409 a_33249_34067.n19 VSS 1.10607f
C410 a_33249_34067.n22 VSS 1.4803f
C411 a_33249_34067.n25 VSS 1.47288f
C412 a_33249_34067.n26 VSS 1.24188f
C413 a_33249_34067.n28 VSS 1.38796f
C414 a_33249_34067.n30 VSS 1.09797f
C415 a_33249_34067.n34 VSS 2.82575f
C416 a_33249_34067.n54 VSS 4.90658f
C417 a_33249_34067.n55 VSS 7.56734f
C418 a_33249_34067.n56 VSS 1.24177f
C419 a_33249_34067.n60 VSS 1.14141f
C420 a_33249_34067.n61 VSS 5.40296f
C421 a_33249_34067.n63 VSS 1.62793f
C422 a_33249_34067.n64 VSS 1.13624f
C423 a_33249_34067.n68 VSS 1.05092f
C424 a_33249_34067.n74 VSS 1.03839f
C425 a_33249_34067.n75 VSS 1.04549f
C426 a_33249_34067.n76 VSS 4.76973f
C427 a_33249_34067.n77 VSS 1.24553f
C428 a_33249_34067.n79 VSS 1.16921f
C429 a_33249_34067.n84 VSS 5.1877f
C430 a_33249_34067.n86 VSS 1.51427f
C431 a_33249_34067.n92 VSS 1.06142f
C432 a_33249_34067.n97 VSS 4.38744f
C433 a_33249_34067.n98 VSS 5.63217f
C434 a_33249_34067.n101 VSS 3.23788f
C435 a_33249_34067.n104 VSS 1.12528f
C436 a_33249_34067.n106 VSS 1.45399f
C437 a_33249_34067.n107 VSS 3.01461f
C438 a_33249_34067.n109 VSS 1.44297f
C439 a_33249_34067.n113 VSS 8.876969f
C440 a_33249_34067.n114 VSS 12.1615f
C441 a_33249_34067.n121 VSS 3.96945f
C442 a_33249_34067.n122 VSS 3.16582f
C443 a_33249_34067.n123 VSS 1.46267f
C444 a_33249_34067.n125 VSS 1.38796f
C445 a_33249_34067.n130 VSS 3.64644f
C446 a_33249_34067.n132 VSS 1.09797f
C447 a_33249_34067.n147 VSS 2.82575f
C448 a_33249_34067.n148 VSS 3.14342f
C449 a_33249_34067.n151 VSS 3.14342f
C450 a_33249_34067.n152 VSS 4.42596f
C451 a_33249_34067.n153 VSS 1.46262f
C452 a_33249_34067.n154 VSS 1.14136f
C453 a_33379_34007.n0 VSS 1.38521f
C454 a_33379_34007.t27 VSS 0.215533p
C455 a_33379_34007.n351 VSS 1.46779f
C456 a_60677_10448.t2 VSS 56.4126f
C457 a_60677_10448.t0 VSS 31.6335f
C458 a_71281_n10073.n0 VSS 3.63047f
C459 a_71281_n10073.n491 VSS 2.21256f
C460 a_71281_n10073.n783 VSS 2.36947f
C461 a_71281_n10073.n784 VSS 5.12344f
C462 a_45445_n19595.t1 VSS 68.227104f
C463 a_45445_n19595.t2 VSS 2.67562f
C464 a_45445_n19595.t0 VSS 18.1973f
C465 a_33379_34917.n0 VSS 3.81673f
C466 a_33379_34917.n1 VSS 1.71606f
C467 a_33379_34917.t0 VSS 1.07595f
C468 a_33379_34917.t68 VSS 0.221873p
C469 a_33379_34917.n9 VSS 1.76731f
C470 a_51711_n5344.t1 VSS 1.26787f
C471 a_51711_n5344.t0 VSS 1.23213f
C472 a_31831_n5342.t1 VSS 6.1634f
C473 a_31831_n5342.t2 VSS 48.951797f
C474 a_31831_n5342.t0 VSS 31.4848f
C475 a_32913_n8930.t1 VSS 63.4564f
C476 a_32913_n8930.t2 VSS 2.38382f
C477 a_32913_n8930.t0 VSS 26.3598f
C478 a_30152_10448.t3 VSS 20.5853f
C479 a_30152_10448.t1 VSS 1.77451f
C480 a_71342_4481.n0 VSS 9.956611f
C481 a_71496_10388.n0 VSS 2.53786f
C482 a_71496_10388.n1 VSS 9.92737f
C483 a_71496_10388.n3 VSS 1.60401f
C484 a_71496_10388.n4 VSS 5.88445f
C485 a_71496_10388.n5 VSS 7.950201f
C486 a_100992_4421.t0 VSS 25.151001f
C487 a_100992_4421.t1 VSS 13.2043f
C488 a_100992_4421.t2 VSS 1.14464f
C489 a_38097_n5342.t1 VSS 6.118411f
C490 a_38097_n5342.t2 VSS 45.5543f
C491 a_38097_n5342.t0 VSS 34.8273f
C492 a_100992_n29313.t0 VSS 23.122198f
C493 a_100992_n29313.t2 VSS 8.80583f
C494 a_100992_n29313.t1 VSS 7.57194f
C495 a_31284_n30339.t2 VSS 7.04722f
C496 a_31284_n30339.t1 VSS 49.8859f
C497 a_31284_n30339.t0 VSS 26.6669f
C498 a_30324_n30399.t1 VSS 45.1766f
C499 a_30324_n30399.t2 VSS 1.60691f
C500 a_30324_n30399.t0 VSS 6.01645f
C501 OUT.n11 VSS 1.93161f
C502 OUT.t109 VSS 7.241391f
C503 OUT.t108 VSS 10.055799f
C504 OUT.n12 VSS 21.947802f
C505 OUT.n13 VSS 20.055302f
C506 OUT.n14 VSS 40.5919f
C507 OUT.n15 VSS 1.90125f
C508 OUT.n17 VSS 1.13405f
C509 OUT.n19 VSS 1.13405f
C510 OUT.n20 VSS 1.17727f
C511 OUT.n29 VSS 2.86532f
C512 OUT.n57 VSS 2.62673f
C513 OUT.n76 VSS 1.66662f
C514 OUT.n77 VSS 1.61549f
C515 OUT.n82 VSS 1.78572f
C516 OUT.n115 VSS 1.93161f
C517 OUT.n116 VSS 2.24452f
C518 OUT.n117 VSS 5.82271f
C519 OUT.n135 VSS 3.11177f
C520 OUT.n137 VSS 1.31092f
C521 OUT.n138 VSS 2.17189f
C522 OUT.n139 VSS 2.93552f
C523 OUT.n140 VSS 2.98586f
C524 a_33249_48695.n20 VSS 1.77855f
C525 a_33249_48695.n21 VSS 1.25797f
C526 a_33249_48695.n22 VSS 1.19957f
C527 a_33249_48695.n23 VSS 1.77855f
C528 a_33249_48695.n24 VSS 1.25797f
C529 a_33249_48695.n26 VSS 1.70465f
C530 a_33249_48695.n27 VSS 1.49105f
C531 a_33249_48695.n29 VSS 1.70465f
C532 a_33249_48695.n30 VSS 1.49105f
C533 a_33249_48695.n38 VSS 1.18777f
C534 a_33249_48695.n39 VSS 1.05609f
C535 a_33249_48695.n45 VSS 1.18777f
C536 a_33249_48695.n51 VSS 2.69004f
C537 a_33249_48695.n52 VSS 1.06267f
C538 a_33249_48695.n66 VSS 3.12051f
C539 a_33249_48695.n71 VSS 2.09974f
C540 a_33249_48695.n76 VSS 2.10814f
C541 a_33249_48695.n77 VSS 2.64144f
C542 a_33249_48695.n80 VSS 1.18974f
C543 a_33249_48695.n85 VSS 2.52449f
C544 a_33249_48695.n86 VSS 2.89625f
C545 a_33249_48695.n89 VSS 2.49893f
C546 a_33249_48695.n90 VSS 1.39244f
C547 a_33249_48695.n106 VSS 1.49372f
C548 a_33249_48695.n108 VSS 1.70039f
C549 a_33249_48695.n109 VSS 1.7652f
C550 a_33249_48695.n110 VSS 3.93851f
C551 a_33249_48695.n129 VSS 4.29625f
C552 a_33249_48695.n132 VSS 1.25177f
C553 a_33249_48695.n133 VSS 2.87631f
C554 a_33249_48695.n134 VSS 2.6775f
C555 a_33249_48695.n137 VSS 1.49372f
C556 a_33249_48695.n139 VSS 1.70039f
C557 a_33249_48695.n140 VSS 1.25245f
C558 a_33249_48695.n141 VSS 2.42226f
C559 a_33249_48695.n174 VSS 2.89625f
C560 a_33249_48695.n175 VSS 2.84854f
C561 a_33249_48695.n176 VSS 1.25177f
C562 a_33249_48695.n177 VSS 3.2993f
C563 a_33249_48695.n178 VSS 2.73275f
C564 a_33249_48695.n179 VSS 3.19912f
C565 a_33249_48695.n183 VSS 1.78511f
C566 a_33249_48695.n185 VSS 4.43096f
C567 a_33249_48695.n218 VSS 3.8908f
C568 a_33249_48695.n221 VSS 1.24524f
C569 a_33249_48695.n223 VSS 1.78417f
C570 a_33249_48695.n224 VSS 1.25132f
C571 a_33249_48695.n225 VSS 2.79169f
C572 a_33249_48695.n226 VSS 2.50126f
C573 a_33249_48695.n227 VSS 1.25252f
C574 a_33249_48695.n228 VSS 2.77274f
C575 a_33249_48695.n261 VSS 2.54509f
C576 a_33249_48695.n262 VSS 3.86208f
C577 a_33249_48695.n265 VSS 1.24524f
C578 a_33249_48695.n267 VSS 1.78417f
C579 a_33249_48695.n268 VSS 1.25132f
C580 a_33249_48695.n269 VSS 3.1335f
C581 a_33249_48695.n270 VSS 2.00968f
C582 a_33249_48695.n271 VSS 2.08409f
C583 a_33249_48695.n272 VSS 2.79169f
C584 a_33249_48695.n283 VSS 1.02196f
C585 a_33249_48695.n285 VSS 1.17271f
C586 a_33249_48695.n294 VSS 1.13487f
C587 a_33249_48695.n295 VSS 3.83834f
C588 a_33249_48695.n296 VSS 1.25143f
C589 a_33249_48695.n300 VSS 1.08733f
C590 a_33249_48695.n303 VSS 4.22418f
C591 a_33249_48695.n306 VSS 1.18974f
C592 a_33249_48695.n320 VSS 2.81996f
C593 a_33249_48695.n321 VSS 2.71764f
C594 a_33249_48695.n323 VSS 2.6883f
C595 a_33249_48695.n326 VSS 1.02196f
C596 a_33249_48695.n328 VSS 1.17271f
C597 a_33249_48695.n334 VSS 1.08733f
C598 a_33249_48695.n335 VSS 1.25143f
C599 a_33249_48695.n336 VSS 2.33745f
C600 a_33249_48695.n337 VSS 3.07641f
C601 a_33249_48695.n347 VSS 3.43055f
C602 a_33249_48695.n348 VSS 2.84218f
C603 a_33249_48695.n349 VSS 3.04283f
C604 a_33249_48695.n352 VSS 3.0578f
C605 a_33249_48695.n353 VSS 1.06267f
C606 a_33249_48695.n363 VSS 1.18777f
C607 a_33249_48695.n364 VSS 1.2517f
C608 a_33249_48695.n365 VSS 2.70921f
C609 a_33249_48695.n366 VSS 2.41819f
C610 a_33249_48695.n379 VSS 2.41819f
C611 a_33249_48695.n386 VSS 2.69004f
C612 a_33249_48695.n387 VSS 4.1989f
C613 a_33249_48695.n393 VSS 1.18777f
C614 a_33249_48695.n394 VSS 1.2517f
C615 a_33249_48695.n395 VSS 3.7876f
C616 a_106809_n17715.t1 VSS 1.00453f
C617 a_71342_n30339.n0 VSS 10.6245f
C618 a_65486_n36322.n0 VSS 11.550099f
C619 a_65486_n36322.n2 VSS 11.477901f
C620 a_52635_48695.n1 VSS 1.21873f
C621 a_52635_48695.n2 VSS 1.21872f
C622 a_52635_48695.n3 VSS 1.18681f
C623 a_52635_48695.n5 VSS 1.21873f
C624 a_52635_48695.n6 VSS 1.71719f
C625 a_52635_48695.n7 VSS 1.52681f
C626 a_52635_48695.n8 VSS 1.21873f
C627 a_52635_48695.n9 VSS 1.21872f
C628 a_52635_48695.n10 VSS 1.18681f
C629 a_52635_48695.n12 VSS 1.21873f
C630 a_52635_48695.n13 VSS 1.71719f
C631 a_52635_48695.n14 VSS 1.2057f
C632 a_52635_48695.n15 VSS 1.0473f
C633 a_52635_48695.n16 VSS 1.14869f
C634 a_52635_48695.n18 VSS 1.16549f
C635 a_52635_48695.n19 VSS 1.16549f
C636 a_52635_48695.n21 VSS 1.0473f
C637 a_52635_48695.n22 VSS 1.14869f
C638 a_52635_48695.n23 VSS 1.36844f
C639 a_52635_48695.n24 VSS 1.2057f
C640 a_52635_48695.n25 VSS 1.0473f
C641 a_52635_48695.n26 VSS 1.14869f
C642 a_52635_48695.n28 VSS 1.16549f
C643 a_52635_48695.n29 VSS 1.16549f
C644 a_52635_48695.n31 VSS 1.0473f
C645 a_52635_48695.n32 VSS 1.14869f
C646 a_52635_48695.n33 VSS 1.36844f
C647 a_52635_48695.n35 VSS 1.21985f
C648 a_52635_48695.n38 VSS 1.72003f
C649 a_52635_48695.n40 VSS 1.21988f
C650 a_52635_48695.n43 VSS 6.43054f
C651 a_52635_48695.n44 VSS 3.88654f
C652 a_52635_48695.n47 VSS 1.47747f
C653 a_52635_48695.n49 VSS 1.69542f
C654 a_52635_48695.n50 VSS 4.5114f
C655 a_52635_48695.n52 VSS 3.88906f
C656 a_52635_48695.n54 VSS 1.35842f
C657 a_52635_48695.n55 VSS 1.14974f
C658 a_52635_48695.n56 VSS 1.04175f
C659 a_52635_48695.n58 VSS 1.21146f
C660 a_52635_48695.n60 VSS 1.21146f
C661 a_52635_48695.n62 VSS 1.53633f
C662 a_52635_48695.n66 VSS 1.41217f
C663 a_52635_48695.n68 VSS 1.35842f
C664 a_52635_48695.n69 VSS 1.14974f
C665 a_52635_48695.n70 VSS 1.04175f
C666 a_52635_48695.n71 VSS 1.04175f
C667 a_52635_48695.n72 VSS 1.14974f
C668 a_52635_48695.n75 VSS 1.157f
C669 a_52635_48695.n76 VSS 1.16648f
C670 a_52635_48695.n80 VSS 5.47584f
C671 a_52635_48695.n81 VSS 1.80962f
C672 a_52635_48695.n83 VSS 1.71719f
C673 a_52635_48695.n87 VSS 1.12283f
C674 a_52635_48695.n88 VSS 6.07046f
C675 a_52635_48695.n95 VSS 3.88906f
C676 a_52635_48695.n96 VSS 3.49604f
C677 a_52635_48695.n98 VSS 1.04175f
C678 a_52635_48695.n99 VSS 1.14974f
C679 a_52635_48695.n102 VSS 1.157f
C680 a_52635_48695.n103 VSS 1.16648f
C681 a_52635_48695.n107 VSS 3.49604f
C682 a_52635_48695.n108 VSS 1.53633f
C683 a_52635_48695.n112 VSS 1.41217f
C684 a_52635_48695.n116 VSS 1.12283f
C685 a_52635_48695.n118 VSS 1.71719f
C686 a_52635_48695.n119 VSS 1.80962f
C687 a_52635_48695.n120 VSS 3.91678f
C688 a_52635_48695.n121 VSS 4.55814f
C689 a_52635_48695.n127 VSS 4.10938f
C690 a_52635_48695.n128 VSS 6.28374f
C691 a_52635_48695.n130 VSS 1.21988f
C692 a_52635_48695.n133 VSS 5.24514f
C693 a_52635_48695.n134 VSS 6.10701f
C694 a_52635_48695.n137 VSS 1.72003f
C695 a_52635_48695.n139 VSS 1.21988f
C696 a_52635_48695.n150 VSS 1.64071f
C697 a_52635_48695.n153 VSS 1.47747f
C698 a_52635_48695.n155 VSS 1.69542f
C699 a_52635_48695.n157 VSS 1.02404f
C700 a_52635_48695.n161 VSS 1.57198f
C701 a_52635_48695.n162 VSS 1.80922f
C702 a_52635_48695.n163 VSS 5.54919f
C703 a_52635_48695.n164 VSS 4.03603f
C704 a_52635_48695.n167 VSS 1.1884f
C705 a_52635_48695.n169 VSS 1.21985f
C706 a_52635_48695.n171 VSS 1.21988f
C707 a_52635_48695.n174 VSS 4.07689f
C708 a_52635_48695.n184 VSS 3.92896f
C709 a_52635_48695.n185 VSS 3.8188f
C710 a_52635_48695.n187 VSS 1.02404f
C711 a_52635_48695.n191 VSS 1.57198f
C712 a_52635_48695.n192 VSS 1.80922f
C713 a_52635_48695.n193 VSS 3.37931f
C714 a_52635_48695.n194 VSS 4.6906f
C715 a_52635_48695.n196 VSS 1.1884f
C716 a_35922_19591.n0 VSS 4.07049f
C717 a_35922_19591.n31 VSS 1.84527f
C718 a_35922_19591.n34 VSS 1.84527f
C719 a_35922_19591.n39 VSS 1.84527f
C720 a_35922_19591.n43 VSS 1.84527f
C721 a_35922_19591.n48 VSS 1.8766f
C722 a_35922_19591.n50 VSS 1.88001f
C723 a_35922_19591.n54 VSS 1.8766f
C724 a_35922_19591.n56 VSS 1.88001f
C725 a_35922_19591.n63 VSS 4.32896f
C726 a_35922_19591.n64 VSS 1.31313f
C727 a_35922_19591.n66 VSS 1.31313f
C728 a_35922_19591.n68 VSS 1.31313f
C729 a_35922_19591.n70 VSS 1.31313f
C730 a_35922_19591.n72 VSS 1.78373f
C731 a_35922_19591.n74 VSS 1.78373f
C732 a_35922_19591.n76 VSS 1.37036f
C733 a_35922_19591.n78 VSS 1.37036f
C734 a_35922_19591.n80 VSS 1.37036f
C735 a_35922_19591.n82 VSS 1.37036f
C736 a_35922_19591.n84 VSS 1.80279f
C737 a_35922_19591.n86 VSS 1.80279f
C738 a_35922_19591.n90 VSS 1.78304f
C739 a_35922_19591.n91 VSS 1.78304f
C740 a_35922_19591.n93 VSS 1.01659f
C741 a_35922_19591.n94 VSS 1.79407f
C742 a_35922_19591.n99 VSS 1.79407f
C743 a_35922_19591.n127 VSS 2.45557f
C744 a_35922_19591.n128 VSS 2.42356f
C745 a_35922_19591.n139 VSS 1.02835f
C746 a_35922_19591.n163 VSS 3.64752f
C747 a_35922_19591.n208 VSS 3.64752f
C748 a_35922_19591.n214 VSS 2.42356f
C749 a_35922_19591.n215 VSS 2.42356f
C750 a_35922_19591.n216 VSS 3.78794f
C751 a_35922_19591.n217 VSS 3.78794f
C752 a_35922_19591.n218 VSS 2.42356f
C753 a_35922_19591.n219 VSS 2.03211f
C754 a_35922_19591.n221 VSS 2.26597f
C755 a_35922_19591.n222 VSS 2.92955f
C756 a_35922_19591.n223 VSS 2.13722f
C757 a_35922_19591.n229 VSS 2.13722f
C758 a_35922_19591.n230 VSS 8.488879f
C759 a_35922_19591.n237 VSS 10.4498f
C760 a_35922_19591.n239 VSS 3.23651f
C761 a_71281_n8397.n0 VSS 1.83357f
C762 a_71281_n8397.n1 VSS 5.784431f
C763 a_71281_n8397.n292 VSS 2.23771f
C764 a_71281_n8397.n584 VSS 2.75402f
C765 a_71281_n8397.n585 VSS 8.049689f
C766 a_41891_4481.t0 VSS 3.64456f
C767 a_41891_4481.n1 VSS 7.74464f
C768 a_35502_24538.n79 VSS 2.41886f
C769 a_35502_24538.n129 VSS 2.23998f
C770 a_35502_24538.n130 VSS 4.67369f
C771 a_35502_24538.n131 VSS 4.46256f
C772 a_35502_24538.n132 VSS 2.59861f
C773 a_31699_20742.n83 VSS 1.05167f
C774 a_31699_20742.n86 VSS 1.07804f
C775 a_31699_20742.n87 VSS 1.05555f
C776 a_31699_20742.n90 VSS 2.03605f
C777 a_31699_20742.n92 VSS 1.07804f
C778 a_31699_20742.n93 VSS 1.05167f
C779 a_31699_20742.n96 VSS 1.07804f
C780 a_31699_20742.n97 VSS 1.05555f
C781 a_31699_20742.n100 VSS 2.03605f
C782 a_31699_20742.n102 VSS 1.07386f
C783 a_31699_20742.n103 VSS 1.0203f
C784 a_31699_20742.n106 VSS 1.07386f
C785 a_31699_20742.n107 VSS 1.0203f
C786 a_31699_20742.n110 VSS 1.0203f
C787 a_31699_20742.n113 VSS 1.0203f
C788 a_31699_20742.n121 VSS 1.07386f
C789 a_31699_20742.n124 VSS 1.07386f
C790 a_31699_20742.n127 VSS 1.07386f
C791 a_31699_20742.n131 VSS 1.07386f
C792 a_31699_20742.n134 VSS 1.00324f
C793 a_31699_20742.n136 VSS 1.00324f
C794 a_31699_20742.n153 VSS 1.07804f
C795 a_31699_20742.n159 VSS 1.07804f
C796 a_31699_20742.n162 VSS 1.07804f
C797 a_31699_20742.n165 VSS 1.0203f
C798 a_31699_20742.n168 VSS 1.0203f
C799 a_31699_20742.n173 VSS 1.02306f
C800 a_31699_20742.n176 VSS 1.02306f
C801 a_31699_20742.n179 VSS 1.02306f
C802 a_31699_20742.n182 VSS 1.02306f
C803 a_31699_20742.n197 VSS 1.06707f
C804 a_31699_20742.n198 VSS 1.06813f
C805 a_31699_20742.n201 VSS 1.06813f
C806 a_31699_20742.n204 VSS 1.06813f
C807 a_31699_20742.n206 VSS 1.06813f
C808 a_31699_20742.n208 VSS 1.04026f
C809 a_31699_20742.n209 VSS 2.17076f
C810 a_31699_20742.n237 VSS 1.07595f
C811 a_31699_20742.n251 VSS 3.58253f
C812 a_31699_20742.n252 VSS 2.7071f
C813 a_31699_20742.n253 VSS 2.75045f
C814 a_31699_20742.n254 VSS 4.29884f
C815 a_31699_20742.n256 VSS 4.29884f
C816 a_31699_20742.n258 VSS 2.75045f
C817 a_31699_20742.n259 VSS 2.75045f
C818 a_31699_20742.n265 VSS 1.06707f
C819 a_31699_20742.n280 VSS 4.13948f
C820 a_31699_20742.n288 VSS 4.13948f
C821 a_31699_20742.n296 VSS 2.75045f
C822 a_31699_20742.n297 VSS 2.49429f
C823 a_31699_20742.n308 VSS 2.74435f
C824 a_31699_20742.n309 VSS 3.41548f
C825 a_31699_20742.n310 VSS 2.37271f
C826 a_31699_20742.n312 VSS 2.37271f
C827 a_31699_20742.n313 VSS 16.538599f
C828 a_31699_20742.n334 VSS 1.54854f
C829 a_31699_20742.n345 VSS 1.03208f
C830 a_31699_20742.n388 VSS 13.563499f
C831 a_31699_20742.t0 VSS 1.11866f
C832 a_31699_20742.n389 VSS 3.50557f
C833 a_31699_20742.n390 VSS 2.18128f
C834 a_31953_n19727.n321 VSS 1.21075f
C835 a_33249_35053.n0 VSS 1.83524f
C836 a_33249_35053.n1 VSS 1.4665f
C837 a_33249_35053.n2 VSS 1.57152f
C838 a_33249_35053.n3 VSS 1.92894f
C839 a_33249_35053.n4 VSS 1.68723f
C840 a_33249_35053.n5 VSS 1.08952f
C841 a_33249_35053.n6 VSS 1.92894f
C842 a_33249_35053.n7 VSS 1.68723f
C843 a_33249_35053.n8 VSS 1.08952f
C844 a_33249_35053.n9 VSS 2.09988f
C845 a_33249_35053.n10 VSS 4.85677f
C846 a_33249_35053.n14 VSS 7.50995f
C847 a_33249_35053.n15 VSS 3.02979f
C848 a_33249_35053.n30 VSS 4.45672f
C849 a_33249_35053.n32 VSS 1.92412f
C850 a_33249_35053.n33 VSS 1.99746f
C851 a_33249_35053.n35 VSS 1.69025f
C852 a_33249_35053.n36 VSS 1.57565f
C853 a_33249_35053.n69 VSS 4.86153f
C854 a_33249_35053.n70 VSS 3.25477f
C855 a_33249_35053.n73 VSS 1.41648f
C856 a_33249_35053.n74 VSS 2.82773f
C857 a_33249_35053.n75 VSS 1.11142f
C858 a_33249_35053.n77 VSS 1.69025f
C859 a_33249_35053.n79 VSS 1.92412f
C860 a_33249_35053.n80 VSS 1.41725f
C861 a_33249_35053.n81 VSS 2.74097f
C862 a_33249_35053.n82 VSS 3.27733f
C863 a_33249_35053.n101 VSS 3.27733f
C864 a_33249_35053.n104 VSS 1.41648f
C865 a_33249_35053.n105 VSS 4.42321f
C866 a_33249_35053.n106 VSS 12.737201f
C867 a_33249_35053.n108 VSS 2.09739f
C868 a_33249_35053.n109 VSS 9.46617f
C869 a_33249_35053.n121 VSS 2.86645f
C870 a_33249_35053.n123 VSS 3.53981f
C871 a_33249_35053.n124 VSS 5.24967f
C872 a_33249_35053.n126 VSS 1.84327f
C873 a_33249_35053.n127 VSS 1.20691f
C874 a_33249_35053.n129 VSS 1.48873f
C875 a_33249_35053.n130 VSS 1.06366f
C876 a_33249_35053.n131 VSS 4.2966f
C877 a_33249_35053.n133 VSS 5.31934f
C878 a_33249_35053.n155 VSS 4.69303f
C879 a_33249_35053.n156 VSS 1.94054f
C880 a_35502_25545.n143 VSS 1.05169f
C881 a_35502_25545.n210 VSS 1.68497f
C882 a_35502_25545.n220 VSS 1.79682f
C883 a_35502_25545.n221 VSS 1.28081f
C884 a_35502_25545.n272 VSS 1.66281f
C885 a_35502_25545.n325 VSS 1.66281f
C886 a_35502_25545.n326 VSS 2.38102f
C887 a_35502_25545.n341 VSS 2.05391f
C888 a_35502_25545.n342 VSS 3.03378f
C889 a_36032_n36322.n0 VSS 8.13687f
C890 a_36032_n36322.n1 VSS 8.260099f
C891 a_53829_n36382.n0 VSS 2.53786f
C892 a_53829_n36382.n1 VSS 9.92737f
C893 a_53829_n36382.n3 VSS 1.60401f
C894 a_53829_n36382.n4 VSS 5.88446f
C895 a_53829_n36382.n5 VSS 7.95021f
C896 a_100820_10448.n0 VSS 7.87162f
C897 a_100820_10448.t0 VSS 13.622499f
C898 a_31284_4481.t1 VSS 5.04925f
C899 a_31284_4481.t2 VSS 40.732197f
C900 a_31284_4481.t0 VSS 37.7185f
C901 a_30324_4421.t0 VSS 25.4694f
C902 a_30324_4421.t1 VSS 13.3715f
C903 a_30324_4421.t2 VSS 1.15913f
C904 a_100820_11614.n1 VSS 11.477901f
C905 a_100820_11614.n2 VSS 11.550099f
C906 a_57977_n12421.t0 VSS 59.2863f
C907 a_57977_n12421.t2 VSS 2.43373f
C908 a_57977_n12421.t1 VSS 31.18f
C909 a_52635_49681.n0 VSS 2.5012f
C910 a_52635_49681.n1 VSS 2.18773f
C911 a_52635_49681.n2 VSS 2.5012f
C912 a_52635_49681.n3 VSS 2.18779f
C913 a_52635_49681.n4 VSS 1.41275f
C914 a_52635_49681.n5 VSS 2.60963f
C915 a_52635_49681.n6 VSS 1.8458f
C916 a_52635_49681.n7 VSS 1.76011f
C917 a_52635_49681.n8 VSS 2.60963f
C918 a_52635_49681.n9 VSS 1.8458f
C919 a_52635_49681.n10 VSS 1.34268f
C920 a_52635_49681.n11 VSS 1.41272f
C921 a_52635_49681.n13 VSS 5.77891f
C922 a_52635_49681.n14 VSS 4.24962f
C923 a_52635_49681.n16 VSS 2.49496f
C924 a_52635_49681.n17 VSS 2.59005f
C925 a_52635_49681.n19 VSS 2.1917f
C926 a_52635_49681.n20 VSS 2.0431f
C927 a_52635_49681.n21 VSS 1.03037f
C928 a_52635_49681.n26 VSS 1.02935f
C929 a_52635_49681.n53 VSS 6.30381f
C930 a_52635_49681.n54 VSS 4.22046f
C931 a_52635_49681.n55 VSS 6.23036f
C932 a_52635_49681.n58 VSS 3.70414f
C933 a_52635_49681.n59 VSS 4.69402f
C934 a_52635_49681.n63 VSS 2.61926f
C935 a_52635_49681.n65 VSS 6.50148f
C936 a_52635_49681.n73 VSS 1.04211f
C937 a_52635_49681.n77 VSS 1.04214f
C938 a_52635_49681.n81 VSS 1.02776f
C939 a_52635_49681.n88 VSS 1.34555f
C940 a_52635_49681.n92 VSS 1.04211f
C941 a_52635_49681.n98 VSS 5.7089f
C942 a_52635_49681.n100 VSS 1.41191f
C943 a_52635_49681.n101 VSS 1.82711f
C944 a_52635_49681.n103 VSS 2.61788f
C945 a_52635_49681.n104 VSS 1.83604f
C946 a_52635_49681.n105 VSS 4.09621f
C947 a_52635_49681.n106 VSS 3.67005f
C948 a_52635_49681.n107 VSS 1.83781f
C949 a_52635_49681.n108 VSS 4.06839f
C950 a_52635_49681.n115 VSS 1.34555f
C951 a_52635_49681.n119 VSS 1.04211f
C952 a_52635_49681.n128 VSS 1.02776f
C953 a_52635_49681.n132 VSS 1.04214f
C954 a_52635_49681.n136 VSS 1.04211f
C955 a_52635_49681.n141 VSS 3.73436f
C956 a_52635_49681.n142 VSS 5.4662f
C957 a_52635_49681.n144 VSS 1.41191f
C958 a_52635_49681.n145 VSS 1.82711f
C959 a_52635_49681.n147 VSS 2.61788f
C960 a_52635_49681.n148 VSS 1.83604f
C961 a_52635_49681.n149 VSS 4.41262f
C962 a_52635_49681.n150 VSS 6.29237f
C963 a_52635_49681.n151 VSS 4.92683f
C964 a_52635_49681.n152 VSS 1.8367f
C965 a_52635_49681.n153 VSS 5.00434f
C966 a_52635_49681.n154 VSS 1.03037f
C967 a_52635_49681.n159 VSS 1.02935f
C968 a_52635_49681.n186 VSS 4.24962f
C969 a_52635_49681.n187 VSS 3.92865f
C970 a_52635_49681.n188 VSS 1.44115f
C971 a_52635_49681.n190 VSS 2.1917f
C972 a_52635_49681.n192 VSS 2.49496f
C973 a_52635_49681.n193 VSS 1.8377f
C974 a_52635_49681.n194 VSS 3.55414f
C975 a_52635_49681.n195 VSS 3.66664f
C976 a_52635_49681.n196 VSS 1.8367f
C977 VDD.n6 VSS 2.53555f
C978 VDD.n7 VSS 1.05204f
C979 VDD.n13 VSS 1.05032f
C980 VDD.t833 VSS 1.45905f
C981 VDD.t1481 VSS 1.96535f
C982 VDD.t538 VSS 1.96535f
C983 VDD.t536 VSS 1.36987f
C984 VDD.t1218 VSS 1.45794f
C985 VDD.t1570 VSS 1.96535f
C986 VDD.t1290 VSS 1.96535f
C987 VDD.t1540 VSS 1.36987f
C988 VDD.t845 VSS 1.31955f
C989 VDD.t1904 VSS 1.96535f
C990 VDD.t1155 VSS 1.96535f
C991 VDD.t1884 VSS 1.45794f
C992 VDD.t635 VSS 1.45794f
C993 VDD.t625 VSS 1.96535f
C994 VDD.t1996 VSS 1.96535f
C995 VDD.t2240 VSS 1.36987f
C996 VDD.t1424 VSS 1.45794f
C997 VDD.t1653 VSS 1.96535f
C998 VDD.t550 VSS 1.96535f
C999 VDD.t549 VSS 1.36987f
C1000 VDD.t547 VSS 1.31955f
C1001 VDD.t548 VSS 1.96535f
C1002 VDD.t828 VSS 1.96535f
C1003 VDD.t619 VSS 1.45794f
C1004 VDD.t1052 VSS 1.45794f
C1005 VDD.t1787 VSS 1.96535f
C1006 VDD.t501 VSS 1.96535f
C1007 VDD.t2382 VSS 1.36987f
C1008 VDD.t1127 VSS 1.45794f
C1009 VDD.t432 VSS 3.20156f
C1010 VDD.t423 VSS 7.65735f
C1011 VDD.t427 VSS 7.734359f
C1012 VDD.t472 VSS 9.533171f
C1013 VDD.t683 VSS 7.54182f
C1014 VDD.n690 VSS 3.54262f
C1015 VDD.t470 VSS 9.533171f
C1016 VDD.t742 VSS 7.54182f
C1017 VDD.n709 VSS 3.4106f
C1018 VDD.t429 VSS 7.65735f
C1019 VDD.t313 VSS 3.20156f
C1020 VDD.t320 VSS 7.65735f
C1021 VDD.t310 VSS 9.533171f
C1022 VDD.t574 VSS 7.54182f
C1023 VDD.n763 VSS 3.58663f
C1024 VDD.t557 VSS 7.54182f
C1025 VDD.t563 VSS 7.54182f
C1026 VDD.t471 VSS 9.533171f
C1027 VDD.t656 VSS 7.54182f
C1028 VDD.n874 VSS 3.4106f
C1029 VDD.t316 VSS 9.533171f
C1030 VDD.t314 VSS 7.734359f
C1031 VDD.t318 VSS 3.20156f
C1032 VDD.n1084 VSS 3.4106f
C1033 VDD.t700 VSS 7.54182f
C1034 VDD.t315 VSS 9.533171f
C1035 VDD.t341 VSS 7.734359f
C1036 VDD.t319 VSS 3.18057f
C1037 VDD.t312 VSS 7.65735f
C1038 VDD.t306 VSS 9.533171f
C1039 VDD.t653 VSS 7.54182f
C1040 VDD.t309 VSS 7.734359f
C1041 VDD.t311 VSS 9.533171f
C1042 VDD.t661 VSS 7.54182f
C1043 VDD.n1345 VSS 3.4106f
C1044 VDD.n1346 VSS 3.4106f
C1045 VDD.n1349 VSS 3.12105f
C1046 VDD.n1354 VSS 3.4106f
C1047 VDD.t818 VSS 7.54182f
C1048 VDD.t307 VSS 9.533171f
C1049 VDD.t317 VSS 7.65735f
C1050 VDD.n1356 VSS 3.12455f
C1051 VDD.t469 VSS 9.533171f
C1052 VDD.t434 VSS 7.65735f
C1053 VDD.n1414 VSS 3.12455f
C1054 VDD.t444 VSS 3.20156f
C1055 VDD.t439 VSS 7.734359f
C1056 VDD.t474 VSS 9.533171f
C1057 VDD.t878 VSS 7.54182f
C1058 VDD.n1415 VSS 3.4106f
C1059 VDD.n1428 VSS 3.4106f
C1060 VDD.n1429 VSS 3.4106f
C1061 VDD.n1442 VSS 1.16761f
C1062 VDD.n1480 VSS 1.50435f
C1063 VDD.n1521 VSS 1.52188f
C1064 VDD.n1549 VSS 1.52159f
C1065 VDD.t920 VSS 3.32223f
C1066 VDD.t1665 VSS 3.93704f
C1067 VDD.t692 VSS 2.74191f
C1068 VDD.t2299 VSS 3.32223f
C1069 VDD.t994 VSS 3.93704f
C1070 VDD.t1188 VSS 2.7319f
C1071 VDD.n1551 VSS 2.04987f
C1072 VDD.n1610 VSS 1.50435f
C1073 VDD.n1652 VSS 3.12455f
C1074 VDD.n1718 VSS 3.12105f
C1075 VDD.t442 VSS 3.18057f
C1076 VDD.t425 VSS 7.734359f
C1077 VDD.t468 VSS 9.533171f
C1078 VDD.t689 VSS 7.54182f
C1079 VDD.n1719 VSS 3.4106f
C1080 VDD.n1742 VSS 3.12455f
C1081 VDD.n1761 VSS 2.45645f
C1082 VDD.n1762 VSS 1.92254f
C1083 VDD.n1771 VSS 1.05032f
C1084 VDD.t965 VSS 1.45905f
C1085 VDD.t1099 VSS 1.96535f
C1086 VDD.t338 VSS 1.96535f
C1087 VDD.t335 VSS 1.36987f
C1088 VDD.t336 VSS 1.31955f
C1089 VDD.t337 VSS 1.96535f
C1090 VDD.t1419 VSS 1.96535f
C1091 VDD.t1642 VSS 1.45794f
C1092 VDD.t852 VSS 1.45794f
C1093 VDD.t2485 VSS 1.96535f
C1094 VDD.t322 VSS 1.96535f
C1095 VDD.t298 VSS 1.36987f
C1096 VDD.t789 VSS 1.45794f
C1097 VDD.t917 VSS 1.96535f
C1098 VDD.t500 VSS 1.96535f
C1099 VDD.t499 VSS 1.36987f
C1100 VDD.t498 VSS 1.31955f
C1101 VDD.t497 VSS 1.96535f
C1102 VDD.t2777 VSS 1.96535f
C1103 VDD.t1142 VSS 1.45794f
C1104 VDD.t1658 VSS 1.45794f
C1105 VDD.t801 VSS 1.96535f
C1106 VDD.t643 VSS 1.96535f
C1107 VDD.t1442 VSS 1.36987f
C1108 VDD.t855 VSS 1.45794f
C1109 VDD.t2118 VSS 1.96535f
C1110 VDD.t1841 VSS 1.96535f
C1111 VDD.t571 VSS 1.36987f
C1112 VDD.t3570 VSS 1.31955f
C1113 VDD.t2924 VSS 1.96535f
C1114 VDD.t1183 VSS 1.96535f
C1115 VDD.t905 VSS 1.45794f
C1116 VDD.t1936 VSS 1.45794f
C1117 VDD.t875 VSS 1.96535f
C1118 VDD.t1378 VSS 1.96535f
C1119 VDD.t866 VSS 1.36987f
C1120 VDD.t798 VSS 1.45794f
C1121 VDD.t638 VSS 1.96535f
C1122 VDD.t1512 VSS 1.96535f
C1123 VDD.t3013 VSS 1.36987f
C1124 VDD.t664 VSS 1.31955f
C1125 VDD.t2542 VSS 1.96535f
C1126 VDD.t2573 VSS 1.96535f
C1127 VDD.t1373 VSS 1.45794f
C1128 VDD.t674 VSS 1.45794f
C1129 VDD.t1549 VSS 1.96535f
C1130 VDD.t496 VSS 1.96535f
C1131 VDD.t508 VSS 1.36987f
C1132 VDD.t1164 VSS 1.45794f
C1133 VDD.t1714 VSS 1.96535f
C1134 VDD.t287 VSS 1.96535f
C1135 VDD.t290 VSS 1.36987f
C1136 VDD.t289 VSS 1.31955f
C1137 VDD.t288 VSS 1.96535f
C1138 VDD.t1206 VSS 1.96535f
C1139 VDD.t1081 VSS 1.45794f
C1140 VDD.n2025 VSS 1.049f
C1141 VDD.n2123 VSS 1.83791f
C1142 VDD.t962 VSS 3.35165f
C1143 VDD.t390 VSS 4.24765f
C1144 VDD.t407 VSS 2.51852f
C1145 VDD.t402 VSS 2.42329f
C1146 VDD.n2188 VSS 1.94948f
C1147 VDD.t27 VSS 3.42569f
C1148 VDD.t925 VSS 3.43836f
C1149 VDD.t34 VSS 3.66626f
C1150 VDD.t20 VSS 2.8468f
C1151 VDD.t25 VSS 2.8468f
C1152 VDD.t32 VSS 3.52342f
C1153 VDD.t14 VSS 3.52342f
C1154 VDD.t23 VSS 1.52113f
C1155 VDD.t593 VSS 9.19382f
C1156 VDD.n2317 VSS 1.26071f
C1157 VDD.t883 VSS 9.19382f
C1158 VDD.t49 VSS 9.81076f
C1159 VDD.t66 VSS 7.617919f
C1160 VDD.t134 VSS 7.617919f
C1161 VDD.t62 VSS 9.428519f
C1162 VDD.t76 VSS 9.213929f
C1163 VDD.t55 VSS 9.81076f
C1164 VDD.t122 VSS 7.617919f
C1165 VDD.t51 VSS 7.617919f
C1166 VDD.t120 VSS 9.428519f
C1167 VDD.t58 VSS 9.428519f
C1168 VDD.t73 VSS 4.02355f
C1169 VDD.t78 VSS 9.213929f
C1170 VDD.t405 VSS 3.66626f
C1171 VDD.t568 VSS 3.43571f
C1172 VDD.n2354 VSS 1.55371f
C1173 VDD.n2355 VSS 1.55371f
C1174 VDD.t910 VSS 3.43571f
C1175 VDD.t12 VSS 3.66626f
C1176 VDD.t38 VSS 1.73916f
C1177 VDD.t16 VSS 3.52342f
C1178 VDD.t18 VSS 2.53105f
C1179 VDD.n2356 VSS 4.61542f
C1180 VDD.t583 VSS 8.89875f
C1181 VDD.t70 VSS 9.81076f
C1182 VDD.t115 VSS 7.617919f
C1183 VDD.t53 VSS 7.617919f
C1184 VDD.t47 VSS 9.428519f
C1185 VDD.t64 VSS 9.428519f
C1186 VDD.t96 VSS 4.02355f
C1187 VDD.n5268 VSS 12.0304f
C1188 VDD.t404 VSS 9.213929f
C1189 VDD.t613 VSS 9.19382f
C1190 VDD.t398 VSS 9.81076f
C1191 VDD.t411 VSS 7.617919f
C1192 VDD.t408 VSS 7.617919f
C1193 VDD.t400 VSS 9.428519f
C1194 VDD.t396 VSS 9.428519f
C1195 VDD.t409 VSS 4.02355f
C1196 VDD.t410 VSS 9.213929f
C1197 VDD.t413 VSS 4.02355f
C1198 VDD.t401 VSS 9.428519f
C1199 VDD.t397 VSS 9.428519f
C1200 VDD.t412 VSS 7.617919f
C1201 VDD.t399 VSS 7.617919f
C1202 VDD.t395 VSS 9.81076f
C1203 VDD.t839 VSS 9.19382f
C1204 VDD.n5376 VSS 4.15767f
C1205 VDD.t403 VSS 9.428519f
C1206 VDD.t392 VSS 7.617919f
C1207 VDD.t415 VSS 7.617919f
C1208 VDD.t391 VSS 9.81076f
C1209 VDD.t616 VSS 9.19382f
C1210 VDD.n5488 VSS 1.75925f
C1211 VDD.n5912 VSS 2.44316f
C1212 VDD.t406 VSS 9.428519f
C1213 VDD.t394 VSS 7.617919f
C1214 VDD.t416 VSS 7.617919f
C1215 VDD.t393 VSS 9.81076f
C1216 VDD.t586 VSS 9.19382f
C1217 VDD.n6013 VSS 1.84672f
C1218 VDD.n6266 VSS 1.1439f
C1219 VDD.n6311 VSS 4.50638f
C1220 VDD.n6326 VSS 2.86995f
C1221 VDD.n6327 VSS 1.64177f
C1222 VDD.n6370 VSS 4.15767f
C1223 VDD.n6396 VSS 3.80896f
C1224 VDD.n6577 VSS 3.80896f
C1225 VDD.t60 VSS 9.428519f
C1226 VDD.t68 VSS 7.617919f
C1227 VDD.t137 VSS 7.617919f
C1228 VDD.t82 VSS 9.81076f
C1229 VDD.t886 VSS 9.19382f
C1230 VDD.n6633 VSS 12.0304f
C1231 VDD.n6685 VSS 1.78684f
C1232 VDD.n6713 VSS 1.39946f
C1233 VDD.n7040 VSS 3.80896f
C1234 VDD.n7048 VSS 1.1439f
C1235 VDD.n7086 VSS 3.80896f
C1236 VDD.n7133 VSS 4.15767f
C1237 VDD.n7834 VSS 4.4125f
C1238 VDD.n7995 VSS 1.4234f
C1239 VDD.n8077 VSS 1.4234f
C1240 VDD.n8089 VSS 1.8928f
C1241 VDD.t2127 VSS 1.36987f
C1242 VDD.t603 VSS 1.45794f
C1243 VDD.t2254 VSS 1.96535f
C1244 VDD.t680 VSS 1.96535f
C1245 VDD.t2302 VSS 1.31955f
C1246 VDD.t2061 VSS 1.36987f
C1247 VDD.t1893 VSS 1.96535f
C1248 VDD.t2155 VSS 1.96535f
C1249 VDD.t1917 VSS 1.45794f
C1250 VDD.t2447 VSS 1.45794f
C1251 VDD.t2160 VSS 1.96535f
C1252 VDD.t560 VSS 1.96535f
C1253 VDD.t2189 VSS 1.31955f
C1254 VDD.t707 VSS 1.36987f
C1255 VDD.t367 VSS 1.36987f
C1256 VDD.t2325 VSS 1.96535f
C1257 VDD.t842 VSS 1.96535f
C1258 VDD.t1251 VSS 1.45794f
C1259 VDD.t979 VSS 1.45794f
C1260 VDD.t667 VSS 1.96535f
C1261 VDD.t417 VSS 1.96535f
C1262 VDD.t301 VSS 1.31955f
C1263 VDD.t544 VSS 1.36987f
C1264 VDD.t6 VSS 1.36987f
C1265 VDD.t546 VSS 1.96535f
C1266 VDD.t2464 VSS 1.96535f
C1267 VDD.t1265 VSS 1.45794f
C1268 VDD.t1333 VSS 1.45794f
C1269 VDD.t1489 VSS 1.96535f
C1270 VDD.t0 VSS 1.96535f
C1271 VDD.t2 VSS 1.31955f
C1272 VDD.t792 VSS 1.96535f
C1273 VDD.t2058 VSS 1.96535f
C1274 VDD.t2812 VSS 1.36987f
C1275 VDD.t2021 VSS 1.31955f
C1276 VDD.t2251 VSS 1.96535f
C1277 VDD.t1408 VSS 1.96535f
C1278 VDD.t810 VSS 1.45794f
C1279 VDD.t1 VSS 1.96535f
C1280 VDD.t898 VSS 1.96535f
C1281 VDD.t1195 VSS 1.45794f
C1282 VDD.t297 VSS 1.96535f
C1283 VDD.t630 VSS 1.96535f
C1284 VDD.t1818 VSS 1.45794f
C1285 VDD.t1015 VSS 1.45794f
C1286 VDD.t2099 VSS 1.96535f
C1287 VDD.t543 VSS 1.96535f
C1288 VDD.t545 VSS 1.31955f
C1289 VDD.t1796 VSS 1.96535f
C1290 VDD.t2079 VSS 1.96535f
C1291 VDD.t1824 VSS 1.45794f
C1292 VDD.t1042 VSS 1.45794f
C1293 VDD.t836 VSS 1.96535f
C1294 VDD.t2559 VSS 1.96535f
C1295 VDD.t2288 VSS 1.31955f
C1296 VDD.t1867 VSS 1.45794f
C1297 VDD.t2142 VSS 1.96535f
C1298 VDD.t551 VSS 1.96535f
C1299 VDD.t2088 VSS 1.36987f
C1300 VDD.t2228 VSS 1.31955f
C1301 VDD.t622 VSS 1.96535f
C1302 VDD.t2399 VSS 1.96535f
C1303 VDD.t720 VSS 1.45905f
C1304 VDD.n9182 VSS 1.049f
C1305 VDD.t598 VSS 1.45794f
C1306 VDD.t2349 VSS 1.96535f
C1307 VDD.t305 VSS 1.96535f
C1308 VDD.t303 VSS 1.36987f
C1309 VDD.t755 VSS 1.45905f
C1310 VDD.t1349 VSS 1.96535f
C1311 VDD.t302 VSS 1.96535f
C1312 VDD.t326 VSS 1.31955f
C1313 VDD.t930 VSS 1.45794f
C1314 VDD.t677 VSS 1.96535f
C1315 VDD.t3423 VSS 1.96535f
C1316 VDD.t3613 VSS 1.31955f
C1317 VDD.t1711 VSS 1.36987f
C1318 VDD.t1494 VSS 1.96535f
C1319 VDD.t1177 VSS 1.96535f
C1320 VDD.t1322 VSS 1.45794f
C1321 VDD.t1439 VSS 1.45794f
C1322 VDD.t648 VSS 1.96535f
C1323 VDD.t507 VSS 1.96535f
C1324 VDD.t510 VSS 1.31955f
C1325 VDD.t1180 VSS 1.45794f
C1326 VDD.t1370 VSS 1.96535f
C1327 VDD.t3678 VSS 1.96535f
C1328 VDD.t1405 VSS 1.31955f
C1329 VDD.t2921 VSS 1.36987f
C1330 VDD.t3747 VSS 1.96535f
C1331 VDD.t955 VSS 1.96535f
C1332 VDD.t813 VSS 1.45794f
C1333 VDD.t1209 VSS 1.45794f
C1334 VDD.t1262 VSS 1.96535f
C1335 VDD.t2261 VSS 1.96535f
C1336 VDD.t1338 VSS 1.31955f
C1337 VDD.t1957 VSS 1.45794f
C1338 VDD.t1799 VSS 1.96535f
C1339 VDD.t351 VSS 1.96535f
C1340 VDD.t353 VSS 1.31955f
C1341 VDD.t363 VSS 1.36987f
C1342 VDD.t352 VSS 1.96535f
C1343 VDD.t1365 VSS 1.96535f
C1344 VDD.t2570 VSS 1.45794f
C1345 VDD.t2680 VSS 1.45794f
C1346 VDD.t1049 VSS 1.96535f
C1347 VDD.t2774 VSS 1.96535f
C1348 VDD.t3354 VSS 1.31955f
C1349 VDD.t780 VSS 1.45794f
C1350 VDD.t697 VSS 1.96535f
C1351 VDD.t552 VSS 1.96535f
C1352 VDD.t554 VSS 1.31955f
C1353 VDD.t555 VSS 1.36987f
C1354 VDD.t553 VSS 1.96535f
C1355 VDD.t893 VSS 1.96535f
C1356 VDD.t935 VSS 1.45794f
C1357 VDD.t745 VSS 1.45794f
C1358 VDD.t944 VSS 1.96535f
C1359 VDD.t321 VSS 1.96535f
C1360 VDD.t293 VSS 1.31955f
C1361 VDD.t1112 VSS 1.45794f
C1362 VDD.t2231 VSS 1.96535f
C1363 VDD.t522 VSS 1.96535f
C1364 VDD.t519 VSS 1.31955f
C1365 VDD.t520 VSS 1.36987f
C1366 VDD.t521 VSS 1.96535f
C1367 VDD.t1747 VSS 1.96535f
C1368 VDD.t1354 VSS 1.45794f
C1369 VDD.t823 VSS 1.45794f
C1370 VDD.t610 VSS 1.96535f
C1371 VDD.t2344 VSS 1.96535f
C1372 VDD.t502 VSS 1.31955f
C1373 VDD.t2076 VSS 1.45794f
C1374 VDD.t1821 VSS 1.96535f
C1375 VDD.t2729 VSS 1.96535f
C1376 VDD.t1850 VSS 1.31955f
C1377 VDD.t1708 VSS 1.36987f
C1378 VDD.t1486 VSS 1.96535f
C1379 VDD.t725 VSS 1.96535f
C1380 VDD.t1505 VSS 1.45794f
C1381 VDD.t976 VSS 1.45794f
C1382 VDD.t748 VSS 1.96535f
C1383 VDD.t795 VSS 1.96535f
C1384 VDD.t2422 VSS 1.31955f
C1385 VDD.t686 VSS 1.45794f
C1386 VDD.t1611 VSS 1.96535f
C1387 VDD.t523 VSS 1.96535f
C1388 VDD.t529 VSS 1.31955f
C1389 VDD.t524 VSS 1.36987f
C1390 VDD.t532 VSS 1.96535f
C1391 VDD.t1515 VSS 1.96535f
C1392 VDD.t1299 VSS 1.45794f
C1393 VDD.t1780 VSS 1.45794f
C1394 VDD.t1086 VSS 1.96535f
C1395 VDD.t535 VSS 1.96535f
C1396 VDD.t537 VSS 1.31955f
C1397 VDD.n12633 VSS 1.76802f
C1398 VDD.n12634 VSS 2.45351f
C1399 a_52635_34067.n1 VSS 1.05429f
C1400 a_52635_34067.n4 VSS 1.05429f
C1401 a_52635_34067.n6 VSS 1.04685f
C1402 a_52635_34067.n10 VSS 1.04685f
C1403 a_52635_34067.n12 VSS 1.05549f
C1404 a_52635_34067.n19 VSS 1.35551f
C1405 a_52635_34067.n21 VSS 1.35551f
C1406 a_52635_34067.n25 VSS 1.05549f
C1407 a_52635_34067.n27 VSS 1.05056f
C1408 a_52635_34067.n30 VSS 1.05056f
C1409 a_52635_34067.n33 VSS 1.34521f
C1410 a_52635_34067.n36 VSS 1.34521f
C1411 a_52635_34067.n44 VSS 1.50271f
C1412 a_52635_34067.n55 VSS 2.60562f
C1413 a_52635_34067.n57 VSS 1.10968f
C1414 a_52635_34067.n58 VSS 1.8542f
C1415 a_52635_34067.n60 VSS 2.60562f
C1416 a_52635_34067.n61 VSS 1.05782f
C1417 a_52635_34067.n64 VSS 2.60562f
C1418 a_52635_34067.n67 VSS 1.05782f
C1419 a_52635_34067.n68 VSS 2.60562f
C1420 a_52635_34067.n70 VSS 1.3574f
C1421 a_52635_34067.n71 VSS 1.04844f
C1422 a_52635_34067.n74 VSS 2.64985f
C1423 a_52635_34067.n75 VSS 2.65467f
C1424 a_52635_34067.n79 VSS 2.65467f
C1425 a_52635_34067.n80 VSS 1.04847f
C1426 a_52635_34067.n82 VSS 2.64985f
C1427 a_52635_34067.n86 VSS 1.8542f
C1428 a_52635_34067.n88 VSS 1.8542f
C1429 a_52635_34067.n90 VSS 1.8542f
C1430 a_52635_34067.n92 VSS 2.51871f
C1431 a_52635_34067.n93 VSS 1.36384f
C1432 a_52635_34067.n94 VSS 1.36384f
C1433 a_52635_34067.n95 VSS 2.51871f
C1434 a_52635_34067.n96 VSS 1.93502f
C1435 a_52635_34067.n98 VSS 1.93502f
C1436 a_52635_34067.n100 VSS 1.93502f
C1437 a_52635_34067.n102 VSS 1.93502f
C1438 a_52635_34067.n104 VSS 2.54563f
C1439 a_52635_34067.n105 VSS 1.38682f
C1440 a_52635_34067.n106 VSS 1.38682f
C1441 a_52635_34067.n107 VSS 2.54563f
C1442 a_52635_34067.n109 VSS 2.51775f
C1443 a_52635_34067.n110 VSS 1.10968f
C1444 a_52635_34067.n111 VSS 2.51775f
C1445 a_52635_34067.n112 VSS 2.53332f
C1446 a_52635_34067.n113 VSS 1.11217f
C1447 a_52635_34067.n114 VSS 1.38815f
C1448 a_52635_34067.n115 VSS 1.11218f
C1449 a_52635_34067.n116 VSS 2.53332f
C1450 a_52635_34067.n138 VSS 1.16767f
C1451 a_52635_34067.t40 VSS 1.50638f
C1452 a_52635_34067.n140 VSS 2.01071f
C1453 a_52635_34067.n145 VSS 2.65583f
C1454 a_52635_34067.n146 VSS 2.3552f
C1455 a_52635_34067.t35 VSS 1.08042f
C1456 a_52635_34067.t12 VSS 3.04611f
C1457 a_52635_34067.n147 VSS 3.51664f
C1458 a_52635_34067.n148 VSS 3.42219f
C1459 a_52635_34067.n149 VSS 1.45207f
C1460 a_52635_34067.n156 VSS 5.15047f
C1461 a_52635_34067.n159 VSS 5.15047f
C1462 a_52635_34067.n164 VSS 3.42219f
C1463 a_52635_34067.n165 VSS 3.42219f
C1464 a_52635_34067.n166 VSS 5.34875f
C1465 a_52635_34067.n167 VSS 5.34875f
C1466 a_52635_34067.n168 VSS 3.42219f
C1467 a_52635_34067.n169 VSS 3.48946f
C1468 a_52635_34067.n170 VSS 3.8813f
C1469 a_52635_34067.n171 VSS 2.83365f
C1470 a_52635_34067.n172 VSS 3.65877f
C1471 a_52635_34067.n178 VSS 3.65877f
C1472 a_52635_34067.n179 VSS 2.14406f
C1473 a_52635_34067.n180 VSS 2.39757f
C1474 a_52635_34067.n181 VSS 2.73209f
C1475 a_52635_34067.n186 VSS 1.28863f
C1476 a_52635_34067.t57 VSS 2.58185f
C1477 a_52635_34067.n187 VSS 3.88688f
C1478 a_52635_34067.t59 VSS 1.9214f
C1479 a_52635_34067.n189 VSS 2.80961f
C1480 a_52635_34067.n190 VSS 4.57473f
C1481 a_52635_34067.n191 VSS 3.72315f
C1482 a_52635_34067.n194 VSS 3.69214f
C1483 a_52635_34067.t39 VSS 1.08042f
C1484 a_52635_34067.t22 VSS 3.04611f
C1485 a_52635_34067.t16 VSS 1.21614f
C1486 a_52635_34067.n195 VSS 1.5238f
C1487 a_52635_34067.n196 VSS 2.37199f
C1488 a_52635_34067.n197 VSS 2.11719f
C1489 a_52635_34067.n207 VSS 2.11719f
C1490 a_52635_34067.n210 VSS 2.3552f
C1491 a_52635_34067.n211 VSS 2.73209f
C1492 a_52635_34067.t8 VSS 1.21614f
C1493 a_52635_34067.n212 VSS 1.5238f
C1494 a_52635_34067.n213 VSS 2.37199f
C1495 a_52635_34067.n214 VSS 2.13513f
.ends

