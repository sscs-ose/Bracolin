* NGSPICE file created from CM_input.ext - technology: gf180mcuD

.subckt CM_input ISBCS INP INP2 INN INN2 VDD VSS
X0 a_3930_2285# ISBCS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X1 a_948_n291# ISBCS ISBCS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X2 INN a_n389_6663# a_3947_7622# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3 a_3930_609# ISBCS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X4 INN2 a_n389_6663# a_3947_5704# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X5 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X6 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X7 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X8 a_n389_6663# ISBCS a_3930_609# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X9 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X10 VSS ISBCS a_948_1385# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X11 a_n389_6663# a_n389_6663# a_3947_6663# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X12 a_3930_n291# ISBCS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X13 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X14 VSS ISBCS a_948_609# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X15 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X16 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X17 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X18 a_3947_7622# a_n389_6663# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X19 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X20 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X21 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X22 a_3947_5704# a_n389_6663# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X23 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X24 VSS ISBCS a_948_2285# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X25 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X26 a_948_609# ISBCS INP2 VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X27 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X28 a_941_7622# a_n389_6663# INN2 VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X29 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X30 a_n389_6663# ISBCS a_3930_1385# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X31 a_3947_6663# a_n389_6663# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X32 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X33 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X34 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X35 a_941_5704# a_n389_6663# INN VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X36 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X37 a_948_1385# ISBCS INP2 VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X38 VDD a_n389_6663# a_941_7622# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X39 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X40 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X41 VSS ISBCS a_948_n291# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X42 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X43 a_941_6663# a_n389_6663# a_n389_6663# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X44 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X45 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X46 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X47 VDD a_n389_6663# a_941_5704# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X48 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X49 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X50 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X51 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X52 VDD a_n389_6663# a_941_6663# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X53 ISBCS ISBCS a_3930_2285# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X54 a_3930_1385# ISBCS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X55 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X56 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X57 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X58 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X59 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X60 a_948_2285# ISBCS INP VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X61 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X62 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X63 INP ISBCS a_3930_n291# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X64 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X65 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
.ends

