* Extracted by KLayout with GF180MCU LVS runset on : 18/02/2024 19:49

.SUBCKT neg_bottom_plate VSSD CK11 VDDD
M$1 \$2 CK11 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$2 \$8 \$2 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$3 \$6 \$5 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$4 \$4 \$8 \$3 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$5 \$5 \$2 \$3 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$6 \$4 \$2 \$6 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$7 \$4 \$2 \$3 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$8 \$5 \$8 \$3 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$9 \$4 \$8 \$6 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$10 \$2 CK11 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$11 \$8 \$2 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$12 \$6 \$5 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
.ENDS neg_bottom_plate
