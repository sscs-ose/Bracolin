* NGSPICE file created from Filter_TOP.ext - technology: gf180mcuD

.subckt Filter_TOP VCM IN_POS IN_NEG VSS I1U VDD I1N IBNOUT OUT IBPOUT
X0 VSS.t3638 VSS.t3637 VSS.t3638 VSS.t1109 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1 a_52635_49681.t175 a_52635_34067.t65 VDD.t4983 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2 VDD.t4745 VDD.t4744 VDD.t4745 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3 VDD.t4743 VDD.t4742 VDD.t4743 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4 VDD.t4741 VDD.t4740 VDD.t4741 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5 VDD.t4739 VDD.t4738 VDD.t4739 VDD.t318 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6 a_100820_11614.t5 a_57977_n12421.t0 a_102796_6405# VSS.t173 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X7 a_31284_4481.t2 a_30324_4421.t0 a_30724_6405# VSS.t146 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X8 VDD.t4737 VDD.t4736 VDD.t4737 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X9 a_102756_12380# a_100820_10448.t12 VDD.t369 VDD.t325 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X10 a_36032_n36322.t2 a_53829_n36382.t8 a_55635_n36322# VDD.t334 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X11 a_33249_35053.t141 a_35502_25545.t28 VSS.t164 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X12 VSS.t3636 VSS.t3635 VSS.t3636 VSS.t576 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X13 VSS.t3634 VSS.t3633 VSS.t3634 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X14 a_101350_10448# a_100820_10448.t4 a_100820_10448.t5 VDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X15 a_52635_49681.t174 a_52635_34067.t66 VDD.t4982 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X16 a_38619_n2651# a_31953_n19727.t74 a_38097_n2651# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X17 VDD.t4735 VDD.t4734 VDD.t4735 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X18 VSS.t3632 VSS.t3631 VSS.t3632 VSS.t910 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X19 VSS.t3630 VSS.t3629 VSS.t3630 VSS.t171 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X20 VDD.t48 a_31699_20742.t45 a_35502_24538.t23 VDD.t17 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X21 VSS.t3628 VSS.t3627 VSS.t3628 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X22 a_43817_6405# a_41891_4481.t11 VSS.t179 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X23 VSS.t3626 VSS.t3625 VSS.t3626 VSS.t458 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X24 VSS.t3624 VSS.t3623 VSS.t3624 VSS.t984 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X25 VDD.t4733 VDD.t4732 VDD.t4733 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X26 a_105365_n7865# a_71281_n8397.t74 a_104527_n7865# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X27 VDD.t49 a_31699_20742.t46 a_35502_25545.t0 VDD.t41 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X28 a_52635_34067.t5 a_35922_19591.t6 a_52635_48695.t87 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X29 a_58851_n7138# a_50751_n19729.t74 a_58329_n8035# VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X30 a_53145_n19597# a_50751_n19729.t75 a_52585_n19597# VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X31 a_71864_n30339# a_65486_n36322.t8 a_71342_n30339.t3 VSS.t153 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X32 VDD.t4731 VDD.t4730 VDD.t4731 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X33 VSS.t3622 VSS.t3621 VSS.t3622 VSS.t563 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X34 a_106809_n17715.t0 a_71281_n8397.t75 a_106501_n21335# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X35 VSS.t3620 VSS.t3619 VSS.t3620 VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X36 VSS.t3618 VSS.t3617 VSS.t3618 VSS.t426 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X37 VDD.t4729 VDD.t4728 VDD.t4729 VDD.t21 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X38 VDD.t4727 VDD.t4726 VDD.t4727 VDD.t73 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X39 a_105933_n2435# a_71281_n8397.t76 a_105365_n2435# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X40 VSS.t3616 VSS.t3615 VSS.t3616 VSS.t316 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X41 VDD.t4725 VDD.t4724 VDD.t4725 VDD.t3679 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X42 a_52635_34067.t6 a_35922_19591.t7 a_52635_48695.t86 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X43 VDD.t4723 VDD.t4722 VDD.t4723 VDD.t979 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X44 a_33249_48695.t332 a_31699_20742.t47 VDD.t51 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X45 VSS.t3614 VSS.t3613 VSS.t3614 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X46 a_52635_48695.t175 a_52635_34067.t67 VDD.t4981 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X47 VSS.t3612 VSS.t3611 VSS.t3612 VSS.t297 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X48 OUT.t107 a_35922_19591.t8 a_52635_49681.t0 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X49 VDD.t4721 VDD.t4720 VDD.t4721 VDD.t394 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X50 VDD.t4719 VDD.t4718 VDD.t4719 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X51 VSS.t3610 VSS.t3609 VSS.t3610 VSS.t952 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X52 VSS.t3608 VSS.t3607 VSS.t3608 VSS.t913 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X53 VSS.t3606 VSS.t3605 VSS.t3606 VSS.t162 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X54 a_33249_48695.t331 a_31699_20742.t48 VDD.t53 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X55 VDD.t55 a_31699_20742.t49 a_33249_48695.t330 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X56 VDD.t4717 VDD.t4716 VDD.t4717 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X57 VSS.t3604 VSS.t3603 VSS.t3604 VSS.t1827 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X58 a_31284_n30339.t1 a_30324_n30399.t1 a_30724_n30339# VSS.t146 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X59 VSS.t3602 VSS.t3601 VSS.t3602 VSS.t284 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X60 VDD.t4715 VDD.t4714 VDD.t4715 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X61 OUT.t106 a_35922_19591.t9 a_52635_49681.t1 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X62 a_33249_35053.t0 a_35502_24538.t24 OUT.t19 VSS.t159 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X63 VDD.t4713 VDD.t4712 VDD.t4713 VDD.t947 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X64 a_38097_n5342.t0 a_100992_n29313.t0 a_101392_n29181# VSS.t384 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X65 VDD.t466 a_71281_n8397.t72 a_71281_n8397.t73 VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X66 a_101392_6405# a_100992_4421.t0 a_100820_10448.t0 VSS.t175 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X67 VDD.t4711 VDD.t4710 VDD.t4711 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X68 a_52635_48695.t85 a_35922_19591.t10 a_52635_34067.t7 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X69 VDD.t57 a_31699_20742.t50 a_33249_48695.t329 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X70 VSS.t3600 VSS.t3599 VSS.t3600 VSS.t643 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X71 VDD.t4709 VDD.t4708 VDD.t4709 VDD.t2467 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X72 a_100235_n15000# a_71281_n8397.t77 a_99667_n15000# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X73 VDD.t4707 VDD.t4706 VDD.t4707 VDD.t1422 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X74 VSS.t3598 VSS.t3597 VSS.t3598 VSS.t901 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X75 a_73302_13546# a_71496_10388.t8 a_71342_4481.t3 VDD.t491 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X76 a_30724_6405# a_30324_4421.t0 a_30152_10448.t3 VSS.t145 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X77 VDD.t4705 VDD.t4704 VDD.t4705 VDD.t979 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X78 VSS.t3596 VSS.t3595 VSS.t3596 VSS.t191 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X79 VDD.t4703 VDD.t4702 VDD.t4703 VDD.t1749 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X80 VDD.t4701 VDD.t4700 VDD.t4701 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X81 VSS.t3594 VSS.t3593 VSS.t3594 VSS.t655 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X82 a_31831_n5342.t0 a_32913_n8930.t1 a_83725_n28415# VSS.t366 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X83 a_45445_n18698# a_31953_n19727.t75 a_44885_n17801# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X84 VSS.t3592 VSS.t3591 VSS.t3592 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X85 VDD.t59 a_31699_20742.t51 a_33249_48695.t328 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X86 OUT.t105 a_35922_19591.t11 a_52635_49681.t2 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X87 VDD.t4699 VDD.t4698 VDD.t4699 VDD.t947 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X88 VSS.t3590 VSS.t3589 VSS.t3590 VSS.t527 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X89 VDD.t4697 VDD.t4696 VDD.t4697 VDD.t311 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X90 VDD.t4695 VDD.t4694 VDD.t4695 VDD.t2450 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X91 VSS.t3588 VSS.t3587 VSS.t3588 VSS.t251 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X92 a_51711_n5344.t1 a_50751_n19729.t76 a_51151_n5344# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X93 a_66551_n17803# a_50751_n19729.t77 a_66029_n18700# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X94 a_33249_35053.t1 a_33379_34917.t3 a_33249_48695.t18 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X95 VSS.t3586 VSS.t3585 VSS.t3586 VSS.t692 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X96 a_33249_35053.t2 a_33379_34917.t4 a_33249_48695.t19 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X97 a_98829_n17715# a_71281_n8397.t78 a_98299_n16810# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X98 OUT.t104 a_35922_19591.t12 a_52635_49681.t3 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X99 VSS.t3584 VSS.t3583 VSS.t3584 VSS.t1543 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X100 a_73302_11614# a_71496_10388.t9 VSS.t347 VDD.t491 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X101 a_73268_n29181# a_65486_n36322.t9 a_45445_n19595.t1 VSS.t156 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X102 a_90245_n6055# a_71281_n10073.t74 a_60677_10448.t4 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X103 VDD.t4693 VDD.t4692 VDD.t4693 VDD.t545 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X104 VSS.t3582 VSS.t3581 VSS.t3582 VSS.t889 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X105 a_98829_n15000# a_71281_n8397.t79 a_98299_n15905# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X106 a_51711_n14215# a_50751_n19729.t78 a_51151_n14215# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X107 VDD.t4691 VDD.t4690 VDD.t4691 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X108 VDD.t4689 VDD.t4688 VDD.t4689 VDD.t79 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X109 VSS.t3580 VSS.t3579 VSS.t3580 VSS.t94 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X110 VSS.t3578 VSS.t3577 VSS.t3578 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X111 a_33249_48695.t339 a_33379_34007.t4 a_33249_34067.t105 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X112 VDD.t4687 VDD.t4686 VDD.t4687 VDD.t572 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X113 VDD.t4685 VDD.t4684 VDD.t4685 VDD.t933 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X114 a_65486_n35156.t3 a_65486_n35156.t2 a_67422_n36322# VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X115 a_60285_n2653# a_50751_n19729.t79 a_59763_n3550# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X116 a_71281_n8397.t71 a_71281_n8397.t70 VDD.t465 VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X117 VDD.t4683 VDD.t4682 VDD.t4683 VDD.t1497 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X118 a_105365_n15000# a_71281_n8397.t80 a_104527_n15000# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X119 VDD.t4681 VDD.t4680 VDD.t4681 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X120 a_106676_n30339.t1 a_100820_n36322.t8 a_108602_n27257# VSS.t350 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X121 VDD.t4679 VDD.t4678 VDD.t4679 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X122 VSS.t3576 VSS.t3575 VSS.t3576 VSS.t686 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X123 a_40613_n8930# a_31953_n19727.t76 a_40053_n8930# VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X124 a_33249_48695.t340 a_33379_34007.t5 a_33249_34067.t104 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X125 VDD.t4677 VDD.t4676 VDD.t4677 VDD.t488 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X126 VDD.t4675 VDD.t4674 VDD.t4675 VDD.t332 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X127 OUT.t103 a_35922_19591.t13 a_52635_49681.t4 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X128 VSS.t3574 VSS.t3573 VSS.t3574 VSS.t839 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X129 VSS.t3572 VSS.t3571 VSS.t3572 VSS.t822 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X130 a_110225_n1530# a_71281_n8397.t81 a_109695_n5150# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X131 a_52635_48695.t84 a_35922_19591.t14 a_52635_34067.t8 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X132 a_88271_n3340# a_71281_n10073.t75 a_87433_n3340# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X133 VDD.t4768 a_83153_11614.t8 a_90935_5639# VSS.t398 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X134 VDD.t4673 VDD.t4672 VDD.t4673 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X135 VDD.t4671 VDD.t4670 VDD.t4671 VDD.t318 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X136 VSS.t3570 VSS.t3569 VSS.t3570 VSS.t214 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X137 a_114516_10448# a_86903_n14095.t3 a_89715_n17715.t2 VDD.t373 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X138 VDD.t4669 VDD.t4668 VDD.t4669 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X139 a_39179_n8033# a_31953_n19727.t77 a_38619_n8033# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X140 VDD.t60 a_31699_20742.t52 a_35502_25545.t1 VDD.t30 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X141 VSS.t3568 VSS.t3567 VSS.t3568 VSS.t658 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X142 VDD.t4667 VDD.t4666 VDD.t4667 VDD.t1716 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X143 VSS.t248 a_50751_n19729.t70 a_50751_n19729.t71 VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X144 VDD.t4665 VDD.t4664 VDD.t4665 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X145 a_84547_n15000# a_71281_n10073.t76 a_83709_n14095# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X146 VDD.t4663 VDD.t4662 VDD.t4663 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X147 a_100235_n20430# a_71281_n8397.t82 a_99667_n20430# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X148 VDD.t4661 VDD.t4660 VDD.t4661 VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X149 a_52635_49681.t5 a_35922_19591.t15 OUT.t102 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X150 VDD.t2 a_65486_n35156.t12 a_66016_n36322# VDD.t1 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X151 a_67111_n2653# a_50751_n19729.t80 a_66551_n1756# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X152 VDD.t4659 VDD.t4658 VDD.t4659 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X153 VDD.t4657 VDD.t4656 VDD.t4657 VDD.t1869 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X154 VDD.t4655 VDD.t4654 VDD.t4655 VDD.t313 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X155 VDD.t4653 VDD.t4652 VDD.t4653 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X156 a_54579_n4447# a_50751_n19729.t81 a_54019_n4447# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X157 a_32353_n7136# a_31953_n19727.t78 a_31831_n7136# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X158 VSS.t3566 VSS.t3565 VSS.t3566 VSS.t105 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X159 VSS.t288 a_112559_4481.t11 a_113081_5639# VSS.t287 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X160 a_30324_n30399.t1 a_30152_n36322.t8 a_36530_n29181# VSS.t325 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X161 VDD.t4651 VDD.t4650 VDD.t4651 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X162 VDD.t4649 VDD.t4648 VDD.t4649 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X163 VSS.t3564 VSS.t3563 VSS.t3564 VSS.t873 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X164 a_34347_n7136# a_31953_n19727.t79 a_33787_n7136# VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X165 VDD.t4647 VDD.t4646 VDD.t4647 VDD.t2402 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X166 a_48349_n35156# a_47819_n35156.t2 a_47819_n35156.t3 VDD.t2561 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X167 VSS.t3562 VSS.t3561 VSS.t3562 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X168 a_51711_n12421.t0 a_83153_11614.t9 a_89531_6405# VSS.t399 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X169 a_101350_n34390# a_100820_n35156.t11 a_100820_n36322.t0 VDD.t529 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X170 VSS.t3560 VSS.t3559 VSS.t3560 VSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X171 VSS.t3558 VSS.t3557 VSS.t3558 VSS.t1366 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X172 a_77225_4481.t1 a_77225_4481.t0 a_79151_5639# VSS.t335 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X173 a_106676_4481.t2 a_106830_10388.t8 a_107230_10448# VDD.t524 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X174 VDD.t4645 VDD.t4644 VDD.t4645 VDD.t901 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X175 VSS.t3556 VSS.t3555 VSS.t3556 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X176 a_33249_48695.t335 a_33379_34007.t6 a_33249_34067.t103 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X177 VSS.t3554 VSS.t3553 VSS.t3554 VSS.t63 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X178 VSS.t3552 VSS.t3551 VSS.t3552 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X179 a_57417_n8932# a_50751_n19729.t82 a_56895_n8932# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X180 VDD.t4643 VDD.t4642 VDD.t4643 VDD.t2779 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X181 a_98829_n20430# a_71281_n8397.t83 a_36032_n35156.t0 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X182 VDD.t4641 VDD.t4640 VDD.t4641 VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X183 VDD.t4639 VDD.t4638 VDD.t4639 VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X184 VSS.t3550 VSS.t3549 VSS.t3550 VSS.t126 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X185 VDD.t4637 VDD.t4636 VDD.t4637 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X186 VDD.t4635 VDD.t4634 VDD.t4635 VDD.t496 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X187 a_30152_n35156.t1 a_30152_n35156.t0 a_32088_n34390# VDD.t554 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X188 VSS.t3548 VSS.t3547 VSS.t3548 VSS.t542 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X189 VDD.t4633 VDD.t4632 VDD.t4633 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X190 a_89563_13546# a_89163_10388.t8 a_89033_13546.t0 VDD.t556 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X191 a_67422_13546# a_65486_10448.t11 VDD.t4748 VDD.t869 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X192 VDD.t4631 VDD.t4630 VDD.t4631 VDD.t2385 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X193 a_51151_n17803# a_50751_n19729.t83 a_50629_n17803# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X194 VSS.t3546 VSS.t3545 VSS.t3546 VSS.t858 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X195 VDD.t4629 VDD.t4628 VDD.t4629 VDD.t1660 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X196 a_43010_10448.t2 a_36032_11614.t3 a_42442_13546# VDD.t292 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X197 VSS.t3544 VSS.t3543 VSS.t3544 VSS.t847 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X198 a_52635_34067.t9 a_35922_19591.t16 a_52635_48695.t83 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X199 a_48349_n33224# a_47819_n35156.t6 a_47819_n35156.t7 VDD.t2561 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X200 a_42047_n19595# a_31953_n19727.t80 a_41487_n19595# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X201 a_30682_10448# a_30152_10448.t4 a_30152_10448.t5 VDD.t351 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X202 VDD.t4627 VDD.t4626 VDD.t4627 VDD.t575 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X203 VDD.t4625 VDD.t4624 VDD.t4625 VDD.t958 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X204 a_32088_n36322# a_30152_n35156.t12 VDD.t4746 VDD.t2091 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X205 VDD.t4623 VDD.t4622 VDD.t4623 VDD.t858 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X206 a_105365_n20430# a_71281_n8397.t84 a_104527_n20430# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X207 VDD.t4621 VDD.t4620 VDD.t4621 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X208 VSS.t3542 VSS.t3541 VSS.t3542 VSS.t15 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X209 VDD.t4980 a_52635_34067.t68 a_52635_48695.t174 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X210 OUT.t101 a_35922_19591.t17 a_52635_49681.t6 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X211 VDD.t4619 VDD.t4618 VDD.t4619 VDD.t901 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X212 VDD.t4617 VDD.t4616 VDD.t4617 VDD.t351 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X213 a_52635_34067.t10 a_35922_19591.t18 a_52635_48695.t82 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X214 VDD.t4615 VDD.t4614 VDD.t4615 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X215 VDD.t47 a_31699_20742.t43 a_31699_20742.t44 VDD.t41 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X216 a_33249_48695.t327 a_31699_20742.t53 VDD.t62 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X217 VSS.t3540 VSS.t3539 VSS.t3540 VSS.t385 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X218 VSS.t3538 VSS.t3537 VSS.t3538 VSS.t842 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X219 OUT.t100 a_35922_19591.t19 a_52635_49681.t7 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X220 a_52635_34067.t11 a_35922_19591.t20 a_52635_48695.t81 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X221 VDD.t4613 VDD.t4612 VDD.t4613 VDD.t1820 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X222 a_89563_11614# a_89163_10388.t9 a_81205_n14095.t1 VDD.t556 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X223 a_67422_11614# a_65486_10448.t12 VDD.t4749 VDD.t869 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X224 VDD.t4611 VDD.t4610 VDD.t4611 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X225 a_44885_n6239# a_31953_n19727.t81 a_44363_n7136# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X226 a_52635_49681.t8 a_35922_19591.t21 OUT.t99 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X227 VDD.t4609 VDD.t4608 VDD.t4609 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X228 a_31953_n19727.t71 a_31953_n19727.t70 VSS.t93 VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X229 a_43010_10448.t3 a_36032_11614.t4 a_42442_11614# VDD.t292 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X230 VSS.t3536 VSS.t3535 VSS.t3536 VSS.t563 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X231 VDD.t4607 VDD.t4606 VDD.t4607 VDD.t748 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X232 VSS.t354 a_89163_n36382.t8 a_89563_n35156# VDD.t548 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X233 VSS.t3534 VSS.t3533 VSS.t3534 VSS.t1432 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X234 VDD.t4605 VDD.t4604 VDD.t4605 VDD.t2347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X235 VDD.t4603 VDD.t4602 VDD.t4603 VDD.t858 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X236 a_31953_n19727.t69 a_31953_n19727.t68 VSS.t92 VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X237 a_47753_n15110# a_31953_n19727.t82 a_47231_n16904# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X238 VDD.t4601 VDD.t4600 VDD.t4601 VDD.t816 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X239 VDD.t4599 VDD.t4598 VDD.t4599 VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X240 VDD.t4597 VDD.t4596 VDD.t4597 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X241 VSS.t3532 VSS.t3531 VSS.t3532 VSS.t282 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X242 a_89531_6405# a_83153_11614.t10 VDD.t4769 VSS.t400 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X243 a_107339_n6055# a_71281_n8397.t85 a_106809_n5150.t0 VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X244 VSS.t3530 VSS.t3529 VSS.t3530 VSS.t768 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X245 VDD.t4595 VDD.t4594 VDD.t4595 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X246 VDD.t4593 VDD.t4592 VDD.t4593 VDD.t433 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X247 a_52635_34067.t2 a_35502_24538.t25 a_33249_34067.t17 VSS.t159 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X248 VSS.t372 a_41891_n29181.t11 a_42413_n27257# VSS.t171 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X249 VDD.t4591 VDD.t4590 VDD.t4591 VDD.t670 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X250 VDD.t4589 VDD.t4588 VDD.t4589 VDD.t923 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X251 VDD.t4587 VDD.t4586 VDD.t4587 VDD.t1789 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X252 VDD.t4585 VDD.t4584 VDD.t4585 VDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X253 VDD.t4583 VDD.t4582 VDD.t4583 VDD.t422 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X254 VSS.t3528 VSS.t3527 VSS.t3528 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X255 a_33249_48695.t336 a_33379_34007.t7 a_33249_34067.t102 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X256 a_89407_n6960# a_71281_n10073.t77 a_88839_n6960# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X257 VSS.t3526 VSS.t3525 VSS.t3526 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X258 VSS.t3524 VSS.t3523 VSS.t3524 VSS.t536 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X259 VDD.t4581 VDD.t4580 VDD.t4581 VDD.t845 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X260 a_89009_n27257.t0 a_89163_n36382.t9 a_89563_n33224# VDD.t548 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X261 a_89033_13546.t1 a_89163_10388.t10 a_90969_10448# VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X262 a_31699_20742.t42 a_31699_20742.t41 VDD.t46 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X263 VDD.t4579 VDD.t4578 VDD.t4579 VDD.t50 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X264 a_53699_n36322.t1 a_71496_n36382.t8 a_73302_n36322# VDD.t2061 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X265 VDD.t4577 VDD.t4576 VDD.t4577 VDD.t816 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X266 VSS.t3522 VSS.t3521 VSS.t3522 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X267 VDD.t4575 VDD.t4574 VDD.t4575 VDD.t831 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X268 a_100235_n15905# a_71281_n8397.t86 a_99667_n15905# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X269 VSS.t3520 VSS.t3519 VSS.t3520 VSS.t1800 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X270 VDD.t4573 VDD.t4572 VDD.t4573 VDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X271 VDD.t4571 VDD.t4570 VDD.t4571 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X272 a_33249_48695.t20 a_33379_34917.t5 a_33249_35053.t3 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X273 VDD.t64 a_31699_20742.t54 a_33249_48695.t326 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X274 a_40613_n14213# a_31953_n19727.t83 a_40053_n14213# VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X275 VSS.t3518 VSS.t3517 VSS.t3518 VSS.t283 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X276 a_67462_n29181# a_45445_n19595.t2 a_44363_n16007.t1 VSS.t412 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X277 a_31699_20742.t40 a_31699_20742.t39 VDD.t45 VDD.t26 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X278 VDD.t4569 VDD.t4568 VDD.t4569 VDD.t2305 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X279 VDD.t4567 VDD.t4566 VDD.t4567 VDD.t438 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X280 a_94537_n9675# a_71281_n10073.t78 a_93969_n9675# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X281 VDD.t4565 VDD.t4564 VDD.t4565 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X282 a_78344_n36322.t3 a_71366_n35156.t5 a_77776_n36322# VDD.t2046 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X283 a_33249_34067.t101 a_33379_34007.t8 a_33249_48695.t337 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X284 a_52635_34067.t12 a_35922_19591.t22 a_52635_48695.t80 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X285 VDD.t4563 VDD.t4562 VDD.t4563 VDD.t488 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X286 VSS.t3516 VSS.t3515 VSS.t3516 VSS.t381 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X287 VDD.t4561 VDD.t4560 VDD.t4561 VDD.t1644 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X288 VSS.t3514 VSS.t3513 VSS.t3514 VSS.t1472 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X289 VSS.t3512 VSS.t3511 VSS.t3512 VSS.t816 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X290 VDD.t4559 VDD.t4558 VDD.t4559 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X291 VDD.t4557 VDD.t4556 VDD.t4557 VDD.t845 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X292 a_39179_n19595.t1 a_31953_n19727.t84 a_38619_n19595# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X293 VSS.t3510 VSS.t3509 VSS.t3510 VSS.t313 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X294 VDD.t4555 VDD.t4554 VDD.t4555 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X295 VSS.t3508 VSS.t3507 VSS.t3508 VSS.t643 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X296 VSS.t3506 VSS.t3505 VSS.t3506 VSS.t813 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X297 a_60845_n19597# a_50751_n19729.t84 a_60285_n18700# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X298 VDD.t4553 VDD.t4552 VDD.t4553 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X299 VDD.t4551 VDD.t4550 VDD.t4551 VDD.t639 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X300 VDD.t4549 VDD.t4548 VDD.t4549 VDD.t831 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X301 VDD.t4547 VDD.t4546 VDD.t4547 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X302 VSS.t3504 VSS.t3503 VSS.t3504 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X303 a_71342_n30339.t0 a_71496_n36382.t9 a_71896_n36322# VDD.t2023 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X304 VDD.t4545 VDD.t4544 VDD.t4545 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X305 VSS.t3502 VSS.t3501 VSS.t3502 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X306 VDD.t4543 VDD.t4542 VDD.t4543 VDD.t402 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X307 VSS.t3500 VSS.t3499 VSS.t3500 VSS.t1391 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X308 VSS.t3498 VSS.t3497 VSS.t3498 VSS.t290 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X309 a_60285_n19597# a_50751_n19729.t85 a_57977_n19597# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X310 a_98829_n15905# a_71281_n8397.t87 a_98299_n15905# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X311 VSS.t3496 VSS.t3495 VSS.t3496 VSS.t260 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X312 VSS.t3494 VSS.t3493 VSS.t3494 VSS.t864 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X313 VSS.t3492 VSS.t3491 VSS.t3492 VSS.t1109 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X314 a_61484_4481# a_59558_4481.t11 VSS.t402 VSS.t314 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X315 VDD.t4541 VDD.t4540 VDD.t4541 VDD.t2257 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X316 a_54229_n35156# a_53829_n36382.t9 a_53699_n35156.t1 VDD.t322 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X317 a_82573_n13190# a_71281_n10073.t79 a_81735_n13190# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X318 VDD.t4539 VDD.t4538 VDD.t4539 VDD.t2682 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X319 VDD.t4537 VDD.t4536 VDD.t4537 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X320 VDD.t4535 VDD.t4534 VDD.t4535 VDD.t614 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X321 VSS.t3490 VSS.t3489 VSS.t3490 VSS.t692 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X322 VSS.t3488 VSS.t3487 VSS.t3488 VSS.t797 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X323 a_105365_n15905# a_71281_n8397.t88 a_104527_n15905# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X324 VSS.t3486 VSS.t3485 VSS.t3486 VSS.t822 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X325 VSS.t3484 VSS.t3483 VSS.t3484 VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X326 VSS.t194 a_35502_25545.t29 a_33249_35053.t140 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X327 VDD.t4533 VDD.t4532 VDD.t4533 VDD.t795 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X328 VSS.t3482 VSS.t3481 VSS.t3482 VSS.t558 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X329 a_39179_n3548# a_31953_n19727.t85 a_38619_n3548# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X330 a_94892_n29181.t10 a_83325_n29313.t1 a_96849_n36322# VDD.t1998 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X331 VDD.t4531 VDD.t4530 VDD.t4531 VDD.t792 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X332 VDD.t4529 VDD.t4528 VDD.t4529 VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X333 a_54579_n19597# a_50751_n19729.t86 a_54019_n18700# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X334 a_32353_n15110# a_31953_n19727.t86 a_31831_n15110# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X335 VSS.t3480 VSS.t3479 VSS.t3480 VSS.t214 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X336 VDD.t4527 VDD.t4526 VDD.t4527 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X337 a_64243_n18700# a_50751_n19729.t87 a_63683_n18700# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X338 a_54019_n4447# a_50751_n19729.t88 a_53497_n6241# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X339 VSS.t247 a_50751_n19729.t68 a_50751_n19729.t69 VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X340 VSS.t3478 VSS.t3477 VSS.t3478 VSS.t418 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X341 a_54229_n33224# a_53829_n36382.t10 a_36032_n36322.t3 VDD.t322 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X342 VSS.t3476 VSS.t3475 VSS.t3476 VSS.t259 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X343 a_88271_n2435# a_71281_n10073.t80 a_87433_n2435# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X344 a_31699_19142# I1U.t2 a_30377_18342# VSS.t362 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X345 VSS.t3474 VSS.t3473 VSS.t3474 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X346 a_79151_n29181# a_77225_n29181.t11 VSS.t388 VSS.t387 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X347 a_52635_34067.t13 a_35922_19591.t23 a_52635_48695.t79 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X348 VDD.t4525 VDD.t4524 VDD.t4525 VDD.t795 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X349 VSS.t3472 VSS.t3471 VSS.t3472 VSS.t780 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X350 a_52635_34067.t14 a_35922_19591.t24 a_52635_48695.t78 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X351 VSS.t3470 VSS.t3469 VSS.t3470 VSS.t414 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X352 VDD.t4523 VDD.t4522 VDD.t4523 VDD.t923 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X353 VDD.t4521 VDD.t4520 VDD.t4521 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X354 VDD.t4519 VDD.t4518 VDD.t4519 VDD.t758 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X355 a_81735_n8770# a_71281_n10073.t81 VDD.t307 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X356 VSS.t3468 VSS.t3467 VSS.t3468 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X357 VSS.t3466 VSS.t3465 VSS.t3466 VSS.t341 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X358 a_48313_n13316# a_31953_n19727.t87 a_47753_n13316# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X359 OUT.t98 a_35922_19591.t25 a_52635_49681.t9 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X360 VDD.t4517 VDD.t4516 VDD.t4517 VDD.t2814 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X361 a_63161_n5344.t1 a_64243_n1756.t1 a_66058_7563# VSS.t411 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X362 VSS.t3464 VSS.t3463 VSS.t3464 VSS.t658 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X363 VDD.t4515 VDD.t4514 VDD.t4515 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X364 VSS.t3462 VSS.t3461 VSS.t3462 VSS.t412 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X365 VDD.t4513 VDD.t4512 VDD.t4513 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X366 OUT.t97 a_35922_19591.t26 a_52635_49681.t10 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X367 a_33249_35053.t4 a_33379_34917.t6 a_33249_48695.t21 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X368 VSS.t3460 VSS.t3459 VSS.t3460 VSS.t1437 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X369 VDD.t4511 VDD.t4510 VDD.t4511 VDD.t318 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X370 VSS.t3458 VSS.t3457 VSS.t3458 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X371 VSS.t3456 VSS.t3455 VSS.t3456 VSS.t800 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X372 VDD.t66 a_31699_20742.t55 a_33249_48695.t325 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X373 a_36008_4481.t0 a_30152_11614.t8 a_37934_7563# VSS.t323 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X374 a_33249_48695.t338 a_33379_34007.t9 a_33249_34067.t100 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X375 a_58851_n14215# a_50751_n19729.t89 a_58329_n14215# VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X376 a_102796_n30339# a_100992_n29313.t0 a_38097_n5342.t1 VSS.t383 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X377 a_96011_n36322.t1 a_83325_n29313.t1 a_95443_n35156# VDD.t2425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X378 a_98829_n8770# a_71281_n8397.t89 a_89033_n35156.t0 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X379 a_83725_n29181# a_83325_n29313.t0 a_83153_n35156.t10 VSS.t367 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X380 VSS.t3454 VSS.t3453 VSS.t3454 VSS.t323 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X381 VDD.t4509 VDD.t4508 VDD.t4509 VDD.t748 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X382 a_52635_34067.t15 a_35922_19591.t27 a_52635_48695.t77 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X383 a_77747_7563# a_77225_4481.t11 a_71496_10388.t0 VSS.t336 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X384 a_57977_n18700# a_50751_n19729.t90 a_57417_n18700# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X385 VSS.t3452 VSS.t3451 VSS.t3452 VSS.t24 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X386 VSS.t3450 VSS.t3449 VSS.t3450 VSS.t1349 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X387 VDD.t68 a_31699_20742.t56 a_33249_48695.t324 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X388 VSS.t3448 VSS.t3447 VSS.t3448 VSS.t1258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X389 VDD.t4507 VDD.t4506 VDD.t4507 VDD.t81 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X390 VDD.t4979 a_52635_34067.t69 a_52635_48695.t173 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X391 VSS.t3446 VSS.t3445 VSS.t3446 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X392 VDD.t4505 VDD.t4504 VDD.t4505 VDD.t758 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X393 VSS.t3444 VSS.t3443 VSS.t3444 VSS.t738 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X394 a_108636_13546# a_106830_10388.t9 a_106676_4481.t3 VDD.t525 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X395 VSS.t3442 VSS.t3441 VSS.t3442 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X396 VDD.t4503 VDD.t4502 VDD.t4503 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X397 VSS.t3440 VSS.t3439 VSS.t3440 VSS.t596 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X398 a_57417_n16009# a_50751_n19729.t91 a_56895_n16009.t1 VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X399 VDD.t4501 VDD.t4500 VDD.t4501 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X400 a_87433_n9675# a_71281_n10073.t82 a_86903_n9675# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X401 a_33787_n17801# a_31953_n19727.t88 a_33265_n18698# VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X402 a_96011_n36322.t1 a_83325_n29313.t1 a_95443_n33224# VDD.t2425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X403 VDD.t4499 VDD.t4498 VDD.t4499 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X404 VDD.t4497 VDD.t4496 VDD.t4497 VDD.t748 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X405 VSS.t3438 VSS.t3437 VSS.t3438 VSS.t503 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X406 VSS.t3436 VSS.t3435 VSS.t3436 VSS.t1069 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X407 VSS.t3434 VSS.t3433 VSS.t3434 VSS.t251 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X408 VDD.t4495 VDD.t4494 VDD.t4495 VDD.t1373 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X409 VDD.t4493 VDD.t4492 VDD.t4493 VDD.t81 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X410 VDD.t4491 VDD.t4490 VDD.t4491 VDD.t751 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X411 VSS.t91 a_31953_n19727.t66 a_31953_n19727.t67 VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X412 VSS.t3432 VSS.t3431 VSS.t3432 VSS.t254 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X413 VSS.t3430 VSS.t3429 VSS.t3430 VSS.t753 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X414 a_33249_34067.t99 a_33379_34007.t10 a_33249_48695.t115 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X415 VSS.t3428 VSS.t3427 VSS.t3428 VSS.t151 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X416 VSS.t3426 VSS.t3425 VSS.t3426 VSS.t325 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X417 VDD.t4489 VDD.t4488 VDD.t4489 VDD.t1551 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X418 a_108636_11614# a_106830_10388.t10 VSS.t331 VDD.t525 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X419 a_64243_n8932# a_50751_n19729.t92 a_63683_n8932# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X420 a_32128_7563# a_30324_4421.t0 a_31284_4481.t2 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X421 VDD.t4487 VDD.t4486 VDD.t4487 VDD.t2193 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X422 a_66551_n4447# a_50751_n19729.t93 a_66029_n6241# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X423 a_52635_48695.t172 a_52635_34067.t70 VDD.t4978 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X424 VSS.t3424 VSS.t3423 VSS.t3424 VSS.t768 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X425 VDD.t70 a_31699_20742.t57 a_33249_48695.t323 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X426 VSS.t3422 VSS.t3421 VSS.t3422 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X427 VSS.t3420 VSS.t3419 VSS.t3420 VSS.t300 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X428 a_30152_n35156.t9 a_30324_n29313.t0 a_32128_n28415# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X429 VDD.t4485 VDD.t4484 VDD.t4485 VDD.t728 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X430 a_33249_48695.t322 a_31699_20742.t58 VDD.t72 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X431 VSS.t3418 VSS.t3417 VSS.t3418 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X432 a_52635_48695.t171 a_52635_34067.t71 VDD.t4977 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X433 VDD.t74 a_31699_20742.t59 a_33249_48695.t321 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X434 VDD.t4976 a_52635_34067.t72 a_52635_49681.t173 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X435 VDD.t4483 VDD.t4482 VDD.t4483 VDD.t751 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X436 VSS.t3416 VSS.t3415 VSS.t3416 VSS.t765 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X437 VDD.t4481 VDD.t4480 VDD.t4481 VDD.t37 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X438 VSS.t3414 VSS.t3413 VSS.t3414 VSS.t1227 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X439 VSS.t3412 VSS.t3411 VSS.t3412 VSS.t1258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X440 a_33249_35053.t5 a_33379_34917.t7 a_33249_48695.t22 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X441 OUT.t96 a_35922_19591.t28 a_52635_49681.t11 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X442 a_48313_n7136# a_31953_n19727.t89 a_47753_n7136# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X443 a_45706_22884# a_35922_19591.t29 a_45138_22884# VDD.t401 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X444 VSS.t417 a_112559_n29181.t11 a_113081_n28415# VSS.t416 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X445 a_107339_n6960# a_71281_n8397.t90 a_106501_n4245# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X446 VSS.t3410 VSS.t3409 VSS.t3410 VSS.t689 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X447 VDD.t4479 VDD.t4478 VDD.t4479 VDD.t123 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X448 VDD.t4477 VDD.t4476 VDD.t4477 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X449 a_49755_12380# a_47819_10448.t11 VDD.t499 VDD.t498 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X450 VDD.t4975 a_52635_34067.t73 a_52635_48695.t170 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X451 VSS.t3408 VSS.t3407 VSS.t3408 VSS.t1311 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X452 VSS.t3406 VSS.t3405 VSS.t3406 VSS.t1308 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X453 VSS.t3404 VSS.t3403 VSS.t3404 VSS.t581 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X454 a_43848_13546# a_30324_4421.t1 a_43010_10448.t2 VDD.t293 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X455 VDD.t4475 VDD.t4474 VDD.t4475 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X456 VDD.t4473 VDD.t4472 VDD.t4473 VDD.t2164 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X457 VDD.t4471 VDD.t4470 VDD.t4471 VDD.t728 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X458 a_47819_n36322.t5 a_39179_n19595.t0 a_49795_n27257# VSS.t282 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X459 VSS.t3402 VSS.t3401 VSS.t3402 VSS.t620 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X460 a_93131_n8770# a_71281_n10073.t83 VDD.t310 VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X461 VDD.t4469 VDD.t4468 VDD.t4469 VDD.t2159 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X462 VSS.t279 a_53829_n36382.t11 a_54229_n34390# VDD.t420 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X463 a_35502_25545.t2 a_31699_20742.t60 VDD.t75 VDD.t15 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X464 VSS.t3400 VSS.t3399 VSS.t3400 VSS.t676 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X465 VSS.t3398 VSS.t3397 VSS.t3398 VSS.t1299 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X466 a_33249_35053.t139 a_35502_25545.t30 VSS.t200 VSS.t142 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X467 a_84017_n17715.t2 a_83325_4421.t1 a_95443_12380# VDD.t501 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X468 VDD.t4467 VDD.t4466 VDD.t4467 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X469 OUT.t95 a_35922_19591.t30 a_52635_49681.t12 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X470 VSS.t3396 VSS.t3395 VSS.t3396 VSS.t105 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X471 VSS.t3394 VSS.t3393 VSS.t3394 VSS.t1292 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X472 VSS.t3392 VSS.t3391 VSS.t3392 VSS.t312 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X473 VDD.t4465 VDD.t4464 VDD.t4465 VDD.t2146 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X474 VSS.t3390 VSS.t3389 VSS.t3390 VSS.t614 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X475 VSS.t3388 VSS.t3387 VSS.t3388 VSS.t327 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X476 VDD.t464 a_71281_n8397.t68 a_71281_n8397.t69 VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X477 a_105365_n1530# a_71281_n8397.t91 a_104527_n1530# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X478 OUT.t94 a_35922_19591.t31 a_52635_49681.t13 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X479 VDD.t77 a_31699_20742.t61 a_33249_48695.t320 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X480 a_43848_11614# a_30324_4421.t1 a_43010_10448.t1 VDD.t293 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X481 a_35502_25545.t3 a_31699_20742.t62 VDD.t78 VDD.t30 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X482 a_38619_n12419# a_31953_n19727.t90 a_38097_n13316# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X483 VDD.t4974 a_52635_34067.t74 a_52635_48695.t169 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X484 VSS.t3386 VSS.t3385 VSS.t3386 VSS.t147 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X485 a_105933_n15000# a_71281_n8397.t92 a_105365_n15000# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X486 VSS.t3384 VSS.t3383 VSS.t3384 VSS.t326 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X487 VSS.t3382 VSS.t3381 VSS.t3382 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X488 a_90935_n30339# a_83153_n36322.t8 a_83325_n29313.t0 VSS.t457 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X489 VDD.t4973 a_52635_34067.t75 a_52635_48695.t168 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X490 VSS.t246 a_50751_n19729.t66 a_50751_n19729.t67 VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X491 VDD.t4463 VDD.t4462 VDD.t4463 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X492 a_47819_n36322.t3 a_47819_n35156.t11 a_49755_n35156# VDD.t2328 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X493 VDD.t4461 VDD.t4460 VDD.t4461 VDD.t2131 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X494 a_52635_49681.t172 a_52635_34067.t76 VDD.t4972 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X495 VDD.t4459 VDD.t4458 VDD.t4459 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X496 VSS.t3380 VSS.t3379 VSS.t3380 VSS.t299 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X497 VDD.t4457 VDD.t4456 VDD.t4457 VDD.t652 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X498 VDD.t4971 a_52635_34067.t77 a_52635_49681.t171 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X499 a_101392_n27257# a_100992_n29313.t1 a_100820_n35156.t1 VSS.t381 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X500 VDD.t4455 VDD.t4454 VDD.t4455 VDD.t2731 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X501 a_41891_n29181.t10 a_41891_n29181.t9 a_43817_n28415# VSS.t181 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X502 a_83153_10448.t9 a_83153_10448.t8 a_85089_13546# VDD.t647 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X503 a_47991_4421.t0 a_47819_11614.t8 a_54197_7563# VSS.t327 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X504 VDD.t4453 VDD.t4452 VDD.t4453 VDD.t527 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X505 VDD.t4451 VDD.t4450 VDD.t4451 VDD.t3614 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X506 VDD.t4449 VDD.t4448 VDD.t4449 VDD.t2575 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X507 VDD.t4447 VDD.t4446 VDD.t4447 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X508 a_63683_n19597# a_50751_n19729.t94 a_63161_n19597# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X509 VSS.t3378 VSS.t3377 VSS.t3378 VSS.t643 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X510 a_52635_48695.t76 a_35922_19591.t32 a_52635_34067.t16 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X511 VDD.t4445 VDD.t4444 VDD.t4445 VDD.t2572 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X512 a_106501_n6960# a_71281_n8397.t93 a_105933_n6960# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X513 a_104527_n17715# a_71281_n8397.t94 a_103997_n16810# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X514 a_71281_n8397.t67 a_71281_n8397.t66 VDD.t463 VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X515 a_58851_n1756# a_50751_n19729.t95 a_57977_n5344.t1 VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X516 VDD.t4443 VDD.t4442 VDD.t4443 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X517 OUT.t93 a_35922_19591.t33 a_52635_49681.t14 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X518 a_104527_n15000# a_71281_n8397.t95 a_103997_n15905# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X519 a_47819_n36322.t2 a_47819_n35156.t12 a_49755_n33224# VDD.t2328 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X520 VDD.t4441 VDD.t4440 VDD.t4441 VDD.t623 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X521 a_44885_n5342# a_31953_n19727.t91 VSS.t102 VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X522 VDD.t4439 VDD.t4438 VDD.t4439 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X523 VDD.t4437 VDD.t4436 VDD.t4437 VDD.t497 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X524 a_112199_n18620# a_71281_n8397.t96 a_111631_n18620# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X525 VDD.t4435 VDD.t4434 VDD.t4435 VDD.t1869 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X526 VDD.t4433 VDD.t4432 VDD.t4433 VDD.t498 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X527 VDD.t4431 VDD.t4430 VDD.t4431 VDD.t652 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X528 VSS.t3376 VSS.t3375 VSS.t3376 VSS.t533 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X529 OUT.t18 a_35502_24538.t26 a_33249_35053.t89 VSS.t162 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X530 VDD.t4800 a_47819_n35156.t13 a_48349_n35156# VDD.t2291 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X531 a_33249_48695.t116 a_33379_34007.t11 a_33249_34067.t98 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X532 VSS.t3374 VSS.t3373 VSS.t3374 VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X533 a_104527_n8770# a_71281_n8397.t97 a_103997_n8770.t0 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X534 VDD.t4429 VDD.t4428 VDD.t4429 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X535 a_83153_10448.t11 a_83153_10448.t10 a_85089_11614# VDD.t647 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X536 a_31953_n19727.t65 a_31953_n19727.t64 VSS.t90 VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X537 a_52635_49681.t15 a_35922_19591.t34 OUT.t92 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X538 VDD.t4427 VDD.t4426 VDD.t4427 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X539 VDD.t4425 VDD.t4424 VDD.t4425 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X540 VSS.t3372 VSS.t3371 VSS.t3372 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X541 a_111631_n9675# a_71281_n8397.t98 a_111063_n9675# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X542 a_47753_n14213# a_31953_n19727.t92 a_47231_n14213# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X543 VSS.t3370 VSS.t3369 VSS.t3370 VSS.t984 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X544 VSS.t3368 VSS.t3367 VSS.t3368 VSS.t686 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X545 VDD.t4423 VDD.t4422 VDD.t4423 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X546 a_46879_n19595# a_31953_n19727.t93 a_46319_n18698# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X547 VDD.t80 a_31699_20742.t63 a_33249_48695.t319 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X548 VDD.t4421 VDD.t4420 VDD.t4421 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X549 a_49795_4481# a_47991_5507.t0 a_48951_4481.t2 VSS.t281 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X550 VDD.t4970 a_52635_34067.t78 a_52635_48695.t167 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X551 a_83709_n19525# a_71281_n10073.t84 a_83141_n19525# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X552 VDD.t4419 VDD.t4418 VDD.t4419 VDD.t394 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X553 a_101350_n36322# a_100820_n35156.t12 a_100820_n36322.t1 VDD.t529 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X554 VSS.t3366 VSS.t3365 VSS.t3366 VSS.t558 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X555 VDD.t4417 VDD.t4416 VDD.t4417 VDD.t2103 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X556 VDD.t4415 VDD.t4414 VDD.t4415 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X557 VDD.t4413 VDD.t4412 VDD.t4413 VDD.t642 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X558 a_52635_34067.t17 a_35922_19591.t35 a_52635_48695.t75 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X559 VSS.t3364 VSS.t3363 VSS.t3364 VSS.t873 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X560 VDD.t4411 VDD.t4410 VDD.t4411 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X561 VSS.t3362 VSS.t3361 VSS.t3362 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X562 a_33249_48695.t318 a_31699_20742.t64 VDD.t82 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X563 VDD.t4409 VDD.t4408 VDD.t4409 VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X564 VDD.t4969 a_52635_34067.t79 a_52635_49681.t170 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X565 VDD.t4407 VDD.t4406 VDD.t4407 VDD.t2100 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X566 a_42047_n4445# a_31953_n19727.t94 a_41487_n4445# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X567 VDD.t4405 VDD.t4404 VDD.t4405 VDD.t629 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X568 VSS.t3360 VSS.t3359 VSS.t3360 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X569 a_106830_10388.t6 a_112559_4481.t12 a_114485_6405# VSS.t286 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X570 VDD.t4801 a_47819_n35156.t14 a_48349_n33224# VDD.t2291 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X571 VSS.t178 a_41891_4481.t12 a_42413_6405# VSS.t171 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X572 a_114485_n27257# a_112559_n29181.t12 VSS.t419 VSS.t418 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X573 a_30152_n35156.t7 a_30152_n35156.t6 a_32088_n36322# VDD.t554 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X574 a_54019_n17803# a_50751_n19729.t96 a_53497_n18700# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X575 a_71896_n35156# a_71496_n36382.t10 a_71366_n35156.t3 VDD.t2254 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X576 a_81735_n7865# a_71281_n10073.t85 a_81205_n7865# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X577 a_105933_n20430# a_71281_n8397.t99 a_105365_n20430# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X578 VDD.t4403 VDD.t4402 VDD.t4403 VDD.t647 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X579 VSS.t3358 VSS.t3357 VSS.t3358 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X580 a_59558_n29181.t9 a_47991_n29313.t1 a_61515_n34390# VDD.t547 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X581 a_32913_n6239# a_31953_n19727.t95 a_32353_n6239# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X582 VDD.t4401 VDD.t4400 VDD.t4401 VDD.t1613 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X583 a_33249_34067.t97 a_33379_34007.t12 a_33249_48695.t110 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X584 a_54197_n30339# a_47819_n36322.t8 a_53675_n30339.t1 VSS.t329 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X585 VDD.t4399 VDD.t4398 VDD.t4399 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X586 a_98829_n7865# a_71281_n8397.t100 a_98299_n7865# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X587 VSS.t3356 VSS.t3355 VSS.t3356 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X588 VDD.t4397 VDD.t4396 VDD.t4397 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X589 VDD.t4395 VDD.t4394 VDD.t4395 VDD.t602 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X590 VSS.t3354 VSS.t3353 VSS.t3354 VSS.t427 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X591 a_33249_34067.t96 a_33379_34007.t13 a_33249_48695.t111 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X592 VDD.t4393 VDD.t4392 VDD.t4393 VDD.t65 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X593 VSS.t3352 VSS.t3351 VSS.t3352 VSS.t704 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X594 VDD.t4391 VDD.t4390 VDD.t4391 VDD.t629 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X595 a_33249_48695.t317 a_31699_20742.t65 VDD.t83 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X596 VSS.t3350 VSS.t3349 VSS.t3350 VSS.t366 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X597 VSS.t3348 VSS.t3347 VSS.t3348 VSS.t1600 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X598 a_71896_n33224# a_71496_n36382.t11 a_53699_n36322.t0 VDD.t2254 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X599 VSS.t3346 VSS.t3345 VSS.t3346 VSS.t1249 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X600 VSS.t3344 VSS.t3343 VSS.t3344 VSS.t695 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X601 VDD.t4389 VDD.t4388 VDD.t4389 VDD.t1820 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X602 a_96849_n35156# a_89033_n35156.t5 a_96011_n36322.t3 VDD.t2243 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X603 VDD.t4387 VDD.t4386 VDD.t4387 VDD.t61 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X604 VSS.t3342 VSS.t3341 VSS.t3342 VSS.t649 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X605 VSS.t3340 VSS.t3339 VSS.t3340 VSS.t1320 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X606 a_33249_35053.t6 a_33379_34917.t8 a_33249_48695.t23 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X607 a_84547_n6960# a_71281_n10073.t86 a_83709_n6960# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X608 VSS.t3338 VSS.t3337 VSS.t3338 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X609 a_104527_n20430# a_71281_n8397.t101 a_53699_n35156.t0 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X610 a_93131_n19525# a_71281_n10073.t87 a_92601_n19525# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X611 a_52635_48695.t166 a_52635_34067.t80 VDD.t4968 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X612 VDD.t4385 VDD.t4384 VDD.t4385 VDD.t2082 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X613 a_60677_n36322.t1 a_53699_n35156.t5 a_60109_n34390# VDD.t546 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X614 a_56895_n16009.t0 a_100992_4421.t0 a_101392_6405# VSS.t174 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X615 VSS.t3336 VSS.t3335 VSS.t3336 VSS.t681 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X616 a_88271_n19525# a_71281_n10073.t88 a_87433_n19525# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X617 VDD.t4383 VDD.t4382 VDD.t4383 VDD.t2079 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X618 VSS.t3334 VSS.t3333 VSS.t3334 VSS.t252 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X619 VDD.t4381 VDD.t4380 VDD.t4381 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X620 VDD.t4791 a_30152_n35156.t13 a_30682_n35156# VDD.t552 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X621 VDD.t520 a_47819_n36322.t9 a_55601_n29181# VSS.t328 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X622 a_108602_n30339# a_100820_n36322.t9 a_100992_n29313.t0 VSS.t351 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X623 a_45445_n14213# a_31953_n19727.t96 a_44885_n13316# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X624 VSS.t3332 VSS.t3331 VSS.t3332 VSS.t260 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X625 VSS.t3330 VSS.t3329 VSS.t3330 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X626 VDD.t4379 VDD.t4378 VDD.t4379 VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X627 a_113081_6405# a_112559_4481.t9 a_112559_4481.t10 VSS.t285 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X628 a_52635_34067.t18 a_35922_19591.t36 a_52635_48695.t74 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X629 a_96849_n33224# a_89033_n35156.t6 a_96011_n36322.t1 VDD.t2243 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X630 VSS.t3328 VSS.t3327 VSS.t3328 VSS.t726 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X631 a_100235_n14095# a_71281_n8397.t102 a_99667_n14095# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X632 a_65486_11614.t5 a_64243_n1756.t1 a_67462_6405# VSS.t413 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X633 VDD.t4377 VDD.t4376 VDD.t4377 VDD.t1789 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X634 VSS.t3326 VSS.t3325 VSS.t3326 VSS.t503 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X635 a_66551_n13318# a_50751_n19729.t97 a_66029_n14215# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X636 a_39179_n3548# a_31953_n19727.t97 a_38619_n2651# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X637 a_42413_6405# a_41891_4481.t2 a_41891_4481.t3 VSS.t177 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X638 VDD.t4375 VDD.t4374 VDD.t4375 VDD.t26 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X639 VSS.t3324 VSS.t3323 VSS.t3324 VSS.t686 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X640 a_32353_n14213# a_31953_n19727.t98 a_31831_n15110# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X641 VDD.t4373 VDD.t4372 VDD.t4373 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X642 a_79151_6405# a_77225_4481.t12 VSS.t338 VSS.t337 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X643 VDD.t4371 VDD.t4370 VDD.t4371 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X644 VDD.t4757 a_30152_n35156.t14 a_30682_n33224# VDD.t552 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X645 a_54229_13546# a_53829_10388.t8 a_53699_13546.t1 VDD.t3679 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X646 OUT.t91 a_35922_19591.t37 a_52635_49681.t16 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X647 a_53699_n35156.t4 a_53829_n36382.t12 a_55635_n35156# VDD.t334 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X648 VDD.t4369 VDD.t4368 VDD.t4369 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X649 VDD.t4367 VDD.t4366 VDD.t4367 VDD.t2064 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X650 a_32353_n1754# a_31953_n19727.t99 a_31831_n2651# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X651 VSS.t3322 VSS.t3321 VSS.t3322 VSS.t428 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X652 VDD.t4365 VDD.t4364 VDD.t4365 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X653 VSS.t3320 VSS.t3319 VSS.t3320 VSS.t614 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X654 VSS.t3318 VSS.t3317 VSS.t3318 VSS.t9 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X655 VSS.t3316 VSS.t3315 VSS.t3316 VSS.t163 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X656 VDD.t4363 VDD.t4362 VDD.t4363 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X657 a_34347_n2651# a_31953_n19727.t100 a_33787_n1754# VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X658 a_90935_4481# a_83153_11614.t11 a_83325_4421.t0 VSS.t401 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X659 a_41487_n16904# a_31953_n19727.t101 a_40965_n16904# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X660 a_35781_n7136# a_31953_n19727.t102 a_35221_n6239# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X661 a_33249_48695.t316 a_31699_20742.t66 VDD.t84 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X662 VSS.t3314 VSS.t3313 VSS.t3314 VSS.t913 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X663 a_52635_49681.t169 a_52635_34067.t81 VDD.t4967 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X664 a_52635_34067.t19 a_35922_19591.t38 a_52635_48695.t73 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X665 a_113037_n17715# a_71281_n8397.t103 a_78344_n36322.t0 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X666 VDD.t4361 VDD.t4360 VDD.t4361 VDD.t35 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X667 a_98829_n14095# a_71281_n8397.t104 VDD.t472 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X668 a_93131_n7865# a_71281_n10073.t89 a_92601_n7865# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X669 a_50751_n19729.t65 a_50751_n19729.t64 VSS.t245 VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X670 VSS.t3312 VSS.t3311 VSS.t3312 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X671 VDD.t4359 VDD.t4358 VDD.t4359 VDD.t1422 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X672 a_52635_34067.t20 a_35922_19591.t39 a_52635_48695.t72 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X673 a_113037_n15000# a_71281_n8397.t105 a_112199_n15000# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X674 a_33249_48695.t315 a_31699_20742.t67 VDD.t86 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X675 VDD.t4357 VDD.t4356 VDD.t4357 VDD.t2488 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X676 a_54229_11614# a_53829_10388.t9 a_53699_11614.t1 VDD.t3679 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X677 VSS.t3310 VSS.t3309 VSS.t3310 VSS.t447 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X678 a_52635_48695.t165 a_52635_34067.t82 VDD.t4966 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X679 a_53699_n36322.t3 a_53829_n36382.t13 a_55635_n33224# VDD.t334 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X680 VDD.t4355 VDD.t4354 VDD.t4355 VDD.t979 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X681 VSS.t3308 VSS.t3307 VSS.t3308 VSS.t1162 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X682 VDD.t87 a_31699_20742.t68 a_33249_48695.t314 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X683 a_83141_n18620# a_71281_n10073.t90 a_82573_n18620# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X684 VSS.t3306 VSS.t3305 VSS.t3306 VSS.t558 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X685 a_105365_n14095# a_71281_n8397.t106 a_104527_n14095# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X686 a_66058_4481# a_65658_4421.t1 a_65486_10448.t10 VSS.t410 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X687 VDD.t4353 VDD.t4352 VDD.t4353 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X688 VDD.t4351 VDD.t4350 VDD.t4351 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X689 a_83153_n35156.t9 a_83325_n29313.t0 a_85129_n30339# VSS.t365 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X690 a_105933_n15905# a_71281_n8397.t107 a_105365_n15905# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X691 a_72603_n10073# I1N.t4 a_71281_n10073.t1 VSS.t302 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X692 a_95105_n13190# a_71281_n10073.t91 a_94537_n13190# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X693 VDD.t88 a_31699_20742.t69 a_33249_48695.t313 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X694 VDD.t4349 VDD.t4348 VDD.t4349 VDD.t1422 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X695 a_52635_34067.t21 a_35922_19591.t40 a_52635_48695.t71 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X696 a_89715_n16810.t1 a_71281_n10073.t92 a_89407_n13190# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X697 VDD.t4347 VDD.t4346 VDD.t4347 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X698 VDD.t4345 VDD.t4344 VDD.t4345 VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X699 a_57417_n15112# a_50751_n19729.t98 a_56895_n15112# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X700 a_53829_n36382.t0 a_59558_n29181.t11 a_61484_n27257# VSS.t312 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X701 a_95943_n6960# a_71281_n10073.t93 a_95105_n6960# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X702 VDD.t4343 VDD.t4342 VDD.t4343 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X703 VSS.t3304 VSS.t3303 VSS.t3304 VSS.t99 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X704 a_44885_n16904# a_31953_n19727.t103 a_44363_n17801# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X705 VDD.t44 a_31699_20742.t37 a_31699_20742.t38 VDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X706 VDD.t4341 VDD.t4340 VDD.t4341 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X707 VDD.t89 a_31699_20742.t70 a_33249_48695.t312 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X708 VDD.t4339 VDD.t4338 VDD.t4339 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X709 a_52635_34067.t22 a_35922_19591.t41 a_52635_48695.t70 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X710 OUT.t90 a_35922_19591.t42 a_52635_49681.t17 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X711 VSS.t3302 VSS.t3301 VSS.t3302 VSS.t63 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X712 a_81735_n18620# a_71281_n10073.t94 a_81205_n19525# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X713 VDD.t4337 VDD.t4336 VDD.t4337 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X714 VSS.t89 a_31953_n19727.t62 a_31953_n19727.t63 VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X715 VSS.t3300 VSS.t3299 VSS.t3300 VSS.t620 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X716 VDD.t4335 VDD.t4334 VDD.t4335 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X717 a_57417_n4447# a_50751_n19729.t99 a_56895_n4447# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X718 VDD.t4333 VDD.t4332 VDD.t4333 VDD.t642 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X719 a_33249_35053.t7 a_33379_34917.t9 a_33249_48695.t24 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X720 a_93969_n8770# a_71281_n10073.t95 a_93131_n8770# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X721 VDD.t4331 VDD.t4330 VDD.t4331 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X722 VDD.t4329 VDD.t4328 VDD.t4329 VDD.t1517 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X723 a_104527_n15905# a_71281_n8397.t108 a_103997_n15905# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X724 a_112199_n4245# a_71281_n8397.t109 a_111631_n4245# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X725 VSS.t3298 VSS.t3297 VSS.t3298 VSS.t1261 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X726 VDD.t4327 VDD.t4326 VDD.t4327 VDD.t947 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X727 VDD.t4325 VDD.t4324 VDD.t4325 VDD.t1376 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X728 VDD.t4766 a_30152_10448.t12 a_30682_12380# VDD.t13 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X729 VDD.t4323 VDD.t4322 VDD.t4323 VDD.t1373 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X730 a_51151_n13318# a_50751_n19729.t100 a_50629_n13318# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X731 a_71896_13546# a_71496_10388.t10 a_71366_13546.t3 VDD.t488 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X732 VDD.t4321 VDD.t4320 VDD.t4321 VDD.t1368 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X733 VSS.t3296 VSS.t3295 VSS.t3296 VSS.t800 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X734 a_94537_n3340# a_71281_n10073.t96 a_93969_n3340# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X735 a_96849_12380# a_81205_n14095.t3 a_84017_n17715.t0 VDD.t502 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X736 VDD.t4319 VDD.t4318 VDD.t4319 VDD.t81 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X737 a_42413_n30339# a_41891_n29181.t12 a_36162_n36382.t5 VSS.t177 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X738 a_88839_n13190# a_71281_n10073.t97 a_88271_n13190# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X739 a_73302_10448# a_71496_10388.t11 a_71342_7563.t2 VDD.t491 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X740 VDD.t4317 VDD.t4316 VDD.t4317 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X741 VDD.t462 a_71281_n8397.t64 a_71281_n8397.t65 VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X742 VDD.t4315 VDD.t4314 VDD.t4315 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X743 VSS.t3294 VSS.t3293 VSS.t3294 VSS.t609 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X744 a_104527_n7865# a_71281_n8397.t110 a_103997_n7865# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X745 a_52635_34067.t23 a_35922_19591.t43 a_52635_48695.t69 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X746 a_82573_n9675# a_71281_n10073.t98 a_81735_n9675# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X747 OUT.t89 a_35922_19591.t44 a_52635_49681.t18 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X748 a_75585_n9297# I1N.t5 VSS.t441 VSS.t303 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X749 VSS.t3292 VSS.t3291 VSS.t3292 VSS.t249 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X750 a_113037_n20430# a_71281_n8397.t111 a_112199_n20430# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X751 a_65486_n36322.t0 a_65486_n35156.t13 a_67422_n35156# VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X752 VDD.t4313 VDD.t4312 VDD.t4313 VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X753 VDD.t4311 VDD.t4310 VDD.t4311 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X754 VDD.t4309 VDD.t4308 VDD.t4309 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X755 a_50751_n19729.t63 a_50751_n19729.t62 VSS.t244 VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X756 OUT.t88 a_35922_19591.t45 a_52635_49681.t19 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X757 VDD.t4307 VDD.t4306 VDD.t4307 VDD.t1357 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X758 a_99667_n9675# a_71281_n8397.t112 a_98829_n9675# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X759 a_71896_11614# a_71496_10388.t12 a_71366_11614.t0 VDD.t488 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X760 a_102756_n34390# a_100820_n35156.t13 VDD.t531 VDD.t530 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X761 a_34347_n13316# a_31953_n19727.t104 a_33787_n12419# VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X762 a_52635_48695.t68 a_35922_19591.t46 a_52635_34067.t24 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X763 a_33249_35053.t8 a_33379_34917.t10 a_33249_48695.t25 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X764 a_95414_n28415# a_94892_n29181.t11 a_89163_n36382.t4 VSS.t446 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X765 VDD.t4305 VDD.t4304 VDD.t4305 VDD.t1352 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X766 a_94892_n29181.t3 a_94892_n29181.t2 a_96818_n30339# VSS.t445 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X767 a_33249_34067.t95 a_33379_34007.t14 a_33249_48695.t333 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X768 VSS.t3290 VSS.t3289 VSS.t3290 VSS.t984 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X769 VSS.t3288 VSS.t3287 VSS.t3288 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X770 VDD.t4303 VDD.t4302 VDD.t4303 VDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X771 VDD.t4301 VDD.t4300 VDD.t4301 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X772 a_30152_10448.t2 a_30324_4421.t0 a_32128_5639# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X773 a_35502_25545.t4 a_31699_20742.t71 VDD.t90 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X774 a_33249_35053.t9 a_33379_34917.t11 a_33249_48695.t26 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X775 VDD.t508 a_47819_11614.t9 a_55601_6405# VSS.t328 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X776 VDD.t4299 VDD.t4298 VDD.t4299 VDD.t1713 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X777 VDD.t4297 VDD.t4296 VDD.t4297 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X778 VDD.t4295 VDD.t4294 VDD.t4295 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X779 VSS.t3286 VSS.t3285 VSS.t3286 VSS.t555 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X780 VDD.t360 a_71281_n10073.t72 a_71281_n10073.t73 VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X781 a_46319_n17801# a_31953_n19727.t105 a_45797_n18698# VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X782 a_65486_n36322.t1 a_65486_n35156.t14 a_67422_n33224# VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X783 a_40613_n8930# a_31953_n19727.t106 a_40053_n8033# VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X784 VDD.t4293 VDD.t4292 VDD.t4293 VDD.t2779 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X785 VSS.t3284 VSS.t3283 VSS.t3284 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X786 VDD.t4 a_65486_n35156.t15 a_66016_n35156# VDD.t1 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X787 VSS.t3282 VSS.t3281 VSS.t3282 VSS.t95 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X788 VSS.t3280 VSS.t3279 VSS.t3280 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X789 a_33249_35053.t10 a_33379_34917.t12 a_33249_48695.t27 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X790 VDD.t4291 VDD.t4290 VDD.t4291 VDD.t2561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X791 a_57977_n8932# a_50751_n19729.t101 a_57417_n8932# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X792 a_79182_13546# a_65658_4421.t2 a_78344_10448.t0 VDD.t575 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X793 VDD.t4289 VDD.t4288 VDD.t4289 VDD.t958 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X794 VSS.t3278 VSS.t3277 VSS.t3278 VSS.t1131 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X795 VSS.t3276 VSS.t3275 VSS.t3276 VSS.t1039 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X796 VSS.t3274 VSS.t3273 VSS.t3274 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X797 a_43817_n29181# a_41891_n29181.t13 VSS.t373 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X798 VDD.t4287 VDD.t4286 VDD.t4287 VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X799 VDD.t4285 VDD.t4284 VDD.t4285 VDD.t52 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X800 VDD.t4283 VDD.t4282 VDD.t4283 VDD.t901 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X801 a_33249_48695.t334 a_33379_34007.t15 a_33249_34067.t94 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X802 VDD.t91 a_31699_20742.t72 a_35502_24538.t22 VDD.t28 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X803 VSS.t3272 VSS.t3271 VSS.t3272 VSS.t150 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X804 VDD.t4281 VDD.t4280 VDD.t4281 VDD.t2779 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X805 VDD.t4279 VDD.t4278 VDD.t4279 VDD.t390 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X806 a_40053_n7136# a_31953_n19727.t107 a_39531_n8033# VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X807 a_49795_n29181# a_39179_n19595.t2 a_38097_n16007.t1 VSS.t281 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X808 VDD.t5 a_65486_n35156.t16 a_66016_n33224# VDD.t1 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X809 a_71281_n10073.t71 a_71281_n10073.t70 VDD.t370 VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X810 VDD.t4965 a_52635_34067.t83 a_52635_49681.t168 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X811 a_31831_n5342.t1 a_83325_n29313.t2 a_83725_n27257# VSS.t366 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X812 VSS.t3270 VSS.t3269 VSS.t3270 VSS.t22 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X813 VDD.t4964 a_52635_34067.t84 a_52635_48695.t164 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X814 OUT.t87 a_35922_19591.t47 a_52635_49681.t20 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X815 VDD.t4277 VDD.t4276 VDD.t4277 VDD.t15 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X816 VDD.t4275 VDD.t4274 VDD.t4275 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X817 VDD.t92 a_31699_20742.t73 a_33249_48695.t311 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X818 VSS.t3268 VSS.t3267 VSS.t3268 VSS.t1116 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X819 VSS.t3266 VSS.t3265 VSS.t3266 VSS.t469 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X820 a_60080_n30339# a_59558_n29181.t12 a_53829_n36382.t1 VSS.t313 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X821 a_54197_4481# a_47819_11614.t10 a_53675_4481.t0 VSS.t329 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X822 a_112199_n21335# a_71281_n8397.t113 a_111631_n21335# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X823 a_102796_5639# a_100992_4421.t0 a_56895_n16009.t0 VSS.t144 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X824 VSS.t3264 VSS.t3263 VSS.t3264 VSS.t11 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X825 VSS.t3262 VSS.t3261 VSS.t3262 VSS.t166 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X826 a_93969_n19525# a_71281_n10073.t99 a_93131_n19525# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X827 VDD.t4273 VDD.t4272 VDD.t4273 VDD.t958 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X828 VDD.t4271 VDD.t4270 VDD.t4271 VDD.t1919 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X829 a_79182_11614# a_65658_4421.t2 a_78344_10448.t1 VDD.t575 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X830 a_52635_34067.t25 a_35922_19591.t48 a_52635_48695.t67 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X831 OUT.t86 a_35922_19591.t49 a_52635_49681.t21 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X832 a_40613_n14213# a_31953_n19727.t108 a_41487_n16007# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X833 VDD.t4269 VDD.t4268 VDD.t4269 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X834 a_41487_n7136# a_31953_n19727.t109 a_40965_n8033# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X835 a_35781_n19595# a_31953_n19727.t110 a_35221_n18698# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X836 VSS.t3260 VSS.t3259 VSS.t3260 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X837 a_32088_n35156# a_30152_n35156.t15 VDD.t4790 VDD.t2091 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X838 a_35221_n6239# a_31953_n19727.t111 a_34699_n6239# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X839 a_53675_n30339.t2 a_53829_n36382.t14 a_54229_n36322# VDD.t420 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X840 a_55601_6405# a_47819_11614.t11 a_47991_5507.t0 VSS.t330 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X841 VDD.t4267 VDD.t4266 VDD.t4267 VDD.t1906 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X842 VDD.t4265 VDD.t4264 VDD.t4265 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X843 a_71281_n8397.t63 a_71281_n8397.t62 VDD.t461 VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X844 VSS.t3258 VSS.t3257 VSS.t3258 VSS.t596 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X845 VSS.t3256 VSS.t3255 VSS.t3256 VSS.t480 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X846 a_87433_n3340# a_71281_n10073.t100 a_86903_n4245# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X847 VSS.t3254 VSS.t3253 VSS.t3254 VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X848 VDD.t4263 VDD.t4262 VDD.t4263 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X849 a_106501_n15000# a_71281_n8397.t114 a_105933_n15000# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X850 a_89563_10448# a_89163_10388.t11 a_71366_13546.t1 VDD.t556 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X851 a_67422_10448# a_65486_10448.t13 VDD.t4750 VDD.t869 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X852 VSS.t3252 VSS.t3251 VSS.t3252 VSS.t593 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X853 a_36162_10388.t4 a_36032_11614.t5 a_43848_12380# VDD.t290 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X854 VDD.t4261 VDD.t4260 VDD.t4261 VDD.t548 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X855 VDD.t4259 VDD.t4258 VDD.t4259 VDD.t2352 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X856 VSS.t3250 VSS.t3249 VSS.t3250 VSS.t1621 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X857 VSS.t3248 VSS.t3247 VSS.t3248 VSS.t500 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X858 VSS.t3246 VSS.t3245 VSS.t3246 VSS.t686 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X859 a_43010_10448.t0 a_30324_4421.t1 a_42442_10448# VDD.t292 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X860 a_101641_n6960# a_71281_n8397.t115 a_100803_n6960# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X861 a_32088_n33224# a_30152_n35156.t16 VDD.t4747 VDD.t2091 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X862 VSS.t3244 VSS.t3243 VSS.t3244 VSS.t1827 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X863 VDD.t4257 VDD.t4256 VDD.t4257 VDD.t1895 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X864 VDD.t4255 VDD.t4254 VDD.t4255 VDD.t858 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X865 a_113037_n18620# a_71281_n8397.t116 a_112199_n15905# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X866 VSS.t243 a_50751_n19729.t60 a_50751_n19729.t61 VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X867 OUT.t85 a_35922_19591.t50 a_52635_49681.t22 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X868 VDD.t371 a_71281_n10073.t68 a_71281_n10073.t69 VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X869 a_32913_n5342.t0 a_31953_n19727.t112 a_32353_n5342# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X870 VSS.t3242 VSS.t3241 VSS.t3242 VSS.t483 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X871 a_52635_48695.t163 a_52635_34067.t85 VDD.t4963 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X872 VSS.t3240 VSS.t3239 VSS.t3240 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X873 a_33249_48695.t0 a_33379_34007.t16 a_33249_34067.t93 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X874 a_52635_34067.t0 a_35502_24538.t27 a_33249_34067.t16 VSS.t162 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X875 VDD.t4253 VDD.t4252 VDD.t4253 VDD.t1886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X876 VDD.t361 a_71281_n10073.t66 a_71281_n10073.t67 VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X877 a_50751_n19729.t59 a_50751_n19729.t58 VSS.t242 VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X878 VDD.t4251 VDD.t4250 VDD.t4251 VDD.t845 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X879 VDD.t4249 VDD.t4248 VDD.t4249 VDD.t670 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X880 VSS.t3238 VSS.t3237 VSS.t3238 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X881 VSS.t3236 VSS.t3235 VSS.t3236 VSS.t58 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X882 VDD.t4247 VDD.t4246 VDD.t4247 VDD.t831 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X883 VDD.t4245 VDD.t4244 VDD.t4245 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X884 a_71366_n35156.t2 a_71496_n36382.t12 a_73302_n35156# VDD.t2061 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X885 VDD.t4243 VDD.t4242 VDD.t4243 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X886 VDD.t4241 VDD.t4240 VDD.t4241 VDD.t816 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X887 a_45138_23609# a_35922_19591.t51 a_44608_22884# VDD.t404 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X888 VDD.t4239 VDD.t4238 VDD.t4239 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X889 VSS.t3234 VSS.t3233 VSS.t3234 VSS.t506 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X890 a_41891_4481.t5 a_41891_4481.t4 a_43817_7563# VSS.t181 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X891 VSS.t3232 VSS.t3231 VSS.t3232 VSS.t1162 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X892 VDD.t4237 VDD.t4236 VDD.t4237 VDD.t670 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X893 VDD.t4235 VDD.t4234 VDD.t4235 VDD.t2682 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X894 OUT.t84 a_35922_19591.t52 a_52635_49681.t23 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X895 VDD.t4233 VDD.t4232 VDD.t4233 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X896 VSS.t3230 VSS.t3229 VSS.t3230 VSS.t981 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X897 a_78344_n36322.t2 a_65658_n29313.t1 a_77776_n35156# VDD.t2046 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X898 VSS.t3228 VSS.t3227 VSS.t3228 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X899 a_66058_n29181# a_65658_n29313.t0 a_65486_n35156.t8 VSS.t410 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X900 VSS.t3226 VSS.t3225 VSS.t3226 VSS.t495 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X901 a_81735_n17715# a_71281_n10073.t101 a_81205_n21335# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X902 a_39179_n16007.t0 a_31953_n19727.t113 a_38619_n16007# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X903 a_33249_34067.t92 a_33379_34007.t17 a_33249_48695.t1 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X904 a_33249_48695.t310 a_31699_20742.t74 VDD.t93 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X905 a_71366_n36322.t3 a_71496_n36382.t13 a_73302_n33224# VDD.t2061 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X906 a_52635_49681.t167 a_52635_34067.t86 VDD.t4962 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X907 VDD.t4231 VDD.t4230 VDD.t4231 VDD.t639 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X908 a_93969_n7865# a_71281_n10073.t102 a_93131_n7865# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X909 a_33249_48695.t309 a_31699_20742.t75 VDD.t94 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X910 VSS.t3224 VSS.t3223 VSS.t3224 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X911 VSS.t88 a_31953_n19727.t60 a_31953_n19727.t61 VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X912 a_33249_34067.t91 a_33379_34007.t18 a_33249_48695.t120 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X913 VSS.t3222 VSS.t3221 VSS.t3222 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X914 VSS.t368 a_71496_n36382.t14 a_71896_n35156# VDD.t2023 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X915 a_48313_n2651# a_31953_n19727.t114 a_47753_n1754# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X916 a_106501_n20430# a_71281_n8397.t117 a_105933_n20430# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X917 a_33787_n13316# a_31953_n19727.t115 a_33265_n14213# VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X918 VSS.t3220 VSS.t3219 VSS.t3220 VSS.t154 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X919 a_66551_n12421# a_50751_n19729.t102 VSS.t261 VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X920 VSS.t3218 VSS.t3217 VSS.t3218 VSS.t539 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X921 a_60285_n16009# a_50751_n19729.t103 a_59411_n14215# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X922 a_94537_n2435# a_71281_n10073.t103 a_93969_n2435# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X923 VDD.t4229 VDD.t4228 VDD.t4229 VDD.t1852 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X924 VDD.t4227 VDD.t4226 VDD.t4227 VDD.t322 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X925 VSS.t3216 VSS.t3215 VSS.t3216 VSS.t149 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X926 a_45445_n6239# a_31953_n19727.t116 a_44885_n4445# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X927 VDD.t4225 VDD.t4224 VDD.t4225 VDD.t2682 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X928 a_78344_n36322.t2 a_65658_n29313.t1 a_77776_n33224# VDD.t2046 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X929 VSS.t3214 VSS.t3213 VSS.t3214 VSS.t536 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X930 VDD.t4223 VDD.t4222 VDD.t4223 VDD.t375 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X931 a_59558_n29181.t10 a_47991_n29313.t1 a_61515_n36322# VDD.t547 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X932 VDD.t4221 VDD.t4220 VDD.t4221 VDD.t1613 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X933 VDD.t4219 VDD.t4218 VDD.t4219 VDD.t795 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X934 VDD.t4217 VDD.t4216 VDD.t4217 VDD.t614 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X935 VDD.t4215 VDD.t4214 VDD.t4215 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X936 a_64243_n6241# a_50751_n19729.t104 a_63683_n4447# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X937 VDD.t4213 VDD.t4212 VDD.t4213 VDD.t639 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X938 a_51711_n19597# a_50751_n19729.t105 a_51151_n19597# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X939 a_100820_10448.t1 a_100992_4421.t0 a_102796_7563# VSS.t173 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X940 VDD.t4211 VDD.t4210 VDD.t4211 VDD.t497 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X941 a_31284_4481.t2 a_30324_5507.t1 a_30724_7563# VSS.t146 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X942 VSS.t3212 VSS.t3211 VSS.t3212 VSS.t416 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X943 VSS.t3210 VSS.t3209 VSS.t3210 VSS.t126 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X944 a_71342_n27257.t2 a_71496_n36382.t15 a_71896_n33224# VDD.t2023 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X945 a_33249_34067.t90 a_33379_34007.t19 a_33249_48695.t121 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X946 a_34347_n3548# a_31953_n19727.t117 a_35221_n5342# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X947 VSS.t3208 VSS.t3207 VSS.t3208 VSS.t148 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X948 a_89163_n36382.t2 a_89033_n35156.t7 a_96849_n35156# VDD.t1998 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X949 VSS.t3206 VSS.t3205 VSS.t3206 VSS.t483 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X950 a_40613_n3548# a_31953_n19727.t118 a_40053_n3548# VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X951 VDD.t4209 VDD.t4208 VDD.t4209 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X952 VDD.t4207 VDD.t4206 VDD.t4207 VDD.t695 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X953 a_83141_n21335# a_71281_n10073.t104 a_82573_n21335# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X954 VDD.t4205 VDD.t4204 VDD.t4205 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X955 a_50751_n19729.t57 a_50751_n19729.t56 VSS.t241 VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X956 VDD.t4203 VDD.t4202 VDD.t4203 VDD.t1826 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X957 a_52635_34067.t17 a_35922_19591.t53 a_52635_48695.t66 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X958 VDD.t4201 VDD.t4200 VDD.t4201 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X959 VDD.t4199 VDD.t4198 VDD.t4199 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X960 VDD.t4197 VDD.t4196 VDD.t4197 VDD.t1823 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X961 VSS.t3204 VSS.t3203 VSS.t3204 VSS.t464 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X962 a_52635_34067.t26 a_35922_19591.t54 a_52635_48695.t65 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X963 a_33249_34067.t89 a_33379_34007.t20 a_33249_48695.t122 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X964 a_111063_n8770# a_71281_n8397.t118 a_110225_n8770# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X965 VSS.t3202 VSS.t3201 VSS.t3202 VSS.t223 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X966 a_85129_5639# a_83325_4421.t0 a_50629_n16009.t0 VSS.t298 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X967 VDD.t4195 VDD.t4194 VDD.t4195 VDD.t614 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X968 VDD.t4193 VDD.t4192 VDD.t4193 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X969 a_43817_7563# a_41891_4481.t13 VSS.t192 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X970 VDD.t4191 VDD.t4190 VDD.t4191 VDD.t2234 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X971 VDD.t95 a_31699_20742.t76 a_33249_48695.t308 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X972 a_60677_n36322.t2 a_53699_n35156.t6 a_60109_n36322# VDD.t546 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X973 a_83709_n4245# a_71281_n10073.t105 a_83141_n4245# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X974 a_32088_12380# a_30152_10448.t13 VDD.t4767 VDD.t304 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X975 OUT.t83 a_35922_19591.t55 a_52635_49681.t24 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X976 a_38097_n5342.t1 a_39179_n8930.t1 a_101392_n30339# VSS.t384 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X977 VSS.t3200 VSS.t3199 VSS.t3200 VSS.t1042 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X978 a_111631_n3340# a_71281_n8397.t119 a_111063_n3340# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X979 VDD.t4189 VDD.t4188 VDD.t4189 VDD.t328 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X980 a_89163_n36382.t3 a_89033_n35156.t8 a_96849_n33224# VDD.t1998 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X981 VSS.t3198 VSS.t3197 VSS.t3198 VSS.t492 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X982 VSS.t3196 VSS.t3195 VSS.t3196 VSS.t326 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X983 VDD.t4187 VDD.t4186 VDD.t4187 VDD.t1212 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X984 VDD.t4185 VDD.t4184 VDD.t4185 VDD.t758 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X985 VDD.t4183 VDD.t4182 VDD.t4183 VDD.t2425 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X986 VSS.t3194 VSS.t3193 VSS.t3194 VSS.t952 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X987 a_81735_n21335# a_71281_n10073.t106 a_81205_n21335# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X988 VSS.t3192 VSS.t3191 VSS.t3192 VSS.t942 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X989 VDD.t4181 VDD.t4180 VDD.t4181 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X990 VDD.t4179 VDD.t4178 VDD.t4179 VDD.t1798 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X991 a_87433_n19525# a_71281_n10073.t107 a_86903_n19525# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X992 VSS.t3190 VSS.t3189 VSS.t3190 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X993 VSS.t3188 VSS.t3187 VSS.t3188 VSS.t223 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X994 VSS.t3186 VSS.t3185 VSS.t3186 VSS.t1030 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X995 a_101392_7563# a_57977_n12421.t0 a_100820_11614.t7 VSS.t175 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X996 a_33249_34067.t141 a_35502_25545.t31 VSS.t275 VSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X997 VSS.t3184 VSS.t3183 VSS.t3184 VSS.t181 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X998 VDD.t4177 VDD.t4176 VDD.t4177 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X999 a_81735_n1530# a_71281_n10073.t108 a_81205_n5150# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1000 a_33249_48695.t112 a_33379_34007.t21 a_33249_34067.t88 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1001 a_45445_n19595.t1 a_65486_n36322.t10 a_71864_n28415# VSS.t155 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1002 VDD.t4175 VDD.t4174 VDD.t4175 VDD.t758 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1003 VSS.t3182 VSS.t3181 VSS.t3182 VSS.t873 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1004 a_33249_35053.t11 a_33379_34917.t13 a_33249_48695.t28 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1005 a_30724_7563# a_30324_5507.t1 a_30152_11614.t1 VSS.t145 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1006 VDD.t4173 VDD.t4172 VDD.t4173 VDD.t1782 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1007 a_73268_n30339# a_65486_n36322.t11 a_65658_n29313.t0 VSS.t156 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1008 VDD.t4961 a_52635_34067.t87 a_52635_48695.t162 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1009 a_98829_n1530# a_71281_n8397.t120 a_98299_n5150# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1010 a_51151_n12421# a_50751_n19729.t106 a_50629_n13318# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1011 VDD.t4171 VDD.t4170 VDD.t4171 VDD.t1336 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1012 VDD.t4169 VDD.t4168 VDD.t4169 VDD.t1265 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1013 a_71281_n8397.t61 a_71281_n8397.t60 VDD.t460 VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1014 a_52635_49681.t166 a_52635_34067.t88 VDD.t4960 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1015 VDD.t4167 VDD.t4166 VDD.t4167 VDD.t751 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1016 VDD.t4165 VDD.t4164 VDD.t4165 VDD.t1341 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1017 a_65677_n17803# a_50751_n19729.t107 a_65117_n17803# VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1018 VDD.t4163 VDD.t4162 VDD.t4163 VDD.t748 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1019 VDD.t4161 VDD.t4160 VDD.t4161 VDD.t1186 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1020 a_33249_48695.t307 a_31699_20742.t77 VDD.t96 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1021 a_52635_49681.t165 a_52635_34067.t89 VDD.t4959 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1022 a_105933_n14095# a_71281_n8397.t121 a_105365_n14095# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1023 VSS.t3180 VSS.t3179 VSS.t3180 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1024 VDD.t4159 VDD.t4158 VDD.t4159 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1025 VDD.t4157 VDD.t4156 VDD.t4157 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1026 a_52635_48695.t161 a_52635_34067.t90 VDD.t4958 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1027 a_30724_n28415# a_30324_n30399.t1 a_30152_n36322.t2 VSS.t145 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1028 VSS.t3178 VSS.t3177 VSS.t3178 VSS.t103 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1029 a_106501_n15905# a_71281_n8397.t122 a_105933_n15905# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1030 a_61484_n29181# a_59558_n29181.t13 VSS.t315 VSS.t314 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1031 a_108636_10448# a_106830_10388.t11 a_106676_7563.t2 VDD.t525 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1032 a_33249_34067.t140 a_35502_25545.t32 VSS.t170 VSS.t33 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1033 VDD.t4155 VDD.t4154 VDD.t4155 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1034 a_87433_n2435# a_71281_n10073.t109 a_53699_11614.t2 VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1035 VDD.t4153 VDD.t4152 VDD.t4153 VDD.t1180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1036 VSS.t3176 VSS.t3175 VSS.t3176 VSS.t162 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1037 VDD.t4151 VDD.t4150 VDD.t4151 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1038 a_52635_48695.t160 a_52635_34067.t91 VDD.t4957 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1039 a_100820_n36322.t6 a_39179_n8930.t1 a_102796_n29181# VSS.t382 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1040 VDD.t4149 VDD.t4148 VDD.t4149 VDD.t728 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1041 VSS.t3174 VSS.t3173 VSS.t3174 VSS.t1003 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1042 VDD.t4147 VDD.t4146 VDD.t4147 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1043 VSS.t3172 VSS.t3171 VSS.t3172 VSS.t249 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1044 a_60285_n8932# a_50751_n19729.t108 a_57977_n8932# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1045 VDD.t4956 a_52635_34067.t92 a_52635_49681.t164 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1046 VDD.t4145 VDD.t4144 VDD.t4145 VDD.t1376 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1047 a_35221_n17801# a_31953_n19727.t119 a_34699_n18698# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1048 VDD.t4143 VDD.t4142 VDD.t4143 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1049 VDD.t459 a_71281_n8397.t58 a_71281_n8397.t59 VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1050 VSS.t3170 VSS.t3169 VSS.t3170 VSS.t842 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1051 VSS.t3168 VSS.t3167 VSS.t3168 VSS.t593 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1052 a_104527_n14095# a_71281_n8397.t123 VDD.t474 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1053 VDD.t4141 VDD.t4140 VDD.t4141 VDD.t428 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1054 VDD.t4139 VDD.t4138 VDD.t4139 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1055 a_95105_n4245# a_71281_n10073.t110 a_94537_n4245# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1056 a_33249_48695.t306 a_31699_20742.t78 VDD.t97 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1057 VDD.t4137 VDD.t4136 VDD.t4137 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1058 a_30324_n29313.t0 a_30152_n36322.t9 a_36530_n30339# VSS.t325 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1059 VDD.t4135 VDD.t4134 VDD.t4135 VDD.t1302 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1060 VSS.t3166 VSS.t3165 VSS.t3166 VSS.t839 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1061 VSS.t3164 VSS.t3163 VSS.t3164 VSS.t1069 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1062 VDD.t98 a_31699_20742.t79 a_33249_48695.t305 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1063 VDD.t4133 VDD.t4132 VDD.t4133 VDD.t73 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1064 VDD.t4131 VDD.t4130 VDD.t4131 VDD.t700 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1065 VDD.t4955 a_52635_34067.t93 a_52635_49681.t163 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1066 VDD.t4129 VDD.t4128 VDD.t4129 VDD.t1517 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1067 a_89407_n13190# a_71281_n10073.t111 a_88839_n13190# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1068 a_54019_n13318# a_50751_n19729.t109 a_53497_n14215# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1069 VSS.t3162 VSS.t3161 VSS.t3162 VSS.t1366 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1070 VSS.t3160 VSS.t3159 VSS.t3160 VSS.t95 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1071 VDD.t4127 VDD.t4126 VDD.t4127 VDD.t2779 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1072 VSS.t3158 VSS.t3157 VSS.t3158 VSS.t66 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1073 VDD.t100 a_31699_20742.t80 a_33249_48695.t304 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1074 a_103997_n8770.t1 a_106830_n36382.t8 a_108636_n34390# VDD.t1293 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1075 VDD.t4125 VDD.t4124 VDD.t4125 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1076 a_36008_7563.t1 a_36162_10388.t8 a_36562_13546# VDD.t3614 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1077 VDD.t4123 VDD.t4122 VDD.t4123 VDD.t2575 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1078 VDD.t4121 VDD.t4120 VDD.t4121 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1079 a_100803_n13190# a_71281_n8397.t124 a_100235_n13190# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1080 a_32913_n8930.t1 a_83153_n36322.t9 a_89531_n28415# VSS.t458 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1081 VDD.t4119 VDD.t4118 VDD.t4119 VDD.t2572 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1082 VDD.t4954 a_52635_34067.t94 a_52635_48695.t159 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1083 a_40613_n19595# a_31953_n19727.t120 a_40053_n19595# VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1084 VSS.t3156 VSS.t3155 VSS.t3156 VSS.t542 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1085 a_93131_n1530# a_71281_n10073.t112 a_92601_n5150# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1086 a_43848_10448# a_36032_11614.t6 a_43010_10448.t0 VDD.t293 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1087 VDD.t4117 VDD.t4116 VDD.t4117 VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1088 a_107198_n29181# a_100820_n36322.t10 VDD.t540 VSS.t352 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1089 a_83325_4421.t0 a_83153_11614.t12 a_89531_7563# VSS.t399 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1090 VDD.t4115 VDD.t4114 VDD.t4115 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1091 a_73268_5639# a_65486_11614.t8 a_64243_n1756.t1 VSS.t426 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1092 VDD.t4113 VDD.t4112 VDD.t4113 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1093 VDD.t4111 VDD.t4110 VDD.t4111 VDD.t2328 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1094 VDD.t4109 VDD.t4108 VDD.t4109 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1095 VSS.t277 a_71496_10388.t13 a_71896_12380# VDD.t489 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1096 VSS.t3154 VSS.t3153 VSS.t3154 VSS.t1827 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1097 VDD.t101 a_31699_20742.t81 a_35502_25545.t5 VDD.t37 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1098 a_52635_34067.t1 a_35502_24538.t28 a_33249_34067.t15 VSS.t163 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1099 VDD.t4107 VDD.t4106 VDD.t4107 VDD.t291 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1100 a_102756_n36322# a_100820_n35156.t14 VDD.t532 VDD.t530 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1101 a_52635_34067.t22 a_35922_19591.t56 a_52635_48695.t64 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1102 VSS.t3152 VSS.t3151 VSS.t3152 VSS.t105 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1103 VSS.t3150 VSS.t3149 VSS.t3150 VSS.t726 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1104 VDD.t4105 VDD.t4104 VDD.t4105 VDD.t2122 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1105 VDD.t4103 VDD.t4102 VDD.t4103 VDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1106 VDD.t4101 VDD.t4100 VDD.t4101 VDD.t2575 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1107 VSS.t437 a_36162_10388.t9 a_36562_11614# VDD.t3614 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1108 VSS.t3148 VSS.t3147 VSS.t3148 VSS.t839 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1109 a_48391_n28415# a_39179_n19595.t0 a_47819_n36322.t6 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1110 a_35221_n5342# a_31953_n19727.t121 a_34347_n7136# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1111 VDD.t4099 VDD.t4098 VDD.t4099 VDD.t2572 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1112 VDD.t4097 VDD.t4096 VDD.t4097 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1113 VDD.t4095 VDD.t4094 VDD.t4095 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1114 a_32913_n16904# a_31953_n19727.t122 a_32353_n16904# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1115 a_33249_35053.t12 a_33379_34917.t14 a_33249_48695.t29 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1116 a_63683_n16009# a_50751_n19729.t110 VSS.t262 VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1117 VDD.t4093 VDD.t4092 VDD.t4093 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1118 VDD.t4091 VDD.t4090 VDD.t4091 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1119 VDD.t4770 a_83153_11614.t13 a_90935_6405# VSS.t398 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1120 VSS.t3146 VSS.t3145 VSS.t3146 VSS.t813 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1121 VDD.t4089 VDD.t4088 VDD.t4089 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1122 VDD.t102 a_31699_20742.t82 a_35502_24538.t21 VDD.t28 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1123 VSS.t3144 VSS.t3143 VSS.t3144 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1124 VDD.t4087 VDD.t4086 VDD.t4087 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1125 a_95943_n20430# a_71281_n10073.t113 a_95105_n19525# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1126 VDD.t4085 VDD.t4084 VDD.t4085 VDD.t1268 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1127 a_84547_n6055# a_71281_n10073.t114 a_43010_10448.t4 VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1128 a_52635_49681.t25 a_35922_19591.t57 OUT.t82 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1129 VDD.t4083 VDD.t4082 VDD.t4083 VDD.t2291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1130 VDD.t4081 VDD.t4080 VDD.t4081 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1131 VDD.t4079 VDD.t4078 VDD.t4079 VDD.t1710 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1132 a_51151_n8035# a_50751_n19729.t111 a_50629_n8932# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1133 a_30152_n36322.t4 a_30324_n30399.t1 a_32128_n27257# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1134 VDD.t4077 VDD.t4076 VDD.t4077 VDD.t1869 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1135 VDD.t4075 VDD.t4074 VDD.t4075 VDD.t652 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1136 VSS.t3142 VSS.t3141 VSS.t3142 VSS.t655 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1137 VDD.t103 a_31699_20742.t83 a_33249_48695.t303 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1138 VSS.t289 a_112559_4481.t13 a_113081_6405# VSS.t287 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1139 VDD.t4073 VDD.t4072 VDD.t4073 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1140 a_45706_24920# a_35922_19591.t58 a_45138_24920# VDD.t401 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X1141 VDD.t4953 a_52635_34067.t95 a_52635_48695.t158 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1142 a_83153_11614.t4 a_83153_10448.t12 a_85089_10448# VDD.t647 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1143 VDD.t4071 VDD.t4070 VDD.t4071 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1144 a_53145_n8932# a_50751_n19729.t112 a_52585_n8035# VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1145 VDD.t4069 VDD.t4068 VDD.t4069 VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1146 VDD.t4067 VDD.t4066 VDD.t4067 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1147 a_31953_n19727.t59 a_31953_n19727.t58 VSS.t87 VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1148 VSS.t420 a_112559_n29181.t13 a_113081_n27257# VSS.t416 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1149 VSS.t3140 VSS.t3139 VSS.t3140 VSS.t563 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1150 a_101350_n35156# a_100820_n35156.t5 a_100820_n35156.t6 VDD.t529 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1151 VSS.t3138 VSS.t3137 VSS.t3138 VSS.t386 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1152 VSS.t3136 VSS.t3135 VSS.t3136 VSS.t1543 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1153 a_111063_n7865# a_71281_n8397.t125 a_110225_n7865# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1154 a_33249_35053.t13 a_33379_34917.t15 a_33249_48695.t30 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1155 VSS.t3134 VSS.t3133 VSS.t3134 VSS.t536 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1156 a_71496_10388.t1 a_77225_4481.t13 a_79151_6405# VSS.t335 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1157 VSS.t3132 VSS.t3131 VSS.t3132 VSS.t460 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1158 VDD.t4065 VDD.t4064 VDD.t4065 VDD.t629 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1159 a_41487_n12419# a_31953_n19727.t123 a_39179_n12419# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1160 VSS.t3130 VSS.t3129 VSS.t3130 VSS.t429 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1161 VSS.t3128 VSS.t3127 VSS.t3128 VSS.t861 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1162 VDD.t4063 VDD.t4062 VDD.t4063 VDD.t1869 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1163 a_94537_n19525# a_71281_n10073.t115 a_93969_n19525# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1164 a_89531_7563# a_83153_11614.t14 a_89009_7563.t1 VSS.t400 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1165 VDD.t4061 VDD.t4060 VDD.t4061 VDD.t2254 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1166 a_104527_n1530# a_71281_n8397.t126 a_103997_n5150# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1167 a_33249_35053.t14 a_33379_34917.t16 a_33249_48695.t31 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1168 a_111631_n2435# a_71281_n8397.t127 a_111063_n2435# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1169 a_82573_n3340# a_71281_n10073.t116 a_81735_n3340# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1170 VDD.t4059 VDD.t4058 VDD.t4059 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1171 VDD.t4057 VDD.t4056 VDD.t4057 VDD.t1115 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1172 VSS.t203 a_35502_25545.t33 a_33249_34067.t139 VSS.t26 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1173 a_71496_10388.t4 a_71366_11614.t3 a_79182_12380# VDD.t1843 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1174 VSS.t3126 VSS.t3125 VSS.t3126 VSS.t514 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1175 a_30152_n36322.t0 a_30152_n35156.t17 a_32088_n35156# VDD.t554 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1176 a_33249_34067.t138 a_35502_25545.t34 VSS.t157 VSS.t134 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1177 a_33249_48695.t302 a_31699_20742.t84 VDD.t104 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1178 a_67462_n30339# a_65658_n29313.t0 a_44363_n16007.t2 VSS.t412 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1179 VDD.t4055 VDD.t4054 VDD.t4055 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1180 VDD.t4053 VDD.t4052 VDD.t4053 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1181 a_33249_48695.t32 a_33379_34917.t17 a_33249_35053.t15 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1182 a_47753_n4445# a_31953_n19727.t124 a_47231_n6239# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1183 a_99667_n3340# a_71281_n8397.t128 a_98829_n3340# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1184 a_101350_n33224# a_100820_n35156.t9 a_100820_n35156.t10 VDD.t529 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1185 a_48313_n19595# a_31953_n19727.t125 a_47753_n18698# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1186 a_33249_34067.t87 a_33379_34007.t22 a_33249_48695.t113 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1187 VSS.t3124 VSS.t3123 VSS.t3124 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1188 VDD.t105 a_31699_20742.t85 a_35502_25545.t6 VDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1189 VSS.t3122 VSS.t3121 VSS.t3122 VSS.t780 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1190 VSS.t3120 VSS.t3119 VSS.t3120 VSS.t847 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1191 a_52635_48695.t157 a_52635_34067.t96 VDD.t4952 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1192 VDD.t106 a_31699_20742.t86 a_33249_48695.t301 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1193 a_35502_25545.t27 a_35502_25545.t26 VSS.t165 VSS.t37 nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X1194 VDD.t4051 VDD.t4050 VDD.t4051 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1195 a_58851_n19597# a_50751_n19729.t113 VSS.t263 VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1196 VSS.t3118 VSS.t3117 VSS.t3118 VSS.t692 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1197 VDD.t4049 VDD.t4048 VDD.t4049 VDD.t2243 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1198 a_113037_n15000# a_71281_n8397.t129 a_112199_n14095# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1199 a_90245_n8770# a_71281_n10073.t117 a_89407_n8770# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1200 a_63161_n5344.t2 a_65658_4421.t1 a_66058_4481# VSS.t411 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1201 a_60845_n15112# a_50751_n19729.t114 a_60285_n14215# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1202 a_63683_n7138# a_50751_n19729.t115 a_63161_n7138# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1203 a_30152_n36322.t6 a_30152_n35156.t18 a_32088_n33224# VDD.t554 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1204 VDD.t4047 VDD.t4046 VDD.t4047 VDD.t1820 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1205 VSS.t3116 VSS.t3115 VSS.t3116 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1206 a_52635_49681.t26 a_35922_19591.t59 OUT.t81 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1207 VDD.t4045 VDD.t4044 VDD.t4045 VDD.t1221 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1208 a_36008_7563.t2 a_30152_11614.t9 a_37934_4481# VSS.t323 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1209 a_65677_n7138# a_50751_n19729.t116 a_65117_n7138# VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1210 a_44885_n12419# a_31953_n19727.t126 a_44363_n13316# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1211 a_77747_4481# a_77225_4481.t2 a_77225_4481.t3 VSS.t336 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1212 VDD.t4043 VDD.t4042 VDD.t4043 VDD.t552 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1213 a_60285_n15112# a_50751_n19729.t117 a_59763_n16906# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1214 a_36162_n36382.t7 a_41891_n29181.t14 a_43817_n27257# VSS.t181 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1215 a_100803_n4245# a_71281_n8397.t130 a_100235_n4245# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1216 VDD.t4041 VDD.t4040 VDD.t4041 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1217 VDD.t4039 VDD.t4038 VDD.t4039 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1218 a_52635_34067.t27 a_35922_19591.t60 a_52635_48695.t63 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1219 VDD.t4037 VDD.t4036 VDD.t4037 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1220 VSS.t3114 VSS.t3113 VSS.t3114 VSS.t676 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1221 VDD.t107 a_31699_20742.t87 a_33249_48695.t300 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1222 a_71281_n10073.t65 a_71281_n10073.t64 VDD.t362 VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1223 VDD.t4035 VDD.t4034 VDD.t4035 VDD.t2488 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1224 a_95943_n6055# a_71281_n10073.t118 a_78344_10448.t4 VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1225 VSS.t3112 VSS.t3111 VSS.t3112 VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1226 VDD.t4033 VDD.t4032 VDD.t4033 VDD.t1820 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1227 VDD.t4031 VDD.t4030 VDD.t4031 VDD.t1789 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1228 VDD.t4029 VDD.t4028 VDD.t4029 VDD.t1084 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1229 VDD.t4027 VDD.t4026 VDD.t4027 VDD.t63 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1230 a_84547_n18620# a_71281_n10073.t119 a_83709_n18620# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1231 VDD.t4025 VDD.t4024 VDD.t4025 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1232 VDD.t4023 VDD.t4022 VDD.t4023 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1233 a_40613_n2651# a_31953_n19727.t127 a_40053_n2651# VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1234 VSS.t3110 VSS.t3109 VSS.t3110 VSS.t314 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1235 VDD.t4021 VDD.t4020 VDD.t4021 VDD.t2488 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1236 a_54579_n15112# a_50751_n19729.t118 a_54019_n14215# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1237 VDD.t4019 VDD.t4018 VDD.t4019 VDD.t334 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1238 VSS.t3108 VSS.t3107 VSS.t3108 VSS.t446 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1239 VSS.t3106 VSS.t3105 VSS.t3106 VSS.t182 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1240 VDD.t4017 VDD.t4016 VDD.t4017 VDD.t1655 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1241 a_64243_n14215# a_50751_n19729.t119 a_63683_n14215# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1242 a_79151_n30339# a_77225_n29181.t12 VSS.t389 VSS.t387 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1243 VDD.t4015 VDD.t4014 VDD.t4015 VDD.t405 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1244 VSS.t196 a_35502_25545.t35 a_33249_34067.t137 VSS.t18 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1245 a_33249_48695.t299 a_31699_20742.t88 VDD.t108 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1246 a_32128_4481# a_30324_5507.t1 a_31284_4481.t1 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1247 a_52635_49681.t162 a_52635_34067.t97 VDD.t4951 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1248 a_32353_n8930# a_31953_n19727.t128 a_31831_n8930# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1249 VDD.t4013 VDD.t4012 VDD.t4013 VDD.t63 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1250 VDD.t4011 VDD.t4010 VDD.t4011 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1251 VDD.t4009 VDD.t4008 VDD.t4009 VDD.t1789 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1252 VSS.t3104 VSS.t3103 VSS.t3104 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1253 VDD.t4007 VDD.t4006 VDD.t4007 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1254 a_34347_n8930# a_31953_n19727.t129 a_33787_n8930# VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1255 VDD.t4005 VDD.t4004 VDD.t4005 VDD.t79 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1256 VDD.t4003 VDD.t4002 VDD.t4003 VDD.t2488 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1257 a_45706_24195# a_35922_19591.t61 a_45138_24195# VDD.t401 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X1258 a_33249_35053.t16 a_33379_34917.t18 a_33249_48695.t33 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1259 a_77747_n28415# a_77225_n29181.t13 a_71496_n36382.t0 VSS.t385 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1260 VDD.t4001 VDD.t4000 VDD.t4001 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1261 a_40053_n1754# a_31953_n19727.t130 VSS.t107 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1262 a_35502_24538.t20 a_31699_20742.t89 VDD.t109 VDD.t17 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1263 a_83725_n30339# a_32913_n8930.t1 a_83153_n36322.t2 VSS.t367 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1264 VDD.t3999 VDD.t3998 VDD.t3999 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1265 a_54229_10448# a_53829_10388.t10 a_36032_13546.t2 VDD.t3679 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1266 a_33249_34067.t86 a_33379_34007.t23 a_33249_48695.t114 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1267 VDD.t3997 VDD.t3996 VDD.t3997 VDD.t550 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1268 VDD.t43 a_31699_20742.t35 a_31699_20742.t36 VDD.t37 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1269 a_52635_49681.t161 a_52635_34067.t98 VDD.t4950 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1270 a_33249_34067.t14 a_35502_24538.t29 a_52635_34067.t3 VSS.t166 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1271 VDD.t3995 VDD.t3994 VDD.t3995 VDD.t390 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1272 a_46319_n13316# a_31953_n19727.t131 a_45797_n14213# VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1273 VSS.t3102 VSS.t3101 VSS.t3102 VSS.t1258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1274 VSS.t3100 VSS.t3099 VSS.t3100 VSS.t1432 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1275 VDD.t3993 VDD.t3992 VDD.t3993 VDD.t1052 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1276 a_33249_48695.t298 a_31699_20742.t90 VDD.t110 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1277 VDD.t3991 VDD.t3990 VDD.t3991 VDD.t50 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1278 VSS.t3098 VSS.t3097 VSS.t3098 VSS.t106 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1279 a_57977_n14215# a_50751_n19729.t120 a_57417_n14215# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1280 VSS.t3096 VSS.t3095 VSS.t3096 VSS.t864 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1281 VSS.t3094 VSS.t3093 VSS.t3094 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1282 VDD.t3989 VDD.t3988 VDD.t3989 VDD.t1183 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1283 VSS.t3092 VSS.t3091 VSS.t3092 VSS.t2042 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X1284 VDD.t111 a_31699_20742.t91 a_33249_48695.t297 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1285 a_52635_49681.t27 a_35922_19591.t62 OUT.t80 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1286 a_52635_34067.t27 a_35922_19591.t63 a_52635_48695.t62 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1287 a_41487_n1754# a_31953_n19727.t132 a_39179_n1754# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1288 VDD.t3987 VDD.t3986 VDD.t3987 VDD.t928 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1289 VDD.t3985 VDD.t3984 VDD.t3985 VDD.t559 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1290 VSS.t3090 VSS.t3089 VSS.t3090 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1291 VSS.t3088 VSS.t3087 VSS.t3088 VSS.t800 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1292 a_89715_n17715.t1 a_100992_4421.t1 a_113110_12380# VDD.t374 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1293 VSS.t3086 VSS.t3085 VSS.t3086 VSS.t223 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1294 VDD.t3983 VDD.t3982 VDD.t3983 VDD.t1422 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1295 a_57977_n6241# a_50751_n19729.t121 a_57417_n4447# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1296 VDD.t3981 VDD.t3980 VDD.t3981 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1297 VSS.t3084 VSS.t3083 VSS.t3084 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1298 VSS.t3082 VSS.t3081 VSS.t3082 VSS.t1621 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1299 a_71281_n10073.t63 a_71281_n10073.t62 VDD.t354 VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1300 VDD.t3979 VDD.t3978 VDD.t3979 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1301 a_51151_n3550# a_50751_n19729.t122 a_50629_n4447# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1302 VSS.t3080 VSS.t3079 VSS.t3080 VSS.t882 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1303 VDD.t3977 VDD.t3976 VDD.t3977 VDD.t1368 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1304 a_35502_25545.t7 a_31699_20742.t92 VDD.t112 VDD.t35 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1305 VSS.t3078 VSS.t3077 VSS.t3078 VSS.t596 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1306 VDD.t3975 VDD.t3974 VDD.t3975 VDD.t1158 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1307 VSS.t3076 VSS.t3075 VSS.t3076 VSS.t949 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1308 VDD.t458 a_71281_n8397.t56 a_71281_n8397.t57 VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1309 a_53145_n3550# a_50751_n19729.t123 a_52585_n3550# VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1310 VDD.t3973 VDD.t3972 VDD.t3973 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1311 a_52635_34067.t28 a_35922_19591.t64 a_52635_48695.t61 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1312 VDD.t3971 VDD.t3970 VDD.t3971 VDD.t123 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1313 VSS.t3074 VSS.t3073 VSS.t3074 VSS.t188 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1314 VSS.t3072 VSS.t3071 VSS.t3072 VSS.t596 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1315 VSS.t3070 VSS.t3069 VSS.t3070 VSS.t726 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1316 VDD.t3969 VDD.t3968 VDD.t3969 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1317 VSS.t3068 VSS.t3067 VSS.t3068 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1318 VDD.t3967 VDD.t3966 VDD.t3967 VDD.t913 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1319 a_110225_n9675# a_71281_n8397.t131 a_109695_n9675# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1320 a_52635_34067.t29 a_35922_19591.t65 a_52635_48695.t60 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1321 VDD.t3965 VDD.t3964 VDD.t3965 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1322 a_33249_48695.t117 a_33379_34007.t24 a_33249_34067.t85 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1323 VSS.t3066 VSS.t3065 VSS.t3066 VSS.t593 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1324 VDD.t3963 VDD.t3962 VDD.t3963 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1325 VSS.t3064 VSS.t3063 VSS.t3064 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1326 VSS.t3062 VSS.t3061 VSS.t3062 VSS.t0 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1327 VSS.t3060 VSS.t3059 VSS.t3060 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1328 a_37968_13546# a_36162_10388.t10 a_36008_4481.t2 VDD.t1713 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1329 a_47991_4421.t0 a_47819_11614.t12 a_54197_4481# VSS.t327 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1330 VDD.t4949 a_52635_34067.t99 a_52635_49681.t160 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1331 VSS.t3058 VSS.t3057 VSS.t3058 VSS.t1227 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1332 VSS.t3056 VSS.t3055 VSS.t3056 VSS.t1472 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1333 a_33249_34067.t84 a_33379_34007.t25 a_33249_48695.t118 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1334 a_33249_35053.t17 a_33379_34917.t19 a_33249_48695.t34 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1335 a_85129_n29181# a_32913_n8930.t2 a_31831_n5342.t0 VSS.t278 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1336 VDD.t3961 VDD.t3960 VDD.t3961 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1337 VDD.t3959 VDD.t3958 VDD.t3959 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1338 VDD.t3957 VDD.t3956 VDD.t3957 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1339 a_93969_n1530# a_71281_n10073.t120 a_93131_n1530# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1340 VSS.t3054 VSS.t3053 VSS.t3054 VSS.t500 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1341 a_99667_n13190# a_71281_n8397.t132 a_98829_n13190# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1342 a_33249_34067.t83 a_33379_34007.t26 a_33249_48695.t119 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1343 VDD.t3955 VDD.t3954 VDD.t3955 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1344 VDD.t3953 VDD.t3952 VDD.t3953 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1345 VSS.t358 a_89163_10388.t12 a_89563_12380# VDD.t558 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1346 VSS.t3052 VSS.t3051 VSS.t3052 VSS.t1391 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1347 a_114485_5639# a_112559_4481.t14 VSS.t291 VSS.t290 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1348 a_47753_n19595# a_31953_n19727.t133 VSS.t108 VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1349 VSS.t3050 VSS.t3049 VSS.t3050 VSS.t620 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1350 a_111063_n13190# a_71281_n8397.t133 a_110225_n13190# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1351 a_71896_10448# a_71496_10388.t14 a_53699_13546.t2 VDD.t488 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1352 VDD.t3951 VDD.t3950 VDD.t3951 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1353 VDD.t3949 VDD.t3948 VDD.t3949 VDD.t920 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1354 a_113037_n6055# a_71281_n8397.t134 VDD.t475 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1355 VSS.t3048 VSS.t3047 VSS.t3048 VSS.t765 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1356 VDD.t3947 VDD.t3946 VDD.t3947 VDD.t376 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1357 VDD.t3945 VDD.t3944 VDD.t3945 VDD.t1572 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1358 VDD.t3943 VDD.t3942 VDD.t3943 VDD.t968 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1359 a_37968_11614# a_36162_10388.t11 VSS.t438 VDD.t1713 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1360 VSS.t3046 VSS.t3045 VSS.t3046 VSS.t762 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1361 VSS.t3044 VSS.t3043 VSS.t3044 VSS.t686 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1362 a_82573_n2435# a_71281_n10073.t121 a_81735_n2435# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1363 VSS.t3042 VSS.t3041 VSS.t3042 VSS.t1600 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1364 a_54019_n12421# a_50751_n19729.t124 VSS.t264 VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1365 VDD.t3941 VDD.t3940 VDD.t3941 VDD.t1959 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1366 VSS.t3040 VSS.t3039 VSS.t3040 VSS.t689 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1367 a_52635_34067.t30 a_35922_19591.t66 a_52635_48695.t59 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1368 a_52635_48695.t58 a_35922_19591.t67 a_52635_34067.t31 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1369 VDD.t3939 VDD.t3938 VDD.t3939 VDD.t290 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1370 a_89531_n29181# a_83153_n36322.t10 VDD.t4786 VSS.t459 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1371 VDD.t3937 VDD.t3936 VDD.t3937 VDD.t1336 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1372 a_106501_n14095# a_71281_n8397.t135 a_105933_n14095# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1373 VDD.t3935 VDD.t3934 VDD.t3935 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1374 VSS.t86 a_31953_n19727.t56 a_31953_n19727.t57 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1375 a_99667_n2435# a_71281_n8397.t136 a_98829_n2435# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1376 VSS.t3038 VSS.t3037 VSS.t3038 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1377 VDD.t3933 VDD.t3932 VDD.t3933 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1378 a_33249_35053.t18 a_33379_34917.t20 a_33249_48695.t35 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1379 a_65117_n7138# a_50751_n19729.t125 a_64595_n8035# VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1380 VDD.t3931 VDD.t3930 VDD.t3931 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1381 VDD.t3929 VDD.t3928 VDD.t3929 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1382 a_101641_n6055# a_71281_n8397.t137 a_101111_n6055.t0 VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1383 VDD.t3927 VDD.t3926 VDD.t3927 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1384 VSS.t3036 VSS.t3035 VSS.t3036 VSS.t66 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1385 VSS.t3034 VSS.t3033 VSS.t3034 VSS.t676 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1386 VSS.t3032 VSS.t3031 VSS.t3032 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1387 VDD.t3925 VDD.t3924 VDD.t3925 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1388 a_52635_49681.t159 a_52635_34067.t100 VDD.t4948 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1389 VDD.t3923 VDD.t3922 VDD.t3923 VDD.t1938 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1390 a_38097_n16007.t1 a_47991_n29313.t0 a_48391_n29181# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1391 VSS.t3030 VSS.t3029 VSS.t3030 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1392 a_90245_n8770# a_71281_n10073.t122 a_89407_n7865# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1393 VDD.t3921 VDD.t3920 VDD.t3921 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1394 VDD.t3919 VDD.t3918 VDD.t3919 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1395 VDD.t3917 VDD.t3916 VDD.t3917 VDD.t1542 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1396 VDD.t3915 VDD.t3914 VDD.t3915 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1397 VDD.t113 a_31699_20742.t93 a_33249_48695.t296 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1398 VSS.t3028 VSS.t3027 VSS.t3028 VSS.t614 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1399 VDD.t3913 VDD.t3912 VDD.t3913 VDD.t1212 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1400 VDD.t4947 a_52635_34067.t101 a_52635_48695.t156 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1401 a_112559_n29181.t10 a_112559_n29181.t9 a_114485_n28415# VSS.t414 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1402 a_33379_34007.t27 IN_POS.t1 cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
X1403 VDD.t3911 VDD.t3910 VDD.t3911 VDD.t2779 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1404 VSS.t3026 VSS.t3025 VSS.t3026 VSS.t539 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1405 VDD.t3909 VDD.t3908 VDD.t3909 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1406 VDD.t3907 VDD.t3906 VDD.t3907 VDD.t494 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1407 a_67111_n8932# a_50751_n19729.t126 a_66551_n8035# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1408 a_67462_5639# a_65658_4421.t0 a_63161_n5344.t1 VSS.t412 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1409 VDD.t3905 VDD.t3904 VDD.t3905 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1410 a_63683_n15112# a_50751_n19729.t127 a_63161_n15112# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1411 VSS.t3024 VSS.t3023 VSS.t3024 VSS.t330 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1412 VSS.t3022 VSS.t3021 VSS.t3022 VSS.t1437 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1413 VDD.t3903 VDD.t3902 VDD.t3903 VDD.t2352 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1414 a_33249_35053.t19 a_33379_34917.t21 a_33249_48695.t36 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1415 a_33249_34067.t13 a_35502_24538.t30 a_52635_34067.t4 VSS.t167 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1416 VDD.t3901 VDD.t3900 VDD.t3901 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1417 VSS.t3020 VSS.t3019 VSS.t3020 VSS.t649 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1418 a_88839_n4245# a_71281_n10073.t123 a_88271_n4245# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1419 VDD.t4772 a_30152_n36322.t10 a_37934_n28415# VSS.t323 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1420 VDD.t3899 VDD.t3898 VDD.t3899 VDD.t2091 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1421 a_79182_10448# a_71366_11614.t4 a_78344_10448.t2 VDD.t575 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1422 VDD.t3897 VDD.t3896 VDD.t3897 VDD.t958 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1423 VDD.t3895 VDD.t3894 VDD.t3895 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1424 VDD.t3893 VDD.t3892 VDD.t3893 VDD.t1302 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1425 a_45445_n18698# a_31953_n19727.t134 a_44885_n18698# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1426 VDD.t3891 VDD.t3890 VDD.t3891 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1427 a_33249_35053.t20 a_33379_34917.t22 a_33249_48695.t37 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1428 VSS.t3018 VSS.t3017 VSS.t3018 VSS.t822 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1429 VSS.t3016 VSS.t3015 VSS.t3016 VSS.t896 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1430 a_35781_n15110# a_31953_n19727.t135 a_35221_n15110# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1431 a_94892_4481.t1 a_94892_4481.t0 a_96818_5639# VSS.t1349 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1432 a_84547_n17715# a_71281_n10073.t124 a_84017_n17715.t4 VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1433 VSS.t3014 VSS.t3013 VSS.t3014 VSS.t2481 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X1434 VSS.t3012 VSS.t3011 VSS.t3012 VSS.t643 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1435 VSS.t380 a_53829_n36382.t15 a_54229_n35156# VDD.t420 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1436 VDD.t3889 VDD.t3888 VDD.t3889 VDD.t3748 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1437 a_33249_48695.t295 a_31699_20742.t94 VDD.t114 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1438 VSS.t3010 VSS.t3009 VSS.t3010 VSS.t483 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1439 VSS.t3008 VSS.t3007 VSS.t3008 VSS.t738 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1440 OUT.t17 a_35502_24538.t31 a_33249_35053.t98 VSS.t163 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1441 a_66551_n18700# a_50751_n19729.t128 a_66029_n18700# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1442 VSS.t3006 VSS.t3005 VSS.t3006 VSS.t489 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1443 VSS.t3004 VSS.t3003 VSS.t3004 VSS.t1249 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1444 a_52635_34067.t30 a_35922_19591.t68 a_52635_48695.t57 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1445 VDD.t3887 VDD.t3886 VDD.t3887 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1446 a_46879_n14213# a_31953_n19727.t136 a_46319_n14213# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1447 VDD.t3885 VDD.t3884 VDD.t3885 VDD.t1938 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1448 a_89033_n36322.t1 a_106830_n36382.t9 a_108636_n36322# VDD.t1293 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1449 VDD.t3883 VDD.t3882 VDD.t3883 VDD.t968 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1450 VDD.t3881 VDD.t3880 VDD.t3881 VDD.t2352 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1451 VSS.t3002 VSS.t3001 VSS.t3002 VSS.t58 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1452 a_32353_n19595# a_31953_n19727.t137 a_31831_n19595# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1453 VDD.t42 a_31699_20742.t33 a_31699_20742.t34 VDD.t41 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1454 VDD.t4946 a_52635_34067.t102 a_52635_49681.t158 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1455 VDD.t3879 VDD.t3878 VDD.t3879 VDD.t1508 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1456 VDD.t3877 VDD.t3876 VDD.t3877 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1457 VSS.t3000 VSS.t2999 VSS.t3000 VSS.t1069 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1458 a_95414_n27257# a_94892_n29181.t4 a_94892_n29181.t5 VSS.t446 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1459 VDD.t3875 VDD.t3874 VDD.t3875 VDD.t923 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X1460 VSS.t2998 VSS.t2997 VSS.t2998 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1461 VDD.t3873 VDD.t3872 VDD.t3873 VDD.t1089 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1462 a_38619_n4445# a_31953_n19727.t138 a_38097_n4445# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1463 a_53675_n27257.t3 a_53829_n36382.t16 a_54229_n33224# VDD.t420 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1464 VSS.t2996 VSS.t2995 VSS.t2996 VSS.t281 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1465 a_33249_34067.t136 a_35502_25545.t36 VSS.t202 VSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1466 VDD.t3871 VDD.t3870 VDD.t3871 VDD.t965 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1467 VDD.t3869 VDD.t3868 VDD.t3869 VDD.t670 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1468 VDD.t421 a_100820_10448.t13 a_101350_12380# VDD.t301 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1469 VSS.t2994 VSS.t2993 VSS.t2994 VSS.t514 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1470 VDD.t457 a_71281_n8397.t54 a_71281_n8397.t55 VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1471 a_33249_34067.t135 a_35502_25545.t37 VSS.t193 VSS.t134 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1472 a_112559_4481.t8 a_112559_4481.t7 a_114485_7563# VSS.t286 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1473 a_50629_n16009.t0 a_51711_n12421.t0 a_83725_5639# VSS.t300 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1474 VSS.t176 a_41891_4481.t14 a_42413_7563# VSS.t171 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1475 VDD.t3867 VDD.t3866 VDD.t3867 VDD.t1492 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1476 VDD.t3865 VDD.t3864 VDD.t3865 VDD.t1167 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1477 VDD.t3863 VDD.t3862 VDD.t3863 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1478 VDD.t3861 VDD.t3860 VDD.t3861 VDD.t2061 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1479 VSS.t2992 VSS.t2991 VSS.t2992 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1480 a_52635_34067.t32 a_35922_19591.t69 a_52635_48695.t56 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1481 VSS.t2990 VSS.t2989 VSS.t2990 VSS.t1258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1482 VDD.t3859 VDD.t3858 VDD.t3859 VDD.t1489 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1483 a_31699_20742.t32 a_31699_20742.t31 VDD.t40 VDD.t35 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1484 a_71281_n8397.t0 I1N.t6 a_75585_n10973# VSS.t301 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X1485 a_33249_35053.t21 a_33379_34917.t23 a_33249_48695.t38 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1486 VDD.t3857 VDD.t3856 VDD.t3857 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1487 a_63683_n6241# a_50751_n19729.t129 a_63161_n7138# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1488 a_33249_48695.t294 a_31699_20742.t95 VDD.t115 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1489 VDD.t3855 VDD.t3854 VDD.t3855 VDD.t1268 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1490 a_52635_48695.t155 a_52635_34067.t103 VDD.t4945 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1491 VSS.t2988 VSS.t2987 VSS.t2988 VSS.t155 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1492 a_33249_48695.t293 a_31699_20742.t96 VDD.t116 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1493 VSS.t2986 VSS.t2985 VSS.t2986 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1494 VSS.t2984 VSS.t2983 VSS.t2984 VSS.t1311 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1495 a_96818_5639# a_94892_4481.t11 VSS.t3642 VSS.t1308 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1496 VSS.t2982 VSS.t2981 VSS.t2982 VSS.t581 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1497 a_33249_35053.t22 a_33379_34917.t24 a_33249_48695.t39 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1498 VDD.t3853 VDD.t3852 VDD.t3853 VDD.t1484 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1499 VDD.t3851 VDD.t3850 VDD.t3851 VDD.t2046 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1500 a_50751_n19729.t55 a_50751_n19729.t54 VSS.t240 VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1501 a_53675_n27257.t0 a_47819_n36322.t10 a_55601_n30339# VSS.t328 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1502 a_113110_13546# a_86903_n14095.t4 a_106830_10388.t0 VDD.t375 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1503 a_33249_34067.t134 a_35502_25545.t38 VSS.t180 VSS.t33 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1504 a_83141_n4245# a_71281_n10073.t125 a_82573_n4245# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1505 VSS.t2980 VSS.t2979 VSS.t2980 VSS.t695 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1506 a_52635_49681.t157 a_52635_34067.t104 VDD.t4944 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1507 VDD.t3849 VDD.t3848 VDD.t3849 VDD.t311 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1508 VDD.t3847 VDD.t3846 VDD.t3847 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1509 VDD.t3845 VDD.t3844 VDD.t3845 VDD.t792 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1510 VDD.t3843 VDD.t3842 VDD.t3843 VDD.t639 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1511 VSS.t2978 VSS.t2977 VSS.t2978 VSS.t1299 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1512 a_48349_13546# a_47819_10448.t12 a_47819_11614.t0 VDD.t497 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1513 VDD.t378 a_71281_n10073.t126 a_83709_n21335# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1514 VDD.t3841 VDD.t3840 VDD.t3841 VDD.t2023 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1515 a_100235_n4245# a_71281_n8397.t138 a_99667_n4245# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1516 VDD.t3839 VDD.t3838 VDD.t3839 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1517 a_56895_n16009.t0 a_57977_n12421.t0 a_101392_7563# VSS.t174 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1518 VSS.t2976 VSS.t2975 VSS.t2976 VSS.t681 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1519 VSS.t2974 VSS.t2973 VSS.t2974 VSS.t145 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1520 VSS.t2972 VSS.t2971 VSS.t2972 VSS.t1292 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1521 VSS.t2970 VSS.t2969 VSS.t2970 VSS.t495 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1522 a_39179_n19595.t0 a_47819_n36322.t11 a_54197_n28415# VSS.t327 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1523 VSS.t2968 VSS.t2967 VSS.t2968 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1524 a_59411_n7138# a_50751_n19729.t130 a_60285_n5344# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1525 VSS.t2966 VSS.t2965 VSS.t2966 VSS.t250 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1526 a_107339_n6960# a_71281_n8397.t139 a_106501_n6960# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1527 a_33249_35053.t23 a_33379_34917.t25 a_33249_48695.t40 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1528 VDD.t3837 VDD.t3836 VDD.t3837 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1529 VDD.t3835 VDD.t3834 VDD.t3835 VDD.t19 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1530 VSS.t2964 VSS.t2963 VSS.t2964 VSS.t768 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1531 a_65677_n13318# a_50751_n19729.t131 a_65117_n13318# VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1532 a_113110_11614# a_86903_n14095.t5 a_106830_10388.t1 VDD.t375 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1533 VDD.t3833 VDD.t3832 VDD.t3833 VDD.t1045 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1534 a_101641_n20430# a_71281_n8397.t140 a_100803_n19525# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1535 a_48313_n8930# a_31953_n19727.t139 a_47753_n8930# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1536 a_113081_7563# a_112559_4481.t15 a_106830_10388.t4 VSS.t285 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1537 a_51151_n18700# a_50751_n19729.t132 a_50629_n19597# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1538 a_51711_n8035# a_50751_n19729.t133 a_51151_n7138# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1539 VDD.t3831 VDD.t3830 VDD.t3831 VDD.t2682 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1540 VDD.t3829 VDD.t3828 VDD.t3829 VDD.t329 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1541 VDD.t3827 VDD.t3826 VDD.t3827 VDD.t614 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1542 a_65486_10448.t8 a_65658_4421.t0 a_67462_7563# VSS.t413 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1543 VDD.t3825 VDD.t3824 VDD.t3825 VDD.t2234 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1544 VSS.t2962 VSS.t2961 VSS.t2962 VSS.t596 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1545 VSS.t2960 VSS.t2959 VSS.t2960 VSS.t673 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1546 VDD.t3823 VDD.t3822 VDD.t3823 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1547 a_53829_n36382.t4 a_53699_n35156.t7 a_61515_n35156# VDD.t547 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1548 a_86903_n14095.t0 a_106830_10388.t12 a_108636_12380# VDD.t526 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1549 a_48349_11614# a_47819_10448.t13 a_47819_11614.t1 VDD.t497 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1550 VDD.t3821 VDD.t3820 VDD.t3821 VDD.t1613 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1551 a_67422_n34390# a_65486_n35156.t17 VDD.t7 VDD.t6 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1552 a_83725_5639# a_51711_n12421.t0 a_83153_11614.t3 VSS.t299 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1553 a_42413_7563# a_41891_4481.t15 a_36162_10388.t3 VSS.t177 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1554 a_51711_n16009.t1 a_50751_n19729.t134 a_51151_n16009# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1555 VSS.t2958 VSS.t2957 VSS.t2958 VSS.t593 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1556 VDD.t3819 VDD.t3818 VDD.t3819 VDD.t1998 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1557 VDD.t3817 VDD.t3816 VDD.t3817 VDD.t426 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1558 VSS.t2956 VSS.t2955 VSS.t2956 VSS.t312 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1559 a_52635_49681.t28 a_35922_19591.t70 OUT.t79 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1560 VDD.t117 a_31699_20742.t97 a_33249_48695.t292 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1561 a_79151_7563# a_77225_4481.t14 VSS.t339 VSS.t337 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1562 a_33249_34067.t133 a_35502_25545.t39 VSS.t19 VSS.t18 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1563 VSS.t41 a_35502_25545.t40 a_33249_35053.t138 VSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1564 a_60285_n4447# a_50751_n19729.t135 a_59763_n6241# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1565 a_33249_48695.t291 a_31699_20742.t98 VDD.t119 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1566 a_113037_n6960# a_71281_n8397.t141 a_112199_n4245# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1567 VSS.t2954 VSS.t2953 VSS.t2954 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1568 a_35221_n13316# a_31953_n19727.t140 a_34699_n14213# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1569 VDD.t4943 a_52635_34067.t105 a_52635_49681.t156 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1570 VDD.t3815 VDD.t3814 VDD.t3815 VDD.t908 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1571 VDD.t3813 VDD.t3812 VDD.t3813 VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1572 VDD.t3811 VDD.t3810 VDD.t3811 VDD.t2234 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1573 VDD.t3809 VDD.t3808 VDD.t3809 VDD.t63 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1574 VDD.t3807 VDD.t3806 VDD.t3807 VDD.t1221 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1575 VDD.t3805 VDD.t3804 VDD.t3805 VDD.t896 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1576 VDD.t3803 VDD.t3802 VDD.t3803 VDD.t389 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1577 a_53829_n36382.t5 a_53699_n35156.t8 a_61515_n33224# VDD.t547 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1578 VDD.t3801 VDD.t3800 VDD.t3801 VDD.t1613 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1579 VSS.t2952 VSS.t2951 VSS.t2952 VSS.t401 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1580 VDD.t3799 VDD.t3798 VDD.t3799 VDD.t313 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1581 VSS.t2950 VSS.t2949 VSS.t2950 VSS.t533 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1582 a_60677_n36322.t1 a_47991_n29313.t1 a_60109_n35156# VDD.t546 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1583 VSS.t2948 VSS.t2947 VSS.t2948 VSS.t458 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1584 VSS.t274 a_35502_25545.t41 a_33249_35053.t137 VSS.t15 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1585 a_107339_n20430# a_71281_n8397.t142 a_106501_n19525# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1586 a_110225_n13190# a_71281_n8397.t143 a_109695_n16810# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1587 a_33249_48695.t41 a_33379_34917.t26 a_33249_35053.t24 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1588 a_67111_n4447# a_50751_n19729.t136 a_66551_n3550# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1589 VSS.t2946 VSS.t2945 VSS.t2946 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1590 VDD.t3797 VDD.t3796 VDD.t3797 VDD.t1801 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1591 VSS.t2944 VSS.t2943 VSS.t2944 VSS.t873 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1592 VDD.t356 a_71281_n10073.t60 a_71281_n10073.t61 VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1593 VSS.t2942 VSS.t2941 VSS.t2942 VSS.t558 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1594 VDD.t3795 VDD.t3794 VDD.t3795 VDD.t1427 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1595 a_111063_n1530# a_71281_n8397.t144 a_110225_n1530# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1596 VSS.t2940 VSS.t2939 VSS.t2940 VSS.t555 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1597 VSS.t2938 VSS.t2937 VSS.t2938 VSS.t410 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1598 VSS.t2936 VSS.t2935 VSS.t2936 VSS.t819 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1599 VDD.t3793 VDD.t3792 VDD.t3793 VDD.t65 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1600 VDD.t4942 a_52635_34067.t106 a_52635_49681.t155 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1601 VDD.t3791 VDD.t3790 VDD.t3791 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1602 OUT.t16 a_35502_24538.t32 a_33249_35053.t99 VSS.t167 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1603 VDD.t3789 VDD.t3788 VDD.t3789 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1604 a_82573_n15000# a_71281_n10073.t127 a_81735_n15000# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1605 a_60677_n36322.t1 a_47991_n29313.t1 a_60109_n33224# VDD.t546 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1606 a_51151_n2653# a_50751_n19729.t137 a_50629_n2653# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1607 VSS.t2934 VSS.t2933 VSS.t2934 VSS.t284 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1608 VDD.t3787 VDD.t3786 VDD.t3787 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1609 VSS.t2932 VSS.t2931 VSS.t2932 VSS.t9 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1610 VSS.t2930 VSS.t2929 VSS.t2930 VSS.t163 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1611 VDD.t4941 a_52635_34067.t107 a_52635_48695.t154 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1612 a_33249_35053.t93 a_35502_24538.t33 OUT.t15 VSS.t166 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1613 VDD.t3785 VDD.t3784 VDD.t3785 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1614 a_52635_49681.t154 a_52635_34067.t108 VDD.t4940 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1615 VSS.t2928 VSS.t2927 VSS.t2928 VSS.t800 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1616 a_53145_n2653# a_50751_n19729.t138 a_52585_n2653# VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1617 a_52635_49681.t153 a_52635_34067.t109 VDD.t4939 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1618 VDD.t3783 VDD.t3782 VDD.t3783 VDD.t1411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1619 VSS.t2926 VSS.t2925 VSS.t2926 VSS.t623 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1620 VDD.t3781 VDD.t3780 VDD.t3781 VDD.t928 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1621 VSS.t2924 VSS.t2923 VSS.t2924 VSS.t1600 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1622 a_52635_49681.t152 a_52635_34067.t110 VDD.t4938 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1623 VSS.t317 a_59558_n29181.t14 a_60080_n29181# VSS.t316 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1624 VDD.t3779 VDD.t3778 VDD.t3779 VDD.t855 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1625 VSS.t2922 VSS.t2921 VSS.t2922 VSS.t539 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1626 VDD.t4782 a_65486_11614.t9 a_73268_5639# VSS.t427 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1627 VSS.t2920 VSS.t2919 VSS.t2920 VSS.t738 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1628 VDD.t3777 VDD.t3776 VDD.t3777 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1629 VSS.t2918 VSS.t2917 VSS.t2918 VSS.t620 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1630 VDD.t3775 VDD.t3774 VDD.t3775 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1631 VDD.t3773 VDD.t3772 VDD.t3773 VDD.t551 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1632 VSS.t2916 VSS.t2915 VSS.t2916 VSS.t655 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1633 VDD.t3771 VDD.t3770 VDD.t3771 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1634 a_32913_n12419# a_31953_n19727.t141 a_32353_n12419# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1635 VDD.t3769 VDD.t3768 VDD.t3769 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1636 a_46274_23609# a_35922_19591.t71 a_45706_23609# VDD.t406 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X1637 VSS.t2914 VSS.t2913 VSS.t2914 VSS.t1320 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1638 VDD.t3767 VDD.t3766 VDD.t3767 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1639 VSS.t2912 VSS.t2911 VSS.t2912 VSS.t1621 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1640 VSS.t198 a_35502_25545.t42 a_33249_34067.t132 VSS.t26 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1641 VSS.t190 a_35502_24538.t34 a_41100_19075# VSS.t189 nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X1642 VSS.t2910 VSS.t2909 VSS.t2910 VSS.t609 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1643 VSS.t2908 VSS.t2907 VSS.t2908 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1644 VDD.t3765 VDD.t3764 VDD.t3765 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1645 a_33249_48695.t290 a_31699_20742.t99 VDD.t120 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1646 VDD.t3763 VDD.t3762 VDD.t3763 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1647 VDD.t3761 VDD.t3760 VDD.t3761 VDD.t700 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1648 VDD.t3759 VDD.t3758 VDD.t3759 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1649 VDD.t3757 VDD.t3756 VDD.t3757 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1650 VSS.t2906 VSS.t2905 VSS.t2906 VSS.t1543 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1651 VSS.t2904 VSS.t2903 VSS.t2904 VSS.t483 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1652 VDD.t3755 VDD.t3754 VDD.t3755 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1653 VDD.t3753 VDD.t3752 VDD.t3753 VDD.t913 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1654 VDD.t3751 VDD.t3750 VDD.t3751 VDD.t3571 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1655 VDD.t3749 VDD.t3747 VDD.t3749 VDD.t3748 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1656 a_33249_48695.t289 a_31699_20742.t100 VDD.t121 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1657 a_67111_n17803# a_50751_n19729.t139 a_66551_n17803# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1658 a_52635_49681.t151 a_52635_34067.t111 VDD.t4937 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1659 a_105365_n9675# a_71281_n8397.t145 a_104527_n9675# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1660 a_63683_n1756# a_50751_n19729.t140 a_63161_n2653# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1661 VSS.t2902 VSS.t2901 VSS.t2902 VSS.t777 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1662 VDD.t122 a_31699_20742.t101 a_33249_48695.t288 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1663 VDD.t3746 VDD.t3745 VDD.t3746 VDD.t982 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1664 a_105933_n4245# a_71281_n8397.t146 a_105365_n4245# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1665 VSS.t239 a_50751_n19729.t52 a_50751_n19729.t53 VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1666 a_82573_n20430# a_71281_n10073.t128 a_81735_n20430# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1667 a_53675_4481.t1 a_47819_11614.t13 a_55601_7563# VSS.t328 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1668 VDD.t3744 VDD.t3743 VDD.t3744 VDD.t700 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1669 VDD.t3742 VDD.t3741 VDD.t3742 VDD.t1158 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1670 VDD.t3740 VDD.t3739 VDD.t3740 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1671 a_65677_n2653# a_50751_n19729.t141 a_65117_n1756# VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1672 VSS.t2900 VSS.t2899 VSS.t2900 VSS.t709 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1673 VSS.t2898 VSS.t2897 VSS.t2898 VSS.t1039 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1674 a_71864_5639# a_65486_11614.t10 VDD.t4783 VSS.t428 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1675 VDD.t3738 VDD.t3737 VDD.t3738 VDD.t804 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1676 a_43817_n30339# a_41891_n29181.t15 VSS.t374 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1677 a_42442_13546# a_36032_11614.t7 a_36162_10388.t5 VDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1678 VDD.t3736 VDD.t3735 VDD.t3736 VDD.t1517 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1679 VDD.t3734 VDD.t3733 VDD.t3734 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1680 VSS.t2896 VSS.t2895 VSS.t2896 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1681 VDD.t3732 VDD.t3731 VDD.t3732 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1682 a_53829_10388.t6 a_53699_11614.t3 a_61515_12380# VDD.t493 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1683 VDD.t3730 VDD.t3729 VDD.t3730 VDD.t2122 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1684 VDD.t3728 VDD.t3727 VDD.t3728 VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1685 a_38619_n17801# a_31953_n19727.t142 a_38097_n17801# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1686 VSS.t2894 VSS.t2893 VSS.t2894 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1687 a_100235_n18620# a_71281_n8397.t147 a_99667_n18620# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1688 VSS.t2892 VSS.t2891 VSS.t2892 VSS.t573 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1689 VDD.t3726 VDD.t3725 VDD.t3726 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1690 VSS.t2890 VSS.t2889 VSS.t2890 VSS.t913 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1691 a_49795_n30339# a_47991_n29313.t0 a_38097_n16007.t2 VSS.t281 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1692 VDD.t3724 VDD.t3723 VDD.t3724 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1693 VSS.t2888 VSS.t2887 VSS.t2888 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1694 VSS.t2886 VSS.t2885 VSS.t2886 VSS.t411 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1695 a_31953_n19727.t55 a_31953_n19727.t54 VSS.t85 VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1696 a_52635_48695.t55 a_35922_19591.t72 a_52635_34067.t33 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1697 a_52635_34067.t61 a_35502_24538.t35 a_33249_34067.t12 VSS.t182 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1698 VDD.t3722 VDD.t3721 VDD.t3722 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1699 a_33249_34067.t82 a_33379_34007.t28 a_33249_48695.t106 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1700 a_96818_n28415# a_94892_n29181.t12 VSS.t448 VSS.t447 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1701 a_111631_n13190# a_71281_n8397.t148 a_111063_n13190# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1702 a_65658_n29313.t0 a_65486_n36322.t12 a_71864_n27257# VSS.t155 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1703 a_33249_48695.t287 a_31699_20742.t102 VDD.t124 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1704 a_42442_11614# a_36032_11614.t8 a_36162_10388.t6 VDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1705 VDD.t3720 VDD.t3719 VDD.t3720 VDD.t1517 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1706 VSS.t2884 VSS.t2883 VSS.t2884 VSS.t1162 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1707 VDD.t3718 VDD.t3717 VDD.t3718 VDD.t2122 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1708 VDD.t3716 VDD.t3715 VDD.t3716 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1709 VDD.t3714 VDD.t3713 VDD.t3714 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1710 a_36032_11614.t0 a_36162_10388.t12 a_37968_12380# VDD.t1497 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1711 VDD.t3712 VDD.t3711 VDD.t3712 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1712 a_33249_48695.t286 a_31699_20742.t103 VDD.t126 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1713 a_102756_n35156# a_100820_n35156.t15 VDD.t533 VDD.t530 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1714 VSS.t2882 VSS.t2881 VSS.t2882 VSS.t573 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1715 VSS.t2880 VSS.t2879 VSS.t2880 VSS.t415 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1716 a_36162_10388.t2 a_41891_4481.t16 a_43817_4481# VSS.t181 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1717 a_35781_n15110# a_31953_n19727.t143 a_35221_n14213# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1718 VDD.t3710 VDD.t3709 VDD.t3710 VDD.t2575 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1719 a_36008_4481.t3 a_36162_10388.t13 a_36562_10448# VDD.t3614 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1720 VDD.t3708 VDD.t3707 VDD.t3708 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1721 VDD.t3706 VDD.t3705 VDD.t3706 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1722 VSS.t2878 VSS.t2877 VSS.t2878 VSS.t106 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1723 a_98829_n18620# a_71281_n8397.t149 a_98299_n19525# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1724 a_30152_11614.t3 a_30324_5507.t1 a_32128_6405# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1725 VDD.t3704 VDD.t3703 VDD.t3704 VDD.t2572 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1726 VDD.t3702 VDD.t3701 VDD.t3702 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1727 VDD.t3700 VDD.t3699 VDD.t3700 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1728 VSS.t2876 VSS.t2875 VSS.t2876 VSS.t469 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1729 VSS.t2874 VSS.t2873 VSS.t2874 VSS.t329 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1730 a_33249_34067.t131 a_35502_25545.t43 VSS.t205 VSS.t142 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1731 a_33787_n18698# a_31953_n19727.t144 a_33265_n18698# VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1732 a_30724_n27257# a_30324_n29313.t1 a_30152_n35156.t11 VSS.t145 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1733 VSS.t2872 VSS.t2871 VSS.t2872 VSS.t550 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1734 VDD.t3698 VDD.t3697 VDD.t3698 VDD.t490 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1735 VDD.t3696 VDD.t3695 VDD.t3696 VDD.t1869 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1736 VSS.t2870 VSS.t2869 VSS.t2870 VSS.t655 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1737 VDD.t3694 VDD.t3693 VDD.t3694 VDD.t375 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1738 a_105365_n18620# a_71281_n8397.t150 a_104527_n18620# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1739 a_55601_7563# a_47819_11614.t14 a_47991_4421.t0 VSS.t330 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1740 VSS.t2868 VSS.t2867 VSS.t2868 VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1741 a_102756_n33224# a_100820_n35156.t16 VDD.t534 VDD.t530 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1742 VSS.t2866 VSS.t2865 VSS.t2866 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1743 VSS.t2864 VSS.t2863 VSS.t2864 VSS.t58 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1744 VDD.t3692 VDD.t3691 VDD.t3692 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1745 VDD.t3690 VDD.t3689 VDD.t3690 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1746 a_33249_35053.t136 a_35502_25545.t44 VSS.t195 VSS.t24 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1747 VDD.t3688 VDD.t3687 VDD.t3688 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1748 a_33249_48695.t285 a_31699_20742.t104 VDD.t127 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1749 VSS.t2862 VSS.t2861 VSS.t2862 VSS.t646 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1750 VDD.t3686 VDD.t3685 VDD.t3686 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1751 a_52635_48695.t54 a_35922_19591.t73 a_52635_34067.t34 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1752 VDD.t3684 VDD.t3683 VDD.t3684 VDD.t402 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1753 VDD.t3682 VDD.t3681 VDD.t3682 VDD.t529 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1754 VSS.t2860 VSS.t2859 VSS.t2860 VSS.t1261 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1755 VDD.t39 a_31699_20742.t29 a_31699_20742.t30 VDD.t17 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1756 VSS.t2858 VSS.t2857 VSS.t2858 VSS.t385 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1757 VDD.t3680 VDD.t3678 VDD.t3680 VDD.t3679 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1758 VDD.t3677 VDD.t3676 VDD.t3677 VDD.t2923 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1759 a_110225_n3340# a_71281_n8397.t151 a_109695_n4245# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1760 a_100820_11614.t6 a_57977_n12421.t0 a_102796_4481# VSS.t173 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1761 a_33249_48695.t107 a_33379_34007.t29 a_33249_34067.t81 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1762 a_31284_4481.t1 a_30324_4421.t2 a_30724_4481# VSS.t146 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1763 VDD.t372 a_71281_n10073.t58 a_71281_n10073.t59 VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1764 a_58851_n8035# a_50751_n19729.t142 a_58329_n8035# VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1765 a_52635_49681.t150 a_52635_34067.t112 VDD.t4936 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1766 VSS.t2856 VSS.t2855 VSS.t2856 VSS.t282 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1767 VSS.t2854 VSS.t2853 VSS.t2854 VSS.t390 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1768 VDD.t128 a_31699_20742.t105 a_33249_48695.t284 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1769 a_52635_49681.t149 a_52635_34067.t113 VDD.t4935 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1770 VDD.t3675 VDD.t3674 VDD.t3675 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1771 VDD.t3673 VDD.t3672 VDD.t3673 VDD.t554 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1772 VDD.t3671 VDD.t3670 VDD.t3671 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1773 VDD.t3669 VDD.t3668 VDD.t3669 VDD.t318 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1774 VDD.t3667 VDD.t3666 VDD.t3667 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1775 a_57417_n16906# a_50751_n19729.t143 a_56895_n17803# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1776 VSS.t2852 VSS.t2851 VSS.t2852 VSS.t11 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1777 VSS.t2850 VSS.t2849 VSS.t2850 VSS.t166 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1778 VDD.t3665 VDD.t3664 VDD.t3665 VDD.t402 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1779 VDD.t3663 VDD.t3662 VDD.t3663 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1780 a_102796_6405# a_57977_n12421.t2 a_56895_n16009.t0 VSS.t144 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1781 VDD.t3661 VDD.t3660 VDD.t3661 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1782 VDD.t3659 VDD.t3658 VDD.t3659 VDD.t315 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1783 VDD.t129 a_31699_20742.t106 a_33249_48695.t283 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1784 VDD.t3657 VDD.t3656 VDD.t3657 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1785 a_82573_n15905# a_71281_n10073.t129 a_81735_n15905# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1786 a_43817_4481# a_41891_4481.t17 VSS.t161 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1787 a_33249_35053.t25 a_33379_34917.t27 a_33249_48695.t42 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1788 VSS.t2848 VSS.t2847 VSS.t2848 VSS.t981 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1789 a_66058_n30339# a_45445_n19595.t1 a_65486_n36322.t4 VSS.t410 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1790 a_48313_n15110# a_31953_n19727.t145 a_47753_n15110# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1791 a_112199_n6960# a_71281_n8397.t152 a_111631_n6960# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1792 a_83325_n29313.t0 a_83153_n36322.t11 a_89531_n27257# VSS.t458 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1793 VDD.t3655 VDD.t3654 VDD.t3655 VDD.t557 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1794 VDD.t3653 VDD.t3652 VDD.t3653 VDD.t123 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1795 VSS.t238 a_50751_n19729.t50 a_50751_n19729.t51 VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1796 a_89563_n34390# a_89163_n36382.t10 a_89033_n35156.t1 VDD.t549 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1797 a_52635_49681.t29 a_35922_19591.t74 OUT.t78 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1798 VDD.t3651 VDD.t3650 VDD.t3651 VDD.t1820 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1799 VDD.t3649 VDD.t3648 VDD.t3649 VDD.t527 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1800 VSS.t2846 VSS.t2845 VSS.t2846 VSS.t506 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1801 VDD.t3647 VDD.t3646 VDD.t3647 VDD.t52 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1802 VSS.t2844 VSS.t2843 VSS.t2844 VSS.t952 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1803 VSS.t2842 VSS.t2841 VSS.t2842 VSS.t1621 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1804 VDD.t3645 VDD.t3644 VDD.t3645 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1805 VDD.t3643 VDD.t3642 VDD.t3643 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1806 VDD.t130 a_31699_20742.t107 a_33249_48695.t282 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1807 VSS.t2840 VSS.t2839 VSS.t2840 VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1808 VSS.t2838 VSS.t2837 VSS.t2838 VSS.t49 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1809 VDD.t3641 VDD.t3640 VDD.t3641 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1810 VSS.t2836 VSS.t2835 VSS.t2836 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1811 VDD.t3639 VDD.t3638 VDD.t3639 VDD.t1089 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1812 a_41100_19075# a_35502_24538.t36 a_40578_19075# VSS.t184 nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X1813 VDD.t3637 VDD.t3636 VDD.t3637 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1814 VSS.t2834 VSS.t2833 VSS.t2834 VSS.t495 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1815 a_35502_24538.t19 a_31699_20742.t108 VDD.t131 VDD.t21 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1816 a_48391_n27257# a_47991_n29313.t2 a_47819_n35156.t8 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1817 a_101392_4481# a_100992_4421.t2 a_100820_10448.t3 VSS.t175 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1818 VDD.t3635 VDD.t3634 VDD.t3635 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1819 a_65677_n13318# a_50751_n19729.t144 a_65117_n12421# VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1820 VSS.t2832 VSS.t2831 VSS.t2832 VSS.t1472 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1821 VDD.t3633 VDD.t3632 VDD.t3633 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1822 a_51711_n6241# a_50751_n19729.t145 a_51151_n6241# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1823 a_89715_n5150.t1 a_71281_n10073.t130 a_89407_n1530# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1824 VSS.t2830 VSS.t2829 VSS.t2830 VSS.t1131 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1825 VSS.t2828 VSS.t2827 VSS.t2828 VSS.t284 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1826 a_65486_n36322.t6 a_45445_n19595.t1 a_67462_n29181# VSS.t413 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1827 VSS.t2826 VSS.t2825 VSS.t2826 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1828 a_30724_4481# a_30324_4421.t2 a_30152_10448.t0 VSS.t145 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1829 VDD.t3631 VDD.t3630 VDD.t3631 VDD.t1789 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1830 VDD.t3629 VDD.t3628 VDD.t3629 VDD.t502 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1831 a_51711_n16906# a_50751_n19729.t146 a_51151_n15112# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1832 a_107198_5639# a_100820_11614.t8 VDD.t294 VSS.t150 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1833 VSS.t2824 VSS.t2823 VSS.t2824 VSS.t655 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1834 a_33249_48695.t43 a_33379_34917.t28 a_33249_35053.t26 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1835 VDD.t3627 VDD.t3626 VDD.t3627 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1836 VSS.t2822 VSS.t2821 VSS.t2822 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1837 a_65117_n1756# a_50751_n19729.t147 a_64243_n5344.t0 VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1838 VSS.t2820 VSS.t2819 VSS.t2820 VSS.t1116 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1839 a_33249_34067.t80 a_33379_34007.t30 a_33249_48695.t108 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1840 VSS.t2818 VSS.t2817 VSS.t2818 VSS.t253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1841 VSS.t2816 VSS.t2815 VSS.t2816 VSS.t98 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1842 VDD.t4934 a_52635_34067.t114 a_52635_49681.t148 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1843 VSS.t2814 VSS.t2813 VSS.t2814 VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1844 VDD.t3625 VDD.t3624 VDD.t3625 VDD.t1183 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1845 a_33249_35053.t27 a_33379_34917.t29 a_33249_48695.t44 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1846 VSS.t2812 VSS.t2811 VSS.t2812 VSS.t1543 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1847 a_52635_48695.t153 a_52635_34067.t115 VDD.t4933 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1848 VDD.t3623 VDD.t3622 VDD.t3623 VDD.t81 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1849 a_90969_13546# a_89163_10388.t13 a_89009_4481.t2 VDD.t559 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1850 a_33249_48695.t281 a_31699_20742.t109 VDD.t132 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1851 VSS.t2810 VSS.t2809 VSS.t2810 VSS.t464 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1852 VDD.t3621 VDD.t3620 VDD.t3621 VDD.t2488 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1853 VSS.t237 a_50751_n19729.t48 a_50751_n19729.t49 VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1854 VSS.t442 a_106830_n36382.t10 a_107230_n34390# VDD.t848 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1855 VSS.t2808 VSS.t2807 VSS.t2808 VSS.t503 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1856 a_89407_n8770# a_71281_n10073.t131 a_88839_n8770# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1857 VSS.t2806 VSS.t2805 VSS.t2806 VSS.t942 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1858 a_67111_n2653# a_50751_n19729.t148 a_66551_n2653# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1859 VDD.t3619 VDD.t3618 VDD.t3619 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1860 VDD.t3617 VDD.t3616 VDD.t3617 VDD.t839 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1861 VDD.t3615 VDD.t3613 VDD.t3615 VDD.t3614 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1862 VDD.t3612 VDD.t3611 VDD.t3612 VDD.t1254 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1863 a_32353_n8033# a_31953_n19727.t146 a_31831_n8930# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1864 a_53145_n7138# a_50751_n19729.t149 a_54019_n5344# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1865 a_40053_n8930# a_31953_n19727.t147 a_39179_n5342.t0 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1866 VDD.t3610 VDD.t3609 VDD.t3610 VDD.t1183 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1867 a_71281_n8397.t53 a_71281_n8397.t52 VDD.t456 VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1868 a_54019_n18700# a_50751_n19729.t150 a_53497_n18700# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1869 a_40053_n12419# a_31953_n19727.t148 VSS.t109 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1870 VSS.t2804 VSS.t2803 VSS.t2804 VSS.t652 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1871 VDD.t3608 VDD.t3607 VDD.t3608 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1872 a_90969_11614# a_89163_10388.t14 VSS.t359 VDD.t559 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1873 VDD.t3606 VDD.t3605 VDD.t3606 VDD.t1045 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1874 VDD.t3604 VDD.t3603 VDD.t3604 VDD.t2302 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X1875 a_34347_n8930# a_31953_n19727.t149 a_33787_n8033# VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1876 VSS.t2802 VSS.t2801 VSS.t2802 VSS.t414 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1877 VSS.t2800 VSS.t2799 VSS.t2800 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1878 VSS.t2798 VSS.t2797 VSS.t2798 VSS.t353 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1879 VDD.t513 a_47819_10448.t14 a_48349_12380# VDD.t512 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1880 VSS.t2796 VSS.t2795 VSS.t2796 VSS.t362 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1881 VDD.t3602 VDD.t3601 VDD.t3602 VDD.t826 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1882 VSS.t2794 VSS.t2793 VSS.t2794 VSS.t259 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1883 VSS.t2792 VSS.t2791 VSS.t2792 VSS.t536 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1884 VDD.t3600 VDD.t3599 VDD.t3600 VDD.t426 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1885 a_67422_n36322# a_65486_n35156.t18 VDD.t8 VDD.t6 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1886 VDD.t3598 VDD.t3597 VDD.t3598 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1887 a_41487_n8930# a_31953_n19727.t150 VSS.t110 VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1888 a_33249_48695.t280 a_31699_20742.t110 VDD.t133 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1889 VSS.t2790 VSS.t2789 VSS.t2790 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1890 VSS.t2788 VSS.t2787 VSS.t2788 VSS.t1437 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1891 VSS.t2786 VSS.t2785 VSS.t2786 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1892 VDD.t3596 VDD.t3595 VDD.t3596 VDD.t813 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1893 VSS.t2784 VSS.t2783 VSS.t2784 VSS.t323 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1894 VSS.t2782 VSS.t2781 VSS.t2782 VSS.t576 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1895 VDD.t3594 VDD.t3593 VDD.t3594 VDD.t3355 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1896 a_33249_48695.t45 a_33379_34917.t30 a_33249_35053.t28 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1897 VDD.t4932 a_52635_34067.t116 a_52635_49681.t147 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1898 VSS.t2780 VSS.t2779 VSS.t2780 VSS.t638 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1899 VDD.t4931 a_52635_34067.t117 a_52635_48695.t152 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1900 a_61484_n30339# a_59558_n29181.t15 VSS.t318 VSS.t314 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1901 a_83325_4421.t0 a_83153_11614.t15 a_89531_4481# VSS.t399 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1902 VSS.t2778 VSS.t2777 VSS.t2778 VSS.t873 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1903 a_98829_n17715# a_71281_n8397.t153 a_98299_n21335# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1904 VSS.t2776 VSS.t2775 VSS.t2776 VSS.t847 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1905 a_100820_n35156.t2 a_100992_n29313.t0 a_102796_n30339# VSS.t382 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1906 VSS.t2774 VSS.t2773 VSS.t2774 VSS.t738 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1907 VSS.t2772 VSS.t2771 VSS.t2772 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1908 VDD.t3592 VDD.t3591 VDD.t3592 VDD.t376 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1909 a_85129_6405# a_51711_n12421.t2 a_50629_n16009.t0 VSS.t298 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1910 VDD.t3590 VDD.t3589 VDD.t3590 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1911 VDD.t3588 VDD.t3587 VDD.t3588 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1912 VDD.t3586 VDD.t3585 VDD.t3586 VDD.t920 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1913 a_52635_49681.t30 a_35922_19591.t75 OUT.t77 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1914 VSS.t2770 VSS.t2769 VSS.t2770 VSS.t324 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1915 VSS.t2768 VSS.t2767 VSS.t2768 VSS.t1162 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1916 VDD.t134 a_31699_20742.t111 a_35502_25545.t8 VDD.t41 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1917 VDD.t3584 VDD.t3583 VDD.t3584 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1918 VSS.t2766 VSS.t2765 VSS.t2766 VSS.t563 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1919 VDD.t455 a_71281_n8397.t50 a_71281_n8397.t51 VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1920 VDD.t3582 VDD.t3581 VDD.t3582 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1921 a_58851_n3550# a_50751_n19729.t151 a_58329_n3550# VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1922 VSS.t2764 VSS.t2763 VSS.t2764 VSS.t492 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1923 VDD.t3580 VDD.t3579 VDD.t3580 VDD.t1959 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1924 a_95443_n34390# a_89033_n35156.t9 a_89163_n36382.t0 VDD.t798 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1925 VDD.t3578 VDD.t3577 VDD.t3578 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1926 a_95443_12380# a_83325_4421.t1 a_94892_4481.t8 VDD.t500 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1927 VSS.t2762 VSS.t2761 VSS.t2762 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1928 VSS.t2760 VSS.t2759 VSS.t2760 VSS.t542 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1929 a_44885_n7136# a_31953_n19727.t151 a_44363_n7136# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1930 VSS.t2758 VSS.t2757 VSS.t2758 VSS.t704 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1931 VSS.t2756 VSS.t2755 VSS.t2756 VSS.t35 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1932 a_34347_n17801# a_31953_n19727.t152 a_33787_n17801# VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1933 VDD.t363 a_71281_n10073.t56 a_71281_n10073.t57 VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1934 VDD.t3576 VDD.t3575 VDD.t3576 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1935 VDD.t3574 VDD.t3573 VDD.t3574 VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1936 a_52635_49681.t31 a_35922_19591.t76 OUT.t76 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1937 a_52635_49681.t32 a_35922_19591.t77 OUT.t75 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1938 a_90245_n17715# a_71281_n10073.t132 a_89715_n16810.t0 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1939 a_46879_n7136# a_31953_n19727.t153 a_46319_n7136# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1940 VDD.t3572 VDD.t3570 VDD.t3572 VDD.t3571 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1941 VSS.t2754 VSS.t2753 VSS.t2754 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1942 VDD.t3569 VDD.t3568 VDD.t3569 VDD.t1843 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1943 VDD.t300 a_65486_n36322.t13 a_73268_n28415# VSS.t154 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1944 VDD.t3567 VDD.t3566 VDD.t3567 VDD.t920 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1945 a_95105_n15000# a_71281_n10073.t133 a_94537_n15000# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1946 a_47753_n16007# a_31953_n19727.t154 a_46879_n17801# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1947 a_110225_n2435# a_71281_n8397.t154 VDD.t476 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1948 a_88271_n4245# a_71281_n10073.t134 a_87433_n4245# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1949 VSS.t2752 VSS.t2751 VSS.t2752 VSS.t617 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1950 a_90245_n15000# a_71281_n10073.t135 a_89407_n15000# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1951 VDD.t3565 VDD.t3564 VDD.t3565 VDD.t1938 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1952 VDD.t3563 VDD.t3562 VDD.t3563 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1953 VDD.t3561 VDD.t3560 VDD.t3561 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1954 a_37968_10448# a_36162_10388.t14 a_36008_7563.t0 VDD.t1713 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1955 VDD.t3559 VDD.t3558 VDD.t3559 VDD.t1198 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1956 VDD.t3557 VDD.t3556 VDD.t3557 VDD.t1959 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1957 VSS.t2750 VSS.t2749 VSS.t2750 VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1958 a_77747_n27257# a_77225_n29181.t2 a_77225_n29181.t3 VSS.t385 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1959 a_100235_n21335# a_71281_n8397.t155 a_99667_n21335# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1960 VSS.t2748 VSS.t2747 VSS.t2748 VSS.t842 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1961 VDD.t3555 VDD.t3554 VDD.t3555 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1962 VDD.t3553 VDD.t3552 VDD.t3553 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1963 VSS.t2746 VSS.t2745 VSS.t2746 VSS.t324 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1964 a_42047_n7136# a_31953_n19727.t155 a_41487_n6239# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1965 VDD.t4751 a_65486_10448.t14 a_66016_12380# VDD.t1341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1966 VSS.t2744 VSS.t2743 VSS.t2744 VSS.t52 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1967 VSS.t2742 VSS.t2741 VSS.t2742 VSS.t563 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1968 VDD.t135 a_31699_20742.t112 a_33249_48695.t279 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1969 VDD.t3551 VDD.t3550 VDD.t3551 VDD.t3424 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1970 VDD.t3549 VDD.t3548 VDD.t3549 VDD.t1336 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1971 a_112559_n29181.t2 a_100992_n29313.t2 a_114516_n34390# VDD.t331 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1972 a_60677_10448.t5 a_53699_11614.t4 a_60109_13546# VDD.t494 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1973 a_32128_n28415# a_30324_n29313.t0 a_31284_n30339.t0 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1974 VSS.t2740 VSS.t2739 VSS.t2740 VSS.t44 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1975 VSS.t2738 VSS.t2737 VSS.t2738 VSS.t187 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1976 a_107198_n30339# a_100820_n36322.t11 a_106676_n30339.t0 VSS.t352 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1977 a_52635_49681.t146 a_52635_34067.t118 VDD.t4930 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1978 VSS.t2736 VSS.t2735 VSS.t2736 VSS.t527 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1979 a_89531_4481# a_83153_11614.t16 a_89009_4481.t0 VSS.t400 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1980 a_71281_n10073.t55 a_71281_n10073.t54 VDD.t336 VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1981 VDD.t3547 VDD.t3546 VDD.t3547 VDD.t1938 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1982 VDD.t3545 VDD.t3544 VDD.t3545 VDD.t394 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1983 VDD.t3543 VDD.t3542 VDD.t3543 VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1984 a_88839_n15000# a_71281_n10073.t136 a_88271_n15000# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1985 VDD.t3541 VDD.t3540 VDD.t3541 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1986 a_30324_5507.t0 a_50751_n19729.t152 a_51151_n1756# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1987 a_33249_34067.t79 a_33379_34007.t31 a_33249_48695.t109 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1988 a_98829_n21335# a_71281_n8397.t156 a_98299_n21335# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1989 VDD.t3539 VDD.t3538 VDD.t3539 VDD.t1336 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1990 VDD.t3537 VDD.t3536 VDD.t3537 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1991 VSS.t3643 a_94892_4481.t12 a_95414_5639# VSS.t1042 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1992 a_60677_10448.t2 a_53699_11614.t5 a_60109_11614# VDD.t494 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1993 VSS.t2734 VSS.t2733 VSS.t2734 VSS.t327 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1994 a_60845_n19597# a_50751_n19729.t153 a_60285_n19597# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1995 a_101350_12380# a_100820_10448.t6 a_100820_10448.t7 VDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1996 a_33249_34067.t78 a_33379_34007.t32 a_33249_48695.t15 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1997 VSS.t2732 VSS.t2731 VSS.t2732 VSS.t450 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1998 VDD.t3535 VDD.t3534 VDD.t3535 VDD.t394 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1999 a_36530_n28415# a_30152_n36322.t11 VDD.t4773 VSS.t326 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2000 a_106809_n5150.t2 a_103997_n8770.t5 a_113110_n34390# VDD.t330 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2001 a_33249_48695.t278 a_31699_20742.t113 VDD.t136 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2002 VSS.t199 a_35502_25545.t45 a_33249_35053.t135 VSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2003 VDD.t3533 VDD.t3532 VDD.t3533 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2004 a_105365_n21335# a_71281_n8397.t157 a_104527_n21335# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2005 VDD.t541 a_100820_n36322.t12 a_108602_n29181# VSS.t350 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2006 VSS.t2730 VSS.t2729 VSS.t2730 VSS.t106 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2007 VSS.t2728 VSS.t2727 VSS.t2728 VSS.t581 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2008 a_33249_34067.t130 a_35502_25545.t46 VSS.t349 VSS.t142 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2009 VDD.t3531 VDD.t3530 VDD.t3531 VDD.t982 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2010 a_45445_n16904# a_31953_n19727.t156 a_44885_n15110# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2011 VDD.t3529 VDD.t3528 VDD.t3529 VDD.t1302 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2012 VSS.t2726 VSS.t2725 VSS.t2726 VSS.t1030 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2013 VDD.t3527 VDD.t3526 VDD.t3527 VDD.t420 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2014 a_95105_n20430# a_71281_n10073.t137 a_94537_n20430# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2015 a_50751_n19729.t47 a_50751_n19729.t46 VSS.t236 VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2016 OUT.t14 a_35502_24538.t37 a_33249_35053.t90 VSS.t182 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2017 a_89009_4481.t1 a_83153_11614.t17 a_90935_7563# VSS.t398 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2018 VSS.t2724 VSS.t2723 VSS.t2724 VSS.t1472 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2019 VDD.t3525 VDD.t3524 VDD.t3525 VDD.t503 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2020 a_90245_n20430# a_71281_n10073.t138 a_89407_n20430# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2021 VDD.t3523 VDD.t3522 VDD.t3523 VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2022 a_83709_n6960# a_71281_n10073.t139 a_83141_n6960# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2023 VSS.t2722 VSS.t2721 VSS.t2722 VSS.t813 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2024 a_39179_n6239# a_31953_n19727.t157 a_38619_n4445# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2025 VDD.t3521 VDD.t3520 VDD.t3521 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2026 VDD.t3519 VDD.t3518 VDD.t3519 VDD.t723 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2027 VDD.t3517 VDD.t3516 VDD.t3517 VDD.t1167 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2028 VDD.t3515 VDD.t3514 VDD.t3515 VDD.t61 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2029 a_103997_n8770.t2 a_106830_n36382.t11 a_108636_n35156# VDD.t1293 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2030 a_54579_n19597# a_50751_n19729.t154 a_54019_n19597# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2031 VDD.t3513 VDD.t3512 VDD.t3513 VDD.t2352 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2032 a_32353_n16007# a_31953_n19727.t158 a_31284_n30339.t2 VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2033 VSS.t16 a_35502_25545.t47 a_33249_35053.t134 VSS.t15 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2034 a_33249_48695.t16 a_33379_34007.t33 a_33249_34067.t77 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2035 VSS.t2720 VSS.t2719 VSS.t2720 VSS.t861 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2036 VSS.t292 a_112559_4481.t16 a_113081_7563# VSS.t287 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2037 VDD.t3511 VDD.t3510 VDD.t3511 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2038 a_54019_n5344# a_50751_n19729.t155 a_53145_n3550# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2039 a_64243_n19597# a_50751_n19729.t156 a_63683_n19597# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2040 a_49755_n34390# a_47819_n35156.t15 VDD.t4802 VDD.t710 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2041 a_107339_n6055# a_71281_n8397.t158 a_106809_n6055.t1 VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2042 a_32353_n3548# a_31953_n19727.t159 a_31831_n4445# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2043 VDD.t3509 VDD.t3508 VDD.t3509 VDD.t1302 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2044 a_73268_6405# a_65486_11614.t11 a_64243_n1756.t1 VSS.t426 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2045 VSS.t2718 VSS.t2717 VSS.t2718 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2046 a_34347_n3548# a_31953_n19727.t160 a_33787_n3548# VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2047 a_77225_4481.t7 a_77225_4481.t6 a_79151_7563# VSS.t335 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2048 I1U.t1 I1U.t0 VSS.t363 VSS.t362 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X2049 a_88839_n20430# a_71281_n10073.t140 a_88271_n20430# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2050 VDD.t3507 VDD.t3506 VDD.t3507 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2051 a_89407_n7865# a_71281_n10073.t141 a_88839_n7865# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2052 a_33249_48695.t277 a_31699_20742.t114 VDD.t138 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2053 VDD.t3505 VDD.t3504 VDD.t3505 VDD.t1167 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2054 a_95414_5639# a_94892_4481.t13 a_89163_10388.t0 VSS.t1003 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2055 VSS.t2716 VSS.t2715 VSS.t2716 VSS.t873 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2056 VCM.t0 a_106830_n36382.t12 a_108636_n33224# VDD.t1293 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2057 VDD.t3503 VDD.t3502 VDD.t3503 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2058 VSS.t2714 VSS.t2713 VSS.t2714 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2059 a_48313_n15110# a_31953_n19727.t161 a_47753_n14213# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2060 a_52635_48695.t53 a_35922_19591.t78 a_52635_34067.t35 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2061 VDD.t3501 VDD.t3500 VDD.t3501 VDD.t402 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2062 VDD.t3499 VDD.t3498 VDD.t3499 VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2063 a_52635_48695.t151 a_52635_34067.t119 VDD.t4929 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2064 a_46319_n18698# a_31953_n19727.t162 a_45797_n18698# VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2065 a_105933_n18620# a_71281_n8397.t159 a_105365_n18620# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2066 a_105365_n3340# a_71281_n8397.t160 a_104527_n3340# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2067 VSS.t2712 VSS.t2711 VSS.t2712 VSS.t1249 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X2068 VSS.t235 a_50751_n19729.t44 a_50751_n19729.t45 VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2069 a_35922_19591.t5 a_35502_25545.t48 VSS.t38 VSS.t37 nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X2070 VSS.t2710 VSS.t2709 VSS.t2710 VSS.t593 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2071 a_57977_n19597# a_50751_n19729.t157 a_57417_n19597# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2072 VDD.t3497 VDD.t3496 VDD.t3497 VDD.t1268 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2073 VDD.t3495 VDD.t3494 VDD.t3495 VDD.t17 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2074 VSS.t2708 VSS.t2707 VSS.t2708 VSS.t780 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2075 VSS.t2706 VSS.t2705 VSS.t2706 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2076 VDD.t3493 VDD.t3492 VDD.t3493 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2077 VDD.t3491 VDD.t3490 VDD.t3491 VDD.t324 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2078 VDD.t3489 VDD.t3488 VDD.t3489 VDD.t933 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2079 a_106830_n36382.t2 a_112559_n29181.t14 a_114485_n27257# VSS.t414 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2080 VSS.t2704 VSS.t2703 VSS.t2704 VSS.t260 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2081 VSS.t2702 VSS.t2701 VSS.t2702 VSS.t1069 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2082 VDD.t3487 VDD.t3486 VDD.t3487 VDD.t1130 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2083 VSS.t2700 VSS.t2699 VSS.t2700 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2084 VSS.t2698 VSS.t2697 VSS.t2698 VSS.t676 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2085 VSS.t2696 VSS.t2695 VSS.t2696 VSS.t533 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2086 VDD.t3485 VDD.t3484 VDD.t3485 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2087 VSS.t2694 VSS.t2693 VSS.t2694 VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2088 VSS.t2692 VSS.t2691 VSS.t2692 VSS.t411 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2089 VSS.t2690 VSS.t2689 VSS.t2690 VSS.t209 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2090 VSS.t2688 VSS.t2687 VSS.t2688 VSS.t800 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2091 VDD.t3483 VDD.t3482 VDD.t3483 VDD.t405 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2092 VSS.t2686 VSS.t2685 VSS.t2686 VSS.t1437 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2093 VSS.t2684 VSS.t2683 VSS.t2684 VSS.t323 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2094 VDD.t3481 VDD.t3480 VDD.t3481 VDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2095 VDD.t3479 VDD.t3478 VDD.t3479 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2096 a_36008_n30339.t2 a_30152_n36322.t12 a_37934_n27257# VSS.t323 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2097 a_106501_n8770# a_71281_n8397.t161 a_105933_n8770# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2098 VSS.t2682 VSS.t2681 VSS.t2682 VSS.t1320 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2099 a_104527_n18620# a_71281_n8397.t162 a_103997_n19525# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2100 VSS.t2680 VSS.t2679 VSS.t2680 VSS.t336 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2101 VDD.t3477 VDD.t3476 VDD.t3477 VDD.t1268 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2102 a_46319_n7136# a_31953_n19727.t163 a_45797_n8033# VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2103 VSS.t2678 VSS.t2677 VSS.t2678 VSS.t316 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2104 VDD.t3475 VDD.t3474 VDD.t3475 VDD.t572 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X2105 VDD.t3473 VDD.t3472 VDD.t3473 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2106 a_82573_n14095# a_71281_n10073.t142 a_81735_n14095# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2107 a_52635_48695.t52 a_35922_19591.t79 a_52635_34067.t36 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2108 VDD.t139 a_31699_20742.t115 a_33249_48695.t276 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2109 VDD.t141 a_31699_20742.t116 a_33249_48695.t275 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2110 VSS.t2676 VSS.t2675 VSS.t2676 VSS.t297 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2111 a_114516_12380# a_86903_n14095.t6 a_89715_n17715.t3 VDD.t373 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2112 a_95105_n6960# a_71281_n10073.t143 a_94537_n6960# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2113 VSS.t2674 VSS.t2673 VSS.t2674 VSS.t913 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2114 a_52635_49681.t145 a_52635_34067.t120 VDD.t4928 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2115 a_113110_10448# a_100992_4421.t1 a_112559_4481.t1 VDD.t375 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2116 VSS.t2672 VSS.t2671 VSS.t2672 VSS.t738 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2117 VSS.t375 a_41891_n29181.t16 a_42413_n29181# VSS.t171 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2118 VDD.t3471 VDD.t3470 VDD.t3471 VDD.t547 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2119 VSS.t2670 VSS.t2669 VSS.t2670 VSS.t596 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2120 a_33249_48695.t274 a_31699_20742.t117 VDD.t142 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2121 VDD.t3469 VDD.t3468 VDD.t3469 VDD.t1613 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2122 a_66551_n5344# a_50751_n19729.t158 a_65677_n3550# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2123 VDD.t4927 a_52635_34067.t121 a_52635_48695.t150 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2124 VSS.t2668 VSS.t2667 VSS.t2668 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2125 a_35502_24538.t18 a_31699_20742.t118 VDD.t143 VDD.t21 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2126 VSS.t2666 VSS.t2665 VSS.t2666 VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2127 a_48349_10448# a_47819_10448.t7 a_47819_10448.t8 VDD.t497 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2128 a_95105_n15905# a_71281_n10073.t144 a_94537_n15905# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2129 VSS.t2664 VSS.t2663 VSS.t2664 VSS.t839 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2130 a_90245_n18620# a_71281_n10073.t145 a_89407_n15905# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2131 VSS.t2662 VSS.t2661 VSS.t2662 VSS.t253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2132 VDD.t4926 a_52635_34067.t122 a_52635_49681.t144 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2133 VDD.t3467 VDD.t3466 VDD.t3467 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2134 VDD.t3465 VDD.t3464 VDD.t3465 VDD.t1442 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2135 VSS.t2660 VSS.t2659 VSS.t2660 VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2136 a_48313_n8930# a_31953_n19727.t164 a_47753_n8033# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2137 VDD.t3463 VDD.t3462 VDD.t3463 VDD.t1801 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2138 a_89563_n36322# a_89163_n36382.t11 a_89033_n36322.t3 VDD.t549 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2139 OUT.t13 a_35502_24538.t38 a_33249_35053.t91 VSS.t183 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2140 a_59411_n7138# a_50751_n19729.t159 a_58851_n7138# VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2141 VDD.t3461 VDD.t3460 VDD.t3461 VDD.t634 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2142 VDD.t3459 VDD.t3458 VDD.t3459 VDD.t1445 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2143 VDD.t3457 VDD.t3456 VDD.t3457 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2144 VSS.t2658 VSS.t2657 VSS.t2658 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2145 VSS.t332 a_106830_10388.t13 a_107230_12380# VDD.t524 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2146 a_33249_35053.t133 a_35502_25545.t49 VSS.t23 VSS.t22 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2147 VDD.t3455 VDD.t3454 VDD.t3455 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2148 VSS.t2656 VSS.t2655 VSS.t2656 VSS.t148 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2149 a_30682_n34390# a_30152_n35156.t19 a_30152_n36322.t7 VDD.t626 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2150 a_67111_n13318# a_50751_n19729.t160 a_66551_n13318# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2151 VDD.t3453 VDD.t3452 VDD.t3453 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2152 VDD.t3451 VDD.t3450 VDD.t3451 VDD.t2234 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2153 VDD.t3449 VDD.t3448 VDD.t3449 VDD.t1221 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2154 a_33249_35053.t29 a_33379_34917.t31 a_33249_48695.t46 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2155 VDD.t3447 VDD.t3446 VDD.t3447 VDD.t546 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2156 VSS.t2654 VSS.t2653 VSS.t2654 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2157 a_81735_n9675# a_71281_n10073.t146 a_81205_n9675# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2158 VDD.t3445 VDD.t3444 VDD.t3445 VDD.t2302 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X2159 VSS.t2652 VSS.t2651 VSS.t2652 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2160 VSS.t2650 VSS.t2649 VSS.t2650 VSS.t643 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2161 VSS.t2648 VSS.t2647 VSS.t2648 VSS.t913 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2162 a_72603_n10973# I1N.t2 I1N.t3 VSS.t302 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X2163 VSS.t2646 VSS.t2645 VSS.t2646 VSS.t765 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2164 VDD.t144 a_31699_20742.t119 a_33249_48695.t273 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2165 a_98829_n9675# a_71281_n8397.t163 a_98299_n9675# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2166 a_88839_n15905# a_71281_n10073.t147 a_88271_n15905# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2167 VSS.t2644 VSS.t2643 VSS.t2644 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2168 VDD.t3443 VDD.t3442 VDD.t3443 VDD.t1801 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2169 a_30682_12380# a_30152_10448.t10 a_30152_10448.t11 VDD.t351 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2170 VDD.t3441 VDD.t3440 VDD.t3441 VDD.t607 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2171 VDD.t4925 a_52635_34067.t123 a_52635_49681.t143 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2172 VSS.t2642 VSS.t2641 VSS.t2642 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2173 a_42047_n17801# a_31953_n19727.t165 a_41487_n16904# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2174 VSS.t2640 VSS.t2639 VSS.t2640 VSS.t447 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2175 a_77225_n29181.t7 a_77225_n29181.t6 a_79151_n28415# VSS.t386 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2176 VSS.t2638 VSS.t2637 VSS.t2638 VSS.t864 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2177 VDD.t4787 a_83153_n36322.t12 a_90935_n28415# VSS.t460 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2178 a_55635_n34390# a_53829_n36382.t17 VSS.t152 VDD.t296 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2179 VDD.t3439 VDD.t3438 VDD.t3439 VDD.t1221 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2180 VSS.t2636 VSS.t2635 VSS.t2636 VSS.t259 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2181 a_52635_48695.t149 a_52635_34067.t124 VDD.t4924 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2182 VDD.t3437 VDD.t3436 VDD.t3437 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2183 VDD.t3435 VDD.t3434 VDD.t3435 VDD.t311 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2184 a_38619_n13316# a_31953_n19727.t166 a_38097_n13316# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2185 VSS.t2634 VSS.t2633 VSS.t2634 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2186 VDD.t3433 VDD.t3432 VDD.t3433 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2187 VDD.t3431 VDD.t3430 VDD.t3431 VDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2188 a_64243_n1756.t1 a_65486_11614.t12 a_71864_5639# VSS.t429 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2189 a_52585_n17803# a_50751_n19729.t161 a_52063_n18700# VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2190 VSS.t2632 VSS.t2631 VSS.t2632 VSS.t182 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2191 VCM.t2 a_33379_34007.t0 cap_mim_2f0_m4m5_noshield c_width=9.8u c_length=9.8u
X2192 VSS.t2630 VSS.t2629 VSS.t2630 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2193 VDD.t3429 VDD.t3428 VDD.t3429 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2194 a_84547_n8770# a_71281_n10073.t148 a_83709_n8770# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2195 VDD.t3427 VDD.t3426 VDD.t3427 VDD.t933 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2196 VSS.t2628 VSS.t2627 VSS.t2628 VSS.t692 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2197 VDD.t3425 VDD.t3423 VDD.t3425 VDD.t3424 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2198 a_52635_49681.t33 a_35922_19591.t80 OUT.t74 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2199 VDD.t3422 VDD.t3421 VDD.t3422 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2200 a_60109_n34390# a_53699_n35156.t9 a_53829_n36382.t6 VDD.t544 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2201 VDD.t3420 VDD.t3419 VDD.t3420 VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2202 a_33249_35053.t132 a_35502_25545.t50 VSS.t168 VSS.t24 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2203 a_47991_n29313.t0 a_47819_n36322.t12 a_54197_n27257# VSS.t327 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2204 VDD.t3418 VDD.t3417 VDD.t3418 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2205 VDD.t3416 VDD.t3415 VDD.t3416 VDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2206 a_85129_n30339# a_83325_n29313.t0 a_31831_n5342.t1 VSS.t278 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2207 VDD.t3414 VDD.t3413 VDD.t3414 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2208 VDD.t3412 VDD.t3411 VDD.t3412 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2209 a_78344_10448.t3 a_71366_11614.t5 a_77776_13546# VDD.t3571 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2210 a_36032_13546.t3 a_53829_10388.t11 a_55635_13546# VDD.t3748 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2211 a_33249_48695.t47 a_33379_34917.t32 a_33249_35053.t30 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2212 VSS.t2626 VSS.t2625 VSS.t2626 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2213 a_58851_n2653# a_50751_n19729.t162 a_58329_n3550# VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2214 VSS.t2624 VSS.t2623 VSS.t2624 VSS.t692 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2215 a_106676_n30339.t3 a_106830_n36382.t13 a_107230_n36322# VDD.t848 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2216 VDD.t3410 VDD.t3409 VDD.t3410 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2217 VDD.t3408 VDD.t3407 VDD.t3408 VDD.t839 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2218 a_33249_48695.t272 a_31699_20742.t120 VDD.t145 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2219 VDD.t3406 VDD.t3405 VDD.t3406 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2220 a_52635_48695.t148 a_52635_34067.t125 VDD.t4923 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2221 VSS.t2622 VSS.t2621 VSS.t2622 VSS.t1261 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2222 a_81205_n14095.t0 a_89163_10388.t15 a_90969_12380# VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2223 VDD.t3404 VDD.t3403 VDD.t3404 VDD.t1801 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2224 VDD.t3402 VDD.t3401 VDD.t3402 VDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2225 VSS.t2620 VSS.t2619 VSS.t2620 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2226 VDD.t3400 VDD.t3399 VDD.t3400 VDD.t489 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2227 VDD.t3398 VDD.t3397 VDD.t3398 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2228 VDD.t3396 VDD.t3395 VDD.t3396 VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2229 VSS.t2618 VSS.t2617 VSS.t2618 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2230 VDD.t3394 VDD.t3393 VDD.t3394 VDD.t1055 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2231 VSS.t2616 VSS.t2615 VSS.t2616 VSS.t1432 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2232 VDD.t3392 VDD.t3391 VDD.t3392 VDD.t495 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2233 VSS.t2614 VSS.t2613 VSS.t2614 VSS.t762 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2234 VDD.t3390 VDD.t3389 VDD.t3390 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2235 VSS.t2612 VSS.t2611 VSS.t2612 VSS.t327 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2236 VDD.t3388 VDD.t3387 VDD.t3388 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2237 VSS.t2610 VSS.t2609 VSS.t2610 VSS.t658 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2238 a_46879_n19595# a_31953_n19727.t167 a_46319_n19595# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2239 a_78344_10448.t0 a_71366_11614.t6 a_77776_11614# VDD.t3571 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2240 a_53699_11614.t0 a_53829_10388.t12 a_55635_11614# VDD.t3748 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2241 VDD.t3386 VDD.t3385 VDD.t3386 VDD.t826 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2242 a_35922_19591.t1 a_35922_19591.t0 a_46274_24920# VDD.t389 pfet_03v3 ad=0.78p pd=3.7u as=0.78p ps=3.7u w=1.2u l=2u
X2243 VSS.t2608 VSS.t2607 VSS.t2608 VSS.t910 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2244 a_89531_n30339# a_83153_n36322.t13 a_89009_n30339.t0 VSS.t459 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2245 a_113037_n18620# a_71281_n8397.t164 a_112199_n18620# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2246 VSS.t2606 VSS.t2605 VSS.t2606 VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2247 a_40613_n3548# a_31953_n19727.t168 a_41487_n5342# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2248 a_93131_n9675# a_71281_n10073.t149 a_92601_n9675# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2249 VSS.t2604 VSS.t2603 VSS.t2604 VSS.t153 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2250 VDD.t3384 VDD.t3383 VDD.t3384 VDD.t813 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2251 VSS.t2602 VSS.t2601 VSS.t2602 VSS.t223 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2252 VDD.t3382 VDD.t3381 VDD.t3382 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2253 VDD.t3380 VDD.t3379 VDD.t3380 VDD.t79 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2254 VSS.t2600 VSS.t2599 VSS.t2600 VSS.t858 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2255 VDD.t3378 VDD.t3377 VDD.t3378 VDD.t41 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2256 a_39179_n16904# a_31953_n19727.t169 a_38619_n16904# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2257 a_38097_n16007.t2 a_39179_n19595.t0 a_48391_n30339# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2258 a_32913_n8033# a_31953_n19727.t170 a_32353_n7136# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2259 VSS.t2598 VSS.t2597 VSS.t2598 VSS.t686 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2260 VDD.t3376 VDD.t3375 VDD.t3376 VDD.t700 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2261 VDD.t3374 VDD.t3373 VDD.t3374 VDD.t1158 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2262 VDD.t3372 VDD.t3371 VDD.t3372 VDD.t1517 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2263 VDD.t3370 VDD.t3369 VDD.t3370 VDD.t2926 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2264 VDD.t3368 VDD.t3367 VDD.t3368 VDD.t12 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2265 VDD.t3366 VDD.t3365 VDD.t3366 VDD.t1408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2266 VDD.t3364 VDD.t3363 VDD.t3364 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2267 VSS.t2596 VSS.t2595 VSS.t2596 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2268 a_52635_49681.t34 a_35922_19591.t81 OUT.t73 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2269 VSS.t2594 VSS.t2593 VSS.t2594 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2270 VSS.t2592 VSS.t2591 VSS.t2592 VSS.t207 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2271 a_100803_n6960# a_71281_n8397.t165 a_100235_n6960# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2272 a_71281_n8397.t49 a_71281_n8397.t48 VDD.t454 VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2273 VDD.t146 a_31699_20742.t121 a_33249_48695.t271 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2274 a_105365_n2435# a_71281_n8397.t166 a_104527_n2435# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2275 VSS.t2590 VSS.t2589 VSS.t2590 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2276 VSS.t2588 VSS.t2587 VSS.t2588 VSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2277 VSS.t2586 VSS.t2585 VSS.t2586 VSS.t146 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2278 VSS.t2584 VSS.t2583 VSS.t2584 VSS.t873 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2279 a_33249_48695.t270 a_31699_20742.t122 VDD.t147 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2280 a_60285_n16906# a_50751_n19729.t163 a_59763_n16906# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2281 VSS.t2582 VSS.t2581 VSS.t2582 VSS.t0 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2282 a_106830_10388.t7 a_112559_4481.t17 a_114485_4481# VSS.t286 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2283 VSS.t172 a_41891_4481.t18 a_42413_4481# VSS.t171 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2284 a_33249_48695.t269 a_31699_20742.t123 VDD.t148 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2285 a_95443_n36322# a_89033_n35156.t10 a_89163_n36382.t1 VDD.t798 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2286 a_95943_n8770# a_71281_n10073.t150 a_95105_n8770# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2287 VDD.t3362 VDD.t3361 VDD.t3362 VDD.t2467 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2288 VDD.t3360 VDD.t3359 VDD.t3360 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2289 VSS.t2580 VSS.t2579 VSS.t2580 VSS.t901 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2290 VDD.t3358 VDD.t3357 VDD.t3358 VDD.t1158 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2291 VDD.t3356 VDD.t3354 VDD.t3356 VDD.t3355 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2292 a_53699_13546.t3 a_71496_10388.t15 a_73302_13546# VDD.t490 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2293 VDD.t3353 VDD.t3352 VDD.t3353 VDD.t792 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2294 VDD.t3351 VDD.t3350 VDD.t3351 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2295 a_42442_10448# a_30324_4421.t1 a_41891_4481.t8 VDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2296 VDD.t3349 VDD.t3348 VDD.t3349 VDD.t1018 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2297 VDD.t3347 VDD.t3346 VDD.t3347 VDD.t530 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2298 a_114485_6405# a_112559_4481.t18 VSS.t293 VSS.t290 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2299 VSS.t2578 VSS.t2577 VSS.t2578 VSS.t1391 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2300 VDD.t3345 VDD.t3344 VDD.t3345 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2301 VDD.t3343 VDD.t3342 VDD.t3343 VDD.t321 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2302 VSS.t2576 VSS.t2575 VSS.t2576 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2303 VDD.t3341 VDD.t3340 VDD.t3341 VDD.t2122 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2304 VDD.t3339 VDD.t3338 VDD.t3339 VDD.t394 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2305 a_106501_n7865# a_71281_n8397.t167 a_105933_n7865# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2306 a_45445_n14213# a_31953_n19727.t171 a_44885_n14213# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2307 a_104527_n17715# a_71281_n8397.t168 a_103997_n21335# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2308 VDD.t453 a_71281_n8397.t46 a_71281_n8397.t47 VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2309 VDD.t3337 VDD.t3336 VDD.t3337 VDD.t2450 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2310 VSS.t2574 VSS.t2573 VSS.t2574 VSS.t695 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2311 a_71281_n10073.t53 a_71281_n10073.t52 VDD.t340 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2312 VSS.t84 a_31953_n19727.t52 a_31953_n19727.t53 VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2313 a_48313_n4445# a_31953_n19727.t172 a_47753_n3548# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2314 a_112199_n19525# a_71281_n8397.t169 a_111631_n19525# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2315 VSS.t83 a_31953_n19727.t50 a_31953_n19727.t51 VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2316 VDD.t149 a_31699_20742.t124 a_33249_48695.t268 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2317 a_66551_n14215# a_50751_n19729.t164 a_66029_n14215# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2318 a_71366_11614.t1 a_71496_10388.t16 a_73302_11614# VDD.t490 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2319 a_61515_n34390# a_47991_n29313.t1 a_60677_n36322.t1 VDD.t545 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2320 VSS.t2572 VSS.t2571 VSS.t2572 VSS.t649 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2321 VSS.t2570 VSS.t2569 VSS.t2570 VSS.t1320 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2322 a_52635_34067.t62 a_35502_24538.t39 a_33249_34067.t11 VSS.t183 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2323 a_52635_49681.t35 a_35922_19591.t82 OUT.t72 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2324 VSS.t2568 VSS.t2567 VSS.t2568 VSS.t889 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2325 VDD.t333 a_71281_n10073.t50 a_71281_n10073.t51 VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2326 a_104527_n9675# a_71281_n8397.t170 a_103997_n9675# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2327 a_65677_n19597# a_50751_n19729.t165 a_65117_n18700# VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2328 a_112559_n29181.t0 a_100992_n29313.t2 a_114516_n36322# VDD.t331 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2329 a_56895_n16009.t0 a_100992_4421.t2 a_101392_4481# VSS.t174 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2330 VSS.t2566 VSS.t2565 VSS.t2566 VSS.t681 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2331 a_45445_n6239# a_31953_n19727.t173 a_44885_n6239# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2332 a_47819_n36322.t4 a_39179_n19595.t0 a_49795_n29181# VSS.t282 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2333 a_89407_n15000# a_71281_n10073.t151 a_88839_n15000# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2334 VDD.t3335 VDD.t3334 VDD.t3335 VDD.t1325 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2335 a_33249_34067.t76 a_33379_34007.t34 a_33249_48695.t17 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2336 a_32353_n2651# a_31953_n19727.t174 a_31831_n2651# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2337 VSS.t2564 VSS.t2563 VSS.t2564 VSS.t882 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2338 VSS.t2562 VSS.t2561 VSS.t2562 VSS.t283 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2339 a_71281_n8397.t45 a_71281_n8397.t44 VDD.t452 VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2340 a_52635_48695.t147 a_52635_34067.t126 VDD.t4922 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2341 VDD.t3333 VDD.t3332 VDD.t3333 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2342 a_113081_4481# a_112559_4481.t3 a_112559_4481.t4 VSS.t285 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2343 VDD.t3331 VDD.t3330 VDD.t3331 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2344 VSS.t2560 VSS.t2559 VSS.t2560 VSS.t949 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2345 VSS.t2558 VSS.t2557 VSS.t2558 VSS.t489 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X2346 a_100803_n15000# a_71281_n8397.t171 a_100235_n15000# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2347 a_34347_n2651# a_31953_n19727.t175 a_33787_n2651# VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2348 a_65486_11614.t4 a_64243_n1756.t1 a_67462_4481# VSS.t413 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2349 VDD.t3329 VDD.t3328 VDD.t3329 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2350 a_41487_n17801# a_31953_n19727.t176 a_40965_n18698# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2351 a_35781_n7136# a_31953_n19727.t177 a_35221_n7136# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2352 VSS.t2556 VSS.t2555 VSS.t2556 VSS.t816 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2353 a_57977_n12421.t0 a_100820_11614.t9 a_107198_5639# VSS.t188 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2354 VSS.t2554 VSS.t2553 VSS.t2554 VSS.t313 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2355 a_33249_48695.t267 a_31699_20742.t125 VDD.t150 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2356 a_52635_49681.t142 a_52635_34067.t127 VDD.t4921 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2357 VSS.t2552 VSS.t2551 VSS.t2552 VSS.t94 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2358 a_42413_4481# a_41891_4481.t0 a_41891_4481.t1 VSS.t177 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2359 a_35221_n18698# a_31953_n19727.t178 a_34699_n18698# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2360 VDD.t151 a_31699_20742.t126 a_33249_48695.t266 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2361 a_33249_34067.t75 a_33379_34007.t35 a_33249_48695.t341 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2362 a_105933_n21335# a_71281_n8397.t172 a_105365_n21335# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2363 a_79151_4481# a_77225_4481.t15 VSS.t340 VSS.t337 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2364 a_107230_13546# a_106830_10388.t14 OUT.t0 VDD.t527 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2365 a_106809_n5150.t1 a_103997_n8770.t6 a_113110_n36322# VDD.t330 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2366 a_67462_6405# a_64243_n1756.t2 a_63161_n5344.t1 VSS.t412 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2367 VSS.t2550 VSS.t2549 VSS.t2550 VSS.t251 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2368 VDD.t3327 VDD.t3326 VDD.t3327 VDD.t389 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X2369 VSS.t2548 VSS.t2547 VSS.t2548 VSS.t500 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2370 a_33249_48695.t342 a_33379_34007.t36 a_33249_34067.t74 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2371 VSS.t2546 VSS.t2545 VSS.t2546 VSS.t530 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2372 a_35502_25545.t9 a_31699_20742.t127 VDD.t152 VDD.t26 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2373 a_101392_n29181# a_100992_n29313.t0 a_100820_n35156.t1 VSS.t381 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2374 a_72603_n8397# I1N.t7 a_71281_n8397.t1 VSS.t302 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X2375 VSS.t2544 VSS.t2543 VSS.t2544 VSS.t913 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2376 VSS.t2542 VSS.t2541 VSS.t2542 VSS.t797 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2377 a_89163_10388.t1 a_94892_4481.t14 a_96818_6405# VSS.t1349 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2378 VDD.t3325 VDD.t3324 VDD.t3325 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2379 VDD.t3323 VDD.t3322 VDD.t3323 VDD.t2402 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2380 a_107230_11614# a_106830_10388.t15 a_86903_n14095.t1 VDD.t527 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2381 VDD.t3321 VDD.t3320 VDD.t3321 VDD.t2575 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2382 a_84547_n8770# a_71281_n10073.t152 a_83709_n7865# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2383 VDD.t3319 VDD.t3318 VDD.t3319 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2384 a_96818_n27257# a_94892_n29181.t13 VSS.t449 VSS.t447 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2385 VDD.t3317 VDD.t3316 VDD.t3317 VDD.t524 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2386 VDD.t3315 VDD.t3314 VDD.t3315 VDD.t723 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2387 a_104527_n21335# a_71281_n8397.t173 a_103997_n21335# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2388 VDD.t3313 VDD.t3312 VDD.t3313 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2389 a_44885_n17801# a_31953_n19727.t179 a_44363_n17801# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2390 VDD.t3311 VDD.t3310 VDD.t3311 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2391 a_44885_n1754# a_31953_n19727.t180 a_44363_n2651# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2392 a_49755_n36322# a_47819_n35156.t16 VDD.t4803 VDD.t710 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2393 VSS.t2540 VSS.t2539 VSS.t2540 VSS.t704 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2394 VSS.t2538 VSS.t2537 VSS.t2538 VSS.t1069 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2395 VSS.t2536 VSS.t2535 VSS.t2536 VSS.t1162 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2396 VDD.t3309 VDD.t3308 VDD.t3309 VDD.t1089 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2397 a_57417_n5344# a_50751_n19729.t166 a_48951_4481.t0 VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2398 a_46879_n2651# a_31953_n19727.t181 a_46319_n1754# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2399 a_79182_n34390# a_65658_n29313.t1 a_78344_n36322.t2 VDD.t2385 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2400 VSS.t2534 VSS.t2533 VSS.t2534 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2401 a_89407_n20430# a_71281_n10073.t153 a_88839_n20430# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2402 VSS.t2532 VSS.t2531 VSS.t2532 VSS.t673 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2403 VDD.t3307 VDD.t3306 VDD.t3307 VDD.t1145 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2404 VDD.t3305 VDD.t3304 VDD.t3305 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2405 VSS.t2530 VSS.t2529 VSS.t2530 VSS.t558 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2406 a_33249_48695.t343 a_33379_34007.t37 a_33249_34067.t73 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2407 a_51151_n14215# a_50751_n19729.t167 a_50629_n15112# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2408 VSS.t2528 VSS.t2527 VSS.t2528 VSS.t341 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2409 a_100803_n20430# a_71281_n8397.t174 a_100235_n20430# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2410 VSS.t2526 VSS.t2525 VSS.t2526 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2411 VSS.t2524 VSS.t2523 VSS.t2524 VSS.t98 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2412 VSS.t2522 VSS.t2521 VSS.t2522 VSS.t249 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2413 a_50629_n16009.t0 a_83325_4421.t0 a_83725_6405# VSS.t300 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2414 VDD.t4920 a_52635_34067.t128 a_52635_48695.t146 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2415 a_106501_n18620# a_71281_n8397.t175 a_105933_n18620# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2416 VDD.t3303 VDD.t3302 VDD.t3303 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2417 a_114485_n29181# a_112559_n29181.t15 VSS.t421 VSS.t418 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2418 VDD.t3301 VDD.t3300 VDD.t3301 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2419 a_87433_n6055# a_71281_n10073.t154 a_86903_n5150# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2420 OUT.t12 a_35502_24538.t40 a_33249_35053.t92 VSS.t187 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2421 VSS.t2520 VSS.t2519 VSS.t2520 VSS.t620 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2422 VSS.t2518 VSS.t2517 VSS.t2518 VSS.t154 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2423 VDD.t3299 VDD.t3298 VDD.t3299 VDD.t1089 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2424 VSS.t2516 VSS.t2515 VSS.t2516 VSS.t1258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2425 VDD.t4919 a_52635_34067.t129 a_52635_49681.t141 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2426 a_55601_n28415# a_47819_n36322.t13 a_39179_n19595.t0 VSS.t330 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2427 a_50751_n19729.t43 a_50751_n19729.t42 VSS.t234 VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2428 VDD.t3297 VDD.t3296 VDD.t3297 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2429 a_101641_n8770# a_71281_n8397.t176 a_100803_n8770# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2430 VSS.t2514 VSS.t2513 VSS.t2514 VSS.t1261 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2431 a_77776_n34390# a_71366_n35156.t6 a_71496_n36382.t4 VDD.t2347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2432 a_34347_n13316# a_31953_n19727.t182 a_33787_n13316# VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2433 a_67111_n13318# a_50751_n19729.t168 a_66551_n12421# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2434 VDD.t3295 VDD.t3294 VDD.t3295 VDD.t1265 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2435 a_113037_n17715# a_71281_n8397.t177 a_112507_n17715.t1 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2436 VSS.t2512 VSS.t2511 VSS.t2512 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2437 VSS.t2510 VSS.t2509 VSS.t2510 VSS.t1311 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2438 a_96818_6405# a_94892_4481.t15 VSS.t3644 VSS.t1308 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2439 VSS.t2508 VSS.t2507 VSS.t2508 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2440 VSS.t2506 VSS.t2505 VSS.t2506 VSS.t581 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2441 VSS.t2504 VSS.t2503 VSS.t2504 VSS.t896 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2442 VSS.t2502 VSS.t2501 VSS.t2502 VSS.t609 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2443 VDD.t3293 VDD.t3292 VDD.t3293 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2444 VSS.t2500 VSS.t2499 VSS.t2500 VSS.t148 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2445 a_83141_n19525# a_71281_n10073.t155 a_82573_n19525# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2446 VSS.t2498 VSS.t2497 VSS.t2498 VSS.t1299 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2447 VDD.t3291 VDD.t3290 VDD.t3291 VDD.t512 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2448 VSS.t2496 VSS.t2495 VSS.t2496 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2449 VSS.t2494 VSS.t2493 VSS.t2494 VSS.t151 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2450 VSS.t2492 VSS.t2491 VSS.t2492 VSS.t753 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2451 VSS.t2490 VSS.t2489 VSS.t2490 VSS.t1292 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2452 VSS.t2488 VSS.t2487 VSS.t2488 VSS.t325 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2453 VDD.t4792 a_83153_10448.t13 a_83683_13546# VDD.t3355 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2454 VDD.t3289 VDD.t3288 VDD.t3289 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2455 VDD.t153 a_31699_20742.t128 a_33249_48695.t265 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2456 a_95105_n14095# a_71281_n10073.t156 a_94537_n14095# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2457 VDD.t3287 VDD.t3286 VDD.t3287 VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2458 VSS.t2486 VSS.t2485 VSS.t2486 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2459 VSS.t2484 VSS.t2483 VSS.t2484 VSS.t103 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2460 VDD.t3285 VDD.t3284 VDD.t3285 VDD.t1183 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2461 VSS.t2482 VSS.t2480 VSS.t2482 VSS.t2481 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X2462 VDD.t3283 VDD.t3282 VDD.t3283 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2463 a_63683_n16906# a_50751_n19729.t169 a_63161_n17803# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2464 a_90245_n15000# a_71281_n10073.t157 a_89407_n14095# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2465 a_88839_n6960# a_71281_n10073.t158 a_88271_n6960# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2466 VDD.t154 a_31699_20742.t129 a_33249_48695.t264 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2467 a_53675_7563.t0 a_47819_11614.t15 a_55601_4481# VSS.t328 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2468 a_90969_10448# a_89163_10388.t16 a_89009_7563.t3 VDD.t559 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2469 VDD.t3281 VDD.t3280 VDD.t3281 VDD.t1045 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2470 VDD.t38 a_31699_20742.t27 a_31699_20742.t28 VDD.t37 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2471 a_95943_n8770# a_71281_n10073.t159 a_95105_n7865# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2472 a_112559_4481.t2 a_100992_4421.t1 a_114516_13546# VDD.t376 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2473 a_33249_48695.t263 a_31699_20742.t130 VDD.t155 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2474 VDD.t4918 a_52635_34067.t130 a_52635_48695.t145 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2475 VDD.t3279 VDD.t3278 VDD.t3279 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2476 a_33249_35053.t31 a_33379_34917.t33 a_33249_48695.t48 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2477 VSS.t3640 a_36162_n36382.t8 a_36562_n34390# VDD.t2305 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2478 VDD.t4917 a_52635_34067.t131 a_52635_48695.t144 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2479 VSS.t2479 VSS.t2478 VSS.t2479 VSS.t326 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2480 VSS.t2477 VSS.t2476 VSS.t2477 VSS.t503 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2481 VSS.t2475 VSS.t2474 VSS.t2475 VSS.t623 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2482 a_89407_n1530# a_71281_n10073.t160 a_88839_n1530# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2483 VSS.t2473 VSS.t2472 VSS.t2473 VSS.t555 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2484 a_67422_n35156# a_65486_n35156.t19 VDD.t9 VDD.t6 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2485 a_83725_6405# a_83325_4421.t0 a_83153_10448.t1 VSS.t299 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2486 VSS.t319 a_59558_n29181.t16 a_60080_n30339# VSS.t316 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2487 a_81735_n19525# a_71281_n10073.t161 a_81205_n19525# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2488 a_51151_n8932# a_50751_n19729.t170 a_50629_n8932# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2489 a_40053_n8033# a_31953_n19727.t183 a_39531_n8033# VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2490 VDD.t4793 a_83153_10448.t14 a_83683_11614# VDD.t3355 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2491 a_52635_48695.t51 a_35922_19591.t83 a_52635_34067.t37 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2492 a_93969_n9675# a_71281_n10073.t162 a_93131_n9675# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2493 a_53145_n8932# a_50751_n19729.t171 a_52585_n8932# VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2494 VDD.t3277 VDD.t3276 VDD.t3277 VDD.t634 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2495 VDD.t3275 VDD.t3274 VDD.t3275 VDD.t642 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2496 VSS.t2471 VSS.t2470 VSS.t2471 VSS.t822 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X2497 VDD.t3273 VDD.t3272 VDD.t3273 VDD.t1045 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2498 VDD.t3271 VDD.t3270 VDD.t3271 VDD.t73 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2499 VDD.t3269 VDD.t3268 VDD.t3269 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2500 a_112559_4481.t0 a_100992_4421.t1 a_114516_11614# VDD.t376 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2501 VDD.t3267 VDD.t3266 VDD.t3267 VDD.t496 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2502 a_94537_n4245# a_71281_n10073.t163 a_93969_n4245# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2503 a_30682_n36322# a_30152_n35156.t20 a_30152_n36322.t5 VDD.t626 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2504 a_88839_n14095# a_71281_n10073.t164 a_88271_n14095# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2505 a_35781_n19595# a_31953_n19727.t184 a_35221_n19595# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2506 a_41487_n8033# a_31953_n19727.t185 a_40965_n8033# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2507 VDD.t3265 VDD.t3264 VDD.t3265 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2508 VDD.t3263 VDD.t3262 VDD.t3263 VDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2509 VSS.t2469 VSS.t2468 VSS.t2469 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2510 a_35221_n7136# a_31953_n19727.t186 a_34699_n8033# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2511 a_67422_n33224# a_65486_n35156.t20 VDD.t10 VDD.t6 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2512 a_89407_n15905# a_71281_n10073.t165 a_88839_n15905# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2513 VDD.t3261 VDD.t3260 VDD.t3261 VDD.t2257 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2514 VSS.t2467 VSS.t2466 VSS.t2467 VSS.t533 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2515 VDD.t3259 VDD.t3258 VDD.t3259 VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2516 a_112507_n17715.t0 a_71281_n8397.t178 a_112199_n21335# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2517 VDD.t3257 VDD.t3256 VDD.t3257 VDD.t1209 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2518 VDD.t3255 VDD.t3254 VDD.t3255 VDD.t607 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2519 a_100803_n15905# a_71281_n8397.t179 a_100235_n15905# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2520 a_36562_13546# a_36162_10388.t15 a_36032_13546.t1 VDD.t3424 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2521 VSS.t2465 VSS.t2464 VSS.t2465 VSS.t147 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2522 VSS.t2463 VSS.t2462 VSS.t2463 VSS.t326 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2523 VDD.t3253 VDD.t3252 VDD.t3253 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2524 VDD.t3251 VDD.t3250 VDD.t3251 VDD.t602 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2525 a_55635_n36322# a_53829_n36382.t18 a_53675_n27257.t2 VDD.t296 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2526 VSS.t2461 VSS.t2460 VSS.t2461 VSS.t495 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2527 VDD.t3249 VDD.t3248 VDD.t3249 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2528 VDD.t3247 VDD.t3246 VDD.t3247 VDD.t920 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2529 a_41660_19698# a_35502_24538.t41 a_41100_20251# VSS.t189 nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X2530 VSS.t2459 VSS.t2458 VSS.t2459 VSS.t530 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2531 a_65117_n17803# a_50751_n19729.t172 a_64595_n18700# VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2532 a_55601_4481# a_47819_11614.t16 a_47991_4421.t0 VSS.t330 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2533 a_35502_24538.t17 a_31699_20742.t131 VDD.t156 VDD.t15 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2534 VDD.t3245 VDD.t3244 VDD.t3245 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2535 VDD.t3243 VDD.t3242 VDD.t3243 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2536 a_71281_n10073.t49 a_71281_n10073.t48 VDD.t337 VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2537 a_53829_n36382.t2 a_59558_n29181.t17 a_61484_n29181# VSS.t312 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2538 VSS.t2457 VSS.t2456 VSS.t2457 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2539 VDD.t3241 VDD.t3240 VDD.t3241 VDD.t1959 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2540 a_60109_n36322# a_53699_n35156.t10 a_53829_n36382.t7 VDD.t544 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2541 a_59411_n17803# a_50751_n19729.t173 a_58851_n17803# VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2542 VDD.t451 a_71281_n8397.t42 a_71281_n8397.t43 VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2543 a_83141_n6960# a_71281_n10073.t166 a_82573_n6960# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2544 a_36562_11614# a_36162_10388.t16 a_36032_11614.t1 VDD.t3424 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2545 VDD.t3239 VDD.t3238 VDD.t3239 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2546 VDD.t3237 VDD.t3236 VDD.t3237 VDD.t1336 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2547 a_33379_34007.t27 IN_POS.t0 cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
X2548 a_59558_4481.t8 a_59558_4481.t7 a_61484_5639# VSS.t312 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2549 VDD.t3235 VDD.t3234 VDD.t3235 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2550 a_33249_35053.t104 a_35502_24538.t42 OUT.t11 VSS.t191 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2551 VDD.t4784 a_65486_11614.t13 a_73268_6405# VSS.t427 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2552 VDD.t3233 VDD.t3232 VDD.t3233 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2553 a_100235_n6960# a_71281_n8397.t180 a_99667_n6960# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2554 a_83709_n13190# a_71281_n10073.t167 a_83141_n13190# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2555 a_46319_n1754# a_31953_n19727.t187 VSS.t111 VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2556 VDD.t3231 VDD.t3230 VDD.t3231 VDD.t405 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2557 VDD.t3229 VDD.t3228 VDD.t3229 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2558 VSS.t2455 VSS.t2454 VSS.t2455 VSS.t1069 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2559 a_47753_n6239# a_31953_n19727.t188 a_47231_n6239# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2560 VSS.t2453 VSS.t2452 VSS.t2453 VSS.t383 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2561 VDD.t3227 VDD.t3226 VDD.t3227 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2562 VDD.t3225 VDD.t3224 VDD.t3225 VDD.t1938 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2563 a_52635_49681.t36 a_35922_19591.t84 OUT.t71 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2564 VDD.t3223 VDD.t3222 VDD.t3223 VDD.t602 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2565 VSS.t2451 VSS.t2450 VSS.t2451 VSS.t61 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2566 VDD.t3221 VDD.t3220 VDD.t3221 VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2567 VSS.t2449 VSS.t2448 VSS.t2449 VSS.t573 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2568 a_81735_n3340# a_71281_n10073.t168 a_81205_n4245# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2569 a_52635_48695.t143 a_52635_34067.t132 VDD.t4916 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2570 VDD.t3219 VDD.t3218 VDD.t3219 VDD.t836 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2571 a_71281_n8397.t41 a_71281_n8397.t40 VDD.t450 VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2572 VDD.t3217 VDD.t3216 VDD.t3217 VDD.t801 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2573 VSS.t2447 VSS.t2446 VSS.t2447 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2574 a_94892_4481.t9 a_83325_4421.t1 a_96849_13546# VDD.t503 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2575 VDD.t3215 VDD.t3214 VDD.t3215 VDD.t1381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2576 a_99667_n15000# a_71281_n8397.t181 a_98829_n15000# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2577 a_59411_n17803# a_50751_n19729.t174 a_60285_n16009# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2578 a_60677_10448.t3 a_47991_4421.t1 a_60109_10448# VDD.t494 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2579 a_71281_n8397.t39 a_71281_n8397.t38 VDD.t449 VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2580 a_98829_n3340# a_71281_n8397.t182 a_98299_n4245# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2581 VDD.t3213 VDD.t3212 VDD.t3213 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2582 VSS.t82 a_31953_n19727.t48 a_31953_n19727.t49 VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2583 VSS.t2445 VSS.t2444 VSS.t2445 VSS.t61 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2584 VSS.t2443 VSS.t2442 VSS.t2443 VSS.t550 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2585 VSS.t2441 VSS.t2440 VSS.t2441 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2586 VSS.t2439 VSS.t2438 VSS.t2439 VSS.t768 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X2587 a_48313_n2651# a_31953_n19727.t189 a_47753_n2651# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2588 a_111063_n15000# a_71281_n8397.t183 a_110225_n15000# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2589 a_33787_n14213# a_31953_n19727.t190 a_33265_n14213# VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2590 VSS.t2437 VSS.t2436 VSS.t2437 VSS.t506 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2591 a_59411_n2653# a_50751_n19729.t175 a_58851_n1756# VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2592 VDD.t3211 VDD.t3210 VDD.t3211 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2593 a_113037_n6960# a_71281_n8397.t184 a_112199_n6960# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2594 VSS.t2435 VSS.t2434 VSS.t2435 VSS.t819 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2595 VSS.t2433 VSS.t2432 VSS.t2433 VSS.t984 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2596 VDD.t3209 VDD.t3208 VDD.t3209 VDD.t1302 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2597 VSS.t2431 VSS.t2430 VSS.t2431 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2598 VSS.t2429 VSS.t2428 VSS.t2429 VSS.t181 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2599 VDD.t3207 VDD.t3206 VDD.t3207 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2600 VSS.t2427 VSS.t2426 VSS.t2427 VSS.t1162 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2601 a_45445_n5342.t1 a_31953_n19727.t191 a_44885_n5342# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2602 VDD.t3205 VDD.t3204 VDD.t3205 VDD.t1180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2603 VDD.t3203 VDD.t3202 VDD.t3203 VDD.t2682 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2604 a_33249_48695.t49 a_33379_34917.t34 a_33249_35053.t32 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2605 a_30152_10448.t1 a_30324_4421.t0 a_32128_7563# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2606 VDD.t3201 VDD.t3200 VDD.t3201 VDD.t2776 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2607 a_94892_4481.t10 a_83325_4421.t1 a_96849_11614# VDD.t503 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2608 VDD.t3199 VDD.t3198 VDD.t3199 VDD.t982 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2609 VDD.t448 a_71281_n8397.t36 a_71281_n8397.t37 VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2610 VDD.t3197 VDD.t3196 VDD.t3197 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2611 a_33249_35053.t131 a_35502_25545.t51 VSS.t206 VSS.t22 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2612 VSS.t2425 VSS.t2424 VSS.t2425 VSS.t495 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2613 VSS.t2423 VSS.t2422 VSS.t2423 VSS.t839 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2614 a_87433_n4245# a_71281_n10073.t169 a_86903_n4245# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2615 VDD.t3195 VDD.t3194 VDD.t3195 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2616 a_43010_n36322.t2 a_36032_n35156.t5 a_42442_n34390# VDD.t2193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2617 VDD.t3193 VDD.t3192 VDD.t3193 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2618 a_64243_n5344.t1 a_50751_n19729.t176 a_63683_n5344# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2619 a_71864_6405# a_65486_11614.t14 VDD.t4785 VSS.t428 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2620 a_33249_48695.t344 a_33379_34007.t38 a_33249_34067.t72 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2621 VDD.t157 a_31699_20742.t132 a_33249_48695.t262 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2622 a_93131_n13190# a_71281_n10073.t170 a_92601_n16810# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2623 VDD.t3191 VDD.t3190 VDD.t3191 VDD.t1293 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2624 a_101641_n8770# a_71281_n8397.t185 a_100803_n7865# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2625 a_88271_n13190# a_71281_n10073.t171 a_87433_n13190# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2626 a_31953_n19727.t47 a_31953_n19727.t46 VSS.t81 VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2627 a_53145_n17803# a_50751_n19729.t177 a_54019_n16009# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2628 VSS.t2421 VSS.t2420 VSS.t2421 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2629 VDD.t4915 a_52635_34067.t133 a_52635_48695.t142 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2630 a_71342_n30339.t2 a_65486_n36322.t14 a_73268_n27257# VSS.t154 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2631 VDD.t3189 VDD.t3188 VDD.t3189 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2632 a_33249_48695.t261 a_31699_20742.t133 VDD.t158 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2633 VSS.t2419 VSS.t2418 VSS.t2419 VSS.t738 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2634 VDD.t3187 VDD.t3186 VDD.t3187 VDD.t2467 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2635 a_64243_n16009.t1 a_50751_n19729.t178 a_63683_n16009# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2636 VDD.t3185 VDD.t3184 VDD.t3185 VDD.t982 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2637 a_71281_n10073.t47 a_71281_n10073.t46 VDD.t347 VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2638 VSS.t2417 VSS.t2416 VSS.t2417 VSS.t94 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2639 a_52635_49681.t37 a_35922_19591.t85 OUT.t70 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2640 VDD.t3183 VDD.t3182 VDD.t3183 VDD.t2572 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2641 VDD.t3181 VDD.t3180 VDD.t3181 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2642 VSS.t2415 VSS.t2414 VSS.t2415 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2643 VSS.t2413 VSS.t2412 VSS.t2413 VSS.t1162 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2644 a_45138_22884# a_35922_19591.t86 a_44608_22884# VDD.t404 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X2645 a_100820_10448.t11 a_100820_10448.t10 a_102756_13546# VDD.t324 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2646 VDD.t3179 VDD.t3178 VDD.t3179 VDD.t2164 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2647 VSS.t2411 VSS.t2410 VSS.t2411 VSS.t173 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2648 VSS.t2409 VSS.t2408 VSS.t2409 VSS.t146 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2649 VDD.t3177 VDD.t3176 VDD.t3177 VDD.t2159 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2650 a_31831_n5342.t0 a_83325_n29313.t0 a_83725_n29181# VSS.t366 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2651 VSS.t2407 VSS.t2406 VSS.t2407 VSS.t386 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2652 VDD.t3175 VDD.t3174 VDD.t3175 VDD.t1167 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2653 a_32128_n27257# a_30324_n30399.t1 a_31284_n30339.t1 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2654 VSS.t2405 VSS.t2404 VSS.t2405 VSS.t1109 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2655 VDD.t3173 VDD.t3172 VDD.t3173 VDD.t2450 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2656 a_40053_n3548# a_31953_n19727.t192 a_39531_n3548# VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2657 VDD.t3171 VDD.t3170 VDD.t3171 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2658 VSS.t2403 VSS.t2402 VSS.t2403 VSS.t460 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2659 VDD.t3169 VDD.t3168 VDD.t3169 VDD.t947 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2660 a_99667_n20430# a_71281_n8397.t186 a_98829_n20430# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2661 a_102796_7563# a_100992_4421.t0 a_56895_n16009.t0 VSS.t144 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2662 VSS.t2401 VSS.t2400 VSS.t2401 VSS.t464 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2663 VDD.t3167 VDD.t3166 VDD.t3167 VDD.t2146 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2664 a_61515_n36322# a_47991_n29313.t1 a_60677_n36322.t2 VDD.t545 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2665 VSS.t80 a_31953_n19727.t44 a_31953_n19727.t45 VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2666 VDD.t3165 VDD.t3164 VDD.t3165 VDD.t1268 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2667 VSS.t2399 VSS.t2398 VSS.t2399 VSS.t7 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2668 VDD.t3163 VDD.t3162 VDD.t3163 VDD.t63 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2669 a_93131_n3340# a_71281_n10073.t172 a_92601_n4245# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2670 a_73302_12380# a_71496_10388.t17 VSS.t280 VDD.t491 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2671 a_57977_n16009.t1 a_50751_n19729.t179 a_57417_n16009# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2672 VSS.t2397 VSS.t2396 VSS.t2397 VSS.t160 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2673 VSS.t2395 VSS.t2394 VSS.t2395 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2674 VDD.t3161 VDD.t3160 VDD.t3161 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2675 a_111063_n20430# a_71281_n8397.t187 a_110225_n20430# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2676 VSS.t2393 VSS.t2392 VSS.t2393 VSS.t777 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2677 VDD.t3159 VDD.t3158 VDD.t3159 VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2678 a_42047_n13316# a_31953_n19727.t193 a_41487_n12419# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2679 a_100820_10448.t9 a_100820_10448.t8 a_102756_11614# VDD.t324 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2680 a_41487_n3548# a_31953_n19727.t194 a_40965_n3548# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2681 VSS.t2391 VSS.t2390 VSS.t2391 VSS.t457 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2682 a_31699_20742.t26 a_31699_20742.t25 VDD.t36 VDD.t35 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2683 VSS.t2389 VSS.t2388 VSS.t2389 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2684 a_37968_n34390# a_36162_n36382.t9 VSS.t3641 VDD.t2131 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2685 a_52585_n13318# a_50751_n19729.t180 a_52063_n14215# VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2686 VSS.t2387 VSS.t2386 VSS.t2387 VSS.t709 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2687 VDD.t159 a_31699_20742.t134 a_35502_25545.t10 VDD.t26 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2688 a_65486_n35156.t9 a_65658_n29313.t0 a_67462_n30339# VSS.t413 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2689 a_52635_48695.t141 a_52635_34067.t134 VDD.t4914 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2690 VDD.t160 a_31699_20742.t135 a_33249_48695.t260 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2691 a_36530_n27257# a_30152_n36322.t13 a_36008_n27257.t2 VSS.t326 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2692 a_52635_48695.t140 a_52635_34067.t135 VDD.t4913 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2693 a_106501_n21335# a_71281_n8397.t188 a_105933_n21335# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2694 VDD.t3157 VDD.t3156 VDD.t3157 VDD.t390 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2695 VSS.t2385 VSS.t2384 VSS.t2385 VSS.t952 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2696 a_52635_49681.t140 a_52635_34067.t136 VDD.t4912 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2697 VSS.t2383 VSS.t2382 VSS.t2383 VSS.t686 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2698 a_33249_35053.t130 a_35502_25545.t52 VSS.t201 VSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2699 VSS.t2381 VSS.t2380 VSS.t2381 VSS.t573 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2700 VDD.t3155 VDD.t3154 VDD.t3155 VDD.t1442 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2701 VDD.t3153 VDD.t3152 VDD.t3153 VDD.t528 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2702 a_52635_49681.t139 a_52635_34067.t137 VDD.t4911 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2703 a_44363_n16007.t1 a_45445_n19595.t1 a_66058_n28415# VSS.t411 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2704 VSS.t2379 VSS.t2378 VSS.t2379 VSS.t175 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2705 a_85089_13546# a_83153_10448.t15 VDD.t4794 VDD.t1445 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2706 a_41100_20251# a_35502_24538.t0 a_35502_24538.t1 VSS.t184 nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X2707 VDD.t3151 VDD.t3150 VDD.t3151 VDD.t50 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2708 VDD.t4910 a_52635_34067.t138 a_52635_48695.t139 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2709 VDD.t3149 VDD.t3148 VDD.t3149 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2710 VDD.t3147 VDD.t3146 VDD.t3147 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2711 VDD.t3145 VDD.t3144 VDD.t3145 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2712 a_105933_n6960# a_71281_n8397.t189 a_105365_n6960# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2713 a_32913_n1754# a_31953_n19727.t195 a_32353_n1754# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2714 VSS.t2377 VSS.t2376 VSS.t2377 VSS.t145 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2715 VDD.t3143 VDD.t3142 VDD.t3143 VDD.t390 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2716 VSS.t2375 VSS.t2374 VSS.t2375 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2717 a_52635_49681.t38 a_35922_19591.t87 OUT.t69 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2718 VDD.t3141 VDD.t3140 VDD.t3141 VDD.t947 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2719 VDD.t3139 VDD.t3138 VDD.t3139 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2720 a_106501_n1530# a_71281_n8397.t190 a_105933_n1530# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2721 a_113081_n28415# a_112559_n29181.t16 a_106830_n36382.t3 VSS.t415 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2722 VDD.t3137 VDD.t3136 VDD.t3137 VDD.t428 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2723 a_33249_34067.t71 a_33379_34007.t39 a_33249_48695.t345 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2724 VDD.t3135 VDD.t3134 VDD.t3135 VDD.t2402 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2725 VDD.t3133 VDD.t3132 VDD.t3133 VDD.t1442 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2726 a_33249_35053.t129 a_35502_25545.t53 VSS.t276 VSS.t33 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2727 a_85089_11614# a_83153_10448.t16 VDD.t4795 VDD.t1445 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2728 VDD.t3131 VDD.t3130 VDD.t3131 VDD.t2103 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2729 a_52635_34067.t63 a_35502_24538.t43 a_33249_34067.t10 VSS.t191 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2730 a_111063_n9675# a_71281_n8397.t191 a_110225_n9675# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2731 VDD.t3129 VDD.t3128 VDD.t3129 VDD.t535 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2732 VDD.t3127 VDD.t3126 VDD.t3127 VDD.t1102 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2733 a_89563_n35156# a_89163_n36382.t12 a_89033_n35156.t2 VDD.t549 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2734 a_33249_48695.t259 a_31699_20742.t136 VDD.t161 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2735 VDD.t3125 VDD.t3124 VDD.t3125 VDD.t1221 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2736 a_104527_n3340# a_71281_n8397.t192 a_103997_n4245# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2737 a_77225_n29181.t10 a_65658_n29313.t1 a_79182_n34390# VDD.t2100 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2738 VDD.t3123 VDD.t3122 VDD.t3123 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2739 VDD.t3121 VDD.t3120 VDD.t3121 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2740 VDD.t349 a_71281_n10073.t44 a_71281_n10073.t45 VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2741 VSS.t2373 VSS.t2372 VSS.t2373 VSS.t49 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2742 a_111631_n4245# a_71281_n8397.t193 a_111063_n4245# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2743 VSS.t2371 VSS.t2370 VSS.t2371 VSS.t655 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2744 a_52635_34067.t4 a_35502_24538.t44 a_33249_34067.t9 VSS.t187 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2745 VDD.t162 a_31699_20742.t137 a_33249_48695.t258 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2746 a_79182_n36322# a_65658_n29313.t1 a_78344_n36322.t3 VDD.t2385 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2747 VDD.t3119 VDD.t3118 VDD.t3119 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2748 a_67111_n8932# a_50751_n19729.t181 a_66551_n8932# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2749 VSS.t2369 VSS.t2368 VSS.t2369 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2750 a_54019_n14215# a_50751_n19729.t182 a_53497_n14215# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2751 VDD.t3117 VDD.t3116 VDD.t3117 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2752 VSS.t2367 VSS.t2366 VSS.t2367 VSS.t249 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2753 a_71281_n8397.t35 a_71281_n8397.t34 VDD.t447 VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2754 VSS.t2365 VSS.t2364 VSS.t2365 VSS.t329 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2755 VDD.t3115 VDD.t3114 VDD.t3115 VDD.t1115 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2756 VSS.t2363 VSS.t2362 VSS.t2363 VSS.t66 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2757 a_39179_n12419# a_31953_n19727.t196 a_38619_n12419# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2758 VSS.t2361 VSS.t2360 VSS.t2361 VSS.t646 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2759 VSS.t2359 VSS.t2358 VSS.t2359 VSS.t1131 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2760 VDD.t3113 VDD.t3112 VDD.t3113 VDD.t1801 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2761 a_89563_n33224# a_89163_n36382.t13 a_71366_n36322.t0 VDD.t549 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2762 VSS.t2357 VSS.t2356 VSS.t2357 VSS.t211 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2763 VSS.t2355 VSS.t2354 VSS.t2355 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2764 VDD.t3111 VDD.t3110 VDD.t3111 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2765 a_52635_48695.t50 a_35922_19591.t88 a_52635_34067.t38 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2766 VDD.t3109 VDD.t3108 VDD.t3109 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2767 VSS.t2353 VSS.t2352 VSS.t2353 VSS.t576 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2768 VSS.t2351 VSS.t2350 VSS.t2351 VSS.t95 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2769 a_81735_n2435# a_71281_n10073.t173 a_36032_11614.t2 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2770 a_99667_n15905# a_71281_n8397.t194 a_98829_n15905# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2771 a_107198_6405# a_100820_11614.t10 VDD.t416 VSS.t150 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2772 VSS.t2349 VSS.t2348 VSS.t2349 VSS.t1069 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2773 a_47819_10448.t2 a_47991_4421.t0 a_49795_5639# VSS.t282 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2774 VDD.t3107 VDD.t3106 VDD.t3107 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2775 OUT.t68 a_35922_19591.t89 a_52635_49681.t39 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2776 VSS.t391 a_77225_n29181.t14 a_77747_n28415# VSS.t390 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2777 VSS.t2347 VSS.t2346 VSS.t2347 VSS.t536 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2778 VDD.t3105 VDD.t3104 VDD.t3105 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2779 a_33249_48695.t346 a_33379_34007.t40 a_33249_34067.t70 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2780 VDD.t3103 VDD.t3102 VDD.t3103 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2781 a_98829_n2435# a_71281_n8397.t195 VDD.t477 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2782 VSS.t2345 VSS.t2344 VSS.t2345 VSS.t1116 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2783 a_89563_12380# a_89163_10388.t17 a_81205_n14095.t1 VDD.t556 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2784 a_67422_12380# a_65486_10448.t15 VDD.t4752 VDD.t869 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2785 a_111063_n15905# a_71281_n8397.t196 a_110225_n15905# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2786 a_71266_n4019.t1 a_71266_n4019.t0 a_75602_n4019# VDD.t1667 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X2787 a_77776_n36322# a_71366_n35156.t7 a_71496_n36382.t5 VDD.t2347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2788 VDD.t3101 VDD.t3100 VDD.t3101 VDD.t2082 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2789 VDD.t446 a_71281_n8397.t32 a_71281_n8397.t33 VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2790 a_43010_10448.t0 a_30324_4421.t1 a_42442_12380# VDD.t292 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2791 a_61515_13546# a_47991_4421.t1 a_60677_10448.t0 VDD.t495 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2792 VDD.t3099 VDD.t3098 VDD.t3099 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2793 VDD.t3097 VDD.t3096 VDD.t3097 VDD.t2079 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2794 a_33249_48695.t50 a_33379_34917.t35 a_33249_35053.t33 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2795 VSS.t2343 VSS.t2342 VSS.t2343 VSS.t351 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2796 VDD.t3095 VDD.t3094 VDD.t3095 VDD.t858 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2797 VDD.t3093 VDD.t3092 VDD.t3093 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2798 VSS.t2341 VSS.t2340 VSS.t2341 VSS.t563 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2799 a_35781_n2651# a_31953_n19727.t197 a_35221_n1754# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2800 a_32913_n18698# a_31953_n19727.t198 a_32353_n17801# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2801 VDD.t3091 VDD.t3090 VDD.t3091 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2802 a_84017_n5150.t0 a_71281_n10073.t174 a_83709_n1530# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2803 VSS.t2339 VSS.t2338 VSS.t2339 VSS.t399 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2804 VDD.t3089 VDD.t3088 VDD.t3089 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2805 VSS.t2337 VSS.t2336 VSS.t2337 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2806 I1N.t1 I1N.t0 a_75585_n8397# VSS.t301 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X2807 a_85129_7563# a_83325_4421.t0 a_50629_n16009.t1 VSS.t298 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2808 VSS.t443 a_106830_n36382.t14 a_107230_n35156# VDD.t848 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2809 VDD.t3087 VDD.t3086 VDD.t3087 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2810 VSS.t2335 VSS.t2334 VSS.t2335 VSS.t949 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2811 VDD.t3085 VDD.t3084 VDD.t3085 VDD.t839 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2812 a_110225_n17715# a_71281_n8397.t197 a_109695_n16810# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2813 a_61515_11614# a_47991_4421.t1 a_60677_10448.t1 VDD.t495 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2814 VSS.t2333 VSS.t2332 VSS.t2333 VSS.t492 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2815 VDD.t3083 VDD.t3082 VDD.t3083 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2816 VSS.t2331 VSS.t2330 VSS.t2331 VSS.t839 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2817 a_43848_n34390# a_30324_n29313.t2 a_43010_n36322.t2 VDD.t2064 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2818 a_30152_10448.t7 a_30152_10448.t6 a_32088_13546# VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2819 a_110225_n15000# a_71281_n8397.t198 a_109695_n15905# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2820 a_53675_7563.t3 a_53829_10388.t13 a_54229_13546# VDD.t1408 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2821 VSS.t2329 VSS.t2328 VSS.t2329 VSS.t614 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2822 VDD.t3081 VDD.t3080 VDD.t3081 VDD.t816 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2823 a_35502_24538.t16 a_31699_20742.t138 VDD.t163 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2824 a_33249_34067.t69 a_33379_34007.t41 a_33249_48695.t347 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2825 a_31953_n19727.t43 a_31953_n19727.t42 VSS.t79 VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2826 a_89009_7563.t0 a_83153_11614.t18 a_90935_4481# VSS.t398 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2827 a_93969_n13190# a_71281_n10073.t175 a_93131_n13190# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2828 a_78344_10448.t2 a_65658_4421.t2 a_77776_10448# VDD.t3571 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2829 a_53699_13546.t0 a_53829_10388.t14 a_55635_10448# VDD.t3748 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2830 a_36008_n30339.t1 a_36162_n36382.t10 a_36562_n36322# VDD.t2305 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2831 VSS.t2327 VSS.t2326 VSS.t2327 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2832 VDD.t3079 VDD.t3078 VDD.t3079 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2833 VDD.t3077 VDD.t3076 VDD.t3077 VDD.t826 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2834 a_48391_5639# a_47991_5507.t0 a_47819_11614.t7 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2835 VDD.t3075 VDD.t3074 VDD.t3075 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2836 a_52635_48695.t138 a_52635_34067.t139 VDD.t4909 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2837 a_106676_n27257.t2 a_106830_n36382.t15 a_107230_n33224# VDD.t848 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2838 VDD.t3073 VDD.t3072 VDD.t3073 VDD.t81 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2839 VSS.t2325 VSS.t2324 VSS.t2325 VSS.t500 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2840 a_41487_n13316# a_31953_n19727.t199 a_40965_n14213# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2841 VDD.t164 a_31699_20742.t139 a_33249_48695.t257 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2842 VDD.t3071 VDD.t3070 VDD.t3071 VDD.t839 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2843 VSS.t2323 VSS.t2322 VSS.t2323 VSS.t527 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2844 a_38619_n6239# a_31953_n19727.t200 a_38097_n7136# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2845 VSS.t294 a_112559_4481.t19 a_113081_4481# VSS.t287 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2846 VSS.t2321 VSS.t2320 VSS.t2321 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2847 VDD.t3069 VDD.t3068 VDD.t3069 VDD.t938 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2848 VDD.t3067 VDD.t3066 VDD.t3067 VDD.t813 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2849 a_89407_n14095# a_71281_n10073.t176 a_88839_n14095# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2850 VDD.t3065 VDD.t3064 VDD.t3065 VDD.t1158 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2851 VSS.t433 a_53829_10388.t15 a_54229_11614# VDD.t1408 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2852 a_30152_10448.t9 a_30152_10448.t8 a_32088_11614# VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2853 VDD.t3063 VDD.t3062 VDD.t3063 VDD.t28 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2854 VDD.t3061 VDD.t3060 VDD.t3061 VDD.t2302 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X2855 a_52635_49681.t138 a_52635_34067.t140 VDD.t4908 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2856 VDD.t165 a_31699_20742.t140 a_33249_48695.t256 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2857 VDD.t4907 a_52635_34067.t141 a_52635_48695.t137 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2858 a_47753_n5342# a_31953_n19727.t201 a_46879_n7136# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2859 VDD.t3059 VDD.t3058 VDD.t3059 VDD.t826 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2860 a_100803_n14095# a_71281_n8397.t199 a_100235_n14095# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2861 VDD.t3057 VDD.t3056 VDD.t3057 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2862 VSS.t2319 VSS.t2318 VSS.t2319 VSS.t365 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2863 a_48313_n19595# a_31953_n19727.t202 a_47753_n19595# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2864 a_35502_24538.t15 a_31699_20742.t141 VDD.t166 VDD.t15 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2865 VSS.t2317 VSS.t2316 VSS.t2317 VSS.t214 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2866 VSS.t2315 VSS.t2314 VSS.t2315 VSS.t563 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2867 a_33249_48695.t51 a_33379_34917.t36 a_33249_35053.t34 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2868 a_71496_10388.t2 a_77225_4481.t16 a_79151_4481# VSS.t335 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2869 a_71496_n36382.t1 a_77225_n29181.t15 a_79151_n27257# VSS.t386 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2870 VDD.t3055 VDD.t3054 VDD.t3055 VDD.t2257 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2871 VSS.t48 a_35502_25545.t54 a_33249_35053.t128 VSS.t26 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2872 a_93131_n2435# a_71281_n10073.t177 a_71366_11614.t2 VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2873 a_89009_n30339.t1 a_83153_n36322.t14 a_90935_n27257# VSS.t460 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2874 VDD.t3053 VDD.t3052 VDD.t3053 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2875 VSS.t2313 VSS.t2312 VSS.t2313 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2876 VDD.t34 a_31699_20742.t23 a_31699_20742.t24 VDD.t30 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2877 VDD.t3051 VDD.t3050 VDD.t3051 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2878 VSS.t2311 VSS.t2310 VSS.t2311 VSS.t400 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2879 VDD.t3049 VDD.t3048 VDD.t3049 VDD.t813 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2880 a_95443_n35156# a_83325_n29313.t1 a_94892_n29181.t9 VDD.t798 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2881 a_60845_n15112# a_50751_n19729.t183 a_60285_n15112# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2882 VSS.t2309 VSS.t2308 VSS.t2309 VSS.t500 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2883 a_63683_n8035# a_50751_n19729.t184 a_63161_n8932# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2884 VSS.t2307 VSS.t2306 VSS.t2307 VSS.t35 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2885 a_106676_n27257.t1 a_100820_n36322.t13 a_108602_n30339# VSS.t350 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2886 VSS.t2305 VSS.t2304 VSS.t2305 VSS.t503 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2887 a_51711_n16906# a_50751_n19729.t185 a_51151_n16906# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2888 a_44885_n13316# a_31953_n19727.t203 a_44363_n13316# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2889 a_65677_n8932# a_50751_n19729.t186 a_65117_n8035# VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2890 VDD.t3047 VDD.t3046 VDD.t3047 VDD.t61 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2891 VDD.t3045 VDD.t3044 VDD.t3045 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2892 VDD.t3043 VDD.t3042 VDD.t3043 VDD.t1325 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2893 VDD.t3041 VDD.t3040 VDD.t3041 VDD.t304 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2894 VDD.t3039 VDD.t3038 VDD.t3039 VDD.t2352 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2895 VSS.t2303 VSS.t2302 VSS.t2303 VSS.t61 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2896 VSS.t2301 VSS.t2300 VSS.t2301 VSS.t483 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2897 VSS.t2299 VSS.t2298 VSS.t2299 VSS.t652 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2898 a_52635_48695.t49 a_35922_19591.t90 a_52635_34067.t39 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2899 VSS.t2297 VSS.t2296 VSS.t2297 VSS.t1082 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X2900 a_95413_n5150.t0 a_71281_n10073.t178 a_95105_n1530# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2901 VDD.t3037 VDD.t3036 VDD.t3037 VDD.t1352 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2902 a_39179_n8930.t1 a_100820_n36322.t14 a_107198_n28415# VSS.t353 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2903 a_110225_n20430# a_71281_n8397.t200 a_71366_n35156.t0 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2904 a_33249_48695.t52 a_33379_34917.t37 a_33249_35053.t35 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2905 a_95443_n33224# a_83325_n29313.t1 a_94892_n29181.t9 VDD.t798 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2906 VDD.t3035 VDD.t3034 VDD.t3035 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2907 a_60845_n7138# a_50751_n19729.t187 a_60285_n7138# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2908 VSS.t2295 VSS.t2294 VSS.t2295 VSS.t177 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2909 VSS.t2293 VSS.t2292 VSS.t2293 VSS.t330 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2910 a_71366_13546.t2 a_71496_10388.t18 a_73302_10448# VDD.t490 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2911 VDD.t3033 VDD.t3032 VDD.t3033 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2912 VSS.t2291 VSS.t2290 VSS.t2291 VSS.t44 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2913 VSS.t2289 VSS.t2288 VSS.t2289 VSS.t187 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2914 a_33249_48695.t255 a_31699_20742.t142 VDD.t167 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2915 a_54579_n15112# a_50751_n19729.t188 a_54019_n15112# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2916 a_52635_48695.t136 a_52635_34067.t142 VDD.t4906 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2917 a_106830_n36382.t4 a_103997_n8770.t7 a_114516_n35156# VDD.t331 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2918 VDD.t3031 VDD.t3030 VDD.t3031 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2919 VSS.t2287 VSS.t2286 VSS.t2287 VSS.t250 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2920 VDD.t3029 VDD.t3028 VDD.t3029 VDD.t1325 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2921 a_93969_n3340# a_71281_n10073.t179 a_93131_n3340# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2922 VDD.t3027 VDD.t3026 VDD.t3027 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2923 VDD.t3025 VDD.t3024 VDD.t3025 VDD.t564 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2924 a_64243_n16906# a_50751_n19729.t189 a_63683_n15112# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2925 VSS.t2285 VSS.t2284 VSS.t2285 VSS.t896 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2926 VSS.t2283 VSS.t2282 VSS.t2283 VSS.t638 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2927 VDD.t3023 VDD.t3022 VDD.t3023 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2928 VSS.t2281 VSS.t2280 VSS.t2281 VSS.t445 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2929 a_33249_48695.t53 a_33379_34917.t38 a_33249_35053.t36 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2930 a_33249_34067.t129 a_35502_25545.t55 VSS.t29 VSS.t9 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2931 VDD.t445 a_71281_n8397.t30 a_71281_n8397.t31 VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2932 a_37934_n28415# a_30152_n36322.t14 a_30324_n30399.t1 VSS.t324 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2933 a_104527_n2435# a_71281_n8397.t201 VDD.t478 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2934 a_82573_n4245# a_71281_n10073.t180 a_81735_n4245# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2935 a_35221_n15110# a_31953_n19727.t204 a_34699_n16904# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2936 a_106830_n36382.t7 a_103997_n8770.t8 a_114516_n33224# VDD.t331 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2937 VSS.t3645 a_94892_4481.t16 a_95414_6405# VSS.t1042 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2938 a_111631_n15000# a_71281_n8397.t202 a_111063_n15000# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2939 a_73268_7563# a_65486_11614.t15 a_65658_4421.t0 VSS.t426 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2940 VDD.t3021 VDD.t3020 VDD.t3021 VDD.t758 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2941 VDD.t3019 VDD.t3018 VDD.t3019 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2942 a_40053_n2651# a_31953_n19727.t205 a_39531_n3548# VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2943 a_33249_48695.t348 a_33379_34007.t42 a_33249_34067.t68 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2944 VSS.t2279 VSS.t2278 VSS.t2279 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2945 a_67111_n19597# a_50751_n19729.t190 a_66551_n18700# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2946 VSS.t2277 VSS.t2276 VSS.t2277 VSS.t542 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2947 a_106809_n5150.t2 a_100992_n29313.t2 a_113110_n35156# VDD.t330 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2948 a_99667_n4245# a_71281_n8397.t203 a_98829_n4245# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2949 VDD.t168 a_31699_20742.t143 a_35502_25545.t11 VDD.t37 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2950 a_52635_34067.t40 a_35922_19591.t91 a_52635_48695.t48 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2951 VDD.t3017 VDD.t3016 VDD.t3017 VDD.t2302 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X2952 a_46319_n14213# a_31953_n19727.t206 a_45797_n14213# VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2953 VDD.t3015 VDD.t3014 VDD.t3015 VDD.t495 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2954 a_57977_n16906# a_50751_n19729.t191 a_57417_n15112# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2955 VDD.t3013 VDD.t3012 VDD.t3013 VDD.t748 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2956 VDD.t3011 VDD.t3010 VDD.t3011 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2957 a_41487_n2651# a_31953_n19727.t207 a_40965_n3548# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2958 VSS.t2275 VSS.t2274 VSS.t2275 VSS.t617 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2959 VSS.t2273 VSS.t2272 VSS.t2273 VSS.t1030 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2960 VDD.t3009 VDD.t3008 VDD.t3009 VDD.t1145 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2961 VDD.t379 a_71281_n10073.t181 a_89407_n9675# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2962 a_35221_n1754# a_31953_n19727.t208 a_32913_n1754# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2963 VDD.t3007 VDD.t3006 VDD.t3007 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2964 VSS.t2271 VSS.t2270 VSS.t2271 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2965 a_43010_n36322.t0 a_36032_n35156.t6 a_42442_n36322# VDD.t2193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2966 a_108636_12380# a_106830_10388.t16 VSS.t333 VDD.t525 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2967 a_52585_n12421# a_50751_n19729.t192 a_51711_n16009.t0 VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2968 a_57977_n5344.t0 a_50751_n19729.t193 a_57417_n5344# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2969 a_107230_10448# a_106830_10388.t17 a_89033_13546.t2 VDD.t527 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2970 VDD.t3005 VDD.t3004 VDD.t3005 VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2971 a_106809_n5150.t2 a_100992_n29313.t2 a_113110_n33224# VDD.t330 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2972 a_38619_n18698# a_31953_n19727.t209 a_38097_n19595# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2973 VDD.t3003 VDD.t3002 VDD.t3003 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2974 a_37934_5639# a_30152_11614.t10 a_30324_5507.t1 VSS.t324 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2975 VDD.t3001 VDD.t3000 VDD.t3001 VDD.t723 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2976 a_33249_34067.t67 a_33379_34007.t43 a_33249_48695.t349 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2977 a_30152_n36322.t1 a_30324_n30399.t1 a_32128_n29181# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2978 VDD.t4905 a_52635_34067.t143 a_52635_48695.t135 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2979 VDD.t2999 VDD.t2998 VDD.t2999 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2980 VSS.t2269 VSS.t2268 VSS.t2269 VSS.t864 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2981 a_51151_n4447# a_50751_n19729.t194 a_50629_n4447# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2982 VDD.t2997 VDD.t2996 VDD.t2997 VDD.t1089 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2983 VDD.t2995 VDD.t2994 VDD.t2995 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2984 VSS.t2267 VSS.t2266 VSS.t2267 VSS.t313 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2985 a_49755_n35156# a_47819_n35156.t17 VDD.t4804 VDD.t710 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2986 VSS.t376 a_41891_n29181.t17 a_42413_n30339# VSS.t171 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2987 VSS.t14 a_35502_25545.t56 a_33249_35053.t127 VSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2988 VDD.t2993 VDD.t2992 VDD.t2993 VDD.t1145 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2989 a_44885_n8930# a_31953_n19727.t210 a_44363_n8930# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2990 VDD.t335 a_71281_n10073.t42 a_71281_n10073.t43 VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2991 VDD.t2991 VDD.t2990 VDD.t2991 VDD.t1919 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2992 a_50751_n19729.t41 a_50751_n19729.t40 VSS.t233 VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2993 VSS.t422 a_112559_n29181.t17 a_113081_n29181# VSS.t416 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2994 VSS.t2265 VSS.t2264 VSS.t2265 VSS.t800 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2995 VDD.t2989 VDD.t2988 VDD.t2989 VDD.t1265 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2996 a_88271_n6960# a_71281_n10073.t182 a_87433_n6960# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2997 a_33249_35053.t37 a_33379_34917.t39 a_33249_48695.t54 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2998 a_84547_n20430# a_71281_n10073.t183 a_83709_n19525# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2999 VSS.t2263 VSS.t2262 VSS.t2263 VSS.t104 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3000 a_46879_n8930# a_31953_n19727.t211 a_46319_n8930# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3001 VDD.t4904 a_52635_34067.t144 a_52635_48695.t134 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3002 VDD.t2987 VDD.t2986 VDD.t2987 VDD.t2164 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3003 a_87433_n13190# a_71281_n10073.t184 a_86903_n16810# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3004 VDD.t2985 VDD.t2984 VDD.t2985 VDD.t492 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3005 VDD.t2983 VDD.t2982 VDD.t2983 VDD.t2159 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3006 VDD.t2981 VDD.t2980 VDD.t2981 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3007 VSS.t2261 VSS.t2260 VSS.t2261 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3008 VDD.t2979 VDD.t2978 VDD.t2979 VDD.t723 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3009 VSS.t2259 VSS.t2258 VSS.t2259 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3010 VSS.t2257 VSS.t2256 VSS.t2257 VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3011 a_95414_6405# a_94892_4481.t6 a_94892_4481.t7 VSS.t1003 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3012 a_110225_n15905# a_71281_n8397.t204 a_109695_n15905# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3013 a_107230_n34390# a_106830_n36382.t16 a_103997_n8770.t3 VDD.t1906 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3014 VDD.t2977 VDD.t2976 VDD.t2977 VDD.t65 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3015 VSS.t2255 VSS.t2254 VSS.t2255 VSS.t495 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3016 VSS.t2253 VSS.t2252 VSS.t2253 VSS.t480 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3017 VSS.t451 a_94892_n29181.t14 a_95414_n28415# VSS.t450 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3018 a_49755_n33224# a_47819_n35156.t18 VDD.t4805 VDD.t710 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3019 VDD.t2975 VDD.t2974 VDD.t2975 VDD.t491 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3020 a_111631_n20430# a_71281_n8397.t205 a_111063_n20430# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3021 VDD.t2973 VDD.t2972 VDD.t2973 VDD.t390 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3022 VSS.t2251 VSS.t2250 VSS.t2251 VSS.t596 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3023 VDD.t2971 VDD.t2970 VDD.t2971 VDD.t2146 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3024 VSS.t2249 VSS.t2248 VSS.t2249 VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3025 VSS.t2247 VSS.t2246 VSS.t2247 VSS.t949 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3026 VDD.t2969 VDD.t2968 VDD.t2969 VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3027 VDD.t2967 VDD.t2966 VDD.t2967 VDD.t1265 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3028 VSS.t34 a_35502_25545.t57 a_33249_35053.t126 VSS.t33 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3029 VSS.t2245 VSS.t2244 VSS.t2245 VSS.t593 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3030 VSS.t2243 VSS.t2242 VSS.t2243 VSS.t581 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3031 a_36032_n35156.t1 a_36162_n36382.t11 a_37968_n34390# VDD.t1895 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3032 VDD.t2965 VDD.t2964 VDD.t2965 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3033 VSS.t2241 VSS.t2240 VSS.t2241 VSS.t643 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3034 VSS.t2239 VSS.t2238 VSS.t2239 VSS.t37 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X3035 VSS.t2237 VSS.t2236 VSS.t2237 VSS.t211 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3036 a_43848_12380# a_36032_11614.t9 a_43010_10448.t1 VDD.t293 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3037 VSS.t2235 VSS.t2234 VSS.t2235 VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3038 VDD.t2963 VDD.t2962 VDD.t2963 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3039 a_31953_n19727.t41 a_31953_n19727.t40 VSS.t78 VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3040 a_37968_n36322# a_36162_n36382.t12 a_36008_n27257.t0 VDD.t2131 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3041 VDD.t169 a_31699_20742.t144 a_35502_24538.t14 VDD.t30 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3042 a_65117_n13318# a_50751_n19729.t195 a_64595_n14215# VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3043 VSS.t2233 VSS.t2232 VSS.t2233 VSS.t1827 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X3044 VDD.t170 a_31699_20742.t145 a_33249_48695.t254 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3045 VDD.t2961 VDD.t2960 VDD.t2961 VDD.t1886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3046 a_52635_49681.t40 a_35922_19591.t92 OUT.t67 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3047 VSS.t2231 VSS.t2230 VSS.t2231 VSS.t99 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3048 a_63683_n3550# a_50751_n19729.t196 a_63161_n4447# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3049 VSS.t2229 VSS.t2228 VSS.t2229 VSS.t500 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3050 VDD.t479 a_71281_n8397.t206 a_100803_n1530# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3051 VDD.t171 a_31699_20742.t146 a_33249_48695.t253 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3052 a_40053_n17801# a_31953_n19727.t212 a_39531_n18698# VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3053 a_33249_34067.t66 a_33379_34007.t44 a_33249_48695.t350 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3054 VDD.t4903 a_52635_34067.t145 a_52635_49681.t137 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3055 VSS.t2227 VSS.t2226 VSS.t2227 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3056 a_59411_n13318# a_50751_n19729.t197 a_58851_n13318# VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3057 a_65117_n8035# a_50751_n19729.t198 a_64595_n8035# VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3058 VDD.t2959 VDD.t2958 VDD.t2959 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3059 VDD.t2957 VDD.t2956 VDD.t2957 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3060 a_36162_n36382.t6 a_41891_n29181.t18 a_43817_n29181# VSS.t181 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3061 VDD.t2955 VDD.t2954 VDD.t2955 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3062 a_65677_n3550# a_50751_n19729.t199 a_65117_n3550# VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3063 VDD.t2953 VDD.t2952 VDD.t2953 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3064 VSS.t2225 VSS.t2224 VSS.t2225 VSS.t692 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3065 VDD.t2951 VDD.t2950 VDD.t2951 VDD.t1045 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3066 VSS.t2223 VSS.t2222 VSS.t2223 VSS.t765 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3067 a_47819_10448.t4 a_47819_10448.t3 a_49755_13546# VDD.t496 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3068 VDD.t2949 VDD.t2948 VDD.t2949 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3069 VSS.t2221 VSS.t2220 VSS.t2221 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3070 a_50751_n19729.t73 a_71266_n4019.t0 a_75602_n4978# VDD.t1667 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3071 VDD.t2947 VDD.t2946 VDD.t2947 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3072 VDD.t2945 VDD.t2944 VDD.t2945 VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3073 VDD.t2943 VDD.t2942 VDD.t2943 VDD.t6 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3074 VDD.t2941 VDD.t2940 VDD.t2941 VDD.t428 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3075 VDD.t338 a_71281_n10073.t40 a_71281_n10073.t41 VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3076 VDD.t2939 VDD.t2938 VDD.t2939 VDD.t292 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3077 VDD.t2937 VDD.t2936 VDD.t2937 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3078 VDD.t2935 VDD.t2934 VDD.t2935 VDD.t652 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3079 VDD.t2933 VDD.t2932 VDD.t2933 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3080 VDD.t2931 VDD.t2930 VDD.t2931 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3081 a_83153_11614.t5 a_83153_10448.t17 a_85089_12380# VDD.t647 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3082 VDD.t2929 VDD.t2928 VDD.t2929 VDD.t1209 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3083 VSS.t2219 VSS.t2218 VSS.t2219 VSS.t819 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3084 VDD.t4796 a_83153_10448.t18 a_83683_10448# VDD.t3355 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3085 VDD.t2927 VDD.t2925 VDD.t2927 VDD.t2926 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3086 VDD.t2924 VDD.t2922 VDD.t2924 VDD.t2923 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3087 VDD.t2921 VDD.t2920 VDD.t2921 VDD.t2103 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3088 a_71281_n8397.t29 a_71281_n8397.t28 VDD.t444 VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3089 VDD.t2919 VDD.t2918 VDD.t2919 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3090 a_47819_10448.t6 a_47819_10448.t5 a_49755_11614# VDD.t496 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3091 VDD.t2917 VDD.t2916 VDD.t2917 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3092 VDD.t2915 VDD.t2914 VDD.t2915 VDD.t634 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3093 VSS.t2217 VSS.t2216 VSS.t2217 VSS.t839 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3094 a_107339_n8770# a_71281_n8397.t207 a_106501_n8770# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3095 a_77225_n29181.t8 a_65658_n29313.t1 a_79182_n36322# VDD.t2100 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3096 VDD.t172 a_31699_20742.t147 a_33249_48695.t252 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3097 a_45445_n19595.t0 a_31953_n19727.t213 a_44885_n19595# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3098 a_106830_10388.t2 a_86903_n14095.t7 a_114516_10448# VDD.t376 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3099 a_30682_n35156# a_30152_n35156.t4 a_30152_n35156.t5 VDD.t626 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3100 a_34347_n14213# a_31953_n19727.t214 a_35221_n16007# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3101 VDD.t4758 a_83153_n35156.t12 a_83683_n34390# VDD.t1852 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3102 a_58851_n8932# a_50751_n19729.t200 VSS.t265 VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3103 VSS.t43 a_35502_25545.t58 a_33249_34067.t128 VSS.t11 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3104 OUT.t66 a_35922_19591.t93 a_52635_49681.t41 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3105 VDD.t2913 VDD.t2912 VDD.t2913 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3106 VSS.t2215 VSS.t2214 VSS.t2215 VSS.t658 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3107 VDD.t2911 VDD.t2910 VDD.t2911 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3108 VDD.t2909 VDD.t2908 VDD.t2909 VDD.t1209 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3109 a_93969_n2435# a_71281_n10073.t185 a_93131_n2435# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3110 VSS.t2213 VSS.t2212 VSS.t2213 VSS.t533 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3111 a_99667_n14095# a_71281_n8397.t208 a_98829_n14095# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3112 a_66551_n19597# a_50751_n19729.t201 a_64243_n19597# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3113 VDD.t2907 VDD.t2906 VDD.t2907 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3114 a_55601_n27257# a_47819_n36322.t14 a_47991_n29313.t0 VSS.t330 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3115 VDD.t2905 VDD.t2904 VDD.t2905 VDD.t607 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3116 VDD.t2903 VDD.t2902 VDD.t2903 VDD.t634 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3117 VDD.t2901 VDD.t2900 VDD.t2901 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3118 a_111063_n14095# a_71281_n8397.t209 a_110225_n14095# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3119 VSS.t2211 VSS.t2210 VSS.t2211 VSS.t1432 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3120 VSS.t2209 VSS.t2208 VSS.t2209 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3121 a_30682_n33224# a_30152_n35156.t2 a_30152_n35156.t3 VDD.t626 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3122 a_113037_n6055# a_71281_n8397.t210 a_112507_n6055.t1 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3123 a_55635_n35156# a_53829_n36382.t19 VSS.t348 VDD.t296 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3124 VDD.t2899 VDD.t2898 VDD.t2899 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3125 VSS.t403 a_59558_4481.t12 a_60080_5639# VSS.t316 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3126 a_111631_n15905# a_71281_n8397.t211 a_111063_n15905# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3127 a_31699_17542# I1U.t3 a_30377_18342# VSS.t362 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X3128 VSS.t2207 VSS.t2206 VSS.t2207 VSS.t896 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3129 a_38619_n5342# a_31953_n19727.t215 a_38097_n5342.t2 VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3130 a_64243_n1756.t1 a_65486_11614.t16 a_71864_6405# VSS.t429 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3131 a_33249_48695.t351 a_33379_34007.t45 a_33249_34067.t65 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3132 VDD.t2897 VDD.t2896 VDD.t2897 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3133 VDD.t2895 VDD.t2894 VDD.t2895 VDD.t1826 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3134 VSS.t2205 VSS.t2204 VSS.t2205 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3135 a_83153_10448.t3 a_83325_4421.t0 a_85129_5639# VSS.t297 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3136 VSS.t2203 VSS.t2202 VSS.t2203 VSS.t913 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3137 VDD.t2893 VDD.t2892 VDD.t2893 VDD.t1823 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3138 VSS.t232 a_50751_n19729.t38 a_50751_n19729.t39 VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3139 VDD.t2891 VDD.t2890 VDD.t2891 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3140 a_95413_n16810.t0 a_71281_n10073.t186 a_95105_n13190# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3141 VDD.t2889 VDD.t2888 VDD.t2889 VDD.t324 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3142 VCM.t3 a_33379_34007.t1 cap_mim_2f0_m4m5_noshield c_width=9.8u c_length=9.8u
X3143 VDD.t2887 VDD.t2886 VDD.t2887 VDD.t855 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3144 VDD.t2885 VDD.t2884 VDD.t2885 VDD.t2082 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3145 VDD.t2883 VDD.t2882 VDD.t2883 VDD.t607 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3146 a_52635_48695.t47 a_35922_19591.t94 a_52635_34067.t41 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3147 VDD.t2881 VDD.t2880 VDD.t2881 VDD.t2079 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3148 a_65486_10448.t3 a_65486_10448.t2 a_67422_13546# VDD.t1381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3149 a_60109_n35156# a_47991_n29313.t1 a_59558_n29181.t8 VDD.t544 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3150 VDD.t173 a_31699_20742.t148 a_33249_48695.t251 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3151 VSS.t2201 VSS.t2200 VSS.t2201 VSS.t384 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3152 a_35502_24538.t13 a_31699_20742.t149 VDD.t174 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3153 a_113110_n34390# a_103997_n8770.t9 a_106830_n36382.t6 VDD.t328 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3154 a_36562_10448# a_36162_10388.t17 a_33379_34917.t1 VDD.t3424 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3155 a_33249_34067.t64 a_33379_34007.t46 a_33249_48695.t2 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3156 VDD.t4902 a_52635_34067.t146 a_52635_49681.t136 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3157 a_55635_n33224# a_53829_n36382.t20 a_53675_n30339.t3 VDD.t296 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3158 VDD.t2879 VDD.t2878 VDD.t2879 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3159 VSS.t2199 VSS.t2198 VSS.t2199 VSS.t777 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3160 a_35502_25545.t12 a_31699_20742.t150 VDD.t175 VDD.t35 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3161 a_82573_n18620# a_71281_n10073.t187 a_81735_n18620# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3162 a_111063_n3340# a_71281_n8397.t212 a_110225_n3340# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3163 a_33249_35053.t125 a_35502_25545.t59 VSS.t27 VSS.t26 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3164 VDD.t2877 VDD.t2876 VDD.t2877 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3165 VSS.t2197 VSS.t2196 VSS.t2197 VSS.t692 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3166 a_52635_48695.t133 a_52635_34067.t147 VDD.t4901 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3167 VSS.t2195 VSS.t2194 VSS.t2195 VSS.t726 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3168 VSS.t2193 VSS.t2192 VSS.t2193 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3169 a_41891_n29181.t2 a_30324_n29313.t2 a_43848_n34390# VDD.t1798 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3170 VDD.t2875 VDD.t2874 VDD.t2875 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3171 VDD.t2873 VDD.t2872 VDD.t2873 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3172 VDD.t2871 VDD.t2870 VDD.t2871 VDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3173 a_46319_n8930# a_31953_n19727.t216 a_45445_n5342.t0 VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3174 a_65486_10448.t7 a_65486_10448.t6 a_67422_11614# VDD.t1381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3175 a_60109_n33224# a_47991_n29313.t1 a_59558_n29181.t8 VDD.t544 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3176 a_94537_n13190# a_71281_n10073.t188 a_93969_n13190# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3177 VSS.t2191 VSS.t2190 VSS.t2191 VSS.t286 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3178 VSS.t2189 VSS.t2188 VSS.t2189 VSS.t171 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3179 a_43848_n36322# a_30324_n29313.t2 a_43010_n36322.t0 VDD.t2064 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3180 VDD.t2869 VDD.t2868 VDD.t2869 VDD.t1749 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3181 VDD.t2867 VDD.t2866 VDD.t2867 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3182 VDD.t2865 VDD.t2864 VDD.t2865 VDD.t1782 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3183 a_52635_34067.t34 a_35922_19591.t95 a_52635_48695.t46 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3184 VDD.t2863 VDD.t2862 VDD.t2863 VDD.t402 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3185 VSS.t2187 VSS.t2186 VSS.t2187 VSS.t156 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3186 VSS.t2185 VSS.t2184 VSS.t2185 VSS.t411 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3187 VSS.t2183 VSS.t2182 VSS.t2183 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3188 a_33249_34067.t63 a_33379_34007.t47 a_33249_48695.t3 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3189 VDD.t2861 VDD.t2860 VDD.t2861 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3190 VDD.t2859 VDD.t2858 VDD.t2859 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3191 a_114485_7563# a_112559_4481.t20 VSS.t295 VSS.t290 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3192 VSS.t2181 VSS.t2180 VSS.t2181 VSS.t1391 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3193 VSS.t2179 VSS.t2178 VSS.t2179 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3194 a_60845_n7138# a_50751_n19729.t202 a_60285_n6241# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3195 a_33249_48695.t55 a_33379_34917.t40 a_33249_35053.t38 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3196 a_47819_n35156.t10 a_47991_n29313.t0 a_49795_n30339# VSS.t282 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3197 VDD.t176 a_31699_20742.t151 a_33249_48695.t250 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3198 a_52635_48695.t132 a_52635_34067.t148 VDD.t4900 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3199 VDD.t2857 VDD.t2856 VDD.t2857 VDD.t982 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3200 a_65677_n14215# a_50751_n19729.t203 a_65117_n14215# VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3201 a_51151_n19597# a_50751_n19729.t204 a_50629_n19597# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3202 VDD.t2855 VDD.t2854 VDD.t2855 VDD.t123 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3203 a_51711_n8035# a_50751_n19729.t205 a_51151_n8035# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3204 VDD.t4899 a_52635_34067.t149 a_52635_49681.t135 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3205 VSS.t2177 VSS.t2176 VSS.t2177 VSS.t415 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3206 VDD.t2853 VDD.t2852 VDD.t2853 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3207 a_89163_10388.t4 a_81205_n14095.t4 a_96849_10448# VDD.t503 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3208 VSS.t2175 VSS.t2174 VSS.t2175 VSS.t695 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3209 VDD.t2851 VDD.t2850 VDD.t2851 VDD.t801 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3210 a_54229_12380# a_53829_10388.t16 a_53699_11614.t1 VDD.t3679 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3211 VSS.t2173 VSS.t2172 VSS.t2173 VSS.t250 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3212 VDD.t2849 VDD.t2848 VDD.t2849 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3213 a_33249_48695.t249 a_31699_20742.t152 VDD.t177 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3214 VSS.t2171 VSS.t2170 VSS.t2171 VSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3215 VDD.t4898 a_52635_34067.t150 a_52635_48695.t131 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3216 VDD.t2847 VDD.t2846 VDD.t2847 VDD.t965 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X3217 VDD.t2845 VDD.t2844 VDD.t2845 VDD.t52 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3218 VSS.t2169 VSS.t2168 VSS.t2169 VSS.t174 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3219 VSS.t2167 VSS.t2166 VSS.t2167 VSS.t681 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3220 VSS.t2165 VSS.t2164 VSS.t2165 VSS.t495 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3221 a_60285_n5344# a_50751_n19729.t206 a_59411_n3550# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3222 VDD.t2843 VDD.t2842 VDD.t2843 VDD.t401 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X3223 VSS.t2163 VSS.t2162 VSS.t2163 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3224 a_65117_n3550# a_50751_n19729.t207 a_64595_n3550# VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3225 VDD.t2841 VDD.t2840 VDD.t2841 VDD.t123 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3226 a_35221_n14213# a_31953_n19727.t217 a_34699_n14213# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3227 VDD.t2839 VDD.t2838 VDD.t2839 VDD.t2467 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3228 VSS.t2161 VSS.t2160 VSS.t2161 VSS.t285 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3229 a_34347_n19595# a_31953_n19727.t218 a_33787_n18698# VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3230 VDD.t2837 VDD.t2836 VDD.t2837 VDD.t1422 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3231 VSS.t2159 VSS.t2158 VSS.t2159 VSS.t1249 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X3232 VDD.t2835 VDD.t2834 VDD.t2835 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3233 VDD.t2833 VDD.t2832 VDD.t2833 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3234 a_101392_n30339# a_39179_n8930.t1 a_100820_n36322.t7 VSS.t381 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3235 VSS.t2157 VSS.t2156 VSS.t2157 VSS.t413 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3236 a_71281_n8397.t27 a_71281_n8397.t26 VDD.t442 VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3237 VSS.t2155 VSS.t2154 VSS.t2155 VSS.t325 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3238 VDD.t2831 VDD.t2830 VDD.t2831 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3239 VSS.t46 a_35502_25545.t60 a_33249_34067.t127 VSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3240 a_52635_48695.t45 a_35922_19591.t96 a_52635_34067.t42 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3241 VSS.t2153 VSS.t2152 VSS.t2153 VSS.t177 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3242 VSS.t2151 VSS.t2150 VSS.t2151 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3243 VDD.t178 a_31699_20742.t153 a_35502_24538.t12 VDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3244 VDD.t179 a_31699_20742.t154 a_33249_48695.t248 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3245 VSS.t2149 VSS.t2148 VSS.t2149 VSS.t337 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3246 VSS.t2147 VSS.t2146 VSS.t2147 VSS.t1366 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3247 a_67462_7563# a_65658_4421.t0 a_63161_n5344.t1 VSS.t412 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3248 VDD.t2829 VDD.t2828 VDD.t2829 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3249 a_52585_n7138# a_50751_n19729.t208 a_52063_n8035# VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3250 VDD.t2827 VDD.t2826 VDD.t2827 VDD.t426 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3251 VDD.t2825 VDD.t2824 VDD.t2825 VDD.t2450 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3252 a_67111_n4447# a_50751_n19729.t209 a_66551_n4447# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3253 VSS.t2145 VSS.t2144 VSS.t2145 VSS.t910 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3254 VDD.t2823 VDD.t2822 VDD.t2823 VDD.t2467 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3255 VDD.t2821 VDD.t2820 VDD.t2821 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3256 VSS.t2143 VSS.t2142 VSS.t2143 VSS.t390 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3257 VDD.t2819 VDD.t2818 VDD.t2819 VDD.t2264 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3258 VDD.t2817 VDD.t2816 VDD.t2817 VDD.t783 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3259 a_52635_49681.t134 a_52635_34067.t151 VDD.t4897 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3260 a_54579_n7138# a_50751_n19729.t210 a_54019_n7138# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3261 VSS.t2141 VSS.t2140 VSS.t2141 VSS.t314 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3262 a_33249_48695.t247 a_31699_20742.t155 VDD.t180 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3263 a_61515_n35156# a_53699_n35156.t11 a_60677_n36322.t3 VDD.t545 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3264 a_52635_48695.t130 a_52635_34067.t152 VDD.t4896 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3265 VSS.t2139 VSS.t2138 VSS.t2139 VSS.t542 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3266 a_94892_4481.t5 a_94892_4481.t4 a_96818_7563# VSS.t1349 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3267 VSS.t31 a_35502_25545.t61 a_33249_34067.t126 VSS.t15 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3268 a_71864_n28415# a_65486_n36322.t15 VDD.t297 VSS.t153 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3269 a_100820_11614.t0 a_100820_10448.t14 a_102756_10448# VDD.t324 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3270 VDD.t2815 VDD.t2813 VDD.t2815 VDD.t2814 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3271 VSS.t2137 VSS.t2136 VSS.t2137 VSS.t858 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3272 VSS.t2135 VSS.t2134 VSS.t2135 VSS.t558 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3273 VSS.t2133 VSS.t2132 VSS.t2133 VSS.t882 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3274 a_52635_48695.t129 a_52635_34067.t153 VDD.t4895 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3275 VDD.t2812 VDD.t2811 VDD.t2812 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3276 VDD.t2810 VDD.t2809 VDD.t2810 VDD.t2450 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3277 VSS.t21 a_35502_25545.t62 a_35922_19591.t4 VSS.t20 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X3278 VDD.t2808 VDD.t2807 VDD.t2808 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3279 VDD.t2806 VDD.t2805 VDD.t2806 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3280 VDD.t2804 VDD.t2803 VDD.t2804 VDD.t37 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3281 a_31284_n30339.t0 a_30324_n30399.t1 a_30724_n28415# VSS.t146 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3282 a_107339_n8770# a_71281_n8397.t213 a_106501_n7865# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3283 a_57977_n12421.t0 a_100820_11614.t11 a_107198_6405# VSS.t188 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3284 a_71896_12380# a_71496_10388.t19 a_71366_11614.t1 VDD.t488 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3285 a_47753_n16904# a_31953_n19727.t219 a_47231_n16904# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3286 a_114485_n30339# a_112559_n29181.t18 VSS.t423 VSS.t418 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3287 a_61515_n33224# a_53699_n35156.t12 a_60677_n36322.t1 VDD.t545 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3288 VSS.t2131 VSS.t2130 VSS.t2131 VSS.t1069 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3289 VSS.t2129 VSS.t2128 VSS.t2129 VSS.t819 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3290 a_95414_n29181# a_94892_n29181.t6 a_94892_n29181.t7 VSS.t446 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3291 VDD.t2802 VDD.t2801 VDD.t2802 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3292 a_52635_48695.t44 a_35922_19591.t97 a_52635_34067.t13 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3293 VSS.t2127 VSS.t2126 VSS.t2127 VSS.t94 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3294 VSS.t2125 VSS.t2124 VSS.t2125 VSS.t104 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3295 VDD.t2800 VDD.t2799 VDD.t2800 VDD.t1102 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3296 a_32913_n14213# a_31953_n19727.t220 a_32353_n13316# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3297 VDD.t181 a_31699_20742.t156 a_33249_48695.t246 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3298 VDD.t2798 VDD.t2797 VDD.t2798 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3299 VSS.t2123 VSS.t2122 VSS.t2123 VSS.t901 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3300 VSS.t2121 VSS.t2120 VSS.t2121 VSS.t255 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3301 a_33249_48695.t56 a_33379_34917.t41 a_33249_35053.t39 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3302 VSS.t2119 VSS.t2118 VSS.t2119 VSS.t159 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3303 a_52635_49681.t42 a_35922_19591.t98 OUT.t65 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3304 a_85089_n34390# a_83153_n35156.t13 VDD.t4759 VDD.t1710 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3305 VSS.t2117 VSS.t2116 VSS.t2117 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3306 a_50629_n16009.t1 a_51711_n12421.t0 a_83725_7563# VSS.t300 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3307 a_52635_48695.t128 a_52635_34067.t154 VDD.t4894 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3308 a_32913_n8930.t0 a_31953_n19727.t221 a_32353_n8930# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3309 VSS.t2115 VSS.t2114 VSS.t2115 VSS.t620 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3310 VDD.t2796 VDD.t2795 VDD.t2796 VDD.t2402 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3311 VSS.t2113 VSS.t2112 VSS.t2113 VSS.t1258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3312 VDD.t2794 VDD.t2793 VDD.t2794 VDD.t1442 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3313 a_33249_48695.t245 a_31699_20742.t157 VDD.t182 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3314 VDD.t2792 VDD.t2791 VDD.t2792 VDD.t1102 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3315 VDD.t2790 VDD.t2789 VDD.t2790 VDD.t549 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3316 a_65117_n12421# a_50751_n19729.t211 a_64243_n16009.t0 VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3317 a_45138_24920# a_35922_19591.t99 a_44608_24195# VDD.t404 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X3318 a_110225_n6055# a_71281_n8397.t214 a_109695_n5150# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3319 a_85089_10448# a_83153_10448.t19 VDD.t4797 VDD.t1445 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3320 VDD.t2788 VDD.t2787 VDD.t2788 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3321 VSS.t2111 VSS.t2110 VSS.t2111 VSS.t536 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3322 VDD.t2786 VDD.t2785 VDD.t2786 VDD.t928 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3323 a_63683_n2653# a_50751_n19729.t212 a_63161_n2653# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3324 VSS.t2109 VSS.t2108 VSS.t2109 VSS.t1311 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3325 a_96818_7563# a_94892_4481.t17 VSS.t3646 VSS.t1308 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3326 VSS.t2107 VSS.t2106 VSS.t2107 VSS.t889 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3327 VSS.t2105 VSS.t2104 VSS.t2105 VSS.t581 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3328 a_33249_34067.t62 a_33379_34007.t48 a_33249_48695.t4 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3329 VDD.t2784 VDD.t2783 VDD.t2784 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3330 a_59411_n13318# a_50751_n19729.t213 a_58851_n12421# VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3331 VDD.t2782 VDD.t2781 VDD.t2782 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3332 VDD.t2780 VDD.t2778 VDD.t2780 VDD.t2779 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3333 VDD.t2777 VDD.t2775 VDD.t2777 VDD.t2776 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3334 VSS.t2103 VSS.t2102 VSS.t2103 VSS.t609 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3335 VDD.t2774 VDD.t2773 VDD.t2774 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3336 VSS.t2101 VSS.t2100 VSS.t2101 VSS.t1249 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X3337 VSS.t2099 VSS.t2098 VSS.t2099 VSS.t99 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3338 a_65677_n2653# a_50751_n19729.t214 a_65117_n2653# VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3339 VDD.t2772 VDD.t2771 VDD.t2772 VDD.t401 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X3340 VSS.t2097 VSS.t2096 VSS.t2097 VSS.t412 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3341 a_48951_4481.t1 a_47991_5507.t0 a_48391_5639# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3342 a_110225_n14095# a_71281_n8397.t215 VDD.t480 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3343 VSS.t2095 VSS.t2094 VSS.t2095 VSS.t1299 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3344 VDD.t2770 VDD.t2769 VDD.t2770 VDD.t1919 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3345 a_79182_n35156# a_71366_n35156.t8 a_78344_n36322.t1 VDD.t2385 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3346 VDD.t2768 VDD.t2767 VDD.t2768 VDD.t2402 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3347 VDD.t2766 VDD.t2765 VDD.t2766 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3348 VSS.t2093 VSS.t2092 VSS.t2093 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3349 a_52635_34067.t40 a_35922_19591.t100 a_52635_48695.t43 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3350 a_71281_n10073.t39 a_71281_n10073.t38 VDD.t348 VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3351 VSS.t2091 VSS.t2090 VSS.t2091 VSS.t503 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3352 a_111063_n2435# a_71281_n8397.t216 a_110225_n2435# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3353 VDD.t2764 VDD.t2763 VDD.t2764 VDD.t73 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3354 VDD.t2762 VDD.t2761 VDD.t2762 VDD.t61 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3355 VDD.t2760 VDD.t2759 VDD.t2760 VDD.t958 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3356 a_79182_12380# a_71366_11614.t7 a_78344_10448.t1 VDD.t575 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3357 a_112199_n8770# a_71281_n8397.t217 a_111631_n8770# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3358 VSS.t2089 VSS.t2088 VSS.t2089 VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3359 VSS.t2087 VSS.t2086 VSS.t2087 VSS.t1292 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3360 OUT.t64 a_35922_19591.t101 a_52635_49681.t43 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3361 VSS.t2085 VSS.t2084 VSS.t2085 VSS.t816 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3362 a_60080_5639# a_59558_4481.t13 a_53829_10388.t2 VSS.t313 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3363 a_33249_35053.t40 a_33379_34917.t42 a_33249_48695.t57 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3364 a_33249_48695.t244 a_31699_20742.t158 VDD.t183 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3365 VSS.t2083 VSS.t2082 VSS.t2083 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3366 a_60845_n2653# a_50751_n19729.t215 a_60285_n1756# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3367 VSS.t2081 VSS.t2080 VSS.t2081 VSS.t777 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3368 a_107230_n36322# a_106830_n36382.t17 VCM.t1 VDD.t1906 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3369 VDD.t2758 VDD.t2757 VDD.t2758 VDD.t913 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3370 a_33249_48695.t5 a_33379_34007.t49 a_33249_34067.t61 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3371 VSS.t2079 VSS.t2078 VSS.t2079 VSS.t328 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3372 a_33249_48695.t243 a_31699_20742.t159 VDD.t184 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3373 VDD.t2756 VDD.t2755 VDD.t2756 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3374 VSS.t2077 VSS.t2076 VSS.t2077 VSS.t596 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3375 VSS.t2075 VSS.t2074 VSS.t2075 VSS.t652 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3376 a_79182_n33224# a_71366_n35156.t9 a_78344_n36322.t2 VDD.t2385 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3377 a_51711_n3550# a_50751_n19729.t216 a_51151_n3550# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3378 VDD.t2754 VDD.t2753 VDD.t2754 VDD.t680 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3379 VDD.t2752 VDD.t2751 VDD.t2752 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3380 a_83725_7563# a_51711_n12421.t0 a_83153_11614.t2 VSS.t299 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3381 VSS.t2073 VSS.t2072 VSS.t2073 VSS.t353 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3382 VSS.t2071 VSS.t2070 VSS.t2071 VSS.t593 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3383 VDD.t2750 VDD.t2749 VDD.t2750 VDD.t677 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3384 a_33379_34007.t2 a_36162_n36382.t13 a_37968_n36322# VDD.t1895 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3385 a_77776_n35156# a_65658_n29313.t1 a_77225_n29181.t9 VDD.t2347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3386 a_32353_n16904# a_31953_n19727.t222 a_31831_n17801# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3387 VDD.t413 a_35922_19591.t102 a_45706_22884# VDD.t406 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X3388 VDD.t2748 VDD.t2747 VDD.t2748 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3389 VSS.t2069 VSS.t2068 VSS.t2069 VSS.t689 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3390 VSS.t2067 VSS.t2066 VSS.t2067 VSS.t797 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3391 a_90245_n3340# a_71281_n10073.t189 a_89407_n3340# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3392 VDD.t2746 VDD.t2745 VDD.t2746 VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3393 VDD.t2744 VDD.t2743 VDD.t2744 VDD.t1084 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3394 a_44363_n16007.t2 a_65658_n29313.t2 a_66058_n27257# VSS.t411 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3395 VDD.t2742 VDD.t2741 VDD.t2742 VDD.t291 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3396 a_33249_34067.t125 a_35502_25545.t63 VSS.t28 VSS.t9 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3397 a_33787_n19595# a_31953_n19727.t223 a_32913_n16007.t1 VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3398 VDD.t2740 VDD.t2739 VDD.t2740 VDD.t1886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3399 VDD.t2738 VDD.t2737 VDD.t2738 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3400 a_33249_35053.t41 a_33379_34917.t43 a_33249_48695.t58 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3401 VDD.t2736 VDD.t2735 VDD.t2736 VDD.t848 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3402 a_35781_n8930# a_31953_n19727.t224 a_35221_n8930# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3403 VSS.t2065 VSS.t2064 VSS.t2065 VSS.t638 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3404 VDD.t2734 VDD.t2733 VDD.t2734 VDD.t839 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3405 VDD.t2732 VDD.t2730 VDD.t2732 VDD.t2731 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3406 VSS.t2063 VSS.t2062 VSS.t2063 VSS.t676 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3407 VSS.t2061 VSS.t2060 VSS.t2061 VSS.t533 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3408 VDD.t2729 VDD.t2728 VDD.t2729 VDD.t938 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3409 VDD.t2727 VDD.t2726 VDD.t2727 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3410 a_77776_n33224# a_65658_n29313.t1 a_77225_n29181.t9 VDD.t2347 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3411 a_52635_49681.t133 a_52635_34067.t155 VDD.t4893 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3412 VSS.t2059 VSS.t2058 VSS.t2059 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3413 VDD.t2725 VDD.t2724 VDD.t2725 VDD.t1655 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3414 VDD.t2723 VDD.t2722 VDD.t2723 VDD.t424 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3415 a_61515_10448# a_53699_11614.t6 a_60677_10448.t3 VDD.t495 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3416 a_52635_49681.t44 a_35922_19591.t103 OUT.t63 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3417 a_113081_n27257# a_112559_n29181.t7 a_112559_n29181.t8 VSS.t415 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3418 VSS.t2057 VSS.t2056 VSS.t2057 VSS.t324 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3419 VDD.t2721 VDD.t2720 VDD.t2721 VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3420 VDD.t2719 VDD.t2718 VDD.t2719 VDD.t394 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3421 a_30152_11614.t0 a_30324_5507.t1 a_32128_4481# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3422 VSS.t2055 VSS.t2054 VSS.t2055 VSS.t387 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3423 VSS.t2053 VSS.t2052 VSS.t2053 VSS.t614 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3424 a_59558_n29181.t1 a_59558_n29181.t0 a_61484_n30339# VSS.t312 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3425 VDD.t2717 VDD.t2716 VDD.t2717 VDD.t826 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3426 a_39179_n6239# a_31953_n19727.t225 a_38619_n6239# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3427 a_33249_48695.t242 a_31699_20742.t160 VDD.t185 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3428 a_52635_48695.t127 a_52635_34067.t156 VDD.t4892 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3429 VDD.t2715 VDD.t2714 VDD.t2715 VDD.t623 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3430 VDD.t2713 VDD.t2712 VDD.t2713 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3431 a_52635_48695.t126 a_52635_34067.t157 VDD.t4891 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3432 VSS.t431 a_36162_n36382.t14 a_36562_n35156# VDD.t2305 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3433 VDD.t2711 VDD.t2710 VDD.t2711 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3434 VDD.t186 a_31699_20742.t161 a_33249_48695.t241 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3435 VDD.t4890 a_52635_34067.t158 a_52635_49681.t132 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3436 a_54019_n7138# a_50751_n19729.t217 a_53497_n8035# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3437 VSS.t342 a_77225_4481.t17 a_77747_5639# VSS.t341 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3438 VDD.t2709 VDD.t2708 VDD.t2709 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3439 a_82573_n21335# a_71281_n10073.t190 a_81735_n21335# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3440 VDD.t2707 VDD.t2706 VDD.t2707 VDD.t938 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3441 VDD.t2705 VDD.t2704 VDD.t2705 VDD.t813 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3442 a_33249_34067.t124 a_35502_25545.t64 VSS.t25 VSS.t24 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3443 a_33249_48695.t6 a_33379_34007.t50 a_33249_34067.t60 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3444 VSS.t2051 VSS.t2050 VSS.t2051 VSS.t330 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3445 VSS.t2049 VSS.t2048 VSS.t2049 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3446 VSS.t2047 VSS.t2046 VSS.t2047 VSS.t367 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3447 a_57417_n17803# a_50751_n19729.t218 a_56895_n17803# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3448 VSS.t2045 VSS.t2044 VSS.t2045 VSS.t617 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3449 a_53675_4481.t2 a_53829_10388.t17 a_54229_10448# VDD.t1408 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3450 a_30152_11614.t7 a_30152_10448.t14 a_32088_10448# VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3451 a_90969_n34390# a_89163_n36382.t14 VSS.t355 VDD.t550 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3452 VSS.t2043 VSS.t2041 VSS.t2043 VSS.t2042 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X3453 VDD.t2703 VDD.t2702 VDD.t2703 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3454 a_45138_24195# a_35922_19591.t104 a_44608_24195# VDD.t404 pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X3455 a_33249_48695.t59 a_33379_34917.t44 a_33249_35053.t42 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3456 VDD.t187 a_31699_20742.t162 a_33249_48695.t240 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3457 VSS.t2040 VSS.t2039 VSS.t2040 VSS.t1258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3458 VDD.t2701 VDD.t2700 VDD.t2701 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3459 a_100235_n19525# a_71281_n8397.t218 a_99667_n19525# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3460 VSS.t2038 VSS.t2037 VSS.t2038 VSS.t643 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3461 VDD.t2699 VDD.t2698 VDD.t2699 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3462 a_36008_n27257.t1 a_36162_n36382.t15 a_36562_n33224# VDD.t2305 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3463 VDD.t4760 a_83153_n35156.t14 a_83683_n36322# VDD.t1852 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3464 VSS.t2036 VSS.t2035 VSS.t2036 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3465 VDD.t2697 VDD.t2696 VDD.t2697 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3466 a_46879_n14213# a_31953_n19727.t226 a_47753_n16007# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3467 a_33249_48695.t7 a_33379_34007.t51 a_33249_34067.t59 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3468 a_75585_n10073# I1N.t8 VSS.t304 VSS.t303 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X3469 VSS.t2034 VSS.t2033 VSS.t2034 VSS.t539 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3470 a_71342_4481.t0 a_65486_11614.t17 a_73268_7563# VSS.t427 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3471 VDD.t4889 a_52635_34067.t159 a_52635_49681.t131 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3472 VDD.t2695 VDD.t2694 VDD.t2695 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3473 VDD.t2693 VDD.t2692 VDD.t2693 VDD.t325 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3474 VDD.t2691 VDD.t2690 VDD.t2691 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3475 VDD.t2689 VDD.t2688 VDD.t2689 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3476 VDD.t2687 VDD.t2686 VDD.t2687 VDD.t2257 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3477 VSS.t2032 VSS.t2031 VSS.t2032 VSS.t103 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3478 VDD.t2685 VDD.t2684 VDD.t2685 VDD.t798 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3479 VDD.t2683 VDD.t2681 VDD.t2683 VDD.t2682 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3480 a_111631_n14095# a_71281_n8397.t219 a_111063_n14095# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3481 VSS.t392 a_77225_n29181.t16 a_77747_n27257# VSS.t390 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3482 OUT.t62 a_35922_19591.t105 a_52635_49681.t45 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3483 a_102796_4481# a_57977_n12421.t0 a_56895_n16009.t0 VSS.t144 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3484 VSS.t2030 VSS.t2029 VSS.t2030 VSS.t984 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3485 VDD.t2680 VDD.t2679 VDD.t2680 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3486 VDD.t295 a_100820_11614.t12 a_108602_5639# VSS.t151 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3487 VSS.t2028 VSS.t2027 VSS.t2028 VSS.t753 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3488 VSS.t2026 VSS.t2025 VSS.t2026 VSS.t281 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3489 a_30324_5507.t1 a_30152_11614.t11 a_36530_5639# VSS.t325 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3490 a_52635_34067.t0 a_35502_24538.t45 a_33249_34067.t8 VSS.t162 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3491 a_52635_48695.t42 a_35922_19591.t106 a_52635_34067.t17 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3492 VSS.t2024 VSS.t2023 VSS.t2024 VSS.t483 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3493 a_52585_n18700# a_50751_n19729.t219 a_52063_n18700# VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3494 a_98829_n19525# a_71281_n8397.t220 a_98299_n19525# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3495 VDD.t2678 VDD.t2677 VDD.t2678 VDD.t1826 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3496 VDD.t2676 VDD.t2675 VDD.t2676 VDD.t2257 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3497 VDD.t2674 VDD.t2673 VDD.t2674 VDD.t1823 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3498 VDD.t2672 VDD.t2671 VDD.t2672 VDD.t35 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3499 VDD.t188 a_31699_20742.t163 a_35502_25545.t13 VDD.t28 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3500 VSS.t2022 VSS.t2021 VSS.t2022 VSS.t450 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3501 VSS.t2020 VSS.t2019 VSS.t2020 VSS.t506 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3502 a_105365_n19525# a_71281_n8397.t221 a_104527_n19525# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3503 a_113110_n36322# a_103997_n8770.t10 a_106830_n36382.t5 VDD.t328 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3504 VDD.t2670 VDD.t2669 VDD.t2670 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3505 VDD.t2668 VDD.t2667 VDD.t2668 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3506 VDD.t2666 VDD.t2665 VDD.t2666 VDD.t331 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3507 VSS.t2018 VSS.t2017 VSS.t2018 VSS.t1227 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3508 a_53829_10388.t0 a_59558_4481.t14 a_61484_6405# VSS.t312 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3509 a_52635_34067.t35 a_35922_19591.t107 a_52635_48695.t41 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3510 VSS.t2016 VSS.t2015 VSS.t2016 VSS.t581 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3511 VSS.t2014 VSS.t2013 VSS.t2014 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3512 VSS.t2012 VSS.t2011 VSS.t2012 VSS.t495 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3513 a_65117_n2653# a_50751_n19729.t220 a_64595_n3550# VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3514 VDD.t2664 VDD.t2663 VDD.t2664 VDD.t1325 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3515 a_33249_35053.t43 a_33379_34917.t45 a_33249_48695.t60 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3516 VDD.t2662 VDD.t2661 VDD.t2662 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3517 a_95105_n18620# a_71281_n10073.t191 a_94537_n18620# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3518 a_33249_34067.t58 a_33379_34007.t52 a_33249_48695.t8 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3519 a_71864_7563# a_65486_11614.t18 a_71342_7563.t0 VSS.t428 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3520 a_66551_n7138# a_50751_n19729.t221 a_66029_n8035# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3521 a_52635_49681.t130 a_52635_34067.t160 VDD.t4888 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3522 a_90245_n18620# a_71281_n10073.t192 a_89407_n18620# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3523 a_33249_48695.t61 a_33379_34917.t46 a_33249_35053.t44 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3524 a_41891_n29181.t1 a_30324_n29313.t2 a_43848_n36322# VDD.t1798 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3525 a_110225_n4245# a_71281_n8397.t222 a_109695_n4245# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3526 VSS.t2010 VSS.t2009 VSS.t2010 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3527 VSS.t2008 VSS.t2007 VSS.t2008 VSS.t620 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3528 a_71281_n10073.t37 a_71281_n10073.t36 VDD.t350 VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3529 a_52635_49681.t46 a_35922_19591.t108 OUT.t61 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3530 a_31831_n5342.t1 a_32913_n8930.t1 a_83725_n30339# VSS.t366 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3531 VDD.t2660 VDD.t2659 VDD.t2660 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3532 VDD.t2658 VDD.t2657 VDD.t2658 VDD.t325 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3533 VDD.t2656 VDD.t2655 VDD.t2656 VDD.t123 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3534 VDD.t2654 VDD.t2653 VDD.t2654 VDD.t1572 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3535 VDD.t2652 VDD.t2651 VDD.t2652 VDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3536 VDD.t481 a_71281_n8397.t223 a_100803_n13190# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3537 VDD.t2650 VDD.t2649 VDD.t2650 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3538 VSS.t47 a_35502_25545.t65 a_33249_34067.t123 VSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3539 VDD.t4781 a_71266_n4019.t0 a_72596_n4019# VDD.t1191 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3540 VDD.t2648 VDD.t2647 VDD.t2648 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3541 VDD.t2646 VDD.t2645 VDD.t2646 VDD.t1782 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3542 VDD.t2644 VDD.t2643 VDD.t2644 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3543 VDD.t2642 VDD.t2641 VDD.t2642 VDD.t330 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3544 VSS.t231 a_50751_n19729.t36 a_50751_n19729.t37 VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3545 a_45445_n19595.t1 a_65486_n36322.t16 a_71864_n29181# VSS.t155 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3546 a_40613_n13316# a_31953_n19727.t227 a_40053_n12419# VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3547 VSS.t2006 VSS.t2005 VSS.t2006 VSS.t1162 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3548 VDD.t2640 VDD.t2639 VDD.t2640 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3549 VSS.t2004 VSS.t2003 VSS.t2004 VSS.t1600 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X3550 a_54579_n7138# a_50751_n19729.t222 a_54019_n6241# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3551 a_108602_5639# a_100820_11614.t13 a_57977_n12421.t0 VSS.t147 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3552 a_36530_5639# a_30152_11614.t12 VDD.t504 VSS.t326 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3553 a_112199_n7865# a_71281_n8397.t224 a_111631_n7865# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3554 a_52635_48695.t40 a_35922_19591.t109 a_52635_34067.t18 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3555 a_88839_n18620# a_71281_n10073.t193 a_88271_n18620# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3556 a_54019_n19597# a_50751_n19729.t223 a_51711_n19597# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3557 a_40053_n13316# a_31953_n19727.t228 a_39531_n14213# VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3558 a_33249_48695.t62 a_33379_34917.t47 a_33249_35053.t45 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3559 a_94537_n6960# a_71281_n10073.t194 a_93969_n6960# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3560 VDD.t4887 a_52635_34067.t161 a_52635_49681.t129 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3561 VDD.t2638 VDD.t2637 VDD.t2638 VDD.t50 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3562 VSS.t2002 VSS.t2001 VSS.t2002 VSS.t104 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3563 VDD.t2636 VDD.t2635 VDD.t2636 VDD.t979 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3564 a_108636_n34390# a_106830_n36382.t18 VSS.t444 VDD.t1542 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3565 a_33249_34067.t122 a_35502_25545.t66 VSS.t39 VSS.t15 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3566 a_43010_n36322.t2 a_30324_n29313.t2 a_42442_n35156# VDD.t2193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3567 VSS.t17 a_35502_25545.t67 a_33249_34067.t121 VSS.t11 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3568 a_52635_48695.t39 a_35922_19591.t110 a_52635_34067.t43 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3569 VDD.t2634 VDD.t2633 VDD.t2634 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3570 a_30724_n29181# a_30324_n29313.t0 a_30152_n35156.t8 VSS.t145 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3571 VSS.t2000 VSS.t1999 VSS.t2000 VSS.t464 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3572 a_60109_13546# a_53699_11614.t7 a_53829_10388.t7 VDD.t492 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3573 VDD.t189 a_31699_20742.t164 a_35502_24538.t11 VDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3574 VSS.t1998 VSS.t1997 VSS.t1998 VSS.t686 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3575 VDD.t2632 VDD.t2631 VDD.t2632 VDD.t723 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3576 a_35221_n8930# a_31953_n19727.t229 VSS.t112 VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3577 a_38619_n15110# a_31953_n19727.t230 a_38097_n15110# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3578 VDD.t2630 VDD.t2629 VDD.t2630 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3579 a_33249_34067.t57 a_33379_34007.t53 a_33249_48695.t9 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3580 VDD.t2628 VDD.t2627 VDD.t2628 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3581 VDD.t2626 VDD.t2625 VDD.t2626 VDD.t710 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3582 VDD.t2624 VDD.t2623 VDD.t2624 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3583 VSS.t1996 VSS.t1995 VSS.t1996 VSS.t738 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3584 VSS.t1994 VSS.t1993 VSS.t1994 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3585 VDD.t482 a_71281_n8397.t225 a_106501_n13190# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3586 VSS.t1992 VSS.t1991 VSS.t1992 VSS.t652 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3587 a_90245_n3340# a_71281_n10073.t195 a_89407_n2435# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3588 VSS.t1990 VSS.t1989 VSS.t1990 VSS.t401 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3589 VDD.t2622 VDD.t2621 VDD.t2622 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3590 VSS.t1988 VSS.t1987 VSS.t1988 VSS.t536 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3591 a_100992_n29313.t0 a_100820_n36322.t15 a_107198_n27257# VSS.t353 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3592 VDD.t2620 VDD.t2619 VDD.t2620 VDD.t1145 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3593 a_102796_n28415# a_100992_n29313.t0 a_38097_n5342.t0 VSS.t383 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3594 VSS.t1986 VSS.t1985 VSS.t1986 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3595 VDD.t2618 VDD.t2617 VDD.t2618 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3596 VDD.t2616 VDD.t2615 VDD.t2616 VDD.t374 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3597 VSS.t1984 VSS.t1983 VSS.t1984 VSS.t533 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3598 a_43010_n36322.t2 a_30324_n29313.t2 a_42442_n33224# VDD.t2193 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3599 VDD.t2614 VDD.t2613 VDD.t2614 VDD.t1749 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3600 a_60109_11614# a_53699_11614.t8 a_53829_10388.t4 VDD.t492 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3601 VDD.t2612 VDD.t2611 VDD.t2612 VDD.t2164 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3602 a_83709_n8770# a_71281_n10073.t196 a_83141_n8770# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3603 VDD.t2610 VDD.t2609 VDD.t2610 VDD.t2159 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3604 VDD.t2608 VDD.t2607 VDD.t2608 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3605 VSS.t230 a_50751_n19729.t34 a_50751_n19729.t35 VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3606 VSS.t1982 VSS.t1981 VSS.t1982 VSS.t1109 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3607 a_52635_34067.t44 a_35922_19591.t111 a_52635_48695.t38 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3608 VSS.t1980 VSS.t1979 VSS.t1980 VSS.t558 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3609 VSS.t1978 VSS.t1977 VSS.t1978 VSS.t410 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3610 a_44885_n8033# a_31953_n19727.t231 a_44363_n8930# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3611 a_33249_35053.t124 a_35502_25545.t68 VSS.t32 VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3612 VDD.t2606 VDD.t2605 VDD.t2606 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3613 VDD.t2604 VDD.t2603 VDD.t2604 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3614 VSS.t1976 VSS.t1975 VSS.t1976 VSS.t638 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3615 VDD.t2602 VDD.t2601 VDD.t2602 VDD.t2146 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3616 a_46879_n8930# a_31953_n19727.t232 a_46319_n8033# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3617 a_85129_4481# a_51711_n12421.t0 a_50629_n16009.t0 VSS.t298 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3618 VSS.t1974 VSS.t1973 VSS.t1974 VSS.t7 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3619 VDD.t2600 VDD.t2599 VDD.t2600 VDD.t1508 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3620 VSS.t1972 VSS.t1971 VSS.t1972 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3621 a_52635_48695.t37 a_35922_19591.t112 a_52635_34067.t21 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3622 VDD.t2598 VDD.t2597 VDD.t2598 VDD.t1265 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3623 VDD.t2596 VDD.t2595 VDD.t2596 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3624 VDD.t2594 VDD.t2593 VDD.t2594 VDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3625 VSS.t1970 VSS.t1969 VSS.t1970 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3626 VDD.t2592 VDD.t2591 VDD.t2592 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3627 a_32913_n8930.t1 a_83153_n36322.t15 a_89531_n29181# VSS.t458 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3628 a_37934_n27257# a_30152_n36322.t15 a_30324_n29313.t0 VSS.t324 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3629 VDD.t2590 VDD.t2589 VDD.t2590 VDD.t2164 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3630 VDD.t2588 VDD.t2587 VDD.t2588 VDD.t2159 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3631 VSS.t1968 VSS.t1967 VSS.t1968 VSS.t704 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3632 VSS.t1966 VSS.t1965 VSS.t1966 VSS.t492 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3633 VDD.t2586 VDD.t2585 VDD.t2586 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3634 a_52635_49681.t47 a_35922_19591.t113 OUT.t60 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3635 VDD.t2584 VDD.t2583 VDD.t2584 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3636 a_37968_n35156# a_36162_n36382.t16 VSS.t432 VDD.t2131 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3637 a_89407_n9675# a_71281_n10073.t197 a_88839_n9675# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3638 VSS.t1964 VSS.t1963 VSS.t1964 VSS.t709 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3639 a_41487_n18698# a_31953_n19727.t233 a_40965_n18698# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3640 a_42047_n7136# a_31953_n19727.t234 a_41487_n7136# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3641 VDD.t2582 VDD.t2581 VDD.t2582 VDD.t2146 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3642 VDD.t2580 VDD.t2579 VDD.t2580 VDD.t1492 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3643 VDD.t2578 VDD.t2577 VDD.t2578 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3644 VSS.t1962 VSS.t1961 VSS.t1962 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3645 VDD.t2576 VDD.t2574 VDD.t2576 VDD.t2575 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3646 VSS.t439 a_36162_10388.t18 a_36562_12380# VDD.t3614 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3647 VSS.t1960 VSS.t1959 VSS.t1960 VSS.t573 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3648 a_77776_13546# a_71366_11614.t8 a_71496_10388.t5 VDD.t2926 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3649 a_55635_13546# a_53829_10388.t18 a_53675_4481.t3 VDD.t2923 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3650 a_48391_n29181# a_47991_n29313.t0 a_47819_n35156.t8 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3651 a_33249_35053.t46 a_33379_34917.t48 a_33249_48695.t63 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3652 VDD.t2573 VDD.t2571 VDD.t2573 VDD.t2572 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3653 a_71281_n8397.t25 a_71281_n8397.t24 VDD.t440 VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3654 a_83153_n35156.t1 a_83153_n35156.t0 a_85089_n34390# VDD.t1489 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3655 VSS.t1958 VSS.t1957 VSS.t1958 VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3656 VSS.t1956 VSS.t1955 VSS.t1956 VSS.t617 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3657 a_33249_35053.t47 a_33379_34917.t49 a_33249_48695.t64 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3658 VDD.t2570 VDD.t2569 VDD.t2570 VDD.t1716 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3659 a_33249_35053.t103 a_35502_24538.t46 OUT.t10 VSS.t162 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3660 VDD.t2568 VDD.t2567 VDD.t2568 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3661 VSS.t1954 VSS.t1953 VSS.t1954 VSS.t1131 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3662 VSS.t1952 VSS.t1951 VSS.t1952 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3663 a_52635_49681.t128 a_52635_34067.t162 VDD.t4886 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3664 a_37968_n33224# a_36162_n36382.t17 a_36008_n30339.t0 VDD.t2131 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3665 a_51711_n3550# a_50751_n19729.t224 a_51151_n2653# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3666 a_33249_34067.t56 a_33379_34007.t54 a_33249_48695.t10 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3667 a_85089_n36322# a_83153_n35156.t15 VDD.t4761 VDD.t1710 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3668 VDD.t2566 VDD.t2565 VDD.t2566 VDD.t63 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3669 VDD.t33 a_31699_20742.t21 a_31699_20742.t22 VDD.t28 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3670 a_52635_49681.t127 a_52635_34067.t163 VDD.t4885 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3671 VDD.t2564 VDD.t2563 VDD.t2564 VDD.t1484 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3672 VSS.t1950 VSS.t1949 VSS.t1950 VSS.t328 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3673 a_87433_n6960# a_71281_n10073.t198 a_86903_n7865# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3674 VDD.t190 a_31699_20742.t165 a_33249_48695.t239 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3675 a_107198_7563# a_100820_11614.t14 a_106676_7563.t0 VSS.t150 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3676 VSS.t1948 VSS.t1947 VSS.t1948 VSS.t655 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3677 a_77776_11614# a_71366_11614.t9 a_71496_10388.t6 VDD.t2926 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3678 a_55635_11614# a_53829_10388.t19 VSS.t434 VDD.t2923 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3679 a_52635_34067.t44 a_35922_19591.t114 a_52635_48695.t36 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3680 VDD.t2562 VDD.t2560 VDD.t2562 VDD.t2561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3681 VDD.t2559 VDD.t2558 VDD.t2559 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3682 VDD.t2557 VDD.t2556 VDD.t2557 VDD.t79 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3683 VSS.t1946 VSS.t1945 VSS.t1946 VSS.t1116 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3684 a_44885_n18698# a_31953_n19727.t235 a_44363_n19595# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3685 VDD.t191 a_31699_20742.t166 a_33249_48695.t238 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3686 VDD.t2555 VDD.t2554 VDD.t2555 VDD.t634 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3687 VDD.t2553 VDD.t2552 VDD.t2553 VDD.t2103 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3688 a_47819_11614.t3 a_47819_10448.t15 a_49755_10448# VDD.t496 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3689 VDD.t2551 VDD.t2550 VDD.t2551 VDD.t901 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3690 VDD.t2549 VDD.t2548 VDD.t2549 VDD.t626 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3691 VSS.t1944 VSS.t1943 VSS.t1944 VSS.t1543 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3692 a_71496_n36382.t6 a_71366_n35156.t10 a_79182_n35156# VDD.t2100 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3693 a_45445_n16007.t1 a_31953_n19727.t236 a_44885_n16007# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3694 a_95105_n8770# a_71281_n10073.t199 a_94537_n8770# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3695 VDD.t2547 VDD.t2546 VDD.t2547 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3696 VSS.t1942 VSS.t1941 VSS.t1942 VSS.t655 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3697 a_90935_n28415# a_83153_n36322.t16 a_32913_n8930.t1 VSS.t457 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3698 a_53145_n17803# a_50751_n19729.t225 a_52585_n17803# VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3699 VDD.t2545 VDD.t2544 VDD.t2545 VDD.t492 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3700 a_114516_n34390# a_100992_n29313.t2 a_106809_n5150.t2 VDD.t329 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3701 VDD.t2543 VDD.t2542 VDD.t2543 VDD.t1660 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3702 VSS.t452 a_94892_n29181.t15 a_95414_n27257# VSS.t450 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3703 a_33249_48695.t65 a_33379_34917.t50 a_33249_35053.t48 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3704 VDD.t2541 VDD.t2540 VDD.t2541 VDD.t1209 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3705 VDD.t2539 VDD.t2538 VDD.t2539 VDD.t607 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3706 a_71281_n10073.t35 a_71281_n10073.t34 VDD.t355 VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3707 a_66551_n16009# a_50751_n19729.t226 a_65677_n14215# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3708 a_39179_n5342.t1 a_31953_n19727.t237 a_38619_n5342# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3709 VDD.t2537 VDD.t2536 VDD.t2537 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3710 VSS.t1940 VSS.t1939 VSS.t1940 VSS.t646 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3711 VDD.t2535 VDD.t2534 VDD.t2535 VDD.t2103 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3712 a_90245_n17715# a_71281_n10073.t200 a_89715_n17715.t5 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3713 a_52585_n1756# a_50751_n19729.t227 a_51711_n5344.t0 VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3714 VDD.t483 a_71281_n8397.t226 a_106501_n1530# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3715 VSS.t1938 VSS.t1937 VSS.t1938 VSS.t52 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3716 VDD.t2533 VDD.t2532 VDD.t2533 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3717 VDD.t2531 VDD.t2530 VDD.t2531 VDD.t296 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3718 a_54019_n6241# a_50751_n19729.t228 a_53497_n6241# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3719 VDD.t2529 VDD.t2528 VDD.t2529 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3720 VSS.t1936 VSS.t1935 VSS.t1936 VSS.t581 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3721 a_71496_n36382.t7 a_71366_n35156.t11 a_79182_n33224# VDD.t2100 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3722 a_32353_n4445# a_31953_n19727.t238 a_31831_n4445# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3723 VDD.t192 a_31699_20742.t167 a_33249_48695.t237 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3724 a_54579_n2653# a_50751_n19729.t229 a_54019_n1756# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3725 VDD.t2527 VDD.t2526 VDD.t2527 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3726 a_33249_35053.t49 a_33379_34917.t51 a_33249_48695.t66 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3727 a_33249_48695.t236 a_31699_20742.t168 VDD.t193 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3728 a_47819_11614.t5 a_47991_5507.t0 a_49795_6405# VSS.t282 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3729 VSS.t1934 VSS.t1933 VSS.t1934 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3730 a_31953_n19727.t39 a_31953_n19727.t38 VSS.t77 VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3731 VSS.t1932 VSS.t1931 VSS.t1932 VSS.t398 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3732 a_33249_34067.t120 a_35502_25545.t69 VSS.t42 VSS.t24 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3733 VDD.t194 a_31699_20742.t169 a_33249_48695.t235 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3734 VDD.t2525 VDD.t2524 VDD.t2525 VDD.t548 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3735 VDD.t2523 VDD.t2522 VDD.t2523 VDD.t544 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3736 VDD.t2521 VDD.t2520 VDD.t2521 VDD.t503 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3737 VSS.t1930 VSS.t1929 VSS.t1930 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3738 VSS.t1928 VSS.t1927 VSS.t1928 VSS.t910 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3739 VDD.t2519 VDD.t2518 VDD.t2519 VDD.t2082 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3740 VDD.t4884 a_52635_34067.t164 a_52635_49681.t126 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3741 VSS.t1926 VSS.t1925 VSS.t1926 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3742 VDD.t2517 VDD.t2516 VDD.t2517 VDD.t2079 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3743 VSS.t1924 VSS.t1923 VSS.t1924 VSS.t469 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3744 VSS.t1922 VSS.t1921 VSS.t1922 VSS.t329 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3745 VDD.t377 a_71281_n10073.t32 a_71281_n10073.t33 VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3746 VSS.t1920 VSS.t1919 VSS.t1920 VSS.t287 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3747 VSS.t1918 VSS.t1917 VSS.t1918 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3748 VSS.t1916 VSS.t1915 VSS.t1916 VSS.t153 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3749 a_46319_n19595# a_31953_n19727.t239 a_45445_n16007.t0 VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3750 a_52635_48695.t35 a_35922_19591.t115 a_52635_34067.t45 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3751 a_73268_4481# a_65486_11614.t19 a_65658_4421.t0 VSS.t426 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3752 VDD.t2515 VDD.t2514 VDD.t2515 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3753 VSS.t1914 VSS.t1913 VSS.t1914 VSS.t37 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X3754 VDD.t2513 VDD.t2512 VDD.t2513 VDD.t1427 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3755 VDD.t2511 VDD.t2510 VDD.t2511 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3756 OUT.t59 a_35922_19591.t116 a_52635_49681.t48 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3757 VSS.t1912 VSS.t1911 VSS.t1912 VSS.t103 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3758 a_33249_34067.t7 a_35502_24538.t47 a_52635_34067.t61 VSS.t159 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3759 VDD.t2509 VDD.t2508 VDD.t2509 VDD.t424 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3760 a_31953_n19727.t72 a_71266_n4019.t0 a_75602_n3060# VDD.t1667 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3761 a_33249_35053.t50 a_33379_34917.t52 a_33249_48695.t67 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3762 VDD.t2507 VDD.t2506 VDD.t2507 VDD.t845 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3763 VSS.t1910 VSS.t1909 VSS.t1910 VSS.t335 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3764 VDD.t2505 VDD.t2504 VDD.t2505 VDD.t2082 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3765 VDD.t2503 VDD.t2502 VDD.t2503 VDD.t1655 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3766 VDD.t2501 VDD.t2500 VDD.t2501 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3767 a_65486_11614.t0 a_65486_10448.t16 a_67422_10448# VDD.t1381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3768 VDD.t2499 VDD.t2498 VDD.t2499 VDD.t831 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3769 VDD.t2497 VDD.t2496 VDD.t2497 VDD.t2079 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3770 VSS.t1908 VSS.t1907 VSS.t1908 VSS.t146 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3771 VDD.t2495 VDD.t2494 VDD.t2495 VDD.t801 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3772 VSS.t1906 VSS.t1905 VSS.t1906 VSS.t58 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3773 a_52635_49681.t125 a_52635_34067.t165 VDD.t4883 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3774 a_43848_n35156# a_36032_n35156.t7 a_43010_n36322.t1 VDD.t2064 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3775 a_52635_48695.t125 a_52635_34067.t166 VDD.t4882 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3776 VSS.t1904 VSS.t1903 VSS.t1904 VSS.t800 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3777 a_54197_n28415# a_47819_n36322.t15 VDD.t521 VSS.t329 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3778 VDD.t2493 VDD.t2492 VDD.t2493 VDD.t1411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3779 a_44885_n3548# a_31953_n19727.t240 a_44363_n4445# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3780 VDD.t195 a_31699_20742.t170 a_33249_48695.t234 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3781 a_48391_6405# a_47991_4421.t0 a_47819_10448.t1 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3782 VSS.t1902 VSS.t1901 VSS.t1902 VSS.t901 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3783 a_52635_48695.t124 a_52635_34067.t167 VDD.t4881 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3784 VSS.t1900 VSS.t1899 VSS.t1900 VSS.t1082 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X3785 a_46319_n8033# a_31953_n19727.t241 a_45797_n8033# VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3786 VDD.t2491 VDD.t2490 VDD.t2491 VDD.t1644 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3787 a_33249_48695.t233 a_31699_20742.t171 VDD.t196 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3788 a_95105_n21335# a_71281_n10073.t201 a_94537_n21335# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3789 VSS.t1898 VSS.t1897 VSS.t1898 VSS.t514 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3790 VDD.t4880 a_52635_34067.t168 a_52635_49681.t124 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3791 a_89033_n35156.t4 a_89163_n36382.t15 a_90969_n34390# VDD.t551 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3792 a_57417_n7138# a_50751_n19729.t230 a_56895_n7138# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3793 a_46879_n3548# a_31953_n19727.t242 a_46319_n3548# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3794 VSS.t1896 VSS.t1895 VSS.t1896 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3795 VSS.t1894 VSS.t1893 VSS.t1894 VSS.t134 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3796 a_47753_n12419# a_31953_n19727.t243 a_45445_n12419# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3797 VDD.t380 a_71281_n10073.t202 a_89407_n21335# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3798 a_83709_n7865# a_71281_n10073.t203 a_83141_n7865# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3799 VSS.t1892 VSS.t1891 VSS.t1892 VSS.t256 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3800 VDD.t2489 VDD.t2487 VDD.t2489 VDD.t2488 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3801 VDD.t2486 VDD.t2485 VDD.t2486 VDD.t801 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3802 VDD.t2484 VDD.t2483 VDD.t2484 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3803 a_51151_n16009# a_50751_n19729.t231 a_50629_n16009.t2 VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3804 a_43848_n33224# a_36032_n35156.t8 a_43010_n36322.t2 VDD.t2064 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3805 VDD.t2482 VDD.t2481 VDD.t2482 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3806 VSS.t1890 VSS.t1889 VSS.t1890 VSS.t533 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3807 a_77747_n29181# a_77225_n29181.t0 a_77225_n29181.t1 VSS.t385 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3808 a_90969_n36322# a_89163_n36382.t16 a_89009_n27257.t1 VDD.t550 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3809 a_111631_n6960# a_71281_n8397.t227 a_111063_n6960# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3810 a_33249_35053.t51 a_33379_34917.t53 a_33249_48695.t68 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3811 VSS.t1888 VSS.t1887 VSS.t1888 VSS.t209 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3812 a_66551_n6241# a_50751_n19729.t232 a_66029_n6241# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3813 VDD.t2480 VDD.t2479 VDD.t2480 VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3814 VDD.t197 a_31699_20742.t172 a_35502_25545.t14 VDD.t17 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3815 VDD.t343 a_71281_n10073.t30 a_71281_n10073.t31 VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3816 VDD.t2478 VDD.t2477 VDD.t2478 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3817 VDD.t2476 VDD.t2475 VDD.t2476 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3818 VDD.t4879 a_52635_34067.t169 a_52635_49681.t123 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3819 VDD.t2474 VDD.t2473 VDD.t2474 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3820 a_108602_n28415# a_100820_n36322.t16 a_39179_n8930.t1 VSS.t351 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3821 VSS.t1886 VSS.t1885 VSS.t1886 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3822 VDD.t2472 VDD.t2471 VDD.t2472 VDD.t1716 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3823 a_52635_49681.t49 a_35922_19591.t117 OUT.t58 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3824 a_83709_n15000# a_71281_n10073.t204 a_83141_n15000# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3825 VDD.t4780 a_71266_n4019.t0 a_72596_n4978# VDD.t1191 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3826 VDD.t2470 VDD.t2469 VDD.t2470 VDD.t322 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3827 VSS.t1884 VSS.t1883 VSS.t1884 VSS.t889 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3828 VDD.t2468 VDD.t2466 VDD.t2468 VDD.t2467 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3829 VDD.t198 a_31699_20742.t173 a_33249_48695.t232 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3830 VDD.t2465 VDD.t2464 VDD.t2465 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3831 a_59411_n8932# a_50751_n19729.t233 a_58851_n8035# VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3832 VDD.t2463 VDD.t2462 VDD.t2463 VDD.t73 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3833 a_66016_13546# a_65486_10448.t17 a_65486_11614.t1 VDD.t2264 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3834 VDD.t2461 VDD.t2460 VDD.t2461 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3835 VDD.t2459 VDD.t2458 VDD.t2459 VDD.t783 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3836 VSS.t1882 VSS.t1881 VSS.t1882 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3837 a_33249_34067.t55 a_33379_34007.t55 a_33249_48695.t11 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3838 VDD.t2457 VDD.t2456 VDD.t2457 VDD.t795 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3839 VDD.t2455 VDD.t2454 VDD.t2455 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3840 a_31953_n19727.t37 a_31953_n19727.t36 VSS.t76 VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3841 a_67111_n15112# a_50751_n19729.t234 a_66551_n14215# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3842 a_88839_n21335# a_71281_n10073.t205 a_88271_n21335# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3843 VSS.t1880 VSS.t1879 VSS.t1880 VSS.t503 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3844 VSS.t1878 VSS.t1877 VSS.t1878 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3845 VDD.t199 a_31699_20742.t174 a_33249_48695.t231 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3846 VDD.t4878 a_52635_34067.t170 a_52635_49681.t122 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3847 a_65117_n18700# a_50751_n19729.t235 a_64595_n18700# VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3848 VDD.t2453 VDD.t2452 VDD.t2453 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3849 VSS.t3647 a_94892_4481.t18 a_95414_7563# VSS.t1042 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3850 a_33249_48695.t230 a_31699_20742.t175 VDD.t200 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3851 VSS.t1876 VSS.t1875 VSS.t1876 VSS.t1039 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3852 VSS.t1874 VSS.t1873 VSS.t1874 VSS.t160 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3853 VSS.t1872 VSS.t1871 VSS.t1872 VSS.t614 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3854 VDD.t2451 VDD.t2449 VDD.t2451 VDD.t2450 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3855 a_100803_n8770# a_71281_n8397.t228 a_100235_n8770# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3856 a_33249_34067.t119 a_35502_25545.t70 VSS.t51 VSS.t22 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3857 a_105933_n19525# a_71281_n8397.t229 a_105365_n19525# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3858 a_105365_n4245# a_71281_n8397.t230 a_104527_n4245# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3859 VDD.t2448 VDD.t2447 VDD.t2448 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3860 VDD.t2446 VDD.t2445 VDD.t2446 VDD.t783 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3861 VDD.t2444 VDD.t2443 VDD.t2444 VDD.t858 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3862 a_66016_11614# a_65486_10448.t18 a_65486_11614.t2 VDD.t2264 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3863 VDD.t2442 VDD.t2441 VDD.t2442 VDD.t21 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3864 a_59411_n19597# a_50751_n19729.t236 a_58851_n18700# VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3865 a_42047_n17801# a_31953_n19727.t244 a_41487_n17801# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3866 VSS.t1870 VSS.t1869 VSS.t1870 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3867 VSS.t1868 VSS.t1867 VSS.t1868 VSS.t281 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3868 VDD.t2440 VDD.t2439 VDD.t2440 VDD.t545 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3869 a_30152_n35156.t10 a_30324_n29313.t0 a_32128_n30339# VSS.t149 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3870 a_38619_n14213# a_31953_n19727.t245 a_38097_n15110# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3871 VSS.t1866 VSS.t1865 VSS.t1866 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3872 VSS.t1864 VSS.t1863 VSS.t1864 VSS.t1030 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3873 VDD.t2438 VDD.t2437 VDD.t2438 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3874 VDD.t2436 VDD.t2435 VDD.t2436 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3875 a_35922_19591.t3 a_35502_25545.t71 VSS.t3 VSS.t2 nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X3876 VDD.t2434 VDD.t2433 VDD.t2434 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3877 a_93131_n17715# a_71281_n10073.t206 a_92601_n16810# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3878 VDD.t2432 VDD.t2431 VDD.t2432 VDD.t1667 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X3879 VDD.t2430 VDD.t2429 VDD.t2430 VDD.t572 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X3880 VDD.t2428 VDD.t2427 VDD.t2428 VDD.t65 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3881 VSS.t1862 VSS.t1861 VSS.t1862 VSS.t1472 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3882 VSS.t1860 VSS.t1859 VSS.t1860 VSS.t18 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3883 VDD.t341 a_71281_n10073.t28 a_71281_n10073.t29 VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3884 VSS.t424 a_112559_n29181.t19 a_113081_n30339# VSS.t416 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3885 a_93131_n15000# a_71281_n10073.t207 a_92601_n15905# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3886 VSS.t1858 VSS.t1857 VSS.t1858 VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3887 VDD.t2426 VDD.t2424 VDD.t2426 VDD.t2425 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3888 VDD.t201 a_31699_20742.t176 a_33249_48695.t229 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3889 VDD.t2423 VDD.t2422 VDD.t2423 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3890 a_88271_n15000# a_71281_n10073.t208 a_87433_n15000# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3891 VDD.t2421 VDD.t2420 VDD.t2421 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3892 a_31699_19142# I1U.t4 a_30377_19942# VSS.t362 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X3893 a_106501_n9675# a_71281_n8397.t231 a_105933_n9675# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3894 a_83153_n35156.t8 a_83325_n29313.t0 a_85129_n28415# VSS.t365 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3895 a_104527_n19525# a_71281_n8397.t232 a_103997_n19525# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3896 VDD.t2419 VDD.t2418 VDD.t2419 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3897 a_33249_48695.t12 a_33379_34007.t56 a_33249_34067.t54 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3898 a_52635_48695.t34 a_35922_19591.t118 a_52635_34067.t17 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3899 VDD.t2417 VDD.t2416 VDD.t2417 VDD.t1572 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3900 a_32353_n12419# a_31953_n19727.t246 a_31831_n13316# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3901 VSS.t1856 VSS.t1855 VSS.t1856 VSS.t864 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3902 a_95105_n7865# a_71281_n10073.t209 a_94537_n7865# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3903 VSS.t1854 VSS.t1853 VSS.t1854 VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3904 a_54019_n1756# a_50751_n19729.t237 VSS.t266 VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3905 VDD.t4877 a_52635_34067.t171 a_52635_49681.t121 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3906 a_83709_n20430# a_71281_n10073.t210 a_83141_n20430# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3907 a_37968_12380# a_36162_10388.t19 VSS.t440 VDD.t1713 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3908 VDD.t2415 VDD.t2414 VDD.t2415 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3909 a_52635_49681.t120 a_52635_34067.t172 VDD.t4876 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3910 VSS.t1852 VSS.t1851 VSS.t1852 VSS.t500 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3911 a_89407_n18620# a_71281_n10073.t211 a_88839_n18620# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3912 VSS.t1850 VSS.t1849 VSS.t1850 VSS.t542 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3913 VDD.t2413 VDD.t2412 VDD.t2413 VDD.t965 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X3914 a_83683_13546# a_83153_10448.t20 a_83153_11614.t6 VDD.t2776 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3915 a_95414_7563# a_94892_4481.t19 a_89163_10388.t2 VSS.t1003 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3916 VSS.t1848 VSS.t1847 VSS.t1848 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3917 VDD.t2411 VDD.t2410 VDD.t2411 VDD.t751 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3918 a_100803_n18620# a_71281_n8397.t233 a_100235_n18620# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3919 VDD.t2409 VDD.t2408 VDD.t2409 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3920 VDD.t2407 VDD.t2406 VDD.t2407 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3921 VDD.t2405 VDD.t2404 VDD.t2405 VDD.t1551 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3922 a_33249_35053.t52 a_33379_34917.t54 a_33249_48695.t69 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3923 VDD.t2403 VDD.t2401 VDD.t2403 VDD.t2402 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3924 VSS.t1846 VSS.t1845 VSS.t1846 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3925 VSS.t1844 VSS.t1843 VSS.t1844 VSS.t483 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3926 VDD.t2400 VDD.t2399 VDD.t2400 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3927 VDD.t2398 VDD.t2397 VDD.t2398 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3928 a_108636_n36322# a_106830_n36382.t19 a_106676_n27257.t3 VDD.t1542 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3929 VDD.t2396 VDD.t2395 VDD.t2396 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3930 VSS.t1842 VSS.t1841 VSS.t1842 VSS.t593 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3931 VDD.t2394 VDD.t2393 VDD.t2394 VDD.t1102 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3932 VDD.t2392 VDD.t2391 VDD.t2392 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3933 VDD.t2390 VDD.t2389 VDD.t2390 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3934 a_72596_n4019# a_71266_n4019.t0 a_71266_n4019.t0 VDD.t997 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X3935 VDD.t2388 VDD.t2387 VDD.t2388 VDD.t728 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3936 VSS.t1840 VSS.t1839 VSS.t1840 VSS.t704 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3937 a_52635_49681.t50 a_35922_19591.t119 OUT.t57 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3938 a_42413_n28415# a_41891_n29181.t19 a_36162_n36382.t4 VSS.t177 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3939 a_41891_n29181.t8 a_41891_n29181.t7 a_43817_n30339# VSS.t181 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3940 a_37934_6405# a_30152_11614.t13 a_30324_5507.t1 VSS.t324 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3941 a_83683_11614# a_83153_10448.t21 a_83153_11614.t7 VDD.t2776 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3942 a_52635_34067.t37 a_35922_19591.t120 a_52635_48695.t33 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3943 VSS.t1838 VSS.t1837 VSS.t1838 VSS.t1432 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3944 a_106830_n36382.t0 a_112559_n29181.t20 a_114485_n29181# VSS.t414 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3945 VSS.t1836 VSS.t1835 VSS.t1836 VSS.t873 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3946 a_52635_48695.t123 a_52635_34067.t173 VDD.t4875 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3947 a_33249_34067.t53 a_33379_34007.t57 a_33249_48695.t13 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3948 a_39179_n18698# a_31953_n19727.t247 a_38619_n17801# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3949 a_33249_48695.t228 a_31699_20742.t177 VDD.t202 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3950 VDD.t2386 VDD.t2384 VDD.t2386 VDD.t2385 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3951 a_60845_n17803# a_50751_n19729.t238 a_60285_n16906# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3952 a_32913_n8033# a_31953_n19727.t248 a_32353_n8033# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3953 a_33249_48695.t227 a_31699_20742.t178 VDD.t203 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3954 VDD.t2383 VDD.t2382 VDD.t2383 VDD.t680 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3955 VSS.t1834 VSS.t1833 VSS.t1834 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3956 VDD.t2381 VDD.t2380 VDD.t2381 VDD.t498 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3957 VSS.t1832 VSS.t1831 VSS.t1832 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3958 VSS.t1830 VSS.t1829 VSS.t1830 VSS.t1437 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3959 VDD.t2379 VDD.t2378 VDD.t2379 VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3960 a_57417_n13318# a_50751_n19729.t239 a_56895_n13318# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3961 VDD.t2377 VDD.t2376 VDD.t2377 VDD.t677 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3962 VDD.t2375 VDD.t2374 VDD.t2375 VDD.t1919 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3963 a_93131_n20430# a_71281_n10073.t212 VDD.t381 VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3964 VSS.t1828 VSS.t1826 VSS.t1828 VSS.t1827 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X3965 a_33249_48695.t226 a_31699_20742.t179 VDD.t204 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3966 VSS.t1825 VSS.t1824 VSS.t1825 VSS.t910 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3967 VSS.t1823 VSS.t1822 VSS.t1823 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3968 VDD.t2373 VDD.t2372 VDD.t2373 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3969 VSS.t1821 VSS.t1820 VSS.t1821 VSS.t981 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3970 a_88271_n20430# a_71281_n10073.t213 a_87433_n20430# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3971 a_60285_n17803# a_50751_n19729.t240 a_59763_n18700# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3972 VSS.t1819 VSS.t1818 VSS.t1819 VSS.t410 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3973 VDD.t2371 VDD.t2370 VDD.t2371 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3974 VDD.t4774 a_30152_n36322.t16 a_37934_n29181# VSS.t323 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3975 a_94892_n29181.t1 a_94892_n29181.t0 a_96818_n28415# VSS.t445 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3976 a_71864_n27257# a_65486_n36322.t17 a_71342_n27257.t0 VSS.t153 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3977 VDD.t382 a_71281_n10073.t214 a_83709_n9675# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3978 a_46319_n3548# a_31953_n19727.t249 a_45797_n3548# VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3979 VDD.t2369 VDD.t2368 VDD.t2369 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3980 a_33249_48695.t70 a_33379_34917.t55 a_33249_35053.t53 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3981 a_107230_n35156# a_106830_n36382.t20 a_103997_n8770.t4 VDD.t1906 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3982 VDD.t2367 VDD.t2366 VDD.t2367 VDD.t501 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3983 VDD.t2365 VDD.t2364 VDD.t2365 VDD.t1644 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3984 VSS.t1817 VSS.t1816 VSS.t1817 VSS.t738 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3985 VDD.t2363 VDD.t2362 VDD.t2363 VDD.t680 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3986 VDD.t2361 VDD.t2360 VDD.t2361 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3987 VDD.t2359 VDD.t2358 VDD.t2359 VDD.t908 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3988 VDD.t2357 VDD.t2356 VDD.t2357 VDD.t677 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3989 VDD.t2355 VDD.t2354 VDD.t2355 VDD.t1919 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3990 VDD.t2353 VDD.t2351 VDD.t2353 VDD.t2352 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3991 VDD.t2350 VDD.t2349 VDD.t2350 VDD.t1508 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3992 VDD.t2348 VDD.t2346 VDD.t2348 VDD.t2347 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3993 a_66551_n1756# a_50751_n19729.t241 VSS.t267 VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3994 VDD.t2345 VDD.t2344 VDD.t2345 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3995 VDD.t2343 VDD.t2342 VDD.t2343 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3996 a_112199_n1530# a_71281_n8397.t234 a_111631_n1530# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3997 a_33249_34067.t52 a_33379_34007.t58 a_33249_48695.t14 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3998 VSS.t1815 VSS.t1814 VSS.t1815 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3999 a_33249_35053.t54 a_33379_34917.t56 a_33249_48695.t71 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4000 VDD.t2341 VDD.t2340 VDD.t2341 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4001 a_54579_n17803# a_50751_n19729.t242 a_54019_n16906# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4002 VDD.t2339 VDD.t2338 VDD.t2339 VDD.t928 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4003 a_31284_n30339.t1 a_30324_n29313.t1 a_30724_n27257# VSS.t146 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4004 a_36032_n35156.t2 a_36162_n36382.t18 a_37968_n35156# VDD.t1895 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4005 VDD.t2337 VDD.t2336 VDD.t2337 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4006 VDD.t205 a_31699_20742.t180 a_35502_24538.t10 VDD.t41 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4007 a_64243_n16906# a_50751_n19729.t243 a_63683_n16906# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4008 VSS.t1813 VSS.t1812 VSS.t1813 VSS.t842 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4009 VDD.t2335 VDD.t2334 VDD.t2335 VDD.t405 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4010 VDD.t2333 VDD.t2332 VDD.t2333 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4011 a_33787_n7136# a_31953_n19727.t250 a_33265_n8033# VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4012 VDD.t2331 VDD.t2330 VDD.t2331 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4013 VDD.t2329 VDD.t2327 VDD.t2329 VDD.t2328 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4014 a_107230_n33224# a_106830_n36382.t21 a_89033_n36322.t0 VDD.t1906 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4015 a_52635_48695.t32 a_35922_19591.t121 a_52635_34067.t46 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4016 a_48313_n4445# a_31953_n19727.t251 a_47753_n4445# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4017 VDD.t2326 VDD.t2325 VDD.t2326 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4018 VSS.t1811 VSS.t1810 VSS.t1811 VSS.t901 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4019 VSS.t75 a_31953_n19727.t34 a_31953_n19727.t35 VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4020 a_66551_n15112# a_50751_n19729.t244 a_66029_n16906# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4021 a_59411_n3550# a_50751_n19729.t245 a_58851_n3550# VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4022 a_82573_n6960# a_71281_n10073.t215 a_81735_n6960# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4023 VDD.t2324 VDD.t2323 VDD.t2324 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4024 VSS.t306 I1N.t9 a_72603_n8397# VSS.t305 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X4025 a_33249_48695.t225 a_31699_20742.t181 VDD.t206 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4026 VDD.t2322 VDD.t2321 VDD.t2322 VDD.t1886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4027 a_52635_49681.t119 a_52635_34067.t174 VDD.t4874 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4028 VDD.t2320 VDD.t2319 VDD.t2320 VDD.t1492 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4029 a_65677_n19597# a_50751_n19729.t246 a_65117_n19597# VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4030 VDD.t2318 VDD.t2317 VDD.t2318 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4031 a_45445_n8033# a_31953_n19727.t252 a_44885_n7136# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4032 a_114485_4481# a_112559_4481.t21 VSS.t296 VSS.t290 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4033 VSS.t1809 VSS.t1808 VSS.t1809 VSS.t1391 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4034 VDD.t2316 VDD.t2315 VDD.t2316 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4035 a_83709_n15905# a_71281_n10073.t216 a_83141_n15905# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4036 VDD.t2314 VDD.t2313 VDD.t2314 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4037 a_99667_n6960# a_71281_n8397.t235 a_98829_n6960# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4038 a_36032_n36322.t0 a_36162_n36382.t19 a_37968_n33224# VDD.t1895 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4039 a_83153_n35156.t7 a_83153_n35156.t6 a_85089_n36322# VDD.t1489 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4040 VSS.t1807 VSS.t1806 VSS.t1807 VSS.t822 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4041 a_64243_n8035# a_50751_n19729.t247 a_63683_n7138# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4042 VDD.t2312 VDD.t2311 VDD.t2312 VDD.t405 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4043 a_60080_n28415# a_59558_n29181.t18 a_53829_n36382.t3 VSS.t313 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4044 VSS.t1805 VSS.t1804 VSS.t1805 VSS.t52 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4045 VDD.t2310 VDD.t2309 VDD.t2310 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4046 OUT.t56 a_35922_19591.t122 a_52635_49681.t51 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4047 VDD.t2308 VDD.t2307 VDD.t2308 VDD.t913 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4048 a_113037_n20430# a_71281_n8397.t236 a_112199_n19525# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4049 VSS.t1803 VSS.t1802 VSS.t1803 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4050 VDD.t2306 VDD.t2304 VDD.t2306 VDD.t2305 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4051 VSS.t1801 VSS.t1799 VSS.t1801 VSS.t1800 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4052 a_33249_35053.t55 a_33379_34917.t57 a_33249_48695.t72 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4053 a_35781_n8930# a_31953_n19727.t253 a_35221_n8033# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4054 VDD.t2303 VDD.t2301 VDD.t2303 VDD.t2302 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X4055 VDD.t2300 VDD.t2299 VDD.t2300 VDD.t965 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4056 VDD.t2298 VDD.t2297 VDD.t2298 VDD.t1484 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4057 a_31953_n19727.t33 a_31953_n19727.t32 VSS.t74 VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4058 VDD.t2296 VDD.t2295 VDD.t2296 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4059 VDD.t2294 VDD.t2293 VDD.t2294 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4060 VDD.t2292 VDD.t2290 VDD.t2292 VDD.t2291 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4061 a_33249_48695.t123 a_33379_34007.t59 a_33249_34067.t51 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4062 VDD.t2289 VDD.t2288 VDD.t2289 VDD.t1886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4063 a_57977_n16906# a_50751_n19729.t248 a_57417_n16906# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4064 VDD.t207 a_31699_20742.t182 a_33249_48695.t224 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4065 VSS.t1798 VSS.t1797 VSS.t1798 VSS.t889 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4066 a_35221_n19595# a_31953_n19727.t254 VSS.t113 VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4067 a_65658_4421.t0 a_65486_11614.t20 a_71864_7563# VSS.t429 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4068 VDD.t2287 VDD.t2286 VDD.t2287 VDD.t50 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4069 a_52635_49681.t118 a_52635_34067.t175 VDD.t4873 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4070 VDD.t2285 VDD.t2284 VDD.t2285 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4071 VSS.t1796 VSS.t1795 VSS.t1796 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4072 a_33249_48695.t73 a_33379_34917.t58 a_33249_35053.t56 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4073 VDD.t2283 VDD.t2282 VDD.t2283 VDD.t938 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4074 VDD.t4872 a_52635_34067.t176 a_52635_48695.t122 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4075 VDD.t2281 VDD.t2280 VDD.t2281 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4076 VDD.t2279 VDD.t2278 VDD.t2279 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4077 VSS.t1794 VSS.t1793 VSS.t1794 VSS.t480 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4078 VDD.t2277 VDD.t2276 VDD.t2277 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4079 VDD.t2275 VDD.t2274 VDD.t2275 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4080 VSS.t1792 VSS.t1791 VSS.t1792 VSS.t726 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4081 VSS.t1790 VSS.t1789 VSS.t1790 VSS.t942 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4082 a_100803_n7865# a_71281_n8397.t237 a_100235_n7865# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4083 VDD.t2273 VDD.t2272 VDD.t2273 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4084 OUT.t9 a_35502_24538.t48 a_33249_35053.t100 VSS.t163 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4085 VDD.t2271 VDD.t2270 VDD.t2271 VDD.t1254 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4086 VDD.t2269 VDD.t2268 VDD.t2269 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4087 VDD.t4871 a_52635_34067.t177 a_52635_49681.t117 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4088 VDD.t2267 VDD.t2266 VDD.t2267 VDD.t629 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4089 VDD.t2265 VDD.t2263 VDD.t2265 VDD.t2264 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4090 a_39179_n19595.t0 a_47819_n36322.t16 a_54197_n29181# VSS.t327 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4091 VDD.t2262 VDD.t2261 VDD.t2262 VDD.t869 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4092 VDD.t2260 VDD.t2259 VDD.t2260 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4093 a_88839_n8770# a_71281_n10073.t217 a_88271_n8770# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4094 VSS.t1788 VSS.t1787 VSS.t1788 VSS.t813 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4095 VDD.t2258 VDD.t2256 VDD.t2258 VDD.t2257 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4096 VDD.t4762 a_83153_n35156.t16 a_83683_n35156# VDD.t1852 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4097 VDD.t2255 VDD.t2253 VDD.t2255 VDD.t2254 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4098 VDD.t383 a_71281_n10073.t218 a_95105_n9675# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4099 a_114516_n36322# a_100992_n29313.t2 a_106809_n5150.t1 VDD.t329 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4100 OUT.t55 a_35922_19591.t123 a_52635_49681.t52 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4101 VDD.t2252 VDD.t2251 VDD.t2252 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4102 a_93131_n15905# a_71281_n10073.t219 a_92601_n15905# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4103 a_113110_12380# a_100992_4421.t1 a_112559_4481.t1 VDD.t375 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4104 VSS.t1786 VSS.t1785 VSS.t1786 VSS.t692 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4105 a_89407_n3340# a_71281_n10073.t220 a_88839_n3340# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4106 VSS.t1784 VSS.t1783 VSS.t1784 VSS.t207 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4107 a_67462_4481# a_64243_n1756.t1 a_63161_n5344.t2 VSS.t412 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4108 a_88271_n15905# a_71281_n10073.t221 a_87433_n15905# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4109 a_46274_24920# a_35922_19591.t124 a_45706_24920# VDD.t406 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X4110 a_48349_12380# a_47819_10448.t9 a_47819_10448.t10 VDD.t497 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4111 a_44885_n2651# a_31953_n19727.t255 a_44363_n2651# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4112 VSS.t1782 VSS.t1781 VSS.t1782 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4113 a_52635_49681.t53 a_35922_19591.t125 OUT.t54 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4114 VSS.t1780 VSS.t1779 VSS.t1780 VSS.t383 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4115 VDD.t346 a_71281_n10073.t26 a_71281_n10073.t27 VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4116 VDD.t2250 VDD.t2249 VDD.t2250 VDD.t52 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4117 a_33249_35053.t123 a_35502_25545.t72 VSS.t1 VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4118 VDD.t208 a_31699_20742.t183 a_33249_48695.t223 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4119 VDD.t2248 VDD.t2247 VDD.t2248 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4120 a_57417_n6241# a_50751_n19729.t249 a_56895_n7138# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4121 a_46879_n2651# a_31953_n19727.t256 a_46319_n2651# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4122 a_52635_48695.t31 a_35922_19591.t126 a_52635_34067.t47 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4123 a_93969_n15000# a_71281_n10073.t222 a_93131_n15000# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4124 VSS.t1778 VSS.t1777 VSS.t1778 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4125 a_89163_10388.t3 a_94892_4481.t20 a_96818_4481# VSS.t1349 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4126 VSS.t404 a_59558_4481.t15 a_60080_6405# VSS.t316 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4127 VDD.t4763 a_83153_n35156.t17 a_83683_n33224# VDD.t1852 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4128 VSS.t1776 VSS.t1775 VSS.t1776 VSS.t314 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4129 VDD.t357 a_71281_n10073.t24 a_71281_n10073.t25 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4130 VDD.t2246 VDD.t2245 VDD.t2246 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4131 VDD.t2244 VDD.t2242 VDD.t2244 VDD.t2243 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4132 a_33249_35053.t122 a_35502_25545.t73 VSS.t204 VSS.t49 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4133 VDD.t2241 VDD.t2240 VDD.t2241 VDD.t1826 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4134 OUT.t53 a_35922_19591.t127 a_52635_49681.t54 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4135 VSS.t1774 VSS.t1773 VSS.t1774 VSS.t382 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4136 a_83153_11614.t1 a_51711_n12421.t0 a_85129_6405# VSS.t297 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4137 VDD.t2239 VDD.t2238 VDD.t2239 VDD.t1823 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4138 a_51151_n15112# a_50751_n19729.t250 a_50629_n15112# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4139 VSS.t1772 VSS.t1771 VSS.t1772 VSS.t913 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4140 a_33249_34067.t50 a_33379_34007.t60 a_33249_48695.t124 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4141 a_33249_35053.t96 a_35502_24538.t49 OUT.t8 VSS.t159 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4142 a_33249_35053.t57 a_33379_34917.t59 a_33249_48695.t74 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4143 a_71281_n10073.t23 a_71281_n10073.t22 VDD.t344 VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4144 VDD.t2237 VDD.t2236 VDD.t2237 VDD.t2234 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4145 a_52635_48695.t121 a_52635_34067.t178 VDD.t4870 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4146 a_102756_13546# a_100820_10448.t15 VDD.t368 VDD.t325 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4147 VSS.t1770 VSS.t1769 VSS.t1770 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4148 VDD.t2235 VDD.t2233 VDD.t2235 VDD.t2234 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4149 VDD.t2232 VDD.t2231 VDD.t2232 VDD.t552 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4150 a_32913_n18698# a_31953_n19727.t257 a_32353_n18698# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4151 VSS.t1768 VSS.t1767 VSS.t1768 VSS.t209 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4152 a_42047_n2651# a_31953_n19727.t258 a_41487_n1754# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4153 a_113110_n35156# a_100992_n29313.t2 a_112559_n29181.t1 VDD.t328 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4154 VDD.t439 a_71281_n8397.t22 a_71281_n8397.t23 VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4155 VSS.t1766 VSS.t1765 VSS.t1766 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4156 VSS.t1764 VSS.t1763 VSS.t1764 VSS.t1069 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4157 VDD.t2230 VDD.t2229 VDD.t2230 VDD.t680 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4158 VDD.t2228 VDD.t2227 VDD.t2228 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4159 VSS.t1762 VSS.t1761 VSS.t1762 VSS.t768 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4160 VDD.t2226 VDD.t2225 VDD.t2226 VDD.t1826 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4161 VDD.t2224 VDD.t2223 VDD.t2224 VDD.t1427 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4162 a_32913_n3548# a_31953_n19727.t259 a_32353_n3548# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4163 VSS.t1760 VSS.t1759 VSS.t1760 VSS.t780 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4164 VDD.t2222 VDD.t2221 VDD.t2222 VDD.t1823 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4165 a_34347_n14213# a_31953_n19727.t260 a_33787_n14213# VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4166 VSS.t1758 VSS.t1757 VSS.t1758 VSS.t839 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4167 VSS.t1756 VSS.t1755 VSS.t1756 VSS.t873 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4168 VDD.t2220 VDD.t2219 VDD.t2220 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4169 VDD.t2218 VDD.t2217 VDD.t2218 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4170 a_36162_n36382.t1 a_36032_n35156.t9 a_43848_n35156# VDD.t1798 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4171 a_102756_11614# a_100820_10448.t16 VDD.t326 VDD.t325 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4172 a_50629_n16009.t0 a_83325_4421.t2 a_83725_4481# VSS.t300 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4173 VSS.t1754 VSS.t1753 VSS.t1754 VSS.t411 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4174 OUT.t52 a_35922_19591.t128 a_52635_49681.t55 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4175 VDD.t2216 VDD.t2215 VDD.t2216 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4176 VDD.t2214 VDD.t2213 VDD.t2214 VDD.t334 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4177 a_33249_35053.t58 a_33379_34917.t60 a_33249_48695.t75 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4178 a_113110_n33224# a_100992_n29313.t2 a_112559_n29181.t1 VDD.t328 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4179 VDD.t2212 VDD.t2211 VDD.t2212 VDD.t1198 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4180 a_35502_25545.t15 a_31699_20742.t184 VDD.t209 VDD.t17 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4181 VSS.t1752 VSS.t1751 VSS.t1752 VSS.t323 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4182 a_83141_n8770# a_71281_n10073.t223 a_82573_n8770# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4183 VDD.t2210 VDD.t2209 VDD.t2210 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4184 VDD.t2208 VDD.t2207 VDD.t2208 VDD.t1782 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4185 VSS.t1750 VSS.t1749 VSS.t1750 VSS.t1258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4186 VDD.t2206 VDD.t2205 VDD.t2206 VDD.t1411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4187 VSS.t1748 VSS.t1747 VSS.t1748 VSS.t336 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4188 VDD.t2204 VDD.t2203 VDD.t2204 VDD.t390 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4189 a_52635_48695.t30 a_35922_19591.t129 a_52635_34067.t27 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4190 VSS.t1746 VSS.t1745 VSS.t1746 VSS.t489 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4191 a_52635_49681.t56 a_35922_19591.t130 OUT.t51 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4192 VSS.t1744 VSS.t1743 VSS.t1744 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4193 VSS.t30 a_35502_25545.t74 a_33249_34067.t118 VSS.t22 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4194 VDD.t2202 VDD.t2201 VDD.t2202 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4195 a_100235_n8770# a_71281_n8397.t238 a_99667_n8770# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4196 VSS.t1742 VSS.t1741 VSS.t1742 VSS.t352 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4197 a_36162_n36382.t3 a_36032_n35156.t10 a_43848_n33224# VDD.t1798 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4198 VSS.t1740 VSS.t1739 VSS.t1740 VSS.t218 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4199 a_71366_n36322.t1 a_89163_n36382.t17 a_90969_n36322# VDD.t551 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4200 VSS.t1738 VSS.t1737 VSS.t1738 VSS.t1311 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4201 a_96818_4481# a_94892_4481.t21 VSS.t3648 VSS.t1308 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4202 VDD.t4869 a_52635_34067.t179 a_52635_49681.t116 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4203 VSS.t1736 VSS.t1735 VSS.t1736 VSS.t581 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4204 VSS.t1734 VSS.t1733 VSS.t1734 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4205 VDD.t2200 VDD.t2199 VDD.t2200 VDD.t928 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4206 a_54019_n16009# a_50751_n19729.t251 a_53145_n14215# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4207 a_63683_n17803# a_50751_n19729.t252 a_63161_n17803# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4208 VDD.t2198 VDD.t2197 VDD.t2198 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4209 VSS.t1732 VSS.t1731 VSS.t1732 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4210 VDD.t2196 VDD.t2195 VDD.t2196 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4211 VSS.t1730 VSS.t1729 VSS.t1730 VSS.t253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4212 a_93969_n20430# a_71281_n10073.t224 a_93131_n20430# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4213 VDD.t2194 VDD.t2192 VDD.t2194 VDD.t2193 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4214 VDD.t2191 VDD.t2190 VDD.t2191 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4215 VDD.t2189 VDD.t2188 VDD.t2189 VDD.t321 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4216 VDD.t2187 VDD.t2186 VDD.t2187 VDD.t1749 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4217 VSS.t1728 VSS.t1727 VSS.t1728 VSS.t1299 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4218 a_81735_n6055# a_71281_n10073.t225 a_81205_n5150# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4219 a_99667_n18620# a_71281_n8397.t239 a_98829_n18620# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4220 VDD.t2185 VDD.t2184 VDD.t2185 VDD.t1782 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4221 VSS.t1726 VSS.t1725 VSS.t1726 VSS.t1320 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4222 VDD.t2183 VDD.t2182 VDD.t2183 VDD.t1551 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4223 VDD.t2181 VDD.t2180 VDD.t2181 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4224 a_95414_n30339# a_94892_n29181.t16 a_89163_n36382.t5 VSS.t446 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4225 VSS.t1724 VSS.t1723 VSS.t1724 VSS.t1292 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4226 a_38097_n5342.t0 a_39179_n8930.t1 a_101392_n28415# VSS.t384 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4227 a_33249_35053.t59 a_33379_34917.t61 a_33249_48695.t76 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4228 a_72603_n9297# I1N.t10 a_71281_n10073.t0 VSS.t302 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X4229 a_111063_n18620# a_71281_n8397.t240 a_110225_n18620# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4230 a_98829_n6055# a_71281_n8397.t241 a_98299_n5150# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4231 VDD.t2179 VDD.t2178 VDD.t2179 VDD.t2122 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4232 a_89407_n21335# a_71281_n10073.t226 a_88839_n21335# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4233 VSS.t1722 VSS.t1721 VSS.t1722 VSS.t882 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4234 VSS.t1720 VSS.t1719 VSS.t1720 VSS.t148 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4235 VSS.t197 a_35502_25545.t24 a_35502_25545.t25 VSS.t20 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X4236 VDD.t2177 VDD.t2176 VDD.t2177 VDD.t1186 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4237 VDD.t2175 VDD.t2174 VDD.t2175 VDD.t402 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4238 a_31953_n19727.t31 a_31953_n19727.t30 VSS.t73 VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4239 VSS.t1718 VSS.t1717 VSS.t1718 VSS.t457 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4240 a_113037_n8770# a_71281_n8397.t242 a_112199_n8770# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4241 a_52635_49681.t57 a_35922_19591.t131 OUT.t50 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4242 VDD.t2173 VDD.t2172 VDD.t2173 VDD.t913 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4243 a_100803_n21335# a_71281_n8397.t243 a_100235_n21335# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4244 VDD.t2171 VDD.t2170 VDD.t2171 VDD.t1749 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4245 a_46274_23609# a_35922_19591.t132 a_45706_24195# VDD.t406 pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X4246 VSS.t1716 VSS.t1715 VSS.t1716 VSS.t822 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4247 a_100992_4421.t0 a_100820_11614.t15 a_107198_7563# VSS.t188 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4248 VSS.t1714 VSS.t1713 VSS.t1714 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4249 VDD.t2169 VDD.t2168 VDD.t2169 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4250 VDD.t2167 VDD.t2166 VDD.t2167 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4251 a_35221_n8033# a_31953_n19727.t261 a_34699_n8033# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4252 VDD.t2165 VDD.t2163 VDD.t2165 VDD.t2164 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4253 a_83725_4481# a_83325_4421.t2 a_83153_10448.t2 VSS.t299 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4254 a_106501_n19525# a_71281_n8397.t244 a_105933_n19525# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4255 VDD.t2162 VDD.t2161 VDD.t2162 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4256 a_35781_n4445# a_31953_n19727.t262 a_35221_n3548# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4257 a_60109_10448# a_47991_4421.t1 a_59558_4481.t2 VDD.t492 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4258 VDD.t2160 VDD.t2158 VDD.t2160 VDD.t2159 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4259 a_87433_n6055# a_71281_n10073.t227 a_86903_n9675# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4260 VDD.t2157 VDD.t2156 VDD.t2157 VDD.t700 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4261 a_53145_n13318# a_50751_n19729.t253 a_52585_n13318# VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4262 VSS.t1712 VSS.t1711 VSS.t1712 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4263 VDD.t2155 VDD.t2154 VDD.t2155 VDD.t1376 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4264 a_101111_n6055.t1 a_71281_n8397.t245 a_100803_n9675# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4265 a_72596_n4978# a_71266_n4019.t0 a_31953_n19727.t73 VDD.t997 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X4266 VDD.t2153 VDD.t2152 VDD.t2153 VDD.t1373 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4267 VDD.t2151 VDD.t2150 VDD.t2151 VDD.t13 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4268 a_73268_n28415# a_65486_n36322.t18 a_45445_n19595.t1 VSS.t156 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4269 VDD.t2149 VDD.t2148 VDD.t2149 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4270 a_52635_48695.t29 a_35922_19591.t133 a_52635_34067.t27 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4271 VDD.t2147 VDD.t2145 VDD.t2147 VDD.t2146 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4272 VDD.t2144 VDD.t2143 VDD.t2144 VDD.t502 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4273 VDD.t2142 VDD.t2141 VDD.t2142 VDD.t1368 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4274 VSS.t1710 VSS.t1709 VSS.t1710 VSS.t861 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4275 VDD.t2140 VDD.t2139 VDD.t2140 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4276 a_33249_35053.t97 a_35502_24538.t50 OUT.t7 VSS.t166 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4277 VSS.t1708 VSS.t1707 VSS.t1708 VSS.t913 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4278 VSS.t36 a_35502_25545.t75 a_33249_35053.t121 VSS.t35 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4279 a_52635_34067.t64 a_35502_24538.t51 a_33249_34067.t6 VSS.t163 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4280 VSS.t1706 VSS.t1705 VSS.t1706 VSS.t533 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4281 VDD.t2138 VDD.t2137 VDD.t2138 VDD.t1716 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4282 a_83709_n1530# a_71281_n10073.t228 a_83141_n1530# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4283 VDD.t2136 VDD.t2135 VDD.t2136 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4284 VSS.t1704 VSS.t1703 VSS.t1704 VSS.t858 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4285 VDD.t2134 VDD.t2133 VDD.t2134 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4286 a_33249_34067.t49 a_33379_34007.t61 a_33249_48695.t125 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4287 VDD.t2132 VDD.t2130 VDD.t2132 VDD.t2131 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4288 a_63683_n8932# a_50751_n19729.t254 a_63161_n8932# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4289 a_33249_34067.t48 a_33379_34007.t62 a_33249_48695.t126 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4290 a_96818_n29181# a_94892_n29181.t17 VSS.t453 VSS.t447 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4291 VDD.t2129 VDD.t2128 VDD.t2129 VDD.t1357 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4292 a_57417_n12421# a_50751_n19729.t255 a_56895_n13318# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4293 a_42442_12380# a_30324_4421.t1 a_41891_4481.t8 VDD.t291 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4294 a_41487_n15110# a_31953_n19727.t263 a_40965_n16904# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4295 VDD.t2127 VDD.t2126 VDD.t2127 VDD.t896 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4296 a_65677_n8932# a_50751_n19729.t256 a_65117_n8932# VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4297 VDD.t2125 VDD.t2124 VDD.t2125 VDD.t1352 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4298 a_52635_48695.t120 a_52635_34067.t180 VDD.t4868 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4299 VDD.t2123 VDD.t2121 VDD.t2123 VDD.t2122 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4300 a_33249_35053.t60 a_33379_34917.t62 a_33249_48695.t77 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4301 a_52635_48695.t119 a_52635_34067.t181 VDD.t4867 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4302 VDD.t2120 VDD.t2119 VDD.t2120 VDD.t558 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4303 a_35502_24538.t9 a_31699_20742.t185 VDD.t210 VDD.t30 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4304 VSS.t1702 VSS.t1701 VSS.t1702 VSS.t1621 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4305 a_88839_n7865# a_71281_n10073.t229 a_88271_n7865# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4306 VDD.t211 a_31699_20742.t186 a_33249_48695.t222 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4307 VDD.t2118 VDD.t2117 VDD.t2118 VDD.t1716 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4308 a_87433_n17715# a_71281_n10073.t230 a_86903_n16810# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4309 VSS.t1700 VSS.t1699 VSS.t1700 VSS.t489 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4310 a_46319_n2651# a_31953_n19727.t264 a_45797_n3548# VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4311 VSS.t1698 VSS.t1697 VSS.t1698 VSS.t596 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4312 a_52635_49681.t115 a_52635_34067.t182 VDD.t4866 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4313 a_47753_n7136# a_31953_n19727.t265 a_47231_n8033# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4314 a_57417_n1756# a_50751_n19729.t257 a_56895_n2653# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4315 a_93131_n6055# a_71281_n10073.t231 a_92601_n5150# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4316 VSS.t45 a_35502_25545.t76 a_33249_35053.t120 VSS.t44 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4317 a_33249_48695.t221 a_31699_20742.t187 VDD.t212 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4318 a_52635_49681.t114 a_52635_34067.t183 VDD.t4865 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4319 a_87433_n15000# a_71281_n10073.t232 a_86903_n15905# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4320 a_89407_n2435# a_71281_n10073.t233 a_88839_n2435# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4321 VSS.t1696 VSS.t1695 VSS.t1696 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4322 VSS.t1694 VSS.t1693 VSS.t1694 VSS.t159 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4323 VSS.t1692 VSS.t1691 VSS.t1692 VSS.t593 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4324 VDD.t213 a_31699_20742.t188 a_33249_48695.t220 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4325 VSS.t1690 VSS.t1689 VSS.t1690 VSS.t327 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4326 VDD.t2116 VDD.t2115 VDD.t2116 VDD.t1959 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4327 VDD.t2114 VDD.t2113 VDD.t2114 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4328 VSS.t1688 VSS.t1687 VSS.t1688 VSS.t329 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4329 VDD.t2112 VDD.t2111 VDD.t2112 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4330 a_30324_n30399.t1 a_30152_n36322.t17 a_36530_n28415# VSS.t325 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4331 a_85089_n35156# a_83153_n35156.t18 VDD.t4764 VDD.t1710 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4332 VDD.t2110 VDD.t2109 VDD.t2110 VDD.t1130 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4333 a_93969_n15905# a_71281_n10073.t234 a_93131_n15905# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4334 VSS.t1686 VSS.t1685 VSS.t1686 VSS.t676 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4335 VDD.t2108 VDD.t2107 VDD.t2108 VDD.t1660 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4336 VDD.t2106 VDD.t2105 VDD.t2106 VDD.t81 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4337 a_71342_7563.t1 a_65486_11614.t21 a_73268_4481# VSS.t427 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4338 a_55635_10448# a_53829_10388.t20 a_53675_7563.t2 VDD.t2923 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4339 VSS.t1684 VSS.t1683 VSS.t1684 VSS.t1366 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4340 a_77776_10448# a_65658_4421.t2 a_77225_4481.t8 VDD.t2926 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4341 VDD.t2104 VDD.t2102 VDD.t2104 VDD.t2103 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4342 a_44885_n15110# a_31953_n19727.t266 a_44363_n15110# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4343 a_102796_n27257# a_39179_n8930.t1 a_38097_n5342.t1 VSS.t383 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4344 VSS.t1682 VSS.t1681 VSS.t1682 VSS.t1261 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4345 a_59411_n2653# a_50751_n19729.t258 a_58851_n2653# VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4346 VDD.t2101 VDD.t2099 VDD.t2101 VDD.t2100 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4347 a_61484_5639# a_59558_4481.t16 VSS.t405 VSS.t314 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4348 VSS.t1680 VSS.t1679 VSS.t1680 VSS.t768 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4349 a_85089_n33224# a_83153_n35156.t19 VDD.t4765 VDD.t1710 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4350 VSS.t1678 VSS.t1677 VSS.t1678 VSS.t686 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4351 VSS.t1676 VSS.t1675 VSS.t1676 VSS.t542 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4352 VSS.t1674 VSS.t1673 VSS.t1674 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4353 VDD.t2098 VDD.t2097 VDD.t2098 VDD.t493 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4354 a_105933_n8770# a_71281_n8397.t246 a_105365_n8770# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4355 VDD.t2096 VDD.t2095 VDD.t2096 VDD.t1660 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4356 VSS.t1672 VSS.t1671 VSS.t1672 VSS.t351 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4357 a_33249_48695.t219 a_31699_20742.t189 VDD.t214 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4358 a_52635_48695.t118 a_52635_34067.t184 VDD.t4864 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4359 a_64243_n6241# a_50751_n19729.t259 a_63683_n6241# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4360 a_48951_4481.t1 a_47991_4421.t0 a_48391_6405# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4361 VSS.t1670 VSS.t1669 VSS.t1670 VSS.t66 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4362 a_33249_48695.t218 a_31699_20742.t190 VDD.t215 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4363 a_33249_48695.t217 a_31699_20742.t191 VDD.t216 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4364 VDD.t2094 VDD.t2093 VDD.t2094 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4365 VDD.t217 a_31699_20742.t192 a_35502_24538.t8 VDD.t41 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4366 a_106501_n3340# a_71281_n8397.t247 a_105933_n3340# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4367 VDD.t2092 VDD.t2090 VDD.t2092 VDD.t2091 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4368 VDD.t218 a_31699_20742.t193 a_33249_48695.t216 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4369 a_31953_n19727.t29 a_31953_n19727.t28 VSS.t72 VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4370 VSS.t1668 VSS.t1667 VSS.t1668 VSS.t816 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4371 a_60080_6405# a_59558_4481.t3 a_59558_4481.t4 VSS.t313 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4372 VDD.t2089 VDD.t2088 VDD.t2089 VDD.t405 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4373 a_95105_n1530# a_71281_n10073.t235 a_94537_n1530# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4374 VSS.t1666 VSS.t1665 VSS.t1666 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4375 VSS.t1664 VSS.t1663 VSS.t1664 VSS.t149 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4376 VDD.t2087 VDD.t2086 VDD.t2087 VDD.t389 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4377 a_104527_n6055# a_71281_n8397.t248 a_103997_n5150# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4378 VSS.t1662 VSS.t1661 VSS.t1662 VSS.t258 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4379 a_112199_n13190# a_71281_n8397.t249 a_111631_n13190# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4380 a_71864_4481# a_65486_11614.t22 a_71342_4481.t1 VSS.t428 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4381 a_83141_n7865# a_71281_n10073.t236 a_82573_n7865# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4382 VSS.t1660 VSS.t1659 VSS.t1660 VSS.t614 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4383 a_71281_n8397.t21 a_71281_n8397.t20 VDD.t437 VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4384 VDD.t2085 VDD.t2084 VDD.t2085 VDD.t290 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4385 VSS.t1658 VSS.t1657 VSS.t1658 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4386 a_52635_49681.t58 a_35922_19591.t134 OUT.t49 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4387 VDD.t2083 VDD.t2081 VDD.t2083 VDD.t2082 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4388 a_87433_n20430# a_71281_n10073.t237 VDD.t384 VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4389 VSS.t1656 VSS.t1655 VSS.t1656 VSS.t539 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4390 VDD.t2080 VDD.t2078 VDD.t2080 VDD.t2079 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4391 VDD.t2077 VDD.t2076 VDD.t2077 VDD.t65 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4392 VDD.t2075 VDD.t2074 VDD.t2075 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4393 a_100235_n7865# a_71281_n8397.t250 a_99667_n7865# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4394 VDD.t2073 VDD.t2072 VDD.t2073 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4395 VSS.t71 a_31953_n19727.t26 a_31953_n19727.t27 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4396 VSS.t1654 VSS.t1653 VSS.t1654 VSS.t142 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4397 a_52635_48695.t28 a_35922_19591.t135 a_52635_34067.t48 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4398 a_83709_n14095# a_71281_n10073.t238 a_83141_n14095# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4399 VSS.t1652 VSS.t1651 VSS.t1652 VSS.t797 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4400 VSS.t1650 VSS.t1649 VSS.t1650 VSS.t649 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4401 VSS.t70 a_31953_n19727.t24 a_31953_n19727.t25 VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4402 VDD.t2071 VDD.t2070 VDD.t2071 VDD.t1357 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4403 a_40053_n18698# a_31953_n19727.t267 a_39531_n18698# VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4404 a_52635_49681.t113 a_52635_34067.t185 VDD.t4863 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4405 VDD.t2069 VDD.t2068 VDD.t2069 VDD.t1644 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4406 VSS.t1648 VSS.t1647 VSS.t1648 VSS.t536 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4407 VDD.t2067 VDD.t2066 VDD.t2067 VDD.t670 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4408 a_81735_n4245# a_71281_n10073.t239 a_81205_n4245# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4409 VDD.t436 a_71281_n8397.t18 a_71281_n8397.t19 VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4410 VSS.t1646 VSS.t1645 VSS.t1646 VSS.t1162 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4411 VSS.t1644 VSS.t1643 VSS.t1644 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4412 VDD.t4862 a_52635_34067.t186 a_52635_48695.t117 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4413 a_42047_n13316# a_31953_n19727.t268 a_41487_n13316# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4414 VSS.t1642 VSS.t1641 VSS.t1642 VSS.t483 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4415 VDD.t219 a_31699_20742.t194 a_33249_48695.t215 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4416 a_41487_n4445# a_31953_n19727.t269 a_40965_n6239# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4417 a_52635_49681.t112 a_52635_34067.t187 VDD.t4861 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4418 a_35221_n3548# a_31953_n19727.t270 a_34699_n3548# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4419 VSS.t1640 VSS.t1639 VSS.t1640 VSS.t365 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4420 VDD.t2065 VDD.t2063 VDD.t2065 VDD.t2064 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4421 VDD.t2062 VDD.t2060 VDD.t2062 VDD.t2061 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4422 VDD.t2059 VDD.t2058 VDD.t2059 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4423 VDD.t2057 VDD.t2056 VDD.t2057 VDD.t1655 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4424 VDD.t435 a_71281_n8397.t16 a_71281_n8397.t17 VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4425 a_98829_n4245# a_71281_n8397.t251 a_98299_n4245# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4426 VDD.t2055 VDD.t2054 VDD.t2055 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4427 a_52585_n14215# a_50751_n19729.t260 a_52063_n14215# VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4428 a_57977_n8035# a_50751_n19729.t261 a_57417_n7138# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4429 a_67462_n28415# a_65658_n29313.t0 a_44363_n16007.t1 VSS.t412 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4430 VDD.t2053 VDD.t2052 VDD.t2053 VDD.t677 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4431 VSS.t1638 VSS.t1637 VSS.t1638 VSS.t144 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4432 VDD.t2051 VDD.t2050 VDD.t2051 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4433 a_113037_n8770# a_71281_n8397.t252 a_112199_n7865# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4434 a_33249_34067.t47 a_33379_34007.t63 a_33249_48695.t127 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4435 VDD.t2049 VDD.t2048 VDD.t2049 VDD.t1644 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4436 VSS.t1636 VSS.t1635 VSS.t1636 VSS.t278 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4437 VSS.t343 a_77225_4481.t18 a_77747_6405# VSS.t341 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4438 VDD.t2047 VDD.t2045 VDD.t2047 VDD.t2046 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4439 a_95943_n17715# a_71281_n10073.t240 a_95413_n16810.t1 VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4440 VDD.t2044 VDD.t2043 VDD.t2044 VDD.t1102 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4441 a_84547_n3340# a_71281_n10073.t241 a_83709_n3340# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4442 VDD.t2042 VDD.t2041 VDD.t2042 VDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4443 a_33249_34067.t5 a_35502_24538.t52 a_52635_34067.t62 VSS.t166 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4444 VDD.t2040 VDD.t2039 VDD.t2040 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4445 a_33249_35053.t61 a_33379_34917.t63 a_33249_48695.t78 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4446 a_90935_n27257# a_83153_n36322.t17 a_83325_n29313.t0 VSS.t457 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4447 VDD.t2038 VDD.t2037 VDD.t2038 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4448 VDD.t4860 a_52635_34067.t188 a_52635_48695.t116 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4449 a_95943_n15000# a_71281_n10073.t242 a_95105_n15000# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4450 VDD.t2036 VDD.t2035 VDD.t2036 VDD.t1655 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4451 VDD.t2034 VDD.t2033 VDD.t2034 VDD.t639 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4452 VDD.t2032 VDD.t2031 VDD.t2032 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4453 VDD.t2030 VDD.t2029 VDD.t2030 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4454 VDD.t2028 VDD.t2027 VDD.t2028 VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4455 a_93131_n14095# a_71281_n10073.t243 IBPOUT.t0 VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4456 VDD.t2026 VDD.t2025 VDD.t2026 VDD.t801 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4457 a_110225_n18620# a_71281_n8397.t253 a_109695_n19525# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4458 VDD.t2024 VDD.t2022 VDD.t2024 VDD.t2023 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4459 a_32913_n3548# a_31953_n19727.t271 a_32353_n2651# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4460 VDD.t2021 VDD.t2020 VDD.t2021 VDD.t1254 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4461 a_90969_n35156# a_89163_n36382.t18 VSS.t356 VDD.t550 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4462 a_52635_49681.t111 a_52635_34067.t189 VDD.t4859 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4463 a_88271_n14095# a_71281_n10073.t244 a_87433_n14095# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4464 a_33249_48695.t79 a_33379_34917.t64 a_33249_35053.t62 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4465 VDD.t2019 VDD.t2018 VDD.t2019 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4466 VDD.t2017 VDD.t2016 VDD.t2017 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4467 VSS.t1634 VSS.t1633 VSS.t1634 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4468 VDD.t2015 VDD.t2014 VDD.t2015 VDD.t1055 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4469 a_65117_n8932# a_50751_n19729.t262 VSS.t268 VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4470 VSS.t1632 VSS.t1631 VSS.t1632 VSS.t762 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4471 a_59558_4481.t6 a_59558_4481.t5 a_61484_7563# VSS.t312 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4472 VSS.t1630 VSS.t1629 VSS.t1630 VSS.t250 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4473 VDD.t2013 VDD.t2012 VDD.t2013 VDD.t1183 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4474 VDD.t220 a_31699_20742.t195 a_33249_48695.t214 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4475 VSS.t1628 VSS.t1627 VSS.t1628 VSS.t177 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4476 VDD.t4858 a_52635_34067.t190 a_52635_48695.t115 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4477 VDD.t2011 VDD.t2010 VDD.t2011 VDD.t394 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4478 VSS.t1626 VSS.t1625 VSS.t1626 VSS.t689 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4479 a_90969_12380# a_89163_10388.t18 VSS.t360 VDD.t559 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4480 VDD.t2009 VDD.t2008 VDD.t2009 VDD.t26 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4481 VDD.t2007 VDD.t2006 VDD.t2007 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4482 a_65658_n29313.t0 a_65486_n36322.t19 a_71864_n30339# VSS.t155 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4483 VSS.t1624 VSS.t1623 VSS.t1624 VSS.t459 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4484 VDD.t2005 VDD.t2004 VDD.t2005 VDD.t614 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4485 a_71281_n10073.t21 a_71281_n10073.t20 VDD.t353 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4486 VSS.t1622 VSS.t1620 VSS.t1622 VSS.t1621 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4487 VDD.t2003 VDD.t2002 VDD.t2003 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4488 VDD.t4857 a_52635_34067.t191 a_52635_49681.t110 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4489 a_94537_n15000# a_71281_n10073.t245 a_93969_n15000# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4490 VDD.t2001 VDD.t2000 VDD.t2001 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4491 VDD.t1999 VDD.t1997 VDD.t1999 VDD.t1998 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4492 a_90969_n33224# a_89163_n36382.t19 a_89009_n30339.t2 VDD.t550 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4493 VSS.t1619 VSS.t1618 VSS.t1619 VSS.t676 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4494 VDD.t1996 VDD.t1995 VDD.t1996 VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4495 VSS.t1617 VSS.t1616 VSS.t1617 VSS.t252 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4496 VSS.t1615 VSS.t1614 VSS.t1615 VSS.t753 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4497 VDD.t417 a_100820_11614.t16 a_108602_6405# VSS.t151 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4498 a_30324_5507.t1 a_30152_11614.t14 a_36530_6405# VSS.t325 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4499 VSS.t1613 VSS.t1612 VSS.t1613 VSS.t283 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4500 VSS.t1611 VSS.t1610 VSS.t1611 VSS.t445 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4501 VSS.t1609 VSS.t1608 VSS.t1609 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4502 a_54019_n15112# a_50751_n19729.t263 a_53497_n16906# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4503 a_99667_n21335# a_71281_n8397.t254 a_98829_n21335# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4504 a_30724_n30339# a_30324_n30399.t1 a_30152_n36322.t3 VSS.t145 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4505 a_39179_n14213# a_31953_n19727.t272 a_38619_n13316# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4506 a_79151_n28415# a_77225_n29181.t17 VSS.t393 VSS.t387 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4507 a_87433_n15905# a_71281_n10073.t246 a_86903_n15905# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4508 VSS.t1607 VSS.t1606 VSS.t1607 VSS.t614 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4509 VDD.t1994 VDD.t1993 VDD.t1994 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4510 VDD.t1992 VDD.t1991 VDD.t1992 VDD.t389 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4511 VDD.t1990 VDD.t1989 VDD.t1990 VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4512 VDD.t1988 VDD.t1987 VDD.t1988 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4513 VDD.t1986 VDD.t1985 VDD.t1986 VDD.t428 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4514 a_93131_n4245# a_71281_n10073.t247 a_92601_n4245# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4515 a_33249_48695.t213 a_31699_20742.t196 VDD.t221 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4516 a_33787_n1754# a_31953_n19727.t273 VSS.t114 VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4517 VSS.t1605 VSS.t1604 VSS.t1605 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4518 VDD.t1984 VDD.t1983 VDD.t1984 VDD.t783 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4519 a_66016_10448# a_65486_10448.t4 a_65486_10448.t5 VDD.t2264 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4520 a_111063_n21335# a_71281_n8397.t255 a_110225_n21335# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4521 VDD.t1982 VDD.t1981 VDD.t1982 VDD.t304 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4522 VDD.t1980 VDD.t1979 VDD.t1980 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4523 a_35781_n17801# a_31953_n19727.t274 a_35221_n16904# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4524 a_33249_48695.t212 a_31699_20742.t197 VDD.t222 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4525 VSS.t1603 VSS.t1602 VSS.t1603 VSS.t1162 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4526 a_60285_n13318# a_50751_n19729.t264 a_59763_n14215# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4527 VSS.t1601 VSS.t1599 VSS.t1601 VSS.t1600 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X4528 VDD.t1978 VDD.t1977 VDD.t1978 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4529 a_33249_48695.t211 a_31699_20742.t198 VDD.t223 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4530 a_45445_n1754# a_31953_n19727.t275 a_44885_n1754# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4531 VSS.t1598 VSS.t1597 VSS.t1598 VSS.t106 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4532 VDD.t1976 VDD.t1975 VDD.t1976 VDD.t1212 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4533 a_83141_n13190# a_71281_n10073.t248 a_82573_n13190# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4534 a_100803_n1530# a_71281_n8397.t256 a_100235_n1530# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4535 a_83725_n28415# a_32913_n8930.t1 a_83153_n36322.t0 VSS.t367 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4536 a_95943_n20430# a_71281_n10073.t249 a_95105_n20430# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4537 a_52635_48695.t114 a_52635_34067.t192 VDD.t4856 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4538 a_54197_n27257# a_47819_n36322.t17 a_53675_n27257.t1 VSS.t329 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4539 VDD.t1974 VDD.t1973 VDD.t1974 VDD.t1018 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4540 a_64243_n1756.t0 a_50751_n19729.t265 a_63683_n1756# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4541 VSS.t1596 VSS.t1595 VSS.t1596 VSS.t1131 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4542 VSS.t1594 VSS.t1593 VSS.t1594 VSS.t1258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4543 VSS.t1592 VSS.t1591 VSS.t1592 VSS.t643 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4544 VSS.t1590 VSS.t1589 VSS.t1590 VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4545 VDD.t1972 VDD.t1971 VDD.t1972 VDD.t1551 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4546 VDD.t298 a_65486_n36322.t20 a_73268_n29181# VSS.t154 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4547 a_95943_n3340# a_71281_n10073.t250 a_95105_n3340# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4548 a_35781_n2651# a_31953_n19727.t276 a_35221_n2651# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4549 VDD.t1970 VDD.t1969 VDD.t1970 VDD.t920 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4550 VSS.t1588 VSS.t1587 VSS.t1588 VSS.t738 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4551 VDD.t1968 VDD.t1967 VDD.t1968 VDD.t1572 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4552 a_33249_34067.t46 a_33379_34007.t64 a_33249_48695.t128 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4553 VDD.t1966 VDD.t1965 VDD.t1966 VDD.t1198 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4554 a_107198_4481# a_100820_11614.t17 a_106676_4481.t1 VSS.t150 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4555 VDD.t1964 VDD.t1963 VDD.t1964 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4556 a_105933_n7865# a_71281_n8397.t257 a_105365_n7865# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4557 a_53145_n13318# a_50751_n19729.t266 a_52585_n12421# VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4558 VSS.t1586 VSS.t1585 VSS.t1586 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4559 VDD.t1962 VDD.t1961 VDD.t1962 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4560 VSS.t1584 VSS.t1583 VSS.t1584 VSS.t536 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4561 VSS.t1582 VSS.t1581 VSS.t1582 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4562 VDD.t1960 VDD.t1958 VDD.t1960 VDD.t1959 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4563 VDD.t1957 VDD.t1956 VDD.t1957 VDD.t1442 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4564 VDD.t1955 VDD.t1954 VDD.t1955 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4565 VDD.t1953 VDD.t1952 VDD.t1953 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4566 a_52635_48695.t113 a_52635_34067.t193 VDD.t4855 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4567 VSS.t1580 VSS.t1579 VSS.t1580 VSS.t1116 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4568 VSS.t1578 VSS.t1577 VSS.t1578 VSS.t313 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4569 a_81735_n13190# a_71281_n10073.t251 a_81205_n16810# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4570 VDD.t358 a_71281_n10073.t18 a_71281_n10073.t19 VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4571 VDD.t1951 VDD.t1950 VDD.t1951 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4572 a_35502_25545.t16 a_31699_20742.t199 VDD.t224 VDD.t21 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4573 VDD.t1949 VDD.t1948 VDD.t1949 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4574 a_83325_n29313.t0 a_83153_n36322.t18 a_89531_n30339# VSS.t458 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4575 a_106501_n2435# a_71281_n8397.t258 a_105933_n2435# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4576 a_94537_n20430# a_71281_n10073.t252 a_93969_n20430# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4577 a_108602_6405# a_100820_11614.t18 a_57977_n12421.t0 VSS.t147 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4578 a_36530_6405# a_30152_11614.t15 VDD.t505 VSS.t326 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4579 VDD.t1947 VDD.t1946 VDD.t1947 VDD.t1186 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4580 a_52635_48695.t27 a_35922_19591.t136 a_52635_34067.t6 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4581 a_49795_5639# a_47991_4421.t0 a_48951_4481.t1 VSS.t281 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4582 VDD.t1945 VDD.t1944 VDD.t1945 VDD.t1551 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4583 a_32128_n29181# a_30324_n30399.t2 a_31284_n30339.t0 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4584 VDD.t1943 VDD.t1942 VDD.t1943 VDD.t321 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4585 a_108602_n27257# a_100820_n36322.t17 a_100992_n29313.t0 VSS.t351 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4586 a_49755_13546# a_47819_10448.t16 VDD.t514 VDD.t498 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4587 VDD.t1941 VDD.t1940 VDD.t1941 VDD.t1572 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4588 a_52635_49681.t109 a_52635_34067.t194 VDD.t4854 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4589 VSS.t1576 VSS.t1575 VSS.t1576 VSS.t555 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4590 VDD.t1939 VDD.t1937 VDD.t1939 VDD.t1938 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4591 VDD.t1936 VDD.t1935 VDD.t1936 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4592 VDD.t1934 VDD.t1933 VDD.t1934 VDD.t315 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4593 VDD.t4779 a_71266_n4019.t0 a_72596_n3060# VDD.t1191 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X4594 a_52635_49681.t59 a_35922_19591.t137 OUT.t48 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4595 a_33249_48695.t210 a_31699_20742.t200 VDD.t225 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4596 VDD.t1932 VDD.t1931 VDD.t1932 VDD.t1180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4597 a_108636_n35156# a_106830_n36382.t22 VSS.t430 VDD.t1542 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4598 a_111631_n18620# a_71281_n8397.t259 a_111063_n18620# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4599 a_104527_n4245# a_71281_n8397.t260 a_103997_n4245# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4600 VDD.t1930 VDD.t1929 VDD.t1930 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4601 VSS.t1574 VSS.t1573 VSS.t1574 VSS.t480 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4602 VSS.t1572 VSS.t1571 VSS.t1572 VSS.t98 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4603 a_71281_n10073.t17 a_71281_n10073.t16 VDD.t327 VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4604 VSS.t1570 VSS.t1569 VSS.t1570 VSS.t298 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4605 a_41487_n14213# a_31953_n19727.t277 a_40965_n14213# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4606 a_48391_n30339# a_39179_n19595.t0 a_47819_n36322.t7 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4607 VDD.t4853 a_52635_34067.t195 a_52635_49681.t108 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4608 VDD.t1928 VDD.t1927 VDD.t1928 VDD.t1325 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4609 a_38619_n7136# a_31953_n19727.t278 a_38097_n7136# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4610 VDD.t1926 VDD.t1925 VDD.t1926 VDD.t1052 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4611 VSS.t1568 VSS.t1567 VSS.t1568 VSS.t1227 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4612 VSS.t1566 VSS.t1565 VSS.t1566 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4613 VSS.t1564 VSS.t1563 VSS.t1564 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4614 a_84017_n17715.t3 a_81205_n14095.t5 a_95443_13546# VDD.t501 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4615 a_83683_10448# a_83153_10448.t4 a_83153_10448.t5 VDD.t2776 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4616 a_60677_10448.t2 a_47991_4421.t1 a_60109_12380# VDD.t494 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4617 VDD.t434 a_71281_n8397.t14 a_71281_n8397.t15 VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4618 VSS.t1562 VSS.t1561 VSS.t1562 VSS.t492 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4619 VSS.t1560 VSS.t1559 VSS.t1560 VSS.t709 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4620 a_49755_11614# a_47819_10448.t17 VDD.t515 VDD.t498 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4621 VDD.t1924 VDD.t1923 VDD.t1924 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4622 VSS.t1558 VSS.t1557 VSS.t1558 VSS.t614 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4623 VDD.t1922 VDD.t1921 VDD.t1922 VDD.t79 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4624 VDD.t1920 VDD.t1918 VDD.t1920 VDD.t1919 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4625 a_33249_48695.t129 a_33379_34007.t65 a_33249_34067.t45 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4626 a_36530_n29181# a_30152_n36322.t18 VDD.t4775 VSS.t326 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4627 VSS.t1556 VSS.t1555 VSS.t1556 VSS.t489 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4628 VDD.t1917 VDD.t1916 VDD.t1917 VDD.t52 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4629 a_108636_n33224# a_106830_n36382.t23 a_106676_n30339.t2 VDD.t1542 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4630 VSS.t1554 VSS.t1553 VSS.t1554 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4631 VSS.t1552 VSS.t1551 VSS.t1552 VSS.t620 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4632 VSS.t1550 VSS.t1549 VSS.t1550 VSS.t573 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4633 a_33249_35053.t119 a_35502_25545.t77 VSS.t50 VSS.t49 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4634 VDD.t1915 VDD.t1914 VDD.t1915 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4635 VDD.t1913 VDD.t1912 VDD.t1913 VDD.t572 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4636 VSS.t1548 VSS.t1547 VSS.t1548 VSS.t655 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4637 VDD.t1911 VDD.t1910 VDD.t1911 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4638 a_33249_48695.t80 a_33379_34917.t65 a_33249_35053.t63 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4639 VDD.t1909 VDD.t1908 VDD.t1909 VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4640 a_33249_34067.t44 a_33379_34007.t66 a_33249_48695.t130 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4641 VSS.t1546 VSS.t1545 VSS.t1546 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4642 VDD.t1907 VDD.t1905 VDD.t1907 VDD.t1906 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4643 VSS.t5 a_35502_25545.t78 a_33249_35053.t118 VSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4644 a_84017_n17715.t2 a_81205_n14095.t6 a_95443_11614# VDD.t501 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4645 a_51711_n8932# a_50751_n19729.t267 a_51151_n8932# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4646 VDD.t1904 VDD.t1903 VDD.t1904 VDD.t783 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4647 VDD.t1902 VDD.t1901 VDD.t1902 VDD.t556 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4648 a_33249_34067.t43 a_33379_34007.t67 a_33249_48695.t131 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4649 a_51711_n18700# a_50751_n19729.t268 a_51151_n17803# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4650 VSS.t1544 VSS.t1542 VSS.t1544 VSS.t1543 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4651 VDD.t1900 VDD.t1899 VDD.t1900 VDD.t680 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4652 a_44885_n14213# a_31953_n19727.t279 a_44363_n15110# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4653 VDD.t1898 VDD.t1897 VDD.t1898 VDD.t677 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4654 VDD.t1896 VDD.t1894 VDD.t1896 VDD.t1895 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4655 a_83153_n36322.t3 a_32913_n8930.t1 a_85129_n27257# VSS.t365 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4656 VDD.t1893 VDD.t1892 VDD.t1893 VDD.t1508 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4657 VDD.t1891 VDD.t1890 VDD.t1891 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4658 a_95943_n18620# a_71281_n10073.t253 a_95105_n15905# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4659 VSS.t1541 VSS.t1540 VSS.t1541 VSS.t673 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4660 a_110225_n6960# a_71281_n8397.t261 a_109695_n7865# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4661 a_84547_n3340# a_71281_n10073.t254 a_83709_n2435# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4662 a_88271_n8770# a_71281_n10073.t255 a_87433_n8770# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4663 VDD.t1889 VDD.t1888 VDD.t1889 VDD.t489 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4664 a_52635_49681.t60 a_35922_19591.t138 OUT.t47 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4665 VDD.t1887 VDD.t1885 VDD.t1887 VDD.t1886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4666 a_60845_n8932# a_50751_n19729.t269 a_60285_n8035# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4667 VDD.t1884 VDD.t1883 VDD.t1884 VDD.t15 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4668 VDD.t1882 VDD.t1881 VDD.t1882 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4669 VSS.t1539 VSS.t1538 VSS.t1539 VSS.t218 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4670 a_52635_34067.t41 a_35922_19591.t139 a_52635_48695.t26 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4671 VSS.t307 I1N.t11 a_72603_n10073# VSS.t305 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X4672 a_110225_n17715# a_71281_n8397.t262 a_109695_n21335# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4673 a_33249_34067.t42 a_33379_34007.t68 a_33249_48695.t132 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4674 a_50751_n19729.t33 a_50751_n19729.t32 VSS.t229 VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4675 VSS.t1537 VSS.t1536 VSS.t1537 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4676 VDD.t1880 VDD.t1879 VDD.t1880 VDD.t1492 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4677 VSS.t1535 VSS.t1534 VSS.t1535 VSS.t655 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4678 VDD.t1878 VDD.t1877 VDD.t1878 VDD.t1167 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4679 VDD.t1876 VDD.t1875 VDD.t1876 VDD.t1508 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4680 VDD.t1874 VDD.t1873 VDD.t1874 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4681 VSS.t1533 VSS.t1532 VSS.t1533 VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4682 a_93969_n14095# a_71281_n10073.t256 a_93131_n14095# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4683 a_52635_48695.t112 a_52635_34067.t196 VDD.t4852 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4684 a_83153_n36322.t7 a_83153_n35156.t20 a_85089_n35156# VDD.t1489 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4685 a_90935_5639# a_83153_11614.t19 a_51711_n12421.t0 VSS.t401 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4686 VSS.t1531 VSS.t1530 VSS.t1531 VSS.t646 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4687 a_52635_49681.t107 a_52635_34067.t197 VDD.t4851 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4688 VSS.t1529 VSS.t1528 VSS.t1529 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4689 a_94537_n15905# a_71281_n10073.t257 a_93969_n15905# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4690 a_71266_n4019.t0 I1N.t12 a_75585_n9297# VSS.t301 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X4691 VSS.t1527 VSS.t1526 VSS.t1527 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4692 VDD.t1872 VDD.t1871 VDD.t1872 VDD.t1191 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X4693 VDD.t1870 VDD.t1868 VDD.t1870 VDD.t1869 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4694 VDD.t1867 VDD.t1866 VDD.t1867 VDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4695 a_52635_49681.t106 a_52635_34067.t198 VDD.t4850 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4696 a_60285_n7138# a_50751_n19729.t270 a_59763_n8035# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4697 VDD.t1865 VDD.t1864 VDD.t1865 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4698 a_42413_n27257# a_41891_n29181.t3 a_41891_n29181.t4 VSS.t177 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4699 VDD.t1863 VDD.t1862 VDD.t1863 VDD.t1484 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4700 VDD.t1861 VDD.t1860 VDD.t1861 VDD.t1130 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4701 VDD.t4849 a_52635_34067.t199 a_52635_48695.t111 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4702 VDD.t1859 VDD.t1858 VDD.t1859 VDD.t1492 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4703 a_35221_n16007# a_31953_n19727.t280 a_34347_n17801# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4704 VSS.t1525 VSS.t1524 VSS.t1525 VSS.t167 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4705 a_47819_10448.t0 a_47991_4421.t0 a_49795_7563# VSS.t282 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4706 VSS.t1523 VSS.t1522 VSS.t1523 VSS.t1069 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4707 a_67111_n19597# a_50751_n19729.t271 a_66551_n19597# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4708 a_101641_n3340# a_71281_n8397.t263 a_100803_n3340# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4709 a_66058_5639# a_64243_n1756.t1 a_65486_11614.t7 VSS.t410 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4710 VSS.t1521 VSS.t1520 VSS.t1521 VSS.t558 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4711 VDD.t1857 VDD.t1856 VDD.t1857 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4712 a_33249_34067.t41 a_33379_34007.t69 a_33249_48695.t133 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4713 OUT.t6 a_35502_24538.t53 a_33249_35053.t101 VSS.t182 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4714 VDD.t1855 VDD.t1854 VDD.t1855 VDD.t529 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4715 a_83153_n36322.t6 a_83153_n35156.t21 a_85089_n33224# VDD.t1489 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4716 a_33249_35053.t117 a_35502_25545.t79 VSS.t122 VSS.t9 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4717 VSS.t1519 VSS.t1518 VSS.t1519 VSS.t181 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4718 VDD.t1853 VDD.t1851 VDD.t1853 VDD.t1852 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4719 a_89163_n36382.t6 a_94892_n29181.t18 a_96818_n27257# VSS.t445 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4720 a_31699_20742.t0 I1U.t5 a_30377_19942# VSS.t362 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X4721 a_52635_48695.t25 a_35922_19591.t140 a_52635_34067.t9 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4722 VDD.t1850 VDD.t1849 VDD.t1850 VDD.t1484 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4723 a_35221_n2651# a_31953_n19727.t281 a_34699_n3548# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4724 VDD.t1848 VDD.t1847 VDD.t1848 VDD.t1115 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4725 VDD.t1846 VDD.t1845 VDD.t1846 VDD.t313 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4726 VDD.t1844 VDD.t1842 VDD.t1844 VDD.t1843 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4727 VDD.t1841 VDD.t1840 VDD.t1841 VDD.t123 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4728 VSS.t1517 VSS.t1516 VSS.t1517 VSS.t384 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4729 VSS.t3649 a_94892_4481.t22 a_95414_4481# VSS.t1042 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4730 VDD.t1839 VDD.t1838 VDD.t1839 VDD.t554 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4731 a_33249_48695.t209 a_31699_20742.t201 VDD.t226 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4732 a_114516_n35156# a_103997_n8770.t11 a_106809_n5150.t3 VDD.t329 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4733 a_63683_n13318# a_50751_n19729.t272 a_63161_n13318# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4734 VSS.t1515 VSS.t1514 VSS.t1515 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4735 a_52635_49681.t61 a_35922_19591.t141 OUT.t46 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4736 a_57977_n6241# a_50751_n19729.t273 a_57417_n6241# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4737 VSS.t1513 VSS.t1512 VSS.t1513 VSS.t426 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4738 VDD.t1837 VDD.t1836 VDD.t1837 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4739 VDD.t1835 VDD.t1834 VDD.t1835 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4740 VSS.t1511 VSS.t1510 VSS.t1511 VSS.t623 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4741 VDD.t1833 VDD.t1832 VDD.t1833 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4742 a_38619_n19595# a_31953_n19727.t282 a_38097_n19595# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4743 VSS.t1509 VSS.t1508 VSS.t1509 VSS.t316 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4744 VSS.t1507 VSS.t1506 VSS.t1507 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4745 VDD.t227 a_31699_20742.t202 a_33249_48695.t208 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4746 a_52635_48695.t24 a_35922_19591.t142 a_52635_34067.t11 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4747 a_31699_20742.t20 a_31699_20742.t19 VDD.t32 VDD.t21 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4748 a_51151_n5344# a_50751_n19729.t274 a_31284_4481.t0 VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4749 VDD.t1831 VDD.t1830 VDD.t1831 VDD.t572 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4750 VDD.t1829 VDD.t1828 VDD.t1829 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4751 a_88839_n1530# a_71281_n10073.t258 a_88271_n1530# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4752 VSS.t1505 VSS.t1504 VSS.t1505 VSS.t839 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4753 a_95943_n3340# a_71281_n10073.t259 a_95105_n2435# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4754 VSS.t1503 VSS.t1502 VSS.t1503 VSS.t1030 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4755 a_110225_n21335# a_71281_n8397.t264 a_109695_n21335# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4756 VDD.t1827 VDD.t1825 VDD.t1827 VDD.t1826 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4757 a_77747_n30339# a_77225_n29181.t18 a_71496_n36382.t2 VSS.t385 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4758 a_50751_n19729.t31 a_50751_n19729.t30 VSS.t228 VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4759 VDD.t1824 VDD.t1822 VDD.t1824 VDD.t1823 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4760 VDD.t1821 VDD.t1819 VDD.t1821 VDD.t1820 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4761 VSS.t1501 VSS.t1500 VSS.t1501 VSS.t173 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4762 VDD.t1818 VDD.t1817 VDD.t1818 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4763 VSS.t1499 VSS.t1498 VSS.t1499 VSS.t146 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4764 a_114516_n33224# a_103997_n8770.t12 a_106809_n5150.t2 VDD.t329 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4765 VDD.t1816 VDD.t1815 VDD.t1816 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4766 a_46879_n13316# a_31953_n19727.t283 a_46319_n12419# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4767 a_48391_7563# a_47991_5507.t0 a_47819_11614.t4 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4768 VSS.t121 a_35502_25545.t80 a_33249_35053.t116 VSS.t35 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4769 VSS.t1497 VSS.t1496 VSS.t1497 VSS.t254 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4770 VDD.t1814 VDD.t1813 VDD.t1814 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4771 VSS.t1495 VSS.t1494 VSS.t1495 VSS.t156 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4772 VDD.t522 a_47819_n36322.t18 a_55601_n28415# VSS.t328 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4773 VSS.t1493 VSS.t1492 VSS.t1493 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4774 VDD.t1812 VDD.t1811 VDD.t1812 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4775 VDD.t1810 VDD.t1809 VDD.t1810 VDD.t328 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4776 a_93969_n4245# a_71281_n10073.t260 a_93131_n4245# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4777 VDD.t1808 VDD.t1807 VDD.t1808 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4778 VDD.t1806 VDD.t1805 VDD.t1806 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4779 a_32913_n16904# a_31953_n19727.t284 a_32353_n15110# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4780 VDD.t1804 VDD.t1803 VDD.t1804 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4781 a_33249_34067.t40 a_33379_34007.t70 a_33249_48695.t134 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4782 a_60080_n27257# a_59558_n29181.t4 a_59558_n29181.t5 VSS.t313 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4783 VSS.t1491 VSS.t1490 VSS.t1491 VSS.t160 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4784 a_42047_n8930# a_31953_n19727.t285 a_41487_n8930# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4785 VDD.t1802 VDD.t1800 VDD.t1802 VDD.t1801 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4786 VDD.t1799 VDD.t1797 VDD.t1799 VDD.t1798 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4787 VDD.t1796 VDD.t1795 VDD.t1796 VDD.t1084 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4788 VDD.t1794 VDD.t1793 VDD.t1794 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4789 VDD.t1792 VDD.t1791 VDD.t1792 VDD.t1427 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4790 VDD.t1790 VDD.t1788 VDD.t1790 VDD.t1789 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4791 a_47753_n1754# a_31953_n19727.t286 a_45445_n1754# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4792 a_71281_n8397.t13 a_71281_n8397.t12 VDD.t432 VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4793 a_71496_n36382.t3 a_77225_n29181.t19 a_79151_n29181# VSS.t386 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4794 OUT.t45 a_35922_19591.t143 a_52635_49681.t62 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4795 a_33249_35053.t64 a_33379_34917.t66 a_33249_48695.t81 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4796 VDD.t4788 a_83153_n36322.t19 a_90935_n29181# VSS.t460 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4797 a_102756_10448# a_100820_10448.t17 VDD.t367 VDD.t325 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4798 VSS.t120 a_35502_25545.t81 a_33249_35053.t115 VSS.t44 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4799 a_95414_4481# a_94892_4481.t2 a_94892_4481.t3 VSS.t1003 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4800 VDD.t1787 VDD.t1786 VDD.t1787 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4801 a_40613_n17801# a_31953_n19727.t287 a_40053_n17801# VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4802 VDD.t31 a_31699_20742.t17 a_31699_20742.t18 VDD.t30 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4803 VDD.t4848 a_52635_34067.t200 a_52635_48695.t110 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4804 VDD.t1785 VDD.t1784 VDD.t1785 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4805 a_65117_n14215# a_50751_n19729.t275 a_64595_n14215# VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4806 VSS.t1489 VSS.t1488 VSS.t1489 VSS.t952 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4807 VDD.t1783 VDD.t1781 VDD.t1783 VDD.t1782 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4808 VSS.t1487 VSS.t1486 VSS.t1487 VSS.t480 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4809 VSS.t1485 VSS.t1484 VSS.t1485 VSS.t252 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4810 a_63683_n4447# a_50751_n19729.t276 a_63161_n4447# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4811 VSS.t1483 VSS.t1482 VSS.t1483 VSS.t503 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4812 VDD.t1780 VDD.t1779 VDD.t1780 VDD.t1411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4813 VSS.t1481 VSS.t1480 VSS.t1481 VSS.t593 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4814 a_59411_n14215# a_50751_n19729.t277 a_58851_n14215# VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4815 VSS.t1479 VSS.t1478 VSS.t1479 VSS.t175 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4816 VDD.t1778 VDD.t1777 VDD.t1778 VDD.t1427 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4817 a_50751_n19729.t29 a_50751_n19729.t28 VSS.t227 VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4818 VSS.t1477 VSS.t1476 VSS.t1477 VSS.t514 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4819 VDD.t1776 VDD.t1775 VDD.t1776 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4820 VSS.t1475 VSS.t1474 VSS.t1475 VSS.t134 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4821 VSS.t1473 VSS.t1471 VSS.t1473 VSS.t1472 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4822 a_71281_n8397.t11 a_71281_n8397.t10 VDD.t430 VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4823 VSS.t1470 VSS.t1469 VSS.t1470 VSS.t325 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4824 VDD.t1774 VDD.t1773 VDD.t1774 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4825 a_60285_n12421# a_50751_n19729.t278 VSS.t269 VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4826 a_89033_n35156.t3 a_89163_n36382.t20 a_90969_n35156# VDD.t551 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4827 a_33249_34067.t39 a_33379_34007.t71 a_33249_48695.t135 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4828 a_57417_n18700# a_50751_n19729.t279 a_56895_n19597# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4829 VSS.t1468 VSS.t1467 VSS.t1468 VSS.t1082 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X4830 VSS.t1466 VSS.t1465 VSS.t1466 VSS.t145 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4831 a_83141_n1530# a_71281_n10073.t261 a_82573_n1530# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4832 a_35502_25545.t23 a_35502_25545.t22 VSS.t169 VSS.t2 nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X4833 VSS.t1464 VSS.t1463 VSS.t1464 VSS.t1366 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4834 VSS.t1462 VSS.t1461 VSS.t1462 VSS.t573 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4835 VDD.t1772 VDD.t1771 VDD.t1772 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4836 VDD.t1770 VDD.t1769 VDD.t1770 VDD.t1052 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4837 VDD.t1768 VDD.t1767 VDD.t1768 VDD.t836 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4838 VDD.t1766 VDD.t1765 VDD.t1766 VDD.t1055 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4839 VSS.t1460 VSS.t1459 VSS.t1460 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4840 a_60845_n4447# a_50751_n19729.t280 a_60285_n3550# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4841 VDD.t1764 VDD.t1763 VDD.t1764 VDD.t1411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4842 a_100235_n1530# a_71281_n8397.t265 a_99667_n1530# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4843 VSS.t1458 VSS.t1457 VSS.t1458 VSS.t469 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4844 VDD.t1762 VDD.t1761 VDD.t1762 VDD.t433 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4845 a_54197_5639# a_47819_11614.t17 VDD.t509 VSS.t329 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4846 a_33249_48695.t207 a_31699_20742.t203 VDD.t228 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4847 a_52635_49681.t105 a_52635_34067.t201 VDD.t4847 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4848 VDD.t1760 VDD.t1759 VDD.t1760 VDD.t1376 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4849 VDD.t1758 VDD.t1757 VDD.t1758 VDD.t1373 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4850 VDD.t14 a_30152_10448.t15 a_30682_13546# VDD.t13 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4851 VDD.t1756 VDD.t1755 VDD.t1756 VDD.t374 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4852 a_89033_n36322.t2 a_89163_n36382.t21 a_90969_n33224# VDD.t551 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4853 a_78344_10448.t0 a_65658_4421.t2 a_77776_12380# VDD.t3571 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4854 a_53699_11614.t0 a_53829_10388.t21 a_55635_12380# VDD.t3748 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4855 VSS.t1456 VSS.t1455 VSS.t1456 VSS.t542 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4856 a_96849_13546# a_83325_4421.t1 a_84017_n17715.t2 VDD.t502 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4857 VDD.t1754 VDD.t1753 VDD.t1754 VDD.t1368 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4858 VSS.t1454 VSS.t1453 VSS.t1454 VSS.t550 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4859 a_88271_n7865# a_71281_n10073.t262 a_87433_n7865# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4860 VDD.t1752 VDD.t1751 VDD.t1752 VDD.t61 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4861 a_101641_n17715# a_71281_n8397.t266 a_43010_n36322.t3 VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4862 a_87433_n14095# a_71281_n10073.t263 a_86903_n14095.t2 VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4863 VDD.t1750 VDD.t1748 VDD.t1750 VDD.t1749 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4864 a_101641_n15000# a_71281_n8397.t267 a_100803_n15000# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4865 VSS.t1452 VSS.t1451 VSS.t1452 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4866 VDD.t1747 VDD.t1746 VDD.t1747 VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4867 a_111631_n21335# a_71281_n8397.t268 a_111063_n21335# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4868 VDD.t1745 VDD.t1744 VDD.t1745 VDD.t1376 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4869 VDD.t1743 VDD.t1742 VDD.t1743 VDD.t1373 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4870 VDD.t365 a_30152_10448.t16 a_30682_11614# VDD.t13 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4871 VDD.t1741 VDD.t1740 VDD.t1741 VDD.t1357 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4872 VSS.t1450 VSS.t1449 VSS.t1450 VSS.t542 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4873 VDD.t1739 VDD.t1738 VDD.t1739 VDD.t1368 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4874 VSS.t1448 VSS.t1447 VSS.t1448 VSS.t800 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4875 a_96849_11614# a_83325_4421.t1 a_84017_n17715.t0 VDD.t502 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4876 VDD.t1737 VDD.t1736 VDD.t1737 VDD.t61 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4877 VDD.t1735 VDD.t1734 VDD.t1735 VDD.t1352 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4878 VDD.t484 a_71281_n8397.t269 a_112199_n1530# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4879 VSS.t12 a_35502_25545.t82 a_33249_35053.t114 VSS.t11 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4880 VSS.t1446 VSS.t1445 VSS.t1446 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4881 a_33249_34067.t4 a_35502_24538.t54 a_52635_34067.t63 VSS.t182 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4882 a_48313_n17801# a_31953_n19727.t288 a_47753_n16904# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4883 a_112559_n29181.t4 a_112559_n29181.t3 a_114485_n30339# VSS.t414 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4884 a_33249_48695.t206 a_31699_20742.t204 VDD.t229 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4885 VDD.t1733 VDD.t1732 VDD.t1733 VDD.t12 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4886 VSS.t1444 VSS.t1443 VSS.t1444 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4887 VSS.t1442 VSS.t1441 VSS.t1442 VSS.t98 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4888 VSS.t1440 VSS.t1439 VSS.t1440 VSS.t18 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4889 VDD.t230 a_31699_20742.t205 a_33249_48695.t205 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4890 a_58851_n17803# a_50751_n19729.t281 a_58329_n18700# VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4891 VSS.t1438 VSS.t1436 VSS.t1438 VSS.t1437 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4892 VSS.t1435 VSS.t1434 VSS.t1435 VSS.t362 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4893 VDD.t231 a_31699_20742.t206 a_33249_48695.t204 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4894 VDD.t1731 VDD.t1730 VDD.t1731 VDD.t1357 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4895 VDD.t1729 VDD.t1728 VDD.t1729 VDD.t558 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4896 a_52635_48695.t109 a_52635_34067.t202 VDD.t4846 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4897 VDD.t1727 VDD.t1726 VDD.t1727 VDD.t1018 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4898 a_101641_n3340# a_71281_n8397.t270 a_100803_n2435# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4899 VDD.t1725 VDD.t1724 VDD.t1725 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4900 VDD.t1723 VDD.t1722 VDD.t1723 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4901 VDD.t1721 VDD.t1720 VDD.t1721 VDD.t1352 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4902 a_36008_n27257.t3 a_30152_n36322.t19 a_37934_n30339# VSS.t323 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4903 a_107339_n17715# a_71281_n8397.t271 a_60677_n36322.t0 VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4904 a_47991_5507.t1 a_50751_n19729.t282 a_57417_n1756# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4905 a_37934_7563# a_30152_11614.t16 a_30324_4421.t0 VSS.t324 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4906 a_33249_48695.t203 a_31699_20742.t207 VDD.t232 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4907 a_52635_48695.t108 a_52635_34067.t203 VDD.t4845 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4908 a_107339_n15000# a_71281_n8397.t272 a_106501_n15000# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4909 VSS.t1433 VSS.t1431 VSS.t1433 VSS.t1432 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4910 VSS.t1430 VSS.t1429 VSS.t1430 VSS.t536 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4911 VSS.t1428 VSS.t1427 VSS.t1428 VSS.t399 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4912 VSS.t1426 VSS.t1425 VSS.t1426 VSS.t738 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4913 a_65658_4421.t0 a_65486_11614.t23 a_71864_4481# VSS.t429 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4914 VDD.t1719 VDD.t1718 VDD.t1719 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4915 VDD.t1717 VDD.t1715 VDD.t1717 VDD.t1716 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4916 VDD.t1714 VDD.t1712 VDD.t1714 VDD.t1713 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4917 VSS.t1424 VSS.t1423 VSS.t1424 VSS.t500 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4918 VSS.t1422 VSS.t1421 VSS.t1422 VSS.t412 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4919 VDD.t1711 VDD.t1709 VDD.t1711 VDD.t1710 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4920 a_71366_11614.t1 a_71496_10388.t20 a_73302_12380# VDD.t490 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4921 VDD.t1708 VDD.t1707 VDD.t1708 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4922 VDD.t1706 VDD.t1705 VDD.t1706 VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4923 VDD.t1704 VDD.t1703 VDD.t1704 VDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4924 VDD.t1702 VDD.t1701 VDD.t1702 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4925 a_38097_n5342.t1 a_100992_n29313.t1 a_101392_n27257# VSS.t384 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4926 a_101641_n20430# a_71281_n8397.t273 a_100803_n20430# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4927 VDD.t1700 VDD.t1699 VDD.t1700 VDD.t315 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4928 VSS.t1420 VSS.t1419 VSS.t1420 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4929 VDD.t1698 VDD.t1697 VDD.t1698 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4930 VSS.t1418 VSS.t1417 VSS.t1418 VSS.t413 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4931 VSS.t1416 VSS.t1415 VSS.t1416 VSS.t1039 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4932 VDD.t1696 VDD.t1695 VDD.t1696 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4933 VSS.t1414 VSS.t1413 VSS.t1414 VSS.t483 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4934 a_43817_n28415# a_41891_n29181.t20 VSS.t377 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4935 VDD.t233 a_31699_20742.t208 a_33249_48695.t202 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4936 VDD.t4844 a_52635_34067.t204 a_52635_48695.t107 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4937 VDD.t29 a_31699_20742.t15 a_31699_20742.t16 VDD.t28 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4938 a_106809_n6055.t0 a_71281_n8397.t274 a_106501_n9675# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4939 VSS.t1412 VSS.t1411 VSS.t1412 VSS.t692 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4940 VSS.t1410 VSS.t1409 VSS.t1410 VSS.t949 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4941 a_33249_48695.t201 a_31699_20742.t209 VDD.t234 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4942 a_52635_49681.t104 a_52635_34067.t205 VDD.t4843 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4943 VDD.t1694 VDD.t1693 VDD.t1694 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4944 VSS.t1408 VSS.t1407 VSS.t1408 VSS.t1242 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4945 VDD.t1692 VDD.t1691 VDD.t1692 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4946 a_49795_n28415# a_47991_n29313.t0 a_38097_n16007.t1 VSS.t281 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4947 a_33249_48695.t200 a_31699_20742.t210 VDD.t235 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4948 a_100820_n35156.t8 a_100820_n35156.t7 a_102756_n34390# VDD.t528 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4949 a_50751_n19729.t27 a_50751_n19729.t26 VSS.t226 VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4950 a_41891_4481.t10 a_30324_4421.t1 a_43848_13546# VDD.t290 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4951 VDD.t1690 VDD.t1689 VDD.t1690 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4952 VSS.t1406 VSS.t1405 VSS.t1406 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4953 VSS.t1404 VSS.t1403 VSS.t1404 VSS.t563 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4954 VDD.t1688 VDD.t1687 VDD.t1688 VDD.t1660 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4955 VDD.t1686 VDD.t1685 VDD.t1686 VDD.t424 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4956 VDD.t1684 VDD.t1683 VDD.t1684 VDD.t332 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4957 VSS.t1402 VSS.t1401 VSS.t1402 VSS.t500 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4958 a_73268_n27257# a_65486_n36322.t21 a_65658_n29313.t0 VSS.t156 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4959 VDD.t1682 VDD.t1681 VDD.t1682 VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4960 VSS.t1400 VSS.t1399 VSS.t1400 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4961 VSS.t1398 VSS.t1397 VSS.t1398 VSS.t96 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4962 a_72596_n3060# a_71266_n4019.t0 a_50751_n19729.t72 VDD.t997 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X4963 VSS.t1396 VSS.t1395 VSS.t1396 VSS.t290 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4964 VSS.t1394 VSS.t1393 VSS.t1394 VSS.t400 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4965 VSS.t1392 VSS.t1390 VSS.t1392 VSS.t1391 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4966 a_105365_n6960# a_71281_n8397.t275 a_104527_n6960# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4967 VSS.t1389 VSS.t1388 VSS.t1389 VSS.t257 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4968 a_60285_n6241# a_50751_n19729.t283 a_59763_n6241# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4969 VDD.t1680 VDD.t1679 VDD.t1680 VDD.t422 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4970 VSS.t1387 VSS.t1386 VSS.t1387 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4971 VDD.t1678 VDD.t1677 VDD.t1678 VDD.t420 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4972 VDD.t1676 VDD.t1675 VDD.t1676 VDD.t438 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4973 VSS.t1385 VSS.t1384 VSS.t1385 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4974 VSS.t225 a_50751_n19729.t24 a_50751_n19729.t25 VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4975 a_107339_n20430# a_71281_n8397.t276 a_106501_n20430# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4976 a_95943_n15000# a_71281_n10073.t264 a_95105_n14095# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4977 a_105933_n1530# a_71281_n8397.t277 a_105365_n1530# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4978 a_34347_n19595# a_31953_n19727.t289 a_33787_n19595# VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4979 VDD.t536 a_100820_n35156.t17 a_101350_n34390# VDD.t535 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4980 a_52635_49681.t63 a_35922_19591.t144 OUT.t44 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4981 VDD.t1674 VDD.t1673 VDD.t1674 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4982 a_33249_48695.t199 a_31699_20742.t211 VDD.t236 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4983 a_41891_4481.t9 a_30324_4421.t1 a_43848_11614# VDD.t290 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4984 VDD.t1672 VDD.t1671 VDD.t1672 VDD.t968 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4985 a_107230_12380# a_106830_10388.t18 a_86903_n14095.t1 VDD.t527 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4986 VDD.t1670 VDD.t1669 VDD.t1670 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4987 VSS.t1383 VSS.t1382 VSS.t1383 VSS.t387 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4988 a_47991_n29313.t0 a_47819_n36322.t19 a_54197_n30339# VSS.t327 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4989 VSS.t1381 VSS.t1380 VSS.t1381 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4990 VSS.t1379 VSS.t1378 VSS.t1379 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4991 VSS.t10 a_35502_25545.t83 a_33249_35053.t113 VSS.t9 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4992 VDD.t4842 a_52635_34067.t206 a_52635_49681.t103 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4993 a_75585_n10973# I1N.t13 VSS.t308 VSS.t303 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X4994 VDD.t1668 VDD.t1666 VDD.t1668 VDD.t1667 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X4995 a_82573_n19525# a_71281_n10073.t265 a_81735_n19525# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4996 a_111063_n4245# a_71281_n8397.t278 a_110225_n4245# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4997 a_52585_n8035# a_50751_n19729.t284 a_52063_n8035# VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4998 a_33249_48695.t198 a_31699_20742.t212 VDD.t237 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4999 a_65677_n7138# a_50751_n19729.t285 a_66551_n5344# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5000 a_63683_n12421# a_50751_n19729.t286 a_63161_n13318# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5001 VDD.t1665 VDD.t1664 VDD.t1665 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5002 a_54579_n8932# a_50751_n19729.t287 a_54019_n8035# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5003 VDD.t1663 VDD.t1662 VDD.t1663 VDD.t301 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5004 VSS.t1377 VSS.t1376 VSS.t1377 VSS.t1109 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5005 VSS.t1375 VSS.t1374 VSS.t1375 VSS.t367 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5006 VDD.t1661 VDD.t1659 VDD.t1661 VDD.t1660 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5007 VSS.t1373 VSS.t1372 VSS.t1373 VSS.t576 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5008 VSS.t69 a_31953_n19727.t22 a_31953_n19727.t23 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5009 a_94537_n14095# a_71281_n10073.t266 a_93969_n14095# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5010 a_30324_n29313.t0 a_30152_n36322.t20 a_36530_n27257# VSS.t325 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5011 VDD.t1658 VDD.t1657 VDD.t1658 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5012 VSS.t1371 VSS.t1370 VSS.t1371 VSS.t1258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5013 VDD.t1656 VDD.t1654 VDD.t1656 VDD.t1655 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5014 a_35781_n13316# a_31953_n19727.t290 a_35221_n12419# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5015 VSS.t1369 VSS.t1368 VSS.t1369 VSS.t873 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5016 VDD.t1653 VDD.t1652 VDD.t1653 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5017 VDD.t1651 VDD.t1650 VDD.t1651 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5018 a_33249_34067.t117 a_35502_25545.t84 VSS.t8 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5019 VDD.t1649 VDD.t1648 VDD.t1649 VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5020 a_36562_n34390# a_36162_n36382.t20 a_36032_n35156.t3 VDD.t683 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5021 a_33249_34067.t38 a_33379_34007.t72 a_33249_48695.t136 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5022 VSS.t1367 VSS.t1365 VSS.t1367 VSS.t1366 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5023 VSS.t1364 VSS.t1363 VSS.t1364 VSS.t412 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5024 a_55601_n29181# a_47819_n36322.t20 a_39179_n19595.t0 VSS.t330 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5025 VSS.t1362 VSS.t1361 VSS.t1362 VSS.t218 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5026 a_101641_n18620# a_71281_n8397.t279 a_100803_n15905# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5027 VSS.t1360 VSS.t1359 VSS.t1360 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5028 VDD.t1647 VDD.t1646 VDD.t1647 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5029 a_90245_n6055# a_71281_n10073.t267 a_89715_n5150.t0 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5030 VSS.t1358 VSS.t1357 VSS.t1358 VSS.t563 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5031 VSS.t1356 VSS.t1355 VSS.t1356 VSS.t981 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5032 a_47753_n17801# a_31953_n19727.t291 a_47231_n18698# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5033 a_66058_n28415# a_45445_n19595.t1 a_65486_n36322.t7 VSS.t410 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5034 a_52635_48695.t106 a_52635_34067.t207 VDD.t4841 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5035 VDD.t1645 VDD.t1643 VDD.t1645 VDD.t1644 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5036 VDD.t1642 VDD.t1641 VDD.t1642 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5037 VDD.t1640 VDD.t1639 VDD.t1640 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5038 VSS.t406 a_59558_4481.t17 a_60080_7563# VSS.t316 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5039 VSS.t158 a_35502_25545.t20 a_35502_25545.t21 VSS.t126 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X5040 VSS.t1354 VSS.t1353 VSS.t1354 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5041 VSS.t1352 VSS.t1351 VSS.t1352 VSS.t896 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5042 VSS.t1350 VSS.t1348 VSS.t1350 VSS.t1349 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5043 VDD.t1638 VDD.t1637 VDD.t1638 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5044 VSS.t1347 VSS.t1346 VSS.t1347 VSS.t542 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5045 a_32913_n14213# a_31953_n19727.t292 a_32353_n14213# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5046 VDD.t1636 VDD.t1635 VDD.t1636 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5047 a_83153_10448.t0 a_83325_4421.t0 a_85129_7563# VSS.t297 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5048 VSS.t1345 VSS.t1344 VSS.t1345 VSS.t913 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5049 VSS.t1343 VSS.t1342 VSS.t1343 VSS.t882 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5050 a_38619_n1754# a_31953_n19727.t293 a_38097_n2651# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5051 VDD.t1634 VDD.t1633 VDD.t1634 VDD.t550 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5052 VSS.t1341 VSS.t1340 VSS.t1341 VSS.t873 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5053 VDD.t1632 VDD.t1631 VDD.t1632 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5054 VDD.t1630 VDD.t1629 VDD.t1630 VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5055 VDD.t1628 VDD.t1627 VDD.t1628 VDD.t1254 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5056 a_100992_4421.t0 a_100820_11614.t19 a_107198_4481# VSS.t188 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5057 VDD.t4840 a_52635_34067.t208 a_52635_48695.t105 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5058 a_53145_n19597# a_50751_n19729.t288 a_52585_n18700# VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5059 VDD.t1626 VDD.t1625 VDD.t1626 VDD.t997 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X5060 VSS.t1339 VSS.t1338 VSS.t1339 VSS.t1069 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5061 VDD.t1624 VDD.t1623 VDD.t1624 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5062 VDD.t1622 VDD.t1621 VDD.t1622 VDD.t79 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5063 VSS.t1337 VSS.t1336 VSS.t1337 VSS.t842 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5064 VSS.t1335 VSS.t1334 VSS.t1335 VSS.t1227 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5065 VDD.t1620 VDD.t1619 VDD.t1620 VDD.t547 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5066 VDD.t1618 VDD.t1617 VDD.t1618 VDD.t526 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5067 a_33249_48695.t137 a_33379_34007.t73 a_33249_34067.t37 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5068 VDD.t1616 VDD.t1615 VDD.t1616 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5069 VDD.t1614 VDD.t1612 VDD.t1614 VDD.t1613 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5070 VSS.t1333 VSS.t1332 VSS.t1333 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5071 a_32088_13546# a_30152_10448.t17 VDD.t366 VDD.t304 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5072 VDD.t1611 VDD.t1610 VDD.t1611 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5073 a_84017_n16810.t0 a_71281_n10073.t268 a_83709_n13190# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5074 VDD.t238 a_31699_20742.t213 a_35502_24538.t7 VDD.t37 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5075 VSS.t6 a_35502_25545.t85 a_33249_35053.t112 VSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5076 a_107339_n18620# a_71281_n8397.t280 a_106501_n15905# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5077 a_33249_48695.t197 a_31699_20742.t214 VDD.t239 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5078 VSS.t1331 VSS.t1330 VSS.t1331 VSS.t527 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5079 VDD.t1609 VDD.t1608 VDD.t1609 VDD.t1254 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5080 VDD.t1607 VDD.t1606 VDD.t1607 VDD.t1212 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5081 VSS.t1329 VSS.t1328 VSS.t1329 VSS.t300 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5082 VSS.t1327 VSS.t1326 VSS.t1327 VSS.t620 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5083 a_33249_48695.t196 a_31699_20742.t215 VDD.t240 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5084 VSS.t1325 VSS.t1324 VSS.t1325 VSS.t800 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5085 VDD.t4798 a_83153_10448.t22 a_83683_12380# VDD.t3355 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5086 VDD.t1605 VDD.t1604 VDD.t1605 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5087 a_33249_48695.t195 a_31699_20742.t216 VDD.t241 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5088 VDD.t1603 VDD.t1602 VDD.t1603 VDD.t908 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5089 VDD.t1601 VDD.t1600 VDD.t1601 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5090 VDD.t1599 VDD.t1598 VDD.t1599 VDD.t896 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5091 VSS.t1323 VSS.t1322 VSS.t1323 VSS.t1258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5092 VSS.t1321 VSS.t1319 VSS.t1321 VSS.t1320 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5093 a_106830_10388.t3 a_86903_n14095.t8 a_114516_12380# VDD.t376 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5094 a_32088_11614# a_30152_10448.t18 VDD.t339 VDD.t304 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5095 VDD.t1597 VDD.t1596 VDD.t1597 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5096 VDD.t1595 VDD.t1594 VDD.t1595 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5097 VSS.t1318 VSS.t1317 VSS.t1318 VSS.t536 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5098 VDD.t1593 VDD.t1592 VDD.t1593 VDD.t546 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5099 a_45445_n16904# a_31953_n19727.t294 a_44885_n16904# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5100 VSS.t1316 VSS.t1315 VSS.t1316 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5101 a_60845_n2653# a_50751_n19729.t289 a_60285_n2653# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5102 VSS.t1314 VSS.t1313 VSS.t1314 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5103 VSS.t1312 VSS.t1310 VSS.t1312 VSS.t1311 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5104 VSS.t1309 VSS.t1307 VSS.t1309 VSS.t1308 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5105 VSS.t1306 VSS.t1305 VSS.t1306 VSS.t581 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5106 VSS.t1304 VSS.t1303 VSS.t1304 VSS.t596 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5107 VDD.t1591 VDD.t1590 VDD.t1591 VDD.t1212 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5108 a_33787_n8930# a_31953_n19727.t295 a_32913_n5342.t1 VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5109 VSS.t1302 VSS.t1301 VSS.t1302 VSS.t350 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5110 VDD.t1589 VDD.t1588 VDD.t1589 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5111 a_33249_48695.t82 a_33379_34917.t67 a_33249_35053.t65 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5112 VDD.t1587 VDD.t1586 VDD.t1587 VDD.t30 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5113 a_51711_n6241# a_50751_n19729.t290 a_51151_n4447# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5114 a_67462_n27257# a_45445_n19595.t1 a_44363_n16007.t2 VSS.t412 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5115 a_66551_n16906# a_50751_n19729.t291 a_66029_n16906# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5116 a_31699_20742.t14 a_31699_20742.t13 VDD.t27 VDD.t26 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5117 VSS.t1300 VSS.t1298 VSS.t1300 VSS.t1299 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5118 VSS.t1297 VSS.t1296 VSS.t1297 VSS.t942 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5119 VDD.t1585 VDD.t1584 VDD.t1585 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5120 VDD.t1583 VDD.t1582 VDD.t1583 VDD.t1186 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5121 a_32353_n17801# a_31953_n19727.t296 a_31831_n17801# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5122 VSS.t115 a_31953_n19727.t297 a_44885_n8930# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5123 VDD.t1581 VDD.t1580 VDD.t1581 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5124 VDD.t4839 a_52635_34067.t209 a_52635_49681.t102 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5125 VSS.t1295 VSS.t1294 VSS.t1295 VSS.t839 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5126 VDD.t1579 VDD.t1578 VDD.t1579 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5127 VDD.t1577 VDD.t1576 VDD.t1577 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5128 a_51711_n14215# a_50751_n19729.t292 a_51151_n13318# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5129 VDD.t1575 VDD.t1574 VDD.t1575 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5130 VSS.t1293 VSS.t1291 VSS.t1293 VSS.t1292 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5131 VSS.t1290 VSS.t1289 VSS.t1290 VSS.t495 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5132 VDD.t1573 VDD.t1571 VDD.t1573 VDD.t1572 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5133 VSS.t1288 VSS.t1287 VSS.t1288 VSS.t813 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5134 VDD.t1570 VDD.t1569 VDD.t1570 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5135 VDD.t1568 VDD.t1567 VDD.t1568 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5136 a_60285_n1756# a_50751_n19729.t293 VSS.t270 VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5137 VDD.t1566 VDD.t1565 VDD.t1566 VDD.t1180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5138 a_33249_35053.t95 a_35502_24538.t55 OUT.t5 VSS.t167 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5139 VDD.t1564 VDD.t1563 VDD.t1564 VDD.t1198 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5140 a_52635_48695.t104 a_52635_34067.t210 VDD.t4838 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5141 VDD.t1562 VDD.t1561 VDD.t1562 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5142 a_52635_48695.t23 a_35922_19591.t145 a_52635_34067.t20 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5143 VSS.t1286 VSS.t1285 VSS.t1286 VSS.t913 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5144 VSS.t1284 VSS.t1283 VSS.t1284 VSS.t299 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5145 VDD.t1560 VDD.t1559 VDD.t1560 VDD.t855 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5146 VDD.t1558 VDD.t1557 VDD.t1558 VDD.t1186 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5147 a_36562_12380# a_36162_10388.t20 a_36032_11614.t1 VDD.t3424 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5148 VSS.t1282 VSS.t1281 VSS.t1282 VSS.t765 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5149 VSS.t1280 VSS.t1279 VSS.t1280 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5150 VDD.t1556 VDD.t1555 VDD.t1556 VDD.t526 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5151 VDD.t1554 VDD.t1553 VDD.t1554 VDD.t63 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5152 a_33379_34917.t68 IN_NEG.t1 cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
X5153 a_42442_n34390# a_36032_n35156.t11 a_36162_n36382.t2 VDD.t564 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5154 a_33249_35053.t111 a_35502_25545.t86 VSS.t123 VSS.t11 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5155 VDD.t4837 a_52635_34067.t211 a_52635_48695.t103 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5156 VDD.t1552 VDD.t1550 VDD.t1552 VDD.t1551 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5157 VDD.t1549 VDD.t1548 VDD.t1549 VDD.t61 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5158 a_61484_n28415# a_59558_n29181.t19 VSS.t320 VSS.t314 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5159 a_110225_n6055# a_71281_n8397.t281 a_109695_n9675# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5160 a_39179_n8033# a_31953_n19727.t298 a_38619_n7136# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5161 a_96818_n30339# a_94892_n29181.t19 VSS.t454 VSS.t447 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5162 VDD.t1547 VDD.t1546 VDD.t1547 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5163 VDD.t1545 VDD.t1544 VDD.t1545 VDD.t1180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5164 VDD.t1543 VDD.t1541 VDD.t1543 VDD.t1542 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5165 a_100820_n35156.t0 a_100992_n29313.t0 a_102796_n28415# VSS.t382 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5166 VDD.t1540 VDD.t1539 VDD.t1540 VDD.t1198 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5167 a_52585_n3550# a_50751_n19729.t294 a_52063_n3550# VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5168 VDD.t1538 VDD.t1537 VDD.t1538 VDD.t836 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5169 a_54019_n8035# a_50751_n19729.t295 a_53497_n8035# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5170 VDD.t1536 VDD.t1535 VDD.t1536 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5171 a_32353_n6239# a_31953_n19727.t299 a_31831_n7136# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5172 a_54579_n4447# a_50751_n19729.t296 a_54019_n3550# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5173 VSS.t1278 VSS.t1277 VSS.t1278 VSS.t533 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5174 VSS.t1276 VSS.t1275 VSS.t1276 VSS.t858 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5175 VDD.t1534 VDD.t1533 VDD.t1534 VDD.t81 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5176 VSS.t1274 VSS.t1273 VSS.t1274 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5177 a_31953_n19727.t21 a_31953_n19727.t20 VSS.t68 VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5178 VDD.t1532 VDD.t1531 VDD.t1532 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5179 VSS.t1272 VSS.t1271 VSS.t1272 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5180 a_33249_48695.t194 a_31699_20742.t217 VDD.t242 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5181 VDD.t1530 VDD.t1529 VDD.t1530 VDD.t390 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5182 a_79151_n27257# a_77225_n29181.t20 VSS.t394 VSS.t387 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5183 OUT.t108 a_33379_34917.t0 cap_mim_2f0_m4m5_noshield c_width=9.8u c_length=9.8u
X5184 a_112199_n9675# a_71281_n8397.t282 a_111631_n9675# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5185 a_49755_10448# a_47819_10448.t18 VDD.t516 VDD.t498 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5186 VSS.t1270 VSS.t1269 VSS.t1270 VSS.t780 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5187 VDD.t1528 VDD.t1527 VDD.t1528 VDD.t424 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5188 VSS.t1268 VSS.t1267 VSS.t1268 VSS.t20 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X5189 VSS.t1266 VSS.t1265 VSS.t1266 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5190 a_33249_48695.t83 a_33379_34917.t69 a_33249_35053.t66 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5191 a_94537_n8770# a_71281_n10073.t269 a_93969_n8770# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5192 VDD.t1526 VDD.t1525 VDD.t1526 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5193 VDD.t1524 VDD.t1523 VDD.t1524 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5194 VSS.t1264 VSS.t1263 VSS.t1264 VSS.t819 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5195 a_63161_n5344.t1 a_64243_n1756.t1 a_66058_5639# VSS.t411 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5196 a_71342_7563.t3 a_71496_10388.t21 a_71896_13546# VDD.t489 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5197 a_89163_10388.t5 a_81205_n14095.t7 a_96849_12380# VDD.t503 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5198 VDD.t1522 VDD.t1521 VDD.t1522 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5199 VDD.t1520 VDD.t1519 VDD.t1520 VDD.t804 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5200 a_51151_n16906# a_50751_n19729.t297 a_50629_n17803# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5201 VDD.t1518 VDD.t1516 VDD.t1518 VDD.t1517 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5202 a_84017_n17715.t1 a_83325_4421.t1 a_95443_10448# VDD.t501 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5203 VDD.t506 a_30152_11614.t17 a_37934_5639# VSS.t323 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5204 VDD.t1515 VDD.t1514 VDD.t1515 VDD.t493 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5205 VSS.t1262 VSS.t1260 VSS.t1262 VSS.t1261 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5206 a_42047_n19595# a_31953_n19727.t300 a_41487_n18698# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5207 a_83725_n27257# a_83325_n29313.t2 a_83153_n35156.t11 VSS.t367 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5208 VDD.t1513 VDD.t1512 VDD.t1513 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5209 a_77747_5639# a_77225_4481.t19 a_71496_10388.t3 VSS.t336 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5210 a_52635_48695.t22 a_35922_19591.t146 a_52635_34067.t23 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5211 VDD.t1511 VDD.t1510 VDD.t1511 VDD.t433 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5212 VDD.t1509 VDD.t1507 VDD.t1509 VDD.t1508 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5213 VSS.t1259 VSS.t1257 VSS.t1259 VSS.t1258 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5214 a_90245_n6960# a_71281_n10073.t270 a_89407_n4245# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5215 a_52585_n19597# a_50751_n19729.t298 VSS.t271 VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5216 a_107198_n28415# a_100820_n36322.t18 VDD.t542 VSS.t352 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5217 VSS.t1256 VSS.t1255 VSS.t1256 VSS.t171 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5218 VDD.t1506 VDD.t1505 VDD.t1506 VDD.t422 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5219 VSS.t1254 VSS.t1253 VSS.t1254 VSS.t427 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5220 a_52635_49681.t64 a_35922_19591.t147 OUT.t43 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5221 VSS.t1252 VSS.t1251 VSS.t1252 VSS.t328 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5222 VSS.t397 a_71496_10388.t22 a_71896_11614# VDD.t489 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5223 a_59411_n8932# a_50751_n19729.t299 a_58851_n8932# VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5224 VDD.t1504 VDD.t1503 VDD.t1504 VDD.t323 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5225 VDD.t1502 VDD.t1501 VDD.t1502 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5226 a_52635_48695.t102 a_52635_34067.t212 VDD.t4836 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5227 VSS.t1250 VSS.t1248 VSS.t1250 VSS.t1249 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X5228 a_33249_48695.t84 a_33379_34917.t70 a_33249_35053.t67 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5229 VDD.t1500 VDD.t1499 VDD.t1500 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5230 VDD.t1498 VDD.t1496 VDD.t1498 VDD.t1497 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5231 VDD.t1495 VDD.t1494 VDD.t1495 VDD.t530 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5232 VDD.t1493 VDD.t1491 VDD.t1493 VDD.t1492 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5233 a_52635_48695.t101 a_52635_34067.t213 VDD.t4835 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5234 a_48951_4481.t1 a_47991_5507.t0 a_48391_7563# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5235 VDD.t1490 VDD.t1488 VDD.t1490 VDD.t1489 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5236 a_66551_n8035# a_50751_n19729.t300 a_66029_n8035# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5237 a_32128_5639# a_30324_4421.t0 a_31284_4481.t2 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5238 a_88271_n1530# a_71281_n10073.t271 a_87433_n1530# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5239 VSS.t1247 VSS.t1246 VSS.t1247 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5240 VDD.t1487 VDD.t1486 VDD.t1487 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5241 VSS.t1245 VSS.t1244 VSS.t1245 VSS.t286 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5242 a_33249_48695.t85 a_33379_34917.t71 a_33249_35053.t68 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5243 VSS.t1243 VSS.t1241 VSS.t1243 VSS.t1242 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X5244 VSS.t1240 VSS.t1239 VSS.t1240 VSS.t171 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5245 VSS.t1238 VSS.t1237 VSS.t1238 VSS.t816 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5246 VSS.t1236 VSS.t1235 VSS.t1236 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5247 a_60080_7563# a_59558_4481.t18 a_53829_10388.t1 VSS.t313 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5248 VDD.t1485 VDD.t1483 VDD.t1485 VDD.t1484 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5249 VSS.t1234 VSS.t1233 VSS.t1234 VSS.t253 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5250 VSS.t1232 VSS.t1231 VSS.t1232 VSS.t643 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5251 VDD.t1482 VDD.t1481 VDD.t1482 VDD.t1115 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5252 a_77225_4481.t10 a_65658_4421.t2 a_79182_13546# VDD.t1843 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5253 VSS.t1230 VSS.t1229 VSS.t1230 VSS.t777 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5254 a_100820_11614.t3 a_100820_10448.t18 a_102756_12380# VDD.t324 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5255 a_33249_48695.t138 a_33379_34007.t74 a_33249_34067.t36 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5256 VDD.t1480 VDD.t1479 VDD.t1480 VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5257 a_53829_10388.t3 a_59558_4481.t19 a_61484_4481# VSS.t312 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5258 VSS.t1228 VSS.t1226 VSS.t1228 VSS.t1227 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5259 VDD.t1478 VDD.t1477 VDD.t1478 VDD.t1130 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5260 VSS.t1225 VSS.t1224 VSS.t1225 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5261 a_33249_34067.t35 a_33379_34007.t75 a_33249_48695.t139 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5262 VDD.t1476 VDD.t1475 VDD.t1476 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5263 a_35502_24538.t6 a_31699_20742.t218 VDD.t243 VDD.t35 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5264 a_40613_n13316# a_31953_n19727.t301 a_40053_n13316# VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5265 a_65677_n17803# a_50751_n19729.t301 a_66551_n16009# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5266 VSS.t1223 VSS.t1222 VSS.t1223 VSS.t428 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5267 a_35502_24538.t5 a_31699_20742.t219 VDD.t244 VDD.t26 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5268 a_52635_48695.t100 a_52635_34067.t214 VDD.t4834 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5269 VDD.t4833 a_52635_34067.t215 a_52635_48695.t99 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5270 VSS.t1221 VSS.t1220 VSS.t1221 VSS.t861 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5271 a_100820_n35156.t4 a_100820_n35156.t3 a_102756_n36322# VDD.t528 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5272 a_35502_25545.t17 a_31699_20742.t220 VDD.t245 VDD.t15 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5273 a_40053_n14213# a_31953_n19727.t302 a_39531_n14213# VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5274 a_61484_6405# a_59558_4481.t20 VSS.t407 VSS.t314 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5275 VSS.t1219 VSS.t1218 VSS.t1219 VSS.t620 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5276 VSS.t1217 VSS.t1216 VSS.t1217 VSS.t695 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5277 VDD.t1474 VDD.t1473 VDD.t1474 VDD.t1115 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5278 VSS.t1215 VSS.t1214 VSS.t1215 VSS.t692 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5279 a_77225_4481.t9 a_65658_4421.t2 a_79182_11614# VDD.t1843 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5280 a_39179_n18698# a_31953_n19727.t303 a_38619_n18698# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5281 VSS.t1213 VSS.t1212 VSS.t1213 VSS.t797 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5282 a_33249_48695.t193 a_31699_20742.t221 VDD.t246 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5283 a_52635_49681.t65 a_35922_19591.t148 OUT.t42 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5284 VDD.t1472 VDD.t1471 VDD.t1472 VDD.t332 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5285 VDD.t1470 VDD.t1469 VDD.t1470 VDD.t73 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5286 VDD.t1468 VDD.t1467 VDD.t1468 VDD.t329 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5287 VDD.t1466 VDD.t1465 VDD.t1466 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5288 VDD.t1464 VDD.t1463 VDD.t1464 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5289 a_44363_n16007.t1 a_65658_n29313.t0 a_66058_n29181# VSS.t411 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5290 VDD.t1462 VDD.t1461 VDD.t1462 VDD.t1130 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5291 VSS.t1211 VSS.t1210 VSS.t1211 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5292 VDD.t1460 VDD.t1459 VDD.t1460 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5293 VDD.t1458 VDD.t1457 VDD.t1458 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5294 VDD.t1456 VDD.t1455 VDD.t1456 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5295 a_87433_n8770# a_71281_n10073.t272 VDD.t385 VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5296 VSS.t1209 VSS.t1208 VSS.t1209 VSS.t174 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5297 VSS.t1207 VSS.t1206 VSS.t1207 VSS.t681 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5298 VSS.t1205 VSS.t1204 VSS.t1205 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5299 a_60285_n18700# a_50751_n19729.t302 a_59763_n18700# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5300 VDD.t1454 VDD.t1453 VDD.t1454 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5301 VDD.t1452 VDD.t1451 VDD.t1452 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5302 VDD.t1450 VDD.t1449 VDD.t1450 VDD.t438 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5303 a_38619_n16007# a_31953_n19727.t304 a_38097_n16007.t0 VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5304 VSS.t1203 VSS.t1202 VSS.t1203 VSS.t1162 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5305 VDD.t1448 VDD.t1447 VDD.t1448 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5306 VSS.t1201 VSS.t1200 VSS.t1201 VSS.t259 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5307 VSS.t1199 VSS.t1198 VSS.t1199 VSS.t285 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5308 a_113081_n29181# a_112559_n29181.t5 a_112559_n29181.t6 VSS.t415 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5309 VSS.t1197 VSS.t1196 VSS.t1197 VSS.t822 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X5310 VSS.t1195 VSS.t1194 VSS.t1195 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5311 VSS.t1193 VSS.t1192 VSS.t1193 VSS.t218 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5312 VDD.t1446 VDD.t1444 VDD.t1446 VDD.t1445 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5313 VDD.t1443 VDD.t1441 VDD.t1443 VDD.t1442 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5314 VSS.t1191 VSS.t1190 VSS.t1191 VSS.t413 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5315 VDD.t1440 VDD.t1439 VDD.t1440 VDD.t804 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5316 VDD.t1438 VDD.t1437 VDD.t1438 VDD.t73 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5317 VDD.t537 a_100820_n35156.t18 a_101350_n36322# VDD.t535 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5318 a_85089_12380# a_83153_10448.t23 VDD.t4799 VDD.t1445 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5319 VDD.t1436 VDD.t1435 VDD.t1436 VDD.t1084 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5320 VSS.t1189 VSS.t1188 VSS.t1189 VSS.t177 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5321 a_33249_48695.t192 a_31699_20742.t222 VDD.t247 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5322 VDD.t1434 VDD.t1433 VDD.t1434 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5323 VSS.t1187 VSS.t1186 VSS.t1187 VSS.t337 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5324 VSS.t344 a_77225_4481.t20 a_77747_7563# VSS.t341 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5325 VSS.t1185 VSS.t1184 VSS.t1185 VSS.t800 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5326 a_47991_5507.t0 a_47819_11614.t18 a_54197_5639# VSS.t327 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5327 VSS.t1183 VSS.t1182 VSS.t1183 VSS.t658 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5328 a_54019_n3550# a_50751_n19729.t303 a_53497_n3550# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5329 VSS.t224 a_50751_n19729.t22 a_50751_n19729.t23 VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5330 a_33249_48695.t191 a_31699_20742.t223 VDD.t248 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5331 VSS.t1181 VSS.t1180 VSS.t1181 VSS.t142 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5332 a_95105_n19525# a_71281_n10073.t273 a_94537_n19525# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5333 a_33249_34067.t34 a_33379_34007.t76 a_33249_48695.t140 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5334 VSS.t1179 VSS.t1178 VSS.t1179 VSS.t676 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5335 VSS.t1177 VSS.t1176 VSS.t1177 VSS.t738 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5336 a_41660_19698# a_35502_24538.t56 a_41100_19698# VSS.t189 nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X5337 a_90245_n20430# a_71281_n10073.t274 a_89407_n19525# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5338 VSS.t1175 VSS.t1174 VSS.t1175 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5339 a_107339_n3340# a_71281_n8397.t283 a_106501_n3340# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5340 VDD.t1432 VDD.t1431 VDD.t1432 VDD.t19 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5341 VDD.t1430 VDD.t1429 VDD.t1430 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5342 VDD.t1428 VDD.t1426 VDD.t1428 VDD.t1427 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5343 VDD.t1425 VDD.t1424 VDD.t1425 VDD.t1084 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5344 VDD.t1423 VDD.t1421 VDD.t1423 VDD.t1422 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5345 a_101641_n15000# a_71281_n8397.t284 a_100803_n14095# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5346 VSS.t1173 VSS.t1172 VSS.t1173 VSS.t686 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5347 a_45706_23609# a_35922_19591.t149 a_45138_23609# VDD.t401 pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X5348 a_48313_n13316# a_31953_n19727.t305 a_47753_n12419# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5349 VDD.t1420 VDD.t1419 VDD.t1420 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5350 VDD.t1418 VDD.t1417 VDD.t1418 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5351 a_33249_34067.t116 a_35502_25545.t87 VSS.t131 VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5352 a_36562_n36322# a_36162_n36382.t21 a_36032_n36322.t1 VDD.t683 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5353 a_47753_n8930# a_31953_n19727.t306 VSS.t116 VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5354 VDD.t1416 VDD.t1415 VDD.t1416 VDD.t1209 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5355 VSS.t395 a_77225_n29181.t21 a_77747_n29181# VSS.t390 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5356 a_41487_n19595# a_31953_n19727.t307 VSS.t117 VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5357 VSS.t1171 VSS.t1170 VSS.t1171 VSS.t13 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5358 VDD.t1414 VDD.t1413 VDD.t1414 VDD.t1052 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5359 a_58851_n13318# a_50751_n19729.t304 a_58329_n14215# VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5360 a_42047_n8930# a_31953_n19727.t308 a_41487_n8033# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5361 VDD.t1412 VDD.t1410 VDD.t1412 VDD.t1411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5362 VDD.t1409 VDD.t1407 VDD.t1409 VDD.t1408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5363 VSS.t1169 VSS.t1168 VSS.t1169 VSS.t207 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5364 VSS.t1167 VSS.t1166 VSS.t1167 VSS.t99 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5365 a_88839_n19525# a_71281_n10073.t275 a_88271_n19525# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5366 VSS.t1165 VSS.t1164 VSS.t1165 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5367 VSS.t1163 VSS.t1161 VSS.t1163 VSS.t1162 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5368 VSS.t1160 VSS.t1159 VSS.t1160 VSS.t753 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5369 a_106676_4481.t0 a_100820_11614.t20 a_108602_7563# VSS.t151 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5370 a_30324_4421.t0 a_30152_11614.t18 a_36530_7563# VSS.t325 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5371 a_94537_n7865# a_71281_n10073.t276 a_93969_n7865# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5372 a_89715_n17715.t0 a_86903_n14095.t9 a_113110_13546# VDD.t374 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5373 VDD.t1406 VDD.t1405 VDD.t1406 VDD.t551 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5374 a_33249_48695.t141 a_33379_34007.t77 a_33249_34067.t33 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5375 VSS.t1158 VSS.t1157 VSS.t1158 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5376 VSS.t1156 VSS.t1155 VSS.t1156 VSS.t211 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5377 VDD.t249 a_31699_20742.t224 a_35502_24538.t4 VDD.t37 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5378 a_33249_48695.t190 a_31699_20742.t225 VDD.t250 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5379 a_52635_48695.t98 a_52635_34067.t216 VDD.t4832 VDD.t390 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5380 VSS.t67 a_31953_n19727.t18 a_31953_n19727.t19 VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5381 VSS.t1154 VSS.t1153 VSS.t1154 VSS.t709 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5382 VDD.t1404 VDD.t1403 VDD.t1404 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5383 VSS.t1152 VSS.t1151 VSS.t1152 VSS.t1039 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5384 VSS.t1150 VSS.t1149 VSS.t1150 VSS.t160 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5385 VDD.t1402 VDD.t1401 VDD.t1402 VDD.t1052 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5386 VDD.t251 a_31699_20742.t226 a_35502_25545.t4 VDD.t28 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5387 a_66016_n34390# a_65486_n35156.t21 a_65486_n36322.t2 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5388 VDD.t1400 VDD.t1399 VDD.t1400 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5389 VDD.t1398 VDD.t1397 VDD.t1398 VDD.t928 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5390 VSS.t1148 VSS.t1147 VSS.t1148 VSS.t620 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5391 a_71342_n27257.t1 a_65486_n36322.t22 a_73268_n30339# VSS.t154 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5392 VDD.t1396 VDD.t1395 VDD.t1396 VDD.t1055 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5393 a_51711_n12421.t1 a_50751_n19729.t305 a_51151_n12421# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5394 VSS.t1146 VSS.t1145 VSS.t1146 VSS.t33 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5395 VSS.t1144 VSS.t1143 VSS.t1144 VSS.t183 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5396 a_61515_12380# a_53699_11614.t9 a_60677_10448.t1 VDD.t495 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5397 VSS.t1142 VSS.t1141 VSS.t1142 VSS.t573 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5398 VSS.t1140 VSS.t1139 VSS.t1140 VSS.t281 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5399 a_107339_n15000# a_71281_n8397.t285 a_106501_n14095# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5400 a_89715_n17715.t1 a_86903_n14095.t10 a_113110_11614# VDD.t374 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5401 VDD.t1394 VDD.t1393 VDD.t1394 VDD.t512 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5402 VSS.t1138 VSS.t1137 VSS.t1138 VSS.t689 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5403 a_52635_34067.t4 a_35502_24538.t57 a_33249_34067.t3 VSS.t187 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5404 VSS.t1136 VSS.t1135 VSS.t1136 VSS.t768 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X5405 a_33249_48695.t142 a_33379_34007.t78 a_33249_34067.t32 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5406 a_44885_n19595# a_31953_n19727.t309 a_44363_n19595# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5407 VSS.t1134 VSS.t1133 VSS.t1134 VSS.t649 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5408 a_66551_n3550# a_50751_n19729.t306 a_66029_n3550# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5409 VDD.t1392 VDD.t1391 VDD.t1392 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5410 VSS.t1132 VSS.t1130 VSS.t1132 VSS.t1131 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5411 VSS.t1129 VSS.t1128 VSS.t1129 VSS.t282 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5412 VSS.t1127 VSS.t1126 VSS.t1127 VSS.t609 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5413 a_52635_48695.t21 a_35922_19591.t150 a_52635_34067.t49 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5414 a_83709_n9675# a_71281_n10073.t277 a_83141_n9675# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5415 a_32128_n30339# a_30324_n29313.t0 a_31284_n30339.t1 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5416 VDD.t1390 VDD.t1389 VDD.t1390 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5417 VDD.t1388 VDD.t1387 VDD.t1388 VDD.t301 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5418 a_53675_n30339.t0 a_47819_n36322.t21 a_55601_n27257# VSS.t328 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5419 VSS.t1125 VSS.t1124 VSS.t1125 VSS.t676 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5420 VDD.t1386 VDD.t1385 VDD.t1386 VDD.t1055 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5421 a_111631_n8770# a_71281_n8397.t286 a_111063_n8770# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5422 VSS.t1123 VSS.t1122 VSS.t1123 VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5423 VSS.t1121 VSS.t1120 VSS.t1121 VSS.t150 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5424 a_33249_48695.t189 a_31699_20742.t227 VDD.t252 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5425 a_48313_n7136# a_31953_n19727.t310 a_47753_n6239# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5426 a_89009_7563.t2 a_89163_10388.t19 a_89563_13546# VDD.t558 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5427 VDD.t1384 VDD.t1383 VDD.t1384 VDD.t913 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5428 VDD.t1382 VDD.t1380 VDD.t1382 VDD.t1381 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5429 a_33249_48695.t86 a_33379_34917.t72 a_33249_35053.t69 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5430 VSS.t435 a_53829_10388.t22 a_54229_12380# VDD.t1408 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5431 a_30152_11614.t5 a_30152_10448.t19 a_32088_12380# VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5432 a_83709_n18620# a_71281_n10073.t278 a_83141_n18620# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5433 VDD.t1379 VDD.t1378 VDD.t1379 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5434 VDD.t1377 VDD.t1375 VDD.t1377 VDD.t1376 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5435 VDD.t253 a_31699_20742.t228 a_33249_48695.t188 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5436 VSS.t1119 VSS.t1118 VSS.t1119 VSS.t614 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5437 VDD.t303 a_30152_10448.t20 a_30682_10448# VDD.t13 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5438 VDD.t1374 VDD.t1372 VDD.t1374 VDD.t1373 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5439 a_52585_n2653# a_50751_n19729.t307 a_52063_n3550# VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5440 VSS.t1117 VSS.t1115 VSS.t1117 VSS.t1116 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5441 VDD.t1371 VDD.t1370 VDD.t1371 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5442 a_96849_10448# a_81205_n14095.t8 a_84017_n17715.t1 VDD.t502 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5443 VDD.t1369 VDD.t1367 VDD.t1369 VDD.t1368 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5444 a_108602_7563# a_100820_11614.t21 a_100992_4421.t0 VSS.t147 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5445 a_36530_7563# a_30152_11614.t19 a_36008_7563.t3 VSS.t326 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5446 VSS.t1114 VSS.t1113 VSS.t1114 VSS.t328 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5447 VDD.t1366 VDD.t1365 VDD.t1366 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5448 a_85129_n28415# a_83325_n29313.t0 a_31831_n5342.t0 VSS.t278 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5449 a_54579_n2653# a_50751_n19729.t308 a_54019_n2653# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5450 a_32353_n5342# a_31953_n19727.t311 a_31831_n5342.t2 VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5451 a_31699_20742.t12 a_31699_20742.t11 VDD.t25 VDD.t15 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5452 VDD.t254 a_31699_20742.t229 a_33249_48695.t187 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5453 VSS.t1112 VSS.t1111 VSS.t1112 VSS.t655 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5454 a_33249_34067.t2 a_35502_24538.t58 a_52635_34067.t4 VSS.t167 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5455 VDD.t1364 VDD.t1363 VDD.t1364 VDD.t500 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5456 VSS.t1110 VSS.t1108 VSS.t1110 VSS.t1109 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5457 a_81735_n6960# a_71281_n10073.t279 a_81205_n7865# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5458 a_36530_n30339# a_30152_n36322.t21 a_36008_n30339.t3 VSS.t326 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5459 a_31953_n19727.t17 a_31953_n19727.t16 VSS.t65 VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5460 VSS.t361 a_89163_10388.t20 a_89563_11614# VDD.t558 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5461 VDD.t1362 VDD.t1361 VDD.t1362 VDD.t404 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5462 VSS.t1107 VSS.t1106 VSS.t1107 VSS.t381 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5463 a_75602_n4019# a_71266_n4019.t0 VDD.t4778 VDD.t695 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X5464 VDD.t1360 VDD.t1359 VDD.t1360 VDD.t525 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5465 VSS.t1105 VSS.t1104 VSS.t1105 VSS.t646 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5466 VDD.t1358 VDD.t1356 VDD.t1358 VDD.t1357 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5467 VDD.t1355 VDD.t1354 VDD.t1355 VDD.t1018 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5468 a_98829_n6960# a_71281_n8397.t287 a_98299_n7865# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5469 a_33249_34067.t115 a_35502_25545.t88 VSS.t130 VSS.t7 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5470 VDD.t1353 VDD.t1351 VDD.t1353 VDD.t1352 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5471 VSS.t1103 VSS.t1102 VSS.t1103 VSS.t643 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5472 VSS.t1101 VSS.t1100 VSS.t1101 VSS.t762 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5473 VDD.t1350 VDD.t1349 VDD.t1350 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5474 VDD.t429 a_71281_n8397.t8 a_71281_n8397.t9 VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5475 VSS.t1099 VSS.t1098 VSS.t1099 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5476 VDD.t1348 VDD.t1347 VDD.t1348 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5477 a_52635_34067.t42 a_35922_19591.t151 a_52635_48695.t20 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5478 VDD.t1346 VDD.t1345 VDD.t1346 VDD.t405 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5479 VDD.t1344 VDD.t1343 VDD.t1344 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5480 VSS.t1097 VSS.t1096 VSS.t1097 VSS.t652 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5481 a_47819_11614.t6 a_47991_5507.t0 a_49795_4481# VSS.t282 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5482 a_89531_n28415# a_83153_n36322.t20 VDD.t4789 VSS.t459 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5483 a_39179_n8930.t1 a_100820_n36322.t19 a_107198_n29181# VSS.t353 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5484 VDD.t1342 VDD.t1340 VDD.t1342 VDD.t1341 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5485 VDD.t255 a_31699_20742.t230 a_33249_48695.t186 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5486 VDD.t4831 a_52635_34067.t217 a_52635_49681.t101 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5487 VDD.t1339 VDD.t1338 VDD.t1339 VDD.t400 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5488 a_93131_n18620# a_71281_n10073.t280 a_92601_n19525# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5489 a_87433_n7865# a_71281_n10073.t281 a_86903_n7865# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5490 VDD.t1337 VDD.t1335 VDD.t1337 VDD.t1336 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5491 VDD.t1334 VDD.t1333 VDD.t1334 VDD.t1018 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5492 a_88271_n18620# a_71281_n10073.t282 a_87433_n18620# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5493 VDD.t1332 VDD.t1331 VDD.t1332 VDD.t501 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5494 VDD.t1330 VDD.t1329 VDD.t1330 VDD.t50 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5495 VDD.t1328 VDD.t1327 VDD.t1328 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5496 a_63683_n18700# a_50751_n19729.t309 a_63161_n19597# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5497 a_42442_n36322# a_36032_n35156.t12 a_36162_n36382.t0 VDD.t564 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5498 a_73302_n34390# a_71496_n36382.t16 VSS.t369 VDD.t2814 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5499 VSS.t1095 VSS.t1094 VSS.t1095 VSS.t410 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5500 VSS.t1093 VSS.t1092 VSS.t1093 VSS.t981 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5501 a_49795_6405# a_47991_5507.t2 a_48951_4481.t1 VSS.t281 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5502 VDD.t1326 VDD.t1324 VDD.t1326 VDD.t1325 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5503 VSS.t1091 VSS.t1090 VSS.t1091 VSS.t558 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5504 a_38097_n16007.t1 a_39179_n19595.t0 a_48391_n28415# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5505 VDD.t4830 a_52635_34067.t218 a_52635_48695.t97 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5506 VDD.t1323 VDD.t1322 VDD.t1323 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5507 a_41100_19698# a_35502_24538.t59 a_40578_19075# VSS.t184 nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X5508 VDD.t1321 VDD.t1320 VDD.t1321 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5509 VSS.t1089 VSS.t1088 VSS.t1089 VSS.t638 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5510 a_44885_n4445# a_31953_n19727.t312 a_44363_n4445# VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5511 a_100235_n13190# a_71281_n8397.t288 a_99667_n13190# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5512 a_95105_n9675# a_71281_n10073.t283 a_94537_n9675# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5513 VSS.t1087 VSS.t1086 VSS.t1087 VSS.t418 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5514 VSS.t1085 VSS.t1084 VSS.t1085 VSS.t330 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5515 VSS.t1083 VSS.t1081 VSS.t1083 VSS.t1082 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X5516 a_57417_n8035# a_50751_n19729.t310 a_56895_n8932# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5517 a_31953_n19727.t15 a_31953_n19727.t14 VSS.t64 VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5518 VSS.t1080 VSS.t1079 VSS.t1080 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5519 VDD.t1319 VDD.t1318 VDD.t1319 VDD.t323 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5520 VDD.t1317 VDD.t1316 VDD.t1317 VDD.t50 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5521 a_37934_n29181# a_30152_n36322.t22 a_30324_n30399.t1 VSS.t324 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5522 a_47753_n13316# a_31953_n19727.t313 a_47231_n14213# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5523 VDD.t1315 VDD.t1314 VDD.t1315 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5524 VDD.t1313 VDD.t1312 VDD.t1313 VDD.t968 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5525 VSS.t1078 VSS.t1077 VSS.t1078 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5526 VDD.t1311 VDD.t1310 VDD.t1311 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5527 a_107339_n3340# a_71281_n8397.t289 a_106501_n2435# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5528 VSS.t1076 VSS.t1075 VSS.t1076 VSS.t800 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5529 VSS.t1074 VSS.t1073 VSS.t1074 VSS.t26 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5530 VDD.t1309 VDD.t1308 VDD.t1309 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5531 a_33249_48695.t185 a_31699_20742.t231 VDD.t256 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5532 VDD.t1307 VDD.t1306 VDD.t1307 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5533 a_48391_4481# a_47991_4421.t2 a_47819_10448.t1 VSS.t284 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5534 VDD.t1305 VDD.t1304 VDD.t1305 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5535 a_42047_n4445# a_31953_n19727.t314 a_41487_n3548# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5536 VDD.t1303 VDD.t1301 VDD.t1303 VDD.t1302 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5537 VSS.t1072 VSS.t1071 VSS.t1072 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5538 VDD.t1300 VDD.t1299 VDD.t1300 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5539 VSS.t1070 VSS.t1068 VSS.t1070 VSS.t1069 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5540 a_98829_n13190# a_71281_n8397.t290 a_98299_n16810# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5541 a_54019_n16906# a_50751_n19729.t311 a_53497_n16906# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5542 a_33249_48695.t184 a_31699_20742.t232 VDD.t257 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5543 a_93131_n6960# a_71281_n10073.t284 a_92601_n7865# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5544 VSS.t1067 VSS.t1066 VSS.t1067 VSS.t617 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5545 VDD.t4829 a_52635_34067.t219 a_52635_48695.t96 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5546 VDD.t1298 VDD.t1297 VDD.t1298 VDD.t433 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5547 VDD.t1296 VDD.t1295 VDD.t1296 VDD.t968 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5548 VDD.t419 a_100820_10448.t19 a_101350_13546# VDD.t301 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5549 VSS.t1065 VSS.t1064 VSS.t1065 VSS.t251 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5550 a_31953_n19727.t13 a_31953_n19727.t12 VSS.t62 VSS.t61 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5551 VDD.t258 a_31699_20742.t233 a_33249_48695.t183 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5552 a_67111_n15112# a_50751_n19729.t312 a_66551_n15112# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5553 a_36162_10388.t7 a_36032_11614.t10 a_43848_10448# VDD.t290 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5554 VDD.t1294 VDD.t1292 VDD.t1294 VDD.t1293 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5555 VDD.t1291 VDD.t1290 VDD.t1291 VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5556 a_105365_n13190# a_71281_n8397.t291 a_104527_n13190# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5557 VSS.t1063 VSS.t1062 VSS.t1063 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5558 VDD.t1289 VDD.t1288 VDD.t1289 VDD.t422 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5559 a_65117_n19597# a_50751_n19729.t313 VSS.t272 VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5560 a_35502_25545.t18 a_31699_20742.t234 VDD.t259 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5561 VDD.t1287 VDD.t1286 VDD.t1287 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5562 VSS.t1061 VSS.t1060 VSS.t1061 VSS.t506 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5563 VSS.t1059 VSS.t1058 VSS.t1059 VSS.t503 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5564 VDD.t1285 VDD.t1284 VDD.t1285 VDD.t1145 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5565 VSS.t1057 VSS.t1056 VSS.t1057 VSS.t555 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5566 VDD.t1283 VDD.t1282 VDD.t1283 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5567 VDD.t1281 VDD.t1280 VDD.t1281 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5568 a_59411_n19597# a_50751_n19729.t314 a_58851_n19597# VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5569 VDD.t418 a_100820_10448.t20 a_101350_11614# VDD.t301 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5570 VDD.t1279 VDD.t1278 VDD.t1279 VDD.t404 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5571 VSS.t1055 VSS.t1054 VSS.t1055 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5572 a_33249_35053.t102 a_35502_24538.t60 OUT.t4 VSS.t187 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5573 a_33249_48695.t87 a_33379_34917.t73 a_33249_35053.t70 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5574 a_33249_48695.t143 a_33379_34007.t79 a_33249_34067.t31 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5575 VSS.t1053 VSS.t1052 VSS.t1053 VSS.t503 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5576 VSS.t1051 VSS.t1050 VSS.t1051 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5577 VSS.t1049 VSS.t1048 VSS.t1049 VSS.t495 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5578 VSS.t1047 VSS.t1046 VSS.t1047 VSS.t942 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5579 VDD.t1277 VDD.t1276 VDD.t1277 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5580 VDD.t1275 VDD.t1274 VDD.t1275 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5581 VSS.t1045 VSS.t1044 VSS.t1045 VSS.t839 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5582 a_35502_24538.t3 a_31699_20742.t235 VDD.t260 VDD.t35 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5583 VDD.t1273 VDD.t1272 VDD.t1273 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5584 a_75585_n8397# I1N.t14 VSS.t309 VSS.t303 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X5585 a_45445_n12419# a_31953_n19727.t315 a_44885_n12419# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5586 a_52635_49681.t66 a_35922_19591.t152 OUT.t41 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5587 VDD.t1271 VDD.t1270 VDD.t1271 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5588 VSS.t1043 VSS.t1041 VSS.t1043 VSS.t1042 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5589 VSS.t1040 VSS.t1038 VSS.t1040 VSS.t1039 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5590 VSS.t455 a_94892_n29181.t20 a_95414_n29181# VSS.t450 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5591 a_43817_n27257# a_41891_n29181.t21 VSS.t378 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5592 a_112199_n3340# a_71281_n8397.t292 a_111631_n3340# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5593 a_90935_6405# a_83153_11614.t20 a_51711_n12421.t0 VSS.t401 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5594 a_52635_48695.t95 a_52635_34067.t220 VDD.t4828 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5595 VDD.t1269 VDD.t1267 VDD.t1269 VDD.t1268 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5596 a_39179_n1754# a_31953_n19727.t316 a_38619_n1754# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5597 VDD.t1266 VDD.t1264 VDD.t1266 VDD.t1265 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5598 a_49795_n27257# a_39179_n19595.t0 a_38097_n16007.t2 VSS.t281 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5599 VSS.t1037 VSS.t1036 VSS.t1037 VSS.t581 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5600 a_32353_n13316# a_31953_n19727.t317 a_31831_n13316# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5601 VSS.t1035 VSS.t1034 VSS.t1035 VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5602 VDD.t1263 VDD.t1262 VDD.t1263 VDD.t933 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5603 a_71281_n8397.t7 a_71281_n8397.t6 VDD.t427 VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5604 VDD.t1261 VDD.t1260 VDD.t1261 VDD.t73 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5605 a_54019_n2653# a_50751_n19729.t315 a_53497_n3550# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5606 VSS.t1033 VSS.t1032 VSS.t1033 VSS.t167 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5607 a_104527_n6960# a_71281_n8397.t293 a_103997_n7865# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5608 VDD.t1259 VDD.t1258 VDD.t1259 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5609 a_89033_13546.t3 a_106830_10388.t19 a_108636_13546# VDD.t526 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5610 VSS.t1031 VSS.t1029 VSS.t1031 VSS.t1030 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5611 a_112199_n15000# a_71281_n8397.t294 a_111631_n15000# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5612 a_82573_n8770# a_71281_n10073.t285 a_81735_n8770# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5613 a_111631_n7865# a_71281_n8397.t295 a_111063_n7865# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5614 VSS.t1028 VSS.t1027 VSS.t1028 VSS.t61 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5615 VSS.t1026 VSS.t1025 VSS.t1026 VSS.t530 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5616 a_52635_34067.t45 a_35922_19591.t153 a_52635_48695.t19 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5617 VSS.t1024 VSS.t1023 VSS.t1024 VSS.t558 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5618 a_66058_6405# a_65658_4421.t0 a_65486_10448.t10 VSS.t410 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5619 a_71281_n10073.t15 a_71281_n10073.t14 VDD.t345 VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5620 VSS.t1022 VSS.t1021 VSS.t1022 VSS.t314 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5621 VDD.t1257 VDD.t1256 VDD.t1257 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5622 a_33249_48695.t88 a_33379_34917.t74 a_33249_35053.t71 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5623 VDD.t1255 VDD.t1253 VDD.t1255 VDD.t1254 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5624 a_83683_n34390# a_83153_n35156.t22 a_83153_n36322.t4 VDD.t2731 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5625 a_77225_n29181.t5 a_77225_n29181.t4 a_79151_n30339# VSS.t386 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5626 VDD.t1252 VDD.t1251 VDD.t1252 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5627 VSS.t1020 VSS.t1019 VSS.t1020 VSS.t382 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5628 VDD.t1250 VDD.t1249 VDD.t1250 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5629 a_99667_n8770# a_71281_n8397.t296 a_98829_n8770# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5630 a_89009_n27257.t2 a_83153_n36322.t21 a_90935_n30339# VSS.t460 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5631 VSS.t1018 VSS.t1017 VSS.t1018 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5632 a_38619_n8930# a_31953_n19727.t318 a_38097_n8930# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5633 VDD.t1248 VDD.t1247 VDD.t1248 VDD.t81 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5634 VDD.t1246 VDD.t1245 VDD.t1246 VDD.t403 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5635 VDD.t1244 VDD.t1243 VDD.t1244 VDD.t373 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5636 VDD.t1242 VDD.t1241 VDD.t1242 VDD.t908 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5637 VSS.t1016 VSS.t1015 VSS.t1016 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5638 VDD.t1240 VDD.t1239 VDD.t1240 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5639 VSS.t1014 VSS.t1013 VSS.t1014 VSS.t464 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5640 a_33249_48695.t144 a_33379_34007.t80 a_33249_34067.t30 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5641 VSS.t1012 VSS.t1011 VSS.t1012 VSS.t312 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5642 VSS.t1010 VSS.t1009 VSS.t1010 VSS.t673 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5643 VDD.t1238 VDD.t1237 VDD.t1238 VDD.t896 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5644 a_86903_n14095.t0 a_106830_10388.t20 a_108636_11614# VDD.t526 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5645 VDD.t1236 VDD.t1235 VDD.t1236 VDD.t623 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5646 OUT.t40 a_35922_19591.t154 a_52635_49681.t67 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5647 VDD.t4827 a_52635_34067.t221 a_52635_48695.t94 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5648 a_58851_n12421# a_50751_n19729.t316 a_57977_n16009.t0 VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5649 VSS.t1008 VSS.t1007 VSS.t1008 VSS.t542 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5650 a_33249_34067.t114 a_35502_25545.t89 VSS.t129 VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5651 VDD.t1234 VDD.t1233 VDD.t1234 VDD.t402 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5652 a_33249_48695.t182 a_31699_20742.t236 VDD.t261 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5653 VSS.t1006 VSS.t1005 VSS.t1006 VSS.t260 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5654 VSS.t1004 VSS.t1002 VSS.t1004 VSS.t1003 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5655 a_100803_n9675# a_71281_n8397.t297 a_100235_n9675# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5656 VSS.t1001 VSS.t1000 VSS.t1001 VSS.t207 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5657 a_60845_n17803# a_50751_n19729.t317 a_60285_n17803# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5658 VDD.t1232 VDD.t1231 VDD.t1232 VDD.t908 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5659 VSS.t999 VSS.t998 VSS.t999 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5660 VDD.t1230 VDD.t1229 VDD.t1230 VDD.t896 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5661 a_57417_n14215# a_50751_n19729.t318 a_56895_n15112# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5662 VDD.t1228 VDD.t1227 VDD.t1228 VDD.t524 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5663 a_47819_11614.t2 a_47819_10448.t19 a_49755_12380# VDD.t496 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5664 VDD.t1226 VDD.t1225 VDD.t1226 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5665 VDD.t1224 VDD.t1223 VDD.t1224 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5666 VDD.t1222 VDD.t1220 VDD.t1222 VDD.t1221 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5667 VDD.t1219 VDD.t1218 VDD.t1219 VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5668 VSS.t997 VSS.t996 VSS.t997 VSS.t211 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5669 VSS.t995 VSS.t994 VSS.t995 VSS.t593 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5670 a_32088_10448# a_30152_10448.t21 VDD.t305 VDD.t304 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5671 VSS.t993 VSS.t992 VSS.t993 VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5672 a_37934_4481# a_30152_11614.t20 a_30324_4421.t0 VSS.t324 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5673 a_93131_n17715# a_71281_n10073.t286 a_92601_n21335# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5674 a_33249_48695.t181 a_31699_20742.t237 VDD.t262 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5675 VDD.t1217 VDD.t1216 VDD.t1217 VDD.t123 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5676 VDD.t352 a_71281_n10073.t12 a_71281_n10073.t13 VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5677 VSS.t60 a_31953_n19727.t10 a_31953_n19727.t11 VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5678 a_71281_n10073.t11 a_71281_n10073.t10 VDD.t364 VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5679 VDD.t1215 VDD.t1214 VDD.t1215 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5680 a_57417_n3550# a_50751_n19729.t319 a_56895_n4447# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5681 VSS.t991 VSS.t990 VSS.t991 VSS.t352 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5682 VDD.t1213 VDD.t1211 VDD.t1213 VDD.t1212 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5683 VDD.t1210 VDD.t1208 VDD.t1210 VDD.t1209 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5684 VDD.t1207 VDD.t1206 VDD.t1207 VDD.t351 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5685 VSS.t989 VSS.t988 VSS.t989 VSS.t533 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5686 VDD.t1205 VDD.t1204 VDD.t1205 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5687 a_112199_n20430# a_71281_n8397.t298 a_111631_n20430# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5688 VSS.t987 VSS.t986 VSS.t987 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5689 a_93969_n18620# a_71281_n10073.t287 a_93131_n18620# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5690 VDD.t1203 VDD.t1202 VDD.t1203 VDD.t855 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5691 VDD.t4826 a_52635_34067.t222 a_52635_49681.t100 VDD.t400 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5692 VSS.t985 VSS.t983 VSS.t985 VSS.t984 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5693 a_66551_n2653# a_50751_n19729.t320 a_66029_n3550# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5694 a_41891_4481.t7 a_41891_4481.t6 a_43817_5639# VSS.t181 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5695 VDD.t1201 VDD.t1200 VDD.t1201 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5696 a_54579_n17803# a_50751_n19729.t321 a_54019_n17803# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5697 a_66058_n27257# a_65658_n29313.t2 a_65486_n35156.t11 VSS.t410 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5698 VSS.t982 VSS.t980 VSS.t982 VSS.t981 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5699 a_83709_n21335# a_71281_n10073.t288 a_83141_n21335# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5700 a_64243_n18700# a_50751_n19729.t322 a_63683_n17803# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5701 VDD.t1199 VDD.t1197 VDD.t1199 VDD.t1198 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5702 a_33787_n8033# a_31953_n19727.t319 a_33265_n8033# VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5703 VDD.t1196 VDD.t1195 VDD.t1196 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5704 a_89407_n19525# a_71281_n10073.t289 a_88839_n19525# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5705 a_46879_n3548# a_31953_n19727.t320 a_47753_n5342# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5706 a_50751_n19729.t21 a_50751_n19729.t20 VSS.t222 VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5707 VSS.t979 VSS.t978 VSS.t979 VSS.t623 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5708 VSS.t321 a_59558_n29181.t20 a_60080_n28415# VSS.t316 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5709 VDD.t1194 VDD.t1193 VDD.t1194 VDD.t855 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5710 VSS.t977 VSS.t976 VSS.t977 VSS.t54 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5711 VDD.t1192 VDD.t1190 VDD.t1192 VDD.t1191 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X5712 a_100803_n19525# a_71281_n8397.t299 a_100235_n19525# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5713 a_45445_n8033# a_31953_n19727.t321 a_44885_n8033# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5714 VDD.t1189 VDD.t1188 VDD.t1189 VDD.t28 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5715 VSS.t975 VSS.t974 VSS.t975 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5716 VDD.t1187 VDD.t1185 VDD.t1187 VDD.t1186 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5717 a_33249_48695.t145 a_33379_34007.t81 a_33249_34067.t29 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5718 a_31699_20742.t10 a_31699_20742.t9 VDD.t24 VDD.t23 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5719 a_64243_n8035# a_50751_n19729.t323 a_63683_n8035# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5720 a_75602_n4978# a_71266_n4019.t0 VDD.t4777 VDD.t695 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X5721 VDD.t263 a_31699_20742.t238 a_33249_48695.t180 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5722 VDD.t1184 VDD.t1182 VDD.t1184 VDD.t1183 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5723 a_52635_48695.t18 a_35922_19591.t155 a_52635_34067.t50 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5724 VSS.t59 a_31953_n19727.t8 a_31953_n19727.t9 VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5725 a_100820_10448.t2 a_100992_4421.t0 a_102796_5639# VSS.t173 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5726 a_31284_4481.t2 a_30324_5507.t1 a_30724_5639# VSS.t146 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5727 a_33249_48695.t179 a_31699_20742.t239 VDD.t264 VDD.t118 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5728 a_66016_n36322# a_65486_n35156.t22 a_65486_n36322.t3 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5729 VDD.t1181 VDD.t1179 VDD.t1181 VDD.t1180 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5730 a_40613_n7136# a_31953_n19727.t322 a_40053_n7136# VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5731 VSS.t973 VSS.t972 VSS.t973 VSS.t366 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5732 a_71281_n10073.t9 a_71281_n10073.t8 VDD.t342 VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5733 a_57977_n18700# a_50751_n19729.t324 a_57417_n17803# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5734 VDD.t1178 VDD.t1177 VDD.t1178 VDD.t557 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5735 VSS.t971 VSS.t970 VSS.t971 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5736 VDD.t1176 VDD.t1175 VDD.t1176 VDD.t836 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5737 a_65486_11614.t3 a_65486_10448.t19 a_67422_12380# VDD.t1381 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5738 VDD.t1174 VDD.t1173 VDD.t1174 VDD.t804 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5739 a_83141_n15000# a_71281_n10073.t290 a_82573_n15000# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5740 VSS.t969 VSS.t968 VSS.t969 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5741 VSS.t967 VSS.t966 VSS.t967 VSS.t2 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X5742 VSS.t965 VSS.t964 VSS.t965 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5743 VSS.t963 VSS.t962 VSS.t963 VSS.t861 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5744 VSS.t961 VSS.t960 VSS.t961 VSS.t469 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5745 a_54197_6405# a_47819_11614.t19 VDD.t510 VSS.t329 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5746 a_59558_4481.t0 a_47991_4421.t1 a_61515_13546# VDD.t493 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5747 a_93131_n21335# a_71281_n10073.t291 a_92601_n21335# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5748 VDD.t1172 VDD.t1171 VDD.t1172 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5749 VSS.t959 VSS.t958 VSS.t959 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5750 a_43817_5639# a_41891_4481.t19 VSS.t186 VSS.t160 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5751 a_88271_n21335# a_71281_n10073.t292 a_87433_n21335# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5752 VDD.t1170 VDD.t1169 VDD.t1170 VDD.t409 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5753 a_52635_48695.t17 a_35922_19591.t156 a_52635_34067.t45 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5754 VSS.t957 VSS.t956 VSS.t957 VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5755 VSS.t57 a_31953_n19727.t6 a_31953_n19727.t7 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5756 VDD.t1168 VDD.t1166 VDD.t1168 VDD.t1167 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5757 VDD.t1165 VDD.t1164 VDD.t1165 VDD.t836 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5758 VDD.t1163 VDD.t1162 VDD.t1163 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5759 VDD.t1161 VDD.t1160 VDD.t1161 VDD.t804 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5760 a_81735_n17715# a_71281_n10073.t293 a_81205_n16810# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5761 VSS.t955 VSS.t954 VSS.t955 VSS.t429 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5762 VDD.t1159 VDD.t1157 VDD.t1159 VDD.t1158 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5763 VDD.t1156 VDD.t1155 VDD.t1156 VDD.t979 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5764 VDD.t1154 VDD.t1153 VDD.t1154 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5765 a_59558_4481.t1 a_47991_4421.t1 a_61515_11614# VDD.t493 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5766 VSS.t953 VSS.t951 VSS.t953 VSS.t952 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5767 VSS.t950 VSS.t948 VSS.t950 VSS.t949 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5768 VDD.t1152 VDD.t1151 VDD.t1152 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5769 VSS.t947 VSS.t946 VSS.t947 VSS.t500 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5770 a_52635_48695.t16 a_35922_19591.t157 a_52635_34067.t29 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5771 VDD.t1150 VDD.t1149 VDD.t1150 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5772 VSS.t945 VSS.t944 VSS.t945 VSS.t686 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5773 a_81735_n15000# a_71281_n10073.t294 a_81205_n15905# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5774 a_93969_n6960# a_71281_n10073.t295 a_93131_n6960# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5775 a_33379_34917.t2 a_36162_10388.t21 a_37968_13546# VDD.t1497 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5776 a_112199_n2435# a_71281_n8397.t300 a_111631_n2435# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5777 a_42047_n15110# a_31953_n19727.t323 a_41487_n15110# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5778 VSS.t943 VSS.t941 VSS.t943 VSS.t942 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5779 VSS.t940 VSS.t939 VSS.t940 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5780 a_41487_n6239# a_31953_n19727.t324 a_40965_n6239# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5781 OUT.t39 a_35922_19591.t158 a_52635_49681.t68 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5782 a_52635_34067.t43 a_35922_19591.t159 a_52635_48695.t15 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5783 a_101392_5639# a_57977_n12421.t0 a_100820_11614.t4 VSS.t175 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5784 VDD.t1148 VDD.t1147 VDD.t1148 VDD.t65 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5785 a_94537_n1530# a_71281_n10073.t296 a_93969_n1530# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5786 a_33249_48695.t146 a_33379_34007.t82 a_33249_34067.t28 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5787 VSS.t938 VSS.t937 VSS.t938 VSS.t398 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5788 a_112199_n15905# a_71281_n8397.t301 a_111631_n15905# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5789 VSS.t221 a_50751_n19729.t18 a_50751_n19729.t19 VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5790 VSS.t936 VSS.t935 VSS.t936 VSS.t483 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5791 a_30724_5639# a_30324_5507.t1 a_30152_11614.t2 VSS.t145 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5792 a_82573_n7865# a_71281_n10073.t297 a_81735_n7865# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5793 VSS.t934 VSS.t933 VSS.t934 VSS.t676 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5794 VSS.t932 VSS.t931 VSS.t932 VSS.t692 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5795 VDD.t1146 VDD.t1144 VDD.t1146 VDD.t1145 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5796 a_71342_4481.t2 a_71496_10388.t23 a_71896_10448# VDD.t489 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5797 VSS.t930 VSS.t929 VSS.t930 VSS.t500 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5798 VDD.t1143 VDD.t1142 VDD.t1143 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5799 VDD.t1141 VDD.t1140 VDD.t1141 VDD.t792 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5800 VDD.t1139 VDD.t1138 VDD.t1139 VDD.t500 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5801 a_33249_48695.t89 a_33379_34917.t75 a_33249_35053.t72 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5802 VSS.t928 VSS.t927 VSS.t928 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5803 VSS.t926 VSS.t925 VSS.t926 VSS.t191 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5804 a_36032_11614.t0 a_36162_10388.t22 a_37968_11614# VDD.t1497 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5805 VDD.t1137 VDD.t1136 VDD.t1137 VDD.t50 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5806 VSS.t924 VSS.t923 VSS.t924 VSS.t573 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5807 VSS.t922 VSS.t921 VSS.t922 VSS.t287 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5808 VDD.t1135 VDD.t1134 VDD.t1135 VDD.t65 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5809 a_30324_n30399.t0 a_31953_n19727.t325 a_32353_n19595# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5810 a_99667_n7865# a_71281_n8397.t302 a_98829_n7865# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5811 a_42047_n2651# a_31953_n19727.t326 a_41487_n2651# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5812 a_33249_34067.t113 a_35502_25545.t90 VSS.t128 VSS.t49 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5813 VSS.t408 a_59558_4481.t21 a_60080_4481# VSS.t316 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5814 a_83141_n20430# a_71281_n10073.t298 a_82573_n20430# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5815 VSS.t920 VSS.t919 VSS.t920 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5816 a_33249_48695.t90 a_33379_34917.t76 a_33249_35053.t73 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5817 a_61484_n27257# a_59558_n29181.t21 VSS.t322 VSS.t314 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5818 a_32913_n6239# a_31953_n19727.t327 a_32353_n4445# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5819 a_83153_11614.t0 a_51711_n12421.t0 a_85129_4481# VSS.t297 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5820 a_33249_48695.t91 a_33379_34917.t77 a_33249_35053.t74 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5821 VSS.t918 VSS.t917 VSS.t918 VSS.t335 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5822 VSS.t916 VSS.t915 VSS.t916 VSS.t550 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5823 VSS.t914 VSS.t912 VSS.t914 VSS.t913 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5824 a_100820_n36322.t5 a_39179_n8930.t1 a_102796_n27257# VSS.t382 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5825 VSS.t911 VSS.t909 VSS.t911 VSS.t910 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5826 VDD.t1133 VDD.t1132 VDD.t1133 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5827 VSS.t310 I1N.t15 a_72603_n9297# VSS.t305 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X5828 a_83709_n3340# a_71281_n10073.t299 a_83141_n3340# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5829 VDD.t4825 a_52635_34067.t223 a_52635_49681.t99 VDD.t403 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5830 VDD.t4824 a_52635_34067.t224 a_52635_49681.t98 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5831 a_73302_n36322# a_71496_n36382.t17 a_71342_n27257.t3 VDD.t2814 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5832 VDD.t1131 VDD.t1129 VDD.t1131 VDD.t1130 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5833 VDD.t1128 VDD.t1127 VDD.t1128 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5834 a_71864_n29181# a_65486_n36322.t23 VDD.t299 VSS.t153 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5835 VDD.t1126 VDD.t1125 VDD.t1126 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5836 a_52635_34067.t3 a_35502_24538.t61 a_33249_34067.t1 VSS.t183 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5837 VDD.t1124 VDD.t1123 VDD.t1124 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5838 a_81735_n20430# a_71281_n10073.t300 VDD.t386 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5839 VDD.t1122 VDD.t1121 VDD.t1122 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5840 a_88839_n9675# a_71281_n10073.t301 a_88271_n9675# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5841 a_31284_n30339.t0 a_30324_n29313.t0 a_30724_n29181# VSS.t146 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5842 a_87433_n18620# a_71281_n10073.t302 a_86903_n19525# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5843 VDD.t1120 VDD.t1119 VDD.t1120 VDD.t928 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5844 VSS.t908 VSS.t907 VSS.t908 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5845 a_100820_n36322.t2 a_100820_n35156.t19 a_102756_n35156# VDD.t528 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5846 VDD.t1118 VDD.t1117 VDD.t1118 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5847 VDD.t1116 VDD.t1114 VDD.t1116 VDD.t1115 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5848 a_89407_n4245# a_71281_n10073.t303 a_88839_n4245# VDD.t332 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5849 a_39179_n16904# a_31953_n19727.t328 a_38619_n15110# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5850 a_71496_10388.t7 a_71366_11614.t10 a_79182_10448# VDD.t1843 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5851 VDD.t1113 VDD.t1112 VDD.t1113 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5852 VSS.t906 VSS.t905 VSS.t906 VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5853 a_55601_n30339# a_47819_n36322.t22 a_47991_n29313.t0 VSS.t330 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5854 VSS.t904 VSS.t903 VSS.t904 VSS.t95 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5855 a_33249_48695.t92 a_33379_34917.t78 a_33249_35053.t75 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5856 VDD.t1111 VDD.t1110 VDD.t1111 VDD.t394 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5857 a_33787_n3548# a_31953_n19727.t329 a_33265_n3548# VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5858 VSS.t902 VSS.t900 VSS.t902 VSS.t901 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5859 VSS.t899 VSS.t898 VSS.t899 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5860 a_71281_n10073.t7 a_71281_n10073.t6 VDD.t359 VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5861 a_33787_n12419# a_31953_n19727.t330 VSS.t118 VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5862 a_33249_48695.t178 a_31699_20742.t240 VDD.t265 VDD.t123 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5863 VSS.t897 VSS.t895 VSS.t897 VSS.t896 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5864 a_45445_n3548# a_31953_n19727.t331 a_44885_n3548# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5865 a_107198_n27257# a_100820_n36322.t20 a_106676_n27257.t0 VSS.t352 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5866 a_51711_n12421.t0 a_83153_11614.t21 a_89531_5639# VSS.t399 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5867 VDD.t1109 VDD.t1108 VDD.t1109 VDD.t17 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5868 a_48349_n34390# a_47819_n35156.t19 a_47819_n36322.t1 VDD.t2561 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5869 a_100820_n36322.t3 a_100820_n35156.t20 a_102756_n33224# VDD.t528 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5870 a_105933_n13190# a_71281_n8397.t303 a_105365_n13190# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5871 a_46879_n17801# a_31953_n19727.t332 a_46319_n17801# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5872 VSS.t894 VSS.t893 VSS.t894 VSS.t20 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X5873 a_33249_48695.t177 a_31699_20742.t241 VDD.t266 VDD.t125 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5874 VDD.t1107 VDD.t1106 VDD.t1107 VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5875 VSS.t892 VSS.t891 VSS.t892 VSS.t40 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5876 VDD.t1105 VDD.t1104 VDD.t1105 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5877 VDD.t538 a_100820_n35156.t21 a_101350_n35156# VDD.t535 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5878 a_64243_n3550# a_50751_n19729.t325 a_63683_n3550# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5879 VDD.t1103 VDD.t1101 VDD.t1103 VDD.t1102 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5880 VDD.t1100 VDD.t1099 VDD.t1100 VDD.t913 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5881 a_51711_n18700# a_50751_n19729.t326 a_51151_n18700# VSS.t249 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5882 VDD.t1098 VDD.t1097 VDD.t1098 VDD.t901 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5883 VSS.t127 a_35502_25545.t91 a_35922_19591.t2 VSS.t126 nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X5884 a_87433_n1530# a_71281_n10073.t304 a_86903_n5150# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5885 a_31699_20742.t8 a_31699_20742.t7 VDD.t22 VDD.t21 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5886 VDD.t1096 VDD.t1095 VDD.t1096 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5887 a_35781_n4445# a_31953_n19727.t333 a_35221_n4445# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5888 VSS.t890 VSS.t888 VSS.t890 VSS.t889 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5889 VDD.t1094 VDD.t1093 VDD.t1094 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5890 VDD.t1092 VDD.t1091 VDD.t1092 VDD.t321 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5891 VDD.t1090 VDD.t1088 VDD.t1090 VDD.t1089 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5892 a_53145_n14215# a_50751_n19729.t327 a_52585_n14215# VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5893 VSS.t887 VSS.t886 VSS.t887 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5894 VSS.t885 VSS.t884 VSS.t885 VSS.t278 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5895 a_65486_n35156.t10 a_65658_n29313.t0 a_67462_n28415# VSS.t413 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5896 a_71281_n8397.t5 a_71281_n8397.t4 VDD.t425 VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5897 VSS.t883 VSS.t881 VSS.t883 VSS.t882 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5898 VSS.t880 VSS.t879 VSS.t880 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5899 VDD.t1087 VDD.t1086 VDD.t1087 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5900 VDD.t539 a_100820_n35156.t22 a_101350_n33224# VDD.t535 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5901 a_104527_n13190# a_71281_n8397.t304 a_103997_n16810# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5902 VSS.t878 VSS.t877 VSS.t878 VSS.t15 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5903 a_95105_n3340# a_71281_n10073.t305 a_94537_n3340# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5904 VDD.t1085 VDD.t1083 VDD.t1085 VDD.t1084 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5905 a_31699_17542# I1U.t6 VSS.t364 VSS.t362 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X5906 VSS.t876 VSS.t875 VSS.t876 VSS.t188 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5907 a_83141_n15905# a_71281_n10073.t306 a_82573_n15905# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5908 VDD.t267 a_31699_20742.t242 a_33249_48695.t176 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5909 VDD.t1082 VDD.t1081 VDD.t1082 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5910 a_52635_49681.t69 a_35922_19591.t160 OUT.t38 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5911 a_52635_34067.t51 a_35922_19591.t161 a_52635_48695.t14 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5912 a_83141_n9675# a_71281_n10073.t307 a_82573_n9675# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5913 VSS.t874 VSS.t872 VSS.t874 VSS.t873 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5914 VSS.t871 VSS.t870 VSS.t871 VSS.t762 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5915 VDD.t1080 VDD.t1079 VDD.t1080 VDD.t923 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X5916 VDD.t1078 VDD.t1077 VDD.t1078 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5917 a_33249_48695.t93 a_33379_34917.t79 a_33249_35053.t76 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5918 VDD.t1076 VDD.t1075 VDD.t1076 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5919 VDD.t1074 VDD.t1073 VDD.t1074 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5920 a_36562_n35156# a_36162_n36382.t22 a_36032_n35156.t4 VDD.t683 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5921 VSS.t869 VSS.t868 VSS.t869 VSS.t563 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5922 VSS.t357 a_89163_n36382.t22 a_89563_n34390# VDD.t548 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5923 a_41487_n16007# a_31953_n19727.t334 a_40613_n17801# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5924 VDD.t268 a_31699_20742.t243 a_33249_48695.t175 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5925 VSS.t867 VSS.t866 VSS.t867 VSS.t459 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5926 VDD.t1072 VDD.t1071 VDD.t1072 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5927 VSS.t865 VSS.t863 VSS.t865 VSS.t864 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5928 VSS.t125 a_35502_25545.t92 a_33249_34067.t112 VSS.t35 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5929 a_100235_n9675# a_71281_n8397.t305 a_99667_n9675# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5930 VDD.t1070 VDD.t1069 VDD.t1070 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5931 VDD.t517 a_47819_10448.t20 a_48349_13546# VDD.t512 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5932 a_33249_48695.t147 a_33379_34007.t83 a_33249_34067.t27 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5933 VSS.t862 VSS.t860 VSS.t862 VSS.t861 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5934 a_89531_5639# a_83153_11614.t22 VDD.t4771 VSS.t400 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5935 VDD.t1068 VDD.t1067 VDD.t1068 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5936 a_93969_n21335# a_71281_n10073.t308 a_93131_n21335# VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5937 a_47753_n8033# a_31953_n19727.t335 a_47231_n8033# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5938 a_57417_n2653# a_50751_n19729.t328 a_56895_n2653# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5939 VSS.t859 VSS.t857 VSS.t859 VSS.t858 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5940 VDD.t1066 VDD.t1065 VDD.t1066 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5941 a_81735_n15905# a_71281_n10073.t309 a_81205_n15905# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5942 VSS.t856 VSS.t855 VSS.t856 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5943 a_81735_n6055# a_71281_n10073.t310 a_81205_n9675# VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5944 VSS.t854 VSS.t853 VSS.t854 VSS.t100 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5945 a_99667_n19525# a_71281_n8397.t306 a_98829_n19525# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5946 VDD.t1064 VDD.t1063 VDD.t1064 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5947 VDD.t1062 VDD.t1061 VDD.t1062 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5948 VDD.t1060 VDD.t1059 VDD.t1060 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5949 VSS.t852 VSS.t851 VSS.t852 VSS.t283 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5950 a_36562_n33224# a_36162_n36382.t23 a_33379_34007.t3 VDD.t683 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5951 a_60845_n8932# a_50751_n19729.t329 a_60285_n8932# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5952 a_33249_48695.t94 a_33379_34917.t80 a_33249_35053.t77 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5953 a_83683_n36322# a_83153_n35156.t23 a_83153_n36322.t5 VDD.t2731 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5954 VDD.t1058 VDD.t1057 VDD.t1058 VDD.t845 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5955 VDD.t269 a_31699_20742.t244 a_35502_25545.t19 VDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5956 a_52635_34067.t45 a_35922_19591.t162 a_52635_48695.t13 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5957 VSS.t850 VSS.t849 VSS.t850 VSS.t495 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5958 VSS.t848 VSS.t846 VSS.t848 VSS.t847 nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X5959 VDD.t1056 VDD.t1054 VDD.t1056 VDD.t1055 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5960 VDD.t1053 VDD.t1051 VDD.t1053 VDD.t1052 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5961 a_50751_n19729.t17 a_50751_n19729.t16 VSS.t220 VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5962 a_111063_n19525# a_71281_n8397.t307 a_110225_n19525# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5963 a_98829_n6055# a_71281_n8397.t308 a_98299_n9675# VDD.t468 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5964 VSS.t845 VSS.t844 VSS.t845 VSS.t63 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5965 VDD.t1050 VDD.t1049 VDD.t1050 VDD.t831 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5966 a_52635_49681.t70 a_35922_19591.t163 OUT.t37 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5967 VDD.t518 a_47819_10448.t21 a_48349_11614# VDD.t512 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5968 VDD.t1048 VDD.t1047 VDD.t1048 VDD.t63 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5969 VSS.t124 a_35502_25545.t93 a_33249_34067.t111 VSS.t44 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5970 VDD.t1046 VDD.t1044 VDD.t1046 VDD.t1045 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5971 VDD.t1043 VDD.t1042 VDD.t1043 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5972 VSS.t843 VSS.t841 VSS.t843 VSS.t842 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5973 VDD.t1041 VDD.t1040 VDD.t1041 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5974 a_112507_n6055.t0 a_71281_n8397.t309 a_112199_n9675# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5975 a_89715_n17715.t2 a_100992_4421.t1 a_113110_10448# VDD.t374 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5976 VDD.t1039 VDD.t1038 VDD.t1039 VDD.t623 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5977 a_52635_48695.t12 a_35922_19591.t164 a_52635_34067.t52 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5978 a_44885_n16007# a_31953_n19727.t336 a_44363_n16007.t0 VSS.t99 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5979 a_95943_n18620# a_71281_n10073.t311 a_95105_n18620# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5980 a_33249_48695.t148 a_33379_34007.t84 a_33249_34067.t26 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5981 VDD.t1037 VDD.t1036 VDD.t1037 VDD.t52 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5982 VDD.t1035 VDD.t1034 VDD.t1035 VDD.t6 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5983 VSS.t840 VSS.t838 VSS.t840 VSS.t839 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5984 a_84547_n6055# a_71281_n10073.t312 a_84017_n5150.t1 VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5985 a_52635_49681.t97 a_52635_34067.t225 VDD.t4823 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5986 VSS.t837 VSS.t836 VSS.t837 VSS.t576 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5987 a_95443_13546# a_81205_n14095.t9 a_89163_10388.t6 VDD.t500 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5988 a_33249_48695.t174 a_31699_20742.t245 VDD.t270 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5989 a_35221_n16904# a_31953_n19727.t337 a_34699_n16904# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5990 VSS.t835 VSS.t834 VSS.t835 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5991 VDD.t1033 VDD.t1032 VDD.t1033 VDD.t938 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5992 VDD.t271 a_31699_20742.t246 a_33249_48695.t173 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5993 VSS.t833 VSS.t832 VSS.t833 VSS.t676 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5994 VDD.t1031 VDD.t1030 VDD.t1031 VDD.t642 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5995 VDD.t1029 VDD.t1028 VDD.t1029 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5996 VDD.t1027 VDD.t1026 VDD.t1027 VDD.t965 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5997 VDD.t1025 VDD.t1024 VDD.t1025 VDD.t52 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5998 a_111063_n6960# a_71281_n8397.t310 a_110225_n6960# VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5999 a_33249_48695.t95 a_33379_34917.t81 a_33249_35053.t78 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6000 VSS.t831 VSS.t830 VSS.t831 VSS.t563 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6001 a_54229_n34390# a_53829_n36382.t21 a_53699_n35156.t2 VDD.t322 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6002 VSS.t829 VSS.t828 VSS.t829 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6003 a_83709_n2435# a_71281_n10073.t313 a_83141_n2435# VDD.t311 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6004 a_94537_n18620# a_71281_n10073.t314 a_93969_n18620# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6005 a_95443_11614# a_81205_n14095.t10 a_89163_10388.t7 VDD.t500 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6006 a_111631_n1530# a_71281_n8397.t311 a_111063_n1530# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6007 VSS.t827 VSS.t826 VSS.t827 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6008 VDD.t1023 VDD.t1022 VDD.t1023 VDD.t795 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6009 VDD.t4753 a_65486_10448.t20 a_66016_13546# VDD.t1341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6010 VDD.t1021 VDD.t1020 VDD.t1021 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6011 OUT.t36 a_35922_19591.t165 a_52635_49681.t71 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6012 a_48951_4481.t2 a_47991_4421.t2 a_48391_4481# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6013 VSS.t825 VSS.t824 VSS.t825 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6014 a_89009_4481.t3 a_89163_10388.t21 a_89563_10448# VDD.t558 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6015 VSS.t823 VSS.t821 VSS.t823 VSS.t822 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X6016 VDD.t1019 VDD.t1017 VDD.t1019 VDD.t1018 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6017 VDD.t1016 VDD.t1015 VDD.t1016 VDD.t602 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6018 VSS.t820 VSS.t818 VSS.t820 VSS.t819 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6019 VSS.t817 VSS.t815 VSS.t817 VSS.t816 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6020 a_60080_4481# a_59558_4481.t9 a_59558_4481.t10 VSS.t313 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6021 a_33249_48695.t172 a_31699_20742.t247 VDD.t272 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6022 a_40613_n19595# a_31953_n19727.t338 a_40053_n18698# VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6023 VSS.t56 a_31953_n19727.t4 a_31953_n19727.t5 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6024 a_87433_n17715# a_71281_n10073.t315 a_86903_n21335# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6025 VSS.t814 VSS.t812 VSS.t814 VSS.t813 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6026 VDD.t4822 a_52635_34067.t226 a_52635_49681.t96 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6027 a_93131_n6055# a_71281_n10073.t316 a_92601_n9675# VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6028 VSS.t811 VSS.t810 VSS.t811 VSS.t97 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6029 VDD.t485 a_71281_n8397.t312 a_112199_n13190# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6030 VDD.t4821 a_52635_34067.t227 a_52635_49681.t95 VDD.t415 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6031 VSS.t809 VSS.t808 VSS.t809 VSS.t530 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6032 VDD.t4754 a_65486_10448.t21 a_66016_11614# VDD.t1341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6033 VDD.t1014 VDD.t1013 VDD.t1014 VDD.t41 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6034 a_40053_n19595# a_31953_n19727.t339 a_39179_n16007.t1 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6035 VSS.t807 VSS.t806 VSS.t807 VSS.t149 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6036 VDD.t1012 VDD.t1011 VDD.t1012 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6037 a_101350_13546# a_100820_10448.t21 a_100820_11614.t1 VDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6038 a_42047_n15110# a_31953_n19727.t340 a_41487_n14213# VSS.t98 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6039 a_41487_n5342# a_31953_n19727.t341 a_40613_n7136# VSS.t104 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6040 a_35221_n4445# a_31953_n19727.t342 a_34699_n6239# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6041 VSS.t805 VSS.t804 VSS.t805 VSS.t527 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6042 a_33249_48695.t96 a_33379_34917.t82 a_33249_35053.t79 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6043 a_100803_n3340# a_71281_n8397.t313 a_100235_n3340# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6044 VDD.t1010 VDD.t1009 VDD.t1010 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6045 VDD.t1008 VDD.t1007 VDD.t1008 VDD.t85 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6046 VDD.t1006 VDD.t1005 VDD.t1006 VDD.t396 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6047 VSS.t803 VSS.t802 VSS.t803 VSS.t416 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6048 VSS.t219 a_50751_n19729.t14 a_50751_n19729.t15 VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6049 VSS.t801 VSS.t799 VSS.t801 VSS.t800 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6050 a_42442_n35156# a_30324_n29313.t2 a_41891_n29181.t0 VDD.t564 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6051 a_57977_n8035# a_50751_n19729.t330 a_57417_n8035# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6052 VSS.t798 VSS.t796 VSS.t798 VSS.t797 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6053 a_96011_n36322.t1 a_89033_n35156.t11 a_95443_n34390# VDD.t2425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6054 VSS.t795 VSS.t794 VSS.t795 VSS.t189 nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X6055 a_52635_48695.t11 a_35922_19591.t166 a_52635_34067.t53 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6056 VSS.t793 VSS.t792 VSS.t793 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6057 VDD.t1004 VDD.t1003 VDD.t1004 VDD.t293 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6058 a_95943_n6055# a_71281_n10073.t317 a_95413_n5150.t1 VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6059 VSS.t791 VSS.t790 VSS.t791 VSS.t24 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6060 VDD.t1002 VDD.t1001 VDD.t1002 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6061 VDD.t4820 a_52635_34067.t228 a_52635_49681.t94 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6062 a_51151_n7138# a_50751_n19729.t331 a_50629_n7138# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6063 VSS.t311 I1N.t16 a_72603_n10973# VSS.t305 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X6064 a_101350_11614# a_100820_10448.t22 a_100820_11614.t2 VDD.t323 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6065 VDD.t1000 VDD.t999 VDD.t1000 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6066 a_105933_n9675# a_71281_n8397.t314 a_105365_n9675# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6067 VSS.t789 VSS.t788 VSS.t789 VSS.t596 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6068 a_53145_n7138# a_50751_n19729.t332 a_52585_n7138# VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6069 VDD.t998 VDD.t996 VDD.t998 VDD.t997 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X6070 VDD.t995 VDD.t994 VDD.t995 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6071 VDD.t993 VDD.t992 VDD.t993 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6072 VDD.t991 VDD.t990 VDD.t991 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6073 a_42442_n33224# a_30324_n29313.t2 a_41891_n29181.t0 VDD.t564 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6074 a_33249_48695.t171 a_31699_20742.t248 VDD.t273 VDD.t81 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6075 VDD.t543 a_100820_n36322.t21 a_108602_n28415# VSS.t350 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6076 VSS.t787 VSS.t786 VSS.t787 VSS.t514 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6077 a_106501_n4245# a_71281_n8397.t315 a_105933_n4245# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6078 VSS.t132 a_35502_25545.t94 a_33249_34067.t110 VSS.t49 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X6079 a_33249_35053.t110 a_35502_25545.t95 VSS.t140 VSS.t134 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6080 VSS.t785 VSS.t784 VSS.t785 VSS.t673 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6081 a_52635_49681.t93 a_52635_34067.t229 VDD.t4819 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6082 VDD.t989 VDD.t988 VDD.t989 VDD.t65 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6083 VSS.t783 VSS.t782 VSS.t783 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6084 VSS.t781 VSS.t779 VSS.t781 VSS.t780 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6085 VDD.t987 VDD.t986 VDD.t987 VDD.t751 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6086 VSS.t778 VSS.t776 VSS.t778 VSS.t777 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6087 a_95105_n2435# a_71281_n10073.t318 a_94537_n2435# VDD.t315 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6088 VSS.t345 a_77225_4481.t21 a_77747_4481# VSS.t341 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6089 OUT.t109 a_33379_34917.t0 cap_mim_2f0_m4m5_noshield c_width=9.8u c_length=9.8u
X6090 VDD.t985 VDD.t984 VDD.t985 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6091 VDD.t983 VDD.t981 VDD.t983 VDD.t982 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6092 VDD.t4818 a_52635_34067.t230 a_52635_48695.t93 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6093 a_85129_n27257# a_32913_n8930.t1 a_31831_n5342.t1 VSS.t278 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6094 VDD.t980 VDD.t978 VDD.t980 VDD.t979 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6095 VDD.t977 VDD.t976 VDD.t977 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6096 a_63161_n5344.t1 a_65658_4421.t0 a_66058_6405# VSS.t411 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6097 a_104527_n6055# a_71281_n8397.t316 a_103997_n9675# VDD.t470 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6098 VDD.t975 VDD.t974 VDD.t975 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6099 a_112199_n14095# a_71281_n8397.t317 a_111631_n14095# VDD.t426 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6100 VSS.t775 VSS.t774 VSS.t775 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6101 VDD.t973 VDD.t972 VDD.t973 VDD.t58 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6102 VDD.t507 a_30152_11614.t21 a_37934_6405# VSS.t323 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6103 VDD.t971 VDD.t970 VDD.t971 VDD.t728 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6104 a_47753_n3548# a_31953_n19727.t343 a_47231_n3548# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6105 VDD.t969 VDD.t967 VDD.t969 VDD.t968 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6106 a_87433_n21335# a_71281_n10073.t319 a_86903_n21335# VDD.t308 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6107 VSS.t773 VSS.t772 VSS.t773 VSS.t181 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6108 VDD.t966 VDD.t964 VDD.t966 VDD.t965 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X6109 VSS.t771 VSS.t770 VSS.t771 VSS.t101 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6110 VDD.t963 VDD.t962 VDD.t963 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6111 a_77747_6405# a_77225_4481.t4 a_77225_4481.t5 VSS.t336 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6112 VDD.t20 a_31699_20742.t5 a_31699_20742.t6 VDD.t19 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6113 VSS.t769 VSS.t767 VSS.t769 VSS.t768 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X6114 VDD.t961 VDD.t960 VDD.t961 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6115 a_33249_48695.t149 a_33379_34007.t85 a_33249_34067.t25 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6116 VSS.t766 VSS.t764 VSS.t766 VSS.t765 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6117 a_33249_48695.t97 a_33379_34917.t83 a_33249_35053.t80 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6118 VSS.t763 VSS.t761 VSS.t763 VSS.t762 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6119 VSS.t217 a_50751_n19729.t12 a_50751_n19729.t13 VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6120 OUT.t35 a_35922_19591.t167 a_52635_49681.t72 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6121 VSS.t760 VSS.t759 VSS.t760 VSS.t312 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6122 a_44363_n16007.t2 a_45445_n19595.t1 a_66058_n30339# VSS.t411 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6123 VDD.t959 VDD.t957 VDD.t959 VDD.t958 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6124 a_58851_n18700# a_50751_n19729.t333 a_58329_n18700# VSS.t223 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6125 a_39179_n14213# a_31953_n19727.t344 a_38619_n14213# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6126 a_52635_48695.t10 a_35922_19591.t168 a_52635_34067.t54 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6127 a_33249_48695.t170 a_31699_20742.t249 VDD.t274 VDD.t52 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6128 a_60845_n13318# a_50751_n19729.t334 a_60285_n13318# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6129 VDD.t275 a_31699_20742.t250 a_33249_48695.t169 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6130 a_89531_n27257# a_83153_n36322.t22 a_89009_n27257.t3 VSS.t459 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6131 a_102796_n29181# a_39179_n8930.t2 a_38097_n5342.t0 VSS.t383 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6132 VSS.t758 VSS.t757 VSS.t758 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6133 a_33787_n2651# a_31953_n19727.t345 a_33265_n3548# VSS.t66 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6134 a_50751_n19729.t11 a_50751_n19729.t10 VSS.t216 VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6135 VDD.t956 VDD.t955 VDD.t956 VDD.t933 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6136 VDD.t954 VDD.t953 VDD.t954 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6137 VDD.t302 a_100820_10448.t23 a_101350_10448# VDD.t301 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6138 a_61484_7563# a_59558_4481.t22 VSS.t409 VSS.t314 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6139 a_60109_12380# a_47991_4421.t1 a_59558_4481.t2 VDD.t492 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6140 VDD.t952 VDD.t951 VDD.t952 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6141 a_35781_n17801# a_31953_n19727.t346 a_35221_n17801# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6142 a_52635_49681.t73 a_35922_19591.t169 OUT.t34 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6143 a_60285_n14215# a_50751_n19729.t335 a_59763_n14215# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6144 VDD.t4817 a_52635_34067.t231 a_52635_49681.t92 VDD.t409 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6145 OUT.t3 a_35502_24538.t62 a_33249_35053.t105 VSS.t183 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6146 a_113081_n30339# a_112559_n29181.t21 a_106830_n36382.t1 VSS.t415 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6147 VDD.t950 VDD.t949 VDD.t950 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6148 VSS.t756 VSS.t755 VSS.t756 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6149 VSS.t754 VSS.t752 VSS.t754 VSS.t753 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6150 a_106676_7563.t1 a_100820_11614.t22 a_108602_4481# VSS.t151 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6151 a_45445_n3548# a_31953_n19727.t347 a_44885_n2651# VSS.t95 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6152 a_30324_4421.t0 a_30152_11614.t22 a_36530_4481# VSS.t325 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6153 VDD.t948 VDD.t946 VDD.t948 VDD.t947 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6154 a_38097_n16007.t2 a_47991_n29313.t2 a_48391_n27257# VSS.t283 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6155 a_32128_6405# a_30324_5507.t2 a_31284_4481.t2 VSS.t148 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6156 VDD.t945 VDD.t944 VDD.t945 VDD.t406 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X6157 VDD.t943 VDD.t942 VDD.t943 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6158 a_64243_n3550# a_50751_n19729.t336 a_63683_n2653# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6159 VDD.t941 VDD.t940 VDD.t941 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6160 VDD.t939 VDD.t937 VDD.t939 VDD.t938 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6161 VDD.t936 VDD.t935 VDD.t936 VDD.t491 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6162 OUT.t33 a_35922_19591.t170 a_52635_49681.t74 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6163 VSS.t139 a_35502_25545.t96 a_33249_35053.t109 VSS.t18 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6164 a_95943_n17715# a_71281_n10073.t320 VDD.t387 VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6165 VSS.t751 VSS.t749 VSS.t751 VSS.t750 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6166 VDD.t934 VDD.t932 VDD.t934 VDD.t933 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6167 a_114516_13546# a_100992_4421.t1 a_89715_n17715.t4 VDD.t373 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6168 VSS.t748 VSS.t747 VSS.t748 VSS.t623 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6169 VSS.t746 VSS.t744 VSS.t746 VSS.t745 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6170 a_110225_n8770# a_71281_n8397.t318 VDD.t486 VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6171 a_84547_n6960# a_71281_n10073.t321 a_83709_n4245# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6172 VSS.t743 VSS.t742 VSS.t743 VSS.t316 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6173 a_54579_n13318# a_50751_n19729.t337 a_54019_n13318# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6174 a_40613_n2651# a_31953_n19727.t348 a_40053_n1754# VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6175 VDD.t931 VDD.t930 VDD.t931 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6176 a_33249_48695.t150 a_33379_34007.t86 a_33249_34067.t24 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6177 a_33249_34067.t23 a_33379_34007.t87 a_33249_48695.t151 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6178 a_47819_n35156.t5 a_47819_n35156.t4 a_49755_n34390# VDD.t2328 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6179 a_39179_n8930.t0 a_31953_n19727.t349 a_38619_n8930# VSS.t96 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6180 a_52635_34067.t55 a_35922_19591.t171 a_52635_48695.t9 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6181 VDD.t929 VDD.t927 VDD.t929 VDD.t928 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6182 a_64243_n14215# a_50751_n19729.t338 a_63683_n13318# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6183 VDD.t926 VDD.t925 VDD.t926 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6184 a_110225_n19525# a_71281_n8397.t319 a_109695_n19525# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6185 a_33249_48695.t98 a_33379_34917.t84 a_33249_35053.t81 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6186 a_52635_34067.t46 a_35922_19591.t172 a_52635_48695.t8 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6187 VDD.t4816 a_52635_34067.t232 a_52635_49681.t91 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6188 a_33249_48695.t168 a_31699_20742.t251 VDD.t276 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6189 VSS.t741 VSS.t740 VSS.t741 VSS.t52 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6190 a_114516_11614# a_100992_4421.t1 a_89715_n17715.t3 VDD.t373 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6191 VSS.t379 a_41891_n29181.t22 a_42413_n28415# VSS.t171 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6192 VDD.t924 VDD.t922 VDD.t924 VDD.t923 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X6193 VDD.t921 VDD.t919 VDD.t921 VDD.t920 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6194 VDD.t918 VDD.t917 VDD.t918 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6195 VSS.t396 a_77225_n29181.t22 a_77747_n30339# VSS.t390 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6196 VDD.t4984 a_71281_n10073.t4 a_71281_n10073.t5 VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6197 VSS.t739 VSS.t737 VSS.t739 VSS.t738 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6198 a_106676_7563.t3 a_106830_10388.t21 a_107230_13546# VDD.t524 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6199 a_33249_48695.t99 a_33379_34917.t85 a_33249_35053.t82 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6200 a_82573_n1530# a_71281_n10073.t322 a_81735_n1530# VDD.t321 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6201 OUT.t1 a_106830_10388.t22 a_108636_10448# VDD.t526 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6202 VDD.t4806 a_47819_n35156.t20 a_48349_n34390# VDD.t2291 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6203 VSS.t736 VSS.t734 VSS.t736 VSS.t735 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6204 VDD.t916 VDD.t915 VDD.t916 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6205 a_46319_n12419# a_31953_n19727.t350 VSS.t119 VSS.t58 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6206 VDD.t914 VDD.t912 VDD.t914 VDD.t913 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6207 a_106501_n13190# a_71281_n8397.t320 a_105933_n13190# VDD.t424 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6208 a_52635_49681.t75 a_35922_19591.t173 OUT.t32 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6209 VSS.t733 VSS.t732 VSS.t733 VSS.t104 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6210 a_99667_n1530# a_71281_n8397.t321 a_98829_n1530# VDD.t433 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6211 a_108602_4481# a_100820_11614.t23 a_100992_4421.t0 VSS.t147 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6212 a_57977_n14215# a_50751_n19729.t339 a_57417_n13318# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6213 a_38619_n8033# a_31953_n19727.t351 a_38097_n8930# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6214 a_36530_4481# a_30152_11614.t23 a_36008_4481.t1 VSS.t326 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6215 VSS.t731 VSS.t730 VSS.t731 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6216 a_48349_n36322# a_47819_n35156.t21 a_47819_n36322.t0 VDD.t2561 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6217 a_101641_n6055# a_71281_n8397.t322 a_96011_n36322.t0 VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6218 a_30682_13546# a_30152_10448.t22 a_30152_11614.t4 VDD.t351 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6219 a_33249_34067.t109 a_35502_25545.t97 VSS.t138 VSS.t35 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6220 VDD.t911 VDD.t910 VDD.t911 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6221 a_77776_12380# a_65658_4421.t2 a_77225_4481.t8 VDD.t2926 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6222 a_55635_12380# a_53829_10388.t23 VSS.t436 VDD.t2923 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6223 a_33249_48695.t167 a_31699_20742.t252 VDD.t277 VDD.t137 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6224 VSS.t729 VSS.t728 VSS.t729 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6225 VSS.t727 VSS.t725 VSS.t727 VSS.t726 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6226 VSS.t334 a_106830_10388.t23 a_107230_11614# VDD.t524 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6227 VDD.t909 VDD.t907 VDD.t909 VDD.t908 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6228 VDD.t906 VDD.t905 VDD.t906 VDD.t549 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6229 VDD.t904 VDD.t903 VDD.t904 VDD.t61 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6230 VDD.t902 VDD.t900 VDD.t902 VDD.t901 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6231 VSS.t724 VSS.t723 VSS.t724 VSS.t184 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X6232 VDD.t899 VDD.t898 VDD.t899 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6233 a_57977_n3550# a_50751_n19729.t340 a_57417_n3550# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6234 a_90245_n6960# a_71281_n10073.t323 a_89407_n6960# VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6235 VDD.t897 VDD.t895 VDD.t897 VDD.t896 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6236 VSS.t722 VSS.t720 VSS.t722 VSS.t721 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6237 VDD.t894 VDD.t893 VDD.t894 VDD.t629 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6238 a_112559_4481.t6 a_112559_4481.t5 a_114485_5639# VSS.t286 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6239 VSS.t719 VSS.t717 VSS.t719 VSS.t718 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6240 VSS.t185 a_41891_4481.t20 a_42413_5639# VSS.t171 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6241 a_33249_34067.t0 a_35502_24538.t63 a_52635_34067.t1 VSS.t191 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6242 VSS.t716 VSS.t715 VSS.t716 VSS.t254 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6243 VSS.t714 VSS.t713 VSS.t714 VSS.t643 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6244 a_47991_5507.t0 a_47819_11614.t20 a_54197_6405# VSS.t327 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6245 a_71896_n34390# a_71496_n36382.t18 a_71366_n35156.t1 VDD.t2254 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6246 VDD.t892 VDD.t891 VDD.t892 VDD.t315 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6247 VSS.t712 VSS.t711 VSS.t712 VSS.t209 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6248 VDD.t890 VDD.t888 VDD.t890 VDD.t889 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6249 VDD.t887 VDD.t885 VDD.t887 VDD.t886 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6250 VDD.t884 VDD.t883 VDD.t884 VDD.t316 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6251 a_83141_n14095# a_71281_n10073.t324 a_82573_n14095# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6252 a_90935_n29181# a_83153_n36322.t23 a_32913_n8930.t1 VSS.t457 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6253 a_100803_n2435# a_71281_n8397.t323 a_100235_n2435# VDD.t438 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6254 a_30682_11614# a_30152_10448.t23 a_30152_11614.t6 VDD.t351 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6255 VDD.t388 a_71281_n10073.t325 a_95105_n21335# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6256 VDD.t882 VDD.t880 VDD.t882 VDD.t881 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6257 VSS.t710 VSS.t708 VSS.t710 VSS.t709 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6258 a_33249_34067.t108 a_35502_25545.t98 VSS.t137 VSS.t44 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6259 a_88839_n3340# a_71281_n10073.t326 a_88271_n3340# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6260 a_33379_34917.t68 IN_NEG.t0 cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
X6261 a_95943_n6960# a_71281_n10073.t327 a_95105_n4245# VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6262 VDD.t879 VDD.t877 VDD.t879 VDD.t878 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6263 VSS.t136 a_35502_25545.t99 a_33249_34067.t107 VSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X6264 VSS.t707 VSS.t706 VSS.t707 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6265 VSS.t705 VSS.t703 VSS.t705 VSS.t704 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6266 VSS.t702 VSS.t701 VSS.t702 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6267 VSS.t700 VSS.t699 VSS.t700 VSS.t573 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6268 VDD.t876 VDD.t875 VDD.t876 VDD.t412 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6269 a_84547_n17715# a_71281_n10073.t328 a_84017_n16810.t1 VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6270 VSS.t698 VSS.t697 VSS.t698 VSS.t573 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6271 VSS.t696 VSS.t694 VSS.t696 VSS.t695 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6272 VSS.t693 VSS.t691 VSS.t693 VSS.t692 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6273 a_96849_n34390# a_83325_n29313.t1 a_96011_n36322.t1 VDD.t2243 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6274 OUT.t31 a_35922_19591.t174 a_52635_49681.t76 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6275 VSS.t690 VSS.t688 VSS.t690 VSS.t689 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6276 VSS.t687 VSS.t685 VSS.t687 VSS.t686 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6277 VDD.t874 VDD.t873 VDD.t874 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6278 a_33249_48695.t100 a_33379_34917.t86 a_33249_35053.t83 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6279 a_84547_n15000# a_71281_n10073.t329 a_83709_n15000# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6280 VDD.t872 VDD.t871 VDD.t872 VDD.t556 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6281 VDD.t870 VDD.t868 VDD.t870 VDD.t869 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6282 a_89009_n30339.t3 a_89163_n36382.t23 a_89563_n36322# VDD.t548 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6283 VSS.t684 VSS.t683 VSS.t684 VSS.t13 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6284 a_52635_34067.t47 a_35922_19591.t175 a_52635_48695.t7 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6285 a_71366_13546.t0 a_89163_10388.t22 a_90969_13546# VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6286 VDD.t867 VDD.t866 VDD.t867 VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6287 a_81735_n14095# a_71281_n10073.t330 a_81205_n14095.t2 VDD.t306 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6288 a_71281_n10073.t3 a_71281_n10073.t2 VDD.t487 VDD.t318 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6289 a_56895_n16009.t0 a_57977_n12421.t0 a_101392_5639# VSS.t174 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6290 VSS.t682 VSS.t680 VSS.t682 VSS.t681 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6291 VDD.t865 VDD.t864 VDD.t865 VDD.t292 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6292 VDD.t278 a_31699_20742.t253 a_33249_48695.t166 VDD.t140 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6293 VDD.t863 VDD.t862 VDD.t863 VDD.t406 pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X6294 a_94537_n21335# a_71281_n10073.t331 a_93969_n21335# VDD.t319 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6295 a_47753_n18698# a_31953_n19727.t352 a_47231_n18698# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6296 a_52635_49681.t77 a_35922_19591.t176 OUT.t30 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6297 VDD.t861 VDD.t860 VDD.t861 VDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6298 VDD.t555 a_30152_n35156.t21 a_30682_n34390# VDD.t552 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6299 VDD.t859 VDD.t857 VDD.t859 VDD.t858 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6300 VSS.t679 VSS.t678 VSS.t679 VSS.t550 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6301 VSS.t677 VSS.t675 VSS.t677 VSS.t676 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6302 VDD.t856 VDD.t854 VDD.t856 VDD.t855 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6303 a_113081_5639# a_112559_4481.t22 a_106830_10388.t5 VSS.t285 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6304 a_52585_n8932# a_50751_n19729.t341 VSS.t273 VSS.t218 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6305 a_52635_48695.t6 a_35922_19591.t177 a_52635_34067.t56 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6306 VDD.t853 VDD.t852 VDD.t853 VDD.t395 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6307 a_65486_10448.t9 a_65658_4421.t0 a_67462_5639# VSS.t413 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6308 VDD.t851 VDD.t850 VDD.t851 VDD.t52 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6309 VSS.t674 VSS.t672 VSS.t674 VSS.t673 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6310 VSS.t671 VSS.t670 VSS.t671 VSS.t614 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6311 a_111631_n19525# a_71281_n8397.t324 a_111063_n19525# VDD.t431 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6312 VDD.t849 VDD.t847 VDD.t849 VDD.t848 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6313 a_54579_n8932# a_50751_n19729.t342 a_54019_n8932# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6314 a_42413_5639# a_41891_4481.t21 a_36162_10388.t1 VSS.t177 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6315 VDD.t846 VDD.t844 VDD.t846 VDD.t845 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6316 VSS.t669 VSS.t668 VSS.t669 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6317 a_81205_n14095.t0 a_89163_10388.t23 a_90969_11614# VDD.t557 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6318 VDD.t843 VDD.t841 VDD.t843 VDD.t842 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6319 VDD.t840 VDD.t838 VDD.t840 VDD.t839 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6320 a_60285_n8035# a_50751_n19729.t343 a_59763_n8035# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6321 a_66016_n35156# a_65486_n35156.t4 a_65486_n35156.t5 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6322 VDD.t837 VDD.t835 VDD.t837 VDD.t836 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6323 VDD.t834 VDD.t833 VDD.t834 VDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6324 VSS.t667 VSS.t666 VSS.t667 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6325 a_79151_5639# a_77225_4481.t22 VSS.t346 VSS.t337 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6326 VSS.t665 VSS.t664 VSS.t665 VSS.t189 nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X6327 VDD.t832 VDD.t830 VDD.t832 VDD.t831 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6328 a_52635_49681.t78 a_35922_19591.t178 OUT.t29 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6329 VSS.t663 VSS.t662 VSS.t663 VSS.t33 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6330 VSS.t661 VSS.t660 VSS.t661 VSS.t183 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6331 VSS.t659 VSS.t657 VSS.t659 VSS.t658 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6332 a_53699_n35156.t3 a_53829_n36382.t22 a_55635_n34390# VDD.t334 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6333 VSS.t656 VSS.t654 VSS.t656 VSS.t655 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6334 VSS.t653 VSS.t651 VSS.t653 VSS.t652 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6335 VDD.t829 VDD.t828 VDD.t829 VDD.t816 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6336 a_100992_n29313.t0 a_100820_n36322.t22 a_107198_n30339# VSS.t353 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6337 VDD.t827 VDD.t825 VDD.t827 VDD.t826 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6338 VDD.t824 VDD.t823 VDD.t824 VDD.t399 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6339 VSS.t650 VSS.t648 VSS.t650 VSS.t649 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6340 a_33249_48695.t101 a_33379_34917.t87 a_33249_35053.t84 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6341 a_54197_n29181# a_47819_n36322.t23 VDD.t523 VSS.t329 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6342 VDD.t822 VDD.t820 VDD.t822 VDD.t821 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6343 VSS.t647 VSS.t645 VSS.t647 VSS.t646 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6344 VSS.t644 VSS.t642 VSS.t644 VSS.t643 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6345 VDD.t819 VDD.t818 VDD.t819 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6346 VDD.t817 VDD.t815 VDD.t817 VDD.t816 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6347 a_66016_n33224# a_65486_n35156.t6 a_65486_n35156.t7 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6348 VDD.t279 a_31699_20742.t254 a_33249_48695.t165 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6349 VDD.t814 VDD.t812 VDD.t814 VDD.t813 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6350 a_52635_34067.t57 a_35922_19591.t179 a_52635_48695.t5 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6351 OUT.t28 a_35922_19591.t180 a_52635_49681.t79 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6352 a_83141_n3340# a_71281_n10073.t332 a_82573_n3340# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6353 VDD.t811 VDD.t810 VDD.t811 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6354 a_67111_n7138# a_50751_n19729.t344 a_66551_n7138# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6355 VDD.t809 VDD.t808 VDD.t809 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6356 a_63683_n14215# a_50751_n19729.t345 a_63161_n15112# VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6357 VSS.t641 VSS.t640 VSS.t641 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6358 VDD.t807 VDD.t806 VDD.t807 VDD.t792 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6359 VSS.t639 VSS.t637 VSS.t639 VSS.t638 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6360 VSS.t636 VSS.t635 VSS.t636 VSS.t282 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6361 VDD.t805 VDD.t803 VDD.t805 VDD.t804 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6362 VDD.t802 VDD.t800 VDD.t802 VDD.t801 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6363 a_84547_n20430# a_71281_n10073.t333 a_83709_n20430# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6364 a_33249_35053.t85 a_33379_34917.t88 a_33249_48695.t102 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6365 a_53829_10388.t5 a_53699_11614.t10 a_61515_10448# VDD.t493 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6366 OUT.t27 a_35922_19591.t181 a_52635_49681.t80 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6367 VSS.t634 VSS.t633 VSS.t634 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6368 a_100235_n3340# a_71281_n8397.t325 a_99667_n3340# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6369 VSS.t632 VSS.t631 VSS.t632 VSS.t446 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6370 a_33249_48695.t152 a_33379_34007.t88 a_33249_34067.t22 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6371 a_35502_25545.t8 a_31699_20742.t255 VDD.t280 VDD.t21 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6372 a_37934_n30339# a_30152_n36322.t23 a_30324_n29313.t0 VSS.t324 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6373 a_54229_n36322# a_53829_n36382.t23 a_53699_n36322.t2 VDD.t322 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6374 a_51151_n6241# a_50751_n19729.t346 a_50629_n7138# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6375 VSS.t630 VSS.t629 VSS.t630 VSS.t149 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6376 a_49795_7563# a_47991_4421.t0 a_48951_4481.t1 VSS.t281 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6377 a_110225_n7865# a_71281_n8397.t326 a_109695_n7865# VDD.t469 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6378 a_108602_n29181# a_100820_n36322.t23 a_39179_n8930.t1 VSS.t351 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6379 a_88271_n9675# a_71281_n10073.t334 a_87433_n9675# VDD.t313 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6380 VDD.t799 VDD.t797 VDD.t799 VDD.t798 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6381 a_101641_n18620# a_71281_n8397.t327 a_100803_n18620# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6382 VDD.t796 VDD.t794 VDD.t796 VDD.t795 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6383 a_50751_n19729.t9 a_50751_n19729.t8 VSS.t215 VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6384 VSS.t628 VSS.t627 VSS.t628 VSS.t530 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6385 VDD.t793 VDD.t791 VDD.t793 VDD.t792 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6386 a_46879_n13316# a_31953_n19727.t353 a_46319_n13316# VSS.t63 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6387 VSS.t626 VSS.t625 VSS.t626 VSS.t413 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6388 a_32353_n18698# a_31953_n19727.t354 a_31831_n19595# VSS.t97 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6389 VSS.t624 VSS.t622 VSS.t624 VSS.t623 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6390 VSS.t3639 a_59558_n29181.t22 a_60080_n27257# VSS.t316 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6391 a_36032_13546.t0 a_36162_10388.t23 a_37968_10448# VDD.t1497 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6392 VDD.t790 VDD.t789 VDD.t790 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6393 VSS.t621 VSS.t619 VSS.t621 VSS.t620 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6394 a_32913_n16007.t0 a_31953_n19727.t355 a_32353_n16007# VSS.t103 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6395 VDD.t788 VDD.t787 VDD.t788 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6396 VSS.t618 VSS.t616 VSS.t618 VSS.t617 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6397 a_38619_n3548# a_31953_n19727.t356 a_38097_n4445# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6398 a_113037_n3340# a_71281_n8397.t328 a_112199_n3340# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6399 VSS.t615 VSS.t613 VSS.t615 VSS.t614 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6400 VDD.t786 VDD.t785 VDD.t786 VDD.t311 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6401 VDD.t784 VDD.t782 VDD.t784 VDD.t783 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6402 a_66016_12380# a_65486_10448.t0 a_65486_10448.t1 VDD.t2264 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6403 a_47753_n2651# a_31953_n19727.t357 a_47231_n3548# VSS.t100 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6404 a_47819_n35156.t9 a_47991_n29313.t0 a_49795_n28415# VSS.t282 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6405 a_75602_n3060# a_71266_n4019.t0 VDD.t4776 VDD.t695 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X6406 VSS.t612 VSS.t611 VSS.t612 VSS.t284 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6407 VSS.t610 VSS.t608 VSS.t610 VSS.t609 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6408 VSS.t607 VSS.t605 VSS.t607 VSS.t606 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6409 VSS.t604 VSS.t603 VSS.t604 VSS.t252 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6410 VDD.t781 VDD.t780 VDD.t781 VDD.t331 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6411 VSS.t602 VSS.t600 VSS.t602 VSS.t601 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6412 VDD.t779 VDD.t778 VDD.t779 VDD.t392 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6413 VDD.t777 VDD.t776 VDD.t777 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6414 a_73302_n35156# a_71496_n36382.t19 VSS.t370 VDD.t2814 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6415 VSS.t213 a_50751_n19729.t6 a_50751_n19729.t7 VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6416 a_65486_n35156.t1 a_65486_n35156.t0 a_67422_n34390# VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6417 a_101641_n6960# a_71281_n8397.t329 a_100803_n4245# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6418 a_96011_n36322.t2 a_89033_n35156.t12 a_95443_n36322# VDD.t2425 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6419 VSS.t599 VSS.t598 VSS.t599 VSS.t144 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6420 VDD.t775 VDD.t774 VDD.t775 VDD.t389 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X6421 OUT.t26 a_35922_19591.t182 a_52635_49681.t81 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6422 a_107339_n18620# a_71281_n8397.t330 a_106501_n18620# VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6423 VDD.t773 VDD.t772 VDD.t773 VDD.t652 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6424 OUT.t25 a_35922_19591.t183 a_52635_49681.t82 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6425 VDD.t771 VDD.t770 VDD.t771 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6426 a_60845_n13318# a_50751_n19729.t347 a_60285_n12421# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6427 a_63683_n5344# a_50751_n19729.t348 a_63161_n5344.t0 VSS.t260 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6428 a_33249_48695.t153 a_33379_34007.t89 a_33249_34067.t21 VDD.t54 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6429 a_50751_n19729.t5 a_50751_n19729.t4 VSS.t212 VSS.t211 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6430 VDD.t769 VDD.t768 VDD.t769 VDD.t63 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6431 a_83153_n36322.t1 a_32913_n8930.t1 a_85129_n29181# VSS.t365 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6432 a_50751_n19729.t3 a_50751_n19729.t2 VSS.t210 VSS.t209 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6433 VDD.t767 VDD.t766 VDD.t767 VDD.t528 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6434 VDD.t511 a_47819_11614.t21 a_55601_5639# VSS.t328 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6435 VDD.t765 VDD.t764 VDD.t765 VDD.t405 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6436 VDD.t763 VDD.t762 VDD.t763 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6437 VDD.t761 VDD.t760 VDD.t761 VDD.t79 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6438 VSS.t597 VSS.t595 VSS.t597 VSS.t596 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6439 a_57417_n19597# a_50751_n19729.t349 a_56895_n19597# VSS.t254 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6440 VDD.t759 VDD.t757 VDD.t759 VDD.t758 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6441 a_33249_48695.t103 a_33379_34917.t89 a_33249_35053.t86 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6442 VSS.t456 a_94892_n29181.t21 a_95414_n30339# VSS.t450 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6443 a_73302_n33224# a_71496_n36382.t20 a_71342_n30339.t1 VDD.t2814 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6444 VDD.t281 a_31699_20742.t256 a_35502_24538.t2 VDD.t26 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6445 VDD.t756 VDD.t755 VDD.t756 VDD.t330 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6446 VDD.t754 VDD.t753 VDD.t754 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6447 VSS.t594 VSS.t592 VSS.t594 VSS.t593 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6448 a_101392_n28415# a_39179_n8930.t1 a_100820_n36322.t4 VSS.t381 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6449 VSS.t591 VSS.t589 VSS.t591 VSS.t590 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6450 a_33249_48695.t164 a_31699_20742.t257 VDD.t282 VDD.t67 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6451 VSS.t588 VSS.t587 VSS.t588 VSS.t26 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6452 VSS.t586 VSS.t585 VSS.t586 VSS.t2 nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X6453 VDD.t4815 a_52635_34067.t233 a_52635_49681.t90 VDD.t407 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6454 VDD.t11 a_65486_n35156.t23 a_66016_n34390# VDD.t1 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6455 VDD.t752 VDD.t750 VDD.t752 VDD.t751 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6456 VSS.t584 VSS.t583 VSS.t584 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6457 VSS.t582 VSS.t580 VSS.t582 VSS.t581 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6458 a_60845_n4447# a_50751_n19729.t350 a_60285_n4447# VSS.t256 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6459 VSS.t579 VSS.t578 VSS.t579 VSS.t503 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6460 VDD.t749 VDD.t747 VDD.t749 VDD.t748 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6461 VDD.t746 VDD.t744 VDD.t746 VDD.t745 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6462 VDD.t743 VDD.t742 VDD.t743 VDD.t309 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6463 a_88839_n2435# a_71281_n10073.t335 a_88271_n2435# VDD.t320 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6464 VDD.t741 VDD.t740 VDD.t741 VDD.t426 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6465 VDD.t739 VDD.t738 VDD.t739 VDD.t313 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6466 VDD.t737 VDD.t736 VDD.t737 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6467 VDD.t735 VDD.t734 VDD.t735 VDD.t79 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6468 VSS.t577 VSS.t575 VSS.t577 VSS.t576 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6469 a_54579_n13318# a_50751_n19729.t351 a_54019_n12421# VSS.t253 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6470 a_84547_n18620# a_71281_n10073.t336 a_83709_n15905# VDD.t312 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6471 VDD.t733 VDD.t732 VDD.t733 VDD.t525 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6472 VDD.t731 VDD.t730 VDD.t731 VDD.t535 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6473 IBNOUT.t0 a_50751_n19729.t352 a_63683_n12421# VSS.t257 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6474 a_90935_7563# a_83153_11614.t23 a_83325_4421.t0 VSS.t401 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6475 VDD.t729 VDD.t727 VDD.t729 VDD.t728 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6476 VDD.t726 VDD.t725 VDD.t726 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6477 VDD.t724 VDD.t722 VDD.t724 VDD.t723 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6478 VDD.t721 VDD.t720 VDD.t721 VDD.t317 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6479 VDD.t719 VDD.t718 VDD.t719 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6480 VDD.t717 VDD.t716 VDD.t717 VDD.t402 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6481 VDD.t715 VDD.t714 VDD.t715 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6482 a_54019_n8932# a_50751_n19729.t353 a_51711_n8932# VSS.t258 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6483 VSS.t574 VSS.t572 VSS.t574 VSS.t573 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6484 a_42413_n29181# a_41891_n29181.t5 a_41891_n29181.t6 VSS.t177 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6485 VDD.t713 VDD.t712 VDD.t713 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6486 VSS.t571 VSS.t570 VSS.t571 VSS.t22 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6487 VSS.t569 VSS.t568 VSS.t569 VSS.t184 nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X6488 a_60285_n3550# a_50751_n19729.t354 a_59763_n3550# VSS.t251 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6489 a_83683_12380# a_83153_10448.t6 a_83153_10448.t7 VDD.t2776 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6490 VDD.t711 VDD.t709 VDD.t711 VDD.t710 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6491 VDD.t708 VDD.t707 VDD.t708 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6492 VSS.t567 VSS.t565 VSS.t567 VSS.t566 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6493 VDD.t706 VDD.t705 VDD.t706 VDD.t559 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6494 VDD.t283 a_31699_20742.t258 a_33249_48695.t163 VDD.t58 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6495 VSS.t564 VSS.t562 VSS.t564 VSS.t563 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6496 VSS.t561 VSS.t560 VSS.t561 VSS.t558 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6497 a_52635_48695.t4 a_35922_19591.t184 a_52635_34067.t58 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6498 a_35221_n12419# a_31953_n19727.t358 a_32913_n12419# VSS.t106 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6499 VDD.t704 VDD.t702 VDD.t704 VDD.t703 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6500 VDD.t284 a_31699_20742.t259 a_33249_48695.t162 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6501 VSS.t559 VSS.t557 VSS.t559 VSS.t558 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6502 a_66058_7563# a_64243_n1756.t1 a_65486_11614.t6 VSS.t410 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6503 OUT.t24 a_35922_19591.t185 a_52635_49681.t83 VDD.t399 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6504 VDD.t701 VDD.t699 VDD.t701 VDD.t700 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6505 VSS.t556 VSS.t554 VSS.t556 VSS.t555 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6506 a_32088_n34390# a_30152_n35156.t22 VDD.t4756 VDD.t2091 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6507 a_105365_n8770# a_71281_n8397.t331 a_104527_n8770# VDD.t428 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6508 VSS.t553 VSS.t552 VSS.t553 VSS.t214 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6509 VSS.t551 VSS.t549 VSS.t551 VSS.t550 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6510 VDD.t285 a_31699_20742.t260 a_33249_48695.t161 VDD.t73 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6511 VDD.t698 VDD.t697 VDD.t698 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6512 VDD.t4814 a_52635_34067.t234 a_52635_48695.t92 VDD.t397 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6513 a_48313_n17801# a_31953_n19727.t359 a_47753_n17801# VSS.t101 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6514 a_114485_n28415# a_112559_n29181.t22 VSS.t425 VSS.t418 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6515 a_55601_5639# a_47819_11614.t22 a_47991_5507.t0 VSS.t330 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6516 VDD.t286 a_31699_20742.t261 a_33249_48695.t160 VDD.t65 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6517 a_33249_34067.t20 a_33379_34007.t90 a_33249_48695.t154 VDD.t85 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6518 a_89163_n36382.t7 a_94892_n29181.t22 a_96818_n29181# VSS.t445 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6519 a_52635_34067.t59 a_35922_19591.t186 a_52635_48695.t3 VDD.t396 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6520 a_105933_n3340# a_71281_n8397.t332 a_105365_n3340# VDD.t441 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6521 a_57977_n12421.t1 a_50751_n19729.t355 a_57417_n12421# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6522 VDD.t696 VDD.t694 VDD.t696 VDD.t695 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X6523 a_33249_48695.t104 a_33379_34917.t90 a_33249_35053.t87 VDD.t56 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6524 VDD.t693 VDD.t691 VDD.t693 VDD.t692 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6525 VDD.t690 VDD.t688 VDD.t690 VDD.t689 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6526 VDD.t687 VDD.t685 VDD.t687 VDD.t686 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6527 VDD.t684 VDD.t682 VDD.t684 VDD.t683 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6528 VSS.t548 VSS.t547 VSS.t548 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6529 VDD.t18 a_31699_20742.t3 a_31699_20742.t4 VDD.t17 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6530 VSS.t546 VSS.t544 VSS.t546 VSS.t545 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6531 VDD.t681 VDD.t679 VDD.t681 VDD.t680 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6532 a_57977_n3550# a_50751_n19729.t356 a_57417_n2653# VSS.t259 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6533 VSS.t543 VSS.t541 VSS.t543 VSS.t542 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6534 VSS.t540 VSS.t538 VSS.t540 VSS.t539 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6535 VDD.t678 VDD.t676 VDD.t678 VDD.t677 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6536 VDD.t423 a_71281_n8397.t2 a_71281_n8397.t3 VDD.t422 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6537 VDD.t675 VDD.t674 VDD.t675 VDD.t293 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6538 OUT.t23 a_35922_19591.t187 a_52635_49681.t84 VDD.t391 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6539 VSS.t537 VSS.t535 VSS.t537 VSS.t536 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6540 a_47819_n35156.t1 a_47819_n35156.t0 a_49755_n36322# VDD.t2328 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6541 a_52635_34067.t60 a_35922_19591.t188 a_52635_48695.t2 VDD.t392 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6542 a_51151_n1756# a_50751_n19729.t357 a_50629_n2653# VSS.t255 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6543 VSS.t534 VSS.t532 VSS.t534 VSS.t533 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6544 VDD.t673 VDD.t672 VDD.t673 VDD.t13 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6545 VSS.t531 VSS.t529 VSS.t531 VSS.t530 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6546 VSS.t528 VSS.t526 VSS.t528 VSS.t527 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6547 VSS.t525 VSS.t524 VSS.t525 VSS.t63 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6548 a_83141_n2435# a_71281_n10073.t337 a_82573_n2435# VDD.t314 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6549 VSS.t523 VSS.t522 VSS.t523 VSS.t254 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6550 a_52635_34067.t48 a_35922_19591.t189 a_52635_48695.t1 VDD.t393 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6551 a_53145_n2653# a_50751_n19729.t358 a_52585_n1756# VSS.t214 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6552 VDD.t671 VDD.t669 VDD.t671 VDD.t670 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6553 VDD.t668 VDD.t667 VDD.t668 VDD.t494 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6554 VSS.t521 VSS.t520 VSS.t521 VSS.t483 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6555 a_52635_49681.t85 a_35922_19591.t190 OUT.t22 VDD.t394 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6556 a_83683_n35156# a_83153_n35156.t2 a_83153_n35156.t3 VDD.t2731 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6557 a_100235_n2435# a_71281_n8397.t333 a_99667_n2435# VDD.t443 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6558 VDD.t666 VDD.t664 VDD.t666 VDD.t665 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6559 VDD.t4813 a_52635_34067.t235 a_52635_49681.t89 VDD.t414 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6560 VSS.t519 VSS.t518 VSS.t519 VSS.t324 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6561 a_71366_n35156.t4 a_71496_n36382.t21 a_73302_n34390# VDD.t2061 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6562 VSS.t517 VSS.t516 VSS.t517 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6563 VDD.t663 VDD.t662 VDD.t663 VDD.t642 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6564 VSS.t515 VSS.t513 VSS.t515 VSS.t514 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6565 VSS.t512 VSS.t510 VSS.t512 VSS.t511 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6566 a_33249_35053.t108 a_35502_25545.t100 VSS.t135 VSS.t134 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6567 a_52635_48695.t91 a_52635_34067.t236 VDD.t4812 VDD.t410 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6568 a_52635_48695.t90 a_52635_34067.t237 VDD.t4811 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6569 VDD.t661 VDD.t659 VDD.t661 VDD.t660 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6570 VDD.t519 a_47819_10448.t22 a_48349_10448# VDD.t512 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6571 a_33249_48695.t159 a_31699_20742.t262 VDD.t287 VDD.t71 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6572 a_66551_n8932# a_50751_n19729.t359 a_64243_n8932# VSS.t250 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6573 VDD.t658 VDD.t656 VDD.t658 VDD.t657 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6574 VSS.t133 a_35502_25545.t101 a_33249_34067.t106 VSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X6575 VSS.t509 VSS.t508 VSS.t509 VSS.t298 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6576 a_60080_n29181# a_59558_n29181.t6 a_59558_n29181.t7 VSS.t313 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6577 VSS.t507 VSS.t505 VSS.t507 VSS.t506 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6578 VSS.t504 VSS.t502 VSS.t504 VSS.t503 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6579 a_101641_n17715# a_71281_n8397.t334 a_101111_n17715.t1 VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6580 VDD.t4807 a_47819_n35156.t22 a_48349_n36322# VDD.t2291 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6581 VDD.t655 VDD.t654 VDD.t655 VDD.t623 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6582 VSS.t501 VSS.t499 VSS.t501 VSS.t500 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6583 a_33249_35053.t94 a_35502_24538.t64 OUT.t2 VSS.t191 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6584 a_52635_49681.t86 a_35922_19591.t191 OUT.t21 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6585 VSS.t498 VSS.t497 VSS.t498 VSS.t350 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6586 VDD.t653 VDD.t651 VDD.t653 VDD.t652 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6587 a_78344_n36322.t2 a_71366_n35156.t12 a_77776_n34390# VDD.t2046 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6588 VDD.t650 VDD.t649 VDD.t650 VDD.t390 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6589 VSS.t496 VSS.t494 VSS.t496 VSS.t495 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6590 a_83683_n33224# a_83153_n35156.t4 a_83153_n35156.t5 VDD.t2731 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6591 VSS.t493 VSS.t491 VSS.t493 VSS.t492 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6592 VDD.t648 VDD.t646 VDD.t648 VDD.t647 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6593 a_33249_48695.t155 a_33379_34007.t91 a_33249_34067.t19 VDD.t76 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6594 VDD.t645 VDD.t644 VDD.t645 VDD.t69 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6595 VSS.t490 VSS.t488 VSS.t490 VSS.t489 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X6596 VDD.t643 VDD.t641 VDD.t643 VDD.t642 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6597 VDD.t640 VDD.t638 VDD.t640 VDD.t639 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6598 VSS.t487 VSS.t485 VSS.t487 VSS.t486 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6599 VSS.t484 VSS.t482 VSS.t484 VSS.t483 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6600 a_65486_n36322.t5 a_45445_n19595.t1 a_67462_n27257# VSS.t413 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6601 VSS.t481 VSS.t479 VSS.t481 VSS.t480 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6602 a_67111_n17803# a_50751_n19729.t360 a_66551_n16906# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6603 VDD.t637 VDD.t636 VDD.t637 VDD.t602 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6604 VDD.t635 VDD.t633 VDD.t635 VDD.t634 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6605 VSS.t371 a_71496_n36382.t22 a_71896_n34390# VDD.t2023 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6606 a_113037_n3340# a_71281_n8397.t335 a_112199_n2435# VDD.t471 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6607 VDD.t632 VDD.t631 VDD.t632 VDD.t397 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6608 a_33249_48695.t105 a_33379_34917.t91 a_33249_35053.t88 VDD.t99 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6609 VDD.t630 VDD.t628 VDD.t630 VDD.t629 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6610 a_52635_34067.t39 a_35922_19591.t192 a_52635_48695.t0 VDD.t395 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6611 VDD.t627 VDD.t625 VDD.t627 VDD.t626 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6612 VDD.t624 VDD.t622 VDD.t624 VDD.t623 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6613 a_71896_n36322# a_71496_n36382.t23 a_71366_n36322.t2 VDD.t2254 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6614 VDD.t621 VDD.t619 VDD.t621 VDD.t620 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6615 a_33249_48695.t158 a_31699_20742.t263 VDD.t288 VDD.t79 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6616 VSS.t478 VSS.t476 VSS.t478 VSS.t477 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6617 VDD.t4810 a_52635_34067.t238 a_52635_49681.t88 VDD.t408 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6618 VSS.t208 a_50751_n19729.t0 a_50751_n19729.t1 VSS.t207 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6619 VSS.t475 VSS.t474 VSS.t475 VSS.t155 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6620 VDD.t618 VDD.t616 VDD.t618 VDD.t617 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6621 a_33249_48695.t157 a_31699_20742.t264 VDD.t289 VDD.t61 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6622 VDD.t615 VDD.t613 VDD.t615 VDD.t614 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6623 a_95443_10448# a_83325_4421.t1 a_94892_4481.t8 VDD.t500 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6624 VDD.t612 VDD.t611 VDD.t612 VDD.t490 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6625 VDD.t610 VDD.t609 VDD.t610 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6626 VDD.t4809 a_52635_34067.t239 a_52635_48695.t89 VDD.t411 pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6627 VDD.t608 VDD.t606 VDD.t608 VDD.t607 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6628 VDD.t605 VDD.t604 VDD.t605 VDD.t67 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6629 a_107339_n17715# a_71281_n8397.t336 a_106809_n17715.t1 VDD.t467 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6630 VDD.t603 VDD.t601 VDD.t603 VDD.t602 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6631 a_94892_n29181.t8 a_83325_n29313.t1 a_96849_n34390# VDD.t1998 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6632 a_38619_n16904# a_31953_n19727.t360 a_38097_n17801# VSS.t94 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6633 a_31699_20742.t2 a_31699_20742.t1 VDD.t16 VDD.t15 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6634 a_36162_10388.t0 a_41891_4481.t22 a_43817_6405# VSS.t181 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6635 VDD.t600 VDD.t599 VDD.t600 VDD.t296 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6636 VDD.t598 VDD.t596 VDD.t598 VDD.t597 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6637 VSS.t473 VSS.t471 VSS.t473 VSS.t472 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6638 VSS.t470 VSS.t468 VSS.t470 VSS.t469 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6639 a_96849_n36322# a_83325_n29313.t1 a_96011_n36322.t2 VDD.t2243 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6640 VDD.t595 VDD.t594 VDD.t595 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6641 a_54197_7563# a_47819_11614.t23 a_53675_7563.t1 VSS.t329 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6642 VDD.t593 VDD.t592 VDD.t593 VDD.t332 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6643 a_71266_n4019.t0 I1N.t17 a_75585_n10073# VSS.t301 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X6644 VSS.t467 VSS.t466 VSS.t467 VSS.t145 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6645 a_31953_n19727.t3 a_31953_n19727.t2 VSS.t55 VSS.t54 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6646 VSS.t465 VSS.t463 VSS.t465 VSS.t464 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6647 a_59558_n29181.t3 a_59558_n29181.t2 a_61484_n28415# VSS.t312 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6648 VSS.t141 a_35502_25545.t102 a_33249_35053.t107 VSS.t18 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6649 a_33249_48695.t156 a_33379_34007.t92 a_33249_34067.t18 VDD.t63 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6650 a_67111_n7138# a_50751_n19729.t361 a_66551_n6241# VSS.t252 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6651 VDD.t591 VDD.t589 VDD.t591 VDD.t590 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6652 VDD.t588 VDD.t586 VDD.t588 VDD.t587 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6653 VDD.t585 VDD.t584 VDD.t585 VDD.t373 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6654 a_33249_35053.t106 a_35502_25545.t103 VSS.t143 VSS.t142 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6655 VDD.t583 VDD.t582 VDD.t583 VDD.t438 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6656 a_52635_49681.t87 a_35922_19591.t193 OUT.t20 VDD.t402 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6657 VDD.t581 VDD.t580 VDD.t581 VDD.t544 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6658 VDD.t4755 a_65486_10448.t22 a_66016_10448# VDD.t1341 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6659 VDD.t553 a_30152_n35156.t23 a_30682_n36322# VDD.t552 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6660 VDD.t579 VDD.t577 VDD.t579 VDD.t578 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6661 VSS.t53 a_31953_n19727.t0 a_31953_n19727.t1 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6662 VDD.t576 VDD.t574 VDD.t576 VDD.t575 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6663 VDD.t573 VDD.t571 VDD.t573 VDD.t572 pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X6664 VDD.t570 VDD.t569 VDD.t570 VDD.t398 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6665 a_101111_n17715.t0 a_71281_n8397.t337 a_100803_n21335# VDD.t473 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6666 VSS.t462 VSS.t461 VSS.t462 VSS.t105 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6667 VDD.t4808 a_52635_34067.t240 a_52635_48695.t88 VDD.t405 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6668 VDD.t568 VDD.t566 VDD.t568 VDD.t567 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6669 a_35781_n13316# a_31953_n19727.t361 a_35221_n13316# VSS.t105 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6670 VDD.t565 VDD.t563 VDD.t565 VDD.t564 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6671 VDD.t562 VDD.t560 VDD.t562 VDD.t561 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
R0 VSS.n11299 VSS.n132 320062
R1 VSS.n10846 VSS.n10697 144034
R2 VSS.n11300 VSS.n11299 49361.9
R3 VSS.n9304 VSS.n9302 17249
R4 VSS.n10287 VSS.n132 12232.4
R5 VSS.n10697 VSS.n10287 9171.32
R6 VSS.n10861 VSS.n244 3502.89
R7 VSS.n11301 VSS.t768 757.145
R8 VSS.n11296 VSS.n11293 752.225
R9 VSS.n11285 VSS.n11280 752.225
R10 VSS.n563 VSS.n562 752.225
R11 VSS.n10065 VSS.n512 752.225
R12 VSS.n9891 VSS.n644 752.225
R13 VSS.n10116 VSS.n440 752.225
R14 VSS.n139 VSS.n135 752.225
R15 VSS.n11278 VSS.n144 752.225
R16 VSS.n568 VSS.n564 752.225
R17 VSS.n1181 VSS.n510 752.225
R18 VSS.n9765 VSS.n646 752.225
R19 VSS.n1235 VSS.n438 752.225
R20 VSS.n11296 VSS.n136 750.567
R21 VSS.n11285 VSS.n145 750.567
R22 VSS.n10033 VSS.n562 750.567
R23 VSS.n512 VSS.n508 750.567
R24 VSS.n9891 VSS.n645 750.567
R25 VSS.n440 VSS.n436 750.567
R26 VSS.n11291 VSS.n135 750.567
R27 VSS.n149 VSS.n144 750.567
R28 VSS.n10031 VSS.n568 750.567
R29 VSS.n1181 VSS.n509 750.567
R30 VSS.n9767 VSS.n646 750.567
R31 VSS.n1235 VSS.n437 750.567
R32 VSS.n11293 VSS.n137 750.383
R33 VSS.n11280 VSS.n146 750.383
R34 VSS.n563 VSS.n561 750.383
R35 VSS.n10065 VSS.n511 750.383
R36 VSS.n9522 VSS.n644 750.383
R37 VSS.n10116 VSS.n439 750.383
R38 VSS.n11290 VSS.n139 750.383
R39 VSS.n11278 VSS.n150 750.383
R40 VSS.n567 VSS.n564 750.383
R41 VSS.n9888 VSS.n510 750.383
R42 VSS.n9765 VSS.n797 750.383
R43 VSS.n1389 VSS.n438 750.383
R44 VSS.n137 VSS.n136 748.725
R45 VSS.n146 VSS.n145 748.725
R46 VSS.n10033 VSS.n561 748.725
R47 VSS.n511 VSS.n508 748.725
R48 VSS.n9522 VSS.n645 748.725
R49 VSS.n439 VSS.n436 748.725
R50 VSS.n11291 VSS.n11290 748.725
R51 VSS.n150 VSS.n149 748.725
R52 VSS.n10031 VSS.n567 748.725
R53 VSS.n9888 VSS.n509 748.725
R54 VSS.n9767 VSS.n797 748.725
R55 VSS.n1389 VSS.n437 748.725
R56 VSS.n9464 VSS.n1381 697.422
R57 VSS.n9466 VSS.n1382 693.922
R58 VSS.n9464 VSS.n1382 693.645
R59 VSS.n9466 VSS.n1381 688.856
R60 VSS.t822 VSS.n10847 684.903
R61 VSS.n10598 VSS.n10344 661.869
R62 VSS.n10695 VSS.n10289 661.869
R63 VSS.n10664 VSS.n10340 661.869
R64 VSS.n10661 VSS.n10343 656.895
R65 VSS.n10603 VSS.n10288 656.895
R66 VSS.n10342 VSS.n10341 656.895
R67 VSS.n10661 VSS.n10344 656.434
R68 VSS.n10603 VSS.n10289 656.434
R69 VSS.n10664 VSS.n10341 656.434
R70 VSS.n10598 VSS.n10343 653.672
R71 VSS.n10695 VSS.n10288 653.672
R72 VSS.n10342 VSS.n10340 653.672
R73 VSS.n10849 VSS.n10848 613.597
R74 VSS.n11302 VSS.n130 531.539
R75 VSS.n10845 VSS.n130 530.25
R76 VSS.n11302 VSS.n131 530.067
R77 VSS.n10845 VSS.n131 528.777
R78 VSS.n11346 VSS.n8 523.342
R79 VSS.n11360 VSS.n95 523.342
R80 VSS.n10983 VSS.n183 523.342
R81 VSS.n10928 VSS.n220 523.342
R82 VSS.n867 VSS.n505 523.342
R83 VSS.n9562 VSS.n835 523.342
R84 VSS.n11375 VSS.n5 523.342
R85 VSS.n11362 VSS.n92 523.342
R86 VSS.n10981 VSS.n180 523.342
R87 VSS.n10930 VSS.n216 523.342
R88 VSS.n1185 VSS.n1153 523.342
R89 VSS.n9541 VSS.n832 523.342
R90 VSS.n9528 VSS.n9527 523.342
R91 VSS.n9421 VSS.n1395 523.342
R92 VSS.n432 VSS.n431 523.342
R93 VSS.n10122 VSS.n421 523.342
R94 VSS.n420 VSS.n393 523.342
R95 VSS.n362 VSS.n361 523.342
R96 VSS.n10182 VSS.n349 523.342
R97 VSS.n348 VSS.n321 523.342
R98 VSS.n290 VSS.n289 523.342
R99 VSS.n10242 VSS.n277 523.342
R100 VSS.n276 VSS.n251 523.342
R101 VSS.n9117 VSS.n1532 523.342
R102 VSS.n9093 VSS.n1537 523.342
R103 VSS.n9009 VSS.n1563 523.342
R104 VSS.n9348 VSS.n1482 523.342
R105 VSS.n9298 VSS.n1507 523.342
R106 VSS.n9250 VSS.n1515 523.342
R107 VSS.n9176 VSS.n1525 523.342
R108 VSS.n11467 VSS.n7 521.869
R109 VSS.n11037 VSS.n94 521.869
R110 VSS.n11151 VSS.n182 521.869
R111 VSS.n547 VSS.n219 521.869
R112 VSS.n10068 VSS.n504 521.869
R113 VSS.n9563 VSS.n834 521.869
R114 VSS.n11469 VSS.n4 521.869
R115 VSS.n11263 VSS.n91 521.869
R116 VSS.n11153 VSS.n179 521.869
R117 VSS.n693 VSS.n215 521.869
R118 VSS.n9559 VSS.n507 521.869
R119 VSS.n9565 VSS.n831 521.869
R120 VSS.n1222 VSS.n435 521.869
R121 VSS.n9381 VSS.n1384 521.869
R122 VSS.n10120 VSS.n10119 521.869
R123 VSS.n10127 VSS.n422 521.869
R124 VSS.n10175 VSS.n394 521.869
R125 VSS.n10180 VSS.n10179 521.869
R126 VSS.n10187 VSS.n350 521.869
R127 VSS.n10235 VSS.n322 521.869
R128 VSS.n10240 VSS.n10239 521.869
R129 VSS.n10247 VSS.n278 521.869
R130 VSS.n10285 VSS.n252 521.869
R131 VSS.n9111 VSS.n1531 521.869
R132 VSS.n9090 VSS.n1555 521.869
R133 VSS.n9014 VSS.n1562 521.869
R134 VSS.n9345 VSS.n1497 521.869
R135 VSS.n9308 VSS.n1506 521.869
R136 VSS.n9247 VSS.n1514 521.869
R137 VSS.n9181 VSS.n1524 521.869
R138 VSS.n11346 VSS.n7 519.659
R139 VSS.n11360 VSS.n94 519.659
R140 VSS.n10983 VSS.n182 519.659
R141 VSS.n10928 VSS.n219 519.659
R142 VSS.n867 VSS.n504 519.659
R143 VSS.n835 VSS.n834 519.659
R144 VSS.n11375 VSS.n4 519.659
R145 VSS.n11362 VSS.n91 519.659
R146 VSS.n10981 VSS.n179 519.659
R147 VSS.n10930 VSS.n215 519.659
R148 VSS.n9559 VSS.n1153 519.659
R149 VSS.n9541 VSS.n831 519.659
R150 VSS.n9528 VSS.n1222 519.659
R151 VSS.n9421 VSS.n1384 519.659
R152 VSS.n10120 VSS.n431 519.659
R153 VSS.n10127 VSS.n421 519.659
R154 VSS.n10175 VSS.n393 519.659
R155 VSS.n10180 VSS.n361 519.659
R156 VSS.n10187 VSS.n349 519.659
R157 VSS.n10235 VSS.n321 519.659
R158 VSS.n10240 VSS.n289 519.659
R159 VSS.n10247 VSS.n277 519.659
R160 VSS.n10285 VSS.n251 519.659
R161 VSS.n9111 VSS.n1532 519.659
R162 VSS.n9093 VSS.n1555 519.659
R163 VSS.n9009 VSS.n1562 519.659
R164 VSS.n9348 VSS.n1497 519.659
R165 VSS.n9298 VSS.n1506 519.659
R166 VSS.n9250 VSS.n1514 519.659
R167 VSS.n9176 VSS.n1524 519.659
R168 VSS.n11467 VSS.n8 516.342
R169 VSS.n11037 VSS.n95 516.342
R170 VSS.n11151 VSS.n183 516.342
R171 VSS.n547 VSS.n220 516.342
R172 VSS.n10068 VSS.n505 516.342
R173 VSS.n9563 VSS.n9562 516.342
R174 VSS.n11469 VSS.n5 516.342
R175 VSS.n11263 VSS.n92 516.342
R176 VSS.n11153 VSS.n180 516.342
R177 VSS.n693 VSS.n216 516.342
R178 VSS.n1185 VSS.n507 516.342
R179 VSS.n9565 VSS.n832 516.342
R180 VSS.n9527 VSS.n435 516.342
R181 VSS.n9381 VSS.n1395 516.342
R182 VSS.n10119 VSS.n432 516.342
R183 VSS.n10122 VSS.n422 516.342
R184 VSS.n420 VSS.n394 516.342
R185 VSS.n10179 VSS.n362 516.342
R186 VSS.n10182 VSS.n350 516.342
R187 VSS.n348 VSS.n322 516.342
R188 VSS.n10239 VSS.n290 516.342
R189 VSS.n10242 VSS.n278 516.342
R190 VSS.n276 VSS.n252 516.342
R191 VSS.n9117 VSS.n1531 516.342
R192 VSS.n9090 VSS.n1537 516.342
R193 VSS.n9014 VSS.n1563 516.342
R194 VSS.n9345 VSS.n1482 516.342
R195 VSS.n9308 VSS.n1507 516.342
R196 VSS.n9247 VSS.n1515 516.342
R197 VSS.n9181 VSS.n1525 516.342
R198 VSS.t2 VSS.t1082 412.349
R199 VSS.t126 VSS.t847 412.349
R200 VSS.n10848 VSS.t822 407.188
R201 VSS.t768 VSS.n11300 407.188
R202 VSS.n10851 VSS.n249 383.618
R203 VSS.n10852 VSS.n10851 381.962
R204 VSS.n249 VSS.n248 381.132
R205 VSS.n10852 VSS.n248 379.474
R206 VSS.t1600 VSS.t189 362.154
R207 VSS.t184 VSS.t1827 358.87
R208 VSS.t414 VSS.t861 303.373
R209 VSS.t415 VSS.t910 303.373
R210 VSS.t901 VSS.t350 303.373
R211 VSS.t352 VSS.t1472 303.373
R212 VSS.t382 VSS.t949 303.373
R213 VSS.t762 VSS.t381 303.373
R214 VSS.t777 VSS.t445 303.373
R215 VSS.t446 VSS.t1366 303.269
R216 VSS.t896 VSS.t460 303.269
R217 VSS.t459 VSS.t576 303.269
R218 VSS.t819 VSS.t365 303.269
R219 VSS.t367 VSS.t726 303.269
R220 VSS.t1116 VSS.t1003 300.337
R221 VSS.t469 VSS.t398 300.337
R222 VSS.t400 VSS.t882 300.337
R223 VSS.t297 VSS.t813 300.337
R224 VSS.t299 VSS.t695 300.337
R225 VSS.t286 VSS.t1299 300.236
R226 VSS.t709 VSS.t285 300.236
R227 VSS.t649 VSS.t151 300.236
R228 VSS.t150 VSS.t506 300.236
R229 VSS.t173 VSS.t492 300.236
R230 VSS.t175 VSS.t765 300.236
R231 VSS.t1349 VSS.t816 296.584
R232 VSS.n10858 VSS.n243 267.474
R233 VSS.n10862 VSS.n243 266.829
R234 VSS.n10858 VSS.n242 266.276
R235 VSS.n10862 VSS.n242 265.632
R236 VSS.t20 VSS.t2 262.702
R237 VSS.t37 VSS.t126 262.702
R238 VSS.t336 VSS.t858 256.925
R239 VSS.t745 VSS.t427 256.925
R240 VSS.t428 VSS.t609 256.925
R241 VSS.n9302 VSS.t1391 248.619
R242 VSS.n1564 VSS.n132 244.691
R243 VSS.n10287 VSS.n10286 242.161
R244 VSS.n10861 VSS.t1600 219.544
R245 VSS.t1827 VSS.n10859 219.544
R246 VSS.t1082 VSS.n245 219.544
R247 VSS.t847 VSS.n10849 219.544
R248 VSS.n10697 VSS.n10696 215.996
R249 VSS.t861 VSS.t617 206.678
R250 VSS.t418 VSS.t414 206.678
R251 VSS.t416 VSS.t415 206.678
R252 VSS.t910 VSS.t1261 206.678
R253 VSS.t981 VSS.t901 206.678
R254 VSS.t350 VSS.t351 206.678
R255 VSS.t353 VSS.t352 206.678
R256 VSS.t1472 VSS.t623 206.678
R257 VSS.t949 VSS.t984 206.678
R258 VSS.t383 VSS.t382 206.678
R259 VSS.t381 VSS.t384 206.678
R260 VSS.t942 VSS.t762 206.678
R261 VSS.t1543 VSS.t777 206.678
R262 VSS.t450 VSS.t446 206.607
R263 VSS.t1366 VSS.t550 206.607
R264 VSS.t539 VSS.t896 206.607
R265 VSS.t460 VSS.t457 206.607
R266 VSS.t458 VSS.t459 206.607
R267 VSS.t576 VSS.t1320 206.607
R268 VSS.t1039 VSS.t819 206.607
R269 VSS.t365 VSS.t278 206.607
R270 VSS.t366 VSS.t367 206.607
R271 VSS.t726 VSS.t652 206.607
R272 VSS.t673 VSS.t889 206.607
R273 VSS.t445 VSS.t447 205.131
R274 VSS.t1308 VSS.t1349 204.609
R275 VSS.t1003 VSS.t1042 204.609
R276 VSS.t681 VSS.t1116 204.609
R277 VSS.t864 VSS.t469 204.609
R278 VSS.t398 VSS.t401 204.609
R279 VSS.t399 VSS.t400 204.609
R280 VSS.t882 VSS.t1131 204.609
R281 VSS.t813 VSS.t842 204.609
R282 VSS.t298 VSS.t297 204.609
R283 VSS.t300 VSS.t299 204.609
R284 VSS.t695 VSS.t952 204.609
R285 VSS.t1391 VSS.t1432 204.609
R286 VSS.t1299 VSS.t1030 204.541
R287 VSS.t290 VSS.t286 204.541
R288 VSS.t285 VSS.t287 204.541
R289 VSS.t689 VSS.t709 204.541
R290 VSS.t780 VSS.t649 204.541
R291 VSS.t151 VSS.t147 204.541
R292 VSS.t188 VSS.t150 204.541
R293 VSS.t506 VSS.t464 204.541
R294 VSS.t492 VSS.t1311 204.541
R295 VSS.t144 VSS.t173 204.541
R296 VSS.t174 VSS.t175 204.541
R297 VSS.t765 VSS.t797 204.541
R298 VSS.t816 VSS.t555 204.541
R299 VSS.n10850 VSS.t37 194.681
R300 VSS.n10850 VSS.t20 186.238
R301 VSS.t335 VSS.t337 175.035
R302 VSS.t341 VSS.t336 175.035
R303 VSS.t858 VSS.t646 175.035
R304 VSS.t753 VSS.t745 175.035
R305 VSS.t427 VSS.t426 175.035
R306 VSS.t429 VSS.t428 175.035
R307 VSS.t609 VSS.t1292 175.035
R308 VSS.t617 VSS.n1564 172.355
R309 VSS.t1261 VSS.n9012 172.355
R310 VSS.n9011 VSS.t981 172.355
R311 VSS.t623 VSS.n1533 172.355
R312 VSS.t984 VSS.n9112 172.355
R313 VSS.n9116 VSS.t942 172.355
R314 VSS.n9115 VSS.t1543 172.355
R315 VSS.t550 VSS.n9179 172.296
R316 VSS.n9178 VSS.t539 172.296
R317 VSS.t1320 VSS.n1517 172.296
R318 VSS.n1516 VSS.t1039 172.296
R319 VSS.t652 VSS.n9306 172.296
R320 VSS.n9305 VSS.t673 172.296
R321 VSS.n353 VSS.t681 170.631
R322 VSS.n10186 VSS.t864 170.631
R323 VSS.t1131 VSS.n10183 170.631
R324 VSS.t842 VSS.n354 170.631
R325 VSS.t952 VSS.n10177 170.631
R326 VSS.n10176 VSS.t1432 170.631
R327 VSS.n10286 VSS.t1030 170.572
R328 VSS.n281 VSS.t689 170.572
R329 VSS.n10246 VSS.t780 170.572
R330 VSS.t464 VSS.n10243 170.572
R331 VSS.t1311 VSS.n282 170.572
R332 VSS.t797 VSS.n10237 170.572
R333 VSS.n10236 VSS.t555 170.572
R334 VSS.t18 VSS.t601 163.815
R335 VSS.t24 VSS.t1109 163.815
R336 VSS.t9 VSS.t44 159.155
R337 VSS.t7 VSS.t142 159.155
R338 VSS.t889 VSS.n9304 158.827
R339 VSS.n9010 VSS.t418 148.365
R340 VSS.n9092 VSS.t351 148.365
R341 VSS.n9113 VSS.t383 148.365
R342 VSS.n9177 VSS.t447 148.315
R343 VSS.n9249 VSS.t457 148.315
R344 VSS.n9299 VSS.t278 148.315
R345 VSS.n351 VSS.t1308 146.881
R346 VSS.t401 VSS.n10185 146.881
R347 VSS.n392 VSS.t298 146.881
R348 VSS.n279 VSS.t290 146.832
R349 VSS.t147 VSS.n10245 146.832
R350 VSS.n320 VSS.t144 146.832
R351 VSS.t646 VSS.n423 145.966
R352 VSS.n10126 VSS.t753 145.966
R353 VSS.t1292 VSS.n10123 145.966
R354 VSS.t0 VSS.t1621 145.738
R355 VSS.t704 VSS.t191 145.738
R356 VSS.n9013 VSS.t416 144.674
R357 VSS.n9091 VSS.t353 144.674
R358 VSS.t384 VSS.n9114 144.674
R359 VSS.n9180 VSS.t450 144.625
R360 VSS.n9248 VSS.t458 144.625
R361 VSS.n9307 VSS.t366 144.625
R362 VSS.t1042 VSS.n352 143.227
R363 VSS.n10184 VSS.t399 143.227
R364 VSS.n10178 VSS.t300 143.227
R365 VSS.t287 VSS.n280 143.179
R366 VSS.n10244 VSS.t188 143.179
R367 VSS.n10238 VSS.t174 143.179
R368 VSS.t187 VSS.t35 142.941
R369 VSS.t183 VSS.t13 142.941
R370 VSS.n10860 VSS.t184 134.636
R371 VSS.n10847 VSS.n10846 132.153
R372 VSS.t189 VSS.n10860 128.067
R373 VSS.t337 VSS.n9301 125.65
R374 VSS.t426 VSS.n10125 125.65
R375 VSS.n9300 VSS.t341 122.525
R376 VSS.n10124 VSS.t429 122.525
R377 VSS.n1391 VSS.n424 122.525
R378 VSS.n9116 VSS.n9115 116.626
R379 VSS.n9306 VSS.n9305 116.585
R380 VSS.n10177 VSS.n10176 115.459
R381 VSS.n10237 VSS.n10236 115.419
R382 VSS.t385 VSS.t480 106.296
R383 VSS.t527 VSS.t153 106.296
R384 VSS.t49 VSS.t18 104.365
R385 VSS.t44 VSS.t49 104.365
R386 VSS.t11 VSS.t9 104.365
R387 VSS.t142 VSS.t4 104.365
R388 VSS.t4 VSS.t24 104.365
R389 VSS.n10662 VSS.t7 100.638
R390 VSS.t163 VSS.t22 88.1506
R391 VSS.t166 VSS.t15 88.1506
R392 VSS.n10696 VSS.t601 87.2188
R393 VSS.t1109 VSS.n244 87.2188
R394 VSS.t40 VSS.t159 86.287
R395 VSS.t134 VSS.t182 86.287
R396 VSS.t530 VSS.t26 83.4915
R397 VSS.n10600 VSS.t514 82.3733
R398 VSS.n9012 VSS.n9011 81.5642
R399 VSS.n9179 VSS.n9178 81.5364
R400 VSS.n10186 VSS.n353 80.7481
R401 VSS.n10246 VSS.n281 80.7209
R402 VSS.n10847 VSS.t362 75.9965
R403 VSS.t33 VSS.n10599 73.8006
R404 VSS.n10602 VSS.t162 73.8006
R405 VSS.t390 VSS.t385 72.4152
R406 VSS.n9465 VSS.t154 72.4152
R407 VSS.t1227 VSS.t527 72.4152
R408 VSS.t303 VSS.t1437 69.1825
R409 VSS.n10126 VSS.n423 69.0763
R410 VSS.n10859 VSS.n245 67.5525
R411 VSS.t558 VSS.t145 65.5106
R412 VSS.t386 VSS.n9303 63.4927
R413 VSS.t255 VSS.t282 63.4385
R414 VSS.t658 VSS.n1499 60.3892
R415 VSS.t326 VSS.t105 59.6927
R416 VSS.n1498 VSS.t1800 56.1219
R417 VSS.t313 VSS.t211 53.3171
R418 VSS.n9112 VSS.n1533 53.1461
R419 VSS.n1517 VSS.n1516 53.128
R420 VSS.n10183 VSS.n354 52.6143
R421 VSS.n10243 VSS.n282 52.5966
R422 VSS.n9347 VSS.t387 51.9839
R423 VSS.t156 VSS.n9422 51.9839
R424 VSS.n1394 VSS.t489 51.9839
R425 VSS.t258 VSS.t503 51.3247
R426 VSS.t155 VSS.n1383 50.6908
R427 VSS.t573 VSS.t103 47.579
R428 VSS.n10123 VSS.n424 45.0092
R429 VSS.n9346 VSS.t1249 44.8718
R430 VSS.t593 VSS.t533 44.6302
R431 VSS.t873 VSS.t614 44.6302
R432 VSS.t284 VSS.t283 44.6302
R433 VSS.t100 VSS.t101 44.6302
R434 VSS.t563 VSS.t1258 44.6302
R435 VSS.t686 VSS.t913 44.6302
R436 VSS.t96 VSS.t94 44.6302
R437 VSS.t323 VSS.t324 44.6302
R438 VSS.t839 VSS.t558 44.6302
R439 VSS.t153 VSS.t302 43.8373
R440 VSS.t249 VSS.t483 42.5581
R441 VSS.t750 VSS.t412 42.0799
R442 VSS.t480 VSS.t2042 41.639
R443 VSS.n1393 VSS.n1392 41.639
R444 VSS.t566 VSS.t177 40.8845
R445 VSS.t99 VSS.t181 40.486
R446 VSS.t250 VSS.t410 39.2906
R447 VSS.t495 VSS.t106 38.8124
R448 VSS.t305 VSS.t156 38.1476
R449 VSS.t511 VSS.n9524 37.2982
R450 VSS.t545 VSS.n1182 37.2982
R451 VSS.n9561 VSS.t581 37.2185
R452 VSS.n1183 VSS.t676 37.2185
R453 VSS.n565 VSS.t1069 37.2185
R454 VSS.t800 VSS.n11288 37.2185
R455 VSS.n11298 VSS.t839 37.2185
R456 VSS.t98 VSS.t596 36.3418
R457 VSS.t104 VSS.t500 36.3418
R458 VSS.t1162 VSS.t472 35.4652
R459 VSS.t643 VSS.t207 35.1464
R460 VSS.n1390 VSS.t413 34.7479
R461 VSS.t259 VSS.t692 34.5885
R462 VSS.t254 VSS.t1162 34.5885
R463 VSS.t257 VSS.t643 34.5088
R464 VSS.t325 VSS.t477 34.2697
R465 VSS.n9465 VSS.t1437 33.8803
R466 VSS.n4805 VSS.n4804 33.7899
R467 VSS.t500 VSS.t54 33.3134
R468 VSS.t314 VSS.n833 32.0383
R469 VSS.t148 VSS.n6 32.0383
R470 VSS.n10118 VSS.t411 31.2413
R471 VSS.n10067 VSS.t327 31.2413
R472 VSS.n11152 VSS.t171 31.2413
R473 VSS.t533 VSS.n1390 30.7631
R474 VSS.t253 VSS.t329 30.4443
R475 VSS.t410 VSS.t209 30.3646
R476 VSS.t472 VSS.t328 30.0459
R477 VSS.t181 VSS.t735 29.5677
R478 VSS.n10599 VSS.n10442 29.446
R479 VSS.t177 VSS.t98 29.1692
R480 VSS.n1499 VSS.n1498 28.5785
R481 VSS.t316 VSS.t251 28.2926
R482 VSS.t412 VSS.t252 27.9738
R483 VSS.n10602 VSS.n10601 26.8369
R484 VSS.t154 VSS.t2481 26.7681
R485 VSS.t149 VSS.t97 26.6986
R486 VSS.n11299 VSS.n11298 26.4596
R487 VSS.n9889 VSS.t330 25.9017
R488 VSS.t312 VSS.t606 25.5032
R489 VSS.n9526 VSS.n9525 25.1844
R490 VSS.t1069 VSS.t95 25.025
R491 VSS.t536 VSS.t99 25.025
R492 VSS.t301 VSS.t658 23.2767
R493 VSS.n9766 VSS.t223 23.1123
R494 VSS.n11279 VSS.t52 23.1123
R495 VSS.t738 VSS.t66 22.5544
R496 VSS.t145 VSS.n11297 22.4748
R497 VSS.t160 VSS.n208 22.2357
R498 VSS.n11297 VSS.t146 22.156
R499 VSS.t66 VSS.t573 22.0763
R500 VSS.n9302 VSS.t335 21.8797
R501 VSS.t209 VSS.n10117 21.5184
R502 VSS.t214 VSS.n10066 21.5184
R503 VSS.n10032 VSS.t63 21.5184
R504 VSS.n11292 VSS.t61 21.5184
R505 VSS.n10929 VSS.n217 21.2793
R506 VSS.t1242 VSS.t155 21.0784
R507 VSS.t514 VSS.t187 20.8733
R508 VSS.t13 VSS.t530 20.8733
R509 VSS.t590 VSS.n506 20.6417
R510 VSS.t260 VSS.t873 20.4824
R511 VSS.t95 VSS.t536 19.6057
R512 VSS.t283 VSS.t718 19.2072
R513 VSS.t606 VSS.t314 19.1275
R514 VSS.n1184 VSS.t218 18.8884
R515 VSS.n1394 VSS.n1393 18.6214
R516 VSS.n9013 VSS.n9010 18.4538
R517 VSS.n9092 VSS.n9091 18.4538
R518 VSS.n9114 VSS.n9113 18.4538
R519 VSS.n9180 VSS.n9177 18.4475
R520 VSS.n9249 VSS.n9248 18.4475
R521 VSS.n9307 VSS.n9299 18.4475
R522 VSS.t503 VSS.t214 18.3306
R523 VSS.t218 VSS.t542 18.3306
R524 VSS.n352 VSS.n351 18.2692
R525 VSS.n10185 VSS.n10184 18.2692
R526 VSS.n10178 VSS.n392 18.2692
R527 VSS.n280 VSS.n279 18.263
R528 VSS.n10245 VSS.n10244 18.263
R529 VSS.n10238 VSS.n320 18.263
R530 VSS.t159 VSS.t0 18.0778
R531 VSS.t182 VSS.t40 18.0778
R532 VSS.t191 VSS.t134 18.0778
R533 VSS.t103 VSS.t149 17.9321
R534 VSS.t97 VSS.t148 17.9321
R535 VSS.n566 VSS.t58 17.7727
R536 VSS.n9561 VSS.n9560 17.6133
R537 VSS.n11279 VSS.n148 17.6133
R538 VSS.n9525 VSS.t260 16.7366
R539 VSS.n11286 VSS.n93 16.7366
R540 VSS.n11361 VSS.t721 16.5773
R541 VSS.t256 VSS.t316 16.3382
R542 VSS.t251 VSS.t313 16.3382
R543 VSS.t35 VSS.t163 16.2142
R544 VSS.t22 VSS.t166 16.2142
R545 VSS.t15 VSS.t183 16.2142
R546 VSS.n11468 VSS.t486 16.0991
R547 VSS.n9301 VSS.n9300 15.6285
R548 VSS.n10125 VSS.n10124 15.6285
R549 VSS.t324 VSS.t721 15.4615
R550 VSS.n11287 VSS.t61 15.1427
R551 VSS.t146 VSS.t486 15.1427
R552 VSS.t735 VSS.t160 15.063
R553 VSS.n9564 VSS.t256 14.9036
R554 VSS.n4803 VSS.n1580 14.678
R555 VSS.n8954 VSS.n8953 14.6753
R556 VSS.t1258 VSS.t100 14.6646
R557 VSS.t327 VSS.t253 14.1864
R558 VSS.t329 VSS.t258 14.1864
R559 VSS.t52 VSS.t686 14.1067
R560 VSS.n10117 VSS.t655 13.6285
R561 VSS.t1621 VSS.t33 13.4187
R562 VSS.t162 VSS.t704 13.4187
R563 VSS.t211 VSS.t620 12.194
R564 VSS.t581 VSS.t223 12.194
R565 VSS.t718 VSS.n218 12.0346
R566 VSS.n9523 VSS.t312 11.7955
R567 VSS.n9524 VSS.n9523 11.4767
R568 VSS.n9890 VSS.n9889 11.4767
R569 VSS.n1184 VSS.n1183 11.4767
R570 VSS.n11289 VSS.n11286 11.4767
R571 VSS.n11288 VSS.n11287 11.4767
R572 VSS.t330 VSS.t590 11.397
R573 VSS.t913 VSS.t96 10.9188
R574 VSS.t281 VSS.n217 10.7595
R575 VSS.n8952 VSS.n1580 10.4817
R576 VSS.t63 VSS.t563 10.361
R577 VSS.t477 VSS.t326 10.361
R578 VSS.t692 VSS.t254 10.0422
R579 VSS.t94 VSS.t323 9.96249
R580 VSS.n10982 VSS.n208 9.8031
R581 VSS.t207 VSS.t655 9.48432
R582 VSS.n1353 VSS.t262 9.37419
R583 VSS.n9766 VSS.t620 9.32492
R584 VSS.n9143 VSS.n9142 9.30555
R585 VSS.n1491 VSS.n1490 9.30555
R586 VSS.n1211 VSS.n1210 9.30555
R587 VSS.n10949 VSS.n10948 9.30555
R588 VSS.n10995 VSS.n10994 9.30555
R589 VSS.n8976 VSS.n8975 9.30555
R590 VSS.n981 VSS.n980 9.30555
R591 VSS.n1039 VSS.n1038 9.30555
R592 VSS.n1088 VSS.n1087 9.30555
R593 VSS.n874 VSS.n873 9.30555
R594 VSS.n576 VSS.t102 9.29148
R595 VSS.n9304 VSS.t386 9.05234
R596 VSS.n1392 VSS.n1391 9.05234
R597 VSS.n9303 VSS.t387 8.92303
R598 VSS.n11309 VSS.n128 8.8165
R599 VSS.n10837 VSS.t3119 8.52542
R600 VSS.n10791 VSS.t3543 8.52542
R601 VSS.n10809 VSS.t846 8.52542
R602 VSS.n10828 VSS.t2775 8.52542
R603 VSS.n10773 VSS.t1467 8.52542
R604 VSS.n10855 VSS.t1899 8.52542
R605 VSS.n10742 VSS.t2296 8.52542
R606 VSS.n10746 VSS.t1081 8.52542
R607 VSS.n10813 VSS.t3209 8.52542
R608 VSS.n10815 VSS.t1913 8.52542
R609 VSS.n10749 VSS.t893 8.52542
R610 VSS.n10747 VSS.t585 8.52542
R611 VSS.n10736 VSS.t3549 8.52542
R612 VSS.n10784 VSS.t2238 8.52542
R613 VSS.n10737 VSS.t1267 8.52542
R614 VSS.n10778 VSS.t966 8.52542
R615 VSS.t489 VSS.t1227 8.40578
R616 VSS.t596 VSS.t104 8.28888
R617 VSS.n4803 VSS.n60 8.20625
R618 VSS.n9202 VSS.t631 8.06917
R619 VSS.n9184 VSS.t2731 8.06917
R620 VSS.n9058 VSS.t3309 8.06917
R621 VSS.n9057 VSS.t2280 8.06917
R622 VSS.n9054 VSS.t2901 8.06917
R623 VSS.n9054 VSS.t3583 8.06917
R624 VSS.n9051 VSS.t2080 8.06917
R625 VSS.n9051 VSS.t2811 8.06917
R626 VSS.n9050 VSS.t2392 8.06917
R627 VSS.n9050 VSS.t3135 8.06917
R628 VSS.n9122 VSS.t1229 8.06917
R629 VSS.n9122 VSS.t1943 8.06917
R630 VSS.n9123 VSS.t776 8.06917
R631 VSS.n9123 VSS.t1542 8.06917
R632 VSS.n9127 VSS.t2198 8.06917
R633 VSS.n9127 VSS.t2905 8.06917
R634 VSS.n9054 VSS.t1789 8.06917
R635 VSS.n9054 VSS.t1631 8.06917
R636 VSS.n9051 VSS.t941 8.06917
R637 VSS.n9051 VSS.t761 8.06917
R638 VSS.n9050 VSS.t1296 8.06917
R639 VSS.n9050 VSS.t1100 8.06917
R640 VSS.n9122 VSS.t3191 8.06917
R641 VSS.n9122 VSS.t3045 8.06917
R642 VSS.n9123 VSS.t2805 8.06917
R643 VSS.n9123 VSS.t2613 8.06917
R644 VSS.n9127 VSS.t1046 8.06917
R645 VSS.n9127 VSS.t870 8.06917
R646 VSS.n1543 VSS.t3515 8.06917
R647 VSS.n1542 VSS.t1516 8.06917
R648 VSS.n1549 VSS.t1779 8.06917
R649 VSS.n1541 VSS.t1019 8.06917
R650 VSS.n9171 VSS.t3107 8.06917
R651 VSS.n9137 VSS.t2021 8.06917
R652 VSS.n1526 VSS.t2639 8.06917
R653 VSS.n9133 VSS.t1610 8.06917
R654 VSS.n1512 VSS.t866 8.06917
R655 VSS.n9253 VSS.t2947 8.06917
R656 VSS.n9139 VSS.t1717 8.06917
R657 VSS.n9138 VSS.t2402 8.06917
R658 VSS.n9237 VSS.t2935 8.06917
R659 VSS.n9237 VSS.t1875 8.06917
R660 VSS.n9234 VSS.t2128 8.06917
R661 VSS.n9234 VSS.t1038 8.06917
R662 VSS.n9233 VSS.t2434 8.06917
R663 VSS.n9233 VSS.t1415 8.06917
R664 VSS.n9227 VSS.t1263 8.06917
R665 VSS.n9227 VSS.t3275 8.06917
R666 VSS.n9226 VSS.t818 8.06917
R667 VSS.n9226 VSS.t2897 8.06917
R668 VSS.n9223 VSS.t2218 8.06917
R669 VSS.n9223 VSS.t1151 8.06917
R670 VSS.n9237 VSS.t3339 8.06917
R671 VSS.n9237 VSS.t1372 8.06917
R672 VSS.n9234 VSS.t2569 8.06917
R673 VSS.n9234 VSS.t3635 8.06917
R674 VSS.n9233 VSS.t2913 8.06917
R675 VSS.n9233 VSS.t836 8.06917
R676 VSS.n9227 VSS.t1725 8.06917
R677 VSS.n9227 VSS.t2781 8.06917
R678 VSS.n9226 VSS.t1319 8.06917
R679 VSS.n9226 VSS.t2352 8.06917
R680 VSS.n9223 VSS.t2681 8.06917
R681 VSS.n9223 VSS.t575 8.06917
R682 VSS.n9242 VSS.t1623 8.06917
R683 VSS.n9212 VSS.t3625 8.06917
R684 VSS.n1518 VSS.t2390 8.06917
R685 VSS.n9208 VSS.t3131 8.06917
R686 VSS.n1504 VSS.t2046 8.06917
R687 VSS.n9311 VSS.t972 8.06917
R688 VSS.n9214 VSS.t1635 8.06917
R689 VSS.n9213 VSS.t2318 8.06917
R690 VSS.n9269 VSS.t2567 8.06917
R691 VSS.n9269 VSS.t1540 8.06917
R692 VSS.n9273 VSS.t1797 8.06917
R693 VSS.n9273 VSS.t672 8.06917
R694 VSS.n9274 VSS.t2106 8.06917
R695 VSS.n9274 VSS.t1009 8.06917
R696 VSS.n9282 VSS.t888 8.06917
R697 VSS.n9282 VSS.t2959 8.06917
R698 VSS.n9283 VSS.t3581 8.06917
R699 VSS.n9283 VSS.t2531 8.06917
R700 VSS.n9287 VSS.t1883 8.06917
R701 VSS.n9287 VSS.t784 8.06917
R702 VSS.n9269 VSS.t2803 8.06917
R703 VSS.n9269 VSS.t725 8.06917
R704 VSS.n9273 VSS.t1991 8.06917
R705 VSS.n9273 VSS.t3069 8.06917
R706 VSS.n9274 VSS.t2298 8.06917
R707 VSS.n9274 VSS.t3327 8.06917
R708 VSS.n9282 VSS.t1096 8.06917
R709 VSS.n9282 VSS.t2194 8.06917
R710 VSS.n9283 VSS.t651 8.06917
R711 VSS.n9283 VSS.t1791 8.06917
R712 VSS.n9287 VSS.t2074 8.06917
R713 VSS.n9287 VSS.t3149 8.06917
R714 VSS.n9293 VSS.t1374 8.06917
R715 VSS.n9263 VSS.t3349 8.06917
R716 VSS.n1508 VSS.t884 8.06917
R717 VSS.n9259 VSS.t1639 8.06917
R718 VSS.n1495 VSS.t2857 8.06917
R719 VSS.n9351 VSS.t2142 8.06917
R720 VSS.n9265 VSS.t1382 8.06917
R721 VSS.n9264 VSS.t2406 8.06917
R722 VSS.n9372 VSS.t3459 8.06917
R723 VSS.n9372 VSS.t2779 8.06917
R724 VSS.n9369 VSS.t2685 8.06917
R725 VSS.n9369 VSS.t1975 8.06917
R726 VSS.n9368 VSS.t3021 8.06917
R727 VSS.n9368 VSS.t2282 8.06917
R728 VSS.n9362 VSS.t1829 8.06917
R729 VSS.n9362 VSS.t1088 8.06917
R730 VSS.n9361 VSS.t1436 8.06917
R731 VSS.n9361 VSS.t637 8.06917
R732 VSS.n9358 VSS.t2787 8.06917
R733 VSS.n9358 VSS.t2064 8.06917
R734 VSS.n9372 VSS.t1182 8.06917
R735 VSS.n9372 VSS.t2252 8.06917
R736 VSS.n9369 VSS.t3463 8.06917
R737 VSS.n9369 VSS.t1486 8.06917
R738 VSS.n9368 VSS.t657 8.06917
R739 VSS.n9368 VSS.t1793 8.06917
R740 VSS.n9362 VSS.t2609 8.06917
R741 VSS.n9362 VSS.t479 8.06917
R742 VSS.n9361 VSS.t2214 8.06917
R743 VSS.n9361 VSS.t3255 8.06917
R744 VSS.n9358 VSS.t3567 8.06917
R745 VSS.n9358 VSS.t1573 8.06917
R746 VSS.n9340 VSS.t3539 8.06917
R747 VSS.n9321 VSS.t2853 8.06917
R748 VSS.n1500 VSS.t2054 8.06917
R749 VSS.n9317 VSS.t3137 8.06917
R750 VSS.n1476 VSS.t2603 8.06917
R751 VSS.n9384 VSS.t474 8.06917
R752 VSS.n1477 VSS.t2186 8.06917
R753 VSS.n9377 VSS.t3219 8.06917
R754 VSS.n9392 VSS.t2695 8.06917
R755 VSS.n9392 VSS.t592 8.06917
R756 VSS.n9396 VSS.t1889 8.06917
R757 VSS.n9396 VSS.t2957 8.06917
R758 VSS.n9397 VSS.t2212 8.06917
R759 VSS.n9397 VSS.t3251 8.06917
R760 VSS.n9405 VSS.t988 8.06917
R761 VSS.n9405 VSS.t2070 8.06917
R762 VSS.n9406 VSS.t532 8.06917
R763 VSS.n9406 VSS.t1691 8.06917
R764 VSS.n9410 VSS.t1983 8.06917
R765 VSS.n9410 VSS.t3065 8.06917
R766 VSS.n9392 VSS.t2017 8.06917
R767 VSS.n9392 VSS.t1330 8.06917
R768 VSS.n9396 VSS.t1226 8.06917
R769 VSS.n9396 VSS.t3589 8.06917
R770 VSS.n9397 VSS.t1567 8.06917
R771 VSS.n9397 VSS.t804 8.06917
R772 VSS.n9405 VSS.t3413 8.06917
R773 VSS.n9405 VSS.t2735 8.06917
R774 VSS.n9406 VSS.t3057 8.06917
R775 VSS.n9406 VSS.t2322 8.06917
R776 VSS.n9410 VSS.t1334 8.06917
R777 VSS.n9410 VSS.t526 8.06917
R778 VSS.n9416 VSS.t1915 8.06917
R779 VSS.n1397 VSS.t2987 8.06917
R780 VSS.n1487 VSS.t1494 8.06917
R781 VSS.n1486 VSS.t2517 8.06917
R782 VSS.n1220 VSS.t1094 8.06917
R783 VSS.n9531 VSS.t2184 8.06917
R784 VSS.n1399 VSS.t1421 8.06917
R785 VSS.n1398 VSS.t625 8.06917
R786 VSS.n1435 VSS.t1557 8.06917
R787 VSS.n1435 VSS.t2583 8.06917
R788 VSS.n1434 VSS.t1871 8.06917
R789 VSS.n1434 VSS.t2943 8.06917
R790 VSS.n1229 VSS.t613 8.06917
R791 VSS.n1229 VSS.t1755 8.06917
R792 VSS.n1228 VSS.t3319 8.06917
R793 VSS.n1228 VSS.t1340 8.06917
R794 VSS.n1225 VSS.t1659 8.06917
R795 VSS.n1225 VSS.t2715 8.06917
R796 VSS.n1435 VSS.t3507 8.06917
R797 VSS.n1435 VSS.t2823 8.06917
R798 VSS.n1434 VSS.t713 8.06917
R799 VSS.n1434 VSS.t3141 8.06917
R800 VSS.n1229 VSS.t2649 8.06917
R801 VSS.n1229 VSS.t1947 8.06917
R802 VSS.n1228 VSS.t2240 8.06917
R803 VSS.n1228 VSS.t1547 8.06917
R804 VSS.n1225 VSS.t3599 8.06917
R805 VSS.n1225 VSS.t2915 8.06917
R806 VSS.n11235 VSS.t3207 8.06917
R807 VSS.n11233 VSS.t806 8.06917
R808 VSS.n11229 VSS.t1461 8.06917
R809 VSS.n11224 VSS.t3443 8.06917
R810 VSS.n11202 VSS.t1903 8.06917
R811 VSS.n11200 VSS.t2969 8.06917
R812 VSS.n11257 VSS.t3195 8.06917
R813 VSS.n11196 VSS.t2154 8.06917
R814 VSS.n11181 VSS.t2769 8.06917
R815 VSS.n11179 VSS.t3453 8.06917
R816 VSS.n11175 VSS.t3313 8.06917
R817 VSS.n11173 VSS.t944 8.06917
R818 VSS.n153 VSS.t3053 8.06917
R819 VSS.n11164 VSS.t595 8.06917
R820 VSS.n177 VSS.t2294 8.06917
R821 VSS.n11156 VSS.t1255 8.06917
R822 VSS.n735 VSS.t1873 8.06917
R823 VSS.n731 VSS.t772 8.06917
R824 VSS.n729 VSS.t2110 8.06917
R825 VSS.n746 VSS.t3163 8.06917
R826 VSS.n705 VSS.t1357 8.06917
R827 VSS.n703 VSS.t2039 8.06917
R828 VSS.n699 VSS.t3601 8.06917
R829 VSS.n695 VSS.t1612 8.06917
R830 VSS.n692 VSS.t1867 8.06917
R831 VSS.n9835 VSS.t1128 8.06917
R832 VSS.n9830 VSS.t520 8.06917
R833 VSS.n9824 VSS.t1685 8.06917
R834 VSS.n9818 VSS.t2138 8.06917
R835 VSS.n9811 VSS.t1058 8.06917
R836 VSS.n9807 VSS.t2364 8.06917
R837 VSS.n9801 VSS.t3387 8.06917
R838 VSS.n9797 VSS.t3023 8.06917
R839 VSS.n788 VSS.t1949 8.06917
R840 VSS.n789 VSS.t3231 8.06917
R841 VSS.n9784 VSS.t1214 8.06917
R842 VSS.n9775 VSS.t2727 8.06917
R843 VSS.n9769 VSS.t2007 8.06917
R844 VSS.n9587 VSS.t2266 8.06917
R845 VSS.n9567 VSS.t1508 8.06917
R846 VSS.n830 VSS.t1775 8.06917
R847 VSS.n9600 VSS.t1011 8.06917
R848 VSS.n1442 VSS.t2328 8.06917
R849 VSS.n1440 VSS.t3363 8.06917
R850 VSS.n1453 VSS.t1231 8.06917
R851 VSS.n1455 VSS.t3593 8.06917
R852 VSS.n1424 VSS.t1818 8.06917
R853 VSS.n1467 VSS.t2885 8.06917
R854 VSS.n1471 VSS.t2096 8.06917
R855 VSS.n1417 VSS.t1417 8.06917
R856 VSS.n1154 VSS.t2426 8.06917
R857 VSS.n1154 VSS.t3489 8.06917
R858 VSS.n1155 VSS.t2767 8.06917
R859 VSS.n1155 VSS.t691 8.06917
R860 VSS.n9555 VSS.t1602 8.06917
R861 VSS.n9555 VSS.t2627 8.06917
R862 VSS.n9554 VSS.t1161 8.06917
R863 VSS.n9554 VSS.t2224 8.06917
R864 VSS.n9551 VSS.t2535 8.06917
R865 VSS.n9551 VSS.t3585 8.06917
R866 VSS.n1154 VSS.t1935 8.06917
R867 VSS.n1154 VSS.t1218 8.06917
R868 VSS.n1155 VSS.t2242 8.06917
R869 VSS.n1155 VSS.t1551 8.06917
R870 VSS.n9555 VSS.t1036 8.06917
R871 VSS.n9555 VSS.t3401 8.06917
R872 VSS.n9554 VSS.t580 8.06917
R873 VSS.n9554 VSS.t3049 8.06917
R874 VSS.n9551 VSS.t2015 8.06917
R875 VSS.n9551 VSS.t1326 8.06917
R876 VSS.n1215 VSS.t1577 8.06917
R877 VSS.n9544 VSS.t742 8.06917
R878 VSS.n1216 VSS.t1021 8.06917
R879 VSS.n9537 VSS.t3391 8.06917
R880 VSS.n1201 VSS.t1687 8.06917
R881 VSS.n1163 VSS.t2733 8.06917
R882 VSS.n1207 VSS.t2292 8.06917
R883 VSS.n1162 VSS.t1251 8.06917
R884 VSS.n213 VSS.t2933 8.06917
R885 VSS.n10933 VSS.t851 8.06917
R886 VSS.n1165 VSS.t1139 8.06917
R887 VSS.n1164 VSS.t3531 8.06917
R888 VSS.n10976 VSS.t1627 8.06917
R889 VSS.n10943 VSS.t3629 8.06917
R890 VSS.n209 VSS.t1149 8.06917
R891 VSS.n10939 VSS.t3183 8.06917
R892 VSS.n89 VSS.t2478 8.06917
R893 VSS.n11365 VSS.t1469 8.06917
R894 VSS.n10945 VSS.t2056 8.06917
R895 VSS.n10944 VSS.t2783 8.06917
R896 VSS.n84 VSS.t2973 8.06917
R897 VSS.n11378 VSS.t1907 8.06917
R898 VSS.n85 VSS.t2499 8.06917
R899 VSS.n11371 VSS.t3215 8.06917
R900 VSS.n66 VSS.t2330 8.06917
R901 VSS.n66 VSS.t3365 8.06917
R902 VSS.n67 VSS.t2663 8.06917
R903 VSS.n67 VSS.t560 8.06917
R904 VSS.n73 VSS.t1504 8.06917
R905 VSS.n73 VSS.t2529 8.06917
R906 VSS.n74 VSS.t1044 8.06917
R907 VSS.n74 VSS.t2134 8.06917
R908 VSS.n77 VSS.t2422 8.06917
R909 VSS.n77 VSS.t3481 8.06917
R910 VSS.t3239 VSS.n11458 8.06917
R911 VSS.n11459 VSS.t3239 8.06917
R912 VSS.t2456 VSS.n11456 8.06917
R913 VSS.n11457 VSS.t2456 8.06917
R914 VSS.t2595 VSS.n11454 8.06917
R915 VSS.n11455 VSS.t2595 8.06917
R916 VSS.t1833 VSS.n11452 8.06917
R917 VSS.n11453 VSS.t1833 8.06917
R918 VSS.n23 VSS.t998 8.06917
R919 VSS.t998 VSS.n18 8.06917
R920 VSS.t1157 VSS.n11442 8.06917
R921 VSS.n11443 VSS.t1157 8.06917
R922 VSS.t3441 VSS.n11440 8.06917
R923 VSS.n11441 VSS.t3441 8.06917
R924 VSS.t2699 VSS.n11438 8.06917
R925 VSS.n11439 VSS.t2699 8.06917
R926 VSS.t2991 VSS.n11436 8.06917
R927 VSS.n11437 VSS.t2991 8.06917
R928 VSS.t919 VSS.n11434 8.06917
R929 VSS.n11435 VSS.t919 8.06917
R930 VSS.t1545 VSS.n11427 8.06917
R931 VSS.n11428 VSS.t1545 8.06917
R932 VSS.t2525 VSS.n11425 8.06917
R933 VSS.n11426 VSS.t2525 8.06917
R934 VSS.t1769 VSS.n11423 8.06917
R935 VSS.n11424 VSS.t1769 8.06917
R936 VSS.t927 VSS.n11421 8.06917
R937 VSS.n11422 VSS.t927 8.06917
R938 VSS.t1077 VSS.n11419 8.06917
R939 VSS.n11420 VSS.t1077 8.06917
R940 VSS.n48 VSS.t3361 8.06917
R941 VSS.t3361 VSS.n43 8.06917
R942 VSS.t2771 VSS.n11409 8.06917
R943 VSS.n11410 VSS.t2771 8.06917
R944 VSS.t1985 VSS.n11407 8.06917
R945 VSS.n11408 VSS.t1985 8.06917
R946 VSS.t1405 VSS.n11405 8.06917
R947 VSS.n11406 VSS.t1405 8.06917
R948 VSS.t485 VSS.n11403 8.06917
R949 VSS.n11404 VSS.t485 8.06917
R950 VSS.t1695 VSS.n11401 8.06917
R951 VSS.n11402 VSS.t1695 8.06917
R952 VSS.n63 VSS.t3147 8.06917
R953 VSS.n63 VSS.t1090 8.06917
R954 VSS.n63 VSS.t466 8.06917
R955 VSS.n63 VSS.t2585 8.06917
R956 VSS.n11324 VSS.t2216 8.06917
R957 VSS.n118 VSS.t1979 8.06917
R958 VSS.n11462 VSS.t1465 8.06917
R959 VSS.n11 VSS.t1498 8.06917
R960 VSS.n11091 VSS.t1719 8.06917
R961 VSS.n11089 VSS.t629 8.06917
R962 VSS.n11084 VSS.t2891 8.06917
R963 VSS.n11079 VSS.t2919 8.06917
R964 VSS.n11058 VSS.t1324 8.06917
R965 VSS.n11056 VSS.t1048 8.06917
R966 VSS.n11113 VSS.t2462 8.06917
R967 VSS.n11052 VSS.t2487 8.06917
R968 VSS.n11034 VSS.t2745 8.06917
R969 VSS.n11032 VSS.t1751 8.06917
R970 VSS.n11028 VSS.t2673 8.06917
R971 VSS.n11025 VSS.t1677 8.06917
R972 VSS.n11132 VSS.t2308 8.06917
R973 VSS.n203 VSS.t1303 8.06917
R974 VSS.n11145 VSS.t1188 8.06917
R975 VSS.n186 VSS.t1239 8.06917
R976 VSS.n10880 VSS.t1490 8.06917
R977 VSS.n10885 VSS.t1518 8.06917
R978 VSS.n10889 VSS.t535 8.06917
R979 VSS.n10873 VSS.t3435 8.06917
R980 VSS.n237 VSS.t1403 8.06917
R981 VSS.n557 VSS.t3411 8.06917
R982 VSS.n553 VSS.t2827 8.06917
R983 VSS.n549 VSS.t2561 8.06917
R984 VSS.n10049 VSS.t2025 8.06917
R985 VSS.n544 VSS.t2855 8.06917
R986 VSS.n540 VSS.t2300 8.06917
R987 VSS.n538 VSS.t2062 8.06917
R988 VSS.n514 VSS.t2759 8.06917
R989 VSS.n529 VSS.t2807 8.06917
R990 VSS.n523 VSS.t1921 8.06917
R991 VSS.n518 VSS.t1689 8.06917
R992 VSS.n500 VSS.t1084 8.06917
R993 VSS.n498 VSS.t1113 8.06917
R994 VSS.n495 VSS.t3307 8.06917
R995 VSS.n10080 VSS.t3117 8.06917
R996 VSS.n489 VSS.t3403 8.06917
R997 VSS.n486 VSS.t1147 8.06917
R998 VSS.n478 VSS.t2553 8.06917
R999 VSS.n459 VSS.t2677 8.06917
R1000 VSS.n10098 VSS.t2140 8.06917
R1001 VSS.n456 VSS.t2955 8.06917
R1002 VSS.n452 VSS.t2052 8.06917
R1003 VSS.n450 VSS.t1835 8.06917
R1004 VSS.n10111 VSS.t2037 8.06917
R1005 VSS.n442 VSS.t2869 8.06917
R1006 VSS.n1301 VSS.t1977 8.06917
R1007 VSS.n1308 VSS.t1753 8.06917
R1008 VSS.n1297 VSS.t3461 8.06917
R1009 VSS.n1317 VSS.t1190 8.06917
R1010 VSS.n11335 VSS.t3165 8.06917
R1011 VSS.n11335 VSS.t2941 8.06917
R1012 VSS.n11333 VSS.t838 8.06917
R1013 VSS.n11333 VSS.t557 8.06917
R1014 VSS.n11332 VSS.t1294 8.06917
R1015 VSS.n11332 VSS.t1023 8.06917
R1016 VSS.n11328 VSS.t1757 8.06917
R1017 VSS.n11328 VSS.t1520 8.06917
R1018 VSS.n11327 VSS.t3573 8.06917
R1019 VSS.n11327 VSS.t3305 8.06917
R1020 VSS.n11342 VSS.t2376 8.06917
R1021 VSS.n102 VSS.t2408 8.06917
R1022 VSS.n11349 VSS.t2655 8.06917
R1023 VSS.n101 VSS.t1663 8.06917
R1024 VSS.n11355 VSS.t3383 8.06917
R1025 VSS.n97 VSS.t3425 8.06917
R1026 VSS.n10991 VSS.t518 8.06917
R1027 VSS.n10990 VSS.t2683 8.06917
R1028 VSS.n206 VSS.t2152 8.06917
R1029 VSS.n10986 VSS.t2188 8.06917
R1030 VSS.n10917 VSS.t2396 8.06917
R1031 VSS.n10916 VSS.t2428 8.06917
R1032 VSS.n10635 VSS.t3637 8.06917
R1033 VSS.n10635 VSS.t1376 8.06917
R1034 VSS.n10635 VSS.t1108 8.06917
R1035 VSS.n10635 VSS.t3491 8.06917
R1036 VSS.n10352 VSS.t1981 8.06917
R1037 VSS.n10640 VSS.t2404 8.06917
R1038 VSS.n10351 VSS.t790 8.06917
R1039 VSS.n10645 VSS.t2587 8.06917
R1040 VSS.n10350 VSS.t1653 8.06917
R1041 VSS.n10650 VSS.t2398 8.06917
R1042 VSS.n10346 VSS.t529 8.06917
R1043 VSS.n10516 VSS.t660 8.06917
R1044 VSS.n10508 VSS.t2849 8.06917
R1045 VSS.n10506 VSS.t2929 8.06917
R1046 VSS.n10502 VSS.t2288 8.06917
R1047 VSS.n10532 VSS.t1032 8.06917
R1048 VSS.n10491 VSS.t3175 8.06917
R1049 VSS.n10543 VSS.t3595 8.06917
R1050 VSS.n10487 VSS.t2631 8.06917
R1051 VSS.n10485 VSS.t1693 8.06917
R1052 VSS.n10590 VSS.t2841 8.06917
R1053 VSS.n10348 VSS.t1073 8.06917
R1054 VSS.n10510 VSS.t1170 8.06917
R1055 VSS.n10517 VSS.t877 8.06917
R1056 VSS.n10507 VSS.t570 8.06917
R1057 VSS.n10505 VSS.t2755 8.06917
R1058 VSS.n10500 VSS.t1897 8.06917
R1059 VSS.n10490 VSS.t703 8.06917
R1060 VSS.n10544 VSS.t1893 8.06917
R1061 VSS.n10486 VSS.t891 8.06917
R1062 VSS.n10484 VSS.t3061 8.06917
R1063 VSS.n10591 VSS.t1145 8.06917
R1064 VSS.n10496 VSS.t3125 8.06917
R1065 VSS.n10495 VSS.t786 8.06917
R1066 VSS.n10606 VSS.t513 8.06917
R1067 VSS.n10607 VSS.t2993 8.06917
R1068 VSS.n10609 VSS.t1476 8.06917
R1069 VSS.n10496 VSS.t1967 8.06917
R1070 VSS.n10495 VSS.t2757 8.06917
R1071 VSS.n10606 VSS.t2539 8.06917
R1072 VSS.n10607 VSS.t1839 8.06917
R1073 VSS.n10609 VSS.t3351 8.06917
R1074 VSS.n10412 VSS.t1474 8.06917
R1075 VSS.n10435 VSS.t3559 8.06917
R1076 VSS.n10413 VSS.t2581 8.06917
R1077 VSS.n10414 VSS.t662 8.06917
R1078 VSS.n10427 VSS.t2851 8.06917
R1079 VSS.n10415 VSS.t2931 8.06917
R1080 VSS.n10416 VSS.t2290 8.06917
R1081 VSS.n10420 VSS.t2372 8.06917
R1082 VSS.n10417 VSS.t1439 8.06917
R1083 VSS.n10477 VSS.t3249 8.06917
R1084 VSS.n10479 VSS.t3081 8.06917
R1085 VSS.n10480 VSS.t1701 8.06917
R1086 VSS.n10595 VSS.t2911 8.06917
R1087 VSS.n10594 VSS.t1620 8.06917
R1088 VSS.n10448 VSS.t1143 8.06917
R1089 VSS.n10457 VSS.t3261 8.06917
R1090 VSS.n10447 VSS.t3315 8.06917
R1091 VSS.n10446 VSS.t2737 8.06917
R1092 VSS.n10465 VSS.t1524 8.06917
R1093 VSS.n10445 VSS.t3605 8.06917
R1094 VSS.n10444 VSS.t925 8.06917
R1095 VSS.n10472 VSS.t3105 8.06917
R1096 VSS.n10443 VSS.t2118 8.06917
R1097 VSS.n10452 VSS.t1025 8.06917
R1098 VSS.n10450 VSS.t808 8.06917
R1099 VSS.n10449 VSS.t2545 8.06917
R1100 VSS.n10658 VSS.t627 8.06917
R1101 VSS.n10657 VSS.t2458 8.06917
R1102 VSS.n10585 VSS.t3263 8.06917
R1103 VSS.n10553 VSS.t3317 8.06917
R1104 VSS.n10554 VSS.t2739 8.06917
R1105 VSS.n10578 VSS.t2837 8.06917
R1106 VSS.n10555 VSS.t1859 8.06917
R1107 VSS.n10561 VSS.t1961 8.06917
R1108 VSS.n10559 VSS.t3179 8.06917
R1109 VSS.n10558 VSS.t855 8.06917
R1110 VSS.n10692 VSS.t600 8.06917
R1111 VSS.n10691 VSS.t3067 8.06917
R1112 VSS.n10689 VSS.t1536 8.06917
R1113 VSS.n1573 VSS.t1709 8.06917
R1114 VSS.n1573 VSS.t2751 8.06917
R1115 VSS.n1576 VSS.t860 8.06917
R1116 VSS.n1576 VSS.t1955 8.06917
R1117 VSS.n1577 VSS.t1220 8.06917
R1118 VSS.n1577 VSS.t2274 8.06917
R1119 VSS.n8958 VSS.t3127 8.06917
R1120 VSS.n8958 VSS.t1066 8.06917
R1121 VSS.n8959 VSS.t2719 8.06917
R1122 VSS.n8959 VSS.t616 8.06917
R1123 VSS.n8962 VSS.t962 8.06917
R1124 VSS.n8962 VSS.t2044 8.06917
R1125 VSS.n9035 VSS.t2879 8.06917
R1126 VSS.n9017 VSS.t802 8.06917
R1127 VSS.n1567 VSS.t1086 8.06917
R1128 VSS.n1566 VSS.t3469 8.06917
R1129 VSS.n8980 VSS.t2579 8.06917
R1130 VSS.n8980 VSS.t1820 8.06917
R1131 VSS.n8984 VSS.t1810 8.06917
R1132 VSS.n8984 VSS.t980 8.06917
R1133 VSS.n8985 VSS.t2122 8.06917
R1134 VSS.n8985 VSS.t1355 8.06917
R1135 VSS.n8993 VSS.t900 8.06917
R1136 VSS.n8993 VSS.t3229 8.06917
R1137 VSS.n8994 VSS.t3597 8.06917
R1138 VSS.n8994 VSS.t2847 8.06917
R1139 VSS.n8998 VSS.t1901 8.06917
R1140 VSS.n8998 VSS.t1092 8.06917
R1141 VSS.n8980 VSS.t3297 8.06917
R1142 VSS.n8980 VSS.t2607 8.06917
R1143 VSS.n8984 VSS.t2513 8.06917
R1144 VSS.n8984 VSS.t1824 8.06917
R1145 VSS.n8985 VSS.t2859 8.06917
R1146 VSS.n8985 VSS.t2144 8.06917
R1147 VSS.n8993 VSS.t1681 8.06917
R1148 VSS.n8993 VSS.t909 8.06917
R1149 VSS.n8994 VSS.t1260 8.06917
R1150 VSS.n8994 VSS.t3631 8.06917
R1151 VSS.n8998 VSS.t2621 8.06917
R1152 VSS.n8998 VSS.t1927 8.06917
R1153 VSS.n9004 VSS.t2176 8.06917
R1154 VSS.n8970 VSS.t3211 8.06917
R1155 VSS.n1565 VSS.t3477 8.06917
R1156 VSS.n8966 VSS.t2801 8.06917
R1157 VSS.n1553 VSS.t990 8.06917
R1158 VSS.n9096 VSS.t2072 8.06917
R1159 VSS.n8972 VSS.t1671 8.06917
R1160 VSS.n8971 VSS.t497 8.06917
R1161 VSS.n9080 VSS.t3075 8.06917
R1162 VSS.n9080 VSS.t983 8.06917
R1163 VSS.n9077 VSS.t2246 8.06917
R1164 VSS.n9077 VSS.t3289 8.06917
R1165 VSS.n9076 VSS.t2559 8.06917
R1166 VSS.n9076 VSS.t3623 8.06917
R1167 VSS.n9107 VSS.t1409 8.06917
R1168 VSS.n9107 VSS.t2432 8.06917
R1169 VSS.n9106 VSS.t948 8.06917
R1170 VSS.n9106 VSS.t2029 8.06917
R1171 VSS.n9103 VSS.t2334 8.06917
R1172 VSS.n9103 VSS.t3369 8.06917
R1173 VSS.n9080 VSS.t1510 8.06917
R1174 VSS.n9080 VSS.t3513 8.06917
R1175 VSS.n9077 VSS.t622 8.06917
R1176 VSS.n9077 VSS.t2723 8.06917
R1177 VSS.n9076 VSS.t978 8.06917
R1178 VSS.n9076 VSS.t3055 8.06917
R1179 VSS.n9107 VSS.t2925 8.06917
R1180 VSS.n9107 VSS.t1861 8.06917
R1181 VSS.n9106 VSS.t2474 8.06917
R1182 VSS.n9106 VSS.t1471 8.06917
R1183 VSS.n9103 VSS.t747 8.06917
R1184 VSS.n9103 VSS.t2831 8.06917
R1185 VSS.n9085 VSS.t1741 8.06917
R1186 VSS.n9045 VSS.t2797 8.06917
R1187 VSS.n1556 VSS.t2342 8.06917
R1188 VSS.n9041 VSS.t1301 8.06917
R1189 VSS.n9064 VSS.t1106 8.06917
R1190 VSS.n9047 VSS.t2200 8.06917
R1191 VSS.n9070 VSS.t2452 8.06917
R1192 VSS.n9046 VSS.t1773 8.06917
R1193 VSS.n962 VSS.t1298 8.06917
R1194 VSS.n962 VSS.t1029 8.06917
R1195 VSS.n960 VSS.t2094 8.06917
R1196 VSS.n960 VSS.t1863 8.06917
R1197 VSS.n959 VSS.t2497 8.06917
R1198 VSS.n959 VSS.t2272 8.06917
R1199 VSS.n10282 VSS.t2977 8.06917
R1200 VSS.n10282 VSS.t2725 8.06917
R1201 VSS.n10281 VSS.t1727 8.06917
R1202 VSS.n10281 VSS.t1502 8.06917
R1203 VSS.n10279 VSS.t3397 8.06917
R1204 VSS.n10279 VSS.t3185 8.06917
R1205 VSS.n953 VSS.t2160 8.06917
R1206 VSS.n971 VSS.t1919 8.06917
R1207 VSS.n954 VSS.t1395 8.06917
R1208 VSS.n965 VSS.t2190 8.06917
R1209 VSS.n950 VSS.t2571 8.06917
R1210 VSS.n950 VSS.t2707 8.06917
R1211 VSS.n947 VSS.t3341 8.06917
R1212 VSS.n947 VSS.t3471 8.06917
R1213 VSS.n946 VSS.t648 8.06917
R1214 VSS.n946 VSS.t779 8.06917
R1215 VSS.n10252 VSS.t1133 8.06917
R1216 VSS.n10252 VSS.t1269 8.06917
R1217 VSS.n10253 VSS.t3019 8.06917
R1218 VSS.n10253 VSS.t3121 8.06917
R1219 VSS.n10257 VSS.t1649 8.06917
R1220 VSS.n10257 VSS.t1759 8.06917
R1221 VSS.n950 VSS.t3039 8.06917
R1222 VSS.n950 VSS.t708 8.06917
R1223 VSS.n947 VSS.t688 8.06917
R1224 VSS.n947 VSS.t1559 8.06917
R1225 VSS.n946 VSS.t1137 8.06917
R1226 VSS.n946 VSS.t1963 8.06917
R1227 VSS.n10252 VSS.t1625 8.06917
R1228 VSS.n10252 VSS.t2386 8.06917
R1229 VSS.n10253 VSS.t3409 8.06917
R1230 VSS.n10253 VSS.t1153 8.06917
R1231 VSS.n10257 VSS.t2068 8.06917
R1232 VSS.n10257 VSS.t2899 8.06917
R1233 VSS.n10268 VSS.t1198 8.06917
R1234 VSS.n258 VSS.t921 8.06917
R1235 VSS.n10274 VSS.t3497 8.06917
R1236 VSS.n257 VSS.t1244 8.06917
R1237 VSS.n301 VSS.t3271 8.06917
R1238 VSS.n309 VSS.t3073 8.06917
R1239 VSS.n302 VSS.t2464 8.06917
R1240 VSS.n303 VSS.t2493 8.06917
R1241 VSS.n997 VSS.t1561 8.06917
R1242 VSS.n997 VSS.t1310 8.06917
R1243 VSS.n994 VSS.t2332 8.06917
R1244 VSS.n994 VSS.t2108 8.06917
R1245 VSS.n993 VSS.t2763 8.06917
R1246 VSS.n993 VSS.t2509 8.06917
R1247 VSS.n292 VSS.t3197 8.06917
R1248 VSS.n292 VSS.t2983 8.06917
R1249 VSS.n293 VSS.t1965 8.06917
R1250 VSS.n293 VSS.t1737 8.06917
R1251 VSS.n297 VSS.t491 8.06917
R1252 VSS.n297 VSS.t3407 8.06917
R1253 VSS.n997 VSS.t1999 8.06917
R1254 VSS.n997 VSS.t2019 8.06917
R1255 VSS.n994 VSS.t2809 8.06917
R1256 VSS.n994 VSS.t2845 8.06917
R1257 VSS.n993 VSS.t3203 8.06917
R1258 VSS.n993 VSS.t3233 8.06917
R1259 VSS.n292 VSS.t463 8.06917
R1260 VSS.n292 VSS.t505 8.06917
R1261 VSS.n293 VSS.t2400 8.06917
R1262 VSS.n293 VSS.t2436 8.06917
R1263 VSS.n297 VSS.t1013 8.06917
R1264 VSS.n297 VSS.t1060 8.06917
R1265 VSS.n942 VSS.t1120 8.06917
R1266 VSS.n987 VSS.t875 8.06917
R1267 VSS.n943 VSS.t3385 8.06917
R1268 VSS.n977 VSS.t3427 8.06917
R1269 VSS.n940 VSS.t2378 8.06917
R1270 VSS.n1008 VSS.t2168 8.06917
R1271 VSS.n941 VSS.t1637 8.06917
R1272 VSS.n1002 VSS.t2410 8.06917
R1273 VSS.n937 VSS.t3511 8.06917
R1274 VSS.n937 VSS.t2472 8.06917
R1275 VSS.n934 VSS.t1237 8.06917
R1276 VSS.n934 VSS.t3285 8.06917
R1277 VSS.n933 VSS.t1667 8.06917
R1278 VSS.n933 VSS.t554 8.06917
R1279 VSS.n10231 VSS.t2084 8.06917
R1280 VSS.n10231 VSS.t1056 8.06917
R1281 VSS.n10230 VSS.t815 8.06917
R1282 VSS.n10230 VSS.t2939 8.06917
R1283 VSS.n10227 VSS.t2555 8.06917
R1284 VSS.n10227 VSS.t1575 8.06917
R1285 VSS.n937 VSS.t3487 8.06917
R1286 VSS.n937 VSS.t2222 8.06917
R1287 VSS.n934 VSS.t1212 8.06917
R1288 VSS.n934 VSS.t3047 8.06917
R1289 VSS.n933 VSS.t1651 8.06917
R1290 VSS.n933 VSS.t3415 8.06917
R1291 VSS.n10231 VSS.t2066 8.06917
R1292 VSS.n10231 VSS.t764 8.06917
R1293 VSS.n10230 VSS.t796 8.06917
R1294 VSS.n10230 VSS.t2645 8.06917
R1295 VSS.n10227 VSS.t2541 8.06917
R1296 VSS.n10227 VSS.t1281 8.06917
R1297 VSS.n10218 VSS.t1478 8.06917
R1298 VSS.n10220 VSS.t1208 8.06917
R1299 VSS.n291 VSS.t598 8.06917
R1300 VSS.n315 VSS.t1500 8.06917
R1301 VSS.n10208 VSS.t3173 8.06917
R1302 VSS.n330 VSS.t3199 8.06917
R1303 VSS.n10214 VSS.t3405 8.06917
R1304 VSS.n329 VSS.t3449 8.06917
R1305 VSS.n1030 VSS.t2875 8.06917
R1306 VSS.n1030 VSS.t1855 8.06917
R1307 VSS.n1027 VSS.t468 8.06917
R1308 VSS.n1027 VSS.t2637 8.06917
R1309 VSS.n1026 VSS.t960 8.06917
R1310 VSS.n1026 VSS.t3095 8.06917
R1311 VSS.n10192 VSS.t1457 8.06917
R1312 VSS.n10192 VSS.t3493 8.06917
R1313 VSS.n10193 VSS.t3265 8.06917
R1314 VSS.n10193 VSS.t2268 8.06917
R1315 VSS.n10197 VSS.t1923 8.06917
R1316 VSS.n10197 VSS.t863 8.06917
R1317 VSS.n1030 VSS.t2166 8.06917
R1318 VSS.n1030 VSS.t1115 8.06917
R1319 VSS.n1027 VSS.t2975 8.06917
R1320 VSS.n1027 VSS.t1945 8.06917
R1321 VSS.n1026 VSS.t3335 8.06917
R1322 VSS.n1026 VSS.t2344 8.06917
R1323 VSS.n10192 VSS.t680 8.06917
R1324 VSS.n10192 VSS.t2819 8.06917
R1325 VSS.n10193 VSS.t2565 8.06917
R1326 VSS.n10193 VSS.t1579 8.06917
R1327 VSS.n10197 VSS.t1206 8.06917
R1328 VSS.n10197 VSS.t3267 8.06917
R1329 VSS.n929 VSS.t1002 8.06917
R1330 VSS.n1020 VSS.t1041 8.06917
R1331 VSS.n930 VSS.t1307 8.06917
R1332 VSS.n1014 VSS.t1348 8.06917
R1333 VSS.n927 VSS.t2310 8.06917
R1334 VSS.n1045 VSS.t2338 8.06917
R1335 VSS.n928 VSS.t2951 8.06917
R1336 VSS.n1035 VSS.t1931 8.06917
R1337 VSS.n924 VSS.t2721 8.06917
R1338 VSS.n924 VSS.t2747 8.06917
R1339 VSS.n921 VSS.t3505 8.06917
R1340 VSS.n921 VSS.t3537 8.06917
R1341 VSS.n920 VSS.t812 8.06917
R1342 VSS.n920 VSS.t841 8.06917
R1343 VSS.n376 VSS.t1287 8.06917
R1344 VSS.n376 VSS.t1336 8.06917
R1345 VSS.n377 VSS.t3145 8.06917
R1346 VSS.n377 VSS.t3169 8.06917
R1347 VSS.n381 VSS.t1787 8.06917
R1348 VSS.n381 VSS.t1812 8.06917
R1349 VSS.n924 VSS.t1130 8.06917
R1350 VSS.n924 VSS.t881 8.06917
R1351 VSS.n921 VSS.t1953 8.06917
R1352 VSS.n921 VSS.t1721 8.06917
R1353 VSS.n920 VSS.t2358 8.06917
R1354 VSS.n920 VSS.t2132 8.06917
R1355 VSS.n376 VSS.t2829 8.06917
R1356 VSS.n376 VSS.t2563 8.06917
R1357 VSS.n377 VSS.t1595 8.06917
R1358 VSS.n377 VSS.t1342 8.06917
R1359 VSS.n381 VSS.t3277 8.06917
R1360 VSS.n381 VSS.t3079 8.06917
R1361 VSS.n364 VSS.t1393 8.06917
R1362 VSS.n372 VSS.t1427 8.06917
R1363 VSS.n365 VSS.t1989 8.06917
R1364 VSS.n366 VSS.t937 8.06917
R1365 VSS.n10158 VSS.t3379 8.06917
R1366 VSS.n10160 VSS.t3419 8.06917
R1367 VSS.n363 VSS.t508 8.06917
R1368 VSS.n387 VSS.t2675 8.06917
R1369 VSS.n1067 VSS.t1390 8.06917
R1370 VSS.n1067 VSS.t1431 8.06917
R1371 VSS.n1064 VSS.t2180 8.06917
R1372 VSS.n1064 VSS.t2210 8.06917
R1373 VSS.n1063 VSS.t2577 8.06917
R1374 VSS.n1063 VSS.t2615 8.06917
R1375 VSS.n10171 VSS.t3051 8.06917
R1376 VSS.n10171 VSS.t3099 8.06917
R1377 VSS.n10170 VSS.t1808 8.06917
R1378 VSS.n10170 VSS.t1837 8.06917
R1379 VSS.n10167 VSS.t3499 8.06917
R1380 VSS.n10167 VSS.t3533 8.06917
R1381 VSS.n1067 VSS.t2384 8.06917
R1382 VSS.n1067 VSS.t2174 8.06917
R1383 VSS.n1064 VSS.t3193 8.06917
R1384 VSS.n1064 VSS.t2979 8.06917
R1385 VSS.n1063 VSS.t3609 8.06917
R1386 VSS.n1063 VSS.t3343 8.06917
R1387 VSS.n10171 VSS.t951 8.06917
R1388 VSS.n10171 VSS.t694 8.06917
R1389 VSS.n10170 VSS.t2843 8.06917
R1390 VSS.n10170 VSS.t2573 8.06917
R1391 VSS.n10167 VSS.t1488 8.06917
R1392 VSS.n10167 VSS.t1216 8.06917
R1393 VSS.n916 VSS.t1283 8.06917
R1394 VSS.n1057 VSS.t1328 8.06917
R1395 VSS.n917 VSS.t1569 8.06917
R1396 VSS.n1051 VSS.t3611 8.06917
R1397 VSS.n914 VSS.t2679 8.06917
R1398 VSS.n1078 VSS.t3465 8.06917
R1399 VSS.n915 VSS.t2148 8.06917
R1400 VSS.n1072 VSS.t1909 8.06917
R1401 VSS.n911 VSS.t2651 8.06917
R1402 VSS.n911 VSS.t3429 8.06917
R1403 VSS.n908 VSS.t3417 8.06917
R1404 VSS.n908 VSS.t1159 8.06917
R1405 VSS.n907 VSS.t744 8.06917
R1406 VSS.n907 VSS.t1614 8.06917
R1407 VSS.n10132 VSS.t1235 8.06917
R1408 VSS.n10132 VSS.t2027 8.06917
R1409 VSS.n10133 VSS.t3103 8.06917
R1410 VSS.n10133 VSS.t752 8.06917
R1411 VSS.n10137 VSS.t1713 8.06917
R1412 VSS.n10137 VSS.t2491 8.06917
R1413 VSS.n911 VSS.t645 8.06917
R1414 VSS.n911 VSS.t3545 8.06917
R1415 VSS.n908 VSS.t1530 8.06917
R1416 VSS.n908 VSS.t1275 8.06917
R1417 VSS.n907 VSS.t1939 8.06917
R1418 VSS.n907 VSS.t1703 8.06917
R1419 VSS.n10132 VSS.t2360 8.06917
R1420 VSS.n10132 VSS.t2136 8.06917
R1421 VSS.n10133 VSS.t1104 8.06917
R1422 VSS.n10133 VSS.t857 8.06917
R1423 VSS.n10137 VSS.t2861 8.06917
R1424 VSS.n10137 VSS.t2599 8.06917
R1425 VSS.n10148 VSS.t1747 8.06917
R1426 VSS.n402 VSS.t2527 8.06917
R1427 VSS.n10154 VSS.t1186 8.06917
R1428 VSS.n401 VSS.t917 8.06917
R1429 VSS.n1283 VSS.t3321 8.06917
R1430 VSS.n1291 VSS.t3129 8.06917
R1431 VSS.n1284 VSS.t3617 8.06917
R1432 VSS.n1285 VSS.t3353 8.06917
R1433 VSS.n1104 VSS.t1277 8.06917
R1434 VSS.n1104 VSS.t994 8.06917
R1435 VSS.n1101 VSS.t2060 8.06917
R1436 VSS.n1101 VSS.t1841 8.06917
R1437 VSS.n1100 VSS.t2466 8.06917
R1438 VSS.n1100 VSS.t2244 8.06917
R1439 VSS.n1274 VSS.t2949 8.06917
R1440 VSS.n1274 VSS.t2709 8.06917
R1441 VSS.n1275 VSS.t1705 8.06917
R1442 VSS.n1275 VSS.t1480 8.06917
R1443 VSS.n1279 VSS.t3375 8.06917
R1444 VSS.n1279 VSS.t3167 8.06917
R1445 VSS.n1104 VSS.t1291 8.06917
R1446 VSS.n1104 VSS.t2102 8.06917
R1447 VSS.n1101 VSS.t2086 8.06917
R1448 VSS.n1101 VSS.t2909 8.06917
R1449 VSS.n1100 VSS.t2489 8.06917
R1450 VSS.n1100 VSS.t3293 8.06917
R1451 VSS.n1274 VSS.t2971 8.06917
R1452 VSS.n1274 VSS.t608 8.06917
R1453 VSS.n1275 VSS.t1723 8.06917
R1454 VSS.n1275 VSS.t2501 8.06917
R1455 VSS.n1279 VSS.t3393 8.06917
R1456 VSS.n1279 VSS.t1126 8.06917
R1457 VSS.n903 VSS.t1222 8.06917
R1458 VSS.n1094 VSS.t954 8.06917
R1459 VSS.n904 VSS.t1512 8.06917
R1460 VSS.n1084 VSS.t1253 8.06917
R1461 VSS.n901 VSS.t2937 8.06917
R1462 VSS.n1115 VSS.t2691 8.06917
R1463 VSS.n902 VSS.t1363 8.06917
R1464 VSS.n1109 VSS.t2156 8.06917
R1465 VSS.n878 VSS.t3509 8.06917
R1466 VSS.n1127 VSS.t3615 8.06917
R1467 VSS.n879 VSS.t3109 8.06917
R1468 VSS.n1121 VSS.t759 8.06917
R1469 VSS.n863 VSS.t2873 8.06917
R1470 VSS.n837 VSS.t2611 8.06917
R1471 VSS.n870 VSS.t2050 8.06917
R1472 VSS.n836 VSS.t2078 8.06917
R1473 VSS.n10923 VSS.t611 8.06917
R1474 VSS.n222 VSS.t3517 8.06917
R1475 VSS.n839 VSS.t2995 8.06917
R1476 VSS.n838 VSS.t635 8.06917
R1477 VSS.n858 VSS.t3241 8.06917
R1478 VSS.n858 VSS.t3033 8.06917
R1479 VSS.n855 VSS.t935 8.06917
R1480 VSS.n855 VSS.t675 8.06917
R1481 VSS.n854 VSS.t1413 8.06917
R1482 VSS.n854 VSS.t1124 8.06917
R1483 VSS.n848 VSS.t1843 8.06917
R1484 VSS.n848 VSS.t1618 8.06917
R1485 VSS.n847 VSS.t482 8.06917
R1486 VSS.n847 VSS.t3399 8.06917
R1487 VSS.n858 VSS.t541 8.06917
R1488 VSS.n858 VSS.t578 8.06917
R1489 VSS.n855 VSS.t1449 8.06917
R1490 VSS.n855 VSS.t1482 8.06917
R1491 VSS.n854 VSS.t1849 8.06917
R1492 VSS.n854 VSS.t1879 8.06917
R1493 VSS.n848 VSS.t2276 8.06917
R1494 VSS.n848 VSS.t2304 8.06917
R1495 VSS.n847 VSS.t1007 8.06917
R1496 VSS.n847 VSS.t1052 8.06917
R1497 VSS.n1135 VSS.t1202 8.06917
R1498 VSS.n1135 VSS.t931 8.06917
R1499 VSS.n1139 VSS.t2005 8.06917
R1500 VSS.n1139 VSS.t1785 8.06917
R1501 VSS.n1140 VSS.t2412 8.06917
R1502 VSS.n1140 VSS.t2196 8.06917
R1503 VSS.n1149 VSS.t2883 8.06917
R1504 VSS.n1149 VSS.t2623 8.06917
R1505 VSS.n1148 VSS.t1645 8.06917
R1506 VSS.n1148 VSS.t1411 8.06917
R1507 VSS.n1135 VSS.t1305 8.06917
R1508 VSS.n1135 VSS.t2114 8.06917
R1509 VSS.n1139 VSS.t2104 8.06917
R1510 VSS.n1139 VSS.t2917 8.06917
R1511 VSS.n1140 VSS.t2505 8.06917
R1512 VSS.n1140 VSS.t3299 8.06917
R1513 VSS.n1149 VSS.t2981 8.06917
R1514 VSS.n1149 VSS.t619 8.06917
R1515 VSS.n1148 VSS.t1735 8.06917
R1516 VSS.n1148 VSS.t2519 8.06917
R1517 VSS.n898 VSS.t3027 8.06917
R1518 VSS.n898 VSS.t2777 8.06917
R1519 VSS.n895 VSS.t670 8.06917
R1520 VSS.n895 VSS.t3563 8.06917
R1521 VSS.n894 VSS.t1118 8.06917
R1522 VSS.n894 VSS.t872 8.06917
R1523 VSS.n888 VSS.t1606 8.06917
R1524 VSS.n888 VSS.t1368 8.06917
R1525 VSS.n887 VSS.t3389 8.06917
R1526 VSS.n887 VSS.t3181 8.06917
R1527 VSS.n898 VSS.t3011 8.06917
R1528 VSS.n898 VSS.t654 8.06917
R1529 VSS.n895 VSS.t642 8.06917
R1530 VSS.n895 VSS.t1534 8.06917
R1531 VSS.n894 VSS.t1102 8.06917
R1532 VSS.n894 VSS.t1941 8.06917
R1533 VSS.n888 VSS.t1591 8.06917
R1534 VSS.n888 VSS.t2370 8.06917
R1535 VSS.n887 VSS.t3377 8.06917
R1536 VSS.n887 VSS.t1111 8.06917
R1537 VSS.n10353 VSS.t3451 8.06917
R1538 VSS.n10361 VSS.t2170 8.06917
R1539 VSS.n10354 VSS.t1180 8.06917
R1540 VSS.n10355 VSS.t1973 8.06917
R1541 VSS.n10666 VSS.t587 8.06917
R1542 VSS.n10338 VSS.t683 8.06917
R1543 VSS.n10337 VSS.t3541 8.06917
R1544 VSS.n10673 VSS.t3269 8.06917
R1545 VSS.n10336 VSS.t2306 8.06917
R1546 VSS.n10909 VSS.t1583 8.06917
R1547 VSS.n10909 VSS.t1338 8.06917
R1548 VSS.n10906 VSS.t2346 8.06917
R1549 VSS.n10906 VSS.t2130 8.06917
R1550 VSS.n10905 VSS.t2791 8.06917
R1551 VSS.n10905 VSS.t2537 8.06917
R1552 VSS.n10899 VSS.t3213 8.06917
R1553 VSS.n10899 VSS.t2999 8.06917
R1554 VSS.n10898 VSS.t1987 8.06917
R1555 VSS.n10898 VSS.t1763 8.06917
R1556 VSS.n10909 VSS.t2314 8.06917
R1557 VSS.n10909 VSS.t1322 8.06917
R1558 VSS.n10906 VSS.t3139 8.06917
R1559 VSS.n10906 VSS.t2112 8.06917
R1560 VSS.n10905 VSS.t3535 8.06917
R1561 VSS.n10905 VSS.t2515 8.06917
R1562 VSS.n10899 VSS.t868 8.06917
R1563 VSS.n10899 VSS.t2989 8.06917
R1564 VSS.n10898 VSS.t2741 8.06917
R1565 VSS.n10898 VSS.t1749 8.06917
R1566 VSS.n11003 VSS.t3607 8.06917
R1567 VSS.n11003 VSS.t2597 8.06917
R1568 VSS.n11007 VSS.t1344 8.06917
R1569 VSS.n11007 VSS.t3367 8.06917
R1570 VSS.n11008 VSS.t1771 8.06917
R1571 VSS.n11008 VSS.t685 8.06917
R1572 VSS.n11016 VSS.t2202 8.06917
R1573 VSS.n11016 VSS.t1172 8.06917
R1574 VSS.n11017 VSS.t912 8.06917
R1575 VSS.n11017 VSS.t3043 8.06917
R1576 VSS.n11003 VSS.t3247 8.06917
R1577 VSS.n11003 VSS.t2250 8.06917
R1578 VSS.n11007 VSS.t946 8.06917
R1579 VSS.n11007 VSS.t3077 8.06917
R1580 VSS.n11008 VSS.t1423 8.06917
R1581 VSS.n11008 VSS.t3439 8.06917
R1582 VSS.n11016 VSS.t1851 8.06917
R1583 VSS.n11016 VSS.t788 8.06917
R1584 VSS.n11017 VSS.t499 8.06917
R1585 VSS.n11017 VSS.t2669 8.06917
R1586 VSS.n11060 VSS.t697 8.06917
R1587 VSS.n11060 VSS.t737 8.06917
R1588 VSS.n11064 VSS.t1549 8.06917
R1589 VSS.n11064 VSS.t1587 8.06917
R1590 VSS.n11065 VSS.t1959 8.06917
R1591 VSS.n11065 VSS.t1995 8.06917
R1592 VSS.n11073 VSS.t2380 8.06917
R1593 VSS.n11073 VSS.t2418 8.06917
R1594 VSS.n11074 VSS.t1141 8.06917
R1595 VSS.n11074 VSS.t1176 8.06917
R1596 VSS.n11060 VSS.t2264 8.06917
R1597 VSS.n11060 VSS.t2011 8.06917
R1598 VSS.n11064 VSS.t3087 8.06917
R1599 VSS.n11064 VSS.t2833 8.06917
R1600 VSS.n11065 VSS.t3455 8.06917
R1601 VSS.n11065 VSS.t3225 8.06917
R1602 VSS.n11073 VSS.t799 8.06917
R1603 VSS.n11073 VSS.t494 8.06917
R1604 VSS.n11074 VSS.t2687 8.06917
R1605 VSS.n11074 VSS.t2424 8.06917
R1606 VSS.n1320 VSS.t1993 8.06917
R1607 VSS.t1993 VSS.n1319 8.06917
R1608 VSS.n1322 VSS.t1194 8.06917
R1609 VSS.t1194 VSS.n1321 8.06917
R1610 VSS.n1324 VSS.t1353 8.06917
R1611 VSS.t1353 VSS.n1323 8.06917
R1612 VSS.n1326 VSS.t3633 8.06917
R1613 VSS.t3633 VSS.n1325 8.06917
R1614 VSS.n1333 VSS.t2865 8.06917
R1615 VSS.t2865 VSS.n1332 8.06917
R1616 VSS.t2058 VSS.n9509 8.06917
R1617 VSS.n9510 VSS.t2058 8.06917
R1618 VSS.n9508 VSS.t2208 8.06917
R1619 VSS.t2208 VSS.n9507 8.06917
R1620 VSS.t1445 VSS.n9504 8.06917
R1621 VSS.n9505 VSS.t1445 8.06917
R1622 VSS.t749 VSS.n9501 8.06917
R1623 VSS.n9502 VSS.t749 8.06917
R1624 VSS.t1802 VSS.n9497 8.06917
R1625 VSS.n9498 VSS.t1802 8.06917
R1626 VSS.n1377 VSS.t2192 8.06917
R1627 VSS.t2192 VSS.n1376 8.06917
R1628 VSS.t1765 VSS.n9624 8.06917
R1629 VSS.n9625 VSS.t1765 8.06917
R1630 VSS.t1885 VSS.n9622 8.06917
R1631 VSS.n9623 VSS.t1885 8.06917
R1632 VSS.t1071 VSS.n9620 8.06917
R1633 VSS.n9621 VSS.t1071 8.06917
R1634 VSS.t3359 VSS.n9618 8.06917
R1635 VSS.n9619 VSS.t3359 8.06917
R1636 VSS.n815 VSS.t3525 8.06917
R1637 VSS.t3525 VSS.n810 8.06917
R1638 VSS.t2907 VSS.n9608 8.06917
R1639 VSS.n9609 VSS.t2907 8.06917
R1640 VSS.t2116 VSS.n9606 8.06917
R1641 VSS.n9607 VSS.t2116 8.06917
R1642 VSS.t1526 VSS.n9604 8.06917
R1643 VSS.n9605 VSS.t1526 8.06917
R1644 VSS.t668 VSS.n9602 8.06917
R1645 VSS.n9603 VSS.t668 8.06917
R1646 VSS.n9624 VSS.t547 8.06917
R1647 VSS.n9625 VSS.t547 8.06917
R1648 VSS.n9622 VSS.t728 8.06917
R1649 VSS.n9623 VSS.t728 8.06917
R1650 VSS.n9620 VSS.t3089 8.06917
R1651 VSS.n9621 VSS.t3089 8.06917
R1652 VSS.n9618 VSS.t2270 8.06917
R1653 VSS.n9619 VSS.t2270 8.06917
R1654 VSS.n815 VSS.t2388 8.06917
R1655 VSS.t2388 VSS.n810 8.06917
R1656 VSS.n9608 VSS.t1795 8.06917
R1657 VSS.n9609 VSS.t1795 8.06917
R1658 VSS.n9606 VSS.t968 8.06917
R1659 VSS.n9607 VSS.t968 8.06917
R1660 VSS.n9604 VSS.t3445 8.06917
R1661 VSS.n9605 VSS.t3445 8.06917
R1662 VSS.n9602 VSS.t2705 8.06917
R1663 VSS.n9603 VSS.t2705 8.06917
R1664 VSS.t1743 VSS.n9648 8.06917
R1665 VSS.n9649 VSS.t1743 8.06917
R1666 VSS.t1869 VSS.n9646 8.06917
R1667 VSS.n9647 VSS.t1869 8.06917
R1668 VSS.t1054 VSS.n9644 8.06917
R1669 VSS.n9645 VSS.t1054 8.06917
R1670 VSS.t3337 VSS.n649 8.06917
R1671 VSS.n9643 VSS.t3337 8.06917
R1672 VSS.n9886 VSS.t3501 8.06917
R1673 VSS.t3501 VSS.n9885 8.06917
R1674 VSS.n779 VSS.t2895 8.06917
R1675 VSS.t2895 VSS.n778 8.06917
R1676 VSS.n781 VSS.t2092 8.06917
R1677 VSS.t2092 VSS.n780 8.06917
R1678 VSS.n783 VSS.t1514 8.06917
R1679 VSS.t1514 VSS.n782 8.06917
R1680 VSS.n785 VSS.t640 8.06917
R1681 VSS.t640 VSS.n784 8.06917
R1682 VSS.n9648 VSS.t516 8.06917
R1683 VSS.n9649 VSS.t516 8.06917
R1684 VSS.n9646 VSS.t706 8.06917
R1685 VSS.n9647 VSS.t706 8.06917
R1686 VSS.n9644 VSS.t3063 8.06917
R1687 VSS.n9645 VSS.t3063 8.06917
R1688 VSS.t2260 VSS.n649 8.06917
R1689 VSS.n9643 VSS.t2260 8.06917
R1690 VSS.n9886 VSS.t2374 8.06917
R1691 VSS.n9885 VSS.t2374 8.06917
R1692 VSS.n779 VSS.t1781 8.06917
R1693 VSS.n778 VSS.t1781 8.06917
R1694 VSS.n781 VSS.t939 8.06917
R1695 VSS.n780 VSS.t939 8.06917
R1696 VSS.n783 VSS.t3421 8.06917
R1697 VSS.n782 VSS.t3421 8.06917
R1698 VSS.n785 VSS.t2667 8.06917
R1699 VSS.n784 VSS.t2667 8.06917
R1700 VSS.t1917 VSS.n9692 8.06917
R1701 VSS.n9693 VSS.t1917 8.06917
R1702 VSS.t1098 VSS.n9689 8.06917
R1703 VSS.n9690 VSS.t1098 8.06917
R1704 VSS.t3381 VSS.n9686 8.06917
R1705 VSS.n9687 VSS.t3381 8.06917
R1706 VSS.t3551 VSS.n9683 8.06917
R1707 VSS.n9684 VSS.t3551 8.06917
R1708 VSS.n1179 VSS.t2785 8.06917
R1709 VSS.t2785 VSS.n654 8.06917
R1710 VSS.t2150 VSS.n9852 8.06917
R1711 VSS.n9853 VSS.t2150 8.06917
R1712 VSS.t1378 VSS.n9849 8.06917
R1713 VSS.n9850 VSS.t1378 8.06917
R1714 VSS.t717 VSS.n9846 8.06917
R1715 VSS.n9847 VSS.t717 8.06917
R1716 VSS.t3083 VSS.n9843 8.06917
R1717 VSS.n9844 VSS.t3083 8.06917
R1718 VSS.n9691 VSS.t828 8.06917
R1719 VSS.t828 VSS.n9671 8.06917
R1720 VSS.n9688 VSS.t970 8.06917
R1721 VSS.t970 VSS.n9674 8.06917
R1722 VSS.n9685 VSS.t3283 8.06917
R1723 VSS.t3283 VSS.n9677 8.06917
R1724 VSS.t2495 VSS.n653 8.06917
R1725 VSS.n9680 VSS.t2495 8.06917
R1726 VSS.n1178 VSS.t2641 8.06917
R1727 VSS.t2641 VSS.n1177 8.06917
R1728 VSS.n9851 VSS.t2009 8.06917
R1729 VSS.t2009 VSS.n680 8.06917
R1730 VSS.n9848 VSS.t1246 8.06917
R1731 VSS.t1246 VSS.n683 8.06917
R1732 VSS.n9845 VSS.t544 8.06917
R1733 VSS.t544 VSS.n686 8.06917
R1734 VSS.n9842 VSS.t2945 8.06917
R1735 VSS.t2945 VSS.n689 8.06917
R1736 VSS.n661 VSS.t3473 8.06917
R1737 VSS.t3473 VSS.n578 8.06917
R1738 VSS.n663 VSS.t2717 8.06917
R1739 VSS.t2717 VSS.n662 8.06917
R1740 VSS.n665 VSS.t1933 8.06917
R1741 VSS.t1933 VSS.n664 8.06917
R1742 VSS.n667 VSS.t2048 8.06917
R1743 VSS.t2048 VSS.n666 8.06917
R1744 VSS.n673 VSS.t1273 8.06917
R1745 VSS.t1273 VSS.n668 8.06917
R1746 VSS.t565 VSS.n9870 8.06917
R1747 VSS.n9871 VSS.t565 8.06917
R1748 VSS.t2953 VSS.n9868 8.06917
R1749 VSS.n9869 VSS.t2953 8.06917
R1750 VSS.t2320 VSS.n9866 8.06917
R1751 VSS.n9867 VSS.t2320 8.06917
R1752 VSS.t1563 VSS.n9864 8.06917
R1753 VSS.n9865 VSS.t1563 8.06917
R1754 VSS.n661 VSS.t2354 8.06917
R1755 VSS.t2354 VSS.n578 8.06917
R1756 VSS.n663 VSS.t1604 8.06917
R1757 VSS.n662 VSS.t1604 8.06917
R1758 VSS.n665 VSS.t757 8.06917
R1759 VSS.n664 VSS.t757 8.06917
R1760 VSS.n667 VSS.t898 8.06917
R1761 VSS.n666 VSS.t898 8.06917
R1762 VSS.n673 VSS.t3223 8.06917
R1763 VSS.t3223 VSS.n668 8.06917
R1764 VSS.n9870 VSS.t2593 8.06917
R1765 VSS.n9871 VSS.t2593 8.06917
R1766 VSS.n9868 VSS.t1831 8.06917
R1767 VSS.n9869 VSS.t1831 8.06917
R1768 VSS.n9866 VSS.t1210 8.06917
R1769 VSS.n9867 VSS.t1210 8.06917
R1770 VSS.n9864 VSS.t3503 8.06917
R1771 VSS.n9865 VSS.t3503 8.06917
R1772 VSS.t2414 VSS.n9965 8.06917
R1773 VSS.n9966 VSS.t2414 8.06917
R1774 VSS.t1657 VSS.n9963 8.06917
R1775 VSS.n9964 VSS.t1657 8.06917
R1776 VSS.t824 VSS.n9961 8.06917
R1777 VSS.n9962 VSS.t824 8.06917
R1778 VSS.t958 VSS.n9959 8.06917
R1779 VSS.n9960 VSS.t958 8.06917
R1780 VSS.n141 VSS.t3273 8.06917
R1781 VSS.t3273 VSS.n140 8.06917
R1782 VSS.n11188 VSS.t2657 8.06917
R1783 VSS.t2657 VSS.n11187 8.06917
R1784 VSS.n11190 VSS.t1881 8.06917
R1785 VSS.t1881 VSS.n11189 8.06917
R1786 VSS.n11192 VSS.t1271 8.06917
R1787 VSS.t1271 VSS.n11191 8.06917
R1788 VSS.n11194 VSS.t3561 8.06917
R1789 VSS.t3561 VSS.n11193 8.06917
R1790 VSS.n9965 VSS.t1313 8.06917
R1791 VSS.n9966 VSS.t1313 8.06917
R1792 VSS.n9963 VSS.t3591 8.06917
R1793 VSS.n9964 VSS.t3591 8.06917
R1794 VSS.n9961 VSS.t2835 8.06917
R1795 VSS.n9962 VSS.t2835 8.06917
R1796 VSS.n9959 VSS.t2967 8.06917
R1797 VSS.n9960 VSS.t2967 8.06917
R1798 VSS.n141 VSS.t2178 8.06917
R1799 VSS.t2178 VSS.n140 8.06917
R1800 VSS.n11188 VSS.t1553 8.06917
R1801 VSS.n11187 VSS.t1553 8.06917
R1802 VSS.n11190 VSS.t720 8.06917
R1803 VSS.n11189 VSS.t720 8.06917
R1804 VSS.n11192 VSS.t3221 8.06917
R1805 VSS.n11191 VSS.t3221 8.06917
R1806 VSS.n11194 VSS.t2440 8.06917
R1807 VSS.n11193 VSS.t2440 8.06917
R1808 VSS.n1261 VSS.t2533 8.06917
R1809 VSS.t2533 VSS.n1260 8.06917
R1810 VSS.n1263 VSS.t1777 8.06917
R1811 VSS.t1777 VSS.n1262 8.06917
R1812 VSS.n1265 VSS.t1895 8.06917
R1813 VSS.t1895 VSS.n1264 8.06917
R1814 VSS.n1267 VSS.t1079 8.06917
R1815 VSS.t1079 VSS.n1266 8.06917
R1816 VSS.n9520 VSS.t3371 8.06917
R1817 VSS.t3371 VSS.n9519 8.06917
R1818 VSS.t2617 VSS.n1246 8.06917
R1819 VSS.n1247 VSS.t2617 8.06917
R1820 VSS.t2753 VSS.n1244 8.06917
R1821 VSS.n1245 VSS.t2753 8.06917
R1822 VSS.t1971 VSS.n1242 8.06917
R1823 VSS.n1243 VSS.t1971 8.06917
R1824 VSS.t1359 VSS.n804 8.06917
R1825 VSS.n1241 VSS.t1359 8.06917
R1826 VSS.n1261 VSS.t1419 8.06917
R1827 VSS.n1260 VSS.t1419 8.06917
R1828 VSS.n1263 VSS.t510 8.06917
R1829 VSS.n1262 VSS.t510 8.06917
R1830 VSS.n1265 VSS.t701 8.06917
R1831 VSS.n1264 VSS.t701 8.06917
R1832 VSS.n1267 VSS.t3059 8.06917
R1833 VSS.n1266 VSS.t3059 8.06917
R1834 VSS.n9520 VSS.t2258 8.06917
R1835 VSS.n9519 VSS.t2258 8.06917
R1836 VSS.n1246 VSS.t1492 8.06917
R1837 VSS.n1247 VSS.t1492 8.06917
R1838 VSS.n1244 VSS.t1633 8.06917
R1839 VSS.n1245 VSS.t1633 8.06917
R1840 VSS.n1242 VSS.t782 8.06917
R1841 VSS.n1243 VSS.t782 8.06917
R1842 VSS.t3259 VSS.n804 8.06917
R1843 VSS.n1241 VSS.t3259 8.06917
R1844 VSS.n635 VSS.t2368 8.06917
R1845 VSS.t2368 VSS.n634 8.06917
R1846 VSS.n637 VSS.t1608 8.06917
R1847 VSS.t1608 VSS.n636 8.06917
R1848 VSS.n639 VSS.t1733 8.06917
R1849 VSS.t1733 VSS.n638 8.06917
R1850 VSS.n641 VSS.t907 8.06917
R1851 VSS.t907 VSS.n640 8.06917
R1852 VSS.t3227 VSS.n9893 8.06917
R1853 VSS.n9894 VSS.t3227 8.06917
R1854 VSS.n9655 VSS.t2446 8.06917
R1855 VSS.t2446 VSS.n9654 8.06917
R1856 VSS.n9657 VSS.t2575 8.06917
R1857 VSS.t2575 VSS.n9656 8.06917
R1858 VSS.n9659 VSS.t1814 8.06917
R1859 VSS.t1814 VSS.n9658 8.06917
R1860 VSS.n9661 VSS.t1164 8.06917
R1861 VSS.t1164 VSS.n9660 8.06917
R1862 VSS.n635 VSS.t1224 8.06917
R1863 VSS.n634 VSS.t1224 8.06917
R1864 VSS.n637 VSS.t3521 8.06917
R1865 VSS.n636 VSS.t3521 8.06917
R1866 VSS.n639 VSS.t471 8.06917
R1867 VSS.n638 VSS.t471 8.06917
R1868 VSS.n641 VSS.t2887 8.06917
R1869 VSS.n640 VSS.t2887 8.06917
R1870 VSS.n9893 VSS.t2082 8.06917
R1871 VSS.n9894 VSS.t2082 8.06917
R1872 VSS.n9655 VSS.t1315 8.06917
R1873 VSS.n9654 VSS.t1315 8.06917
R1874 VSS.n9657 VSS.t1459 8.06917
R1875 VSS.n9656 VSS.t1459 8.06917
R1876 VSS.n9659 VSS.t583 8.06917
R1877 VSS.n9658 VSS.t583 8.06917
R1878 VSS.n9661 VSS.t3123 8.06917
R1879 VSS.n9660 VSS.t3123 8.06917
R1880 VSS.n601 VSS.t1665 8.06917
R1881 VSS.t1665 VSS.n546 8.06917
R1882 VSS.t826 VSS.n600 8.06917
R1883 VSS.n606 VSS.t826 8.06917
R1884 VSS.t964 VSS.n599 8.06917
R1885 VSS.n611 VSS.t964 8.06917
R1886 VSS.t3279 VSS.n598 8.06917
R1887 VSS.n616 VSS.t3279 8.06917
R1888 VSS.t2485 VSS.n9905 8.06917
R1889 VSS.n9906 VSS.t2485 8.06917
R1890 VSS.t2633 VSS.n9697 8.06917
R1891 VSS.n9698 VSS.t2633 8.06917
R1892 VSS.t1865 VSS.n9696 8.06917
R1893 VSS.n9703 VSS.t1865 8.06917
R1894 VSS.t1050 VSS.n9695 8.06917
R1895 VSS.n9708 VSS.t1050 8.06917
R1896 VSS.t1380 VSS.n9694 8.06917
R1897 VSS.n9713 VSS.t1380 8.06917
R1898 VSS.n605 VSS.t1506 8.06917
R1899 VSS.t1506 VSS.n604 8.06917
R1900 VSS.n610 VSS.t633 8.06917
R1901 VSS.t633 VSS.n609 8.06917
R1902 VSS.n615 VSS.t792 8.06917
R1903 VSS.t792 VSS.n614 8.06917
R1904 VSS.n620 VSS.t3143 8.06917
R1905 VSS.t3143 VSS.n619 8.06917
R1906 VSS.n9904 VSS.t2336 8.06917
R1907 VSS.t2336 VSS.n622 8.06917
R1908 VSS.n9702 VSS.t1585 8.06917
R1909 VSS.t1585 VSS.n9701 8.06917
R1910 VSS.n9707 VSS.t1711 8.06917
R1911 VSS.t1711 VSS.n9706 8.06917
R1912 VSS.n9712 VSS.t886 8.06917
R1913 VSS.t886 VSS.n9711 8.06917
R1914 VSS.n9717 VSS.t3329 8.06917
R1915 VSS.t3329 VSS.n9716 8.06917
R1916 VSS.n591 VSS.t2204 8.06917
R1917 VSS.t2204 VSS.n590 8.06917
R1918 VSS.n593 VSS.t1443 8.06917
R1919 VSS.t1443 VSS.n592 8.06917
R1920 VSS.n595 VSS.t1565 8.06917
R1921 VSS.t1565 VSS.n594 8.06917
R1922 VSS.n597 VSS.t730 8.06917
R1923 VSS.t730 VSS.n596 8.06917
R1924 VSS.t3093 VSS.n583 8.06917
R1925 VSS.n9917 VSS.t3093 8.06917
R1926 VSS.n9928 VSS.t3189 8.06917
R1927 VSS.t3189 VSS.n9927 8.06917
R1928 VSS.n9930 VSS.t2394 8.06917
R1929 VSS.t2394 VSS.n9929 8.06917
R1930 VSS.n9932 VSS.t1643 8.06917
R1931 VSS.t1643 VSS.n9931 8.06917
R1932 VSS.n9934 VSS.t1929 8.06917
R1933 VSS.t1929 VSS.n9933 8.06917
R1934 VSS.n591 VSS.t1015 8.06917
R1935 VSS.n590 VSS.t1015 8.06917
R1936 VSS.n593 VSS.t3311 8.06917
R1937 VSS.n592 VSS.t3311 8.06917
R1938 VSS.n595 VSS.t3467 8.06917
R1939 VSS.n594 VSS.t3467 8.06917
R1940 VSS.n597 VSS.t2713 8.06917
R1941 VSS.n596 VSS.t2713 8.06917
R1942 VSS.t1925 VSS.n583 8.06917
R1943 VSS.n9917 VSS.t1925 8.06917
R1944 VSS.n9928 VSS.t2035 8.06917
R1945 VSS.n9927 VSS.t2035 8.06917
R1946 VSS.n9930 VSS.t1265 8.06917
R1947 VSS.n9929 VSS.t1265 8.06917
R1948 VSS.n9932 VSS.t3555 8.06917
R1949 VSS.n9931 VSS.t3555 8.06917
R1950 VSS.n9934 VSS.t734 8.06917
R1951 VSS.n9933 VSS.t734 8.06917
R1952 VSS.t2821 VSS.n11049 8.06917
R1953 VSS.n11050 VSS.t2821 8.06917
R1954 VSS.t2013 VSS.n11047 8.06917
R1955 VSS.n11048 VSS.t2013 8.06917
R1956 VSS.t2162 VSS.n11045 8.06917
R1957 VSS.n11046 VSS.t2162 8.06917
R1958 VSS.t1386 VSS.n11043 8.06917
R1959 VSS.n11044 VSS.t1386 8.06917
R1960 VSS.n11282 VSS.t476 8.06917
R1961 VSS.t476 VSS.n11281 8.06917
R1962 VSS.n9948 VSS.t666 8.06917
R1963 VSS.t666 VSS.n9947 8.06917
R1964 VSS.n9950 VSS.t3037 8.06917
R1965 VSS.t3037 VSS.n9949 8.06917
R1966 VSS.n9952 VSS.t2226 8.06917
R1967 VSS.t2226 VSS.n9951 8.06917
R1968 VSS.n9954 VSS.t2511 8.06917
R1969 VSS.t2511 VSS.n9953 8.06917
R1970 VSS.n11049 VSS.t1673 8.06917
R1971 VSS.n11050 VSS.t1673 8.06917
R1972 VSS.n11047 VSS.t834 8.06917
R1973 VSS.n11048 VSS.t834 8.06917
R1974 VSS.n11045 VSS.t974 8.06917
R1975 VSS.n11046 VSS.t974 8.06917
R1976 VSS.n11043 VSS.t3287 8.06917
R1977 VSS.n11044 VSS.t3287 8.06917
R1978 VSS.n11282 VSS.t2507 8.06917
R1979 VSS.t2507 VSS.n11281 8.06917
R1980 VSS.n9948 VSS.t2653 8.06917
R1981 VSS.n9947 VSS.t2653 8.06917
R1982 VSS.n9950 VSS.t1877 8.06917
R1983 VSS.n9949 VSS.t1877 8.06917
R1984 VSS.n9952 VSS.t1062 8.06917
R1985 VSS.n9951 VSS.t1062 8.06917
R1986 VSS.n9954 VSS.t1399 8.06917
R1987 VSS.n9953 VSS.t1399 8.06917
R1988 VSS.t3237 VSS.n9476 8.06917
R1989 VSS.n9486 VSS.t3237 8.06917
R1990 VSS.t3355 VSS.n9484 8.06917
R1991 VSS.n9485 VSS.t3355 8.06917
R1992 VSS.t2589 VSS.n9482 8.06917
R1993 VSS.n9483 VSS.t2589 8.06917
R1994 VSS.t1822 VSS.n9480 8.06917
R1995 VSS.n9481 VSS.t1822 8.06917
R1996 VSS.n1387 VSS.t1951 8.06917
R1997 VSS.t1951 VSS.n1386 8.06917
R1998 VSS.n1409 VSS.t1332 8.06917
R1999 VSS.t1332 VSS.n1408 8.06917
R2000 VSS.n1411 VSS.t3613 8.06917
R2001 VSS.t3613 VSS.n1410 8.06917
R2002 VSS.n1413 VSS.t3029 8.06917
R2003 VSS.t3029 VSS.n1412 8.06917
R2004 VSS.n1415 VSS.t2220 8.06917
R2005 VSS.t2220 VSS.n1414 8.06917
R2006 VSS.n11220 VSS.t572 8.06917
R2007 VSS.n11220 VSS.t2671 8.06917
R2008 VSS.n11219 VSS.t923 8.06917
R2009 VSS.n11219 VSS.t3007 8.06917
R2010 VSS.n11213 VSS.t2881 8.06917
R2011 VSS.n11213 VSS.t1816 8.06917
R2012 VSS.n11212 VSS.t2448 8.06917
R2013 VSS.n11212 VSS.t1425 8.06917
R2014 VSS.n11209 VSS.t699 8.06917
R2015 VSS.n11209 VSS.t2773 8.06917
R2016 VSS.n11220 VSS.t1075 8.06917
R2017 VSS.n11220 VSS.t2164 8.06917
R2018 VSS.n11219 VSS.t1447 8.06917
R2019 VSS.n11219 VSS.t2460 8.06917
R2020 VSS.n11213 VSS.t3295 8.06917
R2021 VSS.n11213 VSS.t1289 8.06917
R2022 VSS.n11212 VSS.t2927 8.06917
R2023 VSS.n11212 VSS.t849 8.06917
R2024 VSS.n11209 VSS.t1184 8.06917
R2025 VSS.n11209 VSS.t2254 8.06917
R2026 VSS.n10956 VSS.t2543 8.06917
R2027 VSS.n10956 VSS.t3245 8.06917
R2028 VSS.n10957 VSS.t2889 8.06917
R2029 VSS.n10957 VSS.t3575 8.06917
R2030 VSS.n10965 VSS.t1707 8.06917
R2031 VSS.n10965 VSS.t2382 8.06917
R2032 VSS.n10966 VSS.t1285 8.06917
R2033 VSS.n10966 VSS.t1997 8.06917
R2034 VSS.n10970 VSS.t2647 8.06917
R2035 VSS.n10970 VSS.t3323 8.06917
R2036 VSS.n10956 VSS.t2228 8.06917
R2037 VSS.n10956 VSS.t2961 8.06917
R2038 VSS.n10957 VSS.t2547 8.06917
R2039 VSS.n10957 VSS.t3257 8.06917
R2040 VSS.n10965 VSS.t1401 8.06917
R2041 VSS.n10965 VSS.t2076 8.06917
R2042 VSS.n10966 VSS.t929 8.06917
R2043 VSS.n10966 VSS.t1697 8.06917
R2044 VSS.n10970 VSS.t2324 8.06917
R2045 VSS.n10970 VSS.t3071 8.06917
R2046 VSS.n722 VSS.t1317 8.06917
R2047 VSS.n722 VSS.t2348 8.06917
R2048 VSS.n721 VSS.t1647 8.06917
R2049 VSS.n721 VSS.t2701 8.06917
R2050 VSS.n715 VSS.t3523 8.06917
R2051 VSS.n715 VSS.t1522 8.06917
R2052 VSS.n714 VSS.t3133 8.06917
R2053 VSS.n714 VSS.t1068 8.06917
R2054 VSS.n711 VSS.t1429 8.06917
R2055 VSS.n711 VSS.t2454 8.06917
R2056 VSS.n722 VSS.t3621 8.06917
R2057 VSS.n722 VSS.t1257 8.06917
R2058 VSS.n721 VSS.t830 8.06917
R2059 VSS.n721 VSS.t1593 8.06917
R2060 VSS.n715 VSS.t2765 8.06917
R2061 VSS.n715 VSS.t3447 8.06917
R2062 VSS.n714 VSS.t2340 8.06917
R2063 VSS.n714 VSS.t3101 8.06917
R2064 VSS.n711 VSS.t562 8.06917
R2065 VSS.n711 VSS.t1370 8.06917
R2066 VSS.n1169 VSS.t2903 8.06917
R2067 VSS.n1169 VSS.t832 8.06917
R2068 VSS.n1170 VSS.t3205 8.06917
R2069 VSS.n1170 VSS.t1178 8.06917
R2070 VSS.n1190 VSS.t2023 8.06917
R2071 VSS.n1190 VSS.t3113 8.06917
R2072 VSS.n1191 VSS.t1641 8.06917
R2073 VSS.n1191 VSS.t2697 8.06917
R2074 VSS.n1195 VSS.t3009 8.06917
R2075 VSS.n1195 VSS.t933 8.06917
R2076 VSS.n1169 VSS.t1346 8.06917
R2077 VSS.n1169 VSS.t3325 8.06917
R2078 VSS.n1170 VSS.t1675 8.06917
R2079 VSS.n1170 VSS.t502 8.06917
R2080 VSS.n1190 VSS.t3547 8.06917
R2081 VSS.n1190 VSS.t2476 8.06917
R2082 VSS.n1191 VSS.t3155 8.06917
R2083 VSS.n1191 VSS.t2090 8.06917
R2084 VSS.n1195 VSS.t1455 8.06917
R2085 VSS.n1195 VSS.t3437 8.06917
R2086 VSS.n9147 VSS.t3015 8.06917
R2087 VSS.n9147 VSS.t538 8.06917
R2088 VSS.n9151 VSS.t2206 8.06917
R2089 VSS.n9151 VSS.t2921 8.06917
R2090 VSS.n9152 VSS.t2503 8.06917
R2091 VSS.n9152 VSS.t3217 8.06917
R2092 VSS.n9160 VSS.t1351 8.06917
R2093 VSS.n9160 VSS.t2033 8.06917
R2094 VSS.n9161 VSS.t895 8.06917
R2095 VSS.n9161 VSS.t1655 8.06917
R2096 VSS.n9165 VSS.t2284 8.06917
R2097 VSS.n9165 VSS.t3025 8.06917
R2098 VSS.n9147 VSS.t1453 8.06917
R2099 VSS.n9147 VSS.t2146 8.06917
R2100 VSS.n9151 VSS.t549 8.06917
R2101 VSS.n9151 VSS.t1365 8.06917
R2102 VSS.n9152 VSS.t915 8.06917
R2103 VSS.n9152 VSS.t1683 8.06917
R2104 VSS.n9160 VSS.t2871 8.06917
R2105 VSS.n9160 VSS.t3557 8.06917
R2106 VSS.n9161 VSS.t2442 8.06917
R2107 VSS.n9161 VSS.t3161 8.06917
R2108 VSS.n9165 VSS.t678 8.06917
R2109 VSS.n9165 VSS.t1463 8.06917
R2110 VSS.t2042 VSS.t301 7.5006
R2111 VSS.t2481 VSS.t305 7.5006
R2112 VSS.t302 VSS.t1242 7.5006
R2113 VSS.n572 VSS.t115 7.42489
R2114 VSS.t58 VSS.n565 7.41222
R2115 VSS.n9890 VSS.t328 7.25283
R2116 VSS.n11391 VSS.n60 7.08065
R2117 VSS.n10308 VSS.t164 6.72766
R2118 VSS.t282 VSS.t545 6.61526
R2119 VSS.n10760 VSS.t2923 6.60917
R2120 VSS.n10760 VSS.t1599 6.60917
R2121 VSS.n10760 VSS.t3347 6.60917
R2122 VSS.n10760 VSS.t2003 6.60917
R2123 VSS.n10760 VSS.t3041 6.60917
R2124 VSS.n10738 VSS.t568 6.60917
R2125 VSS.n10764 VSS.t664 6.60917
R2126 VSS.n10740 VSS.t723 6.60917
R2127 VSS.n10759 VSS.t794 6.60917
R2128 VSS.n10774 VSS.t3153 6.60917
R2129 VSS.n10771 VSS.t1826 6.60917
R2130 VSS.n10856 VSS.t3603 6.60917
R2131 VSS.n10854 VSS.t2232 6.60917
R2132 VSS.n10743 VSS.t3243 6.60917
R2133 VSS.n10388 VSS.t196 6.53862
R2134 VSS.n9347 VSS.n9346 6.4661
R2135 VSS.n9422 VSS.n1383 6.4661
R2136 VSS.t101 VSS.t284 6.21678
R2137 VSS.t1249 VSS.t390 5.81954
R2138 VSS.t105 VSS.t495 5.8183
R2139 VSS.t106 VSS.t800 5.8183
R2140 VSS.n10739 VSS.t190 5.49372
R2141 VSS.n10306 VSS.t276 5.47432
R2142 VSS.t411 VSS.t250 5.34013
R2143 VSS.n10032 VSS.n566 5.34013
R2144 VSS.n10301 VSS.n10300 5.31981
R2145 VSS.n10392 VSS.t25 5.28484
R2146 VSS.n10397 VSS.t125 5.28484
R2147 VSS.n10391 VSS.t157 5.28484
R2148 VSS.n10305 VSS.n10292 5.26136
R2149 VSS.n10761 VSS.t2924 5.2505
R2150 VSS.t2924 VSS.n241 5.2505
R2151 VSS.n10761 VSS.t1601 5.2505
R2152 VSS.t1601 VSS.n241 5.2505
R2153 VSS.n10761 VSS.t3348 5.2505
R2154 VSS.t3348 VSS.n241 5.2505
R2155 VSS.n10761 VSS.t2004 5.2505
R2156 VSS.t2004 VSS.n241 5.2505
R2157 VSS.n10761 VSS.t3042 5.2505
R2158 VSS.t3042 VSS.n241 5.2505
R2159 VSS.n10768 VSS.t569 5.2505
R2160 VSS.n10763 VSS.t665 5.2505
R2161 VSS.t795 VSS.n10739 5.2505
R2162 VSS.t724 VSS.n10755 5.2505
R2163 VSS.n10410 VSS.n10409 5.16888
R2164 VSS.n10374 VSS.n10373 5.15456
R2165 VSS.n10680 VSS.n10679 5.09675
R2166 VSS.t614 VSS.t511 4.94165
R2167 VSS.n10066 VSS.t542 4.78226
R2168 VSS.n10626 VSS.n10623 4.63106
R2169 VSS.n10617 VSS.n10614 4.63106
R2170 VSS.n10381 VSS.n10378 4.63106
R2171 VSS.n10302 VSS.n10301 4.61712
R2172 VSS.n10684 VSS.n10683 4.61712
R2173 VSS.n10806 VSS.n10802 4.61585
R2174 VSS.n10800 VSS.n10796 4.61585
R2175 VSS.n9196 VSS.n9195 4.61205
R2176 VSS.n9191 VSS.n9190 4.61205
R2177 VSS.n9332 VSS.n9331 4.61205
R2178 VSS.n9327 VSS.n9326 4.61205
R2179 VSS.n170 VSS.n169 4.61205
R2180 VSS.n165 VSS.n164 4.61205
R2181 VSS.n9578 VSS.n9577 4.61205
R2182 VSS.n9573 VSS.n9572 4.61205
R2183 VSS.n193 VSS.n192 4.61205
R2184 VSS.n198 VSS.n197 4.61205
R2185 VSS.n471 VSS.n470 4.61205
R2186 VSS.n476 VSS.n475 4.61205
R2187 VSS.n9029 VSS.n9028 4.61205
R2188 VSS.n9024 VSS.n9023 4.61205
R2189 VSS.n264 VSS.n263 4.61205
R2190 VSS.n269 VSS.n268 4.61205
R2191 VSS.n336 VSS.n335 4.61205
R2192 VSS.n341 VSS.n340 4.61205
R2193 VSS.n408 VSS.n407 4.61205
R2194 VSS.n413 VSS.n412 4.61205
R2195 VSS.n10630 VSS.n10628 4.61078
R2196 VSS.n10621 VSS.n10619 4.61078
R2197 VSS.n10385 VSS.n10383 4.61078
R2198 VSS.n10376 VSS.n10374 4.61078
R2199 VSS.n10682 VSS.n10681 4.61078
R2200 VSS.n10631 VSS.n10630 4.60825
R2201 VSS.n10622 VSS.n10621 4.60825
R2202 VSS.n10386 VSS.n10385 4.60825
R2203 VSS.n10377 VSS.n10376 4.60825
R2204 VSS.n10681 VSS.n10680 4.60825
R2205 VSS.n10309 VSS.n10306 4.60439
R2206 VSS.n10807 VSS.n10806 4.60318
R2207 VSS.n10801 VSS.n10800 4.60318
R2208 VSS.n10303 VSS.n10302 4.60191
R2209 VSS.n10685 VSS.n10684 4.60191
R2210 VSS.n10627 VSS.n10626 4.58796
R2211 VSS.n10618 VSS.n10617 4.58796
R2212 VSS.n10382 VSS.n10381 4.58796
R2213 VSS.n9194 VSS.n9193 4.5005
R2214 VSS.n9189 VSS.n9188 4.5005
R2215 VSS.n9330 VSS.n9329 4.5005
R2216 VSS.n9325 VSS.n9324 4.5005
R2217 VSS.n168 VSS.n167 4.5005
R2218 VSS.n163 VSS.n162 4.5005
R2219 VSS.n9576 VSS.n9575 4.5005
R2220 VSS.n9571 VSS.n9570 4.5005
R2221 VSS.n191 VSS.n190 4.5005
R2222 VSS.n196 VSS.n195 4.5005
R2223 VSS.n469 VSS.n468 4.5005
R2224 VSS.n474 VSS.n473 4.5005
R2225 VSS.n10798 VSS.n10795 4.5005
R2226 VSS.n10804 VSS.n10794 4.5005
R2227 VSS.n9027 VSS.n9026 4.5005
R2228 VSS.n9022 VSS.n9021 4.5005
R2229 VSS.n9019 VSS.n9018 4.5005
R2230 VSS.n9019 VSS.n1560 4.5005
R2231 VSS.n9034 VSS.n9033 4.5005
R2232 VSS.n9033 VSS.n9032 4.5005
R2233 VSS.n262 VSS.n261 4.5005
R2234 VSS.n267 VSS.n266 4.5005
R2235 VSS.n334 VSS.n333 4.5005
R2236 VSS.n339 VSS.n338 4.5005
R2237 VSS.n406 VSS.n405 4.5005
R2238 VSS.n411 VSS.n410 4.5005
R2239 VSS.n10144 VSS.n10143 4.5005
R2240 VSS.n10143 VSS.n403 4.5005
R2241 VSS.n10146 VSS.n10145 4.5005
R2242 VSS.n10147 VSS.n10146 4.5005
R2243 VSS.n10204 VSS.n10203 4.5005
R2244 VSS.n10203 VSS.n331 4.5005
R2245 VSS.n10206 VSS.n10205 4.5005
R2246 VSS.n10207 VSS.n10206 4.5005
R2247 VSS.n10264 VSS.n10263 4.5005
R2248 VSS.n10263 VSS.n259 4.5005
R2249 VSS.n10266 VSS.n10265 4.5005
R2250 VSS.n10267 VSS.n10266 4.5005
R2251 VSS.n10571 VSS.n10570 4.5005
R2252 VSS.n10570 VSS.n10569 4.5005
R2253 VSS.n10569 VSS.n10556 4.5005
R2254 VSS.n10563 VSS.n10556 4.5005
R2255 VSS.n10572 VSS.n10563 4.5005
R2256 VSS.n10572 VSS.n10557 4.5005
R2257 VSS.n10572 VSS.n10571 4.5005
R2258 VSS.n10375 VSS.n10372 4.5005
R2259 VSS.n10380 VSS.n10371 4.5005
R2260 VSS.n10384 VSS.n10370 4.5005
R2261 VSS.n10616 VSS.n10369 4.5005
R2262 VSS.n10620 VSS.n10368 4.5005
R2263 VSS.n10625 VSS.n10367 4.5005
R2264 VSS.n10629 VSS.n10366 4.5005
R2265 VSS.n10294 VSS.n10293 4.5005
R2266 VSS.n10297 VSS.n10295 4.5005
R2267 VSS.n10299 VSS.n10298 4.5005
R2268 VSS.n10913 VSS.n226 4.5005
R2269 VSS.n10913 VSS.n229 4.5005
R2270 VSS.n10913 VSS.n225 4.5005
R2271 VSS.n10913 VSS.n10912 4.5005
R2272 VSS.n229 VSS.n223 4.5005
R2273 VSS.n225 VSS.n223 4.5005
R2274 VSS.n10912 VSS.n223 4.5005
R2275 VSS.n11338 VSS.n108 4.5005
R2276 VSS.n11337 VSS.n103 4.5005
R2277 VSS.n11338 VSS.n106 4.5005
R2278 VSS.n11338 VSS.n109 4.5005
R2279 VSS.n11338 VSS.n11337 4.5005
R2280 VSS.n11337 VSS.n11336 4.5005
R2281 VSS.n11336 VSS.n109 4.5005
R2282 VSS.n11336 VSS.n106 4.5005
R2283 VSS.n11336 VSS.n108 4.5005
R2284 VSS.n483 VSS.n482 4.5005
R2285 VSS.n482 VSS.n466 4.5005
R2286 VSS.n480 VSS.n463 4.5005
R2287 VSS.n480 VSS.n479 4.5005
R2288 VSS.n11141 VSS.n11140 4.5005
R2289 VSS.n11140 VSS.n188 4.5005
R2290 VSS.n11143 VSS.n11142 4.5005
R2291 VSS.n11144 VSS.n11143 4.5005
R2292 VSS.n11432 VSS.n11431 4.5005
R2293 VSS.n11431 VSS.n11430 4.5005
R2294 VSS.n11429 VSS.n32 4.5005
R2295 VSS.n11430 VSS.n11429 4.5005
R2296 VSS.n11433 VSS.n32 4.5005
R2297 VSS.n11433 VSS.n30 4.5005
R2298 VSS.n11433 VSS.n11432 4.5005
R2299 VSS.n11400 VSS.n56 4.5005
R2300 VSS.n11400 VSS.n11399 4.5005
R2301 VSS.n11396 VSS.n57 4.5005
R2302 VSS.n57 VSS.n56 4.5005
R2303 VSS.n11399 VSS.n57 4.5005
R2304 VSS.n11398 VSS.n11396 4.5005
R2305 VSS.n11399 VSS.n11398 4.5005
R2306 VSS.n11384 VSS.n62 4.5005
R2307 VSS.n11387 VSS.n11383 4.5005
R2308 VSS.n11383 VSS.n78 4.5005
R2309 VSS.n11388 VSS.n78 4.5005
R2310 VSS.n11386 VSS.n78 4.5005
R2311 VSS.n11388 VSS.n11387 4.5005
R2312 VSS.n11387 VSS.n62 4.5005
R2313 VSS.n11387 VSS.n83 4.5005
R2314 VSS.n11387 VSS.n11386 4.5005
R2315 VSS.n9582 VSS.n9568 4.5005
R2316 VSS.n9583 VSS.n9582 4.5005
R2317 VSS.n9586 VSS.n9585 4.5005
R2318 VSS.n9585 VSS.n9584 4.5005
R2319 VSS.n160 VSS.n159 4.5005
R2320 VSS.n160 VSS.n157 4.5005
R2321 VSS.n176 VSS.n175 4.5005
R2322 VSS.n175 VSS.n174 4.5005
R2323 VSS.n9335 VSS.n9322 4.5005
R2324 VSS.n9336 VSS.n9335 4.5005
R2325 VSS.n9339 VSS.n9338 4.5005
R2326 VSS.n9338 VSS.n9337 4.5005
R2327 VSS.n9186 VSS.n9185 4.5005
R2328 VSS.n9186 VSS.n1522 4.5005
R2329 VSS.n9201 VSS.n9200 4.5005
R2330 VSS.n9200 VSS.n9199 4.5005
R2331 VSS.n11310 VSS.n11309 4.5005
R2332 VSS.n11305 VSS.n122 4.5005
R2333 VSS.n11305 VSS.n124 4.5005
R2334 VSS.n11309 VSS.n11308 4.5005
R2335 VSS.n11308 VSS.n11307 4.5005
R2336 VSS.n11308 VSS.n122 4.5005
R2337 VSS.n11308 VSS.n124 4.5005
R2338 VSS.n10732 VSS.n10731 4.5005
R2339 VSS.n10728 VSS.n10707 4.5005
R2340 VSS.n10729 VSS.n10728 4.5005
R2341 VSS.n10731 VSS.n10730 4.5005
R2342 VSS.n10730 VSS.n10704 4.5005
R2343 VSS.n10730 VSS.n10707 4.5005
R2344 VSS.n10730 VSS.n10729 4.5005
R2345 VSS.n10322 VSS.t195 4.41563
R2346 VSS.n10331 VSS.t36 4.41563
R2347 VSS.n10320 VSS.t140 4.41563
R2348 VSS.n10310 VSS.t139 4.41563
R2349 VSS.t1800 VSS.t638 4.2678
R2350 VSS.n10404 VSS.t8 4.22616
R2351 VSS.n10402 VSS.t170 4.22616
R2352 VSS.n10308 VSS.n10307 4.21432
R2353 VSS.n10305 VSS.n10304 4.21432
R2354 VSS.n9884 VSS.n9883 4.21138
R2355 VSS.n9881 VSS.n9880 4.21138
R2356 VSS.n9879 VSS.n9878 4.21138
R2357 VSS.n9518 VSS.n642 4.21138
R2358 VSS.n9896 VSS.n9895 4.21138
R2359 VSS.n9914 VSS.n9907 4.21138
R2360 VSS.n9919 VSS.n9918 4.21138
R2361 VSS.n678 VSS.n648 4.21074
R2362 VSS.n9859 VSS.n9854 4.21074
R2363 VSS.n9873 VSS.n9872 4.21074
R2364 VSS.n1255 VSS.n1254 4.21074
R2365 VSS.n9902 VSS.n628 4.21074
R2366 VSS.n627 VSS.n584 4.21074
R2367 VSS.n9926 VSS.n9925 4.21074
R2368 VSS.n11450 VSS.n19 4.21074
R2369 VSS.n11445 VSS.n22 4.21074
R2370 VSS.n11417 VSS.n44 4.21074
R2371 VSS.n11412 VSS.n47 4.21074
R2372 VSS.n9617 VSS.n650 4.21074
R2373 VSS.n9610 VSS.n822 4.21074
R2374 VSS.n9616 VSS.n811 4.21074
R2375 VSS.n9611 VSS.n814 4.21074
R2376 VSS.n9517 VSS.n1327 4.21074
R2377 VSS.n9512 VSS.n9511 4.21074
R2378 VSS.n9611 VSS.n9610 4.19858
R2379 VSS.n822 VSS.n648 4.19794
R2380 VSS.n9884 VSS.n650 4.19794
R2381 VSS.n679 VSS.n678 4.19794
R2382 VSS.n9883 VSS.n9882 4.19794
R2383 VSS.n9872 VSS.n9859 4.19794
R2384 VSS.n9880 VSS.n9879 4.19794
R2385 VSS.n9512 VSS.n1255 4.19794
R2386 VSS.n9518 VSS.n9517 4.19794
R2387 VSS.n1254 VSS.n628 4.19794
R2388 VSS.n9895 VSS.n642 4.19794
R2389 VSS.n9903 VSS.n9902 4.19794
R2390 VSS.n9896 VSS.n621 4.19794
R2391 VSS.n9926 VSS.n584 4.19794
R2392 VSS.n9918 VSS.n9914 4.19794
R2393 VSS.n9925 VSS.n22 4.19794
R2394 VSS.n9919 VSS.n19 4.19794
R2395 VSS.n9873 VSS.n47 4.19794
R2396 VSS.n9878 VSS.n44 4.19794
R2397 VSS.n9617 VSS.n9616 4.19794
R2398 VSS.n11445 VSS.n11444 4.19794
R2399 VSS.n11451 VSS.n11450 4.19794
R2400 VSS.n11412 VSS.n11411 4.19794
R2401 VSS.n11418 VSS.n11417 4.19794
R2402 VSS.n9192 VSS.t449 4.16335
R2403 VSS.n9187 VSS.t453 4.16335
R2404 VSS.n9328 VSS.t394 4.16335
R2405 VSS.n9323 VSS.t388 4.16335
R2406 VSS.n166 VSS.t378 4.16335
R2407 VSS.n161 VSS.t373 4.16335
R2408 VSS.n9574 VSS.t322 4.16335
R2409 VSS.n9569 VSS.t315 4.16335
R2410 VSS.n9025 VSS.t419 4.16335
R2411 VSS.n9020 VSS.t421 4.16335
R2412 VSS.n189 VSS.t179 4.16278
R2413 VSS.n194 VSS.t161 4.16278
R2414 VSS.n467 VSS.t407 4.16278
R2415 VSS.n472 VSS.t402 4.16278
R2416 VSS.n260 VSS.t293 4.16278
R2417 VSS.n265 VSS.t296 4.16278
R2418 VSS.n332 VSS.t3644 4.16278
R2419 VSS.n337 VSS.t3648 4.16278
R2420 VSS.n404 VSS.t338 4.16278
R2421 VSS.n409 VSS.t340 4.16278
R2422 VSS.n9195 VSS.t452 4.16103
R2423 VSS.n9190 VSS.t455 4.16103
R2424 VSS.n9331 VSS.t392 4.16103
R2425 VSS.n9326 VSS.t395 4.16103
R2426 VSS.n169 VSS.t372 4.16103
R2427 VSS.n164 VSS.t375 4.16103
R2428 VSS.n9577 VSS.t3639 4.16103
R2429 VSS.n9572 VSS.t317 4.16103
R2430 VSS.n9028 VSS.t420 4.16103
R2431 VSS.n9023 VSS.t422 4.16103
R2432 VSS.n192 VSS.t178 4.15984
R2433 VSS.n197 VSS.t172 4.15984
R2434 VSS.n470 VSS.t404 4.15984
R2435 VSS.n475 VSS.t408 4.15984
R2436 VSS.n263 VSS.t289 4.15984
R2437 VSS.n268 VSS.t294 4.15984
R2438 VSS.n335 VSS.t3645 4.15984
R2439 VSS.n340 VSS.t3649 4.15984
R2440 VSS.n407 VSS.t343 4.15984
R2441 VSS.n412 VSS.t345 4.15984
R2442 VSS.n10565 VSS.n128 4.1417
R2443 VSS.t252 VSS.n434 4.06499
R2444 VSS.n1346 VSS.t1484 4.03583
R2445 VSS.n1371 VSS.t2172 4.03583
R2446 VSS.n1348 VSS.t1767 4.03583
R2447 VSS.n1365 VSS.t1000 4.03583
R2448 VSS.n1351 VSS.t2659 4.03583
R2449 VSS.n1359 VSS.t3331 4.03583
R2450 VSS.n1354 VSS.t2629 4.03583
R2451 VSS.n803 VSS.t605 4.03583
R2452 VSS.n802 VSS.t2693 4.03583
R2453 VSS.n801 VSS.t3433 4.03583
R2454 VSS.n798 VSS.t996 4.03583
R2455 VSS.n800 VSS.t3085 4.03583
R2456 VSS.n9636 VSS.t2635 4.03583
R2457 VSS.n9756 VSS.t522 4.03583
R2458 VSS.n9638 VSS.t2619 4.03583
R2459 VSS.n9662 VSS.t589 4.03583
R2460 VSS.n9663 VSS.t2661 4.03583
R2461 VSS.n9746 VSS.t1957 4.03583
R2462 VSS.n9665 VSS.t3569 4.03583
R2463 VSS.n9740 VSS.t1192 4.03583
R2464 VSS.n9668 VSS.t3171 4.03583
R2465 VSS.n9734 VSS.t2120 4.03583
R2466 VSS.n9670 VSS.t2893 4.03583
R2467 VSS.n9718 VSS.t879 4.03583
R2468 VSS.n9719 VSS.t3253 4.03583
R2469 VSS.n9724 VSS.t853 4.03583
R2470 VSS.n569 VSS.t3553 4.03583
R2471 VSS.n571 VSS.t2863 4.03583
R2472 VSS.n574 VSS.t3159 4.03583
R2473 VSS.n10021 VSS.t2098 4.03583
R2474 VSS.n577 VSS.t1384 4.03583
R2475 VSS.n9935 VSS.t2468 4.03583
R2476 VSS.n9936 VSS.t1441 4.03583
R2477 VSS.n10009 VSS.t2124 4.03583
R2478 VSS.n9938 VSS.t976 4.03583
R2479 VSS.n10003 VSS.t1804 4.03583
R2480 VSS.n9940 VSS.t1397 4.03583
R2481 VSS.n9997 VSS.t2416 4.03583
R2482 VSS.n9942 VSS.t3357 4.03583
R2483 VSS.n9967 VSS.t1451 4.03583
R2484 VSS.n9968 VSS.t3395 4.03583
R2485 VSS.n9987 VSS.t2729 4.03583
R2486 VSS.n9970 VSS.t2302 4.03583
R2487 VSS.n9981 VSS.t3035 4.03583
R2488 VSS.n9972 VSS.t1911 4.03583
R2489 VSS.n9975 VSS.t810 4.03583
R2490 VSS.n1346 VSS.t3333 4.03583
R2491 VSS.n1371 VSS.t1629 4.03583
R2492 VSS.n1348 VSS.t2689 4.03583
R2493 VSS.n1365 VSS.t2591 4.03583
R2494 VSS.n1351 VSS.t1388 4.03583
R2495 VSS.n1359 VSS.t2703 4.03583
R2496 VSS.n1354 VSS.t1174 4.03583
R2497 VSS.n803 VSS.t2326 4.03583
R2498 VSS.n802 VSS.t1891 4.03583
R2499 VSS.n801 VSS.t1064 4.03583
R2500 VSS.n798 VSS.t2236 4.03583
R2501 VSS.n800 VSS.t3201 4.03583
R2502 VSS.n9636 VSS.t1200 4.03583
R2503 VSS.n9756 VSS.t1496 4.03583
R2504 VSS.n9638 VSS.t986 4.03583
R2505 VSS.n9662 VSS.t2182 4.03583
R2506 VSS.n9663 VSS.t1729 4.03583
R2507 VSS.n9746 VSS.t1661 4.03583
R2508 VSS.n9665 VSS.t3479 4.03583
R2509 VSS.n9740 VSS.t1739 4.03583
R2510 VSS.n9668 VSS.t2521 4.03583
R2511 VSS.n9734 VSS.t3483 4.03583
R2512 VSS.n9670 VSS.t1279 4.03583
R2513 VSS.n9718 VSS.t2420 4.03583
R2514 VSS.n9719 VSS.t905 4.03583
R2515 VSS.n9724 VSS.t2248 4.03583
R2516 VSS.n569 VSS.t3301 4.03583
R2517 VSS.n571 VSS.t3235 4.03583
R2518 VSS.n574 VSS.t2350 4.03583
R2519 VSS.n10021 VSS.t3303 4.03583
R2520 VSS.n577 VSS.t1847 4.03583
R2521 VSS.n9935 VSS.t2997 4.03583
R2522 VSS.n9936 VSS.t2523 4.03583
R2523 VSS.n10009 VSS.t732 4.03583
R2524 VSS.n9938 VSS.t1589 4.03583
R2525 VSS.n10003 VSS.t740 4.03583
R2526 VSS.n9940 VSS.t1857 4.03583
R2527 VSS.n9997 VSS.t2126 4.03583
R2528 VSS.n9942 VSS.t2430 4.03583
R2529 VSS.n9967 VSS.t3577 4.03583
R2530 VSS.n9968 VSS.t3151 4.03583
R2531 VSS.n9987 VSS.t3097 4.03583
R2532 VSS.n9970 VSS.t1027 4.03583
R2533 VSS.n9981 VSS.t2362 4.03583
R2534 VSS.n9972 VSS.t3177 4.03583
R2535 VSS.n9975 VSS.t1034 4.03583
R2536 VSS.n1316 VSS.t2985 4.03583
R2537 VSS.n1312 VSS.t603 4.03583
R2538 VSS.n1307 VSS.t2965 4.03583
R2539 VSS.n1303 VSS.t711 4.03583
R2540 VSS.n443 VSS.t1783 4.03583
R2541 VSS.n447 VSS.t1853 4.03583
R2542 VSS.n449 VSS.t1005 4.03583
R2543 VSS.n453 VSS.t1845 4.03583
R2544 VSS.n10099 VSS.t2643 4.03583
R2545 VSS.n461 VSS.t2665 4.03583
R2546 VSS.n460 VSS.t2549 4.03583
R2547 VSS.n485 VSS.t2356 4.03583
R2548 VSS.n488 VSS.t2601 4.03583
R2549 VSS.n492 VSS.t3475 4.03583
R2550 VSS.n10079 VSS.t3431 4.03583
R2551 VSS.n10075 VSS.t3457 4.03583
R2552 VSS.n501 VSS.t1204 4.03583
R2553 VSS.n519 VSS.t1233 4.03583
R2554 VSS.n522 VSS.t2234 4.03583
R2555 VSS.n528 VSS.t2316 4.03583
R2556 VSS.n515 VSS.t1538 4.03583
R2557 VSS.n539 VSS.t2366 4.03583
R2558 VSS.n541 VSS.t2605 4.03583
R2559 VSS.n545 VSS.t2278 4.03583
R2560 VSS.n551 VSS.t3115 4.03583
R2561 VSS.n554 VSS.t770 4.03583
R2562 VSS.n556 VSS.t3111 4.03583
R2563 VSS.n559 VSS.t844 4.03583
R2564 VSS.n10894 VSS.t1905 4.03583
R2565 VSS.n10890 VSS.t903 4.03583
R2566 VSS.n10876 VSS.t1166 4.03583
R2567 VSS.n10879 VSS.t1969 4.03583
R2568 VSS.n187 VSS.t2799 4.03583
R2569 VSS.n11138 VSS.t2815 4.03583
R2570 VSS.n204 VSS.t2001 4.03583
R2571 VSS.n11021 VSS.t2867 4.03583
R2572 VSS.n11024 VSS.t2743 4.03583
R2573 VSS.n11029 VSS.t3619 4.03583
R2574 VSS.n11031 VSS.t3579 4.03583
R2575 VSS.n11035 VSS.t2825 4.03583
R2576 VSS.n11114 VSS.t3627 4.03583
R2577 VSS.n11055 VSS.t461 4.03583
R2578 VSS.n11057 VSS.t1597 4.03583
R2579 VSS.n11082 VSS.t2450 4.03583
R2580 VSS.n11080 VSS.t1669 4.03583
R2581 VSS.n11088 VSS.t2483 4.03583
R2582 VSS.n11090 VSS.t2749 4.03583
R2583 VSS.n10 VSS.t1731 4.03583
R2584 VSS.n1418 VSS.t2312 4.03583
R2585 VSS.n1420 VSS.t1616 4.03583
R2586 VSS.n1466 VSS.t2286 4.03583
R2587 VSS.n1462 VSS.t1887 4.03583
R2588 VSS.n1427 VSS.t1168 4.03583
R2589 VSS.n1429 VSS.t2813 4.03583
R2590 VSS.n1439 VSS.t3495 4.03583
R2591 VSS.n1443 VSS.t2789 4.03583
R2592 VSS.n829 VSS.t774 4.03583
R2593 VSS.n9589 VSS.t2839 4.03583
R2594 VSS.n9588 VSS.t3587 4.03583
R2595 VSS.n9770 VSS.t1155 4.03583
R2596 VSS.n9776 VSS.t3187 4.03583
R2597 VSS.n9782 VSS.t2793 4.03583
R2598 VSS.n790 VSS.t715 4.03583
R2599 VSS.n787 VSS.t2761 4.03583
R2600 VSS.n9796 VSS.t755 4.03583
R2601 VSS.n772 VSS.t2817 4.03583
R2602 VSS.n9806 VSS.t2088 4.03583
R2603 VSS.n770 VSS.t552 4.03583
R2604 VSS.n9817 VSS.t1361 4.03583
R2605 VSS.n765 VSS.t3291 4.03583
R2606 VSS.n9829 VSS.t2256 4.03583
R2607 VSS.n763 VSS.t3031 4.03583
R2608 VSS.n697 VSS.t1017 4.03583
R2609 VSS.n700 VSS.t3373 4.03583
R2610 VSS.n702 VSS.t992 4.03583
R2611 VSS.n706 VSS.t524 4.03583
R2612 VSS.n726 VSS.t3001 4.03583
R2613 VSS.n728 VSS.t3281 4.03583
R2614 VSS.n740 VSS.t2230 4.03583
R2615 VSS.n736 VSS.t1528 4.03583
R2616 VSS.n158 VSS.t2625 4.03583
R2617 VSS.n11162 VSS.t1571 4.03583
R2618 VSS.n155 VSS.t2262 4.03583
R2619 VSS.n154 VSS.t1122 4.03583
R2620 VSS.n11172 VSS.t1937 4.03583
R2621 VSS.n11176 VSS.t1532 4.03583
R2622 VSS.n11178 VSS.t2551 4.03583
R2623 VSS.n11182 VSS.t3527 4.03583
R2624 VSS.n11258 VSS.t1581 4.03583
R2625 VSS.n11199 VSS.t3565 4.03583
R2626 VSS.n11201 VSS.t2877 4.03583
R2627 VSS.n11227 VSS.t2444 4.03583
R2628 VSS.n11225 VSS.t3157 4.03583
R2629 VSS.n11232 VSS.t2031 4.03583
R2630 VSS.n11234 VSS.t956 4.03583
R2631 VSS.n10394 VSS.n10393 4.02484
R2632 VSS.n10396 VSS.n10395 4.02484
R2633 VSS.n10390 VSS.n10389 4.02484
R2634 VSS.n10388 VSS.n10387 4.02484
R2635 VSS.n10404 VSS.t130 4.02247
R2636 VSS.n10402 VSS.t180 4.02247
R2637 VSS.n10299 VSS.t14 4.00471
R2638 VSS.n10294 VSS.t10 4.00471
R2639 VSS.n10118 VSS.n434 3.9853
R2640 VSS.n9564 VSS.n833 3.9853
R2641 VSS.n10067 VSS.n506 3.9853
R2642 VSS.n10929 VSS.n218 3.9853
R2643 VSS.n11361 VSS.n93 3.9853
R2644 VSS.n11468 VSS.n6 3.9853
R2645 VSS.n9197 VSS.n9191 3.98482
R2646 VSS.n9333 VSS.n9327 3.98482
R2647 VSS.n171 VSS.n165 3.98482
R2648 VSS.n9579 VSS.n9573 3.98482
R2649 VSS.n199 VSS.n193 3.98482
R2650 VSS.n477 VSS.n471 3.98482
R2651 VSS.n9030 VSS.n9024 3.98482
R2652 VSS.n270 VSS.n264 3.98482
R2653 VSS.n342 VSS.n336 3.98482
R2654 VSS.n414 VSS.n408 3.98482
R2655 VSS.n10405 VSS.n10365 3.96014
R2656 VSS.n1454 VSS.t272 3.9481
R2657 VSS.n794 VSS.t263 3.9481
R2658 VSS.n9822 VSS.t271 3.9481
R2659 VSS.n11086 VSS.t114 3.9481
R2660 VSS.n11027 VSS.t107 3.9481
R2661 VSS.n10872 VSS.t111 3.9481
R2662 VSS.n1363 VSS.t268 3.9481
R2663 VSS.n9760 VSS.t265 3.9481
R2664 VSS.n9738 VSS.t273 3.9481
R2665 VSS.n9979 VSS.t118 3.9481
R2666 VSS.n10001 VSS.t109 3.9481
R2667 VSS.n10026 VSS.t119 3.9481
R2668 VSS.n189 VSS.t192 3.93054
R2669 VSS.n194 VSS.t186 3.93054
R2670 VSS.n467 VSS.t409 3.93054
R2671 VSS.n472 VSS.t405 3.93054
R2672 VSS.n260 VSS.t295 3.93054
R2673 VSS.n265 VSS.t291 3.93054
R2674 VSS.n332 VSS.t3646 3.93054
R2675 VSS.n337 VSS.t3642 3.93054
R2676 VSS.n404 VSS.t339 3.93054
R2677 VSS.n409 VSS.t346 3.93054
R2678 VSS.n9192 VSS.t448 3.92996
R2679 VSS.n9187 VSS.t454 3.92996
R2680 VSS.n9328 VSS.t393 3.92996
R2681 VSS.n9323 VSS.t389 3.92996
R2682 VSS.n166 VSS.t377 3.92996
R2683 VSS.n161 VSS.t374 3.92996
R2684 VSS.n9574 VSS.t320 3.92996
R2685 VSS.n9569 VSS.t318 3.92996
R2686 VSS.n9025 VSS.t425 3.92996
R2687 VSS.n9020 VSS.t423 3.92996
R2688 VSS.n9194 VSS.t451 3.92774
R2689 VSS.n9189 VSS.t456 3.92774
R2690 VSS.n9330 VSS.t391 3.92774
R2691 VSS.n9325 VSS.t396 3.92774
R2692 VSS.n168 VSS.t379 3.92774
R2693 VSS.n163 VSS.t376 3.92774
R2694 VSS.n9576 VSS.t321 3.92774
R2695 VSS.n9571 VSS.t319 3.92774
R2696 VSS.n191 VSS.t176 3.92774
R2697 VSS.n196 VSS.t185 3.92774
R2698 VSS.n469 VSS.t406 3.92774
R2699 VSS.n474 VSS.t403 3.92774
R2700 VSS.n9027 VSS.t417 3.92774
R2701 VSS.n9022 VSS.t424 3.92774
R2702 VSS.n262 VSS.t292 3.92774
R2703 VSS.n267 VSS.t288 3.92774
R2704 VSS.n334 VSS.t3647 3.92774
R2705 VSS.n339 VSS.t3643 3.92774
R2706 VSS.n406 VSS.t344 3.92774
R2707 VSS.n411 VSS.t342 3.92774
R2708 VSS.t54 VSS.n148 3.9056
R2709 VSS.n10322 VSS.t168 3.833
R2710 VSS.n10331 VSS.t121 3.833
R2711 VSS.n10320 VSS.t135 3.833
R2712 VSS.n10310 VSS.t141 3.833
R2713 VSS.n10629 VSS.t42 3.81405
R2714 VSS.n10620 VSS.t39 3.81405
R2715 VSS.n10384 VSS.t193 3.81405
R2716 VSS.n10375 VSS.t137 3.81405
R2717 VSS.n10390 VSS.n10388 3.80578
R2718 VSS.n10396 VSS.n10394 3.80578
R2719 VSS.n10319 VSS.n10315 3.80578
R2720 VSS.n10330 VSS.n10326 3.80578
R2721 VSS.n754 VSS.t108 3.78612
R2722 VSS.n156 VSS.t117 3.78612
R2723 VSS.n11204 VSS.t113 3.78612
R2724 VSS.n527 VSS.t266 3.78612
R2725 VSS.n464 VSS.t270 3.78612
R2726 VSS.n1300 VSS.t267 3.78612
R2727 VSS.n9722 VSS.t116 3.78612
R2728 VSS.n10007 VSS.t110 3.78612
R2729 VSS.n9985 VSS.t112 3.78612
R2730 VSS.n9744 VSS.t264 3.78612
R2731 VSS.n9634 VSS.t269 3.78612
R2732 VSS.n1369 VSS.t261 3.78612
R2733 VSS.n10686 VSS.n10685 3.76738
R2734 VSS.n11301 VSS.t362 3.75339
R2735 VSS.t171 VSS.t566 3.74621
R2736 VSS.n9140 VSS.t355 3.73318
R2737 VSS.n9141 VSS.t357 3.73318
R2738 VSS.n1488 VSS.t369 3.73318
R2739 VSS.n1489 VSS.t371 3.73318
R2740 VSS.n1208 VSS.t152 3.73318
R2741 VSS.n1209 VSS.t279 3.73318
R2742 VSS.n10946 VSS.t3641 3.73318
R2743 VSS.n10947 VSS.t3640 3.73318
R2744 VSS.n10992 VSS.t438 3.73318
R2745 VSS.n10993 VSS.t437 3.73318
R2746 VSS.n8973 VSS.t444 3.73318
R2747 VSS.n8974 VSS.t442 3.73318
R2748 VSS.n978 VSS.t331 3.73318
R2749 VSS.n979 VSS.t334 3.73318
R2750 VSS.n1036 VSS.t359 3.73318
R2751 VSS.n1037 VSS.t361 3.73318
R2752 VSS.n1085 VSS.t347 3.73318
R2753 VSS.n1086 VSS.t397 3.73318
R2754 VSS.n871 VSS.t434 3.73318
R2755 VSS.n872 VSS.t433 3.73318
R2756 VSS.n10601 VSS.t167 3.72778
R2757 VSS.n9140 VSS.t356 3.4916
R2758 VSS.n9141 VSS.t354 3.4916
R2759 VSS.n1488 VSS.t370 3.4916
R2760 VSS.n1489 VSS.t368 3.4916
R2761 VSS.n1208 VSS.t348 3.4916
R2762 VSS.n1209 VSS.t380 3.4916
R2763 VSS.n10946 VSS.t432 3.4916
R2764 VSS.n10947 VSS.t431 3.4916
R2765 VSS.n10992 VSS.t440 3.4916
R2766 VSS.n10993 VSS.t439 3.4916
R2767 VSS.n8973 VSS.t430 3.4916
R2768 VSS.n8974 VSS.t443 3.4916
R2769 VSS.n978 VSS.t333 3.4916
R2770 VSS.n979 VSS.t332 3.4916
R2771 VSS.n1036 VSS.t360 3.4916
R2772 VSS.n1037 VSS.t358 3.4916
R2773 VSS.n1085 VSS.t280 3.4916
R2774 VSS.n1086 VSS.t277 3.4916
R2775 VSS.n871 VSS.t436 3.4916
R2776 VSS.n872 VSS.t435 3.4916
R2777 VSS.t1807 VSS.n10840 3.40963
R2778 VSS.n10638 VSS.t1982 3.37683
R2779 VSS.n11324 VSS.t2217 3.36554
R2780 VSS.n10823 VSS.t1716 3.3605
R2781 VSS.t1716 VSS.n10821 3.3605
R2782 VSS.n10823 VSS.t3486 3.3605
R2783 VSS.t3486 VSS.n10821 3.3605
R2784 VSS.n10841 VSS.t1807 3.3605
R2785 VSS.n10843 VSS.t2796 3.3605
R2786 VSS.t2796 VSS.n10842 3.3605
R2787 VSS.n10712 VSS.t364 3.3605
R2788 VSS.n10713 VSS.t363 3.3605
R2789 VSS.t1435 VSS.n127 3.3605
R2790 VSS.n9205 VSS.t632 3.3605
R2791 VSS.n9183 VSS.t2732 3.3605
R2792 VSS.t3310 VSS.n1523 3.3605
R2793 VSS.n9061 VSS.t2281 3.3605
R2794 VSS.t3516 VSS.n1527 3.3605
R2795 VSS.n1546 VSS.t1517 3.3605
R2796 VSS.n1548 VSS.t1780 3.3605
R2797 VSS.n1552 VSS.t1020 3.3605
R2798 VSS.n9170 VSS.t3108 3.3605
R2799 VSS.n9174 VSS.t2022 3.3605
R2800 VSS.n9136 VSS.t2640 3.3605
R2801 VSS.n9132 VSS.t1611 3.3605
R2802 VSS.n9256 VSS.t867 3.3605
R2803 VSS.n9252 VSS.t2948 3.3605
R2804 VSS.t1718 VSS.n1513 3.3605
R2805 VSS.n9146 VSS.t2403 3.3605
R2806 VSS.n9241 VSS.t1624 3.3605
R2807 VSS.n9245 VSS.t3626 3.3605
R2808 VSS.n9211 VSS.t2391 3.3605
R2809 VSS.n9207 VSS.t3132 3.3605
R2810 VSS.n9314 VSS.t2047 3.3605
R2811 VSS.n9310 VSS.t973 3.3605
R2812 VSS.t1636 VSS.n1505 3.3605
R2813 VSS.n9217 VSS.t2319 3.3605
R2814 VSS.n9292 VSS.t1375 3.3605
R2815 VSS.n9296 VSS.t3350 3.3605
R2816 VSS.n9262 VSS.t885 3.3605
R2817 VSS.n9258 VSS.t1640 3.3605
R2818 VSS.n9354 VSS.t2858 3.3605
R2819 VSS.n9350 VSS.t2143 3.3605
R2820 VSS.t1383 VSS.n1496 3.3605
R2821 VSS.n9268 VSS.t2407 3.3605
R2822 VSS.t3540 VSS.n1478 3.3605
R2823 VSS.n9343 VSS.t2854 3.3605
R2824 VSS.n9320 VSS.t2055 3.3605
R2825 VSS.n9316 VSS.t3138 3.3605
R2826 VSS.n9387 VSS.t2604 3.3605
R2827 VSS.n9383 VSS.t475 3.3605
R2828 VSS.n9380 VSS.t2187 3.3605
R2829 VSS.n9376 VSS.t3220 3.3605
R2830 VSS.n9415 VSS.t1916 3.3605
R2831 VSS.n9419 VSS.t2988 3.3605
R2832 VSS.t1495 VSS.n1396 3.3605
R2833 VSS.n1494 VSS.t2518 3.3605
R2834 VSS.n9534 VSS.t1095 3.3605
R2835 VSS.n9530 VSS.t2185 3.3605
R2836 VSS.t1422 VSS.n1221 3.3605
R2837 VSS.n1402 VSS.t626 3.3605
R2838 VSS.n11236 VSS.t957 3.3605
R2839 VSS.n11242 VSS.t2032 3.3605
R2840 VSS.n11230 VSS.t3158 3.3605
R2841 VSS.n11248 VSS.t2445 3.3605
R2842 VSS.n11203 VSS.t2878 3.3605
R2843 VSS.n11254 VSS.t3566 3.3605
R2844 VSS.n11256 VSS.t1582 3.3605
R2845 VSS.t1582 VSS.n11197 3.3605
R2846 VSS.n11262 VSS.t3528 3.3605
R2847 VSS.t3528 VSS.n11180 3.3605
R2848 VSS.t2552 VSS.n11268 3.3605
R2849 VSS.t1533 VSS.n11174 3.3605
R2850 VSS.t1938 VSS.n11274 3.3605
R2851 VSS.t1123 VSS.n11171 3.3605
R2852 VSS.n11167 VSS.t2263 3.3605
R2853 VSS.n173 VSS.t1572 3.3605
R2854 VSS.n11158 VSS.t2626 3.3605
R2855 VSS.t2626 VSS.n11157 3.3605
R2856 VSS.n734 VSS.t1529 3.3605
R2857 VSS.t1529 VSS.n732 3.3605
R2858 VSS.n730 VSS.t2231 3.3605
R2859 VSS.n745 VSS.t3282 3.3605
R2860 VSS.t3002 VSS.n747 3.3605
R2861 VSS.t525 VSS.n704 3.3605
R2862 VSS.t993 VSS.n755 3.3605
R2863 VSS.t3374 VSS.n696 3.3605
R2864 VSS.t1018 VSS.n761 3.3605
R2865 VSS.n762 VSS.t1018 3.3605
R2866 VSS.n9837 VSS.t3032 3.3605
R2867 VSS.t3032 VSS.n9836 3.3605
R2868 VSS.n9833 VSS.t2257 3.3605
R2869 VSS.n9825 VSS.t3292 3.3605
R2870 VSS.n9821 VSS.t1362 3.3605
R2871 VSS.n9812 VSS.t553 3.3605
R2872 VSS.n9810 VSS.t2089 3.3605
R2873 VSS.n9802 VSS.t2818 3.3605
R2874 VSS.n9799 VSS.t756 3.3605
R2875 VSS.t756 VSS.n9798 3.3605
R2876 VSS.n9792 VSS.t2762 3.3605
R2877 VSS.t2762 VSS.n9791 3.3605
R2878 VSS.n9787 VSS.t716 3.3605
R2879 VSS.n9780 VSS.t2794 3.3605
R2880 VSS.n9774 VSS.t3188 3.3605
R2881 VSS.t1156 VSS.n9772 3.3605
R2882 VSS.n9581 VSS.t3588 3.3605
R2883 VSS.n9595 VSS.t2840 3.3605
R2884 VSS.t775 VSS.n9598 3.3605
R2885 VSS.n9599 VSS.t775 3.3605
R2886 VSS.t2790 VSS.n1445 3.3605
R2887 VSS.n1446 VSS.t2790 3.3605
R2888 VSS.n1441 VSS.t3496 3.3605
R2889 VSS.n1452 VSS.t2814 3.3605
R2890 VSS.n1458 VSS.t1169 3.3605
R2891 VSS.t1888 VSS.n1425 3.3605
R2892 VSS.n1423 VSS.t2287 3.3605
R2893 VSS.n1470 VSS.t1617 3.3605
R2894 VSS.n1472 VSS.t2313 3.3605
R2895 VSS.t2313 VSS.n1403 3.3605
R2896 VSS.t3208 VSS.n11237 3.3605
R2897 VSS.t807 VSS.n11231 3.3605
R2898 VSS.t1462 VSS.n11243 3.3605
R2899 VSS.t3444 VSS.n11228 3.3605
R2900 VSS.t1904 VSS.n11249 3.3605
R2901 VSS.t2970 VSS.n11198 3.3605
R2902 VSS.n11255 VSS.t3196 3.3605
R2903 VSS.n11261 VSS.t2155 3.3605
R2904 VSS.t2770 VSS.n11265 3.3605
R2905 VSS.t3454 VSS.n11177 3.3605
R2906 VSS.t3314 VSS.n11271 3.3605
R2907 VSS.t945 VSS.n152 3.3605
R2908 VSS.n11170 VSS.t3054 3.3605
R2909 VSS.n11163 VSS.t597 3.3605
R2910 VSS.n11161 VSS.t2295 3.3605
R2911 VSS.n11155 VSS.t1256 3.3605
R2912 VSS.n733 VSS.t1874 3.3605
R2913 VSS.n739 VSS.t773 3.3605
R2914 VSS.n742 VSS.t2111 3.3605
R2915 VSS.n747 VSS.t3164 3.3605
R2916 VSS.t1358 VSS.n751 3.3605
R2917 VSS.t2040 VSS.n701 3.3605
R2918 VSS.t3602 VSS.n758 3.3605
R2919 VSS.t1613 VSS.n698 3.3605
R2920 VSS.n9840 VSS.t1868 3.3605
R2921 VSS.n9834 VSS.t1129 3.3605
R2922 VSS.t521 VSS.n764 3.3605
R2923 VSS.t1686 VSS.n9826 3.3605
R2924 VSS.t2139 VSS.n769 3.3605
R2925 VSS.t1059 VSS.n9813 3.3605
R2926 VSS.t2365 VSS.n771 3.3605
R2927 VSS.t3388 VSS.n9803 3.3605
R2928 VSS.t3024 VSS.n773 3.3605
R2929 VSS.t1950 VSS.n9793 3.3605
R2930 VSS.n9790 VSS.t3232 3.3605
R2931 VSS.n9783 VSS.t1215 3.3605
R2932 VSS.n9779 VSS.t2728 3.3605
R2933 VSS.n9771 VSS.t2008 3.3605
R2934 VSS.t2267 VSS.n796 3.3605
R2935 VSS.t1509 VSS.n9590 3.3605
R2936 VSS.n9597 VSS.t1776 3.3605
R2937 VSS.t1012 VSS.n827 3.3605
R2938 VSS.n1444 VSS.t2329 3.3605
R2939 VSS.n1449 VSS.t3364 3.3605
R2940 VSS.n1428 VSS.t1232 3.3605
R2941 VSS.n1461 VSS.t3594 3.3605
R2942 VSS.t1819 VSS.n1463 3.3605
R2943 VSS.t2886 VSS.n1422 3.3605
R2944 VSS.n1419 VSS.t2097 3.3605
R2945 VSS.n1475 VSS.t1418 3.3605
R2946 VSS.n9547 VSS.t1578 3.3605
R2947 VSS.n9543 VSS.t743 3.3605
R2948 VSS.n9540 VSS.t1022 3.3605
R2949 VSS.n9536 VSS.t3392 3.3605
R2950 VSS.n1200 VSS.t1688 3.3605
R2951 VSS.n1204 VSS.t2734 3.3605
R2952 VSS.n1206 VSS.t2293 3.3605
R2953 VSS.n1214 VSS.t1252 3.3605
R2954 VSS.n10936 VSS.t2934 3.3605
R2955 VSS.n10932 VSS.t852 3.3605
R2956 VSS.t1140 VSS.n214 3.3605
R2957 VSS.n1168 VSS.t3532 3.3605
R2958 VSS.n10975 VSS.t1628 3.3605
R2959 VSS.n10979 VSS.t3630 3.3605
R2960 VSS.n10942 VSS.t1150 3.3605
R2961 VSS.n10938 VSS.t3184 3.3605
R2962 VSS.n11368 VSS.t2479 3.3605
R2963 VSS.n11364 VSS.t1470 3.3605
R2964 VSS.t2057 VSS.n90 3.3605
R2965 VSS.n10952 VSS.t2784 3.3605
R2966 VSS.n11381 VSS.t2974 3.3605
R2967 VSS.n11377 VSS.t1908 3.3605
R2968 VSS.n11374 VSS.t2500 3.3605
R2969 VSS.n11370 VSS.t3216 3.3605
R2970 VSS.t1980 VSS.n13 3.3605
R2971 VSS.n11461 VSS.t1466 3.3605
R2972 VSS.n11465 VSS.t1499 3.3605
R2973 VSS.t1720 VSS.n11093 3.3605
R2974 VSS.t630 VSS.n11087 3.3605
R2975 VSS.t2892 VSS.n11099 3.3605
R2976 VSS.t2920 VSS.n11083 3.3605
R2977 VSS.t1325 VSS.n11105 3.3605
R2978 VSS.t1049 VSS.n11054 3.3605
R2979 VSS.n11111 VSS.t2463 3.3605
R2980 VSS.n11117 VSS.t2488 3.3605
R2981 VSS.n11036 VSS.t2746 3.3605
R2982 VSS.n11122 VSS.t1752 3.3605
R2983 VSS.n11030 VSS.t2674 3.3605
R2984 VSS.n11128 VSS.t1678 3.3605
R2985 VSS.n205 VSS.t2309 3.3605
R2986 VSS.n11137 VSS.t1304 3.3605
R2987 VSS.n11139 VSS.t1189 3.3605
R2988 VSS.n11149 VSS.t1240 3.3605
R2989 VSS.n10882 VSS.t1491 3.3605
R2990 VSS.t1519 VSS.n10877 3.3605
R2991 VSS.n10875 VSS.t537 3.3605
R2992 VSS.n10893 VSS.t3436 3.3605
R2993 VSS.t1404 VSS.n10035 3.3605
R2994 VSS.t3412 VSS.n555 3.3605
R2995 VSS.t2828 VSS.n10042 3.3605
R2996 VSS.t2562 VSS.n552 3.3605
R2997 VSS.n10047 VSS.t2026 3.3605
R2998 VSS.n10053 VSS.t2856 3.3605
R2999 VSS.n542 VSS.t2301 3.3605
R3000 VSS.n10059 VSS.t2063 3.3605
R3001 VSS.n533 VSS.t2760 3.3605
R3002 VSS.t2808 VSS.n531 3.3605
R3003 VSS.t1922 VSS.n516 3.3605
R3004 VSS.t1690 VSS.n503 3.3605
R3005 VSS.n502 VSS.t1085 3.3605
R3006 VSS.n10074 VSS.t1114 3.3605
R3007 VSS.t3308 VSS.n10076 3.3605
R3008 VSS.t3118 VSS.n493 3.3605
R3009 VSS.t3404 VSS.n10084 3.3605
R3010 VSS.t1148 VSS.n484 3.3605
R3011 VSS.t2554 VSS.n10090 3.3605
R3012 VSS.t2678 VSS.n462 3.3605
R3013 VSS.n10096 VSS.t2141 3.3605
R3014 VSS.n10102 VSS.t2956 3.3605
R3015 VSS.n454 VSS.t2053 3.3605
R3016 VSS.n10107 VSS.t1836 3.3605
R3017 VSS.n446 VSS.t2038 3.3605
R3018 VSS.t2870 VSS.n441 3.3605
R3019 VSS.t1978 VSS.n1304 3.3605
R3020 VSS.t1754 VSS.n1298 3.3605
R3021 VSS.t3462 VSS.n1313 3.3605
R3022 VSS.t1191 VSS.n1296 3.3605
R3023 VSS.n12 VSS.t1732 3.3605
R3024 VSS.t1732 VSS.n9 3.3605
R3025 VSS.n11092 VSS.t2750 3.3605
R3026 VSS.n11098 VSS.t2484 3.3605
R3027 VSS.n11085 VSS.t1670 3.3605
R3028 VSS.n11104 VSS.t2451 3.3605
R3029 VSS.n11059 VSS.t1598 3.3605
R3030 VSS.n11110 VSS.t462 3.3605
R3031 VSS.n11112 VSS.t3628 3.3605
R3032 VSS.t3628 VSS.n11053 3.3605
R3033 VSS.t2826 VSS.n11118 3.3605
R3034 VSS.n11119 VSS.t2826 3.3605
R3035 VSS.n11033 VSS.t3580 3.3605
R3036 VSS.n11125 VSS.t3620 3.3605
R3037 VSS.n11026 VSS.t2744 3.3605
R3038 VSS.n11131 VSS.t2868 3.3605
R3039 VSS.n11134 VSS.t2002 3.3605
R3040 VSS.t2816 VSS.n201 3.3605
R3041 VSS.n11146 VSS.t2800 3.3605
R3042 VSS.t2800 VSS.n185 3.3605
R3043 VSS.t1970 VSS.n10883 3.3605
R3044 VSS.n10884 VSS.t1970 3.3605
R3045 VSS.t1167 VSS.n10886 3.3605
R3046 VSS.t904 VSS.n10874 3.3605
R3047 VSS.n10893 VSS.t1906 3.3605
R3048 VSS.t845 VSS.n10870 3.3605
R3049 VSS.t3112 VSS.n10039 3.3605
R3050 VSS.t771 VSS.n550 3.3605
R3051 VSS.t3116 VSS.n10045 3.3605
R3052 VSS.n10046 VSS.t3116 3.3605
R3053 VSS.n10050 VSS.t2279 3.3605
R3054 VSS.t2279 VSS.n543 3.3605
R3055 VSS.t2606 VSS.n10054 3.3605
R3056 VSS.t2367 VSS.n537 3.3605
R3057 VSS.t1539 VSS.n10061 3.3605
R3058 VSS.n530 VSS.t2317 3.3605
R3059 VSS.n526 VSS.t2235 3.3605
R3060 VSS.n517 VSS.t1234 3.3605
R3061 VSS.t1205 VSS.n10070 3.3605
R3062 VSS.n10071 VSS.t1205 3.3605
R3063 VSS.n497 VSS.t3458 3.3605
R3064 VSS.t3458 VSS.n496 3.3605
R3065 VSS.n494 VSS.t3432 3.3605
R3066 VSS.n10083 VSS.t3476 3.3605
R3067 VSS.n490 VSS.t2602 3.3605
R3068 VSS.n10089 VSS.t2357 3.3605
R3069 VSS.n465 VSS.t2550 3.3605
R3070 VSS.n10095 VSS.t2666 3.3605
R3071 VSS.n10097 VSS.t2644 3.3605
R3072 VSS.t2644 VSS.n457 3.3605
R3073 VSS.t1846 VSS.n10103 3.3605
R3074 VSS.n10104 VSS.t1846 3.3605
R3075 VSS.n451 VSS.t1006 3.3605
R3076 VSS.n10110 VSS.t1854 3.3605
R3077 VSS.t1784 VSS.n10112 3.3605
R3078 VSS.n1302 VSS.t712 3.3605
R3079 VSS.n1299 VSS.t2966 3.3605
R3080 VSS.n1311 VSS.t604 3.3605
R3081 VSS.n1273 VSS.t2986 3.3605
R3082 VSS.t2986 VSS.n1272 3.3605
R3083 VSS.n11341 VSS.t2377 3.3605
R3084 VSS.n11345 VSS.t2409 3.3605
R3085 VSS.n11348 VSS.t2656 3.3605
R3086 VSS.n11352 VSS.t1664 3.3605
R3087 VSS.n11354 VSS.t3384 3.3605
R3088 VSS.n11358 VSS.t3426 3.3605
R3089 VSS.t519 VSS.n96 3.3605
R3090 VSS.n10998 VSS.t2684 3.3605
R3091 VSS.n10989 VSS.t2153 3.3605
R3092 VSS.n10985 VSS.t2189 3.3605
R3093 VSS.t2397 VSS.n207 3.3605
R3094 VSS.n10920 VSS.t2429 3.3605
R3095 VSS.n10637 VSS.t1377 3.3605
R3096 VSS.t1377 VSS.n10636 3.3605
R3097 VSS.n10637 VSS.t1110 3.3605
R3098 VSS.n10636 VSS.t1110 3.3605
R3099 VSS.n10637 VSS.t3492 3.3605
R3100 VSS.n10636 VSS.t3492 3.3605
R3101 VSS.t1982 VSS.n10634 3.3605
R3102 VSS.t791 VSS.n10642 3.3605
R3103 VSS.n10648 VSS.t1654 3.3605
R3104 VSS.n10649 VSS.t2399 3.3605
R3105 VSS.t531 VSS.n10347 3.3605
R3106 VSS.n10511 VSS.t531 3.3605
R3107 VSS.n10513 VSS.t661 3.3605
R3108 VSS.t2930 VSS.n10504 3.3605
R3109 VSS.t2289 VSS.n10525 3.3605
R3110 VSS.t3176 VSS.n10489 3.3605
R3111 VSS.n10540 VSS.t3596 3.3605
R3112 VSS.t1694 VSS.n10483 3.3605
R3113 VSS.n10552 VSS.t2842 3.3605
R3114 VSS.t2842 VSS.n10482 3.3605
R3115 VSS.n10512 VSS.t1171 3.3605
R3116 VSS.n10515 VSS.t878 3.3605
R3117 VSS.n10524 VSS.t2756 3.3605
R3118 VSS.n10503 VSS.t1898 3.3605
R3119 VSS.t1898 VSS.n10498 3.3605
R3120 VSS.t705 VSS.n10538 3.3605
R3121 VSS.n10539 VSS.t705 3.3605
R3122 VSS.n10542 VSS.t1894 3.3605
R3123 VSS.n10551 VSS.t3062 3.3605
R3124 VSS.n10589 VSS.t1146 3.3605
R3125 VSS.n10438 VSS.t1475 3.3605
R3126 VSS.t2582 VSS.n10432 3.3605
R3127 VSS.n10431 VSS.t663 3.3605
R3128 VSS.t2932 VSS.n10424 3.3605
R3129 VSS.n10423 VSS.t2291 3.3605
R3130 VSS.t1440 VSS.n10291 3.3605
R3131 VSS.t1144 VSS.n10454 3.3605
R3132 VSS.n10460 VSS.t3316 3.3605
R3133 VSS.t2738 VSS.n10461 3.3605
R3134 VSS.n10468 VSS.t3606 3.3605
R3135 VSS.t926 VSS.n10469 3.3605
R3136 VSS.n10475 VSS.t2119 3.3605
R3137 VSS.t3318 VSS.n10582 3.3605
R3138 VSS.n10581 VSS.t2740 3.3605
R3139 VSS.t1860 VSS.n10575 3.3605
R3140 VSS.n9038 VSS.t2880 3.3605
R3141 VSS.n9016 VSS.t803 3.3605
R3142 VSS.t1087 VSS.n1561 3.3605
R3143 VSS.n1570 VSS.t3470 3.3605
R3144 VSS.n9003 VSS.t2177 3.3605
R3145 VSS.n9007 VSS.t3212 3.3605
R3146 VSS.n8969 VSS.t3478 3.3605
R3147 VSS.n8965 VSS.t2802 3.3605
R3148 VSS.n9099 VSS.t991 3.3605
R3149 VSS.n9095 VSS.t2073 3.3605
R3150 VSS.t1672 VSS.n1554 3.3605
R3151 VSS.n8979 VSS.t498 3.3605
R3152 VSS.n9084 VSS.t1742 3.3605
R3153 VSS.n9088 VSS.t2798 3.3605
R3154 VSS.n9044 VSS.t2343 3.3605
R3155 VSS.n9040 VSS.t1302 3.3605
R3156 VSS.n9063 VSS.t1107 3.3605
R3157 VSS.n9067 VSS.t2201 3.3605
R3158 VSS.n9069 VSS.t2453 3.3605
R3159 VSS.n9073 VSS.t1774 3.3605
R3160 VSS.n974 VSS.t2161 3.3605
R3161 VSS.n970 VSS.t1920 3.3605
R3162 VSS.n968 VSS.t1396 3.3605
R3163 VSS.n964 VSS.t2191 3.3605
R3164 VSS.n10262 VSS.t1199 3.3605
R3165 VSS.n10271 VSS.t922 3.3605
R3166 VSS.n10273 VSS.t3498 3.3605
R3167 VSS.n10277 VSS.t1245 3.3605
R3168 VSS.n312 VSS.t3272 3.3605
R3169 VSS.n308 VSS.t3074 3.3605
R3170 VSS.n306 VSS.t2465 3.3605
R3171 VSS.t2494 VSS.n272 3.3605
R3172 VSS.n990 VSS.t1121 3.3605
R3173 VSS.n986 VSS.t876 3.3605
R3174 VSS.n984 VSS.t3386 3.3605
R3175 VSS.n976 VSS.t3428 3.3605
R3176 VSS.n1011 VSS.t2379 3.3605
R3177 VSS.n1007 VSS.t2169 3.3605
R3178 VSS.n1005 VSS.t1638 3.3605
R3179 VSS.n1001 VSS.t2411 3.3605
R3180 VSS.n10223 VSS.t1479 3.3605
R3181 VSS.n10219 VSS.t1209 3.3605
R3182 VSS.n318 VSS.t599 3.3605
R3183 VSS.n314 VSS.t1501 3.3605
R3184 VSS.n10202 VSS.t3174 3.3605
R3185 VSS.n10211 VSS.t3200 3.3605
R3186 VSS.n10213 VSS.t3406 3.3605
R3187 VSS.n10217 VSS.t3450 3.3605
R3188 VSS.n1023 VSS.t1004 3.3605
R3189 VSS.n1019 VSS.t1043 3.3605
R3190 VSS.n1017 VSS.t1309 3.3605
R3191 VSS.n1013 VSS.t1350 3.3605
R3192 VSS.n1048 VSS.t2311 3.3605
R3193 VSS.n1044 VSS.t2339 3.3605
R3194 VSS.n1042 VSS.t2952 3.3605
R3195 VSS.n1034 VSS.t1932 3.3605
R3196 VSS.n375 VSS.t1394 3.3605
R3197 VSS.n371 VSS.t1428 3.3605
R3198 VSS.n369 VSS.t1990 3.3605
R3199 VSS.t938 VSS.n344 3.3605
R3200 VSS.n10163 VSS.t3380 3.3605
R3201 VSS.n10159 VSS.t3420 3.3605
R3202 VSS.n390 VSS.t509 3.3605
R3203 VSS.n386 VSS.t2676 3.3605
R3204 VSS.n1060 VSS.t1284 3.3605
R3205 VSS.n1056 VSS.t1329 3.3605
R3206 VSS.n1054 VSS.t1570 3.3605
R3207 VSS.n1050 VSS.t3612 3.3605
R3208 VSS.n1081 VSS.t2680 3.3605
R3209 VSS.n1077 VSS.t3466 3.3605
R3210 VSS.n1075 VSS.t2149 3.3605
R3211 VSS.n1071 VSS.t1910 3.3605
R3212 VSS.n10142 VSS.t1748 3.3605
R3213 VSS.n10151 VSS.t2528 3.3605
R3214 VSS.n10153 VSS.t1187 3.3605
R3215 VSS.n10157 VSS.t918 3.3605
R3216 VSS.n1294 VSS.t3322 3.3605
R3217 VSS.n1290 VSS.t3130 3.3605
R3218 VSS.n1288 VSS.t3618 3.3605
R3219 VSS.t3354 VSS.n416 3.3605
R3220 VSS.n1097 VSS.t1223 3.3605
R3221 VSS.n1093 VSS.t955 3.3605
R3222 VSS.n1091 VSS.t1513 3.3605
R3223 VSS.n1083 VSS.t1254 3.3605
R3224 VSS.n1118 VSS.t2938 3.3605
R3225 VSS.n1114 VSS.t2692 3.3605
R3226 VSS.n1112 VSS.t1364 3.3605
R3227 VSS.n1108 VSS.t2157 3.3605
R3228 VSS.n1130 VSS.t3510 3.3605
R3229 VSS.n1126 VSS.t3616 3.3605
R3230 VSS.n1124 VSS.t3110 3.3605
R3231 VSS.n1120 VSS.t760 3.3605
R3232 VSS.n862 VSS.t2874 3.3605
R3233 VSS.n866 VSS.t2612 3.3605
R3234 VSS.n869 VSS.t2051 3.3605
R3235 VSS.n877 VSS.t2079 3.3605
R3236 VSS.n10922 VSS.t612 3.3605
R3237 VSS.n10926 VSS.t3518 3.3605
R3238 VSS.t2996 VSS.n221 3.3605
R3239 VSS.n842 VSS.t636 3.3605
R3240 VSS.n10364 VSS.t3452 3.3605
R3241 VSS.t1181 VSS.n10358 3.3605
R3242 VSS.n10357 VSS.t1974 3.3605
R3243 VSS.n10669 VSS.t684 3.3605
R3244 VSS.t3542 VSS.n10670 3.3605
R3245 VSS.n10676 VSS.t2307 3.3605
R3246 VSS.n9473 VSS.t1408 3.3605
R3247 VSS.n9469 VSS.t3014 3.3605
R3248 VSS.t3520 VSS.n1380 3.3605
R3249 VSS.n9433 VSS.t2043 3.3605
R3250 VSS.n9461 VSS.t306 3.3605
R3251 VSS.n9461 VSS.t309 3.3605
R3252 VSS.n9460 VSS.t310 3.3605
R3253 VSS.n9460 VSS.t441 3.3605
R3254 VSS.n9459 VSS.t307 3.3605
R3255 VSS.n9459 VSS.t304 3.3605
R3256 VSS.n1379 VSS.t311 3.3605
R3257 VSS.n1379 VSS.t308 3.3605
R3258 VSS.n9454 VSS.t1243 3.3605
R3259 VSS.n9458 VSS.t2482 3.3605
R3260 VSS.n9452 VSS.t1801 3.3605
R3261 VSS.n9448 VSS.t3092 3.3605
R3262 VSS.n9974 VSS.t1035 3.3605
R3263 VSS.n9978 VSS.t3178 3.3605
R3264 VSS.n9980 VSS.t2363 3.3605
R3265 VSS.n9984 VSS.t1028 3.3605
R3266 VSS.n9986 VSS.t3098 3.3605
R3267 VSS.n9990 VSS.t3152 3.3605
R3268 VSS.t3578 VSS.n9991 3.3605
R3269 VSS.n9992 VSS.t3578 3.3605
R3270 VSS.t2431 VSS.n9994 3.3605
R3271 VSS.n9995 VSS.t2431 3.3605
R3272 VSS.n9996 VSS.t2127 3.3605
R3273 VSS.n10000 VSS.t1858 3.3605
R3274 VSS.n10002 VSS.t741 3.3605
R3275 VSS.n10006 VSS.t1590 3.3605
R3276 VSS.n10008 VSS.t733 3.3605
R3277 VSS.n10012 VSS.t2524 3.3605
R3278 VSS.t2998 VSS.n10013 3.3605
R3279 VSS.n10014 VSS.t2998 3.3605
R3280 VSS.t1848 VSS.n10016 3.3605
R3281 VSS.n10017 VSS.t1848 3.3605
R3282 VSS.n10019 VSS.t3304 3.3605
R3283 VSS.n10024 VSS.t2351 3.3605
R3284 VSS.t3236 VSS.n10027 3.3605
R3285 VSS.n9721 VSS.t3302 3.3605
R3286 VSS.n9723 VSS.t2249 3.3605
R3287 VSS.n9727 VSS.t906 3.3605
R3288 VSS.t2421 VSS.n9728 3.3605
R3289 VSS.n9729 VSS.t2421 3.3605
R3290 VSS.t1280 VSS.n9731 3.3605
R3291 VSS.n9732 VSS.t1280 3.3605
R3292 VSS.n9733 VSS.t3484 3.3605
R3293 VSS.n9737 VSS.t2522 3.3605
R3294 VSS.n9739 VSS.t1740 3.3605
R3295 VSS.n9743 VSS.t3480 3.3605
R3296 VSS.n9745 VSS.t1662 3.3605
R3297 VSS.n9749 VSS.t1730 3.3605
R3298 VSS.t2183 VSS.n9750 3.3605
R3299 VSS.n9751 VSS.t2183 3.3605
R3300 VSS.t987 VSS.n9753 3.3605
R3301 VSS.n9754 VSS.t987 3.3605
R3302 VSS.n9755 VSS.t1497 3.3605
R3303 VSS.n9759 VSS.t1201 3.3605
R3304 VSS.t3202 VSS.n9761 3.3605
R3305 VSS.t2237 VSS.n9635 3.3605
R3306 VSS.n9633 VSS.t1065 3.3605
R3307 VSS.n9629 VSS.t1892 3.3605
R3308 VSS.n9628 VSS.t2327 3.3605
R3309 VSS.t2327 VSS.n9627 3.3605
R3310 VSS.t1175 VSS.n805 3.3605
R3311 VSS.n1355 VSS.t1175 3.3605
R3312 VSS.n1357 VSS.t2704 3.3605
R3313 VSS.n1362 VSS.t1389 3.3605
R3314 VSS.n1364 VSS.t2592 3.3605
R3315 VSS.n1368 VSS.t2690 3.3605
R3316 VSS.n1370 VSS.t1630 3.3605
R3317 VSS.n1374 VSS.t3334 3.3605
R3318 VSS.n9974 VSS.t811 3.3605
R3319 VSS.n9978 VSS.t1912 3.3605
R3320 VSS.n9980 VSS.t3036 3.3605
R3321 VSS.n9984 VSS.t2303 3.3605
R3322 VSS.n9986 VSS.t2730 3.3605
R3323 VSS.n9990 VSS.t3396 3.3605
R3324 VSS.n9991 VSS.t1452 3.3605
R3325 VSS.n9992 VSS.t1452 3.3605
R3326 VSS.n9994 VSS.t3358 3.3605
R3327 VSS.n9995 VSS.t3358 3.3605
R3328 VSS.n9996 VSS.t2417 3.3605
R3329 VSS.n10000 VSS.t1398 3.3605
R3330 VSS.n10002 VSS.t1805 3.3605
R3331 VSS.n10006 VSS.t977 3.3605
R3332 VSS.n10008 VSS.t2125 3.3605
R3333 VSS.n10012 VSS.t1442 3.3605
R3334 VSS.n10013 VSS.t2469 3.3605
R3335 VSS.n10014 VSS.t2469 3.3605
R3336 VSS.n10016 VSS.t1385 3.3605
R3337 VSS.n10017 VSS.t1385 3.3605
R3338 VSS.n10019 VSS.t2099 3.3605
R3339 VSS.n10024 VSS.t3160 3.3605
R3340 VSS.n10027 VSS.t2864 3.3605
R3341 VSS.n9721 VSS.t3554 3.3605
R3342 VSS.n9723 VSS.t854 3.3605
R3343 VSS.n9727 VSS.t3254 3.3605
R3344 VSS.n9728 VSS.t880 3.3605
R3345 VSS.n9729 VSS.t880 3.3605
R3346 VSS.n9731 VSS.t2894 3.3605
R3347 VSS.n9732 VSS.t2894 3.3605
R3348 VSS.n9733 VSS.t2121 3.3605
R3349 VSS.n9737 VSS.t3172 3.3605
R3350 VSS.n9739 VSS.t1193 3.3605
R3351 VSS.n9743 VSS.t3570 3.3605
R3352 VSS.n9745 VSS.t1958 3.3605
R3353 VSS.n9749 VSS.t2662 3.3605
R3354 VSS.n9750 VSS.t591 3.3605
R3355 VSS.n9751 VSS.t591 3.3605
R3356 VSS.n9753 VSS.t2620 3.3605
R3357 VSS.n9754 VSS.t2620 3.3605
R3358 VSS.n9755 VSS.t523 3.3605
R3359 VSS.n9759 VSS.t2636 3.3605
R3360 VSS.n9761 VSS.t3086 3.3605
R3361 VSS.n9635 VSS.t997 3.3605
R3362 VSS.n9633 VSS.t3434 3.3605
R3363 VSS.t2694 VSS.n9629 3.3605
R3364 VSS.n9628 VSS.t607 3.3605
R3365 VSS.n9627 VSS.t607 3.3605
R3366 VSS.t2630 VSS.n805 3.3605
R3367 VSS.n1355 VSS.t2630 3.3605
R3368 VSS.n1357 VSS.t3332 3.3605
R3369 VSS.n1362 VSS.t2660 3.3605
R3370 VSS.n1364 VSS.t1001 3.3605
R3371 VSS.n1368 VSS.t1768 3.3605
R3372 VSS.n1370 VSS.t2173 3.3605
R3373 VSS.n1374 VSS.t1485 3.3605
R3374 VSS.n10822 VSS.t1435 3.3605
R3375 VSS.n9197 VSS.n9196 3.27473
R3376 VSS.n9333 VSS.n9332 3.27473
R3377 VSS.n171 VSS.n170 3.27473
R3378 VSS.n9579 VSS.n9578 3.27473
R3379 VSS.n199 VSS.n198 3.27473
R3380 VSS.n477 VSS.n476 3.27473
R3381 VSS.n9030 VSS.n9029 3.27473
R3382 VSS.n270 VSS.n269 3.27473
R3383 VSS.n342 VSS.n341 3.27473
R3384 VSS.n414 VSS.n413 3.27473
R3385 VSS.t638 VSS.t303 3.2333
R3386 VSS.n1391 VSS.t593 3.19467
R3387 VSS.n10325 VSS.n10323 3.15563
R3388 VSS.n10329 VSS.n10327 3.15563
R3389 VSS.n10318 VSS.n10316 3.15563
R3390 VSS.n10314 VSS.n10312 3.15563
R3391 VSS.n10757 VSS.n10756 3.1505
R3392 VSS.n10767 VSS.n10766 3.1505
R3393 VSS.n11289 VSS.t325 3.02895
R3394 VSS.n10309 VSS.n10308 3.02463
R3395 VSS.n10408 VSS.n10406 2.96616
R3396 VSS.n10401 VSS.n10399 2.96616
R3397 VSS.n10378 VSS.n10377 2.885
R3398 VSS.n10623 VSS.n10622 2.885
R3399 VSS.n10614 VSS.n10613 2.795
R3400 VSS.n10408 VSS.n10407 2.76247
R3401 VSS.n10401 VSS.n10400 2.76247
R3402 VSS.n10297 VSS.n10296 2.74471
R3403 VSS.n10403 VSS.n10401 2.71914
R3404 VSS.n10326 VSS.n10322 2.71872
R3405 VSS.n9526 VSS.t257 2.71016
R3406 VSS.n10818 VSS.t3210 2.6955
R3407 VSS.n10814 VSS.t1914 2.6955
R3408 VSS.n10748 VSS.t894 2.6955
R3409 VSS.n10752 VSS.t586 2.6955
R3410 VSS.n10787 VSS.t3550 2.6955
R3411 VSS.n10783 VSS.t2239 2.6955
R3412 VSS.n10781 VSS.t1268 2.6955
R3413 VSS.n10777 VSS.t967 2.6955
R3414 VSS.n9193 VSS.n9192 2.68042
R3415 VSS.n9188 VSS.n9187 2.68042
R3416 VSS.n9329 VSS.n9328 2.68042
R3417 VSS.n9324 VSS.n9323 2.68042
R3418 VSS.n167 VSS.n166 2.68042
R3419 VSS.n162 VSS.n161 2.68042
R3420 VSS.n9575 VSS.n9574 2.68042
R3421 VSS.n9570 VSS.n9569 2.68042
R3422 VSS.n9026 VSS.n9025 2.68042
R3423 VSS.n9021 VSS.n9020 2.68042
R3424 VSS.n190 VSS.n189 2.68012
R3425 VSS.n195 VSS.n194 2.68012
R3426 VSS.n468 VSS.n467 2.68012
R3427 VSS.n473 VSS.n472 2.68012
R3428 VSS.n261 VSS.n260 2.68012
R3429 VSS.n266 VSS.n265 2.68012
R3430 VSS.n333 VSS.n332 2.68012
R3431 VSS.n338 VSS.n337 2.68012
R3432 VSS.n405 VSS.n404 2.68012
R3433 VSS.n410 VSS.n409 2.68012
R3434 VSS.n4804 VSS.n4803 2.66637
R3435 VSS.n10866 VSS.n10864 2.65976
R3436 VSS.n9560 VSS.t259 2.63047
R3437 VSS.n10769 VSS.t3154 2.6255
R3438 VSS.n10772 VSS.t1828 2.6255
R3439 VSS.n10770 VSS.t3604 2.6255
R3440 VSS.n10741 VSS.t2233 2.6255
R3441 VSS.n10745 VSS.t3244 2.6255
R3442 VSS.n10663 VSS.n10662 2.60959
R3443 VSS.n9612 VSS.n813 2.58721
R3444 VSS.n9877 VSS.n669 2.58721
R3445 VSS.n656 VSS.n655 2.58721
R3446 VSS.n821 VSS.n820 2.58721
R3447 VSS.n677 VSS.n676 2.58721
R3448 VSS.n11416 VSS.n45 2.58721
R3449 VSS.n11449 VSS.n20 2.58721
R3450 VSS.n9920 VSS.n585 2.58721
R3451 VSS.n9913 VSS.n9908 2.58721
R3452 VSS.n9513 VSS.n1329 2.58721
R3453 VSS.n1253 VSS.n1252 2.58721
R3454 VSS.n9901 VSS.n9900 2.58721
R3455 VSS.n652 VSS.n651 2.58366
R3456 VSS.n817 VSS.n816 2.58366
R3457 VSS.n9858 VSS.n9857 2.58366
R3458 VSS.n9874 VSS.n670 2.58366
R3459 VSS.n11413 VSS.n46 2.58366
R3460 VSS.n11446 VSS.n21 2.58366
R3461 VSS.n9897 VSS.n629 2.58366
R3462 VSS.n1249 VSS.n1248 2.58366
R3463 VSS.n9516 VSS.n1328 2.58366
R3464 VSS.n9910 VSS.n9909 2.58366
R3465 VSS.n9924 VSS.n9923 2.58366
R3466 VSS.n9615 VSS.n812 2.58366
R3467 VSS.n10325 VSS.n10324 2.573
R3468 VSS.n10329 VSS.n10328 2.573
R3469 VSS.n10318 VSS.n10317 2.573
R3470 VSS.n10314 VSS.n10313 2.573
R3471 VSS.n10625 VSS.n10624 2.55405
R3472 VSS.n10616 VSS.n10615 2.55405
R3473 VSS.n10380 VSS.n10379 2.55405
R3474 VSS.t413 VSS.t750 2.55077
R3475 VSS.n10733 VSS.t1761 2.5394
R3476 VSS.t1248 VSS.n9434 2.53859
R3477 VSS.n9447 VSS.t2100 2.53837
R3478 VSS.n11304 VSS.t3423 2.53699
R3479 VSS.t3571 VSS.n10838 2.52844
R3480 VSS.n10839 VSS.t3571 2.52844
R3481 VSS.t821 VSS.n10835 2.52844
R3482 VSS.n10836 VSS.t821 2.52844
R3483 VSS.t2470 VSS.n10832 2.52844
R3484 VSS.n10833 VSS.t2470 2.52844
R3485 VSS.t1196 VSS.n10829 2.52844
R3486 VSS.n10830 VSS.t1196 2.52844
R3487 VSS.t3017 VSS.n10826 2.52844
R3488 VSS.n10827 VSS.t3017 2.52844
R3489 VSS.n10727 VSS.t1761 2.52844
R3490 VSS.t3529 VSS.n10725 2.52844
R3491 VSS.n10726 VSS.t3529 2.52844
R3492 VSS.t767 VSS.n10723 2.52844
R3493 VSS.n10724 VSS.t767 2.52844
R3494 VSS.t2438 VSS.n10721 2.52844
R3495 VSS.n10722 VSS.t2438 2.52844
R3496 VSS.t1135 VSS.n10718 2.52844
R3497 VSS.n10719 VSS.t1135 2.52844
R3498 VSS.n10717 VSS.t2963 2.52844
R3499 VSS.t2963 VSS.n10716 2.52844
R3500 VSS.t1679 VSS.n10714 2.52844
R3501 VSS.n10715 VSS.t1679 2.52844
R3502 VSS.t3423 VSS.n125 2.52844
R3503 VSS.n1338 VSS.t1699 2.52844
R3504 VSS.t1699 VSS.n1337 2.52844
R3505 VSS.n1341 VSS.t2557 2.52844
R3506 VSS.t2557 VSS.n1340 2.52844
R3507 VSS.n9499 VSS.t1745 2.52844
R3508 VSS.t1745 VSS.n1343 2.52844
R3509 VSS.n9496 VSS.t488 2.52844
R3510 VSS.t488 VSS.n9495 2.52844
R3511 VSS.t3005 VSS.n9491 2.52844
R3512 VSS.n9492 VSS.t3005 2.52844
R3513 VSS.t1555 VSS.n9488 2.52844
R3514 VSS.n9489 VSS.t1555 2.52844
R3515 VSS.n9445 VSS.t2100 2.52844
R3516 VSS.t3003 VSS.n9443 2.52844
R3517 VSS.n9444 VSS.t3003 2.52844
R3518 VSS.t2158 VSS.n9441 2.52844
R3519 VSS.n9442 VSS.t2158 2.52844
R3520 VSS.t3345 VSS.n9438 2.52844
R3521 VSS.n9439 VSS.t3345 2.52844
R3522 VSS.t2711 VSS.n9436 2.52844
R3523 VSS.n9437 VSS.t2711 2.52844
R3524 VSS.n9435 VSS.t1248 2.52844
R3525 VSS.n10410 VSS.n10403 2.46014
R3526 VSS.n10796 VSS.n247 2.45973
R3527 VSS.n10808 VSS.n10807 2.45073
R3528 VSS.n10333 VSS.n10321 2.38034
R3529 VSS.n10392 VSS.n10365 2.37491
R3530 VSS.n10398 VSS.n10397 2.32143
R3531 VSS.n11152 VSS.n181 2.31168
R3532 VSS.n10611 VSS.n10610 2.30076
R3533 VSS.n10018 VSS.n576 2.28095
R3534 VSS.n573 VSS.n572 2.28095
R3535 VSS.n1356 VSS.n1353 2.28095
R3536 VSS.n10020 VSS.n576 2.27641
R3537 VSS.n10025 VSS.n572 2.27641
R3538 VSS.n1358 VSS.n1353 2.27641
R3539 VSS.n228 VSS.n227 2.26832
R3540 VSS.n10679 VSS.n10303 2.26738
R3541 VSS.n5468 VSS.n2743 2.2505
R3542 VSS.n5467 VSS.n5466 2.2505
R3543 VSS.n5465 VSS.n2744 2.2505
R3544 VSS.n5464 VSS.n5463 2.2505
R3545 VSS.n5462 VSS.n2745 2.2505
R3546 VSS.n5461 VSS.n5460 2.2505
R3547 VSS.n5459 VSS.n2746 2.2505
R3548 VSS.n5458 VSS.n5457 2.2505
R3549 VSS.n5456 VSS.n2747 2.2505
R3550 VSS.n5455 VSS.n5454 2.2505
R3551 VSS.n5453 VSS.n2748 2.2505
R3552 VSS.n5452 VSS.n5451 2.2505
R3553 VSS.n5450 VSS.n2749 2.2505
R3554 VSS.n5449 VSS.n5448 2.2505
R3555 VSS.n5447 VSS.n2750 2.2505
R3556 VSS.n5446 VSS.n5445 2.2505
R3557 VSS.n5444 VSS.n2751 2.2505
R3558 VSS.n5443 VSS.n5442 2.2505
R3559 VSS.n5441 VSS.n2752 2.2505
R3560 VSS.n5440 VSS.n5439 2.2505
R3561 VSS.n5438 VSS.n2753 2.2505
R3562 VSS.n5437 VSS.n5436 2.2505
R3563 VSS.n5435 VSS.n2754 2.2505
R3564 VSS.n5434 VSS.n5433 2.2505
R3565 VSS.n5432 VSS.n2755 2.2505
R3566 VSS.n5431 VSS.n5430 2.2505
R3567 VSS.n5429 VSS.n2756 2.2505
R3568 VSS.n5428 VSS.n5427 2.2505
R3569 VSS.n5426 VSS.n2757 2.2505
R3570 VSS.n5425 VSS.n5424 2.2505
R3571 VSS.n5423 VSS.n2758 2.2505
R3572 VSS.n5422 VSS.n5421 2.2505
R3573 VSS.n5420 VSS.n2759 2.2505
R3574 VSS.n5419 VSS.n5418 2.2505
R3575 VSS.n5417 VSS.n2760 2.2505
R3576 VSS.n5416 VSS.n5415 2.2505
R3577 VSS.n5414 VSS.n2761 2.2505
R3578 VSS.n5413 VSS.n5412 2.2505
R3579 VSS.n5411 VSS.n2762 2.2505
R3580 VSS.n5410 VSS.n5409 2.2505
R3581 VSS.n5408 VSS.n2763 2.2505
R3582 VSS.n5407 VSS.n5406 2.2505
R3583 VSS.n5405 VSS.n2764 2.2505
R3584 VSS.n5404 VSS.n5403 2.2505
R3585 VSS.n5402 VSS.n2765 2.2505
R3586 VSS.n5401 VSS.n5400 2.2505
R3587 VSS.n5399 VSS.n2766 2.2505
R3588 VSS.n5398 VSS.n5397 2.2505
R3589 VSS.n5396 VSS.n2767 2.2505
R3590 VSS.n5395 VSS.n5394 2.2505
R3591 VSS.n5393 VSS.n2768 2.2505
R3592 VSS.n5392 VSS.n5391 2.2505
R3593 VSS.n5390 VSS.n2769 2.2505
R3594 VSS.n5389 VSS.n5388 2.2505
R3595 VSS.n5387 VSS.n2770 2.2505
R3596 VSS.n5386 VSS.n5385 2.2505
R3597 VSS.n5384 VSS.n2771 2.2505
R3598 VSS.n5383 VSS.n5382 2.2505
R3599 VSS.n5381 VSS.n2772 2.2505
R3600 VSS.n5380 VSS.n5379 2.2505
R3601 VSS.n5378 VSS.n2773 2.2505
R3602 VSS.n5377 VSS.n5376 2.2505
R3603 VSS.n5375 VSS.n2774 2.2505
R3604 VSS.n5374 VSS.n5373 2.2505
R3605 VSS.n5372 VSS.n2775 2.2505
R3606 VSS.n5371 VSS.n5370 2.2505
R3607 VSS.n5369 VSS.n2776 2.2505
R3608 VSS.n5368 VSS.n5367 2.2505
R3609 VSS.n5366 VSS.n2777 2.2505
R3610 VSS.n5365 VSS.n5364 2.2505
R3611 VSS.n5363 VSS.n2778 2.2505
R3612 VSS.n5362 VSS.n5361 2.2505
R3613 VSS.n5360 VSS.n2779 2.2505
R3614 VSS.n5359 VSS.n5358 2.2505
R3615 VSS.n5357 VSS.n2780 2.2505
R3616 VSS.n5356 VSS.n5355 2.2505
R3617 VSS.n5354 VSS.n2781 2.2505
R3618 VSS.n5353 VSS.n5352 2.2505
R3619 VSS.n5351 VSS.n2782 2.2505
R3620 VSS.n5350 VSS.n5349 2.2505
R3621 VSS.n5348 VSS.n2783 2.2505
R3622 VSS.n5347 VSS.n5346 2.2505
R3623 VSS.n5345 VSS.n2784 2.2505
R3624 VSS.n5344 VSS.n5343 2.2505
R3625 VSS.n5342 VSS.n2785 2.2505
R3626 VSS.n5341 VSS.n5340 2.2505
R3627 VSS.n5339 VSS.n2786 2.2505
R3628 VSS.n5338 VSS.n5337 2.2505
R3629 VSS.n5336 VSS.n2787 2.2505
R3630 VSS.n5335 VSS.n5334 2.2505
R3631 VSS.n5333 VSS.n2788 2.2505
R3632 VSS.n5332 VSS.n5331 2.2505
R3633 VSS.n5330 VSS.n2789 2.2505
R3634 VSS.n5329 VSS.n5328 2.2505
R3635 VSS.n5327 VSS.n2790 2.2505
R3636 VSS.n5326 VSS.n5325 2.2505
R3637 VSS.n5324 VSS.n2791 2.2505
R3638 VSS.n5323 VSS.n5322 2.2505
R3639 VSS.n5321 VSS.n2792 2.2505
R3640 VSS.n5320 VSS.n5319 2.2505
R3641 VSS.n5318 VSS.n2793 2.2505
R3642 VSS.n5317 VSS.n5316 2.2505
R3643 VSS.n5315 VSS.n2794 2.2505
R3644 VSS.n5314 VSS.n5313 2.2505
R3645 VSS.n5312 VSS.n2795 2.2505
R3646 VSS.n5311 VSS.n5310 2.2505
R3647 VSS.n5309 VSS.n2796 2.2505
R3648 VSS.n5308 VSS.n5307 2.2505
R3649 VSS.n5306 VSS.n2797 2.2505
R3650 VSS.n5305 VSS.n5304 2.2505
R3651 VSS.n5303 VSS.n2798 2.2505
R3652 VSS.n5302 VSS.n5301 2.2505
R3653 VSS.n5300 VSS.n2799 2.2505
R3654 VSS.n5299 VSS.n5298 2.2505
R3655 VSS.n5297 VSS.n2800 2.2505
R3656 VSS.n5296 VSS.n5295 2.2505
R3657 VSS.n5294 VSS.n2801 2.2505
R3658 VSS.n5293 VSS.n5292 2.2505
R3659 VSS.n5291 VSS.n2802 2.2505
R3660 VSS.n5290 VSS.n5289 2.2505
R3661 VSS.n5288 VSS.n2803 2.2505
R3662 VSS.n5287 VSS.n5286 2.2505
R3663 VSS.n5285 VSS.n2804 2.2505
R3664 VSS.n5284 VSS.n5283 2.2505
R3665 VSS.n5282 VSS.n2805 2.2505
R3666 VSS.n5281 VSS.n5280 2.2505
R3667 VSS.n5279 VSS.n2806 2.2505
R3668 VSS.n5278 VSS.n5277 2.2505
R3669 VSS.n5276 VSS.n2807 2.2505
R3670 VSS.n5275 VSS.n5274 2.2505
R3671 VSS.n5273 VSS.n2808 2.2505
R3672 VSS.n5272 VSS.n5271 2.2505
R3673 VSS.n5270 VSS.n2809 2.2505
R3674 VSS.n5269 VSS.n5268 2.2505
R3675 VSS.n5267 VSS.n2810 2.2505
R3676 VSS.n5266 VSS.n5265 2.2505
R3677 VSS.n5264 VSS.n2811 2.2505
R3678 VSS.n5263 VSS.n5262 2.2505
R3679 VSS.n5261 VSS.n2812 2.2505
R3680 VSS.n5260 VSS.n5259 2.2505
R3681 VSS.n5258 VSS.n2813 2.2505
R3682 VSS.n5257 VSS.n5256 2.2505
R3683 VSS.n5255 VSS.n2814 2.2505
R3684 VSS.n5254 VSS.n5253 2.2505
R3685 VSS.n5252 VSS.n2815 2.2505
R3686 VSS.n5251 VSS.n5250 2.2505
R3687 VSS.n5249 VSS.n2816 2.2505
R3688 VSS.n5248 VSS.n5247 2.2505
R3689 VSS.n5246 VSS.n2817 2.2505
R3690 VSS.n5245 VSS.n5244 2.2505
R3691 VSS.n5243 VSS.n2818 2.2505
R3692 VSS.n5242 VSS.n5241 2.2505
R3693 VSS.n5240 VSS.n2819 2.2505
R3694 VSS.n5239 VSS.n5238 2.2505
R3695 VSS.n5237 VSS.n2820 2.2505
R3696 VSS.n5236 VSS.n5235 2.2505
R3697 VSS.n5234 VSS.n2821 2.2505
R3698 VSS.n5233 VSS.n5232 2.2505
R3699 VSS.n5231 VSS.n2822 2.2505
R3700 VSS.n5230 VSS.n5229 2.2505
R3701 VSS.n5228 VSS.n2823 2.2505
R3702 VSS.n5227 VSS.n5226 2.2505
R3703 VSS.n5225 VSS.n2824 2.2505
R3704 VSS.n5224 VSS.n5223 2.2505
R3705 VSS.n5222 VSS.n2825 2.2505
R3706 VSS.n5221 VSS.n5220 2.2505
R3707 VSS.n5219 VSS.n2826 2.2505
R3708 VSS.n5218 VSS.n5217 2.2505
R3709 VSS.n5216 VSS.n2827 2.2505
R3710 VSS.n5215 VSS.n5214 2.2505
R3711 VSS.n5213 VSS.n2828 2.2505
R3712 VSS.n5212 VSS.n5211 2.2505
R3713 VSS.n5210 VSS.n2829 2.2505
R3714 VSS.n5209 VSS.n5208 2.2505
R3715 VSS.n5207 VSS.n2830 2.2505
R3716 VSS.n5206 VSS.n5205 2.2505
R3717 VSS.n5204 VSS.n2831 2.2505
R3718 VSS.n5203 VSS.n5202 2.2505
R3719 VSS.n5201 VSS.n2832 2.2505
R3720 VSS.n5200 VSS.n5199 2.2505
R3721 VSS.n5198 VSS.n2833 2.2505
R3722 VSS.n5197 VSS.n5196 2.2505
R3723 VSS.n5195 VSS.n2834 2.2505
R3724 VSS.n5194 VSS.n5193 2.2505
R3725 VSS.n5192 VSS.n2835 2.2505
R3726 VSS.n5191 VSS.n5190 2.2505
R3727 VSS.n5189 VSS.n2836 2.2505
R3728 VSS.n5188 VSS.n5187 2.2505
R3729 VSS.n5186 VSS.n2837 2.2505
R3730 VSS.n5185 VSS.n5184 2.2505
R3731 VSS.n5183 VSS.n2838 2.2505
R3732 VSS.n5182 VSS.n5181 2.2505
R3733 VSS.n5180 VSS.n2839 2.2505
R3734 VSS.n5179 VSS.n5178 2.2505
R3735 VSS.n5177 VSS.n2840 2.2505
R3736 VSS.n5176 VSS.n5175 2.2505
R3737 VSS.n5174 VSS.n2841 2.2505
R3738 VSS.n5173 VSS.n5172 2.2505
R3739 VSS.n5171 VSS.n2842 2.2505
R3740 VSS.n5170 VSS.n5169 2.2505
R3741 VSS.n5168 VSS.n2843 2.2505
R3742 VSS.n5167 VSS.n5166 2.2505
R3743 VSS.n5165 VSS.n2844 2.2505
R3744 VSS.n5164 VSS.n5163 2.2505
R3745 VSS.n5162 VSS.n2845 2.2505
R3746 VSS.n5161 VSS.n5160 2.2505
R3747 VSS.n5159 VSS.n2846 2.2505
R3748 VSS.n5158 VSS.n5157 2.2505
R3749 VSS.n5156 VSS.n2847 2.2505
R3750 VSS.n5155 VSS.n5154 2.2505
R3751 VSS.n5153 VSS.n2848 2.2505
R3752 VSS.n5152 VSS.n5151 2.2505
R3753 VSS.n5150 VSS.n2849 2.2505
R3754 VSS.n5149 VSS.n5148 2.2505
R3755 VSS.n5147 VSS.n2850 2.2505
R3756 VSS.n5146 VSS.n5145 2.2505
R3757 VSS.n5144 VSS.n2851 2.2505
R3758 VSS.n5143 VSS.n5142 2.2505
R3759 VSS.n5141 VSS.n2852 2.2505
R3760 VSS.n5140 VSS.n5139 2.2505
R3761 VSS.n5138 VSS.n2853 2.2505
R3762 VSS.n5137 VSS.n5136 2.2505
R3763 VSS.n5135 VSS.n2854 2.2505
R3764 VSS.n5134 VSS.n5133 2.2505
R3765 VSS.n5132 VSS.n2855 2.2505
R3766 VSS.n5131 VSS.n5130 2.2505
R3767 VSS.n5129 VSS.n2856 2.2505
R3768 VSS.n5128 VSS.n5127 2.2505
R3769 VSS.n5126 VSS.n2857 2.2505
R3770 VSS.n5125 VSS.n5124 2.2505
R3771 VSS.n5123 VSS.n2858 2.2505
R3772 VSS.n5122 VSS.n5121 2.2505
R3773 VSS.n5120 VSS.n2859 2.2505
R3774 VSS.n5119 VSS.n5118 2.2505
R3775 VSS.n5117 VSS.n2860 2.2505
R3776 VSS.n5116 VSS.n5115 2.2505
R3777 VSS.n5114 VSS.n2861 2.2505
R3778 VSS.n5113 VSS.n5112 2.2505
R3779 VSS.n5111 VSS.n2862 2.2505
R3780 VSS.n5110 VSS.n5109 2.2505
R3781 VSS.n5108 VSS.n2863 2.2505
R3782 VSS.n5107 VSS.n5106 2.2505
R3783 VSS.n5105 VSS.n2864 2.2505
R3784 VSS.n5104 VSS.n5103 2.2505
R3785 VSS.n5102 VSS.n2865 2.2505
R3786 VSS.n5101 VSS.n5100 2.2505
R3787 VSS.n5099 VSS.n2866 2.2505
R3788 VSS.n5098 VSS.n5097 2.2505
R3789 VSS.n5096 VSS.n2867 2.2505
R3790 VSS.n5095 VSS.n5094 2.2505
R3791 VSS.n5093 VSS.n2868 2.2505
R3792 VSS.n5092 VSS.n5091 2.2505
R3793 VSS.n5090 VSS.n2869 2.2505
R3794 VSS.n5089 VSS.n5088 2.2505
R3795 VSS.n5087 VSS.n2870 2.2505
R3796 VSS.n5086 VSS.n5085 2.2505
R3797 VSS.n5084 VSS.n2871 2.2505
R3798 VSS.n5083 VSS.n5082 2.2505
R3799 VSS.n5081 VSS.n2872 2.2505
R3800 VSS.n5080 VSS.n5079 2.2505
R3801 VSS.n5078 VSS.n2873 2.2505
R3802 VSS.n5077 VSS.n5076 2.2505
R3803 VSS.n5075 VSS.n2874 2.2505
R3804 VSS.n5074 VSS.n5073 2.2505
R3805 VSS.n5072 VSS.n2875 2.2505
R3806 VSS.n5071 VSS.n5070 2.2505
R3807 VSS.n5069 VSS.n2876 2.2505
R3808 VSS.n5068 VSS.n5067 2.2505
R3809 VSS.n5066 VSS.n2877 2.2505
R3810 VSS.n5065 VSS.n5064 2.2505
R3811 VSS.n5063 VSS.n2878 2.2505
R3812 VSS.n5062 VSS.n5061 2.2505
R3813 VSS.n5060 VSS.n2879 2.2505
R3814 VSS.n5059 VSS.n5058 2.2505
R3815 VSS.n5057 VSS.n2880 2.2505
R3816 VSS.n5056 VSS.n5055 2.2505
R3817 VSS.n5054 VSS.n2881 2.2505
R3818 VSS.n5053 VSS.n5052 2.2505
R3819 VSS.n5051 VSS.n2882 2.2505
R3820 VSS.n5050 VSS.n5049 2.2505
R3821 VSS.n5048 VSS.n2883 2.2505
R3822 VSS.n5047 VSS.n5046 2.2505
R3823 VSS.n5045 VSS.n2884 2.2505
R3824 VSS.n5044 VSS.n5043 2.2505
R3825 VSS.n5042 VSS.n2885 2.2505
R3826 VSS.n5041 VSS.n5040 2.2505
R3827 VSS.n5039 VSS.n2886 2.2505
R3828 VSS.n5038 VSS.n5037 2.2505
R3829 VSS.n5036 VSS.n2887 2.2505
R3830 VSS.n5035 VSS.n5034 2.2505
R3831 VSS.n5033 VSS.n2888 2.2505
R3832 VSS.n5032 VSS.n5031 2.2505
R3833 VSS.n5030 VSS.n2889 2.2505
R3834 VSS.n5029 VSS.n5028 2.2505
R3835 VSS.n5027 VSS.n2890 2.2505
R3836 VSS.n5026 VSS.n5025 2.2505
R3837 VSS.n5024 VSS.n2891 2.2505
R3838 VSS.n5023 VSS.n5022 2.2505
R3839 VSS.n5021 VSS.n2892 2.2505
R3840 VSS.n5020 VSS.n5019 2.2505
R3841 VSS.n5018 VSS.n2893 2.2505
R3842 VSS.n5017 VSS.n5016 2.2505
R3843 VSS.n5015 VSS.n2894 2.2505
R3844 VSS.n5014 VSS.n5013 2.2505
R3845 VSS.n5012 VSS.n2895 2.2505
R3846 VSS.n5011 VSS.n5010 2.2505
R3847 VSS.n5009 VSS.n2896 2.2505
R3848 VSS.n5008 VSS.n5007 2.2505
R3849 VSS.n5006 VSS.n2897 2.2505
R3850 VSS.n5005 VSS.n5004 2.2505
R3851 VSS.n5003 VSS.n2898 2.2505
R3852 VSS.n5002 VSS.n5001 2.2505
R3853 VSS.n5000 VSS.n2899 2.2505
R3854 VSS.n4999 VSS.n4998 2.2505
R3855 VSS.n4997 VSS.n2900 2.2505
R3856 VSS.n4996 VSS.n4995 2.2505
R3857 VSS.n4994 VSS.n2901 2.2505
R3858 VSS.n4993 VSS.n4992 2.2505
R3859 VSS.n4991 VSS.n2902 2.2505
R3860 VSS.n4990 VSS.n4989 2.2505
R3861 VSS.n4988 VSS.n2903 2.2505
R3862 VSS.n4987 VSS.n4986 2.2505
R3863 VSS.n4985 VSS.n2904 2.2505
R3864 VSS.n4984 VSS.n4983 2.2505
R3865 VSS.n4982 VSS.n2905 2.2505
R3866 VSS.n4981 VSS.n4980 2.2505
R3867 VSS.n4979 VSS.n2906 2.2505
R3868 VSS.n4978 VSS.n4977 2.2505
R3869 VSS.n4976 VSS.n2907 2.2505
R3870 VSS.n4975 VSS.n4974 2.2505
R3871 VSS.n4973 VSS.n2908 2.2505
R3872 VSS.n4972 VSS.n4971 2.2505
R3873 VSS.n4970 VSS.n2909 2.2505
R3874 VSS.n4969 VSS.n4968 2.2505
R3875 VSS.n4967 VSS.n2910 2.2505
R3876 VSS.n4966 VSS.n4965 2.2505
R3877 VSS.n4964 VSS.n2911 2.2505
R3878 VSS.n4963 VSS.n4962 2.2505
R3879 VSS.n4961 VSS.n2912 2.2505
R3880 VSS.n4960 VSS.n4959 2.2505
R3881 VSS.n4958 VSS.n2913 2.2505
R3882 VSS.n4957 VSS.n4956 2.2505
R3883 VSS.n4955 VSS.n2914 2.2505
R3884 VSS.n4954 VSS.n4953 2.2505
R3885 VSS.n4952 VSS.n2915 2.2505
R3886 VSS.n4951 VSS.n4950 2.2505
R3887 VSS.n4949 VSS.n2916 2.2505
R3888 VSS.n4948 VSS.n4947 2.2505
R3889 VSS.n4946 VSS.n2917 2.2505
R3890 VSS.n4945 VSS.n4944 2.2505
R3891 VSS.n4943 VSS.n2918 2.2505
R3892 VSS.n4942 VSS.n4941 2.2505
R3893 VSS.n4940 VSS.n2919 2.2505
R3894 VSS.n4939 VSS.n4938 2.2505
R3895 VSS.n4937 VSS.n2920 2.2505
R3896 VSS.n4936 VSS.n4935 2.2505
R3897 VSS.n4934 VSS.n2921 2.2505
R3898 VSS.n4933 VSS.n4932 2.2505
R3899 VSS.n4931 VSS.n2922 2.2505
R3900 VSS.n4930 VSS.n4929 2.2505
R3901 VSS.n4928 VSS.n2923 2.2505
R3902 VSS.n4927 VSS.n4926 2.2505
R3903 VSS.n4925 VSS.n2924 2.2505
R3904 VSS.n4924 VSS.n4923 2.2505
R3905 VSS.n4922 VSS.n2925 2.2505
R3906 VSS.n4921 VSS.n4920 2.2505
R3907 VSS.n4919 VSS.n2926 2.2505
R3908 VSS.n4918 VSS.n4917 2.2505
R3909 VSS.n4916 VSS.n2927 2.2505
R3910 VSS.n4915 VSS.n4914 2.2505
R3911 VSS.n4913 VSS.n2928 2.2505
R3912 VSS.n4912 VSS.n4911 2.2505
R3913 VSS.n4910 VSS.n2929 2.2505
R3914 VSS.n4909 VSS.n4908 2.2505
R3915 VSS.n4907 VSS.n2930 2.2505
R3916 VSS.n4906 VSS.n4905 2.2505
R3917 VSS.n4904 VSS.n2931 2.2505
R3918 VSS.n4903 VSS.n4902 2.2505
R3919 VSS.n4901 VSS.n2932 2.2505
R3920 VSS.n4900 VSS.n4899 2.2505
R3921 VSS.n4898 VSS.n2933 2.2505
R3922 VSS.n4897 VSS.n4896 2.2505
R3923 VSS.n4895 VSS.n2934 2.2505
R3924 VSS.n4894 VSS.n4893 2.2505
R3925 VSS.n4892 VSS.n2935 2.2505
R3926 VSS.n4891 VSS.n4890 2.2505
R3927 VSS.n4889 VSS.n2936 2.2505
R3928 VSS.n4888 VSS.n4887 2.2505
R3929 VSS.n4886 VSS.n2937 2.2505
R3930 VSS.n4885 VSS.n4884 2.2505
R3931 VSS.n4883 VSS.n2938 2.2505
R3932 VSS.n4882 VSS.n4881 2.2505
R3933 VSS.n4880 VSS.n2939 2.2505
R3934 VSS.n4879 VSS.n4878 2.2505
R3935 VSS.n4877 VSS.n2940 2.2505
R3936 VSS.n4876 VSS.n4875 2.2505
R3937 VSS.n4874 VSS.n2941 2.2505
R3938 VSS.n4873 VSS.n4872 2.2505
R3939 VSS.n4871 VSS.n2942 2.2505
R3940 VSS.n4870 VSS.n4869 2.2505
R3941 VSS.n4868 VSS.n2943 2.2505
R3942 VSS.n4867 VSS.n4866 2.2505
R3943 VSS.n4865 VSS.n2944 2.2505
R3944 VSS.n4864 VSS.n4863 2.2505
R3945 VSS.n4862 VSS.n2945 2.2505
R3946 VSS.n4861 VSS.n4860 2.2505
R3947 VSS.n4859 VSS.n2946 2.2505
R3948 VSS.n4858 VSS.n4857 2.2505
R3949 VSS.n4856 VSS.n2947 2.2505
R3950 VSS.n4855 VSS.n4854 2.2505
R3951 VSS.n4853 VSS.n2948 2.2505
R3952 VSS.n4852 VSS.n4851 2.2505
R3953 VSS.n4850 VSS.n2949 2.2505
R3954 VSS.n4849 VSS.n4848 2.2505
R3955 VSS.n4847 VSS.n2950 2.2505
R3956 VSS.n4846 VSS.n4845 2.2505
R3957 VSS.n4844 VSS.n2951 2.2505
R3958 VSS.n4843 VSS.n4842 2.2505
R3959 VSS.n4841 VSS.n2952 2.2505
R3960 VSS.n4840 VSS.n4839 2.2505
R3961 VSS.n4838 VSS.n2953 2.2505
R3962 VSS.n4837 VSS.n4836 2.2505
R3963 VSS.n4835 VSS.n2954 2.2505
R3964 VSS.n4834 VSS.n4833 2.2505
R3965 VSS.n4832 VSS.n2955 2.2505
R3966 VSS.n4831 VSS.n4830 2.2505
R3967 VSS.n4829 VSS.n2956 2.2505
R3968 VSS.n4828 VSS.n4827 2.2505
R3969 VSS.n4826 VSS.n2957 2.2505
R3970 VSS.n4825 VSS.n4824 2.2505
R3971 VSS.n4823 VSS.n2958 2.2505
R3972 VSS.n4822 VSS.n4821 2.2505
R3973 VSS.n4820 VSS.n2959 2.2505
R3974 VSS.n4819 VSS.n4818 2.2505
R3975 VSS.n4817 VSS.n2960 2.2505
R3976 VSS.n4816 VSS.n4815 2.2505
R3977 VSS.n4814 VSS.n2961 2.2505
R3978 VSS.n4813 VSS.n4812 2.2505
R3979 VSS.n4811 VSS.n2962 2.2505
R3980 VSS.n4810 VSS.n4809 2.2505
R3981 VSS.n4808 VSS.n2963 2.2505
R3982 VSS.n4807 VSS.n4806 2.2505
R3983 VSS.n4802 VSS.n2964 2.2505
R3984 VSS.n4801 VSS.n4800 2.2505
R3985 VSS.n4799 VSS.n2965 2.2505
R3986 VSS.n4798 VSS.n4797 2.2505
R3987 VSS.n4796 VSS.n2966 2.2505
R3988 VSS.n4795 VSS.n4794 2.2505
R3989 VSS.n4793 VSS.n2967 2.2505
R3990 VSS.n4792 VSS.n4791 2.2505
R3991 VSS.n4790 VSS.n2968 2.2505
R3992 VSS.n4789 VSS.n4788 2.2505
R3993 VSS.n4787 VSS.n2969 2.2505
R3994 VSS.n4786 VSS.n4785 2.2505
R3995 VSS.n4784 VSS.n2970 2.2505
R3996 VSS.n4783 VSS.n4782 2.2505
R3997 VSS.n4781 VSS.n2971 2.2505
R3998 VSS.n4780 VSS.n4779 2.2505
R3999 VSS.n4778 VSS.n2972 2.2505
R4000 VSS.n4777 VSS.n4776 2.2505
R4001 VSS.n4775 VSS.n2973 2.2505
R4002 VSS.n4774 VSS.n4773 2.2505
R4003 VSS.n4772 VSS.n2974 2.2505
R4004 VSS.n4771 VSS.n4770 2.2505
R4005 VSS.n4769 VSS.n2975 2.2505
R4006 VSS.n4768 VSS.n4767 2.2505
R4007 VSS.n4766 VSS.n2976 2.2505
R4008 VSS.n4765 VSS.n4764 2.2505
R4009 VSS.n4763 VSS.n2977 2.2505
R4010 VSS.n4762 VSS.n4761 2.2505
R4011 VSS.n4760 VSS.n2978 2.2505
R4012 VSS.n4759 VSS.n4758 2.2505
R4013 VSS.n4757 VSS.n2979 2.2505
R4014 VSS.n4756 VSS.n4755 2.2505
R4015 VSS.n4754 VSS.n2980 2.2505
R4016 VSS.n4753 VSS.n4752 2.2505
R4017 VSS.n4751 VSS.n2981 2.2505
R4018 VSS.n4750 VSS.n4749 2.2505
R4019 VSS.n4748 VSS.n2982 2.2505
R4020 VSS.n4747 VSS.n4746 2.2505
R4021 VSS.n4745 VSS.n2983 2.2505
R4022 VSS.n4744 VSS.n4743 2.2505
R4023 VSS.n4742 VSS.n2984 2.2505
R4024 VSS.n4741 VSS.n4740 2.2505
R4025 VSS.n4739 VSS.n2985 2.2505
R4026 VSS.n4738 VSS.n4737 2.2505
R4027 VSS.n4736 VSS.n2986 2.2505
R4028 VSS.n4735 VSS.n4734 2.2505
R4029 VSS.n4733 VSS.n2987 2.2505
R4030 VSS.n4732 VSS.n4731 2.2505
R4031 VSS.n4730 VSS.n2988 2.2505
R4032 VSS.n4729 VSS.n4728 2.2505
R4033 VSS.n4727 VSS.n2989 2.2505
R4034 VSS.n4726 VSS.n4725 2.2505
R4035 VSS.n4724 VSS.n2990 2.2505
R4036 VSS.n4723 VSS.n4722 2.2505
R4037 VSS.n4721 VSS.n2991 2.2505
R4038 VSS.n4720 VSS.n4719 2.2505
R4039 VSS.n4718 VSS.n2992 2.2505
R4040 VSS.n4717 VSS.n4716 2.2505
R4041 VSS.n4715 VSS.n2993 2.2505
R4042 VSS.n4714 VSS.n4713 2.2505
R4043 VSS.n4712 VSS.n2994 2.2505
R4044 VSS.n4711 VSS.n4710 2.2505
R4045 VSS.n4709 VSS.n2995 2.2505
R4046 VSS.n4708 VSS.n4707 2.2505
R4047 VSS.n4706 VSS.n2996 2.2505
R4048 VSS.n4705 VSS.n4704 2.2505
R4049 VSS.n4703 VSS.n2997 2.2505
R4050 VSS.n4702 VSS.n4701 2.2505
R4051 VSS.n4700 VSS.n2998 2.2505
R4052 VSS.n4699 VSS.n4698 2.2505
R4053 VSS.n4697 VSS.n2999 2.2505
R4054 VSS.n4696 VSS.n4695 2.2505
R4055 VSS.n4694 VSS.n3000 2.2505
R4056 VSS.n4693 VSS.n4692 2.2505
R4057 VSS.n4691 VSS.n3001 2.2505
R4058 VSS.n4690 VSS.n4689 2.2505
R4059 VSS.n4688 VSS.n3002 2.2505
R4060 VSS.n4687 VSS.n4686 2.2505
R4061 VSS.n4685 VSS.n3003 2.2505
R4062 VSS.n4684 VSS.n4683 2.2505
R4063 VSS.n4682 VSS.n3004 2.2505
R4064 VSS.n4681 VSS.n4680 2.2505
R4065 VSS.n4679 VSS.n3005 2.2505
R4066 VSS.n4678 VSS.n4677 2.2505
R4067 VSS.n4676 VSS.n3006 2.2505
R4068 VSS.n4675 VSS.n4674 2.2505
R4069 VSS.n4673 VSS.n3007 2.2505
R4070 VSS.n4672 VSS.n4671 2.2505
R4071 VSS.n4670 VSS.n3008 2.2505
R4072 VSS.n4669 VSS.n4668 2.2505
R4073 VSS.n4667 VSS.n3009 2.2505
R4074 VSS.n4666 VSS.n4665 2.2505
R4075 VSS.n4664 VSS.n3010 2.2505
R4076 VSS.n4663 VSS.n4662 2.2505
R4077 VSS.n4661 VSS.n3011 2.2505
R4078 VSS.n4660 VSS.n4659 2.2505
R4079 VSS.n4658 VSS.n3012 2.2505
R4080 VSS.n4657 VSS.n4656 2.2505
R4081 VSS.n4655 VSS.n3013 2.2505
R4082 VSS.n4654 VSS.n4653 2.2505
R4083 VSS.n4652 VSS.n3014 2.2505
R4084 VSS.n4651 VSS.n4650 2.2505
R4085 VSS.n4649 VSS.n3015 2.2505
R4086 VSS.n4648 VSS.n4647 2.2505
R4087 VSS.n4646 VSS.n3016 2.2505
R4088 VSS.n4645 VSS.n4644 2.2505
R4089 VSS.n4643 VSS.n3017 2.2505
R4090 VSS.n4642 VSS.n4641 2.2505
R4091 VSS.n4640 VSS.n3018 2.2505
R4092 VSS.n4639 VSS.n4638 2.2505
R4093 VSS.n4637 VSS.n3019 2.2505
R4094 VSS.n4636 VSS.n4635 2.2505
R4095 VSS.n4634 VSS.n3020 2.2505
R4096 VSS.n4633 VSS.n4632 2.2505
R4097 VSS.n4631 VSS.n3021 2.2505
R4098 VSS.n4630 VSS.n4629 2.2505
R4099 VSS.n4628 VSS.n3022 2.2505
R4100 VSS.n4627 VSS.n4626 2.2505
R4101 VSS.n4625 VSS.n3023 2.2505
R4102 VSS.n4624 VSS.n4623 2.2505
R4103 VSS.n4622 VSS.n3024 2.2505
R4104 VSS.n4621 VSS.n4620 2.2505
R4105 VSS.n4619 VSS.n3025 2.2505
R4106 VSS.n4618 VSS.n4617 2.2505
R4107 VSS.n4616 VSS.n3026 2.2505
R4108 VSS.n4615 VSS.n4614 2.2505
R4109 VSS.n4613 VSS.n3027 2.2505
R4110 VSS.n4612 VSS.n4611 2.2505
R4111 VSS.n4610 VSS.n3028 2.2505
R4112 VSS.n4609 VSS.n4608 2.2505
R4113 VSS.n4607 VSS.n3029 2.2505
R4114 VSS.n4606 VSS.n4605 2.2505
R4115 VSS.n4604 VSS.n3030 2.2505
R4116 VSS.n4603 VSS.n4602 2.2505
R4117 VSS.n4601 VSS.n3031 2.2505
R4118 VSS.n4600 VSS.n4599 2.2505
R4119 VSS.n4598 VSS.n3032 2.2505
R4120 VSS.n4597 VSS.n4596 2.2505
R4121 VSS.n4595 VSS.n3033 2.2505
R4122 VSS.n4594 VSS.n4593 2.2505
R4123 VSS.n4592 VSS.n3034 2.2505
R4124 VSS.n4591 VSS.n4590 2.2505
R4125 VSS.n4589 VSS.n3035 2.2505
R4126 VSS.n4588 VSS.n4587 2.2505
R4127 VSS.n4586 VSS.n3036 2.2505
R4128 VSS.n4585 VSS.n4584 2.2505
R4129 VSS.n4583 VSS.n3037 2.2505
R4130 VSS.n4582 VSS.n4581 2.2505
R4131 VSS.n4580 VSS.n3038 2.2505
R4132 VSS.n4579 VSS.n4578 2.2505
R4133 VSS.n4577 VSS.n3039 2.2505
R4134 VSS.n4576 VSS.n4575 2.2505
R4135 VSS.n4574 VSS.n3040 2.2505
R4136 VSS.n4573 VSS.n4572 2.2505
R4137 VSS.n4571 VSS.n3041 2.2505
R4138 VSS.n4570 VSS.n4569 2.2505
R4139 VSS.n4568 VSS.n3042 2.2505
R4140 VSS.n4567 VSS.n4566 2.2505
R4141 VSS.n4565 VSS.n3043 2.2505
R4142 VSS.n4564 VSS.n4563 2.2505
R4143 VSS.n4562 VSS.n3044 2.2505
R4144 VSS.n4561 VSS.n4560 2.2505
R4145 VSS.n4559 VSS.n3045 2.2505
R4146 VSS.n4558 VSS.n4557 2.2505
R4147 VSS.n4556 VSS.n3046 2.2505
R4148 VSS.n4555 VSS.n4554 2.2505
R4149 VSS.n4553 VSS.n3047 2.2505
R4150 VSS.n4552 VSS.n4551 2.2505
R4151 VSS.n4550 VSS.n3048 2.2505
R4152 VSS.n4549 VSS.n4548 2.2505
R4153 VSS.n4547 VSS.n3049 2.2505
R4154 VSS.n4546 VSS.n4545 2.2505
R4155 VSS.n4544 VSS.n3050 2.2505
R4156 VSS.n4543 VSS.n4542 2.2505
R4157 VSS.n4541 VSS.n3051 2.2505
R4158 VSS.n4540 VSS.n4539 2.2505
R4159 VSS.n4538 VSS.n3052 2.2505
R4160 VSS.n4537 VSS.n4536 2.2505
R4161 VSS.n4535 VSS.n3053 2.2505
R4162 VSS.n4534 VSS.n4533 2.2505
R4163 VSS.n4532 VSS.n3054 2.2505
R4164 VSS.n4531 VSS.n4530 2.2505
R4165 VSS.n4529 VSS.n3055 2.2505
R4166 VSS.n4528 VSS.n4527 2.2505
R4167 VSS.n4526 VSS.n3056 2.2505
R4168 VSS.n4525 VSS.n4524 2.2505
R4169 VSS.n4523 VSS.n3057 2.2505
R4170 VSS.n4522 VSS.n4521 2.2505
R4171 VSS.n4520 VSS.n3058 2.2505
R4172 VSS.n4519 VSS.n4518 2.2505
R4173 VSS.n4517 VSS.n3059 2.2505
R4174 VSS.n4516 VSS.n4515 2.2505
R4175 VSS.n4514 VSS.n3060 2.2505
R4176 VSS.n4513 VSS.n4512 2.2505
R4177 VSS.n4511 VSS.n3061 2.2505
R4178 VSS.n4510 VSS.n4509 2.2505
R4179 VSS.n4508 VSS.n3062 2.2505
R4180 VSS.n4507 VSS.n4506 2.2505
R4181 VSS.n4505 VSS.n3063 2.2505
R4182 VSS.n4504 VSS.n4503 2.2505
R4183 VSS.n4502 VSS.n3064 2.2505
R4184 VSS.n4501 VSS.n4500 2.2505
R4185 VSS.n4499 VSS.n3065 2.2505
R4186 VSS.n4498 VSS.n4497 2.2505
R4187 VSS.n4496 VSS.n3066 2.2505
R4188 VSS.n4495 VSS.n4494 2.2505
R4189 VSS.n4493 VSS.n3067 2.2505
R4190 VSS.n4492 VSS.n4491 2.2505
R4191 VSS.n4490 VSS.n3068 2.2505
R4192 VSS.n4489 VSS.n4488 2.2505
R4193 VSS.n4487 VSS.n3069 2.2505
R4194 VSS.n4486 VSS.n4485 2.2505
R4195 VSS.n4484 VSS.n3070 2.2505
R4196 VSS.n4483 VSS.n4482 2.2505
R4197 VSS.n4481 VSS.n3071 2.2505
R4198 VSS.n4480 VSS.n4479 2.2505
R4199 VSS.n4478 VSS.n3072 2.2505
R4200 VSS.n4477 VSS.n4476 2.2505
R4201 VSS.n4475 VSS.n3073 2.2505
R4202 VSS.n4474 VSS.n4473 2.2505
R4203 VSS.n4472 VSS.n3074 2.2505
R4204 VSS.n4471 VSS.n4470 2.2505
R4205 VSS.n4469 VSS.n3075 2.2505
R4206 VSS.n4468 VSS.n4467 2.2505
R4207 VSS.n4466 VSS.n3076 2.2505
R4208 VSS.n4465 VSS.n4464 2.2505
R4209 VSS.n4463 VSS.n3077 2.2505
R4210 VSS.n4462 VSS.n4461 2.2505
R4211 VSS.n4460 VSS.n3078 2.2505
R4212 VSS.n4459 VSS.n4458 2.2505
R4213 VSS.n4457 VSS.n3079 2.2505
R4214 VSS.n4456 VSS.n4455 2.2505
R4215 VSS.n4454 VSS.n3080 2.2505
R4216 VSS.n4453 VSS.n4452 2.2505
R4217 VSS.n4451 VSS.n3081 2.2505
R4218 VSS.n4450 VSS.n4449 2.2505
R4219 VSS.n4448 VSS.n3082 2.2505
R4220 VSS.n4447 VSS.n4446 2.2505
R4221 VSS.n4445 VSS.n3083 2.2505
R4222 VSS.n4444 VSS.n4443 2.2505
R4223 VSS.n4442 VSS.n3084 2.2505
R4224 VSS.n4441 VSS.n4440 2.2505
R4225 VSS.n4439 VSS.n3085 2.2505
R4226 VSS.n4438 VSS.n4437 2.2505
R4227 VSS.n4436 VSS.n3086 2.2505
R4228 VSS.n4435 VSS.n4434 2.2505
R4229 VSS.n4433 VSS.n3087 2.2505
R4230 VSS.n4432 VSS.n4431 2.2505
R4231 VSS.n4430 VSS.n3088 2.2505
R4232 VSS.n4429 VSS.n4428 2.2505
R4233 VSS.n4427 VSS.n3089 2.2505
R4234 VSS.n4426 VSS.n4425 2.2505
R4235 VSS.n4424 VSS.n3090 2.2505
R4236 VSS.n4423 VSS.n4422 2.2505
R4237 VSS.n4421 VSS.n3091 2.2505
R4238 VSS.n4420 VSS.n4419 2.2505
R4239 VSS.n4418 VSS.n3092 2.2505
R4240 VSS.n4417 VSS.n4416 2.2505
R4241 VSS.n4415 VSS.n3093 2.2505
R4242 VSS.n4414 VSS.n4413 2.2505
R4243 VSS.n4412 VSS.n3094 2.2505
R4244 VSS.n4411 VSS.n4410 2.2505
R4245 VSS.n4409 VSS.n3095 2.2505
R4246 VSS.n4408 VSS.n4407 2.2505
R4247 VSS.n4406 VSS.n3096 2.2505
R4248 VSS.n4405 VSS.n4404 2.2505
R4249 VSS.n4403 VSS.n3097 2.2505
R4250 VSS.n4402 VSS.n4401 2.2505
R4251 VSS.n4400 VSS.n3098 2.2505
R4252 VSS.n4399 VSS.n4398 2.2505
R4253 VSS.n4397 VSS.n3099 2.2505
R4254 VSS.n4396 VSS.n4395 2.2505
R4255 VSS.n4394 VSS.n3100 2.2505
R4256 VSS.n4393 VSS.n4392 2.2505
R4257 VSS.n4391 VSS.n3101 2.2505
R4258 VSS.n4390 VSS.n4389 2.2505
R4259 VSS.n4388 VSS.n3102 2.2505
R4260 VSS.n4387 VSS.n4386 2.2505
R4261 VSS.n4385 VSS.n3103 2.2505
R4262 VSS.n4384 VSS.n4383 2.2505
R4263 VSS.n4382 VSS.n3104 2.2505
R4264 VSS.n4381 VSS.n4380 2.2505
R4265 VSS.n4379 VSS.n3105 2.2505
R4266 VSS.n4378 VSS.n4377 2.2505
R4267 VSS.n4376 VSS.n3106 2.2505
R4268 VSS.n4375 VSS.n4374 2.2505
R4269 VSS.n4373 VSS.n3107 2.2505
R4270 VSS.n4372 VSS.n4371 2.2505
R4271 VSS.n4370 VSS.n3108 2.2505
R4272 VSS.n4369 VSS.n4368 2.2505
R4273 VSS.n4367 VSS.n3109 2.2505
R4274 VSS.n4366 VSS.n4365 2.2505
R4275 VSS.n4364 VSS.n3110 2.2505
R4276 VSS.n4363 VSS.n4362 2.2505
R4277 VSS.n4361 VSS.n3111 2.2505
R4278 VSS.n4360 VSS.n4359 2.2505
R4279 VSS.n4358 VSS.n3112 2.2505
R4280 VSS.n4357 VSS.n4356 2.2505
R4281 VSS.n4355 VSS.n3113 2.2505
R4282 VSS.n4354 VSS.n4353 2.2505
R4283 VSS.n4352 VSS.n3114 2.2505
R4284 VSS.n4351 VSS.n4350 2.2505
R4285 VSS.n4349 VSS.n3115 2.2505
R4286 VSS.n4348 VSS.n4347 2.2505
R4287 VSS.n4346 VSS.n3116 2.2505
R4288 VSS.n4345 VSS.n4344 2.2505
R4289 VSS.n4343 VSS.n3117 2.2505
R4290 VSS.n4342 VSS.n4341 2.2505
R4291 VSS.n4340 VSS.n3118 2.2505
R4292 VSS.n4339 VSS.n4338 2.2505
R4293 VSS.n4337 VSS.n3119 2.2505
R4294 VSS.n4336 VSS.n4335 2.2505
R4295 VSS.n4334 VSS.n3120 2.2505
R4296 VSS.n4333 VSS.n4332 2.2505
R4297 VSS.n4331 VSS.n3121 2.2505
R4298 VSS.n4330 VSS.n4329 2.2505
R4299 VSS.n4328 VSS.n3122 2.2505
R4300 VSS.n4327 VSS.n4326 2.2505
R4301 VSS.n4325 VSS.n3123 2.2505
R4302 VSS.n4324 VSS.n4323 2.2505
R4303 VSS.n4322 VSS.n3124 2.2505
R4304 VSS.n4321 VSS.n4320 2.2505
R4305 VSS.n4319 VSS.n3125 2.2505
R4306 VSS.n4318 VSS.n4317 2.2505
R4307 VSS.n4316 VSS.n3126 2.2505
R4308 VSS.n4315 VSS.n4314 2.2505
R4309 VSS.n4313 VSS.n3127 2.2505
R4310 VSS.n4312 VSS.n4311 2.2505
R4311 VSS.n4310 VSS.n3128 2.2505
R4312 VSS.n4309 VSS.n4308 2.2505
R4313 VSS.n4307 VSS.n3129 2.2505
R4314 VSS.n4306 VSS.n4305 2.2505
R4315 VSS.n4304 VSS.n3130 2.2505
R4316 VSS.n4303 VSS.n4302 2.2505
R4317 VSS.n4301 VSS.n3131 2.2505
R4318 VSS.n4300 VSS.n4299 2.2505
R4319 VSS.n4298 VSS.n3132 2.2505
R4320 VSS.n4297 VSS.n4296 2.2505
R4321 VSS.n4295 VSS.n3133 2.2505
R4322 VSS.n4294 VSS.n4293 2.2505
R4323 VSS.n4292 VSS.n3134 2.2505
R4324 VSS.n4291 VSS.n4290 2.2505
R4325 VSS.n4289 VSS.n3135 2.2505
R4326 VSS.n4288 VSS.n4287 2.2505
R4327 VSS.n4286 VSS.n3136 2.2505
R4328 VSS.n4285 VSS.n4284 2.2505
R4329 VSS.n4283 VSS.n3137 2.2505
R4330 VSS.n4282 VSS.n4281 2.2505
R4331 VSS.n4280 VSS.n3138 2.2505
R4332 VSS.n4279 VSS.n4278 2.2505
R4333 VSS.n4277 VSS.n3139 2.2505
R4334 VSS.n4276 VSS.n4275 2.2505
R4335 VSS.n4274 VSS.n3140 2.2505
R4336 VSS.n4273 VSS.n4272 2.2505
R4337 VSS.n4271 VSS.n3141 2.2505
R4338 VSS.n4270 VSS.n4269 2.2505
R4339 VSS.n4268 VSS.n3142 2.2505
R4340 VSS.n4267 VSS.n4266 2.2505
R4341 VSS.n4265 VSS.n3143 2.2505
R4342 VSS.n4264 VSS.n4263 2.2505
R4343 VSS.n4262 VSS.n3144 2.2505
R4344 VSS.n4261 VSS.n4260 2.2505
R4345 VSS.n4259 VSS.n3145 2.2505
R4346 VSS.n4258 VSS.n4257 2.2505
R4347 VSS.n4256 VSS.n3146 2.2505
R4348 VSS.n4255 VSS.n4254 2.2505
R4349 VSS.n4253 VSS.n3147 2.2505
R4350 VSS.n4252 VSS.n4251 2.2505
R4351 VSS.n4250 VSS.n3148 2.2505
R4352 VSS.n4249 VSS.n4248 2.2505
R4353 VSS.n4247 VSS.n3149 2.2505
R4354 VSS.n4246 VSS.n4245 2.2505
R4355 VSS.n4244 VSS.n3150 2.2505
R4356 VSS.n4243 VSS.n4242 2.2505
R4357 VSS.n4241 VSS.n3151 2.2505
R4358 VSS.n4240 VSS.n4239 2.2505
R4359 VSS.n4238 VSS.n3152 2.2505
R4360 VSS.n4237 VSS.n4236 2.2505
R4361 VSS.n4235 VSS.n3153 2.2505
R4362 VSS.n4234 VSS.n4233 2.2505
R4363 VSS.n4232 VSS.n3154 2.2505
R4364 VSS.n4231 VSS.n4230 2.2505
R4365 VSS.n4229 VSS.n3155 2.2505
R4366 VSS.n4228 VSS.n4227 2.2505
R4367 VSS.n4226 VSS.n3156 2.2505
R4368 VSS.n4225 VSS.n4224 2.2505
R4369 VSS.n4223 VSS.n3157 2.2505
R4370 VSS.n4222 VSS.n4221 2.2505
R4371 VSS.n4220 VSS.n3158 2.2505
R4372 VSS.n4219 VSS.n4218 2.2505
R4373 VSS.n4217 VSS.n3159 2.2505
R4374 VSS.n4216 VSS.n4215 2.2505
R4375 VSS.n4214 VSS.n3160 2.2505
R4376 VSS.n4213 VSS.n4212 2.2505
R4377 VSS.n4211 VSS.n3161 2.2505
R4378 VSS.n4210 VSS.n4209 2.2505
R4379 VSS.n4208 VSS.n3162 2.2505
R4380 VSS.n4207 VSS.n4206 2.2505
R4381 VSS.n4205 VSS.n3163 2.2505
R4382 VSS.n4204 VSS.n4203 2.2505
R4383 VSS.n4202 VSS.n3164 2.2505
R4384 VSS.n4201 VSS.n4200 2.2505
R4385 VSS.n4199 VSS.n3165 2.2505
R4386 VSS.n4198 VSS.n4197 2.2505
R4387 VSS.n4196 VSS.n3166 2.2505
R4388 VSS.n4195 VSS.n4194 2.2505
R4389 VSS.n4193 VSS.n3167 2.2505
R4390 VSS.n4192 VSS.n4191 2.2505
R4391 VSS.n4190 VSS.n3168 2.2505
R4392 VSS.n4189 VSS.n4188 2.2505
R4393 VSS.n4187 VSS.n3169 2.2505
R4394 VSS.n4186 VSS.n4185 2.2505
R4395 VSS.n4184 VSS.n3170 2.2505
R4396 VSS.n4183 VSS.n4182 2.2505
R4397 VSS.n4181 VSS.n3171 2.2505
R4398 VSS.n4180 VSS.n4179 2.2505
R4399 VSS.n4178 VSS.n3172 2.2505
R4400 VSS.n4177 VSS.n4176 2.2505
R4401 VSS.n4175 VSS.n3173 2.2505
R4402 VSS.n4174 VSS.n4173 2.2505
R4403 VSS.n4172 VSS.n3174 2.2505
R4404 VSS.n4171 VSS.n4170 2.2505
R4405 VSS.n4169 VSS.n3175 2.2505
R4406 VSS.n4168 VSS.n4167 2.2505
R4407 VSS.n4166 VSS.n3176 2.2505
R4408 VSS.n4165 VSS.n4164 2.2505
R4409 VSS.n4163 VSS.n3177 2.2505
R4410 VSS.n4162 VSS.n4161 2.2505
R4411 VSS.n4160 VSS.n3178 2.2505
R4412 VSS.n4159 VSS.n4158 2.2505
R4413 VSS.n4157 VSS.n3179 2.2505
R4414 VSS.n4156 VSS.n4155 2.2505
R4415 VSS.n4154 VSS.n3180 2.2505
R4416 VSS.n4153 VSS.n4152 2.2505
R4417 VSS.n4151 VSS.n3181 2.2505
R4418 VSS.n4150 VSS.n4149 2.2505
R4419 VSS.n4148 VSS.n3182 2.2505
R4420 VSS.n4147 VSS.n4146 2.2505
R4421 VSS.n4145 VSS.n3183 2.2505
R4422 VSS.n4144 VSS.n4143 2.2505
R4423 VSS.n4142 VSS.n3184 2.2505
R4424 VSS.n6907 VSS.n6906 2.2505
R4425 VSS.n6905 VSS.n2264 2.2505
R4426 VSS.n6904 VSS.n6903 2.2505
R4427 VSS.n6902 VSS.n2265 2.2505
R4428 VSS.n6901 VSS.n6900 2.2505
R4429 VSS.n6899 VSS.n2266 2.2505
R4430 VSS.n6898 VSS.n6897 2.2505
R4431 VSS.n6896 VSS.n2267 2.2505
R4432 VSS.n6895 VSS.n6894 2.2505
R4433 VSS.n6893 VSS.n2268 2.2505
R4434 VSS.n6892 VSS.n6891 2.2505
R4435 VSS.n6890 VSS.n2269 2.2505
R4436 VSS.n6889 VSS.n6888 2.2505
R4437 VSS.n6887 VSS.n2270 2.2505
R4438 VSS.n6886 VSS.n6885 2.2505
R4439 VSS.n6884 VSS.n2271 2.2505
R4440 VSS.n6883 VSS.n6882 2.2505
R4441 VSS.n6881 VSS.n2272 2.2505
R4442 VSS.n6880 VSS.n6879 2.2505
R4443 VSS.n6878 VSS.n2273 2.2505
R4444 VSS.n6877 VSS.n6876 2.2505
R4445 VSS.n6875 VSS.n2274 2.2505
R4446 VSS.n6874 VSS.n6873 2.2505
R4447 VSS.n6872 VSS.n2275 2.2505
R4448 VSS.n6871 VSS.n6870 2.2505
R4449 VSS.n6869 VSS.n2276 2.2505
R4450 VSS.n6868 VSS.n6867 2.2505
R4451 VSS.n6866 VSS.n2277 2.2505
R4452 VSS.n6865 VSS.n6864 2.2505
R4453 VSS.n6863 VSS.n2278 2.2505
R4454 VSS.n6862 VSS.n6861 2.2505
R4455 VSS.n6860 VSS.n2279 2.2505
R4456 VSS.n6859 VSS.n6858 2.2505
R4457 VSS.n6857 VSS.n2280 2.2505
R4458 VSS.n6856 VSS.n6855 2.2505
R4459 VSS.n6854 VSS.n2281 2.2505
R4460 VSS.n6853 VSS.n6852 2.2505
R4461 VSS.n6851 VSS.n2282 2.2505
R4462 VSS.n6850 VSS.n6849 2.2505
R4463 VSS.n6848 VSS.n2283 2.2505
R4464 VSS.n6847 VSS.n6846 2.2505
R4465 VSS.n6845 VSS.n2284 2.2505
R4466 VSS.n6844 VSS.n6843 2.2505
R4467 VSS.n6842 VSS.n2285 2.2505
R4468 VSS.n6841 VSS.n6840 2.2505
R4469 VSS.n6839 VSS.n2286 2.2505
R4470 VSS.n6838 VSS.n6837 2.2505
R4471 VSS.n6836 VSS.n2287 2.2505
R4472 VSS.n6835 VSS.n6834 2.2505
R4473 VSS.n6833 VSS.n2288 2.2505
R4474 VSS.n6832 VSS.n6831 2.2505
R4475 VSS.n6830 VSS.n2289 2.2505
R4476 VSS.n6829 VSS.n6828 2.2505
R4477 VSS.n6827 VSS.n2290 2.2505
R4478 VSS.n6826 VSS.n6825 2.2505
R4479 VSS.n6824 VSS.n2291 2.2505
R4480 VSS.n6823 VSS.n6822 2.2505
R4481 VSS.n6821 VSS.n2292 2.2505
R4482 VSS.n6820 VSS.n6819 2.2505
R4483 VSS.n6818 VSS.n2293 2.2505
R4484 VSS.n6817 VSS.n6816 2.2505
R4485 VSS.n6815 VSS.n2294 2.2505
R4486 VSS.n6814 VSS.n6813 2.2505
R4487 VSS.n6812 VSS.n2295 2.2505
R4488 VSS.n6811 VSS.n6810 2.2505
R4489 VSS.n6809 VSS.n2296 2.2505
R4490 VSS.n6808 VSS.n6807 2.2505
R4491 VSS.n6806 VSS.n2297 2.2505
R4492 VSS.n6805 VSS.n6804 2.2505
R4493 VSS.n6803 VSS.n2298 2.2505
R4494 VSS.n6802 VSS.n6801 2.2505
R4495 VSS.n6800 VSS.n2299 2.2505
R4496 VSS.n6799 VSS.n6798 2.2505
R4497 VSS.n6797 VSS.n2300 2.2505
R4498 VSS.n6796 VSS.n6795 2.2505
R4499 VSS.n6794 VSS.n2301 2.2505
R4500 VSS.n6793 VSS.n6792 2.2505
R4501 VSS.n6791 VSS.n2302 2.2505
R4502 VSS.n6790 VSS.n6789 2.2505
R4503 VSS.n6788 VSS.n2303 2.2505
R4504 VSS.n6787 VSS.n6786 2.2505
R4505 VSS.n6785 VSS.n2304 2.2505
R4506 VSS.n6784 VSS.n6783 2.2505
R4507 VSS.n6782 VSS.n2305 2.2505
R4508 VSS.n6781 VSS.n6780 2.2505
R4509 VSS.n6779 VSS.n2306 2.2505
R4510 VSS.n6778 VSS.n6777 2.2505
R4511 VSS.n6776 VSS.n2307 2.2505
R4512 VSS.n6775 VSS.n6774 2.2505
R4513 VSS.n6773 VSS.n2308 2.2505
R4514 VSS.n6772 VSS.n6771 2.2505
R4515 VSS.n6770 VSS.n2309 2.2505
R4516 VSS.n6769 VSS.n6768 2.2505
R4517 VSS.n6767 VSS.n2310 2.2505
R4518 VSS.n6766 VSS.n6765 2.2505
R4519 VSS.n6764 VSS.n2311 2.2505
R4520 VSS.n6763 VSS.n6762 2.2505
R4521 VSS.n6761 VSS.n2312 2.2505
R4522 VSS.n6760 VSS.n6759 2.2505
R4523 VSS.n6758 VSS.n2313 2.2505
R4524 VSS.n6757 VSS.n6756 2.2505
R4525 VSS.n6755 VSS.n2314 2.2505
R4526 VSS.n6754 VSS.n6753 2.2505
R4527 VSS.n6752 VSS.n2315 2.2505
R4528 VSS.n6751 VSS.n6750 2.2505
R4529 VSS.n6749 VSS.n2316 2.2505
R4530 VSS.n6748 VSS.n6747 2.2505
R4531 VSS.n6746 VSS.n2317 2.2505
R4532 VSS.n6745 VSS.n6744 2.2505
R4533 VSS.n6743 VSS.n2318 2.2505
R4534 VSS.n6742 VSS.n6741 2.2505
R4535 VSS.n6740 VSS.n2319 2.2505
R4536 VSS.n6739 VSS.n6738 2.2505
R4537 VSS.n6737 VSS.n2320 2.2505
R4538 VSS.n6736 VSS.n6735 2.2505
R4539 VSS.n6734 VSS.n2321 2.2505
R4540 VSS.n6733 VSS.n6732 2.2505
R4541 VSS.n6731 VSS.n2322 2.2505
R4542 VSS.n6730 VSS.n6729 2.2505
R4543 VSS.n6728 VSS.n2323 2.2505
R4544 VSS.n6727 VSS.n6726 2.2505
R4545 VSS.n6725 VSS.n2324 2.2505
R4546 VSS.n6724 VSS.n6723 2.2505
R4547 VSS.n6722 VSS.n2325 2.2505
R4548 VSS.n6721 VSS.n6720 2.2505
R4549 VSS.n6719 VSS.n2326 2.2505
R4550 VSS.n6718 VSS.n6717 2.2505
R4551 VSS.n6716 VSS.n2327 2.2505
R4552 VSS.n6715 VSS.n6714 2.2505
R4553 VSS.n6713 VSS.n2328 2.2505
R4554 VSS.n6712 VSS.n6711 2.2505
R4555 VSS.n6710 VSS.n2329 2.2505
R4556 VSS.n6709 VSS.n6708 2.2505
R4557 VSS.n6707 VSS.n2330 2.2505
R4558 VSS.n6706 VSS.n6705 2.2505
R4559 VSS.n6704 VSS.n2331 2.2505
R4560 VSS.n6703 VSS.n6702 2.2505
R4561 VSS.n6701 VSS.n2332 2.2505
R4562 VSS.n6700 VSS.n6699 2.2505
R4563 VSS.n6698 VSS.n2333 2.2505
R4564 VSS.n6697 VSS.n6696 2.2505
R4565 VSS.n6695 VSS.n2334 2.2505
R4566 VSS.n6694 VSS.n6693 2.2505
R4567 VSS.n6692 VSS.n2335 2.2505
R4568 VSS.n6691 VSS.n6690 2.2505
R4569 VSS.n6689 VSS.n2336 2.2505
R4570 VSS.n6688 VSS.n6687 2.2505
R4571 VSS.n6686 VSS.n2337 2.2505
R4572 VSS.n6685 VSS.n6684 2.2505
R4573 VSS.n6683 VSS.n2338 2.2505
R4574 VSS.n6682 VSS.n6681 2.2505
R4575 VSS.n6680 VSS.n2339 2.2505
R4576 VSS.n6679 VSS.n6678 2.2505
R4577 VSS.n6677 VSS.n2340 2.2505
R4578 VSS.n6676 VSS.n6675 2.2505
R4579 VSS.n6674 VSS.n2341 2.2505
R4580 VSS.n6673 VSS.n6672 2.2505
R4581 VSS.n6671 VSS.n2342 2.2505
R4582 VSS.n6670 VSS.n6669 2.2505
R4583 VSS.n6668 VSS.n2343 2.2505
R4584 VSS.n6667 VSS.n6666 2.2505
R4585 VSS.n6665 VSS.n2344 2.2505
R4586 VSS.n6664 VSS.n6663 2.2505
R4587 VSS.n6662 VSS.n2345 2.2505
R4588 VSS.n6661 VSS.n6660 2.2505
R4589 VSS.n6659 VSS.n2346 2.2505
R4590 VSS.n6658 VSS.n6657 2.2505
R4591 VSS.n6656 VSS.n2347 2.2505
R4592 VSS.n6655 VSS.n6654 2.2505
R4593 VSS.n6653 VSS.n2348 2.2505
R4594 VSS.n6652 VSS.n6651 2.2505
R4595 VSS.n6650 VSS.n2349 2.2505
R4596 VSS.n6649 VSS.n6648 2.2505
R4597 VSS.n6647 VSS.n2350 2.2505
R4598 VSS.n6646 VSS.n6645 2.2505
R4599 VSS.n6644 VSS.n2351 2.2505
R4600 VSS.n6643 VSS.n6642 2.2505
R4601 VSS.n6641 VSS.n2352 2.2505
R4602 VSS.n6640 VSS.n6639 2.2505
R4603 VSS.n6638 VSS.n2353 2.2505
R4604 VSS.n6637 VSS.n6636 2.2505
R4605 VSS.n6635 VSS.n2354 2.2505
R4606 VSS.n6634 VSS.n6633 2.2505
R4607 VSS.n6632 VSS.n2355 2.2505
R4608 VSS.n6631 VSS.n6630 2.2505
R4609 VSS.n6629 VSS.n2356 2.2505
R4610 VSS.n6628 VSS.n6627 2.2505
R4611 VSS.n6626 VSS.n2357 2.2505
R4612 VSS.n6625 VSS.n6624 2.2505
R4613 VSS.n6623 VSS.n2358 2.2505
R4614 VSS.n6622 VSS.n6621 2.2505
R4615 VSS.n6620 VSS.n2359 2.2505
R4616 VSS.n6619 VSS.n6618 2.2505
R4617 VSS.n6617 VSS.n2360 2.2505
R4618 VSS.n6616 VSS.n6615 2.2505
R4619 VSS.n6614 VSS.n2361 2.2505
R4620 VSS.n6613 VSS.n6612 2.2505
R4621 VSS.n6611 VSS.n2362 2.2505
R4622 VSS.n6610 VSS.n6609 2.2505
R4623 VSS.n6608 VSS.n2363 2.2505
R4624 VSS.n6607 VSS.n6606 2.2505
R4625 VSS.n6605 VSS.n2364 2.2505
R4626 VSS.n6604 VSS.n6603 2.2505
R4627 VSS.n6602 VSS.n2365 2.2505
R4628 VSS.n6601 VSS.n6600 2.2505
R4629 VSS.n6599 VSS.n2366 2.2505
R4630 VSS.n6598 VSS.n6597 2.2505
R4631 VSS.n6596 VSS.n2367 2.2505
R4632 VSS.n6595 VSS.n6594 2.2505
R4633 VSS.n6593 VSS.n2368 2.2505
R4634 VSS.n6592 VSS.n6591 2.2505
R4635 VSS.n6590 VSS.n2369 2.2505
R4636 VSS.n6589 VSS.n6588 2.2505
R4637 VSS.n6587 VSS.n2370 2.2505
R4638 VSS.n6586 VSS.n6585 2.2505
R4639 VSS.n6584 VSS.n2371 2.2505
R4640 VSS.n6583 VSS.n6582 2.2505
R4641 VSS.n6581 VSS.n2372 2.2505
R4642 VSS.n6580 VSS.n6579 2.2505
R4643 VSS.n6578 VSS.n2373 2.2505
R4644 VSS.n6577 VSS.n6576 2.2505
R4645 VSS.n6575 VSS.n2374 2.2505
R4646 VSS.n6574 VSS.n6573 2.2505
R4647 VSS.n6572 VSS.n2375 2.2505
R4648 VSS.n6571 VSS.n6570 2.2505
R4649 VSS.n6569 VSS.n2376 2.2505
R4650 VSS.n6568 VSS.n6567 2.2505
R4651 VSS.n6566 VSS.n2377 2.2505
R4652 VSS.n6565 VSS.n6564 2.2505
R4653 VSS.n6563 VSS.n2378 2.2505
R4654 VSS.n6562 VSS.n6561 2.2505
R4655 VSS.n6560 VSS.n2379 2.2505
R4656 VSS.n6559 VSS.n6558 2.2505
R4657 VSS.n6557 VSS.n2380 2.2505
R4658 VSS.n6556 VSS.n6555 2.2505
R4659 VSS.n6554 VSS.n2381 2.2505
R4660 VSS.n6553 VSS.n6552 2.2505
R4661 VSS.n6551 VSS.n2382 2.2505
R4662 VSS.n6550 VSS.n6549 2.2505
R4663 VSS.n6548 VSS.n2383 2.2505
R4664 VSS.n6547 VSS.n6546 2.2505
R4665 VSS.n6545 VSS.n2384 2.2505
R4666 VSS.n6544 VSS.n6543 2.2505
R4667 VSS.n6542 VSS.n2385 2.2505
R4668 VSS.n6541 VSS.n6540 2.2505
R4669 VSS.n6539 VSS.n2386 2.2505
R4670 VSS.n6538 VSS.n6537 2.2505
R4671 VSS.n6536 VSS.n2387 2.2505
R4672 VSS.n6535 VSS.n6534 2.2505
R4673 VSS.n6533 VSS.n2388 2.2505
R4674 VSS.n6532 VSS.n6531 2.2505
R4675 VSS.n6530 VSS.n2389 2.2505
R4676 VSS.n6529 VSS.n6528 2.2505
R4677 VSS.n6527 VSS.n2390 2.2505
R4678 VSS.n6526 VSS.n6525 2.2505
R4679 VSS.n6524 VSS.n2391 2.2505
R4680 VSS.n6523 VSS.n6522 2.2505
R4681 VSS.n6521 VSS.n2392 2.2505
R4682 VSS.n6520 VSS.n6519 2.2505
R4683 VSS.n6518 VSS.n2393 2.2505
R4684 VSS.n6517 VSS.n6516 2.2505
R4685 VSS.n6515 VSS.n2394 2.2505
R4686 VSS.n6514 VSS.n6513 2.2505
R4687 VSS.n6512 VSS.n2395 2.2505
R4688 VSS.n6511 VSS.n6510 2.2505
R4689 VSS.n6509 VSS.n2396 2.2505
R4690 VSS.n6508 VSS.n6507 2.2505
R4691 VSS.n6506 VSS.n2397 2.2505
R4692 VSS.n6505 VSS.n6504 2.2505
R4693 VSS.n6503 VSS.n2398 2.2505
R4694 VSS.n6502 VSS.n6501 2.2505
R4695 VSS.n6500 VSS.n2399 2.2505
R4696 VSS.n6499 VSS.n6498 2.2505
R4697 VSS.n6497 VSS.n2400 2.2505
R4698 VSS.n6496 VSS.n6495 2.2505
R4699 VSS.n6494 VSS.n2401 2.2505
R4700 VSS.n6493 VSS.n6492 2.2505
R4701 VSS.n6491 VSS.n2402 2.2505
R4702 VSS.n6490 VSS.n6489 2.2505
R4703 VSS.n6488 VSS.n2403 2.2505
R4704 VSS.n6487 VSS.n6486 2.2505
R4705 VSS.n6485 VSS.n2404 2.2505
R4706 VSS.n6484 VSS.n6483 2.2505
R4707 VSS.n6482 VSS.n2405 2.2505
R4708 VSS.n6481 VSS.n6480 2.2505
R4709 VSS.n6479 VSS.n2406 2.2505
R4710 VSS.n6478 VSS.n6477 2.2505
R4711 VSS.n6476 VSS.n2407 2.2505
R4712 VSS.n6475 VSS.n6474 2.2505
R4713 VSS.n6473 VSS.n2408 2.2505
R4714 VSS.n6472 VSS.n6471 2.2505
R4715 VSS.n6470 VSS.n2409 2.2505
R4716 VSS.n6469 VSS.n6468 2.2505
R4717 VSS.n6467 VSS.n2410 2.2505
R4718 VSS.n6466 VSS.n6465 2.2505
R4719 VSS.n6464 VSS.n2411 2.2505
R4720 VSS.n6463 VSS.n6462 2.2505
R4721 VSS.n6461 VSS.n2412 2.2505
R4722 VSS.n6460 VSS.n6459 2.2505
R4723 VSS.n6458 VSS.n2413 2.2505
R4724 VSS.n6457 VSS.n6456 2.2505
R4725 VSS.n6455 VSS.n2414 2.2505
R4726 VSS.n6454 VSS.n6453 2.2505
R4727 VSS.n6452 VSS.n2415 2.2505
R4728 VSS.n6451 VSS.n6450 2.2505
R4729 VSS.n6449 VSS.n2416 2.2505
R4730 VSS.n6448 VSS.n6447 2.2505
R4731 VSS.n6446 VSS.n2417 2.2505
R4732 VSS.n6445 VSS.n6444 2.2505
R4733 VSS.n6443 VSS.n2418 2.2505
R4734 VSS.n6442 VSS.n6441 2.2505
R4735 VSS.n6440 VSS.n2419 2.2505
R4736 VSS.n6439 VSS.n6438 2.2505
R4737 VSS.n6437 VSS.n2420 2.2505
R4738 VSS.n6436 VSS.n6435 2.2505
R4739 VSS.n6434 VSS.n2421 2.2505
R4740 VSS.n6433 VSS.n6432 2.2505
R4741 VSS.n6431 VSS.n2422 2.2505
R4742 VSS.n6430 VSS.n6429 2.2505
R4743 VSS.n6428 VSS.n2423 2.2505
R4744 VSS.n6427 VSS.n6426 2.2505
R4745 VSS.n6425 VSS.n2424 2.2505
R4746 VSS.n6424 VSS.n6423 2.2505
R4747 VSS.n6422 VSS.n2425 2.2505
R4748 VSS.n6421 VSS.n6420 2.2505
R4749 VSS.n6419 VSS.n2426 2.2505
R4750 VSS.n6418 VSS.n6417 2.2505
R4751 VSS.n6416 VSS.n2427 2.2505
R4752 VSS.n6415 VSS.n6414 2.2505
R4753 VSS.n6413 VSS.n2428 2.2505
R4754 VSS.n6412 VSS.n6411 2.2505
R4755 VSS.n6410 VSS.n2429 2.2505
R4756 VSS.n6409 VSS.n6408 2.2505
R4757 VSS.n6407 VSS.n2430 2.2505
R4758 VSS.n6406 VSS.n6405 2.2505
R4759 VSS.n6404 VSS.n2431 2.2505
R4760 VSS.n6403 VSS.n6402 2.2505
R4761 VSS.n6401 VSS.n2432 2.2505
R4762 VSS.n6400 VSS.n6399 2.2505
R4763 VSS.n6398 VSS.n2433 2.2505
R4764 VSS.n6397 VSS.n6396 2.2505
R4765 VSS.n6395 VSS.n2434 2.2505
R4766 VSS.n6394 VSS.n6393 2.2505
R4767 VSS.n6392 VSS.n2435 2.2505
R4768 VSS.n6391 VSS.n6390 2.2505
R4769 VSS.n6389 VSS.n2436 2.2505
R4770 VSS.n6388 VSS.n6387 2.2505
R4771 VSS.n6386 VSS.n2437 2.2505
R4772 VSS.n6385 VSS.n6384 2.2505
R4773 VSS.n6383 VSS.n2438 2.2505
R4774 VSS.n6382 VSS.n6381 2.2505
R4775 VSS.n6380 VSS.n2439 2.2505
R4776 VSS.n6379 VSS.n6378 2.2505
R4777 VSS.n6377 VSS.n2440 2.2505
R4778 VSS.n6376 VSS.n6375 2.2505
R4779 VSS.n6374 VSS.n2441 2.2505
R4780 VSS.n6373 VSS.n6372 2.2505
R4781 VSS.n6371 VSS.n2442 2.2505
R4782 VSS.n6370 VSS.n6369 2.2505
R4783 VSS.n6368 VSS.n2443 2.2505
R4784 VSS.n6367 VSS.n6366 2.2505
R4785 VSS.n6365 VSS.n2444 2.2505
R4786 VSS.n6364 VSS.n6363 2.2505
R4787 VSS.n6362 VSS.n2445 2.2505
R4788 VSS.n6361 VSS.n6360 2.2505
R4789 VSS.n6359 VSS.n2446 2.2505
R4790 VSS.n6358 VSS.n6357 2.2505
R4791 VSS.n6356 VSS.n2447 2.2505
R4792 VSS.n6355 VSS.n6354 2.2505
R4793 VSS.n6353 VSS.n2448 2.2505
R4794 VSS.n6352 VSS.n6351 2.2505
R4795 VSS.n6350 VSS.n2449 2.2505
R4796 VSS.n6349 VSS.n6348 2.2505
R4797 VSS.n6347 VSS.n2450 2.2505
R4798 VSS.n6346 VSS.n6345 2.2505
R4799 VSS.n6344 VSS.n2451 2.2505
R4800 VSS.n6343 VSS.n6342 2.2505
R4801 VSS.n6341 VSS.n2452 2.2505
R4802 VSS.n6340 VSS.n6339 2.2505
R4803 VSS.n6338 VSS.n2453 2.2505
R4804 VSS.n6337 VSS.n6336 2.2505
R4805 VSS.n6335 VSS.n2454 2.2505
R4806 VSS.n6334 VSS.n6333 2.2505
R4807 VSS.n6332 VSS.n2455 2.2505
R4808 VSS.n6331 VSS.n6330 2.2505
R4809 VSS.n6329 VSS.n2456 2.2505
R4810 VSS.n6328 VSS.n6327 2.2505
R4811 VSS.n6326 VSS.n2457 2.2505
R4812 VSS.n6325 VSS.n6324 2.2505
R4813 VSS.n6323 VSS.n2458 2.2505
R4814 VSS.n6322 VSS.n6321 2.2505
R4815 VSS.n6320 VSS.n2459 2.2505
R4816 VSS.n6319 VSS.n6318 2.2505
R4817 VSS.n6317 VSS.n2460 2.2505
R4818 VSS.n6316 VSS.n6315 2.2505
R4819 VSS.n6314 VSS.n2461 2.2505
R4820 VSS.n6313 VSS.n6312 2.2505
R4821 VSS.n6311 VSS.n2462 2.2505
R4822 VSS.n6310 VSS.n6309 2.2505
R4823 VSS.n6308 VSS.n2463 2.2505
R4824 VSS.n6307 VSS.n6306 2.2505
R4825 VSS.n6305 VSS.n2464 2.2505
R4826 VSS.n6304 VSS.n6303 2.2505
R4827 VSS.n6302 VSS.n2465 2.2505
R4828 VSS.n6301 VSS.n6300 2.2505
R4829 VSS.n6299 VSS.n2466 2.2505
R4830 VSS.n6298 VSS.n6297 2.2505
R4831 VSS.n6296 VSS.n2467 2.2505
R4832 VSS.n6295 VSS.n6294 2.2505
R4833 VSS.n6293 VSS.n2468 2.2505
R4834 VSS.n6292 VSS.n6291 2.2505
R4835 VSS.n6290 VSS.n2469 2.2505
R4836 VSS.n6289 VSS.n6288 2.2505
R4837 VSS.n6287 VSS.n2470 2.2505
R4838 VSS.n6286 VSS.n6285 2.2505
R4839 VSS.n6284 VSS.n2471 2.2505
R4840 VSS.n6283 VSS.n6282 2.2505
R4841 VSS.n6281 VSS.n2472 2.2505
R4842 VSS.n6280 VSS.n6279 2.2505
R4843 VSS.n6278 VSS.n2473 2.2505
R4844 VSS.n6277 VSS.n6276 2.2505
R4845 VSS.n6275 VSS.n2474 2.2505
R4846 VSS.n6274 VSS.n6273 2.2505
R4847 VSS.n6272 VSS.n2475 2.2505
R4848 VSS.n6271 VSS.n6270 2.2505
R4849 VSS.n6269 VSS.n2476 2.2505
R4850 VSS.n6268 VSS.n6267 2.2505
R4851 VSS.n6266 VSS.n2477 2.2505
R4852 VSS.n6265 VSS.n6264 2.2505
R4853 VSS.n6263 VSS.n2478 2.2505
R4854 VSS.n6262 VSS.n6261 2.2505
R4855 VSS.n6260 VSS.n2479 2.2505
R4856 VSS.n6259 VSS.n6258 2.2505
R4857 VSS.n6257 VSS.n2480 2.2505
R4858 VSS.n6256 VSS.n6255 2.2505
R4859 VSS.n6254 VSS.n2481 2.2505
R4860 VSS.n6253 VSS.n6252 2.2505
R4861 VSS.n6251 VSS.n2482 2.2505
R4862 VSS.n6250 VSS.n6249 2.2505
R4863 VSS.n6248 VSS.n2483 2.2505
R4864 VSS.n6247 VSS.n6246 2.2505
R4865 VSS.n6245 VSS.n2484 2.2505
R4866 VSS.n6244 VSS.n6243 2.2505
R4867 VSS.n6242 VSS.n2485 2.2505
R4868 VSS.n6241 VSS.n6240 2.2505
R4869 VSS.n6239 VSS.n2486 2.2505
R4870 VSS.n6238 VSS.n6237 2.2505
R4871 VSS.n6236 VSS.n2487 2.2505
R4872 VSS.n6235 VSS.n6234 2.2505
R4873 VSS.n6233 VSS.n2488 2.2505
R4874 VSS.n6232 VSS.n6231 2.2505
R4875 VSS.n6230 VSS.n2489 2.2505
R4876 VSS.n6229 VSS.n6228 2.2505
R4877 VSS.n6227 VSS.n2490 2.2505
R4878 VSS.n6226 VSS.n6225 2.2505
R4879 VSS.n6224 VSS.n2491 2.2505
R4880 VSS.n6223 VSS.n6222 2.2505
R4881 VSS.n6221 VSS.n2492 2.2505
R4882 VSS.n6220 VSS.n6219 2.2505
R4883 VSS.n6218 VSS.n2493 2.2505
R4884 VSS.n6217 VSS.n6216 2.2505
R4885 VSS.n6215 VSS.n2494 2.2505
R4886 VSS.n6214 VSS.n6213 2.2505
R4887 VSS.n6212 VSS.n2495 2.2505
R4888 VSS.n6211 VSS.n6210 2.2505
R4889 VSS.n6209 VSS.n2496 2.2505
R4890 VSS.n6208 VSS.n6207 2.2505
R4891 VSS.n6206 VSS.n2497 2.2505
R4892 VSS.n6205 VSS.n6204 2.2505
R4893 VSS.n6203 VSS.n2498 2.2505
R4894 VSS.n6202 VSS.n6201 2.2505
R4895 VSS.n6200 VSS.n2499 2.2505
R4896 VSS.n6199 VSS.n6198 2.2505
R4897 VSS.n6197 VSS.n2500 2.2505
R4898 VSS.n6196 VSS.n6195 2.2505
R4899 VSS.n6194 VSS.n2501 2.2505
R4900 VSS.n6193 VSS.n6192 2.2505
R4901 VSS.n6191 VSS.n2502 2.2505
R4902 VSS.n6190 VSS.n6189 2.2505
R4903 VSS.n6188 VSS.n2503 2.2505
R4904 VSS.n6187 VSS.n6186 2.2505
R4905 VSS.n6185 VSS.n2504 2.2505
R4906 VSS.n6184 VSS.n6183 2.2505
R4907 VSS.n6182 VSS.n2505 2.2505
R4908 VSS.n6181 VSS.n6180 2.2505
R4909 VSS.n6179 VSS.n2506 2.2505
R4910 VSS.n6178 VSS.n6177 2.2505
R4911 VSS.n6176 VSS.n2507 2.2505
R4912 VSS.n6175 VSS.n6174 2.2505
R4913 VSS.n6173 VSS.n2508 2.2505
R4914 VSS.n6172 VSS.n6171 2.2505
R4915 VSS.n6170 VSS.n2509 2.2505
R4916 VSS.n6169 VSS.n6168 2.2505
R4917 VSS.n6167 VSS.n2510 2.2505
R4918 VSS.n6166 VSS.n6165 2.2505
R4919 VSS.n6164 VSS.n2511 2.2505
R4920 VSS.n6163 VSS.n6162 2.2505
R4921 VSS.n6161 VSS.n2512 2.2505
R4922 VSS.n6160 VSS.n6159 2.2505
R4923 VSS.n6158 VSS.n2513 2.2505
R4924 VSS.n6157 VSS.n6156 2.2505
R4925 VSS.n6155 VSS.n2514 2.2505
R4926 VSS.n6154 VSS.n6153 2.2505
R4927 VSS.n6152 VSS.n2515 2.2505
R4928 VSS.n6151 VSS.n6150 2.2505
R4929 VSS.n6149 VSS.n2516 2.2505
R4930 VSS.n6148 VSS.n6147 2.2505
R4931 VSS.n6146 VSS.n2517 2.2505
R4932 VSS.n6145 VSS.n6144 2.2505
R4933 VSS.n6143 VSS.n2518 2.2505
R4934 VSS.n6142 VSS.n6141 2.2505
R4935 VSS.n6140 VSS.n2519 2.2505
R4936 VSS.n6139 VSS.n6138 2.2505
R4937 VSS.n6137 VSS.n2520 2.2505
R4938 VSS.n6136 VSS.n6135 2.2505
R4939 VSS.n6134 VSS.n2521 2.2505
R4940 VSS.n6133 VSS.n6132 2.2505
R4941 VSS.n6131 VSS.n2522 2.2505
R4942 VSS.n6130 VSS.n6129 2.2505
R4943 VSS.n6128 VSS.n2523 2.2505
R4944 VSS.n6127 VSS.n6126 2.2505
R4945 VSS.n6125 VSS.n2524 2.2505
R4946 VSS.n6124 VSS.n6123 2.2505
R4947 VSS.n6122 VSS.n2525 2.2505
R4948 VSS.n6121 VSS.n6120 2.2505
R4949 VSS.n6119 VSS.n2526 2.2505
R4950 VSS.n6118 VSS.n6117 2.2505
R4951 VSS.n6116 VSS.n2527 2.2505
R4952 VSS.n6115 VSS.n6114 2.2505
R4953 VSS.n6113 VSS.n2528 2.2505
R4954 VSS.n6112 VSS.n6111 2.2505
R4955 VSS.n6110 VSS.n2529 2.2505
R4956 VSS.n6109 VSS.n6108 2.2505
R4957 VSS.n6107 VSS.n2530 2.2505
R4958 VSS.n6106 VSS.n6105 2.2505
R4959 VSS.n6104 VSS.n2531 2.2505
R4960 VSS.n6103 VSS.n6102 2.2505
R4961 VSS.n6101 VSS.n2532 2.2505
R4962 VSS.n6100 VSS.n6099 2.2505
R4963 VSS.n6098 VSS.n2533 2.2505
R4964 VSS.n6097 VSS.n6096 2.2505
R4965 VSS.n6095 VSS.n2534 2.2505
R4966 VSS.n6094 VSS.n6093 2.2505
R4967 VSS.n6092 VSS.n2535 2.2505
R4968 VSS.n6091 VSS.n6090 2.2505
R4969 VSS.n6089 VSS.n2536 2.2505
R4970 VSS.n6088 VSS.n6087 2.2505
R4971 VSS.n6086 VSS.n2537 2.2505
R4972 VSS.n6085 VSS.n6084 2.2505
R4973 VSS.n6083 VSS.n2538 2.2505
R4974 VSS.n6082 VSS.n6081 2.2505
R4975 VSS.n6080 VSS.n2539 2.2505
R4976 VSS.n6079 VSS.n6078 2.2505
R4977 VSS.n6077 VSS.n2540 2.2505
R4978 VSS.n6076 VSS.n6075 2.2505
R4979 VSS.n6074 VSS.n2541 2.2505
R4980 VSS.n6073 VSS.n6072 2.2505
R4981 VSS.n6071 VSS.n2542 2.2505
R4982 VSS.n6070 VSS.n6069 2.2505
R4983 VSS.n6068 VSS.n2543 2.2505
R4984 VSS.n6067 VSS.n6066 2.2505
R4985 VSS.n6065 VSS.n2544 2.2505
R4986 VSS.n6064 VSS.n6063 2.2505
R4987 VSS.n6062 VSS.n2545 2.2505
R4988 VSS.n6061 VSS.n6060 2.2505
R4989 VSS.n6059 VSS.n2546 2.2505
R4990 VSS.n6058 VSS.n6057 2.2505
R4991 VSS.n6056 VSS.n2547 2.2505
R4992 VSS.n6055 VSS.n6054 2.2505
R4993 VSS.n6053 VSS.n2548 2.2505
R4994 VSS.n6052 VSS.n6051 2.2505
R4995 VSS.n6050 VSS.n2549 2.2505
R4996 VSS.n6049 VSS.n6048 2.2505
R4997 VSS.n6047 VSS.n2550 2.2505
R4998 VSS.n6046 VSS.n6045 2.2505
R4999 VSS.n6044 VSS.n2551 2.2505
R5000 VSS.n6043 VSS.n6042 2.2505
R5001 VSS.n6041 VSS.n2552 2.2505
R5002 VSS.n6040 VSS.n6039 2.2505
R5003 VSS.n6038 VSS.n2553 2.2505
R5004 VSS.n6037 VSS.n6036 2.2505
R5005 VSS.n6035 VSS.n2554 2.2505
R5006 VSS.n6034 VSS.n6033 2.2505
R5007 VSS.n6032 VSS.n2555 2.2505
R5008 VSS.n6031 VSS.n6030 2.2505
R5009 VSS.n6029 VSS.n2556 2.2505
R5010 VSS.n6028 VSS.n6027 2.2505
R5011 VSS.n6026 VSS.n2557 2.2505
R5012 VSS.n6025 VSS.n6024 2.2505
R5013 VSS.n6023 VSS.n2558 2.2505
R5014 VSS.n6022 VSS.n6021 2.2505
R5015 VSS.n6020 VSS.n2559 2.2505
R5016 VSS.n6019 VSS.n6018 2.2505
R5017 VSS.n6017 VSS.n2560 2.2505
R5018 VSS.n6016 VSS.n6015 2.2505
R5019 VSS.n6014 VSS.n2561 2.2505
R5020 VSS.n6013 VSS.n6012 2.2505
R5021 VSS.n6011 VSS.n2562 2.2505
R5022 VSS.n6010 VSS.n6009 2.2505
R5023 VSS.n6008 VSS.n2563 2.2505
R5024 VSS.n6007 VSS.n6006 2.2505
R5025 VSS.n6005 VSS.n2564 2.2505
R5026 VSS.n6004 VSS.n6003 2.2505
R5027 VSS.n6002 VSS.n2565 2.2505
R5028 VSS.n6001 VSS.n6000 2.2505
R5029 VSS.n5999 VSS.n2566 2.2505
R5030 VSS.n5998 VSS.n5997 2.2505
R5031 VSS.n5996 VSS.n2567 2.2505
R5032 VSS.n5995 VSS.n5994 2.2505
R5033 VSS.n5993 VSS.n2568 2.2505
R5034 VSS.n5992 VSS.n5991 2.2505
R5035 VSS.n5990 VSS.n2569 2.2505
R5036 VSS.n5989 VSS.n5988 2.2505
R5037 VSS.n5987 VSS.n2570 2.2505
R5038 VSS.n5986 VSS.n5985 2.2505
R5039 VSS.n5984 VSS.n2571 2.2505
R5040 VSS.n5983 VSS.n5982 2.2505
R5041 VSS.n5981 VSS.n2572 2.2505
R5042 VSS.n5980 VSS.n5979 2.2505
R5043 VSS.n5978 VSS.n2573 2.2505
R5044 VSS.n5977 VSS.n5976 2.2505
R5045 VSS.n5975 VSS.n2574 2.2505
R5046 VSS.n5974 VSS.n5973 2.2505
R5047 VSS.n5972 VSS.n2575 2.2505
R5048 VSS.n5971 VSS.n5970 2.2505
R5049 VSS.n5969 VSS.n2576 2.2505
R5050 VSS.n5968 VSS.n5967 2.2505
R5051 VSS.n5966 VSS.n2577 2.2505
R5052 VSS.n5965 VSS.n5964 2.2505
R5053 VSS.n5963 VSS.n2578 2.2505
R5054 VSS.n5962 VSS.n5961 2.2505
R5055 VSS.n5960 VSS.n2579 2.2505
R5056 VSS.n5959 VSS.n5958 2.2505
R5057 VSS.n5957 VSS.n2580 2.2505
R5058 VSS.n5956 VSS.n5955 2.2505
R5059 VSS.n5954 VSS.n2581 2.2505
R5060 VSS.n5953 VSS.n5952 2.2505
R5061 VSS.n5951 VSS.n2582 2.2505
R5062 VSS.n5950 VSS.n5949 2.2505
R5063 VSS.n5948 VSS.n2583 2.2505
R5064 VSS.n5947 VSS.n5946 2.2505
R5065 VSS.n5945 VSS.n2584 2.2505
R5066 VSS.n5944 VSS.n5943 2.2505
R5067 VSS.n5942 VSS.n2585 2.2505
R5068 VSS.n5941 VSS.n5940 2.2505
R5069 VSS.n5939 VSS.n2586 2.2505
R5070 VSS.n5938 VSS.n5937 2.2505
R5071 VSS.n5936 VSS.n2587 2.2505
R5072 VSS.n5935 VSS.n5934 2.2505
R5073 VSS.n5933 VSS.n2588 2.2505
R5074 VSS.n5932 VSS.n5931 2.2505
R5075 VSS.n5930 VSS.n2589 2.2505
R5076 VSS.n5929 VSS.n5928 2.2505
R5077 VSS.n5927 VSS.n2590 2.2505
R5078 VSS.n5926 VSS.n5925 2.2505
R5079 VSS.n5924 VSS.n2591 2.2505
R5080 VSS.n5923 VSS.n5922 2.2505
R5081 VSS.n5921 VSS.n2592 2.2505
R5082 VSS.n5920 VSS.n5919 2.2505
R5083 VSS.n5918 VSS.n2593 2.2505
R5084 VSS.n5917 VSS.n5916 2.2505
R5085 VSS.n5915 VSS.n2594 2.2505
R5086 VSS.n5914 VSS.n5913 2.2505
R5087 VSS.n5912 VSS.n2595 2.2505
R5088 VSS.n5911 VSS.n5910 2.2505
R5089 VSS.n5909 VSS.n2596 2.2505
R5090 VSS.n5908 VSS.n5907 2.2505
R5091 VSS.n5906 VSS.n2597 2.2505
R5092 VSS.n5905 VSS.n5904 2.2505
R5093 VSS.n5903 VSS.n2598 2.2505
R5094 VSS.n5902 VSS.n5901 2.2505
R5095 VSS.n5900 VSS.n2599 2.2505
R5096 VSS.n5899 VSS.n5898 2.2505
R5097 VSS.n5897 VSS.n2600 2.2505
R5098 VSS.n5896 VSS.n5895 2.2505
R5099 VSS.n5894 VSS.n2601 2.2505
R5100 VSS.n5893 VSS.n5892 2.2505
R5101 VSS.n5891 VSS.n2602 2.2505
R5102 VSS.n5890 VSS.n5889 2.2505
R5103 VSS.n5888 VSS.n2603 2.2505
R5104 VSS.n5887 VSS.n5886 2.2505
R5105 VSS.n5885 VSS.n2604 2.2505
R5106 VSS.n5884 VSS.n5883 2.2505
R5107 VSS.n5882 VSS.n2605 2.2505
R5108 VSS.n5881 VSS.n5880 2.2505
R5109 VSS.n5879 VSS.n2606 2.2505
R5110 VSS.n5878 VSS.n5877 2.2505
R5111 VSS.n5876 VSS.n2607 2.2505
R5112 VSS.n5875 VSS.n5874 2.2505
R5113 VSS.n5873 VSS.n2608 2.2505
R5114 VSS.n5872 VSS.n5871 2.2505
R5115 VSS.n5870 VSS.n2609 2.2505
R5116 VSS.n5869 VSS.n5868 2.2505
R5117 VSS.n5867 VSS.n2610 2.2505
R5118 VSS.n5866 VSS.n5865 2.2505
R5119 VSS.n5864 VSS.n2611 2.2505
R5120 VSS.n5863 VSS.n5862 2.2505
R5121 VSS.n5861 VSS.n2612 2.2505
R5122 VSS.n5860 VSS.n5859 2.2505
R5123 VSS.n5858 VSS.n2613 2.2505
R5124 VSS.n5857 VSS.n5856 2.2505
R5125 VSS.n5855 VSS.n2614 2.2505
R5126 VSS.n5854 VSS.n5853 2.2505
R5127 VSS.n5852 VSS.n2615 2.2505
R5128 VSS.n5851 VSS.n5850 2.2505
R5129 VSS.n5849 VSS.n2616 2.2505
R5130 VSS.n5848 VSS.n5847 2.2505
R5131 VSS.n5846 VSS.n2617 2.2505
R5132 VSS.n5845 VSS.n5844 2.2505
R5133 VSS.n5843 VSS.n2618 2.2505
R5134 VSS.n5842 VSS.n5841 2.2505
R5135 VSS.n5840 VSS.n2619 2.2505
R5136 VSS.n5839 VSS.n5838 2.2505
R5137 VSS.n5837 VSS.n2620 2.2505
R5138 VSS.n5836 VSS.n5835 2.2505
R5139 VSS.n5834 VSS.n2621 2.2505
R5140 VSS.n5833 VSS.n5832 2.2505
R5141 VSS.n5831 VSS.n2622 2.2505
R5142 VSS.n5830 VSS.n5829 2.2505
R5143 VSS.n5828 VSS.n2623 2.2505
R5144 VSS.n5827 VSS.n5826 2.2505
R5145 VSS.n5825 VSS.n2624 2.2505
R5146 VSS.n5824 VSS.n5823 2.2505
R5147 VSS.n5822 VSS.n2625 2.2505
R5148 VSS.n5821 VSS.n5820 2.2505
R5149 VSS.n5819 VSS.n2626 2.2505
R5150 VSS.n5818 VSS.n5817 2.2505
R5151 VSS.n5816 VSS.n2627 2.2505
R5152 VSS.n5815 VSS.n5814 2.2505
R5153 VSS.n5813 VSS.n2628 2.2505
R5154 VSS.n5812 VSS.n5811 2.2505
R5155 VSS.n5810 VSS.n2629 2.2505
R5156 VSS.n5809 VSS.n5808 2.2505
R5157 VSS.n5807 VSS.n2630 2.2505
R5158 VSS.n5806 VSS.n5805 2.2505
R5159 VSS.n5804 VSS.n2631 2.2505
R5160 VSS.n5803 VSS.n5802 2.2505
R5161 VSS.n5801 VSS.n2632 2.2505
R5162 VSS.n5800 VSS.n5799 2.2505
R5163 VSS.n5798 VSS.n2633 2.2505
R5164 VSS.n5797 VSS.n5796 2.2505
R5165 VSS.n5795 VSS.n2634 2.2505
R5166 VSS.n5794 VSS.n5793 2.2505
R5167 VSS.n5792 VSS.n2635 2.2505
R5168 VSS.n5791 VSS.n5790 2.2505
R5169 VSS.n5789 VSS.n2636 2.2505
R5170 VSS.n5788 VSS.n5787 2.2505
R5171 VSS.n5786 VSS.n2637 2.2505
R5172 VSS.n5785 VSS.n5784 2.2505
R5173 VSS.n5783 VSS.n2638 2.2505
R5174 VSS.n5782 VSS.n5781 2.2505
R5175 VSS.n5780 VSS.n2639 2.2505
R5176 VSS.n5779 VSS.n5778 2.2505
R5177 VSS.n5777 VSS.n2640 2.2505
R5178 VSS.n5776 VSS.n5775 2.2505
R5179 VSS.n5774 VSS.n2641 2.2505
R5180 VSS.n5773 VSS.n5772 2.2505
R5181 VSS.n5771 VSS.n2642 2.2505
R5182 VSS.n5770 VSS.n5769 2.2505
R5183 VSS.n5768 VSS.n2643 2.2505
R5184 VSS.n5767 VSS.n5766 2.2505
R5185 VSS.n5765 VSS.n2644 2.2505
R5186 VSS.n5764 VSS.n5763 2.2505
R5187 VSS.n5762 VSS.n2645 2.2505
R5188 VSS.n5761 VSS.n5760 2.2505
R5189 VSS.n5759 VSS.n2646 2.2505
R5190 VSS.n5758 VSS.n5757 2.2505
R5191 VSS.n5756 VSS.n2647 2.2505
R5192 VSS.n5755 VSS.n5754 2.2505
R5193 VSS.n5753 VSS.n2648 2.2505
R5194 VSS.n5752 VSS.n5751 2.2505
R5195 VSS.n5750 VSS.n2649 2.2505
R5196 VSS.n5749 VSS.n5748 2.2505
R5197 VSS.n5747 VSS.n2650 2.2505
R5198 VSS.n5746 VSS.n5745 2.2505
R5199 VSS.n5744 VSS.n2651 2.2505
R5200 VSS.n5743 VSS.n5742 2.2505
R5201 VSS.n5741 VSS.n2652 2.2505
R5202 VSS.n5740 VSS.n5739 2.2505
R5203 VSS.n5738 VSS.n2653 2.2505
R5204 VSS.n5737 VSS.n5736 2.2505
R5205 VSS.n5735 VSS.n2654 2.2505
R5206 VSS.n5734 VSS.n5733 2.2505
R5207 VSS.n5732 VSS.n2655 2.2505
R5208 VSS.n5731 VSS.n5730 2.2505
R5209 VSS.n5729 VSS.n2656 2.2505
R5210 VSS.n5728 VSS.n5727 2.2505
R5211 VSS.n5726 VSS.n2657 2.2505
R5212 VSS.n5725 VSS.n5724 2.2505
R5213 VSS.n5723 VSS.n2658 2.2505
R5214 VSS.n5722 VSS.n5721 2.2505
R5215 VSS.n5720 VSS.n2659 2.2505
R5216 VSS.n5719 VSS.n5718 2.2505
R5217 VSS.n5717 VSS.n2660 2.2505
R5218 VSS.n5716 VSS.n5715 2.2505
R5219 VSS.n5714 VSS.n2661 2.2505
R5220 VSS.n5713 VSS.n5712 2.2505
R5221 VSS.n5711 VSS.n2662 2.2505
R5222 VSS.n5710 VSS.n5709 2.2505
R5223 VSS.n5708 VSS.n2663 2.2505
R5224 VSS.n5707 VSS.n5706 2.2505
R5225 VSS.n5705 VSS.n2664 2.2505
R5226 VSS.n5704 VSS.n5703 2.2505
R5227 VSS.n5702 VSS.n2665 2.2505
R5228 VSS.n5701 VSS.n5700 2.2505
R5229 VSS.n5699 VSS.n2666 2.2505
R5230 VSS.n5698 VSS.n5697 2.2505
R5231 VSS.n5696 VSS.n2667 2.2505
R5232 VSS.n5695 VSS.n5694 2.2505
R5233 VSS.n5693 VSS.n2668 2.2505
R5234 VSS.n5692 VSS.n5691 2.2505
R5235 VSS.n5690 VSS.n2669 2.2505
R5236 VSS.n5689 VSS.n5688 2.2505
R5237 VSS.n5687 VSS.n2670 2.2505
R5238 VSS.n5686 VSS.n5685 2.2505
R5239 VSS.n5684 VSS.n2671 2.2505
R5240 VSS.n5683 VSS.n5682 2.2505
R5241 VSS.n5681 VSS.n2672 2.2505
R5242 VSS.n5680 VSS.n5679 2.2505
R5243 VSS.n5678 VSS.n2673 2.2505
R5244 VSS.n5677 VSS.n5676 2.2505
R5245 VSS.n5675 VSS.n2674 2.2505
R5246 VSS.n5674 VSS.n5673 2.2505
R5247 VSS.n5672 VSS.n2675 2.2505
R5248 VSS.n5671 VSS.n5670 2.2505
R5249 VSS.n5669 VSS.n2676 2.2505
R5250 VSS.n5668 VSS.n5667 2.2505
R5251 VSS.n5666 VSS.n2677 2.2505
R5252 VSS.n5665 VSS.n5664 2.2505
R5253 VSS.n5663 VSS.n2678 2.2505
R5254 VSS.n5662 VSS.n5661 2.2505
R5255 VSS.n5660 VSS.n2679 2.2505
R5256 VSS.n5659 VSS.n5658 2.2505
R5257 VSS.n5657 VSS.n2680 2.2505
R5258 VSS.n5656 VSS.n5655 2.2505
R5259 VSS.n5654 VSS.n2681 2.2505
R5260 VSS.n5653 VSS.n5652 2.2505
R5261 VSS.n5651 VSS.n2682 2.2505
R5262 VSS.n5650 VSS.n5649 2.2505
R5263 VSS.n5648 VSS.n2683 2.2505
R5264 VSS.n5647 VSS.n5646 2.2505
R5265 VSS.n5645 VSS.n2684 2.2505
R5266 VSS.n5644 VSS.n5643 2.2505
R5267 VSS.n5642 VSS.n2685 2.2505
R5268 VSS.n5641 VSS.n5640 2.2505
R5269 VSS.n5639 VSS.n2686 2.2505
R5270 VSS.n5638 VSS.n5637 2.2505
R5271 VSS.n5636 VSS.n2687 2.2505
R5272 VSS.n5635 VSS.n5634 2.2505
R5273 VSS.n5633 VSS.n2688 2.2505
R5274 VSS.n5632 VSS.n5631 2.2505
R5275 VSS.n5630 VSS.n2689 2.2505
R5276 VSS.n5629 VSS.n5628 2.2505
R5277 VSS.n5627 VSS.n2690 2.2505
R5278 VSS.n5626 VSS.n5625 2.2505
R5279 VSS.n5624 VSS.n2691 2.2505
R5280 VSS.n5623 VSS.n5622 2.2505
R5281 VSS.n5621 VSS.n2692 2.2505
R5282 VSS.n5620 VSS.n5619 2.2505
R5283 VSS.n5618 VSS.n2693 2.2505
R5284 VSS.n5617 VSS.n5616 2.2505
R5285 VSS.n5615 VSS.n2694 2.2505
R5286 VSS.n5614 VSS.n5613 2.2505
R5287 VSS.n5612 VSS.n2695 2.2505
R5288 VSS.n5611 VSS.n5610 2.2505
R5289 VSS.n5609 VSS.n2696 2.2505
R5290 VSS.n5608 VSS.n5607 2.2505
R5291 VSS.n5606 VSS.n2697 2.2505
R5292 VSS.n5605 VSS.n5604 2.2505
R5293 VSS.n5603 VSS.n2698 2.2505
R5294 VSS.n5602 VSS.n5601 2.2505
R5295 VSS.n5600 VSS.n2699 2.2505
R5296 VSS.n5599 VSS.n5598 2.2505
R5297 VSS.n5597 VSS.n2700 2.2505
R5298 VSS.n5596 VSS.n5595 2.2505
R5299 VSS.n5594 VSS.n2701 2.2505
R5300 VSS.n5593 VSS.n5592 2.2505
R5301 VSS.n5591 VSS.n2702 2.2505
R5302 VSS.n5590 VSS.n5589 2.2505
R5303 VSS.n5588 VSS.n2703 2.2505
R5304 VSS.n5587 VSS.n5586 2.2505
R5305 VSS.n5585 VSS.n2704 2.2505
R5306 VSS.n5584 VSS.n5583 2.2505
R5307 VSS.n5582 VSS.n2705 2.2505
R5308 VSS.n5581 VSS.n5580 2.2505
R5309 VSS.n5579 VSS.n2706 2.2505
R5310 VSS.n5578 VSS.n5577 2.2505
R5311 VSS.n5576 VSS.n2707 2.2505
R5312 VSS.n5575 VSS.n5574 2.2505
R5313 VSS.n5573 VSS.n2708 2.2505
R5314 VSS.n5572 VSS.n5571 2.2505
R5315 VSS.n5570 VSS.n2709 2.2505
R5316 VSS.n5569 VSS.n5568 2.2505
R5317 VSS.n5567 VSS.n2710 2.2505
R5318 VSS.n5566 VSS.n5565 2.2505
R5319 VSS.n5564 VSS.n2711 2.2505
R5320 VSS.n5563 VSS.n5562 2.2505
R5321 VSS.n5561 VSS.n2712 2.2505
R5322 VSS.n5560 VSS.n5559 2.2505
R5323 VSS.n5558 VSS.n2713 2.2505
R5324 VSS.n5557 VSS.n5556 2.2505
R5325 VSS.n5555 VSS.n2714 2.2505
R5326 VSS.n5554 VSS.n5553 2.2505
R5327 VSS.n5552 VSS.n2715 2.2505
R5328 VSS.n5551 VSS.n5550 2.2505
R5329 VSS.n5549 VSS.n2716 2.2505
R5330 VSS.n5548 VSS.n5547 2.2505
R5331 VSS.n5546 VSS.n2717 2.2505
R5332 VSS.n5545 VSS.n5544 2.2505
R5333 VSS.n5543 VSS.n2718 2.2505
R5334 VSS.n5542 VSS.n5541 2.2505
R5335 VSS.n5540 VSS.n2719 2.2505
R5336 VSS.n5539 VSS.n5538 2.2505
R5337 VSS.n5537 VSS.n2720 2.2505
R5338 VSS.n5536 VSS.n5535 2.2505
R5339 VSS.n5534 VSS.n2721 2.2505
R5340 VSS.n5533 VSS.n5532 2.2505
R5341 VSS.n5531 VSS.n2722 2.2505
R5342 VSS.n5530 VSS.n5529 2.2505
R5343 VSS.n5528 VSS.n2723 2.2505
R5344 VSS.n5527 VSS.n5526 2.2505
R5345 VSS.n5525 VSS.n2724 2.2505
R5346 VSS.n5524 VSS.n5523 2.2505
R5347 VSS.n5522 VSS.n2725 2.2505
R5348 VSS.n5521 VSS.n5520 2.2505
R5349 VSS.n5519 VSS.n2726 2.2505
R5350 VSS.n5518 VSS.n5517 2.2505
R5351 VSS.n5516 VSS.n2727 2.2505
R5352 VSS.n5515 VSS.n5514 2.2505
R5353 VSS.n5513 VSS.n2728 2.2505
R5354 VSS.n5512 VSS.n5511 2.2505
R5355 VSS.n5510 VSS.n2729 2.2505
R5356 VSS.n5509 VSS.n5508 2.2505
R5357 VSS.n5507 VSS.n2730 2.2505
R5358 VSS.n5506 VSS.n5505 2.2505
R5359 VSS.n5504 VSS.n2731 2.2505
R5360 VSS.n5503 VSS.n5502 2.2505
R5361 VSS.n5501 VSS.n2732 2.2505
R5362 VSS.n5500 VSS.n5499 2.2505
R5363 VSS.n5498 VSS.n2733 2.2505
R5364 VSS.n5497 VSS.n5496 2.2505
R5365 VSS.n5495 VSS.n2734 2.2505
R5366 VSS.n5494 VSS.n5493 2.2505
R5367 VSS.n5492 VSS.n2735 2.2505
R5368 VSS.n5491 VSS.n5490 2.2505
R5369 VSS.n5489 VSS.n2736 2.2505
R5370 VSS.n5488 VSS.n5487 2.2505
R5371 VSS.n5486 VSS.n2737 2.2505
R5372 VSS.n5485 VSS.n5484 2.2505
R5373 VSS.n5483 VSS.n2738 2.2505
R5374 VSS.n5482 VSS.n5481 2.2505
R5375 VSS.n5480 VSS.n2739 2.2505
R5376 VSS.n5479 VSS.n5478 2.2505
R5377 VSS.n5477 VSS.n2740 2.2505
R5378 VSS.n5476 VSS.n5475 2.2505
R5379 VSS.n5474 VSS.n2741 2.2505
R5380 VSS.n5473 VSS.n5472 2.2505
R5381 VSS.n5471 VSS.n2742 2.2505
R5382 VSS.n5470 VSS.n5469 2.2505
R5383 VSS.n6908 VSS.n2263 2.2505
R5384 VSS.n6910 VSS.n6909 2.2505
R5385 VSS.n6911 VSS.n2262 2.2505
R5386 VSS.n6913 VSS.n6912 2.2505
R5387 VSS.n6914 VSS.n2261 2.2505
R5388 VSS.n6916 VSS.n6915 2.2505
R5389 VSS.n6917 VSS.n2260 2.2505
R5390 VSS.n6919 VSS.n6918 2.2505
R5391 VSS.n6920 VSS.n2259 2.2505
R5392 VSS.n6922 VSS.n6921 2.2505
R5393 VSS.n6923 VSS.n2258 2.2505
R5394 VSS.n6925 VSS.n6924 2.2505
R5395 VSS.n6926 VSS.n2257 2.2505
R5396 VSS.n6928 VSS.n6927 2.2505
R5397 VSS.n6929 VSS.n2256 2.2505
R5398 VSS.n6931 VSS.n6930 2.2505
R5399 VSS.n6932 VSS.n2255 2.2505
R5400 VSS.n6934 VSS.n6933 2.2505
R5401 VSS.n6935 VSS.n2254 2.2505
R5402 VSS.n6937 VSS.n6936 2.2505
R5403 VSS.n6938 VSS.n2253 2.2505
R5404 VSS.n6940 VSS.n6939 2.2505
R5405 VSS.n6941 VSS.n2252 2.2505
R5406 VSS.n6943 VSS.n6942 2.2505
R5407 VSS.n6944 VSS.n2251 2.2505
R5408 VSS.n6946 VSS.n6945 2.2505
R5409 VSS.n6947 VSS.n2250 2.2505
R5410 VSS.n6949 VSS.n6948 2.2505
R5411 VSS.n6950 VSS.n2249 2.2505
R5412 VSS.n6952 VSS.n6951 2.2505
R5413 VSS.n6953 VSS.n2248 2.2505
R5414 VSS.n6955 VSS.n6954 2.2505
R5415 VSS.n6956 VSS.n2247 2.2505
R5416 VSS.n6958 VSS.n6957 2.2505
R5417 VSS.n6959 VSS.n2246 2.2505
R5418 VSS.n6961 VSS.n6960 2.2505
R5419 VSS.n6962 VSS.n2245 2.2505
R5420 VSS.n6964 VSS.n6963 2.2505
R5421 VSS.n6965 VSS.n2244 2.2505
R5422 VSS.n6967 VSS.n6966 2.2505
R5423 VSS.n6968 VSS.n2243 2.2505
R5424 VSS.n6970 VSS.n6969 2.2505
R5425 VSS.n6971 VSS.n2242 2.2505
R5426 VSS.n6973 VSS.n6972 2.2505
R5427 VSS.n6974 VSS.n2241 2.2505
R5428 VSS.n6976 VSS.n6975 2.2505
R5429 VSS.n6977 VSS.n2240 2.2505
R5430 VSS.n6979 VSS.n6978 2.2505
R5431 VSS.n6980 VSS.n2239 2.2505
R5432 VSS.n6982 VSS.n6981 2.2505
R5433 VSS.n6983 VSS.n2238 2.2505
R5434 VSS.n6985 VSS.n6984 2.2505
R5435 VSS.n6986 VSS.n2237 2.2505
R5436 VSS.n6988 VSS.n6987 2.2505
R5437 VSS.n6989 VSS.n2236 2.2505
R5438 VSS.n6991 VSS.n6990 2.2505
R5439 VSS.n6992 VSS.n2235 2.2505
R5440 VSS.n6994 VSS.n6993 2.2505
R5441 VSS.n6995 VSS.n2234 2.2505
R5442 VSS.n6997 VSS.n6996 2.2505
R5443 VSS.n6998 VSS.n2233 2.2505
R5444 VSS.n7000 VSS.n6999 2.2505
R5445 VSS.n7001 VSS.n2232 2.2505
R5446 VSS.n7003 VSS.n7002 2.2505
R5447 VSS.n7004 VSS.n2231 2.2505
R5448 VSS.n7006 VSS.n7005 2.2505
R5449 VSS.n7007 VSS.n2230 2.2505
R5450 VSS.n7009 VSS.n7008 2.2505
R5451 VSS.n7010 VSS.n2229 2.2505
R5452 VSS.n7012 VSS.n7011 2.2505
R5453 VSS.n7013 VSS.n2228 2.2505
R5454 VSS.n7015 VSS.n7014 2.2505
R5455 VSS.n7016 VSS.n2227 2.2505
R5456 VSS.n7018 VSS.n7017 2.2505
R5457 VSS.n7019 VSS.n2226 2.2505
R5458 VSS.n7021 VSS.n7020 2.2505
R5459 VSS.n7022 VSS.n2225 2.2505
R5460 VSS.n7024 VSS.n7023 2.2505
R5461 VSS.n7025 VSS.n2224 2.2505
R5462 VSS.n7027 VSS.n7026 2.2505
R5463 VSS.n7028 VSS.n2223 2.2505
R5464 VSS.n7030 VSS.n7029 2.2505
R5465 VSS.n7031 VSS.n2222 2.2505
R5466 VSS.n7033 VSS.n7032 2.2505
R5467 VSS.n7034 VSS.n2221 2.2505
R5468 VSS.n7036 VSS.n7035 2.2505
R5469 VSS.n7037 VSS.n2220 2.2505
R5470 VSS.n7039 VSS.n7038 2.2505
R5471 VSS.n7040 VSS.n2219 2.2505
R5472 VSS.n7042 VSS.n7041 2.2505
R5473 VSS.n7043 VSS.n2218 2.2505
R5474 VSS.n7045 VSS.n7044 2.2505
R5475 VSS.n7046 VSS.n2217 2.2505
R5476 VSS.n7048 VSS.n7047 2.2505
R5477 VSS.n7049 VSS.n2216 2.2505
R5478 VSS.n7051 VSS.n7050 2.2505
R5479 VSS.n7052 VSS.n2215 2.2505
R5480 VSS.n7054 VSS.n7053 2.2505
R5481 VSS.n7055 VSS.n2214 2.2505
R5482 VSS.n7057 VSS.n7056 2.2505
R5483 VSS.n7058 VSS.n2213 2.2505
R5484 VSS.n7060 VSS.n7059 2.2505
R5485 VSS.n7061 VSS.n2212 2.2505
R5486 VSS.n7063 VSS.n7062 2.2505
R5487 VSS.n7064 VSS.n2211 2.2505
R5488 VSS.n7066 VSS.n7065 2.2505
R5489 VSS.n7067 VSS.n2210 2.2505
R5490 VSS.n7069 VSS.n7068 2.2505
R5491 VSS.n7070 VSS.n2209 2.2505
R5492 VSS.n7072 VSS.n7071 2.2505
R5493 VSS.n7073 VSS.n2208 2.2505
R5494 VSS.n7075 VSS.n7074 2.2505
R5495 VSS.n7076 VSS.n2207 2.2505
R5496 VSS.n7078 VSS.n7077 2.2505
R5497 VSS.n7079 VSS.n2206 2.2505
R5498 VSS.n7081 VSS.n7080 2.2505
R5499 VSS.n7082 VSS.n2205 2.2505
R5500 VSS.n7084 VSS.n7083 2.2505
R5501 VSS.n7085 VSS.n2204 2.2505
R5502 VSS.n7087 VSS.n7086 2.2505
R5503 VSS.n7088 VSS.n2203 2.2505
R5504 VSS.n7090 VSS.n7089 2.2505
R5505 VSS.n7091 VSS.n2202 2.2505
R5506 VSS.n7093 VSS.n7092 2.2505
R5507 VSS.n7094 VSS.n2201 2.2505
R5508 VSS.n7096 VSS.n7095 2.2505
R5509 VSS.n7097 VSS.n2200 2.2505
R5510 VSS.n7099 VSS.n7098 2.2505
R5511 VSS.n7100 VSS.n2199 2.2505
R5512 VSS.n7102 VSS.n7101 2.2505
R5513 VSS.n7103 VSS.n2198 2.2505
R5514 VSS.n7105 VSS.n7104 2.2505
R5515 VSS.n7106 VSS.n2197 2.2505
R5516 VSS.n7108 VSS.n7107 2.2505
R5517 VSS.n7109 VSS.n2196 2.2505
R5518 VSS.n7111 VSS.n7110 2.2505
R5519 VSS.n7112 VSS.n2195 2.2505
R5520 VSS.n7114 VSS.n7113 2.2505
R5521 VSS.n7115 VSS.n2194 2.2505
R5522 VSS.n7117 VSS.n7116 2.2505
R5523 VSS.n7118 VSS.n2193 2.2505
R5524 VSS.n7120 VSS.n7119 2.2505
R5525 VSS.n7121 VSS.n2192 2.2505
R5526 VSS.n7123 VSS.n7122 2.2505
R5527 VSS.n7124 VSS.n2191 2.2505
R5528 VSS.n7126 VSS.n7125 2.2505
R5529 VSS.n7127 VSS.n2190 2.2505
R5530 VSS.n7129 VSS.n7128 2.2505
R5531 VSS.n7130 VSS.n2189 2.2505
R5532 VSS.n7132 VSS.n7131 2.2505
R5533 VSS.n7133 VSS.n2188 2.2505
R5534 VSS.n7135 VSS.n7134 2.2505
R5535 VSS.n7136 VSS.n2187 2.2505
R5536 VSS.n7138 VSS.n7137 2.2505
R5537 VSS.n7139 VSS.n2186 2.2505
R5538 VSS.n7141 VSS.n7140 2.2505
R5539 VSS.n7142 VSS.n2185 2.2505
R5540 VSS.n7144 VSS.n7143 2.2505
R5541 VSS.n7145 VSS.n2184 2.2505
R5542 VSS.n7147 VSS.n7146 2.2505
R5543 VSS.n7148 VSS.n2183 2.2505
R5544 VSS.n7150 VSS.n7149 2.2505
R5545 VSS.n7151 VSS.n2182 2.2505
R5546 VSS.n7153 VSS.n7152 2.2505
R5547 VSS.n7154 VSS.n2181 2.2505
R5548 VSS.n7156 VSS.n7155 2.2505
R5549 VSS.n7157 VSS.n2180 2.2505
R5550 VSS.n7159 VSS.n7158 2.2505
R5551 VSS.n7160 VSS.n2179 2.2505
R5552 VSS.n7162 VSS.n7161 2.2505
R5553 VSS.n7163 VSS.n2178 2.2505
R5554 VSS.n7165 VSS.n7164 2.2505
R5555 VSS.n7166 VSS.n2177 2.2505
R5556 VSS.n7168 VSS.n7167 2.2505
R5557 VSS.n7169 VSS.n2176 2.2505
R5558 VSS.n7171 VSS.n7170 2.2505
R5559 VSS.n7172 VSS.n2175 2.2505
R5560 VSS.n7174 VSS.n7173 2.2505
R5561 VSS.n7175 VSS.n2174 2.2505
R5562 VSS.n7177 VSS.n7176 2.2505
R5563 VSS.n7178 VSS.n2173 2.2505
R5564 VSS.n7180 VSS.n7179 2.2505
R5565 VSS.n7181 VSS.n2172 2.2505
R5566 VSS.n7183 VSS.n7182 2.2505
R5567 VSS.n7184 VSS.n2171 2.2505
R5568 VSS.n7186 VSS.n7185 2.2505
R5569 VSS.n7187 VSS.n2170 2.2505
R5570 VSS.n7189 VSS.n7188 2.2505
R5571 VSS.n7190 VSS.n2169 2.2505
R5572 VSS.n7192 VSS.n7191 2.2505
R5573 VSS.n7193 VSS.n2168 2.2505
R5574 VSS.n7195 VSS.n7194 2.2505
R5575 VSS.n7196 VSS.n2167 2.2505
R5576 VSS.n7198 VSS.n7197 2.2505
R5577 VSS.n7199 VSS.n2166 2.2505
R5578 VSS.n7201 VSS.n7200 2.2505
R5579 VSS.n7202 VSS.n2165 2.2505
R5580 VSS.n7204 VSS.n7203 2.2505
R5581 VSS.n7205 VSS.n2164 2.2505
R5582 VSS.n7207 VSS.n7206 2.2505
R5583 VSS.n7208 VSS.n2163 2.2505
R5584 VSS.n7210 VSS.n7209 2.2505
R5585 VSS.n7211 VSS.n2162 2.2505
R5586 VSS.n7213 VSS.n7212 2.2505
R5587 VSS.n7214 VSS.n2161 2.2505
R5588 VSS.n7216 VSS.n7215 2.2505
R5589 VSS.n7217 VSS.n2160 2.2505
R5590 VSS.n7219 VSS.n7218 2.2505
R5591 VSS.n7220 VSS.n2159 2.2505
R5592 VSS.n7222 VSS.n7221 2.2505
R5593 VSS.n7223 VSS.n2158 2.2505
R5594 VSS.n7225 VSS.n7224 2.2505
R5595 VSS.n7226 VSS.n2157 2.2505
R5596 VSS.n7228 VSS.n7227 2.2505
R5597 VSS.n7229 VSS.n2156 2.2505
R5598 VSS.n7231 VSS.n7230 2.2505
R5599 VSS.n7232 VSS.n2155 2.2505
R5600 VSS.n7234 VSS.n7233 2.2505
R5601 VSS.n7235 VSS.n2154 2.2505
R5602 VSS.n7237 VSS.n7236 2.2505
R5603 VSS.n7238 VSS.n2153 2.2505
R5604 VSS.n7240 VSS.n7239 2.2505
R5605 VSS.n7241 VSS.n2152 2.2505
R5606 VSS.n7243 VSS.n7242 2.2505
R5607 VSS.n7244 VSS.n2151 2.2505
R5608 VSS.n7246 VSS.n7245 2.2505
R5609 VSS.n7247 VSS.n2150 2.2505
R5610 VSS.n7249 VSS.n7248 2.2505
R5611 VSS.n7250 VSS.n2149 2.2505
R5612 VSS.n7252 VSS.n7251 2.2505
R5613 VSS.n7253 VSS.n2148 2.2505
R5614 VSS.n7255 VSS.n7254 2.2505
R5615 VSS.n7256 VSS.n2147 2.2505
R5616 VSS.n7258 VSS.n7257 2.2505
R5617 VSS.n7259 VSS.n2146 2.2505
R5618 VSS.n7261 VSS.n7260 2.2505
R5619 VSS.n7262 VSS.n2145 2.2505
R5620 VSS.n7264 VSS.n7263 2.2505
R5621 VSS.n7265 VSS.n2144 2.2505
R5622 VSS.n7267 VSS.n7266 2.2505
R5623 VSS.n7268 VSS.n2143 2.2505
R5624 VSS.n7270 VSS.n7269 2.2505
R5625 VSS.n7271 VSS.n2142 2.2505
R5626 VSS.n7273 VSS.n7272 2.2505
R5627 VSS.n7274 VSS.n2141 2.2505
R5628 VSS.n7276 VSS.n7275 2.2505
R5629 VSS.n7277 VSS.n2140 2.2505
R5630 VSS.n7279 VSS.n7278 2.2505
R5631 VSS.n7280 VSS.n2139 2.2505
R5632 VSS.n7282 VSS.n7281 2.2505
R5633 VSS.n7283 VSS.n2138 2.2505
R5634 VSS.n7285 VSS.n7284 2.2505
R5635 VSS.n7286 VSS.n2137 2.2505
R5636 VSS.n7288 VSS.n7287 2.2505
R5637 VSS.n7289 VSS.n2136 2.2505
R5638 VSS.n7291 VSS.n7290 2.2505
R5639 VSS.n7292 VSS.n2135 2.2505
R5640 VSS.n7294 VSS.n7293 2.2505
R5641 VSS.n7295 VSS.n2134 2.2505
R5642 VSS.n7297 VSS.n7296 2.2505
R5643 VSS.n7298 VSS.n2133 2.2505
R5644 VSS.n7300 VSS.n7299 2.2505
R5645 VSS.n7301 VSS.n2132 2.2505
R5646 VSS.n7303 VSS.n7302 2.2505
R5647 VSS.n7304 VSS.n2131 2.2505
R5648 VSS.n7306 VSS.n7305 2.2505
R5649 VSS.n7307 VSS.n2130 2.2505
R5650 VSS.n7309 VSS.n7308 2.2505
R5651 VSS.n7310 VSS.n2129 2.2505
R5652 VSS.n7312 VSS.n7311 2.2505
R5653 VSS.n7313 VSS.n2128 2.2505
R5654 VSS.n7315 VSS.n7314 2.2505
R5655 VSS.n7316 VSS.n2127 2.2505
R5656 VSS.n7318 VSS.n7317 2.2505
R5657 VSS.n7319 VSS.n2126 2.2505
R5658 VSS.n7321 VSS.n7320 2.2505
R5659 VSS.n7322 VSS.n2125 2.2505
R5660 VSS.n7324 VSS.n7323 2.2505
R5661 VSS.n7325 VSS.n2124 2.2505
R5662 VSS.n7327 VSS.n7326 2.2505
R5663 VSS.n7328 VSS.n2123 2.2505
R5664 VSS.n7330 VSS.n7329 2.2505
R5665 VSS.n7331 VSS.n2122 2.2505
R5666 VSS.n7333 VSS.n7332 2.2505
R5667 VSS.n7334 VSS.n2121 2.2505
R5668 VSS.n7336 VSS.n7335 2.2505
R5669 VSS.n7337 VSS.n2120 2.2505
R5670 VSS.n7339 VSS.n7338 2.2505
R5671 VSS.n7340 VSS.n2119 2.2505
R5672 VSS.n7342 VSS.n7341 2.2505
R5673 VSS.n7343 VSS.n2118 2.2505
R5674 VSS.n7345 VSS.n7344 2.2505
R5675 VSS.n7346 VSS.n2117 2.2505
R5676 VSS.n7348 VSS.n7347 2.2505
R5677 VSS.n7349 VSS.n2116 2.2505
R5678 VSS.n7351 VSS.n7350 2.2505
R5679 VSS.n7352 VSS.n2115 2.2505
R5680 VSS.n7354 VSS.n7353 2.2505
R5681 VSS.n7355 VSS.n2114 2.2505
R5682 VSS.n7357 VSS.n7356 2.2505
R5683 VSS.n7358 VSS.n2113 2.2505
R5684 VSS.n7360 VSS.n7359 2.2505
R5685 VSS.n7361 VSS.n2112 2.2505
R5686 VSS.n7363 VSS.n7362 2.2505
R5687 VSS.n7364 VSS.n2111 2.2505
R5688 VSS.n7366 VSS.n7365 2.2505
R5689 VSS.n7367 VSS.n2110 2.2505
R5690 VSS.n7369 VSS.n7368 2.2505
R5691 VSS.n7370 VSS.n2109 2.2505
R5692 VSS.n7372 VSS.n7371 2.2505
R5693 VSS.n7373 VSS.n2108 2.2505
R5694 VSS.n7375 VSS.n7374 2.2505
R5695 VSS.n7376 VSS.n2107 2.2505
R5696 VSS.n7378 VSS.n7377 2.2505
R5697 VSS.n7379 VSS.n2106 2.2505
R5698 VSS.n7381 VSS.n7380 2.2505
R5699 VSS.n7382 VSS.n2105 2.2505
R5700 VSS.n7384 VSS.n7383 2.2505
R5701 VSS.n7385 VSS.n2104 2.2505
R5702 VSS.n7387 VSS.n7386 2.2505
R5703 VSS.n7388 VSS.n2103 2.2505
R5704 VSS.n7390 VSS.n7389 2.2505
R5705 VSS.n7391 VSS.n2102 2.2505
R5706 VSS.n7393 VSS.n7392 2.2505
R5707 VSS.n7394 VSS.n2101 2.2505
R5708 VSS.n7396 VSS.n7395 2.2505
R5709 VSS.n7397 VSS.n2100 2.2505
R5710 VSS.n7399 VSS.n7398 2.2505
R5711 VSS.n7400 VSS.n2099 2.2505
R5712 VSS.n7402 VSS.n7401 2.2505
R5713 VSS.n7403 VSS.n2098 2.2505
R5714 VSS.n7405 VSS.n7404 2.2505
R5715 VSS.n7406 VSS.n2097 2.2505
R5716 VSS.n7408 VSS.n7407 2.2505
R5717 VSS.n7409 VSS.n2096 2.2505
R5718 VSS.n7411 VSS.n7410 2.2505
R5719 VSS.n7412 VSS.n2095 2.2505
R5720 VSS.n7414 VSS.n7413 2.2505
R5721 VSS.n7415 VSS.n2094 2.2505
R5722 VSS.n7417 VSS.n7416 2.2505
R5723 VSS.n7418 VSS.n2093 2.2505
R5724 VSS.n7420 VSS.n7419 2.2505
R5725 VSS.n7421 VSS.n2092 2.2505
R5726 VSS.n7423 VSS.n7422 2.2505
R5727 VSS.n7424 VSS.n2091 2.2505
R5728 VSS.n7426 VSS.n7425 2.2505
R5729 VSS.n7427 VSS.n2090 2.2505
R5730 VSS.n7429 VSS.n7428 2.2505
R5731 VSS.n7430 VSS.n2089 2.2505
R5732 VSS.n7432 VSS.n7431 2.2505
R5733 VSS.n7433 VSS.n2088 2.2505
R5734 VSS.n7435 VSS.n7434 2.2505
R5735 VSS.n7436 VSS.n2087 2.2505
R5736 VSS.n7438 VSS.n7437 2.2505
R5737 VSS.n7439 VSS.n2086 2.2505
R5738 VSS.n7441 VSS.n7440 2.2505
R5739 VSS.n7442 VSS.n2085 2.2505
R5740 VSS.n7444 VSS.n7443 2.2505
R5741 VSS.n7445 VSS.n2084 2.2505
R5742 VSS.n7447 VSS.n7446 2.2505
R5743 VSS.n7448 VSS.n2083 2.2505
R5744 VSS.n7450 VSS.n7449 2.2505
R5745 VSS.n7451 VSS.n2082 2.2505
R5746 VSS.n7453 VSS.n7452 2.2505
R5747 VSS.n7454 VSS.n2081 2.2505
R5748 VSS.n7456 VSS.n7455 2.2505
R5749 VSS.n7457 VSS.n2080 2.2505
R5750 VSS.n7459 VSS.n7458 2.2505
R5751 VSS.n7460 VSS.n2079 2.2505
R5752 VSS.n7462 VSS.n7461 2.2505
R5753 VSS.n7463 VSS.n2078 2.2505
R5754 VSS.n7465 VSS.n7464 2.2505
R5755 VSS.n7466 VSS.n2077 2.2505
R5756 VSS.n7468 VSS.n7467 2.2505
R5757 VSS.n7469 VSS.n2076 2.2505
R5758 VSS.n7471 VSS.n7470 2.2505
R5759 VSS.n7472 VSS.n2075 2.2505
R5760 VSS.n7474 VSS.n7473 2.2505
R5761 VSS.n7475 VSS.n2074 2.2505
R5762 VSS.n7477 VSS.n7476 2.2505
R5763 VSS.n7478 VSS.n2073 2.2505
R5764 VSS.n7480 VSS.n7479 2.2505
R5765 VSS.n7481 VSS.n2072 2.2505
R5766 VSS.n7483 VSS.n7482 2.2505
R5767 VSS.n7484 VSS.n2071 2.2505
R5768 VSS.n7486 VSS.n7485 2.2505
R5769 VSS.n7487 VSS.n2070 2.2505
R5770 VSS.n7489 VSS.n7488 2.2505
R5771 VSS.n7490 VSS.n2069 2.2505
R5772 VSS.n7492 VSS.n7491 2.2505
R5773 VSS.n7493 VSS.n2068 2.2505
R5774 VSS.n7495 VSS.n7494 2.2505
R5775 VSS.n7496 VSS.n2067 2.2505
R5776 VSS.n7498 VSS.n7497 2.2505
R5777 VSS.n7499 VSS.n2066 2.2505
R5778 VSS.n7501 VSS.n7500 2.2505
R5779 VSS.n7502 VSS.n2065 2.2505
R5780 VSS.n7504 VSS.n7503 2.2505
R5781 VSS.n7505 VSS.n2064 2.2505
R5782 VSS.n7507 VSS.n7506 2.2505
R5783 VSS.n7508 VSS.n2063 2.2505
R5784 VSS.n7510 VSS.n7509 2.2505
R5785 VSS.n7511 VSS.n2062 2.2505
R5786 VSS.n7513 VSS.n7512 2.2505
R5787 VSS.n7514 VSS.n2061 2.2505
R5788 VSS.n7516 VSS.n7515 2.2505
R5789 VSS.n7517 VSS.n2060 2.2505
R5790 VSS.n7519 VSS.n7518 2.2505
R5791 VSS.n7520 VSS.n2059 2.2505
R5792 VSS.n7522 VSS.n7521 2.2505
R5793 VSS.n7523 VSS.n2058 2.2505
R5794 VSS.n7525 VSS.n7524 2.2505
R5795 VSS.n7526 VSS.n2057 2.2505
R5796 VSS.n7528 VSS.n7527 2.2505
R5797 VSS.n7529 VSS.n2056 2.2505
R5798 VSS.n7531 VSS.n7530 2.2505
R5799 VSS.n7532 VSS.n2055 2.2505
R5800 VSS.n7534 VSS.n7533 2.2505
R5801 VSS.n7535 VSS.n2054 2.2505
R5802 VSS.n7537 VSS.n7536 2.2505
R5803 VSS.n7538 VSS.n2053 2.2505
R5804 VSS.n7540 VSS.n7539 2.2505
R5805 VSS.n7541 VSS.n2052 2.2505
R5806 VSS.n7543 VSS.n7542 2.2505
R5807 VSS.n7544 VSS.n2051 2.2505
R5808 VSS.n7546 VSS.n7545 2.2505
R5809 VSS.n7547 VSS.n2050 2.2505
R5810 VSS.n7549 VSS.n7548 2.2505
R5811 VSS.n7550 VSS.n2049 2.2505
R5812 VSS.n7552 VSS.n7551 2.2505
R5813 VSS.n7553 VSS.n2048 2.2505
R5814 VSS.n7555 VSS.n7554 2.2505
R5815 VSS.n7556 VSS.n2047 2.2505
R5816 VSS.n7558 VSS.n7557 2.2505
R5817 VSS.n7559 VSS.n2046 2.2505
R5818 VSS.n7561 VSS.n7560 2.2505
R5819 VSS.n7562 VSS.n2045 2.2505
R5820 VSS.n7564 VSS.n7563 2.2505
R5821 VSS.n7565 VSS.n2044 2.2505
R5822 VSS.n7567 VSS.n7566 2.2505
R5823 VSS.n7568 VSS.n2043 2.2505
R5824 VSS.n7570 VSS.n7569 2.2505
R5825 VSS.n7571 VSS.n2042 2.2505
R5826 VSS.n7573 VSS.n7572 2.2505
R5827 VSS.n7574 VSS.n2041 2.2505
R5828 VSS.n7576 VSS.n7575 2.2505
R5829 VSS.n7577 VSS.n2040 2.2505
R5830 VSS.n7579 VSS.n7578 2.2505
R5831 VSS.n7580 VSS.n2039 2.2505
R5832 VSS.n7582 VSS.n7581 2.2505
R5833 VSS.n7583 VSS.n2038 2.2505
R5834 VSS.n7585 VSS.n7584 2.2505
R5835 VSS.n7586 VSS.n2037 2.2505
R5836 VSS.n7588 VSS.n7587 2.2505
R5837 VSS.n7589 VSS.n2036 2.2505
R5838 VSS.n7591 VSS.n7590 2.2505
R5839 VSS.n7592 VSS.n2035 2.2505
R5840 VSS.n7594 VSS.n7593 2.2505
R5841 VSS.n7595 VSS.n2034 2.2505
R5842 VSS.n7597 VSS.n7596 2.2505
R5843 VSS.n7598 VSS.n2033 2.2505
R5844 VSS.n7600 VSS.n7599 2.2505
R5845 VSS.n7601 VSS.n2032 2.2505
R5846 VSS.n7603 VSS.n7602 2.2505
R5847 VSS.n7604 VSS.n2031 2.2505
R5848 VSS.n7606 VSS.n7605 2.2505
R5849 VSS.n7607 VSS.n2030 2.2505
R5850 VSS.n7609 VSS.n7608 2.2505
R5851 VSS.n7610 VSS.n2029 2.2505
R5852 VSS.n7612 VSS.n7611 2.2505
R5853 VSS.n7613 VSS.n2028 2.2505
R5854 VSS.n7615 VSS.n7614 2.2505
R5855 VSS.n7616 VSS.n2027 2.2505
R5856 VSS.n7618 VSS.n7617 2.2505
R5857 VSS.n7619 VSS.n2026 2.2505
R5858 VSS.n7621 VSS.n7620 2.2505
R5859 VSS.n7622 VSS.n2025 2.2505
R5860 VSS.n7624 VSS.n7623 2.2505
R5861 VSS.n7625 VSS.n2024 2.2505
R5862 VSS.n7627 VSS.n7626 2.2505
R5863 VSS.n7628 VSS.n2023 2.2505
R5864 VSS.n7630 VSS.n7629 2.2505
R5865 VSS.n7631 VSS.n2022 2.2505
R5866 VSS.n7633 VSS.n7632 2.2505
R5867 VSS.n7634 VSS.n2021 2.2505
R5868 VSS.n7636 VSS.n7635 2.2505
R5869 VSS.n7637 VSS.n2020 2.2505
R5870 VSS.n7639 VSS.n7638 2.2505
R5871 VSS.n7640 VSS.n2019 2.2505
R5872 VSS.n7642 VSS.n7641 2.2505
R5873 VSS.n7643 VSS.n2018 2.2505
R5874 VSS.n7645 VSS.n7644 2.2505
R5875 VSS.n7646 VSS.n2017 2.2505
R5876 VSS.n7648 VSS.n7647 2.2505
R5877 VSS.n7649 VSS.n2016 2.2505
R5878 VSS.n7651 VSS.n7650 2.2505
R5879 VSS.n7652 VSS.n2015 2.2505
R5880 VSS.n7654 VSS.n7653 2.2505
R5881 VSS.n7655 VSS.n2014 2.2505
R5882 VSS.n7657 VSS.n7656 2.2505
R5883 VSS.n7658 VSS.n2013 2.2505
R5884 VSS.n7660 VSS.n7659 2.2505
R5885 VSS.n7661 VSS.n2012 2.2505
R5886 VSS.n7663 VSS.n7662 2.2505
R5887 VSS.n7664 VSS.n2011 2.2505
R5888 VSS.n7666 VSS.n7665 2.2505
R5889 VSS.n7667 VSS.n2010 2.2505
R5890 VSS.n7669 VSS.n7668 2.2505
R5891 VSS.n7670 VSS.n2009 2.2505
R5892 VSS.n7672 VSS.n7671 2.2505
R5893 VSS.n7673 VSS.n2008 2.2505
R5894 VSS.n7675 VSS.n7674 2.2505
R5895 VSS.n7676 VSS.n2007 2.2505
R5896 VSS.n7678 VSS.n7677 2.2505
R5897 VSS.n7679 VSS.n2006 2.2505
R5898 VSS.n7681 VSS.n7680 2.2505
R5899 VSS.n7682 VSS.n2005 2.2505
R5900 VSS.n7684 VSS.n7683 2.2505
R5901 VSS.n7685 VSS.n2004 2.2505
R5902 VSS.n7687 VSS.n7686 2.2505
R5903 VSS.n7688 VSS.n2003 2.2505
R5904 VSS.n7690 VSS.n7689 2.2505
R5905 VSS.n7691 VSS.n2002 2.2505
R5906 VSS.n7693 VSS.n7692 2.2505
R5907 VSS.n7694 VSS.n2001 2.2505
R5908 VSS.n7696 VSS.n7695 2.2505
R5909 VSS.n7697 VSS.n2000 2.2505
R5910 VSS.n7699 VSS.n7698 2.2505
R5911 VSS.n7700 VSS.n1999 2.2505
R5912 VSS.n7702 VSS.n7701 2.2505
R5913 VSS.n7703 VSS.n1998 2.2505
R5914 VSS.n7705 VSS.n7704 2.2505
R5915 VSS.n7706 VSS.n1997 2.2505
R5916 VSS.n7708 VSS.n7707 2.2505
R5917 VSS.n7709 VSS.n1996 2.2505
R5918 VSS.n7711 VSS.n7710 2.2505
R5919 VSS.n7712 VSS.n1995 2.2505
R5920 VSS.n7714 VSS.n7713 2.2505
R5921 VSS.n7715 VSS.n1994 2.2505
R5922 VSS.n7717 VSS.n7716 2.2505
R5923 VSS.n7718 VSS.n1993 2.2505
R5924 VSS.n7720 VSS.n7719 2.2505
R5925 VSS.n7721 VSS.n1992 2.2505
R5926 VSS.n7723 VSS.n7722 2.2505
R5927 VSS.n7724 VSS.n1991 2.2505
R5928 VSS.n7726 VSS.n7725 2.2505
R5929 VSS.n7727 VSS.n1990 2.2505
R5930 VSS.n7729 VSS.n7728 2.2505
R5931 VSS.n7730 VSS.n1989 2.2505
R5932 VSS.n7732 VSS.n7731 2.2505
R5933 VSS.n7733 VSS.n1988 2.2505
R5934 VSS.n7735 VSS.n7734 2.2505
R5935 VSS.n7736 VSS.n1987 2.2505
R5936 VSS.n7738 VSS.n7737 2.2505
R5937 VSS.n7739 VSS.n1986 2.2505
R5938 VSS.n7741 VSS.n7740 2.2505
R5939 VSS.n7742 VSS.n1985 2.2505
R5940 VSS.n7744 VSS.n7743 2.2505
R5941 VSS.n7745 VSS.n1984 2.2505
R5942 VSS.n7747 VSS.n7746 2.2505
R5943 VSS.n7748 VSS.n1983 2.2505
R5944 VSS.n7750 VSS.n7749 2.2505
R5945 VSS.n7751 VSS.n1982 2.2505
R5946 VSS.n7753 VSS.n7752 2.2505
R5947 VSS.n7754 VSS.n1981 2.2505
R5948 VSS.n7756 VSS.n7755 2.2505
R5949 VSS.n7757 VSS.n1980 2.2505
R5950 VSS.n7759 VSS.n7758 2.2505
R5951 VSS.n7760 VSS.n1979 2.2505
R5952 VSS.n7762 VSS.n7761 2.2505
R5953 VSS.n7763 VSS.n1978 2.2505
R5954 VSS.n7765 VSS.n7764 2.2505
R5955 VSS.n7766 VSS.n1977 2.2505
R5956 VSS.n7768 VSS.n7767 2.2505
R5957 VSS.n7769 VSS.n1976 2.2505
R5958 VSS.n7771 VSS.n7770 2.2505
R5959 VSS.n7772 VSS.n1975 2.2505
R5960 VSS.n7774 VSS.n7773 2.2505
R5961 VSS.n7775 VSS.n1974 2.2505
R5962 VSS.n7777 VSS.n7776 2.2505
R5963 VSS.n7778 VSS.n1973 2.2505
R5964 VSS.n7780 VSS.n7779 2.2505
R5965 VSS.n7781 VSS.n1972 2.2505
R5966 VSS.n7783 VSS.n7782 2.2505
R5967 VSS.n7784 VSS.n1971 2.2505
R5968 VSS.n7786 VSS.n7785 2.2505
R5969 VSS.n7787 VSS.n1970 2.2505
R5970 VSS.n7789 VSS.n7788 2.2505
R5971 VSS.n7790 VSS.n1969 2.2505
R5972 VSS.n7792 VSS.n7791 2.2505
R5973 VSS.n7793 VSS.n1968 2.2505
R5974 VSS.n7795 VSS.n7794 2.2505
R5975 VSS.n7796 VSS.n1967 2.2505
R5976 VSS.n7798 VSS.n7797 2.2505
R5977 VSS.n7799 VSS.n1966 2.2505
R5978 VSS.n7801 VSS.n7800 2.2505
R5979 VSS.n7802 VSS.n1965 2.2505
R5980 VSS.n7804 VSS.n7803 2.2505
R5981 VSS.n7805 VSS.n1964 2.2505
R5982 VSS.n7807 VSS.n7806 2.2505
R5983 VSS.n7808 VSS.n1963 2.2505
R5984 VSS.n7810 VSS.n7809 2.2505
R5985 VSS.n7811 VSS.n1962 2.2505
R5986 VSS.n7813 VSS.n7812 2.2505
R5987 VSS.n7814 VSS.n1961 2.2505
R5988 VSS.n7816 VSS.n7815 2.2505
R5989 VSS.n7817 VSS.n1960 2.2505
R5990 VSS.n7819 VSS.n7818 2.2505
R5991 VSS.n7820 VSS.n1959 2.2505
R5992 VSS.n7822 VSS.n7821 2.2505
R5993 VSS.n7823 VSS.n1958 2.2505
R5994 VSS.n7825 VSS.n7824 2.2505
R5995 VSS.n7826 VSS.n1957 2.2505
R5996 VSS.n7828 VSS.n7827 2.2505
R5997 VSS.n7829 VSS.n1956 2.2505
R5998 VSS.n7831 VSS.n7830 2.2505
R5999 VSS.n7832 VSS.n1955 2.2505
R6000 VSS.n7834 VSS.n7833 2.2505
R6001 VSS.n7835 VSS.n1954 2.2505
R6002 VSS.n7837 VSS.n7836 2.2505
R6003 VSS.n7838 VSS.n1953 2.2505
R6004 VSS.n7840 VSS.n7839 2.2505
R6005 VSS.n7841 VSS.n1952 2.2505
R6006 VSS.n7843 VSS.n7842 2.2505
R6007 VSS.n7844 VSS.n1951 2.2505
R6008 VSS.n7846 VSS.n7845 2.2505
R6009 VSS.n7847 VSS.n1950 2.2505
R6010 VSS.n7849 VSS.n7848 2.2505
R6011 VSS.n7850 VSS.n1949 2.2505
R6012 VSS.n7852 VSS.n7851 2.2505
R6013 VSS.n7853 VSS.n1948 2.2505
R6014 VSS.n7855 VSS.n7854 2.2505
R6015 VSS.n7856 VSS.n1947 2.2505
R6016 VSS.n7858 VSS.n7857 2.2505
R6017 VSS.n7859 VSS.n1946 2.2505
R6018 VSS.n7861 VSS.n7860 2.2505
R6019 VSS.n7862 VSS.n1945 2.2505
R6020 VSS.n7864 VSS.n7863 2.2505
R6021 VSS.n7865 VSS.n1944 2.2505
R6022 VSS.n7867 VSS.n7866 2.2505
R6023 VSS.n7868 VSS.n1943 2.2505
R6024 VSS.n7870 VSS.n7869 2.2505
R6025 VSS.n7871 VSS.n1942 2.2505
R6026 VSS.n7873 VSS.n7872 2.2505
R6027 VSS.n7874 VSS.n1941 2.2505
R6028 VSS.n7876 VSS.n7875 2.2505
R6029 VSS.n7877 VSS.n1940 2.2505
R6030 VSS.n7879 VSS.n7878 2.2505
R6031 VSS.n7880 VSS.n1939 2.2505
R6032 VSS.n7882 VSS.n7881 2.2505
R6033 VSS.n7883 VSS.n1938 2.2505
R6034 VSS.n7885 VSS.n7884 2.2505
R6035 VSS.n7886 VSS.n1937 2.2505
R6036 VSS.n7888 VSS.n7887 2.2505
R6037 VSS.n7889 VSS.n1936 2.2505
R6038 VSS.n7891 VSS.n7890 2.2505
R6039 VSS.n7892 VSS.n1935 2.2505
R6040 VSS.n7894 VSS.n7893 2.2505
R6041 VSS.n7895 VSS.n1934 2.2505
R6042 VSS.n7897 VSS.n7896 2.2505
R6043 VSS.n7898 VSS.n1933 2.2505
R6044 VSS.n7900 VSS.n7899 2.2505
R6045 VSS.n7901 VSS.n1932 2.2505
R6046 VSS.n7903 VSS.n7902 2.2505
R6047 VSS.n7904 VSS.n1931 2.2505
R6048 VSS.n7906 VSS.n7905 2.2505
R6049 VSS.n7907 VSS.n1930 2.2505
R6050 VSS.n7909 VSS.n7908 2.2505
R6051 VSS.n7910 VSS.n1929 2.2505
R6052 VSS.n7912 VSS.n7911 2.2505
R6053 VSS.n7913 VSS.n1928 2.2505
R6054 VSS.n7915 VSS.n7914 2.2505
R6055 VSS.n7916 VSS.n1927 2.2505
R6056 VSS.n7918 VSS.n7917 2.2505
R6057 VSS.n7919 VSS.n1926 2.2505
R6058 VSS.n7921 VSS.n7920 2.2505
R6059 VSS.n7922 VSS.n1925 2.2505
R6060 VSS.n7924 VSS.n7923 2.2505
R6061 VSS.n7925 VSS.n1924 2.2505
R6062 VSS.n7927 VSS.n7926 2.2505
R6063 VSS.n7928 VSS.n1923 2.2505
R6064 VSS.n7930 VSS.n7929 2.2505
R6065 VSS.n7931 VSS.n1922 2.2505
R6066 VSS.n7933 VSS.n7932 2.2505
R6067 VSS.n7934 VSS.n1921 2.2505
R6068 VSS.n7936 VSS.n7935 2.2505
R6069 VSS.n7937 VSS.n1920 2.2505
R6070 VSS.n7939 VSS.n7938 2.2505
R6071 VSS.n7940 VSS.n1919 2.2505
R6072 VSS.n7942 VSS.n7941 2.2505
R6073 VSS.n7943 VSS.n1918 2.2505
R6074 VSS.n7945 VSS.n7944 2.2505
R6075 VSS.n7946 VSS.n1917 2.2505
R6076 VSS.n7948 VSS.n7947 2.2505
R6077 VSS.n7949 VSS.n1916 2.2505
R6078 VSS.n7951 VSS.n7950 2.2505
R6079 VSS.n7952 VSS.n1915 2.2505
R6080 VSS.n7954 VSS.n7953 2.2505
R6081 VSS.n7955 VSS.n1914 2.2505
R6082 VSS.n7957 VSS.n7956 2.2505
R6083 VSS.n7958 VSS.n1913 2.2505
R6084 VSS.n7960 VSS.n7959 2.2505
R6085 VSS.n7961 VSS.n1912 2.2505
R6086 VSS.n7963 VSS.n7962 2.2505
R6087 VSS.n7964 VSS.n1911 2.2505
R6088 VSS.n7966 VSS.n7965 2.2505
R6089 VSS.n7967 VSS.n1910 2.2505
R6090 VSS.n7969 VSS.n7968 2.2505
R6091 VSS.n7970 VSS.n1909 2.2505
R6092 VSS.n7972 VSS.n7971 2.2505
R6093 VSS.n7973 VSS.n1908 2.2505
R6094 VSS.n7975 VSS.n7974 2.2505
R6095 VSS.n7976 VSS.n1907 2.2505
R6096 VSS.n7978 VSS.n7977 2.2505
R6097 VSS.n7979 VSS.n1906 2.2505
R6098 VSS.n7981 VSS.n7980 2.2505
R6099 VSS.n7982 VSS.n1905 2.2505
R6100 VSS.n7984 VSS.n7983 2.2505
R6101 VSS.n7985 VSS.n1904 2.2505
R6102 VSS.n7987 VSS.n7986 2.2505
R6103 VSS.n7988 VSS.n1903 2.2505
R6104 VSS.n7990 VSS.n7989 2.2505
R6105 VSS.n7991 VSS.n1902 2.2505
R6106 VSS.n7993 VSS.n7992 2.2505
R6107 VSS.n7994 VSS.n1901 2.2505
R6108 VSS.n7996 VSS.n7995 2.2505
R6109 VSS.n7997 VSS.n1900 2.2505
R6110 VSS.n7999 VSS.n7998 2.2505
R6111 VSS.n8000 VSS.n1899 2.2505
R6112 VSS.n8002 VSS.n8001 2.2505
R6113 VSS.n8003 VSS.n1898 2.2505
R6114 VSS.n8005 VSS.n8004 2.2505
R6115 VSS.n8006 VSS.n1897 2.2505
R6116 VSS.n8008 VSS.n8007 2.2505
R6117 VSS.n8009 VSS.n1896 2.2505
R6118 VSS.n8011 VSS.n8010 2.2505
R6119 VSS.n8012 VSS.n1895 2.2505
R6120 VSS.n8014 VSS.n8013 2.2505
R6121 VSS.n8015 VSS.n1894 2.2505
R6122 VSS.n8017 VSS.n8016 2.2505
R6123 VSS.n8018 VSS.n1893 2.2505
R6124 VSS.n8020 VSS.n8019 2.2505
R6125 VSS.n8021 VSS.n1892 2.2505
R6126 VSS.n8023 VSS.n8022 2.2505
R6127 VSS.n8024 VSS.n1891 2.2505
R6128 VSS.n8026 VSS.n8025 2.2505
R6129 VSS.n8027 VSS.n1890 2.2505
R6130 VSS.n8029 VSS.n8028 2.2505
R6131 VSS.n8030 VSS.n1889 2.2505
R6132 VSS.n8032 VSS.n8031 2.2505
R6133 VSS.n8033 VSS.n1888 2.2505
R6134 VSS.n8035 VSS.n8034 2.2505
R6135 VSS.n8036 VSS.n1887 2.2505
R6136 VSS.n8038 VSS.n8037 2.2505
R6137 VSS.n8039 VSS.n1886 2.2505
R6138 VSS.n8041 VSS.n8040 2.2505
R6139 VSS.n8042 VSS.n1885 2.2505
R6140 VSS.n8044 VSS.n8043 2.2505
R6141 VSS.n8045 VSS.n1884 2.2505
R6142 VSS.n8047 VSS.n8046 2.2505
R6143 VSS.n8048 VSS.n1883 2.2505
R6144 VSS.n8050 VSS.n8049 2.2505
R6145 VSS.n8051 VSS.n1882 2.2505
R6146 VSS.n8053 VSS.n8052 2.2505
R6147 VSS.n8054 VSS.n1881 2.2505
R6148 VSS.n8056 VSS.n8055 2.2505
R6149 VSS.n8057 VSS.n1880 2.2505
R6150 VSS.n8059 VSS.n8058 2.2505
R6151 VSS.n8060 VSS.n1879 2.2505
R6152 VSS.n8062 VSS.n8061 2.2505
R6153 VSS.n8063 VSS.n1878 2.2505
R6154 VSS.n8065 VSS.n8064 2.2505
R6155 VSS.n8066 VSS.n1877 2.2505
R6156 VSS.n8068 VSS.n8067 2.2505
R6157 VSS.n8069 VSS.n1876 2.2505
R6158 VSS.n8071 VSS.n8070 2.2505
R6159 VSS.n8072 VSS.n1875 2.2505
R6160 VSS.n8074 VSS.n8073 2.2505
R6161 VSS.n8075 VSS.n1874 2.2505
R6162 VSS.n8077 VSS.n8076 2.2505
R6163 VSS.n8078 VSS.n1873 2.2505
R6164 VSS.n8080 VSS.n8079 2.2505
R6165 VSS.n8081 VSS.n1872 2.2505
R6166 VSS.n8083 VSS.n8082 2.2505
R6167 VSS.n8084 VSS.n1871 2.2505
R6168 VSS.n8086 VSS.n8085 2.2505
R6169 VSS.n8087 VSS.n1870 2.2505
R6170 VSS.n8089 VSS.n8088 2.2505
R6171 VSS.n8090 VSS.n1869 2.2505
R6172 VSS.n8092 VSS.n8091 2.2505
R6173 VSS.n8093 VSS.n1868 2.2505
R6174 VSS.n8095 VSS.n8094 2.2505
R6175 VSS.n8096 VSS.n1867 2.2505
R6176 VSS.n8098 VSS.n8097 2.2505
R6177 VSS.n8099 VSS.n1866 2.2505
R6178 VSS.n8101 VSS.n8100 2.2505
R6179 VSS.n8102 VSS.n1865 2.2505
R6180 VSS.n8104 VSS.n8103 2.2505
R6181 VSS.n8105 VSS.n1864 2.2505
R6182 VSS.n8107 VSS.n8106 2.2505
R6183 VSS.n8108 VSS.n1863 2.2505
R6184 VSS.n8110 VSS.n8109 2.2505
R6185 VSS.n8111 VSS.n1862 2.2505
R6186 VSS.n8113 VSS.n8112 2.2505
R6187 VSS.n8114 VSS.n1861 2.2505
R6188 VSS.n8116 VSS.n8115 2.2505
R6189 VSS.n8117 VSS.n1860 2.2505
R6190 VSS.n8119 VSS.n8118 2.2505
R6191 VSS.n8120 VSS.n1859 2.2505
R6192 VSS.n8122 VSS.n8121 2.2505
R6193 VSS.n8123 VSS.n1858 2.2505
R6194 VSS.n8125 VSS.n8124 2.2505
R6195 VSS.n8126 VSS.n1857 2.2505
R6196 VSS.n8128 VSS.n8127 2.2505
R6197 VSS.n8129 VSS.n1856 2.2505
R6198 VSS.n8131 VSS.n8130 2.2505
R6199 VSS.n8132 VSS.n1855 2.2505
R6200 VSS.n8134 VSS.n8133 2.2505
R6201 VSS.n8135 VSS.n1854 2.2505
R6202 VSS.n8137 VSS.n8136 2.2505
R6203 VSS.n8138 VSS.n1853 2.2505
R6204 VSS.n8140 VSS.n8139 2.2505
R6205 VSS.n8141 VSS.n1852 2.2505
R6206 VSS.n8143 VSS.n8142 2.2505
R6207 VSS.n8144 VSS.n1851 2.2505
R6208 VSS.n8146 VSS.n8145 2.2505
R6209 VSS.n8147 VSS.n1850 2.2505
R6210 VSS.n8149 VSS.n8148 2.2505
R6211 VSS.n8150 VSS.n1849 2.2505
R6212 VSS.n8152 VSS.n8151 2.2505
R6213 VSS.n8153 VSS.n1848 2.2505
R6214 VSS.n8155 VSS.n8154 2.2505
R6215 VSS.n8156 VSS.n1847 2.2505
R6216 VSS.n8158 VSS.n8157 2.2505
R6217 VSS.n8159 VSS.n1846 2.2505
R6218 VSS.n8161 VSS.n8160 2.2505
R6219 VSS.n8162 VSS.n1845 2.2505
R6220 VSS.n8164 VSS.n8163 2.2505
R6221 VSS.n8165 VSS.n1844 2.2505
R6222 VSS.n8167 VSS.n8166 2.2505
R6223 VSS.n8168 VSS.n1843 2.2505
R6224 VSS.n8170 VSS.n8169 2.2505
R6225 VSS.n8171 VSS.n1842 2.2505
R6226 VSS.n8173 VSS.n8172 2.2505
R6227 VSS.n8174 VSS.n1841 2.2505
R6228 VSS.n8176 VSS.n8175 2.2505
R6229 VSS.n8177 VSS.n1840 2.2505
R6230 VSS.n8179 VSS.n8178 2.2505
R6231 VSS.n8180 VSS.n1839 2.2505
R6232 VSS.n8182 VSS.n8181 2.2505
R6233 VSS.n8183 VSS.n1838 2.2505
R6234 VSS.n8185 VSS.n8184 2.2505
R6235 VSS.n8186 VSS.n1837 2.2505
R6236 VSS.n8188 VSS.n8187 2.2505
R6237 VSS.n8189 VSS.n1836 2.2505
R6238 VSS.n8191 VSS.n8190 2.2505
R6239 VSS.n8192 VSS.n1835 2.2505
R6240 VSS.n8194 VSS.n8193 2.2505
R6241 VSS.n8195 VSS.n1834 2.2505
R6242 VSS.n8197 VSS.n8196 2.2505
R6243 VSS.n8198 VSS.n1833 2.2505
R6244 VSS.n8200 VSS.n8199 2.2505
R6245 VSS.n8201 VSS.n1832 2.2505
R6246 VSS.n8203 VSS.n8202 2.2505
R6247 VSS.n8204 VSS.n1831 2.2505
R6248 VSS.n8206 VSS.n8205 2.2505
R6249 VSS.n8207 VSS.n1830 2.2505
R6250 VSS.n8209 VSS.n8208 2.2505
R6251 VSS.n8210 VSS.n1829 2.2505
R6252 VSS.n8212 VSS.n8211 2.2505
R6253 VSS.n8213 VSS.n1828 2.2505
R6254 VSS.n8215 VSS.n8214 2.2505
R6255 VSS.n8216 VSS.n1827 2.2505
R6256 VSS.n8218 VSS.n8217 2.2505
R6257 VSS.n8219 VSS.n1826 2.2505
R6258 VSS.n8221 VSS.n8220 2.2505
R6259 VSS.n8222 VSS.n1825 2.2505
R6260 VSS.n8224 VSS.n8223 2.2505
R6261 VSS.n8225 VSS.n1824 2.2505
R6262 VSS.n8227 VSS.n8226 2.2505
R6263 VSS.n8228 VSS.n1823 2.2505
R6264 VSS.n8230 VSS.n8229 2.2505
R6265 VSS.n8231 VSS.n1822 2.2505
R6266 VSS.n4141 VSS.n4140 2.2505
R6267 VSS.n4139 VSS.n3185 2.2505
R6268 VSS.n4138 VSS.n4137 2.2505
R6269 VSS.n4136 VSS.n3186 2.2505
R6270 VSS.n4135 VSS.n4134 2.2505
R6271 VSS.n4133 VSS.n3187 2.2505
R6272 VSS.n4132 VSS.n4131 2.2505
R6273 VSS.n4130 VSS.n3188 2.2505
R6274 VSS.n4129 VSS.n4128 2.2505
R6275 VSS.n4127 VSS.n3189 2.2505
R6276 VSS.n4126 VSS.n4125 2.2505
R6277 VSS.n4124 VSS.n3190 2.2505
R6278 VSS.n4123 VSS.n4122 2.2505
R6279 VSS.n4121 VSS.n3191 2.2505
R6280 VSS.n4120 VSS.n4119 2.2505
R6281 VSS.n4118 VSS.n3192 2.2505
R6282 VSS.n4117 VSS.n4116 2.2505
R6283 VSS.n4115 VSS.n3193 2.2505
R6284 VSS.n4114 VSS.n4113 2.2505
R6285 VSS.n4112 VSS.n3194 2.2505
R6286 VSS.n4111 VSS.n4110 2.2505
R6287 VSS.n4109 VSS.n3195 2.2505
R6288 VSS.n4108 VSS.n4107 2.2505
R6289 VSS.n4106 VSS.n3196 2.2505
R6290 VSS.n4105 VSS.n4104 2.2505
R6291 VSS.n4103 VSS.n3197 2.2505
R6292 VSS.n4102 VSS.n4101 2.2505
R6293 VSS.n4100 VSS.n3198 2.2505
R6294 VSS.n4099 VSS.n4098 2.2505
R6295 VSS.n4097 VSS.n3199 2.2505
R6296 VSS.n4096 VSS.n4095 2.2505
R6297 VSS.n4094 VSS.n3200 2.2505
R6298 VSS.n4093 VSS.n4092 2.2505
R6299 VSS.n4091 VSS.n3201 2.2505
R6300 VSS.n4090 VSS.n4089 2.2505
R6301 VSS.n4088 VSS.n3202 2.2505
R6302 VSS.n4087 VSS.n4086 2.2505
R6303 VSS.n4085 VSS.n3203 2.2505
R6304 VSS.n4084 VSS.n4083 2.2505
R6305 VSS.n4082 VSS.n3204 2.2505
R6306 VSS.n4081 VSS.n4080 2.2505
R6307 VSS.n4079 VSS.n3205 2.2505
R6308 VSS.n4078 VSS.n4077 2.2505
R6309 VSS.n4076 VSS.n3206 2.2505
R6310 VSS.n4075 VSS.n4074 2.2505
R6311 VSS.n4073 VSS.n3207 2.2505
R6312 VSS.n4072 VSS.n4071 2.2505
R6313 VSS.n4070 VSS.n3208 2.2505
R6314 VSS.n4069 VSS.n4068 2.2505
R6315 VSS.n4067 VSS.n3209 2.2505
R6316 VSS.n4066 VSS.n4065 2.2505
R6317 VSS.n4064 VSS.n3210 2.2505
R6318 VSS.n4063 VSS.n4062 2.2505
R6319 VSS.n4061 VSS.n3211 2.2505
R6320 VSS.n4060 VSS.n4059 2.2505
R6321 VSS.n4058 VSS.n3212 2.2505
R6322 VSS.n4057 VSS.n4056 2.2505
R6323 VSS.n4055 VSS.n3213 2.2505
R6324 VSS.n4054 VSS.n4053 2.2505
R6325 VSS.n4052 VSS.n3214 2.2505
R6326 VSS.n4051 VSS.n4050 2.2505
R6327 VSS.n4049 VSS.n3215 2.2505
R6328 VSS.n4048 VSS.n4047 2.2505
R6329 VSS.n4046 VSS.n3216 2.2505
R6330 VSS.n4045 VSS.n4044 2.2505
R6331 VSS.n4043 VSS.n3217 2.2505
R6332 VSS.n4042 VSS.n4041 2.2505
R6333 VSS.n4040 VSS.n3218 2.2505
R6334 VSS.n4039 VSS.n4038 2.2505
R6335 VSS.n4037 VSS.n3219 2.2505
R6336 VSS.n4036 VSS.n4035 2.2505
R6337 VSS.n4034 VSS.n3220 2.2505
R6338 VSS.n4033 VSS.n4032 2.2505
R6339 VSS.n4031 VSS.n3221 2.2505
R6340 VSS.n4030 VSS.n4029 2.2505
R6341 VSS.n4028 VSS.n3222 2.2505
R6342 VSS.n4027 VSS.n4026 2.2505
R6343 VSS.n4025 VSS.n3223 2.2505
R6344 VSS.n4024 VSS.n4023 2.2505
R6345 VSS.n4022 VSS.n3224 2.2505
R6346 VSS.n4021 VSS.n4020 2.2505
R6347 VSS.n4019 VSS.n3225 2.2505
R6348 VSS.n4018 VSS.n4017 2.2505
R6349 VSS.n4016 VSS.n3226 2.2505
R6350 VSS.n4015 VSS.n4014 2.2505
R6351 VSS.n4013 VSS.n3227 2.2505
R6352 VSS.n4012 VSS.n4011 2.2505
R6353 VSS.n4010 VSS.n3228 2.2505
R6354 VSS.n4009 VSS.n4008 2.2505
R6355 VSS.n4007 VSS.n3229 2.2505
R6356 VSS.n4006 VSS.n4005 2.2505
R6357 VSS.n4004 VSS.n3230 2.2505
R6358 VSS.n4003 VSS.n4002 2.2505
R6359 VSS.n4001 VSS.n3231 2.2505
R6360 VSS.n4000 VSS.n3999 2.2505
R6361 VSS.n3998 VSS.n3232 2.2505
R6362 VSS.n3997 VSS.n3996 2.2505
R6363 VSS.n3995 VSS.n3233 2.2505
R6364 VSS.n3994 VSS.n3993 2.2505
R6365 VSS.n3992 VSS.n3234 2.2505
R6366 VSS.n3991 VSS.n3990 2.2505
R6367 VSS.n3989 VSS.n3235 2.2505
R6368 VSS.n3988 VSS.n3987 2.2505
R6369 VSS.n3986 VSS.n3236 2.2505
R6370 VSS.n3985 VSS.n3984 2.2505
R6371 VSS.n3983 VSS.n3237 2.2505
R6372 VSS.n3982 VSS.n3981 2.2505
R6373 VSS.n3980 VSS.n3238 2.2505
R6374 VSS.n3979 VSS.n3978 2.2505
R6375 VSS.n3977 VSS.n3239 2.2505
R6376 VSS.n3976 VSS.n3975 2.2505
R6377 VSS.n3974 VSS.n3240 2.2505
R6378 VSS.n3973 VSS.n3972 2.2505
R6379 VSS.n3971 VSS.n3241 2.2505
R6380 VSS.n3970 VSS.n3969 2.2505
R6381 VSS.n3968 VSS.n3242 2.2505
R6382 VSS.n3967 VSS.n3966 2.2505
R6383 VSS.n3965 VSS.n3243 2.2505
R6384 VSS.n3964 VSS.n3963 2.2505
R6385 VSS.n3962 VSS.n3244 2.2505
R6386 VSS.n3961 VSS.n3960 2.2505
R6387 VSS.n3959 VSS.n3245 2.2505
R6388 VSS.n3958 VSS.n3957 2.2505
R6389 VSS.n3956 VSS.n3246 2.2505
R6390 VSS.n3955 VSS.n3954 2.2505
R6391 VSS.n3953 VSS.n3247 2.2505
R6392 VSS.n3952 VSS.n3951 2.2505
R6393 VSS.n3950 VSS.n3248 2.2505
R6394 VSS.n3949 VSS.n3948 2.2505
R6395 VSS.n3947 VSS.n3249 2.2505
R6396 VSS.n3946 VSS.n3945 2.2505
R6397 VSS.n3944 VSS.n3250 2.2505
R6398 VSS.n3943 VSS.n3942 2.2505
R6399 VSS.n3941 VSS.n3251 2.2505
R6400 VSS.n3940 VSS.n3939 2.2505
R6401 VSS.n3938 VSS.n3252 2.2505
R6402 VSS.n3937 VSS.n3936 2.2505
R6403 VSS.n3935 VSS.n3253 2.2505
R6404 VSS.n3934 VSS.n3933 2.2505
R6405 VSS.n3932 VSS.n3254 2.2505
R6406 VSS.n3931 VSS.n3930 2.2505
R6407 VSS.n3929 VSS.n3255 2.2505
R6408 VSS.n3928 VSS.n3927 2.2505
R6409 VSS.n3926 VSS.n3256 2.2505
R6410 VSS.n3925 VSS.n3924 2.2505
R6411 VSS.n3923 VSS.n3257 2.2505
R6412 VSS.n3922 VSS.n3921 2.2505
R6413 VSS.n3920 VSS.n3258 2.2505
R6414 VSS.n3919 VSS.n3918 2.2505
R6415 VSS.n3917 VSS.n3259 2.2505
R6416 VSS.n3916 VSS.n3915 2.2505
R6417 VSS.n3914 VSS.n3260 2.2505
R6418 VSS.n3913 VSS.n3912 2.2505
R6419 VSS.n3911 VSS.n3261 2.2505
R6420 VSS.n3910 VSS.n3909 2.2505
R6421 VSS.n3908 VSS.n3262 2.2505
R6422 VSS.n3907 VSS.n3906 2.2505
R6423 VSS.n3905 VSS.n3263 2.2505
R6424 VSS.n3904 VSS.n3903 2.2505
R6425 VSS.n3902 VSS.n3264 2.2505
R6426 VSS.n3901 VSS.n3900 2.2505
R6427 VSS.n3899 VSS.n3265 2.2505
R6428 VSS.n3898 VSS.n3897 2.2505
R6429 VSS.n3896 VSS.n3266 2.2505
R6430 VSS.n3895 VSS.n3894 2.2505
R6431 VSS.n3893 VSS.n3267 2.2505
R6432 VSS.n3892 VSS.n3891 2.2505
R6433 VSS.n3890 VSS.n3268 2.2505
R6434 VSS.n3889 VSS.n3888 2.2505
R6435 VSS.n3887 VSS.n3269 2.2505
R6436 VSS.n3886 VSS.n3885 2.2505
R6437 VSS.n3884 VSS.n3270 2.2505
R6438 VSS.n3883 VSS.n3882 2.2505
R6439 VSS.n3881 VSS.n3271 2.2505
R6440 VSS.n3880 VSS.n3879 2.2505
R6441 VSS.n3878 VSS.n3272 2.2505
R6442 VSS.n3877 VSS.n3876 2.2505
R6443 VSS.n3875 VSS.n3273 2.2505
R6444 VSS.n3874 VSS.n3873 2.2505
R6445 VSS.n3872 VSS.n3274 2.2505
R6446 VSS.n3871 VSS.n3870 2.2505
R6447 VSS.n3869 VSS.n3275 2.2505
R6448 VSS.n3868 VSS.n3867 2.2505
R6449 VSS.n3866 VSS.n3276 2.2505
R6450 VSS.n3865 VSS.n3864 2.2505
R6451 VSS.n3863 VSS.n3277 2.2505
R6452 VSS.n3862 VSS.n3861 2.2505
R6453 VSS.n3860 VSS.n3278 2.2505
R6454 VSS.n3859 VSS.n3858 2.2505
R6455 VSS.n3857 VSS.n3279 2.2505
R6456 VSS.n3856 VSS.n3855 2.2505
R6457 VSS.n3854 VSS.n3280 2.2505
R6458 VSS.n3853 VSS.n3852 2.2505
R6459 VSS.n3851 VSS.n3281 2.2505
R6460 VSS.n3850 VSS.n3849 2.2505
R6461 VSS.n3848 VSS.n3282 2.2505
R6462 VSS.n3847 VSS.n3846 2.2505
R6463 VSS.n3845 VSS.n3283 2.2505
R6464 VSS.n3844 VSS.n3843 2.2505
R6465 VSS.n3842 VSS.n3284 2.2505
R6466 VSS.n3841 VSS.n3840 2.2505
R6467 VSS.n3839 VSS.n3285 2.2505
R6468 VSS.n3838 VSS.n3837 2.2505
R6469 VSS.n3836 VSS.n3286 2.2505
R6470 VSS.n3835 VSS.n3834 2.2505
R6471 VSS.n3833 VSS.n3287 2.2505
R6472 VSS.n3832 VSS.n3831 2.2505
R6473 VSS.n3830 VSS.n3288 2.2505
R6474 VSS.n3829 VSS.n3828 2.2505
R6475 VSS.n3827 VSS.n3289 2.2505
R6476 VSS.n3826 VSS.n3825 2.2505
R6477 VSS.n3824 VSS.n3290 2.2505
R6478 VSS.n3823 VSS.n3822 2.2505
R6479 VSS.n3821 VSS.n3291 2.2505
R6480 VSS.n3820 VSS.n3819 2.2505
R6481 VSS.n3818 VSS.n3292 2.2505
R6482 VSS.n3817 VSS.n3816 2.2505
R6483 VSS.n3815 VSS.n3293 2.2505
R6484 VSS.n3814 VSS.n3813 2.2505
R6485 VSS.n3812 VSS.n3294 2.2505
R6486 VSS.n3811 VSS.n3810 2.2505
R6487 VSS.n3809 VSS.n3295 2.2505
R6488 VSS.n3808 VSS.n3807 2.2505
R6489 VSS.n3806 VSS.n3296 2.2505
R6490 VSS.n3805 VSS.n3804 2.2505
R6491 VSS.n3803 VSS.n3297 2.2505
R6492 VSS.n3802 VSS.n3801 2.2505
R6493 VSS.n3800 VSS.n3298 2.2505
R6494 VSS.n3799 VSS.n3798 2.2505
R6495 VSS.n3797 VSS.n3299 2.2505
R6496 VSS.n3796 VSS.n3795 2.2505
R6497 VSS.n3794 VSS.n3300 2.2505
R6498 VSS.n3793 VSS.n3792 2.2505
R6499 VSS.n3791 VSS.n3301 2.2505
R6500 VSS.n3790 VSS.n3789 2.2505
R6501 VSS.n3788 VSS.n3302 2.2505
R6502 VSS.n3787 VSS.n3786 2.2505
R6503 VSS.n3785 VSS.n3303 2.2505
R6504 VSS.n3784 VSS.n3783 2.2505
R6505 VSS.n3782 VSS.n3304 2.2505
R6506 VSS.n3781 VSS.n3780 2.2505
R6507 VSS.n3779 VSS.n3305 2.2505
R6508 VSS.n3778 VSS.n3777 2.2505
R6509 VSS.n3776 VSS.n3306 2.2505
R6510 VSS.n3775 VSS.n3774 2.2505
R6511 VSS.n3773 VSS.n3307 2.2505
R6512 VSS.n3772 VSS.n3771 2.2505
R6513 VSS.n3770 VSS.n3308 2.2505
R6514 VSS.n3769 VSS.n3768 2.2505
R6515 VSS.n3767 VSS.n3309 2.2505
R6516 VSS.n3766 VSS.n3765 2.2505
R6517 VSS.n3764 VSS.n3310 2.2505
R6518 VSS.n3763 VSS.n3762 2.2505
R6519 VSS.n3761 VSS.n3311 2.2505
R6520 VSS.n3760 VSS.n3759 2.2505
R6521 VSS.n3758 VSS.n3312 2.2505
R6522 VSS.n3757 VSS.n3756 2.2505
R6523 VSS.n3755 VSS.n3313 2.2505
R6524 VSS.n3754 VSS.n3753 2.2505
R6525 VSS.n3752 VSS.n3314 2.2505
R6526 VSS.n3751 VSS.n3750 2.2505
R6527 VSS.n3749 VSS.n3315 2.2505
R6528 VSS.n3748 VSS.n3747 2.2505
R6529 VSS.n3746 VSS.n3316 2.2505
R6530 VSS.n3745 VSS.n3744 2.2505
R6531 VSS.n3743 VSS.n3317 2.2505
R6532 VSS.n3742 VSS.n3741 2.2505
R6533 VSS.n3740 VSS.n3318 2.2505
R6534 VSS.n3739 VSS.n3738 2.2505
R6535 VSS.n3737 VSS.n3319 2.2505
R6536 VSS.n3736 VSS.n3735 2.2505
R6537 VSS.n3734 VSS.n3320 2.2505
R6538 VSS.n3733 VSS.n3732 2.2505
R6539 VSS.n3731 VSS.n3321 2.2505
R6540 VSS.n3730 VSS.n3729 2.2505
R6541 VSS.n3728 VSS.n3322 2.2505
R6542 VSS.n3727 VSS.n3726 2.2505
R6543 VSS.n3725 VSS.n3323 2.2505
R6544 VSS.n3724 VSS.n3723 2.2505
R6545 VSS.n3722 VSS.n3324 2.2505
R6546 VSS.n3721 VSS.n3720 2.2505
R6547 VSS.n3719 VSS.n3325 2.2505
R6548 VSS.n3718 VSS.n3717 2.2505
R6549 VSS.n3716 VSS.n3326 2.2505
R6550 VSS.n3715 VSS.n3714 2.2505
R6551 VSS.n3713 VSS.n3327 2.2505
R6552 VSS.n3712 VSS.n3711 2.2505
R6553 VSS.n3710 VSS.n3328 2.2505
R6554 VSS.n3709 VSS.n3708 2.2505
R6555 VSS.n3707 VSS.n3329 2.2505
R6556 VSS.n3706 VSS.n3705 2.2505
R6557 VSS.n3704 VSS.n3330 2.2505
R6558 VSS.n3703 VSS.n3702 2.2505
R6559 VSS.n3701 VSS.n3331 2.2505
R6560 VSS.n3700 VSS.n3699 2.2505
R6561 VSS.n3698 VSS.n3332 2.2505
R6562 VSS.n3697 VSS.n3696 2.2505
R6563 VSS.n3695 VSS.n3333 2.2505
R6564 VSS.n3694 VSS.n3693 2.2505
R6565 VSS.n3692 VSS.n3334 2.2505
R6566 VSS.n3691 VSS.n3690 2.2505
R6567 VSS.n3689 VSS.n3335 2.2505
R6568 VSS.n3688 VSS.n3687 2.2505
R6569 VSS.n3686 VSS.n3336 2.2505
R6570 VSS.n3685 VSS.n3684 2.2505
R6571 VSS.n3683 VSS.n3337 2.2505
R6572 VSS.n3682 VSS.n3681 2.2505
R6573 VSS.n3680 VSS.n3338 2.2505
R6574 VSS.n3679 VSS.n3678 2.2505
R6575 VSS.n3677 VSS.n3339 2.2505
R6576 VSS.n3676 VSS.n3675 2.2505
R6577 VSS.n3674 VSS.n3340 2.2505
R6578 VSS.n3673 VSS.n3672 2.2505
R6579 VSS.n3671 VSS.n3341 2.2505
R6580 VSS.n3670 VSS.n3669 2.2505
R6581 VSS.n3668 VSS.n3342 2.2505
R6582 VSS.n3667 VSS.n3666 2.2505
R6583 VSS.n3665 VSS.n3343 2.2505
R6584 VSS.n3664 VSS.n3663 2.2505
R6585 VSS.n3662 VSS.n3344 2.2505
R6586 VSS.n3661 VSS.n3660 2.2505
R6587 VSS.n3659 VSS.n3345 2.2505
R6588 VSS.n3658 VSS.n3657 2.2505
R6589 VSS.n3656 VSS.n3346 2.2505
R6590 VSS.n3655 VSS.n3654 2.2505
R6591 VSS.n3653 VSS.n3347 2.2505
R6592 VSS.n3652 VSS.n3651 2.2505
R6593 VSS.n3650 VSS.n3348 2.2505
R6594 VSS.n3649 VSS.n3648 2.2505
R6595 VSS.n3647 VSS.n3349 2.2505
R6596 VSS.n3646 VSS.n3645 2.2505
R6597 VSS.n3644 VSS.n3350 2.2505
R6598 VSS.n3643 VSS.n3642 2.2505
R6599 VSS.n3641 VSS.n3351 2.2505
R6600 VSS.n3640 VSS.n3639 2.2505
R6601 VSS.n3638 VSS.n3352 2.2505
R6602 VSS.n3637 VSS.n3636 2.2505
R6603 VSS.n3635 VSS.n3353 2.2505
R6604 VSS.n3634 VSS.n3633 2.2505
R6605 VSS.n3632 VSS.n3354 2.2505
R6606 VSS.n3631 VSS.n3630 2.2505
R6607 VSS.n3629 VSS.n3355 2.2505
R6608 VSS.n3628 VSS.n3627 2.2505
R6609 VSS.n3626 VSS.n3356 2.2505
R6610 VSS.n3625 VSS.n3624 2.2505
R6611 VSS.n3623 VSS.n3357 2.2505
R6612 VSS.n3622 VSS.n3621 2.2505
R6613 VSS.n3620 VSS.n3358 2.2505
R6614 VSS.n3619 VSS.n3618 2.2505
R6615 VSS.n3617 VSS.n3359 2.2505
R6616 VSS.n3616 VSS.n3615 2.2505
R6617 VSS.n3614 VSS.n3360 2.2505
R6618 VSS.n3613 VSS.n3612 2.2505
R6619 VSS.n3611 VSS.n3361 2.2505
R6620 VSS.n3610 VSS.n3609 2.2505
R6621 VSS.n3608 VSS.n3362 2.2505
R6622 VSS.n3607 VSS.n3606 2.2505
R6623 VSS.n3605 VSS.n3363 2.2505
R6624 VSS.n3604 VSS.n3603 2.2505
R6625 VSS.n3602 VSS.n3364 2.2505
R6626 VSS.n3601 VSS.n3600 2.2505
R6627 VSS.n3599 VSS.n3365 2.2505
R6628 VSS.n3598 VSS.n3597 2.2505
R6629 VSS.n3596 VSS.n3366 2.2505
R6630 VSS.n3595 VSS.n3594 2.2505
R6631 VSS.n3593 VSS.n3367 2.2505
R6632 VSS.n3592 VSS.n3591 2.2505
R6633 VSS.n3590 VSS.n3368 2.2505
R6634 VSS.n3589 VSS.n3588 2.2505
R6635 VSS.n3587 VSS.n3369 2.2505
R6636 VSS.n3586 VSS.n3585 2.2505
R6637 VSS.n3584 VSS.n3370 2.2505
R6638 VSS.n3583 VSS.n3582 2.2505
R6639 VSS.n3581 VSS.n3371 2.2505
R6640 VSS.n3580 VSS.n3579 2.2505
R6641 VSS.n3578 VSS.n3372 2.2505
R6642 VSS.n3577 VSS.n3576 2.2505
R6643 VSS.n3575 VSS.n3373 2.2505
R6644 VSS.n3574 VSS.n3573 2.2505
R6645 VSS.n3572 VSS.n3374 2.2505
R6646 VSS.n3571 VSS.n3570 2.2505
R6647 VSS.n3569 VSS.n3375 2.2505
R6648 VSS.n3568 VSS.n3567 2.2505
R6649 VSS.n3566 VSS.n3376 2.2505
R6650 VSS.n3565 VSS.n3564 2.2505
R6651 VSS.n3563 VSS.n3377 2.2505
R6652 VSS.n3562 VSS.n3561 2.2505
R6653 VSS.n3560 VSS.n3378 2.2505
R6654 VSS.n3559 VSS.n3558 2.2505
R6655 VSS.n3557 VSS.n3379 2.2505
R6656 VSS.n3556 VSS.n3555 2.2505
R6657 VSS.n3554 VSS.n3380 2.2505
R6658 VSS.n3553 VSS.n3552 2.2505
R6659 VSS.n3551 VSS.n3381 2.2505
R6660 VSS.n3550 VSS.n3549 2.2505
R6661 VSS.n3548 VSS.n3382 2.2505
R6662 VSS.n3547 VSS.n3546 2.2505
R6663 VSS.n3545 VSS.n3383 2.2505
R6664 VSS.n3544 VSS.n3543 2.2505
R6665 VSS.n3542 VSS.n3384 2.2505
R6666 VSS.n3541 VSS.n3540 2.2505
R6667 VSS.n3539 VSS.n3385 2.2505
R6668 VSS.n3538 VSS.n3537 2.2505
R6669 VSS.n3536 VSS.n3386 2.2505
R6670 VSS.n3535 VSS.n3534 2.2505
R6671 VSS.n3533 VSS.n3387 2.2505
R6672 VSS.n3532 VSS.n3531 2.2505
R6673 VSS.n3530 VSS.n3388 2.2505
R6674 VSS.n3529 VSS.n3528 2.2505
R6675 VSS.n3527 VSS.n3389 2.2505
R6676 VSS.n3526 VSS.n3525 2.2505
R6677 VSS.n3524 VSS.n3390 2.2505
R6678 VSS.n3523 VSS.n3522 2.2505
R6679 VSS.n3521 VSS.n3391 2.2505
R6680 VSS.n3520 VSS.n3519 2.2505
R6681 VSS.n3518 VSS.n3392 2.2505
R6682 VSS.n3517 VSS.n3516 2.2505
R6683 VSS.n3515 VSS.n3393 2.2505
R6684 VSS.n3514 VSS.n3513 2.2505
R6685 VSS.n3512 VSS.n3394 2.2505
R6686 VSS.n3511 VSS.n3510 2.2505
R6687 VSS.n3509 VSS.n3395 2.2505
R6688 VSS.n3508 VSS.n3507 2.2505
R6689 VSS.n3506 VSS.n3396 2.2505
R6690 VSS.n3505 VSS.n3504 2.2505
R6691 VSS.n3503 VSS.n3397 2.2505
R6692 VSS.n3502 VSS.n3501 2.2505
R6693 VSS.n3500 VSS.n3398 2.2505
R6694 VSS.n3499 VSS.n3498 2.2505
R6695 VSS.n3497 VSS.n3399 2.2505
R6696 VSS.n3496 VSS.n3495 2.2505
R6697 VSS.n3494 VSS.n3400 2.2505
R6698 VSS.n3493 VSS.n3492 2.2505
R6699 VSS.n3491 VSS.n3401 2.2505
R6700 VSS.n3490 VSS.n3489 2.2505
R6701 VSS.n3488 VSS.n3402 2.2505
R6702 VSS.n3487 VSS.n3486 2.2505
R6703 VSS.n3485 VSS.n3403 2.2505
R6704 VSS.n3484 VSS.n3483 2.2505
R6705 VSS.n3482 VSS.n3404 2.2505
R6706 VSS.n3481 VSS.n3480 2.2505
R6707 VSS.n3479 VSS.n3405 2.2505
R6708 VSS.n3478 VSS.n3477 2.2505
R6709 VSS.n3476 VSS.n3406 2.2505
R6710 VSS.n3475 VSS.n3474 2.2505
R6711 VSS.n3473 VSS.n3407 2.2505
R6712 VSS.n3472 VSS.n3471 2.2505
R6713 VSS.n3470 VSS.n3408 2.2505
R6714 VSS.n3469 VSS.n3468 2.2505
R6715 VSS.n3467 VSS.n3409 2.2505
R6716 VSS.n3466 VSS.n3465 2.2505
R6717 VSS.n3464 VSS.n3410 2.2505
R6718 VSS.n3463 VSS.n3462 2.2505
R6719 VSS.n3461 VSS.n3411 2.2505
R6720 VSS.n3460 VSS.n3459 2.2505
R6721 VSS.n3458 VSS.n3412 2.2505
R6722 VSS.n3457 VSS.n3456 2.2505
R6723 VSS.n3455 VSS.n3413 2.2505
R6724 VSS.n3454 VSS.n3453 2.2505
R6725 VSS.n3452 VSS.n3414 2.2505
R6726 VSS.n3451 VSS.n3450 2.2505
R6727 VSS.n3449 VSS.n3415 2.2505
R6728 VSS.n3448 VSS.n3447 2.2505
R6729 VSS.n3446 VSS.n3416 2.2505
R6730 VSS.n3445 VSS.n3444 2.2505
R6731 VSS.n3443 VSS.n3417 2.2505
R6732 VSS.n3442 VSS.n3441 2.2505
R6733 VSS.n3440 VSS.n3418 2.2505
R6734 VSS.n3439 VSS.n3438 2.2505
R6735 VSS.n3437 VSS.n3419 2.2505
R6736 VSS.n3436 VSS.n3435 2.2505
R6737 VSS.n3434 VSS.n3420 2.2505
R6738 VSS.n3433 VSS.n3432 2.2505
R6739 VSS.n3431 VSS.n3421 2.2505
R6740 VSS.n3430 VSS.n3429 2.2505
R6741 VSS.n3428 VSS.n3422 2.2505
R6742 VSS.n3427 VSS.n3426 2.2505
R6743 VSS.n3425 VSS.n3423 2.2505
R6744 VSS.n3424 VSS.n1581 2.2505
R6745 VSS.n8951 VSS.n1582 2.2505
R6746 VSS.n8950 VSS.n8949 2.2505
R6747 VSS.n8948 VSS.n1583 2.2505
R6748 VSS.n8947 VSS.n8946 2.2505
R6749 VSS.n8945 VSS.n1584 2.2505
R6750 VSS.n8944 VSS.n8943 2.2505
R6751 VSS.n8942 VSS.n1585 2.2505
R6752 VSS.n8941 VSS.n8940 2.2505
R6753 VSS.n8939 VSS.n1586 2.2505
R6754 VSS.n8938 VSS.n8937 2.2505
R6755 VSS.n8936 VSS.n1587 2.2505
R6756 VSS.n8935 VSS.n8934 2.2505
R6757 VSS.n8933 VSS.n1588 2.2505
R6758 VSS.n8932 VSS.n8931 2.2505
R6759 VSS.n8930 VSS.n1589 2.2505
R6760 VSS.n8929 VSS.n8928 2.2505
R6761 VSS.n8927 VSS.n1590 2.2505
R6762 VSS.n8926 VSS.n8925 2.2505
R6763 VSS.n8924 VSS.n1591 2.2505
R6764 VSS.n8923 VSS.n8922 2.2505
R6765 VSS.n8921 VSS.n1592 2.2505
R6766 VSS.n8920 VSS.n8919 2.2505
R6767 VSS.n8918 VSS.n1593 2.2505
R6768 VSS.n8917 VSS.n8916 2.2505
R6769 VSS.n8915 VSS.n1594 2.2505
R6770 VSS.n8914 VSS.n8913 2.2505
R6771 VSS.n8912 VSS.n1595 2.2505
R6772 VSS.n8911 VSS.n8910 2.2505
R6773 VSS.n8909 VSS.n1596 2.2505
R6774 VSS.n8908 VSS.n8907 2.2505
R6775 VSS.n8906 VSS.n1597 2.2505
R6776 VSS.n8905 VSS.n8904 2.2505
R6777 VSS.n8903 VSS.n1598 2.2505
R6778 VSS.n8902 VSS.n8901 2.2505
R6779 VSS.n8900 VSS.n1599 2.2505
R6780 VSS.n8899 VSS.n8898 2.2505
R6781 VSS.n8897 VSS.n1600 2.2505
R6782 VSS.n8896 VSS.n8895 2.2505
R6783 VSS.n8894 VSS.n1601 2.2505
R6784 VSS.n8893 VSS.n8892 2.2505
R6785 VSS.n8891 VSS.n1602 2.2505
R6786 VSS.n8890 VSS.n8889 2.2505
R6787 VSS.n8888 VSS.n1603 2.2505
R6788 VSS.n8887 VSS.n8886 2.2505
R6789 VSS.n8885 VSS.n1604 2.2505
R6790 VSS.n8884 VSS.n8883 2.2505
R6791 VSS.n8882 VSS.n1605 2.2505
R6792 VSS.n8881 VSS.n8880 2.2505
R6793 VSS.n8879 VSS.n1606 2.2505
R6794 VSS.n8878 VSS.n8877 2.2505
R6795 VSS.n8876 VSS.n1607 2.2505
R6796 VSS.n8875 VSS.n8874 2.2505
R6797 VSS.n8873 VSS.n1608 2.2505
R6798 VSS.n8872 VSS.n8871 2.2505
R6799 VSS.n8870 VSS.n1609 2.2505
R6800 VSS.n8869 VSS.n8868 2.2505
R6801 VSS.n8867 VSS.n1610 2.2505
R6802 VSS.n8866 VSS.n8865 2.2505
R6803 VSS.n8864 VSS.n1611 2.2505
R6804 VSS.n8863 VSS.n8862 2.2505
R6805 VSS.n8861 VSS.n1612 2.2505
R6806 VSS.n8860 VSS.n8859 2.2505
R6807 VSS.n8858 VSS.n1613 2.2505
R6808 VSS.n8857 VSS.n8856 2.2505
R6809 VSS.n8855 VSS.n1614 2.2505
R6810 VSS.n8854 VSS.n8853 2.2505
R6811 VSS.n8852 VSS.n1615 2.2505
R6812 VSS.n8851 VSS.n8850 2.2505
R6813 VSS.n8849 VSS.n1616 2.2505
R6814 VSS.n8848 VSS.n8847 2.2505
R6815 VSS.n8846 VSS.n1617 2.2505
R6816 VSS.n8845 VSS.n8844 2.2505
R6817 VSS.n8843 VSS.n1618 2.2505
R6818 VSS.n8842 VSS.n8841 2.2505
R6819 VSS.n8840 VSS.n1619 2.2505
R6820 VSS.n8839 VSS.n8838 2.2505
R6821 VSS.n8837 VSS.n1620 2.2505
R6822 VSS.n8836 VSS.n8835 2.2505
R6823 VSS.n8834 VSS.n1621 2.2505
R6824 VSS.n8833 VSS.n8832 2.2505
R6825 VSS.n8831 VSS.n1622 2.2505
R6826 VSS.n8830 VSS.n8829 2.2505
R6827 VSS.n8828 VSS.n1623 2.2505
R6828 VSS.n8827 VSS.n8826 2.2505
R6829 VSS.n8825 VSS.n1624 2.2505
R6830 VSS.n8824 VSS.n8823 2.2505
R6831 VSS.n8822 VSS.n1625 2.2505
R6832 VSS.n8821 VSS.n8820 2.2505
R6833 VSS.n8819 VSS.n1626 2.2505
R6834 VSS.n8818 VSS.n8817 2.2505
R6835 VSS.n8816 VSS.n1627 2.2505
R6836 VSS.n8815 VSS.n8814 2.2505
R6837 VSS.n8813 VSS.n1628 2.2505
R6838 VSS.n8812 VSS.n8811 2.2505
R6839 VSS.n8810 VSS.n1629 2.2505
R6840 VSS.n8809 VSS.n8808 2.2505
R6841 VSS.n8807 VSS.n1630 2.2505
R6842 VSS.n8806 VSS.n8805 2.2505
R6843 VSS.n8804 VSS.n1631 2.2505
R6844 VSS.n8803 VSS.n8802 2.2505
R6845 VSS.n8801 VSS.n1632 2.2505
R6846 VSS.n8800 VSS.n8799 2.2505
R6847 VSS.n8798 VSS.n1633 2.2505
R6848 VSS.n8797 VSS.n8796 2.2505
R6849 VSS.n8795 VSS.n1634 2.2505
R6850 VSS.n8794 VSS.n8793 2.2505
R6851 VSS.n8792 VSS.n1635 2.2505
R6852 VSS.n8791 VSS.n8790 2.2505
R6853 VSS.n8789 VSS.n1636 2.2505
R6854 VSS.n8788 VSS.n8787 2.2505
R6855 VSS.n8786 VSS.n1637 2.2505
R6856 VSS.n8785 VSS.n8784 2.2505
R6857 VSS.n8783 VSS.n1638 2.2505
R6858 VSS.n8782 VSS.n8781 2.2505
R6859 VSS.n8780 VSS.n1639 2.2505
R6860 VSS.n8779 VSS.n8778 2.2505
R6861 VSS.n8777 VSS.n1640 2.2505
R6862 VSS.n8776 VSS.n8775 2.2505
R6863 VSS.n8774 VSS.n1641 2.2505
R6864 VSS.n8773 VSS.n8772 2.2505
R6865 VSS.n8771 VSS.n1642 2.2505
R6866 VSS.n8770 VSS.n8769 2.2505
R6867 VSS.n8768 VSS.n1643 2.2505
R6868 VSS.n8767 VSS.n8766 2.2505
R6869 VSS.n8765 VSS.n1644 2.2505
R6870 VSS.n8764 VSS.n8763 2.2505
R6871 VSS.n8762 VSS.n1645 2.2505
R6872 VSS.n8761 VSS.n8760 2.2505
R6873 VSS.n8759 VSS.n1646 2.2505
R6874 VSS.n8758 VSS.n8757 2.2505
R6875 VSS.n8756 VSS.n1647 2.2505
R6876 VSS.n8755 VSS.n8754 2.2505
R6877 VSS.n8753 VSS.n1648 2.2505
R6878 VSS.n8752 VSS.n8751 2.2505
R6879 VSS.n8750 VSS.n1649 2.2505
R6880 VSS.n8749 VSS.n8748 2.2505
R6881 VSS.n8747 VSS.n1650 2.2505
R6882 VSS.n8746 VSS.n8745 2.2505
R6883 VSS.n8744 VSS.n1651 2.2505
R6884 VSS.n8743 VSS.n8742 2.2505
R6885 VSS.n8741 VSS.n1652 2.2505
R6886 VSS.n8740 VSS.n8739 2.2505
R6887 VSS.n8738 VSS.n1653 2.2505
R6888 VSS.n8737 VSS.n8736 2.2505
R6889 VSS.n8735 VSS.n1654 2.2505
R6890 VSS.n8734 VSS.n8733 2.2505
R6891 VSS.n8732 VSS.n1655 2.2505
R6892 VSS.n8731 VSS.n8730 2.2505
R6893 VSS.n8729 VSS.n1656 2.2505
R6894 VSS.n8728 VSS.n8727 2.2505
R6895 VSS.n8726 VSS.n1657 2.2505
R6896 VSS.n8725 VSS.n8724 2.2505
R6897 VSS.n8723 VSS.n1658 2.2505
R6898 VSS.n8722 VSS.n8721 2.2505
R6899 VSS.n8720 VSS.n1659 2.2505
R6900 VSS.n8719 VSS.n8718 2.2505
R6901 VSS.n8717 VSS.n1660 2.2505
R6902 VSS.n8716 VSS.n8715 2.2505
R6903 VSS.n8714 VSS.n1661 2.2505
R6904 VSS.n8713 VSS.n8712 2.2505
R6905 VSS.n8711 VSS.n1662 2.2505
R6906 VSS.n8710 VSS.n8709 2.2505
R6907 VSS.n8708 VSS.n1663 2.2505
R6908 VSS.n8707 VSS.n8706 2.2505
R6909 VSS.n8705 VSS.n1664 2.2505
R6910 VSS.n8704 VSS.n8703 2.2505
R6911 VSS.n8702 VSS.n1665 2.2505
R6912 VSS.n8701 VSS.n8700 2.2505
R6913 VSS.n8699 VSS.n1666 2.2505
R6914 VSS.n8698 VSS.n8697 2.2505
R6915 VSS.n8696 VSS.n1667 2.2505
R6916 VSS.n8695 VSS.n8694 2.2505
R6917 VSS.n8693 VSS.n1668 2.2505
R6918 VSS.n8692 VSS.n8691 2.2505
R6919 VSS.n8690 VSS.n1669 2.2505
R6920 VSS.n8689 VSS.n8688 2.2505
R6921 VSS.n8687 VSS.n1670 2.2505
R6922 VSS.n8686 VSS.n8685 2.2505
R6923 VSS.n8684 VSS.n1671 2.2505
R6924 VSS.n8683 VSS.n8682 2.2505
R6925 VSS.n8681 VSS.n1672 2.2505
R6926 VSS.n8680 VSS.n8679 2.2505
R6927 VSS.n8678 VSS.n1673 2.2505
R6928 VSS.n8677 VSS.n8676 2.2505
R6929 VSS.n8675 VSS.n1674 2.2505
R6930 VSS.n8674 VSS.n8673 2.2505
R6931 VSS.n8672 VSS.n1675 2.2505
R6932 VSS.n8671 VSS.n8670 2.2505
R6933 VSS.n8669 VSS.n1676 2.2505
R6934 VSS.n8668 VSS.n8667 2.2505
R6935 VSS.n8666 VSS.n1677 2.2505
R6936 VSS.n8665 VSS.n8664 2.2505
R6937 VSS.n8663 VSS.n1678 2.2505
R6938 VSS.n8662 VSS.n8661 2.2505
R6939 VSS.n8660 VSS.n1679 2.2505
R6940 VSS.n8659 VSS.n8658 2.2505
R6941 VSS.n8657 VSS.n1680 2.2505
R6942 VSS.n8656 VSS.n8655 2.2505
R6943 VSS.n8654 VSS.n1681 2.2505
R6944 VSS.n8653 VSS.n8652 2.2505
R6945 VSS.n8651 VSS.n1682 2.2505
R6946 VSS.n8650 VSS.n8649 2.2505
R6947 VSS.n8648 VSS.n1683 2.2505
R6948 VSS.n8647 VSS.n8646 2.2505
R6949 VSS.n8645 VSS.n1684 2.2505
R6950 VSS.n8644 VSS.n8643 2.2505
R6951 VSS.n8642 VSS.n1685 2.2505
R6952 VSS.n8641 VSS.n8640 2.2505
R6953 VSS.n8639 VSS.n1686 2.2505
R6954 VSS.n8638 VSS.n8637 2.2505
R6955 VSS.n8636 VSS.n1687 2.2505
R6956 VSS.n8635 VSS.n8634 2.2505
R6957 VSS.n8633 VSS.n1688 2.2505
R6958 VSS.n8632 VSS.n8631 2.2505
R6959 VSS.n8630 VSS.n1689 2.2505
R6960 VSS.n8629 VSS.n8628 2.2505
R6961 VSS.n8627 VSS.n1690 2.2505
R6962 VSS.n8626 VSS.n8625 2.2505
R6963 VSS.n8624 VSS.n1691 2.2505
R6964 VSS.n8623 VSS.n8622 2.2505
R6965 VSS.n8621 VSS.n1692 2.2505
R6966 VSS.n8620 VSS.n8619 2.2505
R6967 VSS.n8618 VSS.n1693 2.2505
R6968 VSS.n8617 VSS.n8616 2.2505
R6969 VSS.n8615 VSS.n1694 2.2505
R6970 VSS.n8614 VSS.n8613 2.2505
R6971 VSS.n8612 VSS.n1695 2.2505
R6972 VSS.n8611 VSS.n8610 2.2505
R6973 VSS.n8609 VSS.n1696 2.2505
R6974 VSS.n8608 VSS.n8607 2.2505
R6975 VSS.n8606 VSS.n1697 2.2505
R6976 VSS.n8605 VSS.n8604 2.2505
R6977 VSS.n8603 VSS.n1698 2.2505
R6978 VSS.n8602 VSS.n8601 2.2505
R6979 VSS.n8600 VSS.n1699 2.2505
R6980 VSS.n8599 VSS.n8598 2.2505
R6981 VSS.n8597 VSS.n1700 2.2505
R6982 VSS.n8596 VSS.n8595 2.2505
R6983 VSS.n8594 VSS.n1701 2.2505
R6984 VSS.n8593 VSS.n8592 2.2505
R6985 VSS.n8591 VSS.n1702 2.2505
R6986 VSS.n8590 VSS.n8589 2.2505
R6987 VSS.n8588 VSS.n1703 2.2505
R6988 VSS.n8587 VSS.n8586 2.2505
R6989 VSS.n8585 VSS.n1704 2.2505
R6990 VSS.n8584 VSS.n8583 2.2505
R6991 VSS.n8582 VSS.n1705 2.2505
R6992 VSS.n8581 VSS.n8580 2.2505
R6993 VSS.n8579 VSS.n1706 2.2505
R6994 VSS.n8578 VSS.n8577 2.2505
R6995 VSS.n8576 VSS.n1707 2.2505
R6996 VSS.n8575 VSS.n8574 2.2505
R6997 VSS.n8573 VSS.n1708 2.2505
R6998 VSS.n8572 VSS.n8571 2.2505
R6999 VSS.n8570 VSS.n1709 2.2505
R7000 VSS.n8569 VSS.n8568 2.2505
R7001 VSS.n8567 VSS.n1710 2.2505
R7002 VSS.n8566 VSS.n8565 2.2505
R7003 VSS.n8564 VSS.n1711 2.2505
R7004 VSS.n8563 VSS.n8562 2.2505
R7005 VSS.n8561 VSS.n1712 2.2505
R7006 VSS.n8560 VSS.n8559 2.2505
R7007 VSS.n8558 VSS.n1713 2.2505
R7008 VSS.n8557 VSS.n8556 2.2505
R7009 VSS.n8555 VSS.n1714 2.2505
R7010 VSS.n8554 VSS.n8553 2.2505
R7011 VSS.n8552 VSS.n1715 2.2505
R7012 VSS.n8551 VSS.n8550 2.2505
R7013 VSS.n8549 VSS.n1716 2.2505
R7014 VSS.n8548 VSS.n8547 2.2505
R7015 VSS.n8546 VSS.n1717 2.2505
R7016 VSS.n8545 VSS.n8544 2.2505
R7017 VSS.n8543 VSS.n1718 2.2505
R7018 VSS.n8542 VSS.n8541 2.2505
R7019 VSS.n8540 VSS.n1719 2.2505
R7020 VSS.n8539 VSS.n8538 2.2505
R7021 VSS.n8537 VSS.n1720 2.2505
R7022 VSS.n8536 VSS.n8535 2.2505
R7023 VSS.n8534 VSS.n1721 2.2505
R7024 VSS.n8533 VSS.n8532 2.2505
R7025 VSS.n8531 VSS.n1722 2.2505
R7026 VSS.n8530 VSS.n8529 2.2505
R7027 VSS.n8528 VSS.n1723 2.2505
R7028 VSS.n8527 VSS.n8526 2.2505
R7029 VSS.n8525 VSS.n1724 2.2505
R7030 VSS.n8524 VSS.n8523 2.2505
R7031 VSS.n8522 VSS.n1725 2.2505
R7032 VSS.n8521 VSS.n8520 2.2505
R7033 VSS.n8519 VSS.n1726 2.2505
R7034 VSS.n8518 VSS.n8517 2.2505
R7035 VSS.n8516 VSS.n1727 2.2505
R7036 VSS.n8515 VSS.n8514 2.2505
R7037 VSS.n8513 VSS.n1728 2.2505
R7038 VSS.n8512 VSS.n8511 2.2505
R7039 VSS.n8510 VSS.n1729 2.2505
R7040 VSS.n8509 VSS.n8508 2.2505
R7041 VSS.n8507 VSS.n1730 2.2505
R7042 VSS.n8506 VSS.n8505 2.2505
R7043 VSS.n8504 VSS.n1731 2.2505
R7044 VSS.n8503 VSS.n8502 2.2505
R7045 VSS.n8501 VSS.n1732 2.2505
R7046 VSS.n8500 VSS.n8499 2.2505
R7047 VSS.n8498 VSS.n1733 2.2505
R7048 VSS.n8497 VSS.n8496 2.2505
R7049 VSS.n8495 VSS.n1734 2.2505
R7050 VSS.n8494 VSS.n8493 2.2505
R7051 VSS.n8492 VSS.n1735 2.2505
R7052 VSS.n8491 VSS.n8490 2.2505
R7053 VSS.n8489 VSS.n1736 2.2505
R7054 VSS.n8488 VSS.n8487 2.2505
R7055 VSS.n8486 VSS.n1737 2.2505
R7056 VSS.n8485 VSS.n8484 2.2505
R7057 VSS.n8483 VSS.n1738 2.2505
R7058 VSS.n8482 VSS.n8481 2.2505
R7059 VSS.n8480 VSS.n1739 2.2505
R7060 VSS.n8479 VSS.n8478 2.2505
R7061 VSS.n8477 VSS.n1740 2.2505
R7062 VSS.n8476 VSS.n8475 2.2505
R7063 VSS.n8474 VSS.n1741 2.2505
R7064 VSS.n8473 VSS.n8472 2.2505
R7065 VSS.n8471 VSS.n1742 2.2505
R7066 VSS.n8470 VSS.n8469 2.2505
R7067 VSS.n8468 VSS.n1743 2.2505
R7068 VSS.n8467 VSS.n8466 2.2505
R7069 VSS.n8465 VSS.n1744 2.2505
R7070 VSS.n8464 VSS.n8463 2.2505
R7071 VSS.n8462 VSS.n1745 2.2505
R7072 VSS.n8461 VSS.n8460 2.2505
R7073 VSS.n8459 VSS.n1746 2.2505
R7074 VSS.n8458 VSS.n8457 2.2505
R7075 VSS.n8456 VSS.n1747 2.2505
R7076 VSS.n8455 VSS.n8454 2.2505
R7077 VSS.n8453 VSS.n1748 2.2505
R7078 VSS.n8452 VSS.n8451 2.2505
R7079 VSS.n8450 VSS.n1749 2.2505
R7080 VSS.n8449 VSS.n8448 2.2505
R7081 VSS.n8447 VSS.n1750 2.2505
R7082 VSS.n8446 VSS.n8445 2.2505
R7083 VSS.n8444 VSS.n1751 2.2505
R7084 VSS.n8443 VSS.n8442 2.2505
R7085 VSS.n8441 VSS.n1752 2.2505
R7086 VSS.n8440 VSS.n8439 2.2505
R7087 VSS.n8438 VSS.n1753 2.2505
R7088 VSS.n8437 VSS.n8436 2.2505
R7089 VSS.n8435 VSS.n1754 2.2505
R7090 VSS.n8434 VSS.n8433 2.2505
R7091 VSS.n8432 VSS.n1755 2.2505
R7092 VSS.n8431 VSS.n8430 2.2505
R7093 VSS.n8429 VSS.n1756 2.2505
R7094 VSS.n8428 VSS.n8427 2.2505
R7095 VSS.n8426 VSS.n1757 2.2505
R7096 VSS.n8425 VSS.n8424 2.2505
R7097 VSS.n8423 VSS.n1758 2.2505
R7098 VSS.n8422 VSS.n8421 2.2505
R7099 VSS.n8420 VSS.n1759 2.2505
R7100 VSS.n8419 VSS.n8418 2.2505
R7101 VSS.n8417 VSS.n1760 2.2505
R7102 VSS.n8416 VSS.n8415 2.2505
R7103 VSS.n8414 VSS.n1761 2.2505
R7104 VSS.n8413 VSS.n8412 2.2505
R7105 VSS.n8411 VSS.n1762 2.2505
R7106 VSS.n8410 VSS.n8409 2.2505
R7107 VSS.n8408 VSS.n1763 2.2505
R7108 VSS.n8407 VSS.n8406 2.2505
R7109 VSS.n8405 VSS.n1764 2.2505
R7110 VSS.n8404 VSS.n8403 2.2505
R7111 VSS.n8402 VSS.n1765 2.2505
R7112 VSS.n8401 VSS.n8400 2.2505
R7113 VSS.n8399 VSS.n1766 2.2505
R7114 VSS.n8398 VSS.n8397 2.2505
R7115 VSS.n8396 VSS.n1767 2.2505
R7116 VSS.n8395 VSS.n8394 2.2505
R7117 VSS.n8393 VSS.n1768 2.2505
R7118 VSS.n8392 VSS.n8391 2.2505
R7119 VSS.n8390 VSS.n1769 2.2505
R7120 VSS.n8389 VSS.n8388 2.2505
R7121 VSS.n8387 VSS.n1770 2.2505
R7122 VSS.n8386 VSS.n8385 2.2505
R7123 VSS.n8384 VSS.n1771 2.2505
R7124 VSS.n8383 VSS.n8382 2.2505
R7125 VSS.n8381 VSS.n1772 2.2505
R7126 VSS.n8380 VSS.n8379 2.2505
R7127 VSS.n8378 VSS.n1773 2.2505
R7128 VSS.n8377 VSS.n8376 2.2505
R7129 VSS.n8375 VSS.n1774 2.2505
R7130 VSS.n8374 VSS.n8373 2.2505
R7131 VSS.n8372 VSS.n1775 2.2505
R7132 VSS.n8371 VSS.n8370 2.2505
R7133 VSS.n8369 VSS.n1776 2.2505
R7134 VSS.n8368 VSS.n8367 2.2505
R7135 VSS.n8366 VSS.n1777 2.2505
R7136 VSS.n8365 VSS.n8364 2.2505
R7137 VSS.n8363 VSS.n1778 2.2505
R7138 VSS.n8362 VSS.n8361 2.2505
R7139 VSS.n8360 VSS.n1779 2.2505
R7140 VSS.n8359 VSS.n8358 2.2505
R7141 VSS.n8357 VSS.n1780 2.2505
R7142 VSS.n8356 VSS.n8355 2.2505
R7143 VSS.n8354 VSS.n1781 2.2505
R7144 VSS.n8353 VSS.n8352 2.2505
R7145 VSS.n8351 VSS.n1782 2.2505
R7146 VSS.n8350 VSS.n8349 2.2505
R7147 VSS.n8348 VSS.n1783 2.2505
R7148 VSS.n8347 VSS.n8346 2.2505
R7149 VSS.n8345 VSS.n1784 2.2505
R7150 VSS.n8344 VSS.n8343 2.2505
R7151 VSS.n8342 VSS.n1785 2.2505
R7152 VSS.n8341 VSS.n8340 2.2505
R7153 VSS.n8339 VSS.n1786 2.2505
R7154 VSS.n8338 VSS.n8337 2.2505
R7155 VSS.n8336 VSS.n1787 2.2505
R7156 VSS.n8335 VSS.n8334 2.2505
R7157 VSS.n8333 VSS.n1788 2.2505
R7158 VSS.n8332 VSS.n8331 2.2505
R7159 VSS.n8330 VSS.n1789 2.2505
R7160 VSS.n8329 VSS.n8328 2.2505
R7161 VSS.n8327 VSS.n1790 2.2505
R7162 VSS.n8326 VSS.n8325 2.2505
R7163 VSS.n8324 VSS.n1791 2.2505
R7164 VSS.n8323 VSS.n8322 2.2505
R7165 VSS.n8321 VSS.n1792 2.2505
R7166 VSS.n8320 VSS.n8319 2.2505
R7167 VSS.n8318 VSS.n1793 2.2505
R7168 VSS.n8317 VSS.n8316 2.2505
R7169 VSS.n8315 VSS.n1794 2.2505
R7170 VSS.n8314 VSS.n8313 2.2505
R7171 VSS.n8312 VSS.n1795 2.2505
R7172 VSS.n8311 VSS.n8310 2.2505
R7173 VSS.n8309 VSS.n1796 2.2505
R7174 VSS.n8308 VSS.n8307 2.2505
R7175 VSS.n8306 VSS.n1797 2.2505
R7176 VSS.n8305 VSS.n8304 2.2505
R7177 VSS.n8303 VSS.n1798 2.2505
R7178 VSS.n8302 VSS.n8301 2.2505
R7179 VSS.n8300 VSS.n1799 2.2505
R7180 VSS.n8299 VSS.n8298 2.2505
R7181 VSS.n8297 VSS.n1800 2.2505
R7182 VSS.n8296 VSS.n8295 2.2505
R7183 VSS.n8294 VSS.n1801 2.2505
R7184 VSS.n8293 VSS.n8292 2.2505
R7185 VSS.n8291 VSS.n1802 2.2505
R7186 VSS.n8290 VSS.n8289 2.2505
R7187 VSS.n8288 VSS.n1803 2.2505
R7188 VSS.n8287 VSS.n8286 2.2505
R7189 VSS.n8285 VSS.n1804 2.2505
R7190 VSS.n8284 VSS.n8283 2.2505
R7191 VSS.n8282 VSS.n1805 2.2505
R7192 VSS.n8281 VSS.n8280 2.2505
R7193 VSS.n8279 VSS.n1806 2.2505
R7194 VSS.n8278 VSS.n8277 2.2505
R7195 VSS.n8276 VSS.n1807 2.2505
R7196 VSS.n8275 VSS.n8274 2.2505
R7197 VSS.n8273 VSS.n1808 2.2505
R7198 VSS.n8272 VSS.n8271 2.2505
R7199 VSS.n8270 VSS.n1809 2.2505
R7200 VSS.n8269 VSS.n8268 2.2505
R7201 VSS.n8267 VSS.n1810 2.2505
R7202 VSS.n8266 VSS.n8265 2.2505
R7203 VSS.n8264 VSS.n1811 2.2505
R7204 VSS.n8263 VSS.n8262 2.2505
R7205 VSS.n8261 VSS.n1812 2.2505
R7206 VSS.n8260 VSS.n8259 2.2505
R7207 VSS.n8258 VSS.n1813 2.2505
R7208 VSS.n8257 VSS.n8256 2.2505
R7209 VSS.n8255 VSS.n1814 2.2505
R7210 VSS.n8254 VSS.n8253 2.2505
R7211 VSS.n8252 VSS.n1815 2.2505
R7212 VSS.n8251 VSS.n8250 2.2505
R7213 VSS.n8249 VSS.n1816 2.2505
R7214 VSS.n8248 VSS.n8247 2.2505
R7215 VSS.n8246 VSS.n1817 2.2505
R7216 VSS.n8245 VSS.n8244 2.2505
R7217 VSS.n8243 VSS.n1818 2.2505
R7218 VSS.n8242 VSS.n8241 2.2505
R7219 VSS.n8240 VSS.n1819 2.2505
R7220 VSS.n8239 VSS.n8238 2.2505
R7221 VSS.n8237 VSS.n1820 2.2505
R7222 VSS.n8236 VSS.n8235 2.2505
R7223 VSS.n8234 VSS.n1821 2.2505
R7224 VSS.n8233 VSS.n8232 2.2505
R7225 VSS.n36 VSS.n35 2.25016
R7226 VSS.n58 VSS.n54 2.25016
R7227 VSS.n11395 VSS.n11394 2.25016
R7228 VSS.n11312 VSS.n123 2.2497
R7229 VSS.n10705 VSS.n10703 2.24949
R7230 VSS.n111 VSS.n105 2.24922
R7231 VSS.n10567 VSS.n10566 2.24813
R7232 VSS.n10570 VSS.n10568 2.24218
R7233 VSS.n10572 VSS.n10562 2.24218
R7234 VSS.n10564 VSS.n10556 2.24218
R7235 VSS.n227 VSS.n223 2.24218
R7236 VSS.n10910 VSS.n230 2.24218
R7237 VSS.n10911 VSS.n10910 2.24218
R7238 VSS.n107 VSS.n103 2.24218
R7239 VSS.n110 VSS.n103 2.24218
R7240 VSS.n11431 VSS.n37 2.24218
R7241 VSS.n11429 VSS.n33 2.24218
R7242 VSS.n11433 VSS.n29 2.24218
R7243 VSS.n11400 VSS.n55 2.24218
R7244 VSS.n11398 VSS.n11397 2.24218
R7245 VSS.n11385 VSS.n11384 2.24218
R7246 VSS.n11384 VSS.n79 2.24218
R7247 VSS.n82 VSS.n78 2.24218
R7248 VSS.n11311 VSS.n11310 2.24218
R7249 VSS.n11310 VSS.n126 2.24218
R7250 VSS.n11306 VSS.n11305 2.24218
R7251 VSS.n10732 VSS.n10700 2.24218
R7252 VSS.n10732 VSS.n10699 2.24218
R7253 VSS.n10728 VSS.n10702 2.24218
R7254 VSS.n10334 VSS.n10309 2.23722
R7255 VSS.n10804 VSS.n10803 2.15932
R7256 VSS.n10798 VSS.n10797 2.15932
R7257 VSS.n10806 VSS.n10805 2.15458
R7258 VSS.n10800 VSS.n10799 2.15458
R7259 VSS.n10411 VSS.n10398 2.13932
R7260 VSS.n10767 VSS.t665 2.1005
R7261 VSS.t569 VSS.n10767 2.1005
R7262 VSS.n10756 VSS.t795 2.1005
R7263 VSS.n10756 VSS.t724 2.1005
R7264 VSS.n10474 VSS.n10473 2.1005
R7265 VSS.n10471 VSS.n10470 2.1005
R7266 VSS.n10467 VSS.n10466 2.1005
R7267 VSS.n10463 VSS.n10462 2.1005
R7268 VSS.n10459 VSS.n10458 2.1005
R7269 VSS.n10456 VSS.n10455 2.1005
R7270 VSS.n9072 VSS.n9071 2.1005
R7271 VSS.n9066 VSS.n9065 2.1005
R7272 VSS.n9043 VSS.n9042 2.1005
R7273 VSS.n9087 VSS.n9086 2.1005
R7274 VSS.n8978 VSS.n8977 2.1005
R7275 VSS.n9098 VSS.n9097 2.1005
R7276 VSS.n8968 VSS.n8967 2.1005
R7277 VSS.n9006 VSS.n9005 2.1005
R7278 VSS.n1569 VSS.n1568 2.1005
R7279 VSS.n9037 VSS.n9036 2.1005
R7280 VSS.n841 VSS.n840 2.1005
R7281 VSS.n10925 VSS.n10924 2.1005
R7282 VSS.n876 VSS.n875 2.1005
R7283 VSS.n865 VSS.n864 2.1005
R7284 VSS.n1123 VSS.n1122 2.1005
R7285 VSS.n1129 VSS.n1128 2.1005
R7286 VSS.n1111 VSS.n1110 2.1005
R7287 VSS.n1117 VSS.n1116 2.1005
R7288 VSS.n1090 VSS.n1089 2.1005
R7289 VSS.n1096 VSS.n1095 2.1005
R7290 VSS.n1287 VSS.n1286 2.1005
R7291 VSS.n1293 VSS.n1292 2.1005
R7292 VSS.n10156 VSS.n10155 2.1005
R7293 VSS.n10150 VSS.n10149 2.1005
R7294 VSS.n1074 VSS.n1073 2.1005
R7295 VSS.n1080 VSS.n1079 2.1005
R7296 VSS.n1053 VSS.n1052 2.1005
R7297 VSS.n1059 VSS.n1058 2.1005
R7298 VSS.n389 VSS.n388 2.1005
R7299 VSS.n10162 VSS.n10161 2.1005
R7300 VSS.n368 VSS.n367 2.1005
R7301 VSS.n374 VSS.n373 2.1005
R7302 VSS.n1041 VSS.n1040 2.1005
R7303 VSS.n1047 VSS.n1046 2.1005
R7304 VSS.n1016 VSS.n1015 2.1005
R7305 VSS.n1022 VSS.n1021 2.1005
R7306 VSS.n10216 VSS.n10215 2.1005
R7307 VSS.n10210 VSS.n10209 2.1005
R7308 VSS.n317 VSS.n316 2.1005
R7309 VSS.n10222 VSS.n10221 2.1005
R7310 VSS.n1004 VSS.n1003 2.1005
R7311 VSS.n1010 VSS.n1009 2.1005
R7312 VSS.n983 VSS.n982 2.1005
R7313 VSS.n989 VSS.n988 2.1005
R7314 VSS.n305 VSS.n304 2.1005
R7315 VSS.n311 VSS.n310 2.1005
R7316 VSS.n10276 VSS.n10275 2.1005
R7317 VSS.n10270 VSS.n10269 2.1005
R7318 VSS.n967 VSS.n966 2.1005
R7319 VSS.n973 VSS.n972 2.1005
R7320 VSS.n10577 VSS.n10576 2.1005
R7321 VSS.n10580 VSS.n10579 2.1005
R7322 VSS.n10584 VSS.n10583 2.1005
R7323 VSS.n10675 VSS.n10674 2.1005
R7324 VSS.n10672 VSS.n10671 2.1005
R7325 VSS.n10668 VSS.n10667 2.1005
R7326 VSS.n10356 VSS.n10339 2.1005
R7327 VSS.n10360 VSS.n10359 2.1005
R7328 VSS.n10363 VSS.n10362 2.1005
R7329 VSS.n10419 VSS.n10418 2.1005
R7330 VSS.n10422 VSS.n10421 2.1005
R7331 VSS.n10426 VSS.n10425 2.1005
R7332 VSS.n10430 VSS.n10429 2.1005
R7333 VSS.n10434 VSS.n10433 2.1005
R7334 VSS.n10437 VSS.n10436 2.1005
R7335 VSS.n10588 VSS.n10587 2.1005
R7336 VSS.n10550 VSS.n10549 2.1005
R7337 VSS.n10541 VSS.n10488 2.1005
R7338 VSS.n10523 VSS.n10522 2.1005
R7339 VSS.n10514 VSS.n10509 2.1005
R7340 VSS.n10654 VSS.n10653 2.1005
R7341 VSS.n10548 VSS.n10547 2.1005
R7342 VSS.n10546 VSS.n10545 2.1005
R7343 VSS.n10501 VSS.n10492 2.1005
R7344 VSS.n10527 VSS.n10526 2.1005
R7345 VSS.n10521 VSS.n10520 2.1005
R7346 VSS.n10519 VSS.n10518 2.1005
R7347 VSS.n10652 VSS.n10651 2.1005
R7348 VSS.n10647 VSS.n10646 2.1005
R7349 VSS.n10644 VSS.n10643 2.1005
R7350 VSS.n10919 VSS.n10918 2.1005
R7351 VSS.n10988 VSS.n10987 2.1005
R7352 VSS.n10997 VSS.n10996 2.1005
R7353 VSS.n11357 VSS.n11356 2.1005
R7354 VSS.n11351 VSS.n11350 2.1005
R7355 VSS.n11344 VSS.n11343 2.1005
R7356 VSS.n9451 VSS.n9450 2.1005
R7357 VSS.n9457 VSS.n9456 2.1005
R7358 VSS.n9432 VSS.n9431 2.1005
R7359 VSS.n9472 VSS.n9471 2.1005
R7360 VSS.n819 VSS.n818 2.1005
R7361 VSS.n675 VSS.n674 2.1005
R7362 VSS.n9856 VSS.n9855 2.1005
R7363 VSS.n9876 VSS.n9875 2.1005
R7364 VSS.n11415 VSS.n11414 2.1005
R7365 VSS.n11448 VSS.n11447 2.1005
R7366 VSS.n9515 VSS.n9514 2.1005
R7367 VSS.n1251 VSS.n1250 2.1005
R7368 VSS.n9899 VSS.n9898 2.1005
R7369 VSS.n9912 VSS.n9911 2.1005
R7370 VSS.n9922 VSS.n9921 2.1005
R7371 VSS.n1372 VSS.n1347 2.1005
R7372 VSS.n1366 VSS.n1350 2.1005
R7373 VSS.n1360 VSS.n1352 2.1005
R7374 VSS.n9631 VSS.n9630 2.1005
R7375 VSS.n9763 VSS.n799 2.1005
R7376 VSS.n9757 VSS.n9637 2.1005
R7377 VSS.n9747 VSS.n9664 2.1005
R7378 VSS.n9741 VSS.n9667 2.1005
R7379 VSS.n9735 VSS.n9669 2.1005
R7380 VSS.n9725 VSS.n9720 2.1005
R7381 VSS.n10029 VSS.n570 2.1005
R7382 VSS.n10022 VSS.n575 2.1005
R7383 VSS.n10010 VSS.n9937 2.1005
R7384 VSS.n10004 VSS.n9939 2.1005
R7385 VSS.n9998 VSS.n9941 2.1005
R7386 VSS.n9988 VSS.n9969 2.1005
R7387 VSS.n9982 VSS.n9971 2.1005
R7388 VSS.n9976 VSS.n9973 2.1005
R7389 VSS.n1373 VSS.n1372 2.1005
R7390 VSS.n1367 VSS.n1366 2.1005
R7391 VSS.n1361 VSS.n1360 2.1005
R7392 VSS.n9632 VSS.n9631 2.1005
R7393 VSS.n9763 VSS.n9762 2.1005
R7394 VSS.n9758 VSS.n9757 2.1005
R7395 VSS.n9748 VSS.n9747 2.1005
R7396 VSS.n9742 VSS.n9741 2.1005
R7397 VSS.n9736 VSS.n9735 2.1005
R7398 VSS.n9726 VSS.n9725 2.1005
R7399 VSS.n10029 VSS.n10028 2.1005
R7400 VSS.n10023 VSS.n10022 2.1005
R7401 VSS.n10011 VSS.n10010 2.1005
R7402 VSS.n10005 VSS.n10004 2.1005
R7403 VSS.n9999 VSS.n9998 2.1005
R7404 VSS.n9989 VSS.n9988 2.1005
R7405 VSS.n9983 VSS.n9982 2.1005
R7406 VSS.n9977 VSS.n9976 2.1005
R7407 VSS.n9614 VSS.n9613 2.1005
R7408 VSS.n1310 VSS.n1309 2.1005
R7409 VSS.n10114 VSS.n10113 2.1005
R7410 VSS.n10109 VSS.n10108 2.1005
R7411 VSS.n10094 VSS.n10093 2.1005
R7412 VSS.n10088 VSS.n10087 2.1005
R7413 VSS.n10082 VSS.n10081 2.1005
R7414 VSS.n525 VSS.n524 2.1005
R7415 VSS.n10063 VSS.n10062 2.1005
R7416 VSS.n10056 VSS.n10055 2.1005
R7417 VSS.n10041 VSS.n10040 2.1005
R7418 VSS.n10871 VSS.n235 2.1005
R7419 VSS.n10888 VSS.n10887 2.1005
R7420 VSS.n11133 VSS.n202 2.1005
R7421 VSS.n11130 VSS.n11129 2.1005
R7422 VSS.n11124 VSS.n11123 2.1005
R7423 VSS.n11109 VSS.n11108 2.1005
R7424 VSS.n11103 VSS.n11102 2.1005
R7425 VSS.n11097 VSS.n11096 2.1005
R7426 VSS.n1315 VSS.n1314 2.1005
R7427 VSS.n1306 VSS.n1305 2.1005
R7428 VSS.n445 VSS.n444 2.1005
R7429 VSS.n10106 VSS.n10105 2.1005
R7430 VSS.n10101 VSS.n10100 2.1005
R7431 VSS.n10092 VSS.n10091 2.1005
R7432 VSS.n10086 VSS.n10085 2.1005
R7433 VSS.n10078 VSS.n10077 2.1005
R7434 VSS.n10073 VSS.n10072 2.1005
R7435 VSS.n521 VSS.n520 2.1005
R7436 VSS.n532 VSS.n513 2.1005
R7437 VSS.n10058 VSS.n10057 2.1005
R7438 VSS.n10052 VSS.n10051 2.1005
R7439 VSS.n10044 VSS.n10043 2.1005
R7440 VSS.n10037 VSS.n10036 2.1005
R7441 VSS.n10892 VSS.n10891 2.1005
R7442 VSS.n10881 VSS.n10878 2.1005
R7443 VSS.n11148 VSS.n11147 2.1005
R7444 VSS.n11136 VSS.n11135 2.1005
R7445 VSS.n11127 VSS.n11126 2.1005
R7446 VSS.n11121 VSS.n11120 2.1005
R7447 VSS.n11116 VSS.n11115 2.1005
R7448 VSS.n11107 VSS.n11106 2.1005
R7449 VSS.n11101 VSS.n11100 2.1005
R7450 VSS.n11095 VSS.n11094 2.1005
R7451 VSS.n11464 VSS.n11463 2.1005
R7452 VSS.n11323 VSS.n11322 2.1005
R7453 VSS.n11373 VSS.n11372 2.1005
R7454 VSS.n11380 VSS.n11379 2.1005
R7455 VSS.n10951 VSS.n10950 2.1005
R7456 VSS.n11367 VSS.n11366 2.1005
R7457 VSS.n10941 VSS.n10940 2.1005
R7458 VSS.n10978 VSS.n10977 2.1005
R7459 VSS.n1167 VSS.n1166 2.1005
R7460 VSS.n10935 VSS.n10934 2.1005
R7461 VSS.n1213 VSS.n1212 2.1005
R7462 VSS.n1203 VSS.n1202 2.1005
R7463 VSS.n9539 VSS.n9538 2.1005
R7464 VSS.n9546 VSS.n9545 2.1005
R7465 VSS.n1474 VSS.n1473 2.1005
R7466 VSS.n1465 VSS.n1464 2.1005
R7467 VSS.n1460 VSS.n1459 2.1005
R7468 VSS.n1448 VSS.n1447 2.1005
R7469 VSS.n9596 VSS.n828 2.1005
R7470 VSS.n9592 VSS.n9591 2.1005
R7471 VSS.n9778 VSS.n9777 2.1005
R7472 VSS.n9789 VSS.n9788 2.1005
R7473 VSS.n9795 VSS.n9794 2.1005
R7474 VSS.n9805 VSS.n9804 2.1005
R7475 VSS.n9815 VSS.n9814 2.1005
R7476 VSS.n9828 VSS.n9827 2.1005
R7477 VSS.n9839 VSS.n9838 2.1005
R7478 VSS.n760 VSS.n759 2.1005
R7479 VSS.n753 VSS.n752 2.1005
R7480 VSS.n741 VSS.n727 2.1005
R7481 VSS.n738 VSS.n737 2.1005
R7482 VSS.n11160 VSS.n11159 2.1005
R7483 VSS.n11169 VSS.n11168 2.1005
R7484 VSS.n11273 VSS.n11272 2.1005
R7485 VSS.n11267 VSS.n11266 2.1005
R7486 VSS.n11260 VSS.n11259 2.1005
R7487 VSS.n11251 VSS.n11250 2.1005
R7488 VSS.n11245 VSS.n11244 2.1005
R7489 VSS.n11239 VSS.n11238 2.1005
R7490 VSS.n1469 VSS.n1468 2.1005
R7491 VSS.n1457 VSS.n1456 2.1005
R7492 VSS.n1451 VSS.n1450 2.1005
R7493 VSS.n9594 VSS.n9593 2.1005
R7494 VSS.n9773 VSS.n795 2.1005
R7495 VSS.n9786 VSS.n9785 2.1005
R7496 VSS.n9809 VSS.n9808 2.1005
R7497 VSS.n9820 VSS.n9819 2.1005
R7498 VSS.n9832 VSS.n9831 2.1005
R7499 VSS.n757 VSS.n756 2.1005
R7500 VSS.n749 VSS.n748 2.1005
R7501 VSS.n744 VSS.n743 2.1005
R7502 VSS.n11166 VSS.n11165 2.1005
R7503 VSS.n11276 VSS.n11275 2.1005
R7504 VSS.n11270 VSS.n11269 2.1005
R7505 VSS.n11253 VSS.n11252 2.1005
R7506 VSS.n11247 VSS.n11246 2.1005
R7507 VSS.n11241 VSS.n11240 2.1005
R7508 VSS.n1401 VSS.n1400 2.1005
R7509 VSS.n9533 VSS.n9532 2.1005
R7510 VSS.n1493 VSS.n1492 2.1005
R7511 VSS.n9418 VSS.n9417 2.1005
R7512 VSS.n9379 VSS.n9378 2.1005
R7513 VSS.n9386 VSS.n9385 2.1005
R7514 VSS.n9319 VSS.n9318 2.1005
R7515 VSS.n9342 VSS.n9341 2.1005
R7516 VSS.n9267 VSS.n9266 2.1005
R7517 VSS.n9353 VSS.n9352 2.1005
R7518 VSS.n9261 VSS.n9260 2.1005
R7519 VSS.n9295 VSS.n9294 2.1005
R7520 VSS.n9216 VSS.n9215 2.1005
R7521 VSS.n9313 VSS.n9312 2.1005
R7522 VSS.n9210 VSS.n9209 2.1005
R7523 VSS.n9244 VSS.n9243 2.1005
R7524 VSS.n9145 VSS.n9144 2.1005
R7525 VSS.n9255 VSS.n9254 2.1005
R7526 VSS.n9135 VSS.n9134 2.1005
R7527 VSS.n9173 VSS.n9172 2.1005
R7528 VSS.n1551 VSS.n1550 2.1005
R7529 VSS.n1545 VSS.n1544 2.1005
R7530 VSS.n9060 VSS.n9059 2.1005
R7531 VSS.n9204 VSS.n9203 2.1005
R7532 VSS.n11392 VSS.n59 2.08328
R7533 VSS.n11390 VSS.n61 2.08259
R7534 VSS.t676 VSS.t249 2.07259
R7535 VSS.t483 VSS.t255 2.07259
R7536 VSS.n10499 VSS.n128 1.97855
R7537 VSS.n8953 VSS.n8952 1.87288
R7538 VSS.n8953 VSS.n253 1.8724
R7539 VSS.n11318 VSS.n11317 1.8392
R7540 VSS.n10633 VSS.n10632 1.7274
R7541 VSS.n9198 VSS.n9197 1.69669
R7542 VSS.n9334 VSS.n9333 1.69669
R7543 VSS.n172 VSS.n171 1.69669
R7544 VSS.n9580 VSS.n9579 1.69669
R7545 VSS.n200 VSS.n199 1.69669
R7546 VSS.n481 VSS.n477 1.69669
R7547 VSS.n9031 VSS.n9030 1.69669
R7548 VSS.n271 VSS.n270 1.69669
R7549 VSS.n343 VSS.n342 1.69669
R7550 VSS.n415 VSS.n414 1.69669
R7551 VSS.n10735 VSS.t3572 1.6805
R7552 VSS.n10790 VSS.t823 1.6805
R7553 VSS.n10792 VSS.t2471 1.6805
R7554 VSS.n10811 VSS.t1197 1.6805
R7555 VSS.n10820 VSS.t3018 1.6805
R7556 VSS.n10701 VSS.t1762 1.6805
R7557 VSS.n10708 VSS.t3530 1.6805
R7558 VSS.n10709 VSS.t769 1.6805
R7559 VSS.n10710 VSS.t2439 1.6805
R7560 VSS.n10711 VSS.t1136 1.6805
R7561 VSS.n10712 VSS.t2964 1.6805
R7562 VSS.n10713 VSS.t1680 1.6805
R7563 VSS.n127 VSS.t3424 1.6805
R7564 VSS.n14 VSS.t3240 1.6805
R7565 VSS.n15 VSS.t2457 1.6805
R7566 VSS.n16 VSS.t2596 1.6805
R7567 VSS.n17 VSS.t1834 1.6805
R7568 VSS.n11294 VSS.t999 1.6805
R7569 VSS.n24 VSS.t1158 1.6805
R7570 VSS.n25 VSS.t3442 1.6805
R7571 VSS.n26 VSS.t2700 1.6805
R7572 VSS.n27 VSS.t2992 1.6805
R7573 VSS.n28 VSS.t920 1.6805
R7574 VSS.n38 VSS.t1546 1.6805
R7575 VSS.n39 VSS.t2526 1.6805
R7576 VSS.n40 VSS.t1770 1.6805
R7577 VSS.n41 VSS.t928 1.6805
R7578 VSS.n42 VSS.t1078 1.6805
R7579 VSS.n133 VSS.t3362 1.6805
R7580 VSS.n49 VSS.t2772 1.6805
R7581 VSS.n50 VSS.t1986 1.6805
R7582 VSS.n51 VSS.t1406 1.6805
R7583 VSS.n52 VSS.t487 1.6805
R7584 VSS.n53 VSS.t1696 1.6805
R7585 VSS.n10641 VSS.t2405 1.6805
R7586 VSS.n10639 VSS.t3638 1.6805
R7587 VSS.n10497 VSS.t3126 1.6805
R7588 VSS.n10494 VSS.t787 1.6805
R7589 VSS.n10605 VSS.t515 1.6805
R7590 VSS.n10608 VSS.t2994 1.6805
R7591 VSS.n10440 VSS.t1477 1.6805
R7592 VSS.n10497 VSS.t1968 1.6805
R7593 VSS.n10494 VSS.t2758 1.6805
R7594 VSS.n10605 VSS.t2540 1.6805
R7595 VSS.n10608 VSS.t1840 1.6805
R7596 VSS.n10440 VSS.t3352 1.6805
R7597 VSS.n10476 VSS.t3250 1.6805
R7598 VSS.n10478 VSS.t3082 1.6805
R7599 VSS.n10481 VSS.t1702 1.6805
R7600 VSS.n10596 VSS.t2912 1.6805
R7601 VSS.n10593 VSS.t1622 1.6805
R7602 VSS.n10453 VSS.t1026 1.6805
R7603 VSS.n10451 VSS.t809 1.6805
R7604 VSS.n10345 VSS.t2546 1.6805
R7605 VSS.n10659 VSS.t628 1.6805
R7606 VSS.n10656 VSS.t2459 1.6805
R7607 VSS.n10573 VSS.t1962 1.6805
R7608 VSS.n10560 VSS.t3180 1.6805
R7609 VSS.n10290 VSS.t856 1.6805
R7610 VSS.n10693 VSS.t602 1.6805
R7611 VSS.n10690 VSS.t3068 1.6805
R7612 VSS.n10688 VSS.t1537 1.6805
R7613 VSS.n1271 VSS.t1994 1.6805
R7614 VSS.n1270 VSS.t1195 1.6805
R7615 VSS.n1269 VSS.t1354 1.6805
R7616 VSS.n1268 VSS.t3634 1.6805
R7617 VSS.n1331 VSS.t2866 1.6805
R7618 VSS.n1334 VSS.t2059 1.6805
R7619 VSS.n1335 VSS.t2209 1.6805
R7620 VSS.n1339 VSS.t1446 1.6805
R7621 VSS.n1342 VSS.t751 1.6805
R7622 VSS.n9494 VSS.t1803 1.6805
R7623 VSS.n9490 VSS.t2193 1.6805
R7624 VSS.n9487 VSS.t3238 1.6805
R7625 VSS.n9506 VSS.t1700 1.6805
R7626 VSS.n9503 VSS.t2558 1.6805
R7627 VSS.n9500 VSS.t1746 1.6805
R7628 VSS.n1345 VSS.t490 1.6805
R7629 VSS.n1375 VSS.t3006 1.6805
R7630 VSS.n9474 VSS.t1556 1.6805
R7631 VSS.n9446 VSS.t2101 1.6805
R7632 VSS.n9424 VSS.t3004 1.6805
R7633 VSS.n9425 VSS.t2159 1.6805
R7634 VSS.n9426 VSS.t3346 1.6805
R7635 VSS.n9427 VSS.t2712 1.6805
R7636 VSS.n9428 VSS.t1250 1.6805
R7637 VSS.n806 VSS.t1766 1.6805
R7638 VSS.n807 VSS.t1886 1.6805
R7639 VSS.n808 VSS.t1072 1.6805
R7640 VSS.n809 VSS.t3360 1.6805
R7641 VSS.n1233 VSS.t3526 1.6805
R7642 VSS.n823 VSS.t2908 1.6805
R7643 VSS.n824 VSS.t2117 1.6805
R7644 VSS.n825 VSS.t1527 1.6805
R7645 VSS.n826 VSS.t669 1.6805
R7646 VSS.n806 VSS.t548 1.6805
R7647 VSS.n807 VSS.t729 1.6805
R7648 VSS.n808 VSS.t3090 1.6805
R7649 VSS.n809 VSS.t2271 1.6805
R7650 VSS.n1233 VSS.t2389 1.6805
R7651 VSS.n823 VSS.t1796 1.6805
R7652 VSS.n824 VSS.t969 1.6805
R7653 VSS.n825 VSS.t3446 1.6805
R7654 VSS.n826 VSS.t2706 1.6805
R7655 VSS.n9639 VSS.t1744 1.6805
R7656 VSS.n9640 VSS.t1870 1.6805
R7657 VSS.n9641 VSS.t1055 1.6805
R7658 VSS.n9642 VSS.t3338 1.6805
R7659 VSS.n647 VSS.t3502 1.6805
R7660 VSS.n777 VSS.t2896 1.6805
R7661 VSS.n776 VSS.t2093 1.6805
R7662 VSS.n775 VSS.t1515 1.6805
R7663 VSS.n774 VSS.t641 1.6805
R7664 VSS.n9639 VSS.t517 1.6805
R7665 VSS.n9640 VSS.t707 1.6805
R7666 VSS.n9641 VSS.t3064 1.6805
R7667 VSS.n9642 VSS.t2261 1.6805
R7668 VSS.n647 VSS.t2375 1.6805
R7669 VSS.n777 VSS.t1782 1.6805
R7670 VSS.n776 VSS.t940 1.6805
R7671 VSS.n775 VSS.t3422 1.6805
R7672 VSS.n774 VSS.t2668 1.6805
R7673 VSS.n9672 VSS.t1918 1.6805
R7674 VSS.n9675 VSS.t1099 1.6805
R7675 VSS.n9678 VSS.t3382 1.6805
R7676 VSS.n9681 VSS.t3552 1.6805
R7677 VSS.n1175 VSS.t2786 1.6805
R7678 VSS.n681 VSS.t2151 1.6805
R7679 VSS.n684 VSS.t1379 1.6805
R7680 VSS.n687 VSS.t719 1.6805
R7681 VSS.n690 VSS.t3084 1.6805
R7682 VSS.n9673 VSS.t829 1.6805
R7683 VSS.n9676 VSS.t971 1.6805
R7684 VSS.n9679 VSS.t3284 1.6805
R7685 VSS.n9682 VSS.t2496 1.6805
R7686 VSS.n1174 VSS.t2642 1.6805
R7687 VSS.n682 VSS.t2010 1.6805
R7688 VSS.n685 VSS.t1247 1.6805
R7689 VSS.n688 VSS.t546 1.6805
R7690 VSS.n691 VSS.t2946 1.6805
R7691 VSS.n660 VSS.t3474 1.6805
R7692 VSS.n659 VSS.t2718 1.6805
R7693 VSS.n658 VSS.t1934 1.6805
R7694 VSS.n657 VSS.t2049 1.6805
R7695 VSS.n672 VSS.t1274 1.6805
R7696 VSS.n9860 VSS.t567 1.6805
R7697 VSS.n9861 VSS.t2954 1.6805
R7698 VSS.n9862 VSS.t2321 1.6805
R7699 VSS.n9863 VSS.t1564 1.6805
R7700 VSS.n660 VSS.t2355 1.6805
R7701 VSS.n659 VSS.t1605 1.6805
R7702 VSS.n658 VSS.t758 1.6805
R7703 VSS.n657 VSS.t899 1.6805
R7704 VSS.n672 VSS.t3224 1.6805
R7705 VSS.n9860 VSS.t2594 1.6805
R7706 VSS.n9861 VSS.t1832 1.6805
R7707 VSS.n9862 VSS.t1211 1.6805
R7708 VSS.n9863 VSS.t3504 1.6805
R7709 VSS.n9955 VSS.t2415 1.6805
R7710 VSS.n9956 VSS.t1658 1.6805
R7711 VSS.n9957 VSS.t825 1.6805
R7712 VSS.n9958 VSS.t959 1.6805
R7713 VSS.n142 VSS.t3274 1.6805
R7714 VSS.n11186 VSS.t2658 1.6805
R7715 VSS.n11185 VSS.t1882 1.6805
R7716 VSS.n11184 VSS.t1272 1.6805
R7717 VSS.n11183 VSS.t3562 1.6805
R7718 VSS.n9955 VSS.t1314 1.6805
R7719 VSS.n9956 VSS.t3592 1.6805
R7720 VSS.n9957 VSS.t2836 1.6805
R7721 VSS.n9958 VSS.t2968 1.6805
R7722 VSS.n142 VSS.t2179 1.6805
R7723 VSS.n11186 VSS.t1554 1.6805
R7724 VSS.n11185 VSS.t722 1.6805
R7725 VSS.n11184 VSS.t3222 1.6805
R7726 VSS.n11183 VSS.t2441 1.6805
R7727 VSS.n1259 VSS.t2534 1.6805
R7728 VSS.n1258 VSS.t1778 1.6805
R7729 VSS.n1257 VSS.t1896 1.6805
R7730 VSS.n1256 VSS.t1080 1.6805
R7731 VSS.n1236 VSS.t3372 1.6805
R7732 VSS.n1237 VSS.t2618 1.6805
R7733 VSS.n1238 VSS.t2754 1.6805
R7734 VSS.n1239 VSS.t1972 1.6805
R7735 VSS.n1240 VSS.t1360 1.6805
R7736 VSS.n1259 VSS.t1420 1.6805
R7737 VSS.n1258 VSS.t512 1.6805
R7738 VSS.n1257 VSS.t702 1.6805
R7739 VSS.n1256 VSS.t3060 1.6805
R7740 VSS.n1236 VSS.t2259 1.6805
R7741 VSS.n1237 VSS.t1493 1.6805
R7742 VSS.n1238 VSS.t1634 1.6805
R7743 VSS.n1239 VSS.t783 1.6805
R7744 VSS.n1240 VSS.t3260 1.6805
R7745 VSS.n633 VSS.t2369 1.6805
R7746 VSS.n632 VSS.t1609 1.6805
R7747 VSS.n631 VSS.t1734 1.6805
R7748 VSS.n630 VSS.t908 1.6805
R7749 VSS.n643 VSS.t3228 1.6805
R7750 VSS.n9653 VSS.t2447 1.6805
R7751 VSS.n9652 VSS.t2576 1.6805
R7752 VSS.n9651 VSS.t1815 1.6805
R7753 VSS.n9650 VSS.t1165 1.6805
R7754 VSS.n633 VSS.t1225 1.6805
R7755 VSS.n632 VSS.t3522 1.6805
R7756 VSS.n631 VSS.t473 1.6805
R7757 VSS.n630 VSS.t2888 1.6805
R7758 VSS.n643 VSS.t2083 1.6805
R7759 VSS.n9653 VSS.t1316 1.6805
R7760 VSS.n9652 VSS.t1460 1.6805
R7761 VSS.n9651 VSS.t584 1.6805
R7762 VSS.n9650 VSS.t3124 1.6805
R7763 VSS.n603 VSS.t1666 1.6805
R7764 VSS.n608 VSS.t827 1.6805
R7765 VSS.n613 VSS.t965 1.6805
R7766 VSS.n618 VSS.t3280 1.6805
R7767 VSS.n624 VSS.t2486 1.6805
R7768 VSS.n9700 VSS.t2634 1.6805
R7769 VSS.n9705 VSS.t1866 1.6805
R7770 VSS.n9710 VSS.t1051 1.6805
R7771 VSS.n9715 VSS.t1381 1.6805
R7772 VSS.n602 VSS.t1507 1.6805
R7773 VSS.n607 VSS.t634 1.6805
R7774 VSS.n612 VSS.t793 1.6805
R7775 VSS.n617 VSS.t3144 1.6805
R7776 VSS.n625 VSS.t2337 1.6805
R7777 VSS.n9699 VSS.t1586 1.6805
R7778 VSS.n9704 VSS.t1712 1.6805
R7779 VSS.n9709 VSS.t887 1.6805
R7780 VSS.n9714 VSS.t3330 1.6805
R7781 VSS.n589 VSS.t2205 1.6805
R7782 VSS.n588 VSS.t1444 1.6805
R7783 VSS.n587 VSS.t1566 1.6805
R7784 VSS.n586 VSS.t731 1.6805
R7785 VSS.n9915 VSS.t3094 1.6805
R7786 VSS.n582 VSS.t3190 1.6805
R7787 VSS.n581 VSS.t2395 1.6805
R7788 VSS.n580 VSS.t1644 1.6805
R7789 VSS.n579 VSS.t1930 1.6805
R7790 VSS.n589 VSS.t1016 1.6805
R7791 VSS.n588 VSS.t3312 1.6805
R7792 VSS.n587 VSS.t3468 1.6805
R7793 VSS.n586 VSS.t2714 1.6805
R7794 VSS.n9915 VSS.t1926 1.6805
R7795 VSS.n582 VSS.t2036 1.6805
R7796 VSS.n581 VSS.t1266 1.6805
R7797 VSS.n580 VSS.t3556 1.6805
R7798 VSS.n579 VSS.t736 1.6805
R7799 VSS.n11039 VSS.t2822 1.6805
R7800 VSS.n11040 VSS.t2014 1.6805
R7801 VSS.n11041 VSS.t2163 1.6805
R7802 VSS.n11042 VSS.t1387 1.6805
R7803 VSS.n11283 VSS.t478 1.6805
R7804 VSS.n9946 VSS.t667 1.6805
R7805 VSS.n9945 VSS.t3038 1.6805
R7806 VSS.n9944 VSS.t2227 1.6805
R7807 VSS.n9943 VSS.t2512 1.6805
R7808 VSS.n11039 VSS.t1674 1.6805
R7809 VSS.n11040 VSS.t835 1.6805
R7810 VSS.n11041 VSS.t975 1.6805
R7811 VSS.n11042 VSS.t3288 1.6805
R7812 VSS.n11283 VSS.t2508 1.6805
R7813 VSS.n9946 VSS.t2654 1.6805
R7814 VSS.n9945 VSS.t1878 1.6805
R7815 VSS.n9944 VSS.t1063 1.6805
R7816 VSS.n9943 VSS.t1400 1.6805
R7817 VSS.n9477 VSS.t3356 1.6805
R7818 VSS.n9478 VSS.t2590 1.6805
R7819 VSS.n9479 VSS.t1823 1.6805
R7820 VSS.n1385 VSS.t1952 1.6805
R7821 VSS.n1407 VSS.t1333 1.6805
R7822 VSS.n1406 VSS.t3614 1.6805
R7823 VSS.n1405 VSS.t3030 1.6805
R7824 VSS.n1404 VSS.t2221 1.6805
R7825 VSS.n10687 VSS.n10686 1.67828
R7826 VSS.n10678 VSS.n10677 1.67828
R7827 VSS.n10311 VSS.n10292 1.67718
R7828 VSS.n10982 VSS.n181 1.67411
R7829 VSS.n11318 VSS.n11316 1.65519
R7830 VSS.n10632 VSS.n10631 1.60175
R7831 VSS.n10751 VSS.n10750 1.5755
R7832 VSS.n10817 VSS.n10816 1.5755
R7833 VSS.n10780 VSS.n10779 1.5755
R7834 VSS.n10786 VSS.n10785 1.5755
R7835 VSS.n10038 VSS.n238 1.53593
R7836 VSS.n560 VSS.n239 1.53593
R7837 VSS.n11320 VSS.n116 1.53593
R7838 VSS.n10537 VSS.n10536 1.53593
R7839 VSS.n10529 VSS.n10528 1.53593
R7840 VSS.n10613 VSS.n10612 1.5005
R7841 VSS.n10411 VSS.n10410 1.5005
R7842 VSS.n10679 VSS.n10678 1.5005
R7843 VSS.n10334 VSS.n10333 1.5005
R7844 VSS.n10536 VSS.n10535 1.5005
R7845 VSS.n10533 VSS.n10493 1.5005
R7846 VSS.n10530 VSS.n10529 1.5005
R7847 VSS.n558 VSS.n239 1.5005
R7848 VSS.n10869 VSS.n10868 1.5005
R7849 VSS.n238 VSS.n236 1.5005
R7850 VSS.n120 VSS.n117 1.5005
R7851 VSS.n11321 VSS.n11320 1.5005
R7852 VSS.n817 VSS.n650 1.47409
R7853 VSS.n822 VSS.n821 1.47409
R7854 VSS.n9883 VSS.n652 1.47409
R7855 VSS.n678 VSS.n677 1.47409
R7856 VSS.n9880 VSS.n656 1.47409
R7857 VSS.n9859 VSS.n9858 1.47409
R7858 VSS.n9878 VSS.n9877 1.47409
R7859 VSS.n9874 VSS.n9873 1.47409
R7860 VSS.n11413 VSS.n11412 1.47409
R7861 VSS.n11417 VSS.n11416 1.47409
R7862 VSS.n11446 VSS.n11445 1.47409
R7863 VSS.n11450 VSS.n11449 1.47409
R7864 VSS.n9517 VSS.n9516 1.47409
R7865 VSS.n9513 VSS.n9512 1.47409
R7866 VSS.n1249 VSS.n642 1.47409
R7867 VSS.n1254 VSS.n1253 1.47409
R7868 VSS.n9897 VSS.n9896 1.47409
R7869 VSS.n9902 VSS.n9901 1.47409
R7870 VSS.n9914 VSS.n9913 1.47409
R7871 VSS.n9910 VSS.n584 1.47409
R7872 VSS.n9920 VSS.n9919 1.47409
R7873 VSS.n9925 VSS.n9924 1.47409
R7874 VSS.n9612 VSS.n9611 1.47409
R7875 VSS.n9616 VSS.n9615 1.47409
R7876 VSS.n10405 VSS.n10404 1.46537
R7877 VSS.n10409 VSS.n10408 1.46537
R7878 VSS.n10403 VSS.n10402 1.46537
R7879 VSS.n10326 VSS.n10325 1.46537
R7880 VSS.n10330 VSS.n10329 1.46537
R7881 VSS.n10332 VSS.n10331 1.46537
R7882 VSS.n10321 VSS.n10320 1.46537
R7883 VSS.n10319 VSS.n10318 1.46537
R7884 VSS.n10315 VSS.n10314 1.46537
R7885 VSS.n10311 VSS.n10310 1.46537
R7886 VSS.n11316 VSS.n11314 1.37022
R7887 VSS.n10789 VSS.t3120 1.348
R7888 VSS.n10834 VSS.t3544 1.348
R7889 VSS.n10810 VSS.t848 1.348
R7890 VSS.n10812 VSS.t2776 1.348
R7891 VSS.n10775 VSS.t1468 1.348
R7892 VSS.n246 VSS.t1900 1.348
R7893 VSS.n10744 VSS.t2297 1.348
R7894 VSS.n10753 VSS.t1083 1.348
R7895 VSS.n9449 VSS.t3091 1.26547
R7896 VSS.n9423 VSS.t1799 1.26547
R7897 VSS.n9453 VSS.t2480 1.26547
R7898 VSS.n9455 VSS.t1241 1.26547
R7899 VSS.n9429 VSS.t2041 1.26547
R7900 VSS.n9430 VSS.t3519 1.26547
R7901 VSS.n9470 VSS.t3013 1.26547
R7902 VSS.n1378 VSS.t1407 1.26547
R7903 VSS.n129 VSS.t1434 1.26547
R7904 VSS.n10698 VSS.t2795 1.26547
R7905 VSS.n10734 VSS.t1806 1.26547
R7906 VSS.n10824 VSS.t3485 1.26547
R7907 VSS.n10824 VSS.t1715 1.26547
R7908 VSS.n10867 VSS.n10866 1.26528
R7909 VSS.n10802 VSS.n10801 1.265
R7910 VSS.n9204 VSS.t2732 1.2605
R7911 VSS.t632 VSS.n9204 1.2605
R7912 VSS.t2281 VSS.n9060 1.2605
R7913 VSS.n9060 VSS.t3310 1.2605
R7914 VSS.t1517 VSS.n1545 1.2605
R7915 VSS.n1545 VSS.t3516 1.2605
R7916 VSS.t1020 VSS.n1551 1.2605
R7917 VSS.n1551 VSS.t1780 1.2605
R7918 VSS.t2022 VSS.n9173 1.2605
R7919 VSS.n9173 VSS.t3108 1.2605
R7920 VSS.n9135 VSS.t1611 1.2605
R7921 VSS.t2640 VSS.n9135 1.2605
R7922 VSS.n9255 VSS.t2948 1.2605
R7923 VSS.t867 VSS.n9255 1.2605
R7924 VSS.t2403 VSS.n9145 1.2605
R7925 VSS.n9145 VSS.t1718 1.2605
R7926 VSS.t3626 VSS.n9244 1.2605
R7927 VSS.n9244 VSS.t1624 1.2605
R7928 VSS.n9210 VSS.t3132 1.2605
R7929 VSS.t2391 VSS.n9210 1.2605
R7930 VSS.n9313 VSS.t973 1.2605
R7931 VSS.t2047 VSS.n9313 1.2605
R7932 VSS.t2319 VSS.n9216 1.2605
R7933 VSS.n9216 VSS.t1636 1.2605
R7934 VSS.t3350 VSS.n9295 1.2605
R7935 VSS.n9295 VSS.t1375 1.2605
R7936 VSS.n9261 VSS.t1640 1.2605
R7937 VSS.t885 VSS.n9261 1.2605
R7938 VSS.n9353 VSS.t2143 1.2605
R7939 VSS.t2858 VSS.n9353 1.2605
R7940 VSS.t2407 VSS.n9267 1.2605
R7941 VSS.n9267 VSS.t1383 1.2605
R7942 VSS.t2854 VSS.n9342 1.2605
R7943 VSS.n9342 VSS.t3540 1.2605
R7944 VSS.n9319 VSS.t3138 1.2605
R7945 VSS.t2055 VSS.n9319 1.2605
R7946 VSS.n9386 VSS.t475 1.2605
R7947 VSS.t2604 VSS.n9386 1.2605
R7948 VSS.n9379 VSS.t3220 1.2605
R7949 VSS.t2187 VSS.n9379 1.2605
R7950 VSS.t2988 VSS.n9418 1.2605
R7951 VSS.n9418 VSS.t1916 1.2605
R7952 VSS.t2518 VSS.n1493 1.2605
R7953 VSS.n1493 VSS.t1495 1.2605
R7954 VSS.n9533 VSS.t2185 1.2605
R7955 VSS.t1095 VSS.n9533 1.2605
R7956 VSS.t626 VSS.n1401 1.2605
R7957 VSS.n1401 VSS.t1422 1.2605
R7958 VSS.t2032 VSS.n11241 1.2605
R7959 VSS.n11241 VSS.t957 1.2605
R7960 VSS.t2445 VSS.n11247 1.2605
R7961 VSS.n11247 VSS.t3158 1.2605
R7962 VSS.t3566 VSS.n11253 1.2605
R7963 VSS.n11253 VSS.t2878 1.2605
R7964 VSS.n11269 VSS.t1533 1.2605
R7965 VSS.n11269 VSS.t2552 1.2605
R7966 VSS.n11275 VSS.t1123 1.2605
R7967 VSS.n11275 VSS.t1938 1.2605
R7968 VSS.n11166 VSS.t1572 1.2605
R7969 VSS.t2263 VSS.n11166 1.2605
R7970 VSS.t3282 VSS.n744 1.2605
R7971 VSS.n744 VSS.t2231 1.2605
R7972 VSS.n748 VSS.t525 1.2605
R7973 VSS.n748 VSS.t3002 1.2605
R7974 VSS.n756 VSS.t3374 1.2605
R7975 VSS.n756 VSS.t993 1.2605
R7976 VSS.n9832 VSS.t3292 1.2605
R7977 VSS.t2257 VSS.n9832 1.2605
R7978 VSS.n9820 VSS.t553 1.2605
R7979 VSS.t1362 VSS.n9820 1.2605
R7980 VSS.n9809 VSS.t2818 1.2605
R7981 VSS.t2089 VSS.n9809 1.2605
R7982 VSS.n9786 VSS.t2794 1.2605
R7983 VSS.t716 VSS.n9786 1.2605
R7984 VSS.n9773 VSS.t1156 1.2605
R7985 VSS.t3188 VSS.n9773 1.2605
R7986 VSS.t2840 VSS.n9594 1.2605
R7987 VSS.n9594 VSS.t3588 1.2605
R7988 VSS.t2814 VSS.n1451 1.2605
R7989 VSS.n1451 VSS.t3496 1.2605
R7990 VSS.n1457 VSS.t1888 1.2605
R7991 VSS.t1169 VSS.n1457 1.2605
R7992 VSS.t1617 VSS.n1469 1.2605
R7993 VSS.n1469 VSS.t2287 1.2605
R7994 VSS.n11238 VSS.t807 1.2605
R7995 VSS.n11238 VSS.t3208 1.2605
R7996 VSS.n11244 VSS.t3444 1.2605
R7997 VSS.n11244 VSS.t1462 1.2605
R7998 VSS.n11250 VSS.t2970 1.2605
R7999 VSS.n11250 VSS.t1904 1.2605
R8000 VSS.t2155 VSS.n11260 1.2605
R8001 VSS.n11260 VSS.t3196 1.2605
R8002 VSS.n11266 VSS.t3454 1.2605
R8003 VSS.n11266 VSS.t2770 1.2605
R8004 VSS.n11272 VSS.t945 1.2605
R8005 VSS.n11272 VSS.t3314 1.2605
R8006 VSS.n11169 VSS.t597 1.2605
R8007 VSS.t3054 VSS.n11169 1.2605
R8008 VSS.n11160 VSS.t1256 1.2605
R8009 VSS.t2295 VSS.n11160 1.2605
R8010 VSS.t773 VSS.n738 1.2605
R8011 VSS.n738 VSS.t1874 1.2605
R8012 VSS.n741 VSS.t3164 1.2605
R8013 VSS.t2111 VSS.n741 1.2605
R8014 VSS.n752 VSS.t2040 1.2605
R8015 VSS.n752 VSS.t1358 1.2605
R8016 VSS.n759 VSS.t1613 1.2605
R8017 VSS.n759 VSS.t3602 1.2605
R8018 VSS.n9839 VSS.t1129 1.2605
R8019 VSS.t1868 VSS.n9839 1.2605
R8020 VSS.n9827 VSS.t1686 1.2605
R8021 VSS.n9827 VSS.t521 1.2605
R8022 VSS.n9814 VSS.t1059 1.2605
R8023 VSS.n9814 VSS.t2139 1.2605
R8024 VSS.n9804 VSS.t3388 1.2605
R8025 VSS.n9804 VSS.t2365 1.2605
R8026 VSS.n9794 VSS.t1950 1.2605
R8027 VSS.n9794 VSS.t3024 1.2605
R8028 VSS.n9789 VSS.t1215 1.2605
R8029 VSS.t3232 VSS.n9789 1.2605
R8030 VSS.n9778 VSS.t2008 1.2605
R8031 VSS.t2728 VSS.n9778 1.2605
R8032 VSS.n9591 VSS.t1509 1.2605
R8033 VSS.n9591 VSS.t2267 1.2605
R8034 VSS.n9596 VSS.t1012 1.2605
R8035 VSS.t1776 VSS.n9596 1.2605
R8036 VSS.t3364 VSS.n1448 1.2605
R8037 VSS.n1448 VSS.t2329 1.2605
R8038 VSS.t3594 VSS.n1460 1.2605
R8039 VSS.n1460 VSS.t1232 1.2605
R8040 VSS.n1464 VSS.t2886 1.2605
R8041 VSS.n1464 VSS.t1819 1.2605
R8042 VSS.t1418 VSS.n1474 1.2605
R8043 VSS.n1474 VSS.t2097 1.2605
R8044 VSS.n9546 VSS.t743 1.2605
R8045 VSS.t1578 VSS.n9546 1.2605
R8046 VSS.n9539 VSS.t3392 1.2605
R8047 VSS.t1022 VSS.n9539 1.2605
R8048 VSS.t2734 VSS.n1203 1.2605
R8049 VSS.n1203 VSS.t1688 1.2605
R8050 VSS.t1252 VSS.n1213 1.2605
R8051 VSS.n1213 VSS.t2293 1.2605
R8052 VSS.n10935 VSS.t852 1.2605
R8053 VSS.t2934 VSS.n10935 1.2605
R8054 VSS.t3532 VSS.n1167 1.2605
R8055 VSS.n1167 VSS.t1140 1.2605
R8056 VSS.t3630 VSS.n10978 1.2605
R8057 VSS.n10978 VSS.t1628 1.2605
R8058 VSS.n10941 VSS.t3184 1.2605
R8059 VSS.t1150 VSS.n10941 1.2605
R8060 VSS.n11367 VSS.t1470 1.2605
R8061 VSS.t2479 VSS.n11367 1.2605
R8062 VSS.t2784 VSS.n10951 1.2605
R8063 VSS.n10951 VSS.t2057 1.2605
R8064 VSS.n11380 VSS.t1908 1.2605
R8065 VSS.t2974 VSS.n11380 1.2605
R8066 VSS.n11373 VSS.t3216 1.2605
R8067 VSS.t2500 VSS.n11373 1.2605
R8068 VSS.n11323 VSS.t1980 1.2605
R8069 VSS.t2217 VSS.n11323 1.2605
R8070 VSS.t1499 VSS.n11464 1.2605
R8071 VSS.n11464 VSS.t1466 1.2605
R8072 VSS.n11094 VSS.t630 1.2605
R8073 VSS.n11094 VSS.t1720 1.2605
R8074 VSS.n11100 VSS.t2920 1.2605
R8075 VSS.n11100 VSS.t2892 1.2605
R8076 VSS.n11106 VSS.t1049 1.2605
R8077 VSS.n11106 VSS.t1325 1.2605
R8078 VSS.t2488 VSS.n11116 1.2605
R8079 VSS.n11116 VSS.t2463 1.2605
R8080 VSS.t1752 VSS.n11121 1.2605
R8081 VSS.n11121 VSS.t2746 1.2605
R8082 VSS.t1678 VSS.n11127 1.2605
R8083 VSS.n11127 VSS.t2674 1.2605
R8084 VSS.t1304 VSS.n11136 1.2605
R8085 VSS.n11136 VSS.t2309 1.2605
R8086 VSS.t1240 VSS.n11148 1.2605
R8087 VSS.n11148 VSS.t1189 1.2605
R8088 VSS.n10881 VSS.t1519 1.2605
R8089 VSS.t1491 VSS.n10881 1.2605
R8090 VSS.t3436 VSS.n10892 1.2605
R8091 VSS.n10892 VSS.t537 1.2605
R8092 VSS.n10036 VSS.t3412 1.2605
R8093 VSS.n10036 VSS.t1404 1.2605
R8094 VSS.n10043 VSS.t2562 1.2605
R8095 VSS.n10043 VSS.t2828 1.2605
R8096 VSS.t2856 VSS.n10052 1.2605
R8097 VSS.n10052 VSS.t2026 1.2605
R8098 VSS.t2063 VSS.n10058 1.2605
R8099 VSS.n10058 VSS.t2301 1.2605
R8100 VSS.n532 VSS.t2808 1.2605
R8101 VSS.t2760 VSS.n532 1.2605
R8102 VSS.n520 VSS.t1690 1.2605
R8103 VSS.n520 VSS.t1922 1.2605
R8104 VSS.t1114 VSS.n10073 1.2605
R8105 VSS.n10073 VSS.t1085 1.2605
R8106 VSS.n10077 VSS.t3118 1.2605
R8107 VSS.n10077 VSS.t3308 1.2605
R8108 VSS.n10085 VSS.t1148 1.2605
R8109 VSS.n10085 VSS.t3404 1.2605
R8110 VSS.n10091 VSS.t2678 1.2605
R8111 VSS.n10091 VSS.t2554 1.2605
R8112 VSS.t2956 VSS.n10101 1.2605
R8113 VSS.n10101 VSS.t2141 1.2605
R8114 VSS.t1836 VSS.n10106 1.2605
R8115 VSS.n10106 VSS.t2053 1.2605
R8116 VSS.n445 VSS.t2870 1.2605
R8117 VSS.t2038 VSS.n445 1.2605
R8118 VSS.n1305 VSS.t1754 1.2605
R8119 VSS.n1305 VSS.t1978 1.2605
R8120 VSS.n1314 VSS.t1191 1.2605
R8121 VSS.n1314 VSS.t3462 1.2605
R8122 VSS.t2484 VSS.n11097 1.2605
R8123 VSS.n11097 VSS.t2750 1.2605
R8124 VSS.t2451 VSS.n11103 1.2605
R8125 VSS.n11103 VSS.t1670 1.2605
R8126 VSS.t462 VSS.n11109 1.2605
R8127 VSS.n11109 VSS.t1598 1.2605
R8128 VSS.t3620 VSS.n11124 1.2605
R8129 VSS.n11124 VSS.t3580 1.2605
R8130 VSS.t2868 VSS.n11130 1.2605
R8131 VSS.n11130 VSS.t2744 1.2605
R8132 VSS.n11133 VSS.t2816 1.2605
R8133 VSS.t2002 VSS.n11133 1.2605
R8134 VSS.n10887 VSS.t904 1.2605
R8135 VSS.n10887 VSS.t1167 1.2605
R8136 VSS.n10871 VSS.t845 1.2605
R8137 VSS.t1906 VSS.n10871 1.2605
R8138 VSS.n10040 VSS.t771 1.2605
R8139 VSS.n10040 VSS.t3112 1.2605
R8140 VSS.n10055 VSS.t2367 1.2605
R8141 VSS.n10055 VSS.t2606 1.2605
R8142 VSS.n10062 VSS.t2317 1.2605
R8143 VSS.n10062 VSS.t1539 1.2605
R8144 VSS.n525 VSS.t1234 1.2605
R8145 VSS.t2235 VSS.n525 1.2605
R8146 VSS.t3476 VSS.n10082 1.2605
R8147 VSS.n10082 VSS.t3432 1.2605
R8148 VSS.t2357 VSS.n10088 1.2605
R8149 VSS.n10088 VSS.t2602 1.2605
R8150 VSS.t2666 VSS.n10094 1.2605
R8151 VSS.n10094 VSS.t2550 1.2605
R8152 VSS.t1854 VSS.n10109 1.2605
R8153 VSS.n10109 VSS.t1006 1.2605
R8154 VSS.n10113 VSS.t712 1.2605
R8155 VSS.n10113 VSS.t1784 1.2605
R8156 VSS.t604 VSS.n1310 1.2605
R8157 VSS.n1310 VSS.t2966 1.2605
R8158 VSS.t2409 VSS.n11344 1.2605
R8159 VSS.n11344 VSS.t2377 1.2605
R8160 VSS.t1664 VSS.n11351 1.2605
R8161 VSS.n11351 VSS.t2656 1.2605
R8162 VSS.t3426 VSS.n11357 1.2605
R8163 VSS.n11357 VSS.t3384 1.2605
R8164 VSS.t2684 VSS.n10997 1.2605
R8165 VSS.n10997 VSS.t519 1.2605
R8166 VSS.n10988 VSS.t2189 1.2605
R8167 VSS.t2153 VSS.n10988 1.2605
R8168 VSS.t2429 VSS.n10919 1.2605
R8169 VSS.n10919 VSS.t2397 1.2605
R8170 VSS.n10643 VSS.t2588 1.2605
R8171 VSS.n10643 VSS.t791 1.2605
R8172 VSS.t1654 VSS.n10647 1.2605
R8173 VSS.n10647 VSS.t2588 1.2605
R8174 VSS.t1074 VSS.n10652 1.2605
R8175 VSS.n10652 VSS.t2399 1.2605
R8176 VSS.t2850 VSS.n10519 1.2605
R8177 VSS.n10519 VSS.t661 1.2605
R8178 VSS.n10520 VSS.t2930 1.2605
R8179 VSS.n10520 VSS.t2850 1.2605
R8180 VSS.n10526 VSS.t1033 1.2605
R8181 VSS.n10526 VSS.t2289 1.2605
R8182 VSS.n10501 VSS.t3176 1.2605
R8183 VSS.t1033 VSS.n10501 1.2605
R8184 VSS.t2632 VSS.n10546 1.2605
R8185 VSS.n10546 VSS.t3596 1.2605
R8186 VSS.n10547 VSS.t1694 1.2605
R8187 VSS.n10547 VSS.t2632 1.2605
R8188 VSS.n10653 VSS.t1171 1.2605
R8189 VSS.n10653 VSS.t1074 1.2605
R8190 VSS.n10514 VSS.t571 1.2605
R8191 VSS.t878 VSS.n10514 1.2605
R8192 VSS.t2756 VSS.n10523 1.2605
R8193 VSS.n10523 VSS.t571 1.2605
R8194 VSS.n10541 VSS.t892 1.2605
R8195 VSS.t1894 VSS.n10541 1.2605
R8196 VSS.t3062 VSS.n10550 1.2605
R8197 VSS.n10550 VSS.t892 1.2605
R8198 VSS.n10588 VSS.t3264 1.2605
R8199 VSS.t1146 VSS.n10588 1.2605
R8200 VSS.n10437 VSS.t3560 1.2605
R8201 VSS.t1475 VSS.n10437 1.2605
R8202 VSS.n10433 VSS.t2582 1.2605
R8203 VSS.n10433 VSS.t3560 1.2605
R8204 VSS.n10430 VSS.t2852 1.2605
R8205 VSS.t663 VSS.n10430 1.2605
R8206 VSS.n10425 VSS.t2932 1.2605
R8207 VSS.n10425 VSS.t2852 1.2605
R8208 VSS.n10422 VSS.t2373 1.2605
R8209 VSS.t2291 VSS.n10422 1.2605
R8210 VSS.n10418 VSS.t1440 1.2605
R8211 VSS.n10418 VSS.t2373 1.2605
R8212 VSS.n10455 VSS.t3262 1.2605
R8213 VSS.n10455 VSS.t1144 1.2605
R8214 VSS.t3316 VSS.n10459 1.2605
R8215 VSS.n10459 VSS.t3262 1.2605
R8216 VSS.n10462 VSS.t1525 1.2605
R8217 VSS.n10462 VSS.t2738 1.2605
R8218 VSS.t3606 VSS.n10467 1.2605
R8219 VSS.n10467 VSS.t1525 1.2605
R8220 VSS.n10470 VSS.t3106 1.2605
R8221 VSS.n10470 VSS.t926 1.2605
R8222 VSS.t2119 VSS.n10474 1.2605
R8223 VSS.n10474 VSS.t3106 1.2605
R8224 VSS.n10583 VSS.t3318 1.2605
R8225 VSS.n10583 VSS.t3264 1.2605
R8226 VSS.n10580 VSS.t2838 1.2605
R8227 VSS.t2740 VSS.n10580 1.2605
R8228 VSS.n10576 VSS.t1860 1.2605
R8229 VSS.n10576 VSS.t2838 1.2605
R8230 VSS.n9037 VSS.t803 1.2605
R8231 VSS.t2880 VSS.n9037 1.2605
R8232 VSS.t3470 VSS.n1569 1.2605
R8233 VSS.n1569 VSS.t1087 1.2605
R8234 VSS.t3212 VSS.n9006 1.2605
R8235 VSS.n9006 VSS.t2177 1.2605
R8236 VSS.n8968 VSS.t2802 1.2605
R8237 VSS.t3478 VSS.n8968 1.2605
R8238 VSS.n9098 VSS.t2073 1.2605
R8239 VSS.t991 VSS.n9098 1.2605
R8240 VSS.t498 VSS.n8978 1.2605
R8241 VSS.n8978 VSS.t1672 1.2605
R8242 VSS.t2798 VSS.n9087 1.2605
R8243 VSS.n9087 VSS.t1742 1.2605
R8244 VSS.n9043 VSS.t1302 1.2605
R8245 VSS.t2343 VSS.n9043 1.2605
R8246 VSS.t2201 VSS.n9066 1.2605
R8247 VSS.n9066 VSS.t1107 1.2605
R8248 VSS.t1774 VSS.n9072 1.2605
R8249 VSS.n9072 VSS.t2453 1.2605
R8250 VSS.n973 VSS.t1920 1.2605
R8251 VSS.t2161 VSS.n973 1.2605
R8252 VSS.n967 VSS.t2191 1.2605
R8253 VSS.t1396 VSS.n967 1.2605
R8254 VSS.t922 VSS.n10270 1.2605
R8255 VSS.n10270 VSS.t1199 1.2605
R8256 VSS.t1245 VSS.n10276 1.2605
R8257 VSS.n10276 VSS.t3498 1.2605
R8258 VSS.n311 VSS.t3074 1.2605
R8259 VSS.t3272 VSS.n311 1.2605
R8260 VSS.n305 VSS.t2494 1.2605
R8261 VSS.t2465 VSS.n305 1.2605
R8262 VSS.n989 VSS.t876 1.2605
R8263 VSS.t1121 VSS.n989 1.2605
R8264 VSS.n983 VSS.t3428 1.2605
R8265 VSS.t3386 VSS.n983 1.2605
R8266 VSS.n1010 VSS.t2169 1.2605
R8267 VSS.t2379 VSS.n1010 1.2605
R8268 VSS.n1004 VSS.t2411 1.2605
R8269 VSS.t1638 VSS.n1004 1.2605
R8270 VSS.n10222 VSS.t1209 1.2605
R8271 VSS.t1479 VSS.n10222 1.2605
R8272 VSS.n317 VSS.t1501 1.2605
R8273 VSS.t599 VSS.n317 1.2605
R8274 VSS.t3200 VSS.n10210 1.2605
R8275 VSS.n10210 VSS.t3174 1.2605
R8276 VSS.t3450 VSS.n10216 1.2605
R8277 VSS.n10216 VSS.t3406 1.2605
R8278 VSS.n1022 VSS.t1043 1.2605
R8279 VSS.t1004 VSS.n1022 1.2605
R8280 VSS.n1016 VSS.t1350 1.2605
R8281 VSS.t1309 VSS.n1016 1.2605
R8282 VSS.n1047 VSS.t2339 1.2605
R8283 VSS.t2311 VSS.n1047 1.2605
R8284 VSS.n1041 VSS.t1932 1.2605
R8285 VSS.t2952 VSS.n1041 1.2605
R8286 VSS.n374 VSS.t1428 1.2605
R8287 VSS.t1394 VSS.n374 1.2605
R8288 VSS.n368 VSS.t938 1.2605
R8289 VSS.t1990 VSS.n368 1.2605
R8290 VSS.n10162 VSS.t3420 1.2605
R8291 VSS.t3380 VSS.n10162 1.2605
R8292 VSS.n389 VSS.t2676 1.2605
R8293 VSS.t509 VSS.n389 1.2605
R8294 VSS.n1059 VSS.t1329 1.2605
R8295 VSS.t1284 VSS.n1059 1.2605
R8296 VSS.n1053 VSS.t3612 1.2605
R8297 VSS.t1570 VSS.n1053 1.2605
R8298 VSS.n1080 VSS.t3466 1.2605
R8299 VSS.t2680 VSS.n1080 1.2605
R8300 VSS.n1074 VSS.t1910 1.2605
R8301 VSS.t2149 VSS.n1074 1.2605
R8302 VSS.t2528 VSS.n10150 1.2605
R8303 VSS.n10150 VSS.t1748 1.2605
R8304 VSS.t918 VSS.n10156 1.2605
R8305 VSS.n10156 VSS.t1187 1.2605
R8306 VSS.n1293 VSS.t3130 1.2605
R8307 VSS.t3322 VSS.n1293 1.2605
R8308 VSS.n1287 VSS.t3354 1.2605
R8309 VSS.t3618 VSS.n1287 1.2605
R8310 VSS.n1096 VSS.t955 1.2605
R8311 VSS.t1223 VSS.n1096 1.2605
R8312 VSS.n1090 VSS.t1254 1.2605
R8313 VSS.t1513 VSS.n1090 1.2605
R8314 VSS.n1117 VSS.t2692 1.2605
R8315 VSS.t2938 VSS.n1117 1.2605
R8316 VSS.n1111 VSS.t2157 1.2605
R8317 VSS.t1364 VSS.n1111 1.2605
R8318 VSS.n1129 VSS.t3616 1.2605
R8319 VSS.t3510 VSS.n1129 1.2605
R8320 VSS.n1123 VSS.t760 1.2605
R8321 VSS.t3110 VSS.n1123 1.2605
R8322 VSS.t2612 VSS.n865 1.2605
R8323 VSS.n865 VSS.t2874 1.2605
R8324 VSS.t2079 VSS.n876 1.2605
R8325 VSS.n876 VSS.t2051 1.2605
R8326 VSS.t3518 VSS.n10925 1.2605
R8327 VSS.n10925 VSS.t612 1.2605
R8328 VSS.t636 VSS.n841 1.2605
R8329 VSS.n841 VSS.t2996 1.2605
R8330 VSS.n10363 VSS.t2171 1.2605
R8331 VSS.t3452 VSS.n10363 1.2605
R8332 VSS.n10359 VSS.t1181 1.2605
R8333 VSS.n10359 VSS.t2171 1.2605
R8334 VSS.n10356 VSS.t588 1.2605
R8335 VSS.t1974 VSS.n10356 1.2605
R8336 VSS.t684 VSS.n10668 1.2605
R8337 VSS.n10668 VSS.t588 1.2605
R8338 VSS.n10671 VSS.t3270 1.2605
R8339 VSS.n10671 VSS.t3542 1.2605
R8340 VSS.t2307 VSS.n10675 1.2605
R8341 VSS.n10675 VSS.t3270 1.2605
R8342 VSS.n10406 VSS.t275 1.2605
R8343 VSS.n10406 VSS.t203 1.2605
R8344 VSS.n10407 VSS.t202 1.2605
R8345 VSS.n10407 VSS.t198 1.2605
R8346 VSS.n10399 VSS.t29 1.2605
R8347 VSS.n10399 VSS.t43 1.2605
R8348 VSS.n10400 VSS.t28 1.2605
R8349 VSS.n10400 VSS.t17 1.2605
R8350 VSS.n10393 VSS.t205 1.2605
R8351 VSS.n10393 VSS.t136 1.2605
R8352 VSS.n10395 VSS.t51 1.2605
R8353 VSS.n10395 VSS.t31 1.2605
R8354 VSS.n10389 VSS.t131 1.2605
R8355 VSS.n10389 VSS.t46 1.2605
R8356 VSS.n10387 VSS.t128 1.2605
R8357 VSS.n10387 VSS.t124 1.2605
R8358 VSS.n10624 VSS.t349 1.2605
R8359 VSS.n10624 VSS.t133 1.2605
R8360 VSS.n10615 VSS.t138 1.2605
R8361 VSS.n10615 VSS.t30 1.2605
R8362 VSS.n10379 VSS.t129 1.2605
R8363 VSS.n10379 VSS.t47 1.2605
R8364 VSS.n10373 VSS.t19 1.2605
R8365 VSS.n10373 VSS.t132 1.2605
R8366 VSS.n10300 VSS.t27 1.2605
R8367 VSS.n10300 VSS.t194 1.2605
R8368 VSS.n10296 VSS.t123 1.2605
R8369 VSS.n10296 VSS.t34 1.2605
R8370 VSS.n10323 VSS.t143 1.2605
R8371 VSS.n10323 VSS.t5 1.2605
R8372 VSS.n10324 VSS.t200 1.2605
R8373 VSS.n10324 VSS.t6 1.2605
R8374 VSS.n10327 VSS.t23 1.2605
R8375 VSS.n10327 VSS.t274 1.2605
R8376 VSS.n10328 VSS.t206 1.2605
R8377 VSS.n10328 VSS.t16 1.2605
R8378 VSS.n10316 VSS.t32 1.2605
R8379 VSS.n10316 VSS.t41 1.2605
R8380 VSS.n10317 VSS.t1 1.2605
R8381 VSS.n10317 VSS.t199 1.2605
R8382 VSS.n10312 VSS.t204 1.2605
R8383 VSS.n10312 VSS.t45 1.2605
R8384 VSS.n10313 VSS.t50 1.2605
R8385 VSS.n10313 VSS.t120 1.2605
R8386 VSS.n10307 VSS.t201 1.2605
R8387 VSS.n10307 VSS.t48 1.2605
R8388 VSS.n10304 VSS.t122 1.2605
R8389 VSS.n10304 VSS.t12 1.2605
R8390 VSS.n9472 VSS.t3014 1.2605
R8391 VSS.t1408 VSS.n9472 1.2605
R8392 VSS.t2043 VSS.n9432 1.2605
R8393 VSS.n9432 VSS.t3520 1.2605
R8394 VSS.t2482 VSS.n9457 1.2605
R8395 VSS.n9457 VSS.t1243 1.2605
R8396 VSS.n9451 VSS.t3092 1.2605
R8397 VSS.t1801 VSS.n9451 1.2605
R8398 VSS.n9613 VSS.t229 1.2605
R8399 VSS.n9613 VSS.t217 1.2605
R8400 VSS.n813 VSS.t220 1.2605
R8401 VSS.n813 VSS.t243 1.2605
R8402 VSS.t3178 VSS.n9977 1.2605
R8403 VSS.n9977 VSS.t1035 1.2605
R8404 VSS.t1028 VSS.n9983 1.2605
R8405 VSS.n9983 VSS.t2363 1.2605
R8406 VSS.t3152 VSS.n9989 1.2605
R8407 VSS.n9989 VSS.t3098 1.2605
R8408 VSS.t1858 VSS.n9999 1.2605
R8409 VSS.n9999 VSS.t2127 1.2605
R8410 VSS.t1590 VSS.n10005 1.2605
R8411 VSS.n10005 VSS.t741 1.2605
R8412 VSS.t2524 VSS.n10011 1.2605
R8413 VSS.n10011 VSS.t733 1.2605
R8414 VSS.t2351 VSS.n10023 1.2605
R8415 VSS.n10023 VSS.t3304 1.2605
R8416 VSS.n10028 VSS.t3302 1.2605
R8417 VSS.n10028 VSS.t3236 1.2605
R8418 VSS.t906 VSS.n9726 1.2605
R8419 VSS.n9726 VSS.t2249 1.2605
R8420 VSS.t2522 VSS.n9736 1.2605
R8421 VSS.n9736 VSS.t3484 1.2605
R8422 VSS.t3480 VSS.n9742 1.2605
R8423 VSS.n9742 VSS.t1740 1.2605
R8424 VSS.t1730 VSS.n9748 1.2605
R8425 VSS.n9748 VSS.t1662 1.2605
R8426 VSS.t1201 VSS.n9758 1.2605
R8427 VSS.n9758 VSS.t1497 1.2605
R8428 VSS.n9762 VSS.t2237 1.2605
R8429 VSS.n9762 VSS.t3202 1.2605
R8430 VSS.n9632 VSS.t1892 1.2605
R8431 VSS.t1065 VSS.n9632 1.2605
R8432 VSS.t1389 VSS.n1361 1.2605
R8433 VSS.n1361 VSS.t2704 1.2605
R8434 VSS.t2690 VSS.n1367 1.2605
R8435 VSS.n1367 VSS.t2592 1.2605
R8436 VSS.t3334 VSS.n1373 1.2605
R8437 VSS.n1373 VSS.t1630 1.2605
R8438 VSS.n9973 VSS.t1912 1.2605
R8439 VSS.t811 VSS.n9973 1.2605
R8440 VSS.n9971 VSS.t2303 1.2605
R8441 VSS.t3036 VSS.n9971 1.2605
R8442 VSS.n9969 VSS.t3396 1.2605
R8443 VSS.t2730 VSS.n9969 1.2605
R8444 VSS.n9941 VSS.t1398 1.2605
R8445 VSS.t2417 VSS.n9941 1.2605
R8446 VSS.n9939 VSS.t977 1.2605
R8447 VSS.t1805 VSS.n9939 1.2605
R8448 VSS.n9937 VSS.t1442 1.2605
R8449 VSS.t2125 VSS.n9937 1.2605
R8450 VSS.n575 VSS.t3160 1.2605
R8451 VSS.t2099 VSS.n575 1.2605
R8452 VSS.t3554 VSS.n570 1.2605
R8453 VSS.t2864 VSS.n570 1.2605
R8454 VSS.n9720 VSS.t3254 1.2605
R8455 VSS.t854 VSS.n9720 1.2605
R8456 VSS.n9669 VSS.t3172 1.2605
R8457 VSS.t2121 VSS.n9669 1.2605
R8458 VSS.n9667 VSS.t3570 1.2605
R8459 VSS.t1193 VSS.n9667 1.2605
R8460 VSS.n9664 VSS.t2662 1.2605
R8461 VSS.t1958 VSS.n9664 1.2605
R8462 VSS.n9637 VSS.t2636 1.2605
R8463 VSS.t523 VSS.n9637 1.2605
R8464 VSS.t997 VSS.n799 1.2605
R8465 VSS.t3086 VSS.n799 1.2605
R8466 VSS.n9630 VSS.t2694 1.2605
R8467 VSS.n9630 VSS.t3434 1.2605
R8468 VSS.n1352 VSS.t2660 1.2605
R8469 VSS.t3332 VSS.n1352 1.2605
R8470 VSS.n1350 VSS.t1768 1.2605
R8471 VSS.t1001 VSS.n1350 1.2605
R8472 VSS.n1347 VSS.t1485 1.2605
R8473 VSS.t2173 VSS.n1347 1.2605
R8474 VSS.n670 VSS.t78 1.2605
R8475 VSS.n670 VSS.t86 1.2605
R8476 VSS.n9875 VSS.t85 1.2605
R8477 VSS.n9875 VSS.t53 1.2605
R8478 VSS.n669 VSS.t55 1.2605
R8479 VSS.n669 VSS.t69 1.2605
R8480 VSS.n9857 VSS.t73 1.2605
R8481 VSS.n9857 VSS.t59 1.2605
R8482 VSS.n9855 VSS.t79 1.2605
R8483 VSS.n9855 VSS.t70 1.2605
R8484 VSS.n655 VSS.t87 1.2605
R8485 VSS.n655 VSS.t80 1.2605
R8486 VSS.n676 VSS.t236 1.2605
R8487 VSS.n676 VSS.t246 1.2605
R8488 VSS.n674 VSS.t245 1.2605
R8489 VSS.n674 VSS.t221 1.2605
R8490 VSS.n651 VSS.t241 1.2605
R8491 VSS.n651 VSS.t219 1.2605
R8492 VSS.n820 VSS.t242 1.2605
R8493 VSS.n820 VSS.t232 1.2605
R8494 VSS.n818 VSS.t216 1.2605
R8495 VSS.n818 VSS.t238 1.2605
R8496 VSS.n816 VSS.t212 1.2605
R8497 VSS.n816 VSS.t235 1.2605
R8498 VSS.n11414 VSS.t62 1.2605
R8499 VSS.n11414 VSS.t75 1.2605
R8500 VSS.n46 VSS.t93 1.2605
R8501 VSS.n46 VSS.t67 1.2605
R8502 VSS.n45 VSS.t76 1.2605
R8503 VSS.n45 VSS.t83 1.2605
R8504 VSS.n11447 VSS.t65 1.2605
R8505 VSS.n11447 VSS.t82 1.2605
R8506 VSS.n21 VSS.t68 1.2605
R8507 VSS.n21 VSS.t84 1.2605
R8508 VSS.n20 VSS.t77 1.2605
R8509 VSS.n20 VSS.t88 1.2605
R8510 VSS.n9923 VSS.t74 1.2605
R8511 VSS.n9923 VSS.t57 1.2605
R8512 VSS.n9921 VSS.t72 1.2605
R8513 VSS.n9921 VSS.t56 1.2605
R8514 VSS.n585 VSS.t81 1.2605
R8515 VSS.n585 VSS.t71 1.2605
R8516 VSS.n9909 VSS.t92 1.2605
R8517 VSS.n9909 VSS.t91 1.2605
R8518 VSS.n9911 VSS.t90 1.2605
R8519 VSS.n9911 VSS.t89 1.2605
R8520 VSS.n9908 VSS.t64 1.2605
R8521 VSS.n9908 VSS.t60 1.2605
R8522 VSS.n9900 VSS.t215 1.2605
R8523 VSS.n9900 VSS.t231 1.2605
R8524 VSS.n9898 VSS.t228 1.2605
R8525 VSS.n9898 VSS.t237 1.2605
R8526 VSS.n629 VSS.t233 1.2605
R8527 VSS.n629 VSS.t248 1.2605
R8528 VSS.n1252 VSS.t234 1.2605
R8529 VSS.n1252 VSS.t247 1.2605
R8530 VSS.n1250 VSS.t244 1.2605
R8531 VSS.n1250 VSS.t224 1.2605
R8532 VSS.n1248 VSS.t222 1.2605
R8533 VSS.n1248 VSS.t230 1.2605
R8534 VSS.n1329 VSS.t240 1.2605
R8535 VSS.n1329 VSS.t239 1.2605
R8536 VSS.n9514 VSS.t210 1.2605
R8537 VSS.n9514 VSS.t208 1.2605
R8538 VSS.n1328 VSS.t227 1.2605
R8539 VSS.n1328 VSS.t225 1.2605
R8540 VSS.n812 VSS.t226 1.2605
R8541 VSS.n812 VSS.t213 1.2605
R8542 VSS.n10391 VSS.n10390 1.25428
R8543 VSS.n10397 VSS.n10396 1.25428
R8544 VSS.n10394 VSS.n10392 1.25428
R8545 VSS.n10409 VSS.n10405 1.25428
R8546 VSS.n10315 VSS.n10311 1.25428
R8547 VSS.n10321 VSS.n10319 1.25428
R8548 VSS.n10332 VSS.n10330 1.25428
R8549 VSS.n10306 VSS.n10305 1.25428
R8550 VSS.n11392 VSS.n11391 1.21249
R8551 VSS.n10611 VSS.n10439 1.13691
R8552 VSS.n10803 VSS.t38 1.1205
R8553 VSS.n10803 VSS.t127 1.1205
R8554 VSS.n10805 VSS.t165 1.1205
R8555 VSS.n10805 VSS.t158 1.1205
R8556 VSS.n10797 VSS.t169 1.1205
R8557 VSS.n10797 VSS.t197 1.1205
R8558 VSS.n10799 VSS.t3 1.1205
R8559 VSS.n10799 VSS.t21 1.1205
R8560 VSS.n10817 VSS.t1914 1.1205
R8561 VSS.t3210 VSS.n10817 1.1205
R8562 VSS.t586 VSS.n10751 1.1205
R8563 VSS.n10751 VSS.t894 1.1205
R8564 VSS.n10786 VSS.t2239 1.1205
R8565 VSS.t3550 VSS.n10786 1.1205
R8566 VSS.n10780 VSS.t967 1.1205
R8567 VSS.t1268 VSS.n10780 1.1205
R8568 VSS.n10442 VSS.t11 1.11868
R8569 VSS.t167 VSS.n10600 1.11868
R8570 VSS.n10663 VSS.t26 1.11868
R8571 VSS.n10383 VSS.n10382 0.9995
R8572 VSS.n10619 VSS.n10618 0.9995
R8573 VSS.n10628 VSS.n10627 0.9995
R8574 VSS.n10683 VSS.n10682 0.973625
R8575 VSS.n10612 VSS.n10611 0.970331
R8576 VSS.n9048 VSS.t3584 0.918039
R8577 VSS.n9049 VSS.t2812 0.918039
R8578 VSS.n1528 VSS.t3136 0.918039
R8579 VSS.n9119 VSS.t1944 0.918039
R8580 VSS.n9124 VSS.t1544 0.918039
R8581 VSS.n9128 VSS.t2906 0.918039
R8582 VSS.n9055 VSS.t1632 0.918039
R8583 VSS.n9052 VSS.t763 0.918039
R8584 VSS.n1529 VSS.t1101 0.918039
R8585 VSS.n9120 VSS.t3046 0.918039
R8586 VSS.n9125 VSS.t2614 0.918039
R8587 VSS.n9129 VSS.t871 0.918039
R8588 VSS.n9218 VSS.t1876 0.918039
R8589 VSS.n9219 VSS.t1040 0.918039
R8590 VSS.n9220 VSS.t1416 0.918039
R8591 VSS.n9221 VSS.t3276 0.918039
R8592 VSS.n9222 VSS.t2898 0.918039
R8593 VSS.n1509 VSS.t1152 0.918039
R8594 VSS.n9238 VSS.t1373 0.918039
R8595 VSS.n9235 VSS.t3636 0.918039
R8596 VSS.n9231 VSS.t837 0.918039
R8597 VSS.n9228 VSS.t2782 0.918039
R8598 VSS.n9224 VSS.t2353 0.918039
R8599 VSS.n1510 VSS.t577 0.918039
R8600 VSS.n1501 VSS.t1541 0.918039
R8601 VSS.n9270 VSS.t674 0.918039
R8602 VSS.n9275 VSS.t1010 0.918039
R8603 VSS.n9279 VSS.t2960 0.918039
R8604 VSS.n9284 VSS.t2532 0.918039
R8605 VSS.n9288 VSS.t785 0.918039
R8606 VSS.n1502 VSS.t727 0.918039
R8607 VSS.n9271 VSS.t3070 0.918039
R8608 VSS.n9276 VSS.t3328 0.918039
R8609 VSS.n9280 VSS.t2195 0.918039
R8610 VSS.n9285 VSS.t1792 0.918039
R8611 VSS.n9289 VSS.t3150 0.918039
R8612 VSS.n1479 VSS.t2780 0.918039
R8613 VSS.n1480 VSS.t1976 0.918039
R8614 VSS.n1481 VSS.t2283 0.918039
R8615 VSS.n1483 VSS.t1089 0.918039
R8616 VSS.n1484 VSS.t639 0.918039
R8617 VSS.n1485 VSS.t2065 0.918039
R8618 VSS.n9373 VSS.t2253 0.918039
R8619 VSS.n9370 VSS.t1487 0.918039
R8620 VSS.n9366 VSS.t1794 0.918039
R8621 VSS.n9363 VSS.t481 0.918039
R8622 VSS.n9359 VSS.t3256 0.918039
R8623 VSS.n9356 VSS.t1574 0.918039
R8624 VSS.n9389 VSS.t594 0.918039
R8625 VSS.n9393 VSS.t2958 0.918039
R8626 VSS.n9398 VSS.t3252 0.918039
R8627 VSS.n9402 VSS.t2071 0.918039
R8628 VSS.n9407 VSS.t1692 0.918039
R8629 VSS.n9411 VSS.t3066 0.918039
R8630 VSS.n9390 VSS.t1331 0.918039
R8631 VSS.n9394 VSS.t3590 0.918039
R8632 VSS.n9399 VSS.t805 0.918039
R8633 VSS.n9403 VSS.t2736 0.918039
R8634 VSS.n9408 VSS.t2323 0.918039
R8635 VSS.n9412 VSS.t528 0.918039
R8636 VSS.n1430 VSS.t2584 0.918039
R8637 VSS.n1431 VSS.t2944 0.918039
R8638 VSS.n1223 VSS.t1756 0.918039
R8639 VSS.n1224 VSS.t1341 0.918039
R8640 VSS.n1217 VSS.t2716 0.918039
R8641 VSS.n1436 VSS.t2824 0.918039
R8642 VSS.n1432 VSS.t3142 0.918039
R8643 VSS.n1230 VSS.t1948 0.918039
R8644 VSS.n1226 VSS.t1548 0.918039
R8645 VSS.n1218 VSS.t2916 0.918039
R8646 VSS.n791 VSS.t3490 0.918039
R8647 VSS.n1156 VSS.t693 0.918039
R8648 VSS.n1159 VSS.t2628 0.918039
R8649 VSS.n1160 VSS.t2225 0.918039
R8650 VSS.n1161 VSS.t3586 0.918039
R8651 VSS.n792 VSS.t1219 0.918039
R8652 VSS.n1157 VSS.t1552 0.918039
R8653 VSS.n9556 VSS.t3402 0.918039
R8654 VSS.n9552 VSS.t3050 0.918039
R8655 VSS.n9549 VSS.t1327 0.918039
R8656 VSS.n64 VSS.t3366 0.918039
R8657 VSS.n68 VSS.t561 0.918039
R8658 VSS.n71 VSS.t2530 0.918039
R8659 VSS.n75 VSS.t2135 0.918039
R8660 VSS.n80 VSS.t3482 0.918039
R8661 VSS.n1 VSS.t1091 0.918039
R8662 VSS.n2 VSS.t2586 0.918039
R8663 VSS.n104 VSS.t2942 0.918039
R8664 VSS.n112 VSS.t559 0.918039
R8665 VSS.n113 VSS.t1024 0.918039
R8666 VSS.n114 VSS.t1521 0.918039
R8667 VSS.n115 VSS.t3306 0.918039
R8668 VSS.n1571 VSS.t2752 0.918039
R8669 VSS.n1574 VSS.t1956 0.918039
R8670 VSS.n1578 VSS.t2275 0.918039
R8671 VSS.n8956 VSS.t1067 0.918039
R8672 VSS.n8960 VSS.t618 0.918039
R8673 VSS.n8963 VSS.t2045 0.918039
R8674 VSS.n1557 VSS.t1821 0.918039
R8675 VSS.n8981 VSS.t982 0.918039
R8676 VSS.n8986 VSS.t1356 0.918039
R8677 VSS.n8990 VSS.t3230 0.918039
R8678 VSS.n8995 VSS.t2848 0.918039
R8679 VSS.n8999 VSS.t1093 0.918039
R8680 VSS.n1558 VSS.t2608 0.918039
R8681 VSS.n8982 VSS.t1825 0.918039
R8682 VSS.n8987 VSS.t2145 0.918039
R8683 VSS.n8991 VSS.t911 0.918039
R8684 VSS.n8996 VSS.t3632 0.918039
R8685 VSS.n9000 VSS.t1928 0.918039
R8686 VSS.n9074 VSS.t985 0.918039
R8687 VSS.n9075 VSS.t3290 0.918039
R8688 VSS.n1534 VSS.t3624 0.918039
R8689 VSS.n1538 VSS.t2433 0.918039
R8690 VSS.n1539 VSS.t2030 0.918039
R8691 VSS.n1540 VSS.t3370 0.918039
R8692 VSS.n9081 VSS.t3514 0.918039
R8693 VSS.n9078 VSS.t2724 0.918039
R8694 VSS.n1535 VSS.t3056 0.918039
R8695 VSS.n9108 VSS.t1862 0.918039
R8696 VSS.n9104 VSS.t1473 0.918039
R8697 VSS.n9101 VSS.t2832 0.918039
R8698 VSS.n955 VSS.t1031 0.918039
R8699 VSS.n956 VSS.t1864 0.918039
R8700 VSS.n957 VSS.t2273 0.918039
R8701 VSS.n254 VSS.t2726 0.918039
R8702 VSS.n255 VSS.t1503 0.918039
R8703 VSS.n256 VSS.t3186 0.918039
R8704 VSS.n944 VSS.t2708 0.918039
R8705 VSS.n945 VSS.t3472 0.918039
R8706 VSS.n273 VSS.t781 0.918039
R8707 VSS.n10249 VSS.t1270 0.918039
R8708 VSS.n10254 VSS.t3122 0.918039
R8709 VSS.n10258 VSS.t1760 0.918039
R8710 VSS.n951 VSS.t710 0.918039
R8711 VSS.n948 VSS.t1560 0.918039
R8712 VSS.n274 VSS.t1964 0.918039
R8713 VSS.n10250 VSS.t2387 0.918039
R8714 VSS.n10255 VSS.t1154 0.918039
R8715 VSS.n10259 VSS.t2900 0.918039
R8716 VSS.n991 VSS.t1312 0.918039
R8717 VSS.n992 VSS.t2109 0.918039
R8718 VSS.n283 VSS.t2510 0.918039
R8719 VSS.n286 VSS.t2984 0.918039
R8720 VSS.n294 VSS.t1738 0.918039
R8721 VSS.n298 VSS.t3408 0.918039
R8722 VSS.n998 VSS.t2020 0.918039
R8723 VSS.n995 VSS.t2846 0.918039
R8724 VSS.n284 VSS.t3234 0.918039
R8725 VSS.n287 VSS.t507 0.918039
R8726 VSS.n295 VSS.t2437 0.918039
R8727 VSS.n299 VSS.t1061 0.918039
R8728 VSS.n931 VSS.t2473 0.918039
R8729 VSS.n932 VSS.t3286 0.918039
R8730 VSS.n323 VSS.t556 0.918039
R8731 VSS.n326 VSS.t1057 0.918039
R8732 VSS.n327 VSS.t2940 0.918039
R8733 VSS.n328 VSS.t1576 0.918039
R8734 VSS.n938 VSS.t2223 0.918039
R8735 VSS.n935 VSS.t3048 0.918039
R8736 VSS.n324 VSS.t3416 0.918039
R8737 VSS.n10232 VSS.t766 0.918039
R8738 VSS.n10228 VSS.t2646 0.918039
R8739 VSS.n10225 VSS.t1282 0.918039
R8740 VSS.n1024 VSS.t1856 0.918039
R8741 VSS.n1025 VSS.t2638 0.918039
R8742 VSS.n345 VSS.t3096 0.918039
R8743 VSS.n10189 VSS.t3494 0.918039
R8744 VSS.n10194 VSS.t2269 0.918039
R8745 VSS.n10198 VSS.t865 0.918039
R8746 VSS.n1031 VSS.t1117 0.918039
R8747 VSS.n1028 VSS.t1946 0.918039
R8748 VSS.n346 VSS.t2345 0.918039
R8749 VSS.n10190 VSS.t2820 0.918039
R8750 VSS.n10195 VSS.t1580 0.918039
R8751 VSS.n10199 VSS.t3268 0.918039
R8752 VSS.n918 VSS.t2748 0.918039
R8753 VSS.n919 VSS.t3538 0.918039
R8754 VSS.n355 VSS.t843 0.918039
R8755 VSS.n358 VSS.t1337 0.918039
R8756 VSS.n378 VSS.t3170 0.918039
R8757 VSS.n382 VSS.t1813 0.918039
R8758 VSS.n925 VSS.t883 0.918039
R8759 VSS.n922 VSS.t1722 0.918039
R8760 VSS.n356 VSS.t2133 0.918039
R8761 VSS.n359 VSS.t2564 0.918039
R8762 VSS.n379 VSS.t1343 0.918039
R8763 VSS.n383 VSS.t3080 0.918039
R8764 VSS.n1061 VSS.t1433 0.918039
R8765 VSS.n1062 VSS.t2211 0.918039
R8766 VSS.n395 VSS.t2616 0.918039
R8767 VSS.n398 VSS.t3100 0.918039
R8768 VSS.n399 VSS.t1838 0.918039
R8769 VSS.n400 VSS.t3534 0.918039
R8770 VSS.n1068 VSS.t2175 0.918039
R8771 VSS.n1065 VSS.t2980 0.918039
R8772 VSS.n396 VSS.t3344 0.918039
R8773 VSS.n10172 VSS.t696 0.918039
R8774 VSS.n10168 VSS.t2574 0.918039
R8775 VSS.n10165 VSS.t1217 0.918039
R8776 VSS.n905 VSS.t3430 0.918039
R8777 VSS.n906 VSS.t1160 0.918039
R8778 VSS.n417 VSS.t1615 0.918039
R8779 VSS.n10129 VSS.t2028 0.918039
R8780 VSS.n10134 VSS.t754 0.918039
R8781 VSS.n10138 VSS.t2492 0.918039
R8782 VSS.n912 VSS.t3546 0.918039
R8783 VSS.n909 VSS.t1276 0.918039
R8784 VSS.n418 VSS.t1704 0.918039
R8785 VSS.n10130 VSS.t2137 0.918039
R8786 VSS.n10135 VSS.t859 0.918039
R8787 VSS.n10139 VSS.t2600 0.918039
R8788 VSS.n1098 VSS.t995 0.918039
R8789 VSS.n1099 VSS.t1842 0.918039
R8790 VSS.n425 VSS.t2245 0.918039
R8791 VSS.n428 VSS.t2710 0.918039
R8792 VSS.n1276 VSS.t1481 0.918039
R8793 VSS.n1280 VSS.t3168 0.918039
R8794 VSS.n1105 VSS.t2103 0.918039
R8795 VSS.n1102 VSS.t2910 0.918039
R8796 VSS.n426 VSS.t3294 0.918039
R8797 VSS.n429 VSS.t610 0.918039
R8798 VSS.n1277 VSS.t2502 0.918039
R8799 VSS.n1281 VSS.t1127 0.918039
R8800 VSS.n843 VSS.t3034 0.918039
R8801 VSS.n844 VSS.t677 0.918039
R8802 VSS.n845 VSS.t1125 0.918039
R8803 VSS.n846 VSS.t1619 0.918039
R8804 VSS.n534 VSS.t3400 0.918039
R8805 VSS.n859 VSS.t579 0.918039
R8806 VSS.n856 VSS.t1483 0.918039
R8807 VSS.n852 VSS.t1880 0.918039
R8808 VSS.n849 VSS.t2305 0.918039
R8809 VSS.n535 VSS.t1053 0.918039
R8810 VSS.n1132 VSS.t932 0.918039
R8811 VSS.n1136 VSS.t1786 0.918039
R8812 VSS.n1141 VSS.t2197 0.918039
R8813 VSS.n1144 VSS.t2624 0.918039
R8814 VSS.n1145 VSS.t1412 0.918039
R8815 VSS.n1133 VSS.t2115 0.918039
R8816 VSS.n1137 VSS.t2918 0.918039
R8817 VSS.n1142 VSS.t3300 0.918039
R8818 VSS.n1150 VSS.t621 0.918039
R8819 VSS.n1146 VSS.t2520 0.918039
R8820 VSS.n880 VSS.t2778 0.918039
R8821 VSS.n881 VSS.t3564 0.918039
R8822 VSS.n882 VSS.t874 0.918039
R8823 VSS.n883 VSS.t1369 0.918039
R8824 VSS.n884 VSS.t3182 0.918039
R8825 VSS.n899 VSS.t656 0.918039
R8826 VSS.n896 VSS.t1535 0.918039
R8827 VSS.n892 VSS.t1942 0.918039
R8828 VSS.n889 VSS.t2371 0.918039
R8829 VSS.n885 VSS.t1112 0.918039
R8830 VSS.n224 VSS.t1339 0.918039
R8831 VSS.n231 VSS.t2131 0.918039
R8832 VSS.n232 VSS.t2538 0.918039
R8833 VSS.n233 VSS.t3000 0.918039
R8834 VSS.n234 VSS.t1764 0.918039
R8835 VSS.n10914 VSS.t1323 0.918039
R8836 VSS.n10907 VSS.t2113 0.918039
R8837 VSS.n10903 VSS.t2516 0.918039
R8838 VSS.n10900 VSS.t2990 0.918039
R8839 VSS.n10896 VSS.t1750 0.918039
R8840 VSS.n11000 VSS.t2598 0.918039
R8841 VSS.n11004 VSS.t3368 0.918039
R8842 VSS.n11009 VSS.t687 0.918039
R8843 VSS.n11013 VSS.t1173 0.918039
R8844 VSS.n11018 VSS.t3044 0.918039
R8845 VSS.n11001 VSS.t2251 0.918039
R8846 VSS.n11005 VSS.t3078 0.918039
R8847 VSS.n11010 VSS.t3440 0.918039
R8848 VSS.n11014 VSS.t789 0.918039
R8849 VSS.n11019 VSS.t2670 0.918039
R8850 VSS.n98 VSS.t739 0.918039
R8851 VSS.n11061 VSS.t1588 0.918039
R8852 VSS.n11066 VSS.t1996 0.918039
R8853 VSS.n11070 VSS.t2419 0.918039
R8854 VSS.n11075 VSS.t1177 0.918039
R8855 VSS.n99 VSS.t2012 0.918039
R8856 VSS.n11062 VSS.t2834 0.918039
R8857 VSS.n11067 VSS.t3226 0.918039
R8858 VSS.n11071 VSS.t496 0.918039
R8859 VSS.n11076 VSS.t2425 0.918039
R8860 VSS.n11205 VSS.t2672 0.918039
R8861 VSS.n11206 VSS.t3008 0.918039
R8862 VSS.n11207 VSS.t1817 0.918039
R8863 VSS.n11208 VSS.t1426 0.918039
R8864 VSS.n86 VSS.t2774 0.918039
R8865 VSS.n11221 VSS.t2165 0.918039
R8866 VSS.n11217 VSS.t2461 0.918039
R8867 VSS.n11214 VSS.t1290 0.918039
R8868 VSS.n11210 VSS.t850 0.918039
R8869 VSS.n87 VSS.t2255 0.918039
R8870 VSS.n10953 VSS.t3246 0.918039
R8871 VSS.n10958 VSS.t3576 0.918039
R8872 VSS.n10962 VSS.t2383 0.918039
R8873 VSS.n10967 VSS.t1998 0.918039
R8874 VSS.n10971 VSS.t3324 0.918039
R8875 VSS.n10954 VSS.t2962 0.918039
R8876 VSS.n10959 VSS.t3258 0.918039
R8877 VSS.n10963 VSS.t2077 0.918039
R8878 VSS.n10968 VSS.t1698 0.918039
R8879 VSS.n10972 VSS.t3072 0.918039
R8880 VSS.n707 VSS.t2349 0.918039
R8881 VSS.n708 VSS.t2702 0.918039
R8882 VSS.n709 VSS.t1523 0.918039
R8883 VSS.n710 VSS.t1070 0.918039
R8884 VSS.n210 VSS.t2455 0.918039
R8885 VSS.n723 VSS.t1259 0.918039
R8886 VSS.n719 VSS.t1594 0.918039
R8887 VSS.n716 VSS.t3448 0.918039
R8888 VSS.n712 VSS.t3102 0.918039
R8889 VSS.n211 VSS.t1371 0.918039
R8890 VSS.n766 VSS.t833 0.918039
R8891 VSS.n1171 VSS.t1179 0.918039
R8892 VSS.n1187 VSS.t3114 0.918039
R8893 VSS.n1192 VSS.t2698 0.918039
R8894 VSS.n1196 VSS.t934 0.918039
R8895 VSS.n767 VSS.t3326 0.918039
R8896 VSS.n1172 VSS.t504 0.918039
R8897 VSS.n1188 VSS.t2477 0.918039
R8898 VSS.n1193 VSS.t2091 0.918039
R8899 VSS.n1197 VSS.t3438 0.918039
R8900 VSS.n1519 VSS.t540 0.918039
R8901 VSS.n9148 VSS.t2922 0.918039
R8902 VSS.n9153 VSS.t3218 0.918039
R8903 VSS.n9157 VSS.t2034 0.918039
R8904 VSS.n9162 VSS.t1656 0.918039
R8905 VSS.n9166 VSS.t3026 0.918039
R8906 VSS.n1520 VSS.t2147 0.918039
R8907 VSS.n9149 VSS.t1367 0.918039
R8908 VSS.n9154 VSS.t1684 0.918039
R8909 VSS.n9158 VSS.t3558 0.918039
R8910 VSS.n9163 VSS.t3162 0.918039
R8911 VSS.n9167 VSS.t1464 0.918039
R8912 VSS.n9048 VSS.t2902 0.91749
R8913 VSS.n9049 VSS.t2081 0.91749
R8914 VSS.n1528 VSS.t2393 0.91749
R8915 VSS.n9119 VSS.t1230 0.91749
R8916 VSS.n9124 VSS.t778 0.91749
R8917 VSS.n9128 VSS.t2199 0.91749
R8918 VSS.n9055 VSS.t1790 0.91749
R8919 VSS.n9052 VSS.t943 0.91749
R8920 VSS.n1529 VSS.t1297 0.91749
R8921 VSS.n9120 VSS.t3192 0.91749
R8922 VSS.n9125 VSS.t2806 0.91749
R8923 VSS.n9129 VSS.t1047 0.91749
R8924 VSS.n9218 VSS.t2936 0.91749
R8925 VSS.n9219 VSS.t2129 0.91749
R8926 VSS.n9220 VSS.t2435 0.91749
R8927 VSS.n9221 VSS.t1264 0.91749
R8928 VSS.n9222 VSS.t820 0.91749
R8929 VSS.n1509 VSS.t2219 0.91749
R8930 VSS.n9238 VSS.t3340 0.91749
R8931 VSS.n9235 VSS.t2570 0.91749
R8932 VSS.n9231 VSS.t2914 0.91749
R8933 VSS.n9228 VSS.t1726 0.91749
R8934 VSS.n9224 VSS.t1321 0.91749
R8935 VSS.n1510 VSS.t2682 0.91749
R8936 VSS.n1501 VSS.t2568 0.91749
R8937 VSS.n9270 VSS.t1798 0.91749
R8938 VSS.n9275 VSS.t2107 0.91749
R8939 VSS.n9279 VSS.t890 0.91749
R8940 VSS.n9284 VSS.t3582 0.91749
R8941 VSS.n9288 VSS.t1884 0.91749
R8942 VSS.n1502 VSS.t2804 0.91749
R8943 VSS.n9271 VSS.t1992 0.91749
R8944 VSS.n9276 VSS.t2299 0.91749
R8945 VSS.n9280 VSS.t1097 0.91749
R8946 VSS.n9285 VSS.t653 0.91749
R8947 VSS.n9289 VSS.t2075 0.91749
R8948 VSS.n1479 VSS.t3460 0.91749
R8949 VSS.n1480 VSS.t2686 0.91749
R8950 VSS.n1481 VSS.t3022 0.91749
R8951 VSS.n1483 VSS.t1830 0.91749
R8952 VSS.n1484 VSS.t1438 0.91749
R8953 VSS.n1485 VSS.t2788 0.91749
R8954 VSS.n9373 VSS.t1183 0.91749
R8955 VSS.n9370 VSS.t3464 0.91749
R8956 VSS.n9366 VSS.t659 0.91749
R8957 VSS.n9363 VSS.t2610 0.91749
R8958 VSS.n9359 VSS.t2215 0.91749
R8959 VSS.n9356 VSS.t3568 0.91749
R8960 VSS.n9389 VSS.t2696 0.91749
R8961 VSS.n9393 VSS.t1890 0.91749
R8962 VSS.n9398 VSS.t2213 0.91749
R8963 VSS.n9402 VSS.t989 0.91749
R8964 VSS.n9407 VSS.t534 0.91749
R8965 VSS.n9411 VSS.t1984 0.91749
R8966 VSS.n9390 VSS.t2018 0.91749
R8967 VSS.n9394 VSS.t1228 0.91749
R8968 VSS.n9399 VSS.t1568 0.91749
R8969 VSS.n9403 VSS.t3414 0.91749
R8970 VSS.n9408 VSS.t3058 0.91749
R8971 VSS.n9412 VSS.t1335 0.91749
R8972 VSS.n1430 VSS.t1558 0.91749
R8973 VSS.n1431 VSS.t1872 0.91749
R8974 VSS.n1223 VSS.t615 0.91749
R8975 VSS.n1224 VSS.t3320 0.91749
R8976 VSS.n1217 VSS.t1660 0.91749
R8977 VSS.n1436 VSS.t3508 0.91749
R8978 VSS.n1432 VSS.t714 0.91749
R8979 VSS.n1230 VSS.t2650 0.91749
R8980 VSS.n1226 VSS.t2241 0.91749
R8981 VSS.n1218 VSS.t3600 0.91749
R8982 VSS.n791 VSS.t2427 0.91749
R8983 VSS.n1156 VSS.t2768 0.91749
R8984 VSS.n1159 VSS.t1603 0.91749
R8985 VSS.n1160 VSS.t1163 0.91749
R8986 VSS.n1161 VSS.t2536 0.91749
R8987 VSS.n792 VSS.t1936 0.91749
R8988 VSS.n1157 VSS.t2243 0.91749
R8989 VSS.n9556 VSS.t1037 0.91749
R8990 VSS.n9552 VSS.t582 0.91749
R8991 VSS.n9549 VSS.t2016 0.91749
R8992 VSS.n64 VSS.t2331 0.91749
R8993 VSS.n68 VSS.t2664 0.91749
R8994 VSS.n71 VSS.t1505 0.91749
R8995 VSS.n75 VSS.t1045 0.91749
R8996 VSS.n80 VSS.t2423 0.91749
R8997 VSS.n1 VSS.t3148 0.91749
R8998 VSS.n2 VSS.t467 0.91749
R8999 VSS.n104 VSS.t3166 0.91749
R9000 VSS.n112 VSS.t840 0.91749
R9001 VSS.n113 VSS.t1295 0.91749
R9002 VSS.n114 VSS.t1758 0.91749
R9003 VSS.n115 VSS.t3574 0.91749
R9004 VSS.n1571 VSS.t1710 0.91749
R9005 VSS.n1574 VSS.t862 0.91749
R9006 VSS.n1578 VSS.t1221 0.91749
R9007 VSS.n8956 VSS.t3128 0.91749
R9008 VSS.n8960 VSS.t2720 0.91749
R9009 VSS.n8963 VSS.t963 0.91749
R9010 VSS.n1557 VSS.t2580 0.91749
R9011 VSS.n8981 VSS.t1811 0.91749
R9012 VSS.n8986 VSS.t2123 0.91749
R9013 VSS.n8990 VSS.t902 0.91749
R9014 VSS.n8995 VSS.t3598 0.91749
R9015 VSS.n8999 VSS.t1902 0.91749
R9016 VSS.n1558 VSS.t3298 0.91749
R9017 VSS.n8982 VSS.t2514 0.91749
R9018 VSS.n8987 VSS.t2860 0.91749
R9019 VSS.n8991 VSS.t1682 0.91749
R9020 VSS.n8996 VSS.t1262 0.91749
R9021 VSS.n9000 VSS.t2622 0.91749
R9022 VSS.n9074 VSS.t3076 0.91749
R9023 VSS.n9075 VSS.t2247 0.91749
R9024 VSS.n1534 VSS.t2560 0.91749
R9025 VSS.n1538 VSS.t1410 0.91749
R9026 VSS.n1539 VSS.t950 0.91749
R9027 VSS.n1540 VSS.t2335 0.91749
R9028 VSS.n9081 VSS.t1511 0.91749
R9029 VSS.n9078 VSS.t624 0.91749
R9030 VSS.n1535 VSS.t979 0.91749
R9031 VSS.n9108 VSS.t2926 0.91749
R9032 VSS.n9104 VSS.t2475 0.91749
R9033 VSS.n9101 VSS.t748 0.91749
R9034 VSS.n955 VSS.t1300 0.91749
R9035 VSS.n956 VSS.t2095 0.91749
R9036 VSS.n957 VSS.t2498 0.91749
R9037 VSS.n254 VSS.t2978 0.91749
R9038 VSS.n255 VSS.t1728 0.91749
R9039 VSS.n256 VSS.t3398 0.91749
R9040 VSS.n944 VSS.t2572 0.91749
R9041 VSS.n945 VSS.t3342 0.91749
R9042 VSS.n273 VSS.t650 0.91749
R9043 VSS.n10249 VSS.t1134 0.91749
R9044 VSS.n10254 VSS.t3020 0.91749
R9045 VSS.n10258 VSS.t1650 0.91749
R9046 VSS.n951 VSS.t3040 0.91749
R9047 VSS.n948 VSS.t690 0.91749
R9048 VSS.n274 VSS.t1138 0.91749
R9049 VSS.n10250 VSS.t1626 0.91749
R9050 VSS.n10255 VSS.t3410 0.91749
R9051 VSS.n10259 VSS.t2069 0.91749
R9052 VSS.n991 VSS.t1562 0.91749
R9053 VSS.n992 VSS.t2333 0.91749
R9054 VSS.n283 VSS.t2764 0.91749
R9055 VSS.n286 VSS.t3198 0.91749
R9056 VSS.n294 VSS.t1966 0.91749
R9057 VSS.n298 VSS.t493 0.91749
R9058 VSS.n998 VSS.t2000 0.91749
R9059 VSS.n995 VSS.t2810 0.91749
R9060 VSS.n284 VSS.t3204 0.91749
R9061 VSS.n287 VSS.t465 0.91749
R9062 VSS.n295 VSS.t2401 0.91749
R9063 VSS.n299 VSS.t1014 0.91749
R9064 VSS.n931 VSS.t3512 0.91749
R9065 VSS.n932 VSS.t1238 0.91749
R9066 VSS.n323 VSS.t1668 0.91749
R9067 VSS.n326 VSS.t2085 0.91749
R9068 VSS.n327 VSS.t817 0.91749
R9069 VSS.n328 VSS.t2556 0.91749
R9070 VSS.n938 VSS.t3488 0.91749
R9071 VSS.n935 VSS.t1213 0.91749
R9072 VSS.n324 VSS.t1652 0.91749
R9073 VSS.n10232 VSS.t2067 0.91749
R9074 VSS.n10228 VSS.t798 0.91749
R9075 VSS.n10225 VSS.t2542 0.91749
R9076 VSS.n1024 VSS.t2876 0.91749
R9077 VSS.n1025 VSS.t470 0.91749
R9078 VSS.n345 VSS.t961 0.91749
R9079 VSS.n10189 VSS.t1458 0.91749
R9080 VSS.n10194 VSS.t3266 0.91749
R9081 VSS.n10198 VSS.t1924 0.91749
R9082 VSS.n1031 VSS.t2167 0.91749
R9083 VSS.n1028 VSS.t2976 0.91749
R9084 VSS.n346 VSS.t3336 0.91749
R9085 VSS.n10190 VSS.t682 0.91749
R9086 VSS.n10195 VSS.t2566 0.91749
R9087 VSS.n10199 VSS.t1207 0.91749
R9088 VSS.n918 VSS.t2722 0.91749
R9089 VSS.n919 VSS.t3506 0.91749
R9090 VSS.n355 VSS.t814 0.91749
R9091 VSS.n358 VSS.t1288 0.91749
R9092 VSS.n378 VSS.t3146 0.91749
R9093 VSS.n382 VSS.t1788 0.91749
R9094 VSS.n925 VSS.t1132 0.91749
R9095 VSS.n922 VSS.t1954 0.91749
R9096 VSS.n356 VSS.t2359 0.91749
R9097 VSS.n359 VSS.t2830 0.91749
R9098 VSS.n379 VSS.t1596 0.91749
R9099 VSS.n383 VSS.t3278 0.91749
R9100 VSS.n1061 VSS.t1392 0.91749
R9101 VSS.n1062 VSS.t2181 0.91749
R9102 VSS.n395 VSS.t2578 0.91749
R9103 VSS.n398 VSS.t3052 0.91749
R9104 VSS.n399 VSS.t1809 0.91749
R9105 VSS.n400 VSS.t3500 0.91749
R9106 VSS.n1068 VSS.t2385 0.91749
R9107 VSS.n1065 VSS.t3194 0.91749
R9108 VSS.n396 VSS.t3610 0.91749
R9109 VSS.n10172 VSS.t953 0.91749
R9110 VSS.n10168 VSS.t2844 0.91749
R9111 VSS.n10165 VSS.t1489 0.91749
R9112 VSS.n905 VSS.t2652 0.91749
R9113 VSS.n906 VSS.t3418 0.91749
R9114 VSS.n417 VSS.t746 0.91749
R9115 VSS.n10129 VSS.t1236 0.91749
R9116 VSS.n10134 VSS.t3104 0.91749
R9117 VSS.n10138 VSS.t1714 0.91749
R9118 VSS.n912 VSS.t647 0.91749
R9119 VSS.n909 VSS.t1531 0.91749
R9120 VSS.n418 VSS.t1940 0.91749
R9121 VSS.n10130 VSS.t2361 0.91749
R9122 VSS.n10135 VSS.t1105 0.91749
R9123 VSS.n10139 VSS.t2862 0.91749
R9124 VSS.n1098 VSS.t1278 0.91749
R9125 VSS.n1099 VSS.t2061 0.91749
R9126 VSS.n425 VSS.t2467 0.91749
R9127 VSS.n428 VSS.t2950 0.91749
R9128 VSS.n1276 VSS.t1706 0.91749
R9129 VSS.n1280 VSS.t3376 0.91749
R9130 VSS.n1105 VSS.t1293 0.91749
R9131 VSS.n1102 VSS.t2087 0.91749
R9132 VSS.n426 VSS.t2490 0.91749
R9133 VSS.n429 VSS.t2972 0.91749
R9134 VSS.n1277 VSS.t1724 0.91749
R9135 VSS.n1281 VSS.t3394 0.91749
R9136 VSS.n843 VSS.t3242 0.91749
R9137 VSS.n844 VSS.t936 0.91749
R9138 VSS.n845 VSS.t1414 0.91749
R9139 VSS.n846 VSS.t1844 0.91749
R9140 VSS.n534 VSS.t484 0.91749
R9141 VSS.n859 VSS.t543 0.91749
R9142 VSS.n856 VSS.t1450 0.91749
R9143 VSS.n852 VSS.t1850 0.91749
R9144 VSS.n849 VSS.t2277 0.91749
R9145 VSS.n535 VSS.t1008 0.91749
R9146 VSS.n1132 VSS.t1203 0.91749
R9147 VSS.n1136 VSS.t2006 0.91749
R9148 VSS.n1141 VSS.t2413 0.91749
R9149 VSS.n1144 VSS.t2884 0.91749
R9150 VSS.n1145 VSS.t1646 0.91749
R9151 VSS.n1133 VSS.t1306 0.91749
R9152 VSS.n1137 VSS.t2105 0.91749
R9153 VSS.n1142 VSS.t2506 0.91749
R9154 VSS.n1150 VSS.t2982 0.91749
R9155 VSS.n1146 VSS.t1736 0.91749
R9156 VSS.n880 VSS.t3028 0.91749
R9157 VSS.n881 VSS.t671 0.91749
R9158 VSS.n882 VSS.t1119 0.91749
R9159 VSS.n883 VSS.t1607 0.91749
R9160 VSS.n884 VSS.t3390 0.91749
R9161 VSS.n899 VSS.t3012 0.91749
R9162 VSS.n896 VSS.t644 0.91749
R9163 VSS.n892 VSS.t1103 0.91749
R9164 VSS.n889 VSS.t1592 0.91749
R9165 VSS.n885 VSS.t3378 0.91749
R9166 VSS.n224 VSS.t1584 0.91749
R9167 VSS.n231 VSS.t2347 0.91749
R9168 VSS.n232 VSS.t2792 0.91749
R9169 VSS.n233 VSS.t3214 0.91749
R9170 VSS.n234 VSS.t1988 0.91749
R9171 VSS.n10914 VSS.t2315 0.91749
R9172 VSS.n10907 VSS.t3140 0.91749
R9173 VSS.n10903 VSS.t3536 0.91749
R9174 VSS.n10900 VSS.t869 0.91749
R9175 VSS.n10896 VSS.t2742 0.91749
R9176 VSS.n11000 VSS.t3608 0.91749
R9177 VSS.n11004 VSS.t1345 0.91749
R9178 VSS.n11009 VSS.t1772 0.91749
R9179 VSS.n11013 VSS.t2203 0.91749
R9180 VSS.n11018 VSS.t914 0.91749
R9181 VSS.n11001 VSS.t3248 0.91749
R9182 VSS.n11005 VSS.t947 0.91749
R9183 VSS.n11010 VSS.t1424 0.91749
R9184 VSS.n11014 VSS.t1852 0.91749
R9185 VSS.n11019 VSS.t501 0.91749
R9186 VSS.n98 VSS.t698 0.91749
R9187 VSS.n11061 VSS.t1550 0.91749
R9188 VSS.n11066 VSS.t1960 0.91749
R9189 VSS.n11070 VSS.t2381 0.91749
R9190 VSS.n11075 VSS.t1142 0.91749
R9191 VSS.n99 VSS.t2265 0.91749
R9192 VSS.n11062 VSS.t3088 0.91749
R9193 VSS.n11067 VSS.t3456 0.91749
R9194 VSS.n11071 VSS.t801 0.91749
R9195 VSS.n11076 VSS.t2688 0.91749
R9196 VSS.n11205 VSS.t574 0.91749
R9197 VSS.n11206 VSS.t924 0.91749
R9198 VSS.n11207 VSS.t2882 0.91749
R9199 VSS.n11208 VSS.t2449 0.91749
R9200 VSS.n86 VSS.t700 0.91749
R9201 VSS.n11221 VSS.t1076 0.91749
R9202 VSS.n11217 VSS.t1448 0.91749
R9203 VSS.n11214 VSS.t3296 0.91749
R9204 VSS.n11210 VSS.t2928 0.91749
R9205 VSS.n87 VSS.t1185 0.91749
R9206 VSS.n10953 VSS.t2544 0.91749
R9207 VSS.n10958 VSS.t2890 0.91749
R9208 VSS.n10962 VSS.t1708 0.91749
R9209 VSS.n10967 VSS.t1286 0.91749
R9210 VSS.n10971 VSS.t2648 0.91749
R9211 VSS.n10954 VSS.t2229 0.91749
R9212 VSS.n10959 VSS.t2548 0.91749
R9213 VSS.n10963 VSS.t1402 0.91749
R9214 VSS.n10968 VSS.t930 0.91749
R9215 VSS.n10972 VSS.t2325 0.91749
R9216 VSS.n707 VSS.t1318 0.91749
R9217 VSS.n708 VSS.t1648 0.91749
R9218 VSS.n709 VSS.t3524 0.91749
R9219 VSS.n710 VSS.t3134 0.91749
R9220 VSS.n210 VSS.t1430 0.91749
R9221 VSS.n723 VSS.t3622 0.91749
R9222 VSS.n719 VSS.t831 0.91749
R9223 VSS.n716 VSS.t2766 0.91749
R9224 VSS.n712 VSS.t2341 0.91749
R9225 VSS.n211 VSS.t564 0.91749
R9226 VSS.n766 VSS.t2904 0.91749
R9227 VSS.n1171 VSS.t3206 0.91749
R9228 VSS.n1187 VSS.t2024 0.91749
R9229 VSS.n1192 VSS.t1642 0.91749
R9230 VSS.n1196 VSS.t3010 0.91749
R9231 VSS.n767 VSS.t1347 0.91749
R9232 VSS.n1172 VSS.t1676 0.91749
R9233 VSS.n1188 VSS.t3548 0.91749
R9234 VSS.n1193 VSS.t3156 0.91749
R9235 VSS.n1197 VSS.t1456 0.91749
R9236 VSS.n1519 VSS.t3016 0.91749
R9237 VSS.n9148 VSS.t2207 0.91749
R9238 VSS.n9153 VSS.t2504 0.91749
R9239 VSS.n9157 VSS.t1352 0.91749
R9240 VSS.n9162 VSS.t897 0.91749
R9241 VSS.n9166 VSS.t2285 0.91749
R9242 VSS.n1520 VSS.t1454 0.91749
R9243 VSS.n9149 VSS.t551 0.91749
R9244 VSS.n9154 VSS.t916 0.91749
R9245 VSS.n9158 VSS.t2872 0.91749
R9246 VSS.n9163 VSS.t2443 0.91749
R9247 VSS.n9167 VSS.t679 0.91749
R9248 VSS.n10706 VSS.n121 0.823492
R9249 VSS.n120 VSS.n119 0.794733
R9250 VSS.n1182 VSS.t281 0.717763
R9251 VSS.n10612 VSS.n10411 0.585196
R9252 VSS.n10632 VSS.n10365 0.585196
R9253 VSS.n10686 VSS.n10292 0.585196
R9254 VSS.n10678 VSS.n10334 0.585196
R9255 VSS.n9102 VSS.n9101 0.582999
R9256 VSS.n9105 VSS.n9104 0.582999
R9257 VSS.n9109 VSS.n9108 0.582999
R9258 VSS.n1536 VSS.n1535 0.582999
R9259 VSS.n9079 VSS.n9078 0.582999
R9260 VSS.n9082 VSS.n9081 0.582999
R9261 VSS.n9102 VSS.n1540 0.582999
R9262 VSS.n9105 VSS.n1539 0.582999
R9263 VSS.n9109 VSS.n1538 0.582999
R9264 VSS.n1536 VSS.n1534 0.582999
R9265 VSS.n9079 VSS.n9075 0.582999
R9266 VSS.n9082 VSS.n9074 0.582999
R9267 VSS.n9001 VSS.n9000 0.582999
R9268 VSS.n8997 VSS.n8996 0.582999
R9269 VSS.n8992 VSS.n8991 0.582999
R9270 VSS.n8988 VSS.n8987 0.582999
R9271 VSS.n8983 VSS.n8982 0.582999
R9272 VSS.n1559 VSS.n1558 0.582999
R9273 VSS.n9001 VSS.n8999 0.582999
R9274 VSS.n8997 VSS.n8995 0.582999
R9275 VSS.n8992 VSS.n8990 0.582999
R9276 VSS.n8988 VSS.n8986 0.582999
R9277 VSS.n8983 VSS.n8981 0.582999
R9278 VSS.n1559 VSS.n1557 0.582999
R9279 VSS.n8964 VSS.n8963 0.582999
R9280 VSS.n8961 VSS.n8960 0.582999
R9281 VSS.n8957 VSS.n8956 0.582999
R9282 VSS.n1579 VSS.n1578 0.582999
R9283 VSS.n1575 VSS.n1574 0.582999
R9284 VSS.n1572 VSS.n1571 0.582999
R9285 VSS.n536 VSS.n535 0.582999
R9286 VSS.n850 VSS.n849 0.582999
R9287 VSS.n853 VSS.n852 0.582999
R9288 VSS.n857 VSS.n856 0.582999
R9289 VSS.n860 VSS.n859 0.582999
R9290 VSS.n536 VSS.n534 0.582999
R9291 VSS.n850 VSS.n846 0.582999
R9292 VSS.n853 VSS.n845 0.582999
R9293 VSS.n857 VSS.n844 0.582999
R9294 VSS.n860 VSS.n843 0.582999
R9295 VSS.n1147 VSS.n1146 0.582999
R9296 VSS.n1151 VSS.n1150 0.582999
R9297 VSS.n1143 VSS.n1142 0.582999
R9298 VSS.n1138 VSS.n1137 0.582999
R9299 VSS.n1134 VSS.n1133 0.582999
R9300 VSS.n1147 VSS.n1145 0.582999
R9301 VSS.n1151 VSS.n1144 0.582999
R9302 VSS.n1143 VSS.n1141 0.582999
R9303 VSS.n1138 VSS.n1136 0.582999
R9304 VSS.n1134 VSS.n1132 0.582999
R9305 VSS.n886 VSS.n885 0.582999
R9306 VSS.n890 VSS.n889 0.582999
R9307 VSS.n893 VSS.n892 0.582999
R9308 VSS.n897 VSS.n896 0.582999
R9309 VSS.n900 VSS.n899 0.582999
R9310 VSS.n886 VSS.n884 0.582999
R9311 VSS.n890 VSS.n883 0.582999
R9312 VSS.n893 VSS.n882 0.582999
R9313 VSS.n897 VSS.n881 0.582999
R9314 VSS.n900 VSS.n880 0.582999
R9315 VSS.n1282 VSS.n1281 0.582999
R9316 VSS.n1278 VSS.n1277 0.582999
R9317 VSS.n430 VSS.n429 0.582999
R9318 VSS.n427 VSS.n426 0.582999
R9319 VSS.n1103 VSS.n1102 0.582999
R9320 VSS.n1106 VSS.n1105 0.582999
R9321 VSS.n1282 VSS.n1280 0.582999
R9322 VSS.n1278 VSS.n1276 0.582999
R9323 VSS.n430 VSS.n428 0.582999
R9324 VSS.n427 VSS.n425 0.582999
R9325 VSS.n1103 VSS.n1099 0.582999
R9326 VSS.n1106 VSS.n1098 0.582999
R9327 VSS.n10140 VSS.n10139 0.582999
R9328 VSS.n10136 VSS.n10135 0.582999
R9329 VSS.n10131 VSS.n10130 0.582999
R9330 VSS.n419 VSS.n418 0.582999
R9331 VSS.n910 VSS.n909 0.582999
R9332 VSS.n913 VSS.n912 0.582999
R9333 VSS.n10140 VSS.n10138 0.582999
R9334 VSS.n10136 VSS.n10134 0.582999
R9335 VSS.n10131 VSS.n10129 0.582999
R9336 VSS.n419 VSS.n417 0.582999
R9337 VSS.n910 VSS.n906 0.582999
R9338 VSS.n913 VSS.n905 0.582999
R9339 VSS.n10166 VSS.n10165 0.582999
R9340 VSS.n10169 VSS.n10168 0.582999
R9341 VSS.n10173 VSS.n10172 0.582999
R9342 VSS.n397 VSS.n396 0.582999
R9343 VSS.n1066 VSS.n1065 0.582999
R9344 VSS.n1069 VSS.n1068 0.582999
R9345 VSS.n10166 VSS.n400 0.582999
R9346 VSS.n10169 VSS.n399 0.582999
R9347 VSS.n10173 VSS.n398 0.582999
R9348 VSS.n397 VSS.n395 0.582999
R9349 VSS.n1066 VSS.n1062 0.582999
R9350 VSS.n1069 VSS.n1061 0.582999
R9351 VSS.n384 VSS.n383 0.582999
R9352 VSS.n380 VSS.n379 0.582999
R9353 VSS.n360 VSS.n359 0.582999
R9354 VSS.n357 VSS.n356 0.582999
R9355 VSS.n923 VSS.n922 0.582999
R9356 VSS.n926 VSS.n925 0.582999
R9357 VSS.n384 VSS.n382 0.582999
R9358 VSS.n380 VSS.n378 0.582999
R9359 VSS.n360 VSS.n358 0.582999
R9360 VSS.n357 VSS.n355 0.582999
R9361 VSS.n923 VSS.n919 0.582999
R9362 VSS.n926 VSS.n918 0.582999
R9363 VSS.n10200 VSS.n10199 0.582999
R9364 VSS.n10196 VSS.n10195 0.582999
R9365 VSS.n10191 VSS.n10190 0.582999
R9366 VSS.n347 VSS.n346 0.582999
R9367 VSS.n1029 VSS.n1028 0.582999
R9368 VSS.n1032 VSS.n1031 0.582999
R9369 VSS.n10200 VSS.n10198 0.582999
R9370 VSS.n10196 VSS.n10194 0.582999
R9371 VSS.n10191 VSS.n10189 0.582999
R9372 VSS.n347 VSS.n345 0.582999
R9373 VSS.n1029 VSS.n1025 0.582999
R9374 VSS.n1032 VSS.n1024 0.582999
R9375 VSS.n10226 VSS.n10225 0.582999
R9376 VSS.n10229 VSS.n10228 0.582999
R9377 VSS.n10233 VSS.n10232 0.582999
R9378 VSS.n325 VSS.n324 0.582999
R9379 VSS.n936 VSS.n935 0.582999
R9380 VSS.n939 VSS.n938 0.582999
R9381 VSS.n10226 VSS.n328 0.582999
R9382 VSS.n10229 VSS.n327 0.582999
R9383 VSS.n10233 VSS.n326 0.582999
R9384 VSS.n325 VSS.n323 0.582999
R9385 VSS.n936 VSS.n932 0.582999
R9386 VSS.n939 VSS.n931 0.582999
R9387 VSS.n300 VSS.n299 0.582999
R9388 VSS.n296 VSS.n295 0.582999
R9389 VSS.n288 VSS.n287 0.582999
R9390 VSS.n285 VSS.n284 0.582999
R9391 VSS.n996 VSS.n995 0.582999
R9392 VSS.n999 VSS.n998 0.582999
R9393 VSS.n300 VSS.n298 0.582999
R9394 VSS.n296 VSS.n294 0.582999
R9395 VSS.n288 VSS.n286 0.582999
R9396 VSS.n285 VSS.n283 0.582999
R9397 VSS.n996 VSS.n992 0.582999
R9398 VSS.n999 VSS.n991 0.582999
R9399 VSS.n10260 VSS.n10259 0.582999
R9400 VSS.n10256 VSS.n10255 0.582999
R9401 VSS.n10251 VSS.n10250 0.582999
R9402 VSS.n275 VSS.n274 0.582999
R9403 VSS.n949 VSS.n948 0.582999
R9404 VSS.n952 VSS.n951 0.582999
R9405 VSS.n10260 VSS.n10258 0.582999
R9406 VSS.n10256 VSS.n10254 0.582999
R9407 VSS.n10251 VSS.n10249 0.582999
R9408 VSS.n275 VSS.n273 0.582999
R9409 VSS.n949 VSS.n945 0.582999
R9410 VSS.n952 VSS.n944 0.582999
R9411 VSS.n10278 VSS.n256 0.582999
R9412 VSS.n10280 VSS.n255 0.582999
R9413 VSS.n10283 VSS.n254 0.582999
R9414 VSS.n958 VSS.n957 0.582999
R9415 VSS.n961 VSS.n956 0.582999
R9416 VSS.n963 VSS.n955 0.582999
R9417 VSS.n10897 VSS.n10896 0.582999
R9418 VSS.n10901 VSS.n10900 0.582999
R9419 VSS.n10904 VSS.n10903 0.582999
R9420 VSS.n10908 VSS.n10907 0.582999
R9421 VSS.n10915 VSS.n10914 0.582999
R9422 VSS.n10897 VSS.n234 0.582999
R9423 VSS.n10901 VSS.n233 0.582999
R9424 VSS.n10904 VSS.n232 0.582999
R9425 VSS.n10908 VSS.n231 0.582999
R9426 VSS.n10915 VSS.n224 0.582999
R9427 VSS.n11020 VSS.n11019 0.582999
R9428 VSS.n11015 VSS.n11014 0.582999
R9429 VSS.n11011 VSS.n11010 0.582999
R9430 VSS.n11006 VSS.n11005 0.582999
R9431 VSS.n11002 VSS.n11001 0.582999
R9432 VSS.n11020 VSS.n11018 0.582999
R9433 VSS.n11015 VSS.n11013 0.582999
R9434 VSS.n11011 VSS.n11009 0.582999
R9435 VSS.n11006 VSS.n11004 0.582999
R9436 VSS.n11002 VSS.n11000 0.582999
R9437 VSS.n11077 VSS.n11076 0.582999
R9438 VSS.n11072 VSS.n11071 0.582999
R9439 VSS.n11068 VSS.n11067 0.582999
R9440 VSS.n11063 VSS.n11062 0.582999
R9441 VSS.n100 VSS.n99 0.582999
R9442 VSS.n11077 VSS.n11075 0.582999
R9443 VSS.n11072 VSS.n11070 0.582999
R9444 VSS.n11068 VSS.n11066 0.582999
R9445 VSS.n11063 VSS.n11061 0.582999
R9446 VSS.n100 VSS.n98 0.582999
R9447 VSS.n11326 VSS.n115 0.582999
R9448 VSS.n11329 VSS.n114 0.582999
R9449 VSS.n11331 VSS.n113 0.582999
R9450 VSS.n11334 VSS.n112 0.582999
R9451 VSS.n11339 VSS.n104 0.582999
R9452 VSS.n3 VSS.n2 0.582999
R9453 VSS.n3 VSS.n1 0.582999
R9454 VSS.n81 VSS.n80 0.582999
R9455 VSS.n76 VSS.n75 0.582999
R9456 VSS.n72 VSS.n71 0.582999
R9457 VSS.n69 VSS.n68 0.582999
R9458 VSS.n65 VSS.n64 0.582999
R9459 VSS.n88 VSS.n87 0.582999
R9460 VSS.n11211 VSS.n11210 0.582999
R9461 VSS.n11215 VSS.n11214 0.582999
R9462 VSS.n11218 VSS.n11217 0.582999
R9463 VSS.n11222 VSS.n11221 0.582999
R9464 VSS.n88 VSS.n86 0.582999
R9465 VSS.n11211 VSS.n11208 0.582999
R9466 VSS.n11215 VSS.n11207 0.582999
R9467 VSS.n11218 VSS.n11206 0.582999
R9468 VSS.n11222 VSS.n11205 0.582999
R9469 VSS.n10973 VSS.n10972 0.582999
R9470 VSS.n10969 VSS.n10968 0.582999
R9471 VSS.n10964 VSS.n10963 0.582999
R9472 VSS.n10960 VSS.n10959 0.582999
R9473 VSS.n10955 VSS.n10954 0.582999
R9474 VSS.n10973 VSS.n10971 0.582999
R9475 VSS.n10969 VSS.n10967 0.582999
R9476 VSS.n10964 VSS.n10962 0.582999
R9477 VSS.n10960 VSS.n10958 0.582999
R9478 VSS.n10955 VSS.n10953 0.582999
R9479 VSS.n212 VSS.n211 0.582999
R9480 VSS.n713 VSS.n712 0.582999
R9481 VSS.n717 VSS.n716 0.582999
R9482 VSS.n720 VSS.n719 0.582999
R9483 VSS.n724 VSS.n723 0.582999
R9484 VSS.n212 VSS.n210 0.582999
R9485 VSS.n713 VSS.n710 0.582999
R9486 VSS.n717 VSS.n709 0.582999
R9487 VSS.n720 VSS.n708 0.582999
R9488 VSS.n724 VSS.n707 0.582999
R9489 VSS.n1198 VSS.n1197 0.582999
R9490 VSS.n1194 VSS.n1193 0.582999
R9491 VSS.n1189 VSS.n1188 0.582999
R9492 VSS.n1173 VSS.n1172 0.582999
R9493 VSS.n768 VSS.n767 0.582999
R9494 VSS.n1198 VSS.n1196 0.582999
R9495 VSS.n1194 VSS.n1192 0.582999
R9496 VSS.n1189 VSS.n1187 0.582999
R9497 VSS.n1173 VSS.n1171 0.582999
R9498 VSS.n768 VSS.n766 0.582999
R9499 VSS.n9550 VSS.n9549 0.582999
R9500 VSS.n9553 VSS.n9552 0.582999
R9501 VSS.n9557 VSS.n9556 0.582999
R9502 VSS.n1158 VSS.n1157 0.582999
R9503 VSS.n793 VSS.n792 0.582999
R9504 VSS.n9550 VSS.n1161 0.582999
R9505 VSS.n9553 VSS.n1160 0.582999
R9506 VSS.n9557 VSS.n1159 0.582999
R9507 VSS.n1158 VSS.n1156 0.582999
R9508 VSS.n793 VSS.n791 0.582999
R9509 VSS.n1219 VSS.n1218 0.582999
R9510 VSS.n1227 VSS.n1226 0.582999
R9511 VSS.n1231 VSS.n1230 0.582999
R9512 VSS.n1433 VSS.n1432 0.582999
R9513 VSS.n1437 VSS.n1436 0.582999
R9514 VSS.n1219 VSS.n1217 0.582999
R9515 VSS.n1227 VSS.n1224 0.582999
R9516 VSS.n1231 VSS.n1223 0.582999
R9517 VSS.n1433 VSS.n1431 0.582999
R9518 VSS.n1437 VSS.n1430 0.582999
R9519 VSS.n9413 VSS.n9412 0.582999
R9520 VSS.n9409 VSS.n9408 0.582999
R9521 VSS.n9404 VSS.n9403 0.582999
R9522 VSS.n9400 VSS.n9399 0.582999
R9523 VSS.n9395 VSS.n9394 0.582999
R9524 VSS.n9391 VSS.n9390 0.582999
R9525 VSS.n9413 VSS.n9411 0.582999
R9526 VSS.n9409 VSS.n9407 0.582999
R9527 VSS.n9404 VSS.n9402 0.582999
R9528 VSS.n9400 VSS.n9398 0.582999
R9529 VSS.n9395 VSS.n9393 0.582999
R9530 VSS.n9391 VSS.n9389 0.582999
R9531 VSS.n9357 VSS.n9356 0.582999
R9532 VSS.n9360 VSS.n9359 0.582999
R9533 VSS.n9364 VSS.n9363 0.582999
R9534 VSS.n9367 VSS.n9366 0.582999
R9535 VSS.n9371 VSS.n9370 0.582999
R9536 VSS.n9374 VSS.n9373 0.582999
R9537 VSS.n9357 VSS.n1485 0.582999
R9538 VSS.n9360 VSS.n1484 0.582999
R9539 VSS.n9364 VSS.n1483 0.582999
R9540 VSS.n9367 VSS.n1481 0.582999
R9541 VSS.n9371 VSS.n1480 0.582999
R9542 VSS.n9374 VSS.n1479 0.582999
R9543 VSS.n9290 VSS.n9289 0.582999
R9544 VSS.n9286 VSS.n9285 0.582999
R9545 VSS.n9281 VSS.n9280 0.582999
R9546 VSS.n9277 VSS.n9276 0.582999
R9547 VSS.n9272 VSS.n9271 0.582999
R9548 VSS.n1503 VSS.n1502 0.582999
R9549 VSS.n9290 VSS.n9288 0.582999
R9550 VSS.n9286 VSS.n9284 0.582999
R9551 VSS.n9281 VSS.n9279 0.582999
R9552 VSS.n9277 VSS.n9275 0.582999
R9553 VSS.n9272 VSS.n9270 0.582999
R9554 VSS.n1503 VSS.n1501 0.582999
R9555 VSS.n1511 VSS.n1510 0.582999
R9556 VSS.n9225 VSS.n9224 0.582999
R9557 VSS.n9229 VSS.n9228 0.582999
R9558 VSS.n9232 VSS.n9231 0.582999
R9559 VSS.n9236 VSS.n9235 0.582999
R9560 VSS.n9239 VSS.n9238 0.582999
R9561 VSS.n1511 VSS.n1509 0.582999
R9562 VSS.n9225 VSS.n9222 0.582999
R9563 VSS.n9229 VSS.n9221 0.582999
R9564 VSS.n9232 VSS.n9220 0.582999
R9565 VSS.n9236 VSS.n9219 0.582999
R9566 VSS.n9239 VSS.n9218 0.582999
R9567 VSS.n9168 VSS.n9167 0.582999
R9568 VSS.n9164 VSS.n9163 0.582999
R9569 VSS.n9159 VSS.n9158 0.582999
R9570 VSS.n9155 VSS.n9154 0.582999
R9571 VSS.n9150 VSS.n9149 0.582999
R9572 VSS.n1521 VSS.n1520 0.582999
R9573 VSS.n9168 VSS.n9166 0.582999
R9574 VSS.n9164 VSS.n9162 0.582999
R9575 VSS.n9159 VSS.n9157 0.582999
R9576 VSS.n9155 VSS.n9153 0.582999
R9577 VSS.n9150 VSS.n9148 0.582999
R9578 VSS.n1521 VSS.n1519 0.582999
R9579 VSS.n9130 VSS.n9129 0.582999
R9580 VSS.n9126 VSS.n9125 0.582999
R9581 VSS.n9121 VSS.n9120 0.582999
R9582 VSS.n1530 VSS.n1529 0.582999
R9583 VSS.n9053 VSS.n9052 0.582999
R9584 VSS.n9056 VSS.n9055 0.582999
R9585 VSS.n9130 VSS.n9128 0.582999
R9586 VSS.n9126 VSS.n9124 0.582999
R9587 VSS.n9121 VSS.n9119 0.582999
R9588 VSS.n1530 VSS.n1528 0.582999
R9589 VSS.n9053 VSS.n9049 0.582999
R9590 VSS.n9056 VSS.n9048 0.582999
R9591 VSS.n11292 VSS.t738 0.558372
R9592 VSS.n819 VSS.n817 0.489579
R9593 VSS.n675 VSS.n652 0.489579
R9594 VSS.n9858 VSS.n9856 0.489579
R9595 VSS.n9876 VSS.n9874 0.489579
R9596 VSS.n11415 VSS.n11413 0.489579
R9597 VSS.n11448 VSS.n11446 0.489579
R9598 VSS.n9516 VSS.n9515 0.489579
R9599 VSS.n1251 VSS.n1249 0.489579
R9600 VSS.n9899 VSS.n9897 0.489579
R9601 VSS.n9912 VSS.n9910 0.489579
R9602 VSS.n9924 VSS.n9922 0.489579
R9603 VSS.n9615 VSS.n9614 0.489579
R9604 VSS.n821 VSS.n819 0.486026
R9605 VSS.n677 VSS.n675 0.486026
R9606 VSS.n9856 VSS.n656 0.486026
R9607 VSS.n9877 VSS.n9876 0.486026
R9608 VSS.n11416 VSS.n11415 0.486026
R9609 VSS.n11449 VSS.n11448 0.486026
R9610 VSS.n9515 VSS.n9513 0.486026
R9611 VSS.n1253 VSS.n1251 0.486026
R9612 VSS.n9901 VSS.n9899 0.486026
R9613 VSS.n9913 VSS.n9912 0.486026
R9614 VSS.n9922 VSS.n9920 0.486026
R9615 VSS.n9614 VSS.n9612 0.486026
R9616 VSS.n11314 VSS.n121 0.465835
R9617 VSS.n60 VSS.n59 0.46265
R9618 VSS.n11391 VSS.n11390 0.458898
R9619 VSS.n11317 VSS.n34 0.3755
R9620 VSS.n11319 VSS.n11318 0.3755
R9621 VSS.n11393 VSS.n11392 0.3755
R9622 VSS.n11390 VSS.n11389 0.3755
R9623 VSS.n11316 VSS.n11315 0.3755
R9624 VSS.n11314 VSS.n11313 0.3755
R9625 VSS.n10866 VSS.n10865 0.3755
R9626 VSS.n4804 VSS.n121 0.347815
R9627 VSS.n9461 VSS.n9460 0.240145
R9628 VSS.n9459 VSS.n1379 0.240145
R9629 VSS.n10398 VSS.n10391 0.236091
R9630 VSS.n9460 VSS.n9459 0.207127
R9631 VSS.n10863 VSS.n10862 0.186214
R9632 VSS.n10862 VSS.n10861 0.186214
R9633 VSS.n10858 VSS.n10857 0.186214
R9634 VSS.n10859 VSS.n10858 0.186214
R9635 VSS.n10333 VSS.n10332 0.177184
R9636 VSS.n9142 VSS.n9141 0.174974
R9637 VSS.n1490 VSS.n1489 0.174974
R9638 VSS.n1210 VSS.n1209 0.174974
R9639 VSS.n10948 VSS.n10947 0.174974
R9640 VSS.n10994 VSS.n10993 0.174974
R9641 VSS.n8975 VSS.n8974 0.174974
R9642 VSS.n980 VSS.n979 0.174974
R9643 VSS.n1038 VSS.n1037 0.174974
R9644 VSS.n1087 VSS.n1086 0.174974
R9645 VSS.n873 VSS.n872 0.174974
R9646 VSS.n10765 VSS.n242 0.163
R9647 VSS.n10860 VSS.n242 0.163
R9648 VSS.n10758 VSS.n243 0.163
R9649 VSS.n10860 VSS.n243 0.163
R9650 VSS.n9462 VSS.n9461 0.160263
R9651 VSS.n9468 VSS.n1379 0.160263
R9652 VSS.n9196 VSS.n9193 0.157683
R9653 VSS.n9191 VSS.n9188 0.157683
R9654 VSS.n9332 VSS.n9329 0.157683
R9655 VSS.n9327 VSS.n9324 0.157683
R9656 VSS.n170 VSS.n167 0.157683
R9657 VSS.n165 VSS.n162 0.157683
R9658 VSS.n9578 VSS.n9575 0.157683
R9659 VSS.n9573 VSS.n9570 0.157683
R9660 VSS.n193 VSS.n190 0.157683
R9661 VSS.n198 VSS.n195 0.157683
R9662 VSS.n471 VSS.n468 0.157683
R9663 VSS.n476 VSS.n473 0.157683
R9664 VSS.n9029 VSS.n9026 0.157683
R9665 VSS.n9024 VSS.n9021 0.157683
R9666 VSS.n264 VSS.n261 0.157683
R9667 VSS.n269 VSS.n266 0.157683
R9668 VSS.n336 VSS.n333 0.157683
R9669 VSS.n341 VSS.n338 0.157683
R9670 VSS.n408 VSS.n405 0.157683
R9671 VSS.n413 VSS.n410 0.157683
R9672 VSS.n10864 VSS.n240 0.14444
R9673 VSS.n10853 VSS.n10852 0.141041
R9674 VSS.n10852 VSS.n245 0.141041
R9675 VSS.n10793 VSS.n249 0.141041
R9676 VSS.n10849 VSS.n249 0.141041
R9677 VSS.n10796 VSS.n10795 0.14
R9678 VSS.n10801 VSS.n10795 0.14
R9679 VSS.n10802 VSS.n10794 0.14
R9680 VSS.n10807 VSS.n10794 0.14
R9681 VSS.n10374 VSS.n10372 0.14
R9682 VSS.n10377 VSS.n10372 0.14
R9683 VSS.n10378 VSS.n10371 0.14
R9684 VSS.n10382 VSS.n10371 0.14
R9685 VSS.n10383 VSS.n10370 0.14
R9686 VSS.n10386 VSS.n10370 0.14
R9687 VSS.n10614 VSS.n10369 0.14
R9688 VSS.n10618 VSS.n10369 0.14
R9689 VSS.n10619 VSS.n10368 0.14
R9690 VSS.n10622 VSS.n10368 0.14
R9691 VSS.n10623 VSS.n10367 0.14
R9692 VSS.n10627 VSS.n10367 0.14
R9693 VSS.n10628 VSS.n10366 0.14
R9694 VSS.n10631 VSS.n10366 0.14
R9695 VSS.n10685 VSS.n10293 0.14
R9696 VSS.n10683 VSS.n10293 0.14
R9697 VSS.n10682 VSS.n10295 0.14
R9698 VSS.n10680 VSS.n10295 0.14
R9699 VSS.n10303 VSS.n10298 0.14
R9700 VSS.n10301 VSS.n10298 0.14
R9701 VSS.n10762 VSS.n10739 0.132207
R9702 VSS.n9142 VSS.n9140 0.130788
R9703 VSS.n1490 VSS.n1488 0.130788
R9704 VSS.n1210 VSS.n1208 0.130788
R9705 VSS.n10948 VSS.n10946 0.130788
R9706 VSS.n10994 VSS.n10992 0.130788
R9707 VSS.n8975 VSS.n8973 0.130788
R9708 VSS.n980 VSS.n978 0.130788
R9709 VSS.n1038 VSS.n1036 0.130788
R9710 VSS.n1087 VSS.n1085 0.130788
R9711 VSS.n873 VSS.n871 0.130788
R9712 VSS.n6908 VSS.n6907 0.109625
R9713 VSS.n8233 VSS.n1822 0.109625
R9714 VSS.n6906 VSS.n2263 0.109625
R9715 VSS.n8232 VSS.n8231 0.109625
R9716 VSS.n5469 VSS.n5468 0.10925
R9717 VSS.n4140 VSS.n3184 0.10925
R9718 VSS.n4142 VSS.n4141 0.10925
R9719 VSS.n5470 VSS.n2743 0.10925
R9720 VSS.n10782 VSS.n248 0.108833
R9721 VSS.n10850 VSS.n248 0.108833
R9722 VSS.n10851 VSS.n250 0.108833
R9723 VSS.n10851 VSS.n10850 0.108833
R9724 VSS.n10452 VSS.n10451 0.105988
R9725 VSS.n10478 VSS.n10477 0.105988
R9726 VSS.n10561 VSS.n10560 0.105988
R9727 VSS.n10690 VSS.n10689 0.105988
R9728 VSS.n10640 VSS.n10639 0.105988
R9729 VSS.n10656 VSS.n10655 0.102012
R9730 VSS.n10593 VSS.n10592 0.102012
R9731 VSS.n10613 VSS.n10386 0.10175
R9732 VSS.n10762 VSS.n10759 0.100659
R9733 VSS.n10864 VSS.n10863 0.0996408
R9734 VSS.n11303 VSS.n11302 0.0986132
R9735 VSS.n11302 VSS.n11301 0.0986132
R9736 VSS.n10845 VSS.n10844 0.0986132
R9737 VSS.n10846 VSS.n10845 0.0986132
R9738 VSS.n9440 VSS.n1381 0.0933571
R9739 VSS.n9303 VSS.n1381 0.0933571
R9740 VSS.n1382 VSS.n1344 0.0917281
R9741 VSS.n1392 VSS.n1382 0.0917281
R9742 VSS.n9156 VSS.n1525 0.0886356
R9743 VSS.n9179 VSS.n1525 0.0886356
R9744 VSS.n9176 VSS.n9175 0.0886356
R9745 VSS.n9177 VSS.n9176 0.0886356
R9746 VSS.n9156 VSS.n1514 0.0886356
R9747 VSS.n9178 VSS.n1514 0.0886356
R9748 VSS.n9230 VSS.n1515 0.0886356
R9749 VSS.n1517 VSS.n1515 0.0886356
R9750 VSS.n9251 VSS.n9250 0.0886356
R9751 VSS.n9250 VSS.n9249 0.0886356
R9752 VSS.n9230 VSS.n1506 0.0886356
R9753 VSS.n1516 VSS.n1506 0.0886356
R9754 VSS.n9278 VSS.n1507 0.0886356
R9755 VSS.n9306 VSS.n1507 0.0886356
R9756 VSS.n9298 VSS.n9297 0.0886356
R9757 VSS.n9299 VSS.n9298 0.0886356
R9758 VSS.n9278 VSS.n1497 0.0886356
R9759 VSS.n9305 VSS.n1497 0.0886356
R9760 VSS.n8955 VSS.n1562 0.0886356
R9761 VSS.n1564 VSS.n1562 0.0886356
R9762 VSS.n8989 VSS.n1563 0.0886356
R9763 VSS.n9012 VSS.n1563 0.0886356
R9764 VSS.n9009 VSS.n9008 0.0886356
R9765 VSS.n9010 VSS.n9009 0.0886356
R9766 VSS.n8989 VSS.n1555 0.0886356
R9767 VSS.n9011 VSS.n1555 0.0886356
R9768 VSS.n9110 VSS.n1537 0.0886356
R9769 VSS.n1537 VSS.n1533 0.0886356
R9770 VSS.n9094 VSS.n9093 0.0886356
R9771 VSS.n9093 VSS.n9092 0.0886356
R9772 VSS.n9111 VSS.n9110 0.0886356
R9773 VSS.n9112 VSS.n9111 0.0886356
R9774 VSS.n9118 VSS.n9117 0.0886356
R9775 VSS.n9117 VSS.n9116 0.0886356
R9776 VSS.n1547 VSS.n1532 0.0886356
R9777 VSS.n9113 VSS.n1532 0.0886356
R9778 VSS.n9118 VSS.n1524 0.0886356
R9779 VSS.n9115 VSS.n1524 0.0886356
R9780 VSS.n969 VSS.n251 0.0886356
R9781 VSS.n279 VSS.n251 0.0886356
R9782 VSS.n10285 VSS.n10284 0.0886356
R9783 VSS.n10286 VSS.n10285 0.0886356
R9784 VSS.n10248 VSS.n276 0.0886356
R9785 VSS.n281 VSS.n276 0.0886356
R9786 VSS.n985 VSS.n277 0.0886356
R9787 VSS.n10245 VSS.n277 0.0886356
R9788 VSS.n10248 VSS.n10247 0.0886356
R9789 VSS.n10247 VSS.n10246 0.0886356
R9790 VSS.n10242 VSS.n10241 0.0886356
R9791 VSS.n10243 VSS.n10242 0.0886356
R9792 VSS.n1006 VSS.n289 0.0886356
R9793 VSS.n320 VSS.n289 0.0886356
R9794 VSS.n10241 VSS.n10240 0.0886356
R9795 VSS.n10240 VSS.n282 0.0886356
R9796 VSS.n10234 VSS.n290 0.0886356
R9797 VSS.n10237 VSS.n290 0.0886356
R9798 VSS.n10235 VSS.n10234 0.0886356
R9799 VSS.n10236 VSS.n10235 0.0886356
R9800 VSS.n1018 VSS.n321 0.0886356
R9801 VSS.n351 VSS.n321 0.0886356
R9802 VSS.n10188 VSS.n348 0.0886356
R9803 VSS.n353 VSS.n348 0.0886356
R9804 VSS.n1043 VSS.n349 0.0886356
R9805 VSS.n10185 VSS.n349 0.0886356
R9806 VSS.n10188 VSS.n10187 0.0886356
R9807 VSS.n10187 VSS.n10186 0.0886356
R9808 VSS.n10182 VSS.n10181 0.0886356
R9809 VSS.n10183 VSS.n10182 0.0886356
R9810 VSS.n1055 VSS.n361 0.0886356
R9811 VSS.n392 VSS.n361 0.0886356
R9812 VSS.n10181 VSS.n10180 0.0886356
R9813 VSS.n10180 VSS.n354 0.0886356
R9814 VSS.n10174 VSS.n362 0.0886356
R9815 VSS.n10177 VSS.n362 0.0886356
R9816 VSS.n10175 VSS.n10174 0.0886356
R9817 VSS.n10176 VSS.n10175 0.0886356
R9818 VSS.n1076 VSS.n393 0.0886356
R9819 VSS.n9301 VSS.n393 0.0886356
R9820 VSS.n10128 VSS.n420 0.0886356
R9821 VSS.n423 VSS.n420 0.0886356
R9822 VSS.n1092 VSS.n421 0.0886356
R9823 VSS.n10125 VSS.n421 0.0886356
R9824 VSS.n10128 VSS.n10127 0.0886356
R9825 VSS.n10127 VSS.n10126 0.0886356
R9826 VSS.n10122 VSS.n10121 0.0886356
R9827 VSS.n10123 VSS.n10122 0.0886356
R9828 VSS.n10121 VSS.n10120 0.0886356
R9829 VSS.n10120 VSS.n424 0.0886356
R9830 VSS.n9365 VSS.n1482 0.0886356
R9831 VSS.n1499 VSS.n1482 0.0886356
R9832 VSS.n9349 VSS.n9348 0.0886356
R9833 VSS.n9348 VSS.n9347 0.0886356
R9834 VSS.n9365 VSS.n1384 0.0886356
R9835 VSS.n1498 VSS.n1384 0.0886356
R9836 VSS.n9401 VSS.n1395 0.0886356
R9837 VSS.n1395 VSS.n1394 0.0886356
R9838 VSS.n9421 VSS.n9420 0.0886356
R9839 VSS.n9422 VSS.n9421 0.0886356
R9840 VSS.n9401 VSS.n1222 0.0886356
R9841 VSS.n1393 VSS.n1222 0.0886356
R9842 VSS.n9527 VSS.n1232 0.0886356
R9843 VSS.n9527 VSS.n9526 0.0886356
R9844 VSS.n9529 VSS.n9528 0.0886356
R9845 VSS.n9528 VSS.n434 0.0886356
R9846 VSS.n1232 VSS.n831 0.0886356
R9847 VSS.n9525 VSS.n831 0.0886356
R9848 VSS.n9558 VSS.n832 0.0886356
R9849 VSS.n9561 VSS.n832 0.0886356
R9850 VSS.n9542 VSS.n9541 0.0886356
R9851 VSS.n9541 VSS.n833 0.0886356
R9852 VSS.n9559 VSS.n9558 0.0886356
R9853 VSS.n9560 VSS.n9559 0.0886356
R9854 VSS.n1186 VSS.n1185 0.0886356
R9855 VSS.n1185 VSS.n1184 0.0886356
R9856 VSS.n1205 VSS.n1153 0.0886356
R9857 VSS.n1153 VSS.n506 0.0886356
R9858 VSS.n1186 VSS.n215 0.0886356
R9859 VSS.n1183 VSS.n215 0.0886356
R9860 VSS.n718 VSS.n216 0.0886356
R9861 VSS.n566 VSS.n216 0.0886356
R9862 VSS.n10931 VSS.n10930 0.0886356
R9863 VSS.n10930 VSS.n10929 0.0886356
R9864 VSS.n718 VSS.n179 0.0886356
R9865 VSS.n565 VSS.n179 0.0886356
R9866 VSS.n10961 VSS.n180 0.0886356
R9867 VSS.n180 VSS.n148 0.0886356
R9868 VSS.n10981 VSS.n10980 0.0886356
R9869 VSS.n10982 VSS.n10981 0.0886356
R9870 VSS.n10961 VSS.n91 0.0886356
R9871 VSS.n11279 VSS.n91 0.0886356
R9872 VSS.n11216 VSS.n92 0.0886356
R9873 VSS.n11288 VSS.n92 0.0886356
R9874 VSS.n11363 VSS.n11362 0.0886356
R9875 VSS.n11362 VSS.n11361 0.0886356
R9876 VSS.n11216 VSS.n4 0.0886356
R9877 VSS.n11287 VSS.n4 0.0886356
R9878 VSS.n70 VSS.n5 0.0886356
R9879 VSS.n11298 VSS.n5 0.0886356
R9880 VSS.n11376 VSS.n11375 0.0886356
R9881 VSS.n11375 VSS.n6 0.0886356
R9882 VSS.n1113 VSS.n431 0.0886356
R9883 VSS.n434 VSS.n431 0.0886356
R9884 VSS.n891 VSS.n432 0.0886356
R9885 VSS.n9526 VSS.n432 0.0886356
R9886 VSS.n1125 VSS.n835 0.0886356
R9887 VSS.n835 VSS.n833 0.0886356
R9888 VSS.n891 VSS.n834 0.0886356
R9889 VSS.n9525 VSS.n834 0.0886356
R9890 VSS.n9562 VSS.n1152 0.0886356
R9891 VSS.n9562 VSS.n9561 0.0886356
R9892 VSS.n868 VSS.n867 0.0886356
R9893 VSS.n867 VSS.n506 0.0886356
R9894 VSS.n1152 VSS.n504 0.0886356
R9895 VSS.n9560 VSS.n504 0.0886356
R9896 VSS.n851 VSS.n505 0.0886356
R9897 VSS.n1184 VSS.n505 0.0886356
R9898 VSS.n10928 VSS.n10927 0.0886356
R9899 VSS.n10929 VSS.n10928 0.0886356
R9900 VSS.n851 VSS.n219 0.0886356
R9901 VSS.n1183 VSS.n219 0.0886356
R9902 VSS.n10902 VSS.n220 0.0886356
R9903 VSS.n566 VSS.n220 0.0886356
R9904 VSS.n10984 VSS.n10983 0.0886356
R9905 VSS.n10983 VSS.n10982 0.0886356
R9906 VSS.n10902 VSS.n182 0.0886356
R9907 VSS.n565 VSS.n182 0.0886356
R9908 VSS.n11012 VSS.n183 0.0886356
R9909 VSS.n183 VSS.n148 0.0886356
R9910 VSS.n11360 VSS.n11359 0.0886356
R9911 VSS.n11361 VSS.n11360 0.0886356
R9912 VSS.n11012 VSS.n94 0.0886356
R9913 VSS.n11279 VSS.n94 0.0886356
R9914 VSS.n11069 VSS.n95 0.0886356
R9915 VSS.n11288 VSS.n95 0.0886356
R9916 VSS.n11347 VSS.n11346 0.0886356
R9917 VSS.n11346 VSS.n6 0.0886356
R9918 VSS.n11069 VSS.n7 0.0886356
R9919 VSS.n11287 VSS.n7 0.0886356
R9920 VSS.n11330 VSS.n8 0.0886356
R9921 VSS.n11298 VSS.n8 0.0886356
R9922 VSS.n9182 VSS.n9181 0.0871667
R9923 VSS.n9181 VSS.n9180 0.0871667
R9924 VSS.n9247 VSS.n9246 0.0871667
R9925 VSS.n9248 VSS.n9247 0.0871667
R9926 VSS.n9309 VSS.n9308 0.0871667
R9927 VSS.n9308 VSS.n9307 0.0871667
R9928 VSS.n9015 VSS.n9014 0.0871667
R9929 VSS.n9014 VSS.n9013 0.0871667
R9930 VSS.n9090 VSS.n9089 0.0871667
R9931 VSS.n9091 VSS.n9090 0.0871667
R9932 VSS.n9068 VSS.n1531 0.0871667
R9933 VSS.n9114 VSS.n1531 0.0871667
R9934 VSS.n10272 VSS.n252 0.0871667
R9935 VSS.n280 VSS.n252 0.0871667
R9936 VSS.n307 VSS.n278 0.0871667
R9937 VSS.n10244 VSS.n278 0.0871667
R9938 VSS.n10239 VSS.n319 0.0871667
R9939 VSS.n10239 VSS.n10238 0.0871667
R9940 VSS.n10212 VSS.n322 0.0871667
R9941 VSS.n352 VSS.n322 0.0871667
R9942 VSS.n370 VSS.n350 0.0871667
R9943 VSS.n10184 VSS.n350 0.0871667
R9944 VSS.n10179 VSS.n391 0.0871667
R9945 VSS.n10179 VSS.n10178 0.0871667
R9946 VSS.n10152 VSS.n394 0.0871667
R9947 VSS.n9300 VSS.n394 0.0871667
R9948 VSS.n1289 VSS.n422 0.0871667
R9949 VSS.n10124 VSS.n422 0.0871667
R9950 VSS.n9345 VSS.n9344 0.0871667
R9951 VSS.n9346 VSS.n9345 0.0871667
R9952 VSS.n9382 VSS.n9381 0.0871667
R9953 VSS.n9381 VSS.n1383 0.0871667
R9954 VSS.n1421 VSS.n435 0.0871667
R9955 VSS.n10118 VSS.n435 0.0871667
R9956 VSS.n9566 VSS.n9565 0.0871667
R9957 VSS.n9565 VSS.n9564 0.0871667
R9958 VSS.n9800 VSS.n507 0.0871667
R9959 VSS.n10067 VSS.n507 0.0871667
R9960 VSS.n694 VSS.n693 0.0871667
R9961 VSS.n693 VSS.n218 0.0871667
R9962 VSS.n11154 VSS.n11153 0.0871667
R9963 VSS.n11153 VSS.n11152 0.0871667
R9964 VSS.n11264 VSS.n11263 0.0871667
R9965 VSS.n11263 VSS.n93 0.0871667
R9966 VSS.n11470 VSS.n11469 0.0871667
R9967 VSS.n11469 VSS.n11468 0.0871667
R9968 VSS.n10119 VSS.n433 0.0871667
R9969 VSS.n10119 VSS.n10118 0.0871667
R9970 VSS.n9563 VSS.n458 0.0871667
R9971 VSS.n9564 VSS.n9563 0.0871667
R9972 VSS.n10069 VSS.n10068 0.0871667
R9973 VSS.n10068 VSS.n10067 0.0871667
R9974 VSS.n548 VSS.n547 0.0871667
R9975 VSS.n547 VSS.n218 0.0871667
R9976 VSS.n11151 VSS.n11150 0.0871667
R9977 VSS.n11152 VSS.n11151 0.0871667
R9978 VSS.n11038 VSS.n11037 0.0871667
R9979 VSS.n11037 VSS.n93 0.0871667
R9980 VSS.n11467 VSS.n11466 0.0871667
R9981 VSS.n11468 VSS.n11467 0.0871667
R9982 VSS.n1349 VSS.n438 0.08175
R9983 VSS.n10117 VSS.n438 0.08175
R9984 VSS.n1426 VSS.n437 0.08175
R9985 VSS.n10117 VSS.n437 0.08175
R9986 VSS.n9765 VSS.n9764 0.08175
R9987 VSS.n9766 VSS.n9765 0.08175
R9988 VSS.n9768 VSS.n9767 0.08175
R9989 VSS.n9767 VSS.n9766 0.08175
R9990 VSS.n9666 VSS.n510 0.08175
R9991 VSS.n10066 VSS.n510 0.08175
R9992 VSS.n9816 VSS.n509 0.08175
R9993 VSS.n10066 VSS.n509 0.08175
R9994 VSS.n10031 VSS.n10030 0.08175
R9995 VSS.n10032 VSS.n10031 0.08175
R9996 VSS.n750 VSS.n564 0.08175
R9997 VSS.n10032 VSS.n564 0.08175
R9998 VSS.n149 VSS.n147 0.08175
R9999 VSS.n11279 VSS.n149 0.08175
R10000 VSS.n11278 VSS.n11277 0.08175
R10001 VSS.n11279 VSS.n11278 0.08175
R10002 VSS.n11291 VSS.n138 0.08175
R10003 VSS.n11292 VSS.n11291 0.08175
R10004 VSS.n11226 VSS.n139 0.08175
R10005 VSS.n11292 VSS.n139 0.08175
R10006 VSS.n10116 VSS.n10115 0.08175
R10007 VSS.n10117 VSS.n10116 0.08175
R10008 VSS.n1349 VSS.n436 0.08175
R10009 VSS.n10117 VSS.n436 0.08175
R10010 VSS.n644 VSS.n487 0.08175
R10011 VSS.n9766 VSS.n644 0.08175
R10012 VSS.n9764 VSS.n645 0.08175
R10013 VSS.n9766 VSS.n645 0.08175
R10014 VSS.n10065 VSS.n10064 0.08175
R10015 VSS.n10066 VSS.n10065 0.08175
R10016 VSS.n9666 VSS.n508 0.08175
R10017 VSS.n10066 VSS.n508 0.08175
R10018 VSS.n10034 VSS.n10033 0.08175
R10019 VSS.n10033 VSS.n10032 0.08175
R10020 VSS.n10030 VSS.n563 0.08175
R10021 VSS.n10032 VSS.n563 0.08175
R10022 VSS.n11023 VSS.n145 0.08175
R10023 VSS.n11279 VSS.n145 0.08175
R10024 VSS.n11280 VSS.n147 0.08175
R10025 VSS.n11280 VSS.n11279 0.08175
R10026 VSS.n11081 VSS.n136 0.08175
R10027 VSS.n11292 VSS.n136 0.08175
R10028 VSS.n11293 VSS.n138 0.08175
R10029 VSS.n11293 VSS.n11292 0.08175
R10030 VSS.n10695 VSS.n10694 0.0769706
R10031 VSS.n10696 VSS.n10695 0.0769706
R10032 VSS.n10598 VSS.n10597 0.0769706
R10033 VSS.n10599 VSS.n10598 0.0769706
R10034 VSS.n10661 VSS.n10660 0.0769706
R10035 VSS.n10662 VSS.n10661 0.0769706
R10036 VSS.n10604 VSS.n10603 0.0769706
R10037 VSS.n10603 VSS.n10602 0.0769706
R10038 VSS.n10441 VSS.n10340 0.0769706
R10039 VSS.n10601 VSS.n10340 0.0769706
R10040 VSS.n10341 VSS.n240 0.0769706
R10041 VSS.n10341 VSS.n244 0.0769706
R10042 VSS.n10720 VSS.n131 0.0769706
R10043 VSS.n11300 VSS.n131 0.0769706
R10044 VSS.n10831 VSS.n130 0.0769706
R10045 VSS.n10848 VSS.n130 0.0769706
R10046 VSS.n10597 VSS.n10596 0.072814
R10047 VSS.n10694 VSS.n10693 0.072814
R10048 VSS.n9433 VSS.n9429 0.069264
R10049 VSS.n9431 VSS.n9429 0.069264
R10050 VSS.n9431 VSS.n9430 0.069264
R10051 VSS.n9430 VSS.n1380 0.069264
R10052 VSS.n9470 VSS.n9469 0.069264
R10053 VSS.n9471 VSS.n9470 0.069264
R10054 VSS.n9471 VSS.n1378 0.069264
R10055 VSS.n9473 VSS.n1378 0.069264
R10056 VSS.n10822 VSS.n129 0.0686515
R10057 VSS.n10842 VSS.n10698 0.0686515
R10058 VSS.n9449 VSS.n9448 0.0685756
R10059 VSS.n9450 VSS.n9449 0.0685756
R10060 VSS.n9450 VSS.n9423 0.0685756
R10061 VSS.n9452 VSS.n9423 0.0685756
R10062 VSS.n9458 VSS.n9453 0.0685756
R10063 VSS.n9456 VSS.n9453 0.0685756
R10064 VSS.n9456 VSS.n9455 0.0685756
R10065 VSS.n9455 VSS.n9454 0.0685756
R10066 VSS.n10660 VSS.n10345 0.0681047
R10067 VSS.n10660 VSS.n10659 0.0678953
R10068 VSS.n10844 VSS.n10843 0.0678497
R10069 VSS.n10586 VSS.n10288 0.0646975
R10070 VSS.n10442 VSS.n10288 0.0646975
R10071 VSS.n10464 VSS.n10343 0.0646975
R10072 VSS.n10600 VSS.n10343 0.0646975
R10073 VSS.n10665 VSS.n10664 0.0646975
R10074 VSS.n10664 VSS.n10663 0.0646975
R10075 VSS.n10428 VSS.n10289 0.0646975
R10076 VSS.n10442 VSS.n10289 0.0646975
R10077 VSS.n10349 VSS.n10342 0.0646975
R10078 VSS.n10663 VSS.n10342 0.0646975
R10079 VSS.n10531 VSS.n10344 0.0646975
R10080 VSS.n10600 VSS.n10344 0.0646975
R10081 VSS.n11304 VSS.n11303 0.0640412
R10082 VSS.n10597 VSS.n10481 0.063186
R10083 VSS.n10694 VSS.n10290 0.063186
R10084 VSS.n10841 VSS.n10734 0.0583997
R10085 VSS.n10609 VSS.n10608 0.0533671
R10086 VSS.n9464 VSS.n9463 0.0519852
R10087 VSS.n9465 VSS.n9464 0.0519852
R10088 VSS.n9467 VSS.n9466 0.0519852
R10089 VSS.n9466 VSS.n9465 0.0519852
R10090 VSS.n10534 VSS.n10497 0.0513741
R10091 VSS.n1389 VSS.n1388 0.0490981
R10092 VSS.n1390 VSS.n1389 0.0490981
R10093 VSS.n1235 VSS.n1234 0.0490981
R10094 VSS.n9524 VSS.n1235 0.0490981
R10095 VSS.n1234 VSS.n797 0.0490981
R10096 VSS.n9523 VSS.n797 0.0490981
R10097 VSS.n9887 VSS.n646 0.0490981
R10098 VSS.n9890 VSS.n646 0.0490981
R10099 VSS.n9888 VSS.n9887 0.0490981
R10100 VSS.n9889 VSS.n9888 0.0490981
R10101 VSS.n1181 VSS.n1180 0.0490981
R10102 VSS.n1182 VSS.n1181 0.0490981
R10103 VSS.n1176 VSS.n567 0.0490981
R10104 VSS.n567 VSS.n217 0.0490981
R10105 VSS.n671 VSS.n568 0.0490981
R10106 VSS.n568 VSS.n208 0.0490981
R10107 VSS.n671 VSS.n150 0.0490981
R10108 VSS.n181 VSS.n150 0.0490981
R10109 VSS.n144 VSS.n143 0.0490981
R10110 VSS.n11286 VSS.n144 0.0490981
R10111 VSS.n11290 VSS.n143 0.0490981
R10112 VSS.n11290 VSS.n11289 0.0490981
R10113 VSS.n135 VSS.n134 0.0490981
R10114 VSS.n11297 VSS.n135 0.0490981
R10115 VSS.n1330 VSS.n439 0.0490981
R10116 VSS.n1390 VSS.n439 0.0490981
R10117 VSS.n9521 VSS.n440 0.0490981
R10118 VSS.n9524 VSS.n440 0.0490981
R10119 VSS.n9522 VSS.n9521 0.0490981
R10120 VSS.n9523 VSS.n9522 0.0490981
R10121 VSS.n9892 VSS.n9891 0.0490981
R10122 VSS.n9891 VSS.n9890 0.0490981
R10123 VSS.n9892 VSS.n511 0.0490981
R10124 VSS.n9889 VSS.n511 0.0490981
R10125 VSS.n626 VSS.n512 0.0490981
R10126 VSS.n1182 VSS.n512 0.0490981
R10127 VSS.n623 VSS.n561 0.0490981
R10128 VSS.n561 VSS.n217 0.0490981
R10129 VSS.n9916 VSS.n562 0.0490981
R10130 VSS.n562 VSS.n208 0.0490981
R10131 VSS.n9916 VSS.n146 0.0490981
R10132 VSS.n181 VSS.n146 0.0490981
R10133 VSS.n11285 VSS.n11284 0.0490981
R10134 VSS.n11286 VSS.n11285 0.0490981
R10135 VSS.n11284 VSS.n137 0.0490981
R10136 VSS.n11289 VSS.n137 0.0490981
R10137 VSS.n11296 VSS.n11295 0.0490981
R10138 VSS.n11297 VSS.n11296 0.0490981
R10139 VSS.n9475 VSS.n9473 0.0456011
R10140 VSS.n9454 VSS.n1336 0.0451496
R10141 VSS.n10764 VSS.n10763 0.0431396
R10142 VSS.n10766 VSS.n10738 0.0431396
R10143 VSS.n10768 VSS.n10738 0.0431396
R10144 VSS.n10765 VSS.n10764 0.0420736
R10145 VSS.n1319 VSS.n1318 0.0414574
R10146 VSS.n10450 VSS.n10449 0.041314
R10147 VSS.n10480 VSS.n10479 0.041314
R10148 VSS.n10559 VSS.n10558 0.041314
R10149 VSS.n1416 VSS.n1415 0.0412447
R10150 VSS.n10658 VSS.n10657 0.0411047
R10151 VSS.n10595 VSS.n10594 0.0411047
R10152 VSS.n10692 VSS.n10691 0.0411047
R10153 VSS.n5469 VSS.n2742 0.04025
R10154 VSS.n5473 VSS.n2742 0.04025
R10155 VSS.n5474 VSS.n5473 0.04025
R10156 VSS.n5475 VSS.n5474 0.04025
R10157 VSS.n5475 VSS.n2740 0.04025
R10158 VSS.n5479 VSS.n2740 0.04025
R10159 VSS.n5480 VSS.n5479 0.04025
R10160 VSS.n5481 VSS.n5480 0.04025
R10161 VSS.n5481 VSS.n2738 0.04025
R10162 VSS.n5485 VSS.n2738 0.04025
R10163 VSS.n5486 VSS.n5485 0.04025
R10164 VSS.n5487 VSS.n5486 0.04025
R10165 VSS.n5487 VSS.n2736 0.04025
R10166 VSS.n5491 VSS.n2736 0.04025
R10167 VSS.n5492 VSS.n5491 0.04025
R10168 VSS.n5493 VSS.n5492 0.04025
R10169 VSS.n5493 VSS.n2734 0.04025
R10170 VSS.n5497 VSS.n2734 0.04025
R10171 VSS.n5498 VSS.n5497 0.04025
R10172 VSS.n5499 VSS.n5498 0.04025
R10173 VSS.n5499 VSS.n2732 0.04025
R10174 VSS.n5503 VSS.n2732 0.04025
R10175 VSS.n5504 VSS.n5503 0.04025
R10176 VSS.n5505 VSS.n5504 0.04025
R10177 VSS.n5505 VSS.n2730 0.04025
R10178 VSS.n5509 VSS.n2730 0.04025
R10179 VSS.n5510 VSS.n5509 0.04025
R10180 VSS.n5511 VSS.n5510 0.04025
R10181 VSS.n5511 VSS.n2728 0.04025
R10182 VSS.n5515 VSS.n2728 0.04025
R10183 VSS.n5516 VSS.n5515 0.04025
R10184 VSS.n5517 VSS.n5516 0.04025
R10185 VSS.n5517 VSS.n2726 0.04025
R10186 VSS.n5521 VSS.n2726 0.04025
R10187 VSS.n5522 VSS.n5521 0.04025
R10188 VSS.n5523 VSS.n5522 0.04025
R10189 VSS.n5523 VSS.n2724 0.04025
R10190 VSS.n5527 VSS.n2724 0.04025
R10191 VSS.n5528 VSS.n5527 0.04025
R10192 VSS.n5529 VSS.n5528 0.04025
R10193 VSS.n5529 VSS.n2722 0.04025
R10194 VSS.n5533 VSS.n2722 0.04025
R10195 VSS.n5534 VSS.n5533 0.04025
R10196 VSS.n5535 VSS.n5534 0.04025
R10197 VSS.n5535 VSS.n2720 0.04025
R10198 VSS.n5539 VSS.n2720 0.04025
R10199 VSS.n5540 VSS.n5539 0.04025
R10200 VSS.n5541 VSS.n5540 0.04025
R10201 VSS.n5541 VSS.n2718 0.04025
R10202 VSS.n5545 VSS.n2718 0.04025
R10203 VSS.n5546 VSS.n5545 0.04025
R10204 VSS.n5547 VSS.n5546 0.04025
R10205 VSS.n5547 VSS.n2716 0.04025
R10206 VSS.n5551 VSS.n2716 0.04025
R10207 VSS.n5552 VSS.n5551 0.04025
R10208 VSS.n5553 VSS.n5552 0.04025
R10209 VSS.n5553 VSS.n2714 0.04025
R10210 VSS.n5557 VSS.n2714 0.04025
R10211 VSS.n5558 VSS.n5557 0.04025
R10212 VSS.n5559 VSS.n5558 0.04025
R10213 VSS.n5559 VSS.n2712 0.04025
R10214 VSS.n5563 VSS.n2712 0.04025
R10215 VSS.n5564 VSS.n5563 0.04025
R10216 VSS.n5565 VSS.n5564 0.04025
R10217 VSS.n5565 VSS.n2710 0.04025
R10218 VSS.n5569 VSS.n2710 0.04025
R10219 VSS.n5570 VSS.n5569 0.04025
R10220 VSS.n5571 VSS.n5570 0.04025
R10221 VSS.n5571 VSS.n2708 0.04025
R10222 VSS.n5575 VSS.n2708 0.04025
R10223 VSS.n5576 VSS.n5575 0.04025
R10224 VSS.n5577 VSS.n5576 0.04025
R10225 VSS.n5577 VSS.n2706 0.04025
R10226 VSS.n5581 VSS.n2706 0.04025
R10227 VSS.n5582 VSS.n5581 0.04025
R10228 VSS.n5583 VSS.n5582 0.04025
R10229 VSS.n5583 VSS.n2704 0.04025
R10230 VSS.n5587 VSS.n2704 0.04025
R10231 VSS.n5588 VSS.n5587 0.04025
R10232 VSS.n5589 VSS.n5588 0.04025
R10233 VSS.n5589 VSS.n2702 0.04025
R10234 VSS.n5593 VSS.n2702 0.04025
R10235 VSS.n5594 VSS.n5593 0.04025
R10236 VSS.n5595 VSS.n5594 0.04025
R10237 VSS.n5595 VSS.n2700 0.04025
R10238 VSS.n5599 VSS.n2700 0.04025
R10239 VSS.n5600 VSS.n5599 0.04025
R10240 VSS.n5601 VSS.n5600 0.04025
R10241 VSS.n5601 VSS.n2698 0.04025
R10242 VSS.n5605 VSS.n2698 0.04025
R10243 VSS.n5606 VSS.n5605 0.04025
R10244 VSS.n5607 VSS.n5606 0.04025
R10245 VSS.n5607 VSS.n2696 0.04025
R10246 VSS.n5611 VSS.n2696 0.04025
R10247 VSS.n5612 VSS.n5611 0.04025
R10248 VSS.n5613 VSS.n5612 0.04025
R10249 VSS.n5613 VSS.n2694 0.04025
R10250 VSS.n5617 VSS.n2694 0.04025
R10251 VSS.n5618 VSS.n5617 0.04025
R10252 VSS.n5619 VSS.n5618 0.04025
R10253 VSS.n5619 VSS.n2692 0.04025
R10254 VSS.n5623 VSS.n2692 0.04025
R10255 VSS.n5624 VSS.n5623 0.04025
R10256 VSS.n5625 VSS.n5624 0.04025
R10257 VSS.n5625 VSS.n2690 0.04025
R10258 VSS.n5629 VSS.n2690 0.04025
R10259 VSS.n5630 VSS.n5629 0.04025
R10260 VSS.n5631 VSS.n5630 0.04025
R10261 VSS.n5631 VSS.n2688 0.04025
R10262 VSS.n5635 VSS.n2688 0.04025
R10263 VSS.n5636 VSS.n5635 0.04025
R10264 VSS.n5637 VSS.n5636 0.04025
R10265 VSS.n5637 VSS.n2686 0.04025
R10266 VSS.n5641 VSS.n2686 0.04025
R10267 VSS.n5642 VSS.n5641 0.04025
R10268 VSS.n5643 VSS.n5642 0.04025
R10269 VSS.n5643 VSS.n2684 0.04025
R10270 VSS.n5647 VSS.n2684 0.04025
R10271 VSS.n5648 VSS.n5647 0.04025
R10272 VSS.n5649 VSS.n5648 0.04025
R10273 VSS.n5649 VSS.n2682 0.04025
R10274 VSS.n5653 VSS.n2682 0.04025
R10275 VSS.n5654 VSS.n5653 0.04025
R10276 VSS.n5655 VSS.n5654 0.04025
R10277 VSS.n5655 VSS.n2680 0.04025
R10278 VSS.n5659 VSS.n2680 0.04025
R10279 VSS.n5660 VSS.n5659 0.04025
R10280 VSS.n5661 VSS.n5660 0.04025
R10281 VSS.n5661 VSS.n2678 0.04025
R10282 VSS.n5665 VSS.n2678 0.04025
R10283 VSS.n5666 VSS.n5665 0.04025
R10284 VSS.n5667 VSS.n5666 0.04025
R10285 VSS.n5667 VSS.n2676 0.04025
R10286 VSS.n5671 VSS.n2676 0.04025
R10287 VSS.n5672 VSS.n5671 0.04025
R10288 VSS.n5673 VSS.n5672 0.04025
R10289 VSS.n5673 VSS.n2674 0.04025
R10290 VSS.n5677 VSS.n2674 0.04025
R10291 VSS.n5678 VSS.n5677 0.04025
R10292 VSS.n5679 VSS.n5678 0.04025
R10293 VSS.n5679 VSS.n2672 0.04025
R10294 VSS.n5683 VSS.n2672 0.04025
R10295 VSS.n5684 VSS.n5683 0.04025
R10296 VSS.n5685 VSS.n5684 0.04025
R10297 VSS.n5685 VSS.n2670 0.04025
R10298 VSS.n5689 VSS.n2670 0.04025
R10299 VSS.n5690 VSS.n5689 0.04025
R10300 VSS.n5691 VSS.n5690 0.04025
R10301 VSS.n5691 VSS.n2668 0.04025
R10302 VSS.n5695 VSS.n2668 0.04025
R10303 VSS.n5696 VSS.n5695 0.04025
R10304 VSS.n5697 VSS.n5696 0.04025
R10305 VSS.n5697 VSS.n2666 0.04025
R10306 VSS.n5701 VSS.n2666 0.04025
R10307 VSS.n5702 VSS.n5701 0.04025
R10308 VSS.n5703 VSS.n5702 0.04025
R10309 VSS.n5703 VSS.n2664 0.04025
R10310 VSS.n5707 VSS.n2664 0.04025
R10311 VSS.n5708 VSS.n5707 0.04025
R10312 VSS.n5709 VSS.n5708 0.04025
R10313 VSS.n5709 VSS.n2662 0.04025
R10314 VSS.n5713 VSS.n2662 0.04025
R10315 VSS.n5714 VSS.n5713 0.04025
R10316 VSS.n5715 VSS.n5714 0.04025
R10317 VSS.n5715 VSS.n2660 0.04025
R10318 VSS.n5719 VSS.n2660 0.04025
R10319 VSS.n5720 VSS.n5719 0.04025
R10320 VSS.n5721 VSS.n5720 0.04025
R10321 VSS.n5721 VSS.n2658 0.04025
R10322 VSS.n5725 VSS.n2658 0.04025
R10323 VSS.n5726 VSS.n5725 0.04025
R10324 VSS.n5727 VSS.n5726 0.04025
R10325 VSS.n5727 VSS.n2656 0.04025
R10326 VSS.n5731 VSS.n2656 0.04025
R10327 VSS.n5732 VSS.n5731 0.04025
R10328 VSS.n5733 VSS.n5732 0.04025
R10329 VSS.n5733 VSS.n2654 0.04025
R10330 VSS.n5737 VSS.n2654 0.04025
R10331 VSS.n5738 VSS.n5737 0.04025
R10332 VSS.n5739 VSS.n5738 0.04025
R10333 VSS.n5739 VSS.n2652 0.04025
R10334 VSS.n5743 VSS.n2652 0.04025
R10335 VSS.n5744 VSS.n5743 0.04025
R10336 VSS.n5745 VSS.n5744 0.04025
R10337 VSS.n5745 VSS.n2650 0.04025
R10338 VSS.n5749 VSS.n2650 0.04025
R10339 VSS.n5750 VSS.n5749 0.04025
R10340 VSS.n5751 VSS.n5750 0.04025
R10341 VSS.n5751 VSS.n2648 0.04025
R10342 VSS.n5755 VSS.n2648 0.04025
R10343 VSS.n5756 VSS.n5755 0.04025
R10344 VSS.n5757 VSS.n5756 0.04025
R10345 VSS.n5757 VSS.n2646 0.04025
R10346 VSS.n5761 VSS.n2646 0.04025
R10347 VSS.n5762 VSS.n5761 0.04025
R10348 VSS.n5763 VSS.n5762 0.04025
R10349 VSS.n5763 VSS.n2644 0.04025
R10350 VSS.n5767 VSS.n2644 0.04025
R10351 VSS.n5768 VSS.n5767 0.04025
R10352 VSS.n5769 VSS.n5768 0.04025
R10353 VSS.n5769 VSS.n2642 0.04025
R10354 VSS.n5773 VSS.n2642 0.04025
R10355 VSS.n5774 VSS.n5773 0.04025
R10356 VSS.n5775 VSS.n5774 0.04025
R10357 VSS.n5775 VSS.n2640 0.04025
R10358 VSS.n5779 VSS.n2640 0.04025
R10359 VSS.n5780 VSS.n5779 0.04025
R10360 VSS.n5781 VSS.n5780 0.04025
R10361 VSS.n5781 VSS.n2638 0.04025
R10362 VSS.n5785 VSS.n2638 0.04025
R10363 VSS.n5786 VSS.n5785 0.04025
R10364 VSS.n5787 VSS.n5786 0.04025
R10365 VSS.n5787 VSS.n2636 0.04025
R10366 VSS.n5791 VSS.n2636 0.04025
R10367 VSS.n5792 VSS.n5791 0.04025
R10368 VSS.n5793 VSS.n5792 0.04025
R10369 VSS.n5793 VSS.n2634 0.04025
R10370 VSS.n5797 VSS.n2634 0.04025
R10371 VSS.n5798 VSS.n5797 0.04025
R10372 VSS.n5799 VSS.n5798 0.04025
R10373 VSS.n5799 VSS.n2632 0.04025
R10374 VSS.n5803 VSS.n2632 0.04025
R10375 VSS.n5804 VSS.n5803 0.04025
R10376 VSS.n5805 VSS.n5804 0.04025
R10377 VSS.n5805 VSS.n2630 0.04025
R10378 VSS.n5809 VSS.n2630 0.04025
R10379 VSS.n5810 VSS.n5809 0.04025
R10380 VSS.n5811 VSS.n5810 0.04025
R10381 VSS.n5811 VSS.n2628 0.04025
R10382 VSS.n5815 VSS.n2628 0.04025
R10383 VSS.n5816 VSS.n5815 0.04025
R10384 VSS.n5817 VSS.n5816 0.04025
R10385 VSS.n5817 VSS.n2626 0.04025
R10386 VSS.n5821 VSS.n2626 0.04025
R10387 VSS.n5822 VSS.n5821 0.04025
R10388 VSS.n5823 VSS.n5822 0.04025
R10389 VSS.n5823 VSS.n2624 0.04025
R10390 VSS.n5827 VSS.n2624 0.04025
R10391 VSS.n5828 VSS.n5827 0.04025
R10392 VSS.n5829 VSS.n5828 0.04025
R10393 VSS.n5829 VSS.n2622 0.04025
R10394 VSS.n5833 VSS.n2622 0.04025
R10395 VSS.n5834 VSS.n5833 0.04025
R10396 VSS.n5835 VSS.n5834 0.04025
R10397 VSS.n5835 VSS.n2620 0.04025
R10398 VSS.n5839 VSS.n2620 0.04025
R10399 VSS.n5840 VSS.n5839 0.04025
R10400 VSS.n5841 VSS.n5840 0.04025
R10401 VSS.n5841 VSS.n2618 0.04025
R10402 VSS.n5845 VSS.n2618 0.04025
R10403 VSS.n5846 VSS.n5845 0.04025
R10404 VSS.n5847 VSS.n5846 0.04025
R10405 VSS.n5847 VSS.n2616 0.04025
R10406 VSS.n5851 VSS.n2616 0.04025
R10407 VSS.n5852 VSS.n5851 0.04025
R10408 VSS.n5853 VSS.n5852 0.04025
R10409 VSS.n5853 VSS.n2614 0.04025
R10410 VSS.n5857 VSS.n2614 0.04025
R10411 VSS.n5858 VSS.n5857 0.04025
R10412 VSS.n5859 VSS.n5858 0.04025
R10413 VSS.n5859 VSS.n2612 0.04025
R10414 VSS.n5863 VSS.n2612 0.04025
R10415 VSS.n5864 VSS.n5863 0.04025
R10416 VSS.n5865 VSS.n5864 0.04025
R10417 VSS.n5865 VSS.n2610 0.04025
R10418 VSS.n5869 VSS.n2610 0.04025
R10419 VSS.n5870 VSS.n5869 0.04025
R10420 VSS.n5871 VSS.n5870 0.04025
R10421 VSS.n5871 VSS.n2608 0.04025
R10422 VSS.n5875 VSS.n2608 0.04025
R10423 VSS.n5876 VSS.n5875 0.04025
R10424 VSS.n5877 VSS.n5876 0.04025
R10425 VSS.n5877 VSS.n2606 0.04025
R10426 VSS.n5881 VSS.n2606 0.04025
R10427 VSS.n5882 VSS.n5881 0.04025
R10428 VSS.n5883 VSS.n5882 0.04025
R10429 VSS.n5883 VSS.n2604 0.04025
R10430 VSS.n5887 VSS.n2604 0.04025
R10431 VSS.n5888 VSS.n5887 0.04025
R10432 VSS.n5889 VSS.n5888 0.04025
R10433 VSS.n5889 VSS.n2602 0.04025
R10434 VSS.n5893 VSS.n2602 0.04025
R10435 VSS.n5894 VSS.n5893 0.04025
R10436 VSS.n5895 VSS.n5894 0.04025
R10437 VSS.n5895 VSS.n2600 0.04025
R10438 VSS.n5899 VSS.n2600 0.04025
R10439 VSS.n5900 VSS.n5899 0.04025
R10440 VSS.n5901 VSS.n5900 0.04025
R10441 VSS.n5901 VSS.n2598 0.04025
R10442 VSS.n5905 VSS.n2598 0.04025
R10443 VSS.n5906 VSS.n5905 0.04025
R10444 VSS.n5907 VSS.n5906 0.04025
R10445 VSS.n5907 VSS.n2596 0.04025
R10446 VSS.n5911 VSS.n2596 0.04025
R10447 VSS.n5912 VSS.n5911 0.04025
R10448 VSS.n5913 VSS.n5912 0.04025
R10449 VSS.n5913 VSS.n2594 0.04025
R10450 VSS.n5917 VSS.n2594 0.04025
R10451 VSS.n5918 VSS.n5917 0.04025
R10452 VSS.n5919 VSS.n5918 0.04025
R10453 VSS.n5919 VSS.n2592 0.04025
R10454 VSS.n5923 VSS.n2592 0.04025
R10455 VSS.n5924 VSS.n5923 0.04025
R10456 VSS.n5925 VSS.n5924 0.04025
R10457 VSS.n5925 VSS.n2590 0.04025
R10458 VSS.n5929 VSS.n2590 0.04025
R10459 VSS.n5930 VSS.n5929 0.04025
R10460 VSS.n5931 VSS.n5930 0.04025
R10461 VSS.n5931 VSS.n2588 0.04025
R10462 VSS.n5935 VSS.n2588 0.04025
R10463 VSS.n5936 VSS.n5935 0.04025
R10464 VSS.n5937 VSS.n5936 0.04025
R10465 VSS.n5937 VSS.n2586 0.04025
R10466 VSS.n5941 VSS.n2586 0.04025
R10467 VSS.n5942 VSS.n5941 0.04025
R10468 VSS.n5943 VSS.n5942 0.04025
R10469 VSS.n5943 VSS.n2584 0.04025
R10470 VSS.n5947 VSS.n2584 0.04025
R10471 VSS.n5948 VSS.n5947 0.04025
R10472 VSS.n5949 VSS.n5948 0.04025
R10473 VSS.n5949 VSS.n2582 0.04025
R10474 VSS.n5953 VSS.n2582 0.04025
R10475 VSS.n5954 VSS.n5953 0.04025
R10476 VSS.n5955 VSS.n5954 0.04025
R10477 VSS.n5955 VSS.n2580 0.04025
R10478 VSS.n5959 VSS.n2580 0.04025
R10479 VSS.n5960 VSS.n5959 0.04025
R10480 VSS.n5961 VSS.n5960 0.04025
R10481 VSS.n5961 VSS.n2578 0.04025
R10482 VSS.n5965 VSS.n2578 0.04025
R10483 VSS.n5966 VSS.n5965 0.04025
R10484 VSS.n5967 VSS.n5966 0.04025
R10485 VSS.n5967 VSS.n2576 0.04025
R10486 VSS.n5971 VSS.n2576 0.04025
R10487 VSS.n5972 VSS.n5971 0.04025
R10488 VSS.n5973 VSS.n5972 0.04025
R10489 VSS.n5973 VSS.n2574 0.04025
R10490 VSS.n5977 VSS.n2574 0.04025
R10491 VSS.n5978 VSS.n5977 0.04025
R10492 VSS.n5979 VSS.n5978 0.04025
R10493 VSS.n5979 VSS.n2572 0.04025
R10494 VSS.n5983 VSS.n2572 0.04025
R10495 VSS.n5984 VSS.n5983 0.04025
R10496 VSS.n5985 VSS.n5984 0.04025
R10497 VSS.n5985 VSS.n2570 0.04025
R10498 VSS.n5989 VSS.n2570 0.04025
R10499 VSS.n5990 VSS.n5989 0.04025
R10500 VSS.n5991 VSS.n5990 0.04025
R10501 VSS.n5991 VSS.n2568 0.04025
R10502 VSS.n5995 VSS.n2568 0.04025
R10503 VSS.n5996 VSS.n5995 0.04025
R10504 VSS.n5997 VSS.n5996 0.04025
R10505 VSS.n5997 VSS.n2566 0.04025
R10506 VSS.n6001 VSS.n2566 0.04025
R10507 VSS.n6002 VSS.n6001 0.04025
R10508 VSS.n6003 VSS.n6002 0.04025
R10509 VSS.n6003 VSS.n2564 0.04025
R10510 VSS.n6007 VSS.n2564 0.04025
R10511 VSS.n6008 VSS.n6007 0.04025
R10512 VSS.n6009 VSS.n6008 0.04025
R10513 VSS.n6009 VSS.n2562 0.04025
R10514 VSS.n6013 VSS.n2562 0.04025
R10515 VSS.n6014 VSS.n6013 0.04025
R10516 VSS.n6015 VSS.n6014 0.04025
R10517 VSS.n6015 VSS.n2560 0.04025
R10518 VSS.n6019 VSS.n2560 0.04025
R10519 VSS.n6020 VSS.n6019 0.04025
R10520 VSS.n6021 VSS.n6020 0.04025
R10521 VSS.n6021 VSS.n2558 0.04025
R10522 VSS.n6025 VSS.n2558 0.04025
R10523 VSS.n6026 VSS.n6025 0.04025
R10524 VSS.n6027 VSS.n6026 0.04025
R10525 VSS.n6027 VSS.n2556 0.04025
R10526 VSS.n6031 VSS.n2556 0.04025
R10527 VSS.n6032 VSS.n6031 0.04025
R10528 VSS.n6033 VSS.n6032 0.04025
R10529 VSS.n6033 VSS.n2554 0.04025
R10530 VSS.n6037 VSS.n2554 0.04025
R10531 VSS.n6038 VSS.n6037 0.04025
R10532 VSS.n6039 VSS.n6038 0.04025
R10533 VSS.n6039 VSS.n2552 0.04025
R10534 VSS.n6043 VSS.n2552 0.04025
R10535 VSS.n6044 VSS.n6043 0.04025
R10536 VSS.n6045 VSS.n6044 0.04025
R10537 VSS.n6045 VSS.n2550 0.04025
R10538 VSS.n6049 VSS.n2550 0.04025
R10539 VSS.n6050 VSS.n6049 0.04025
R10540 VSS.n6051 VSS.n6050 0.04025
R10541 VSS.n6051 VSS.n2548 0.04025
R10542 VSS.n6055 VSS.n2548 0.04025
R10543 VSS.n6056 VSS.n6055 0.04025
R10544 VSS.n6057 VSS.n6056 0.04025
R10545 VSS.n6057 VSS.n2546 0.04025
R10546 VSS.n6061 VSS.n2546 0.04025
R10547 VSS.n6062 VSS.n6061 0.04025
R10548 VSS.n6063 VSS.n6062 0.04025
R10549 VSS.n6063 VSS.n2544 0.04025
R10550 VSS.n6067 VSS.n2544 0.04025
R10551 VSS.n6068 VSS.n6067 0.04025
R10552 VSS.n6069 VSS.n6068 0.04025
R10553 VSS.n6069 VSS.n2542 0.04025
R10554 VSS.n6073 VSS.n2542 0.04025
R10555 VSS.n6074 VSS.n6073 0.04025
R10556 VSS.n6075 VSS.n6074 0.04025
R10557 VSS.n6075 VSS.n2540 0.04025
R10558 VSS.n6079 VSS.n2540 0.04025
R10559 VSS.n6080 VSS.n6079 0.04025
R10560 VSS.n6081 VSS.n6080 0.04025
R10561 VSS.n6081 VSS.n2538 0.04025
R10562 VSS.n6085 VSS.n2538 0.04025
R10563 VSS.n6086 VSS.n6085 0.04025
R10564 VSS.n6087 VSS.n6086 0.04025
R10565 VSS.n6087 VSS.n2536 0.04025
R10566 VSS.n6091 VSS.n2536 0.04025
R10567 VSS.n6092 VSS.n6091 0.04025
R10568 VSS.n6093 VSS.n6092 0.04025
R10569 VSS.n6093 VSS.n2534 0.04025
R10570 VSS.n6097 VSS.n2534 0.04025
R10571 VSS.n6098 VSS.n6097 0.04025
R10572 VSS.n6099 VSS.n6098 0.04025
R10573 VSS.n6099 VSS.n2532 0.04025
R10574 VSS.n6103 VSS.n2532 0.04025
R10575 VSS.n6104 VSS.n6103 0.04025
R10576 VSS.n6105 VSS.n6104 0.04025
R10577 VSS.n6105 VSS.n2530 0.04025
R10578 VSS.n6109 VSS.n2530 0.04025
R10579 VSS.n6110 VSS.n6109 0.04025
R10580 VSS.n6111 VSS.n6110 0.04025
R10581 VSS.n6111 VSS.n2528 0.04025
R10582 VSS.n6115 VSS.n2528 0.04025
R10583 VSS.n6116 VSS.n6115 0.04025
R10584 VSS.n6117 VSS.n6116 0.04025
R10585 VSS.n6117 VSS.n2526 0.04025
R10586 VSS.n6121 VSS.n2526 0.04025
R10587 VSS.n6122 VSS.n6121 0.04025
R10588 VSS.n6123 VSS.n6122 0.04025
R10589 VSS.n6123 VSS.n2524 0.04025
R10590 VSS.n6127 VSS.n2524 0.04025
R10591 VSS.n6128 VSS.n6127 0.04025
R10592 VSS.n6129 VSS.n6128 0.04025
R10593 VSS.n6129 VSS.n2522 0.04025
R10594 VSS.n6133 VSS.n2522 0.04025
R10595 VSS.n6134 VSS.n6133 0.04025
R10596 VSS.n6135 VSS.n6134 0.04025
R10597 VSS.n6135 VSS.n2520 0.04025
R10598 VSS.n6139 VSS.n2520 0.04025
R10599 VSS.n6140 VSS.n6139 0.04025
R10600 VSS.n6141 VSS.n6140 0.04025
R10601 VSS.n6141 VSS.n2518 0.04025
R10602 VSS.n6145 VSS.n2518 0.04025
R10603 VSS.n6146 VSS.n6145 0.04025
R10604 VSS.n6147 VSS.n6146 0.04025
R10605 VSS.n6147 VSS.n2516 0.04025
R10606 VSS.n6151 VSS.n2516 0.04025
R10607 VSS.n6152 VSS.n6151 0.04025
R10608 VSS.n6153 VSS.n6152 0.04025
R10609 VSS.n6153 VSS.n2514 0.04025
R10610 VSS.n6157 VSS.n2514 0.04025
R10611 VSS.n6158 VSS.n6157 0.04025
R10612 VSS.n6159 VSS.n6158 0.04025
R10613 VSS.n6159 VSS.n2512 0.04025
R10614 VSS.n6163 VSS.n2512 0.04025
R10615 VSS.n6164 VSS.n6163 0.04025
R10616 VSS.n6165 VSS.n6164 0.04025
R10617 VSS.n6165 VSS.n2510 0.04025
R10618 VSS.n6169 VSS.n2510 0.04025
R10619 VSS.n6170 VSS.n6169 0.04025
R10620 VSS.n6171 VSS.n6170 0.04025
R10621 VSS.n6171 VSS.n2508 0.04025
R10622 VSS.n6175 VSS.n2508 0.04025
R10623 VSS.n6176 VSS.n6175 0.04025
R10624 VSS.n6177 VSS.n6176 0.04025
R10625 VSS.n6177 VSS.n2506 0.04025
R10626 VSS.n6181 VSS.n2506 0.04025
R10627 VSS.n6182 VSS.n6181 0.04025
R10628 VSS.n6183 VSS.n6182 0.04025
R10629 VSS.n6183 VSS.n2504 0.04025
R10630 VSS.n6187 VSS.n2504 0.04025
R10631 VSS.n6188 VSS.n6187 0.04025
R10632 VSS.n6189 VSS.n6188 0.04025
R10633 VSS.n6189 VSS.n2502 0.04025
R10634 VSS.n6193 VSS.n2502 0.04025
R10635 VSS.n6194 VSS.n6193 0.04025
R10636 VSS.n6195 VSS.n6194 0.04025
R10637 VSS.n6195 VSS.n2500 0.04025
R10638 VSS.n6199 VSS.n2500 0.04025
R10639 VSS.n6200 VSS.n6199 0.04025
R10640 VSS.n6201 VSS.n6200 0.04025
R10641 VSS.n6201 VSS.n2498 0.04025
R10642 VSS.n6205 VSS.n2498 0.04025
R10643 VSS.n6206 VSS.n6205 0.04025
R10644 VSS.n6207 VSS.n6206 0.04025
R10645 VSS.n6207 VSS.n2496 0.04025
R10646 VSS.n6211 VSS.n2496 0.04025
R10647 VSS.n6212 VSS.n6211 0.04025
R10648 VSS.n6213 VSS.n6212 0.04025
R10649 VSS.n6213 VSS.n2494 0.04025
R10650 VSS.n6217 VSS.n2494 0.04025
R10651 VSS.n6218 VSS.n6217 0.04025
R10652 VSS.n6219 VSS.n6218 0.04025
R10653 VSS.n6219 VSS.n2492 0.04025
R10654 VSS.n6223 VSS.n2492 0.04025
R10655 VSS.n6224 VSS.n6223 0.04025
R10656 VSS.n6225 VSS.n6224 0.04025
R10657 VSS.n6225 VSS.n2490 0.04025
R10658 VSS.n6229 VSS.n2490 0.04025
R10659 VSS.n6230 VSS.n6229 0.04025
R10660 VSS.n6231 VSS.n6230 0.04025
R10661 VSS.n6231 VSS.n2488 0.04025
R10662 VSS.n6235 VSS.n2488 0.04025
R10663 VSS.n6236 VSS.n6235 0.04025
R10664 VSS.n6237 VSS.n6236 0.04025
R10665 VSS.n6237 VSS.n2486 0.04025
R10666 VSS.n6241 VSS.n2486 0.04025
R10667 VSS.n6242 VSS.n6241 0.04025
R10668 VSS.n6243 VSS.n6242 0.04025
R10669 VSS.n6243 VSS.n2484 0.04025
R10670 VSS.n6247 VSS.n2484 0.04025
R10671 VSS.n6248 VSS.n6247 0.04025
R10672 VSS.n6249 VSS.n6248 0.04025
R10673 VSS.n6249 VSS.n2482 0.04025
R10674 VSS.n6253 VSS.n2482 0.04025
R10675 VSS.n6254 VSS.n6253 0.04025
R10676 VSS.n6255 VSS.n6254 0.04025
R10677 VSS.n6255 VSS.n2480 0.04025
R10678 VSS.n6259 VSS.n2480 0.04025
R10679 VSS.n6260 VSS.n6259 0.04025
R10680 VSS.n6261 VSS.n6260 0.04025
R10681 VSS.n6261 VSS.n2478 0.04025
R10682 VSS.n6265 VSS.n2478 0.04025
R10683 VSS.n6266 VSS.n6265 0.04025
R10684 VSS.n6267 VSS.n6266 0.04025
R10685 VSS.n6267 VSS.n2476 0.04025
R10686 VSS.n6271 VSS.n2476 0.04025
R10687 VSS.n6272 VSS.n6271 0.04025
R10688 VSS.n6273 VSS.n6272 0.04025
R10689 VSS.n6273 VSS.n2474 0.04025
R10690 VSS.n6277 VSS.n2474 0.04025
R10691 VSS.n6278 VSS.n6277 0.04025
R10692 VSS.n6279 VSS.n6278 0.04025
R10693 VSS.n6279 VSS.n2472 0.04025
R10694 VSS.n6283 VSS.n2472 0.04025
R10695 VSS.n6284 VSS.n6283 0.04025
R10696 VSS.n6285 VSS.n6284 0.04025
R10697 VSS.n6285 VSS.n2470 0.04025
R10698 VSS.n6289 VSS.n2470 0.04025
R10699 VSS.n6290 VSS.n6289 0.04025
R10700 VSS.n6291 VSS.n6290 0.04025
R10701 VSS.n6291 VSS.n2468 0.04025
R10702 VSS.n6295 VSS.n2468 0.04025
R10703 VSS.n6296 VSS.n6295 0.04025
R10704 VSS.n6297 VSS.n6296 0.04025
R10705 VSS.n6297 VSS.n2466 0.04025
R10706 VSS.n6301 VSS.n2466 0.04025
R10707 VSS.n6302 VSS.n6301 0.04025
R10708 VSS.n6303 VSS.n6302 0.04025
R10709 VSS.n6303 VSS.n2464 0.04025
R10710 VSS.n6307 VSS.n2464 0.04025
R10711 VSS.n6308 VSS.n6307 0.04025
R10712 VSS.n6309 VSS.n6308 0.04025
R10713 VSS.n6309 VSS.n2462 0.04025
R10714 VSS.n6313 VSS.n2462 0.04025
R10715 VSS.n6314 VSS.n6313 0.04025
R10716 VSS.n6315 VSS.n6314 0.04025
R10717 VSS.n6315 VSS.n2460 0.04025
R10718 VSS.n6319 VSS.n2460 0.04025
R10719 VSS.n6320 VSS.n6319 0.04025
R10720 VSS.n6321 VSS.n6320 0.04025
R10721 VSS.n6321 VSS.n2458 0.04025
R10722 VSS.n6325 VSS.n2458 0.04025
R10723 VSS.n6326 VSS.n6325 0.04025
R10724 VSS.n6327 VSS.n6326 0.04025
R10725 VSS.n6327 VSS.n2456 0.04025
R10726 VSS.n6331 VSS.n2456 0.04025
R10727 VSS.n6332 VSS.n6331 0.04025
R10728 VSS.n6333 VSS.n6332 0.04025
R10729 VSS.n6333 VSS.n2454 0.04025
R10730 VSS.n6337 VSS.n2454 0.04025
R10731 VSS.n6338 VSS.n6337 0.04025
R10732 VSS.n6339 VSS.n6338 0.04025
R10733 VSS.n6339 VSS.n2452 0.04025
R10734 VSS.n6343 VSS.n2452 0.04025
R10735 VSS.n6344 VSS.n6343 0.04025
R10736 VSS.n6345 VSS.n6344 0.04025
R10737 VSS.n6345 VSS.n2450 0.04025
R10738 VSS.n6349 VSS.n2450 0.04025
R10739 VSS.n6350 VSS.n6349 0.04025
R10740 VSS.n6351 VSS.n6350 0.04025
R10741 VSS.n6351 VSS.n2448 0.04025
R10742 VSS.n6355 VSS.n2448 0.04025
R10743 VSS.n6356 VSS.n6355 0.04025
R10744 VSS.n6357 VSS.n6356 0.04025
R10745 VSS.n6357 VSS.n2446 0.04025
R10746 VSS.n6361 VSS.n2446 0.04025
R10747 VSS.n6362 VSS.n6361 0.04025
R10748 VSS.n6363 VSS.n6362 0.04025
R10749 VSS.n6363 VSS.n2444 0.04025
R10750 VSS.n6367 VSS.n2444 0.04025
R10751 VSS.n6368 VSS.n6367 0.04025
R10752 VSS.n6369 VSS.n6368 0.04025
R10753 VSS.n6369 VSS.n2442 0.04025
R10754 VSS.n6373 VSS.n2442 0.04025
R10755 VSS.n6374 VSS.n6373 0.04025
R10756 VSS.n6375 VSS.n6374 0.04025
R10757 VSS.n6375 VSS.n2440 0.04025
R10758 VSS.n6379 VSS.n2440 0.04025
R10759 VSS.n6380 VSS.n6379 0.04025
R10760 VSS.n6381 VSS.n6380 0.04025
R10761 VSS.n6381 VSS.n2438 0.04025
R10762 VSS.n6385 VSS.n2438 0.04025
R10763 VSS.n6386 VSS.n6385 0.04025
R10764 VSS.n6387 VSS.n6386 0.04025
R10765 VSS.n6387 VSS.n2436 0.04025
R10766 VSS.n6391 VSS.n2436 0.04025
R10767 VSS.n6392 VSS.n6391 0.04025
R10768 VSS.n6393 VSS.n6392 0.04025
R10769 VSS.n6393 VSS.n2434 0.04025
R10770 VSS.n6397 VSS.n2434 0.04025
R10771 VSS.n6398 VSS.n6397 0.04025
R10772 VSS.n6399 VSS.n6398 0.04025
R10773 VSS.n6399 VSS.n2432 0.04025
R10774 VSS.n6403 VSS.n2432 0.04025
R10775 VSS.n6404 VSS.n6403 0.04025
R10776 VSS.n6405 VSS.n6404 0.04025
R10777 VSS.n6405 VSS.n2430 0.04025
R10778 VSS.n6409 VSS.n2430 0.04025
R10779 VSS.n6410 VSS.n6409 0.04025
R10780 VSS.n6411 VSS.n6410 0.04025
R10781 VSS.n6411 VSS.n2428 0.04025
R10782 VSS.n6415 VSS.n2428 0.04025
R10783 VSS.n6416 VSS.n6415 0.04025
R10784 VSS.n6417 VSS.n6416 0.04025
R10785 VSS.n6417 VSS.n2426 0.04025
R10786 VSS.n6421 VSS.n2426 0.04025
R10787 VSS.n6422 VSS.n6421 0.04025
R10788 VSS.n6423 VSS.n6422 0.04025
R10789 VSS.n6423 VSS.n2424 0.04025
R10790 VSS.n6427 VSS.n2424 0.04025
R10791 VSS.n6428 VSS.n6427 0.04025
R10792 VSS.n6429 VSS.n6428 0.04025
R10793 VSS.n6429 VSS.n2422 0.04025
R10794 VSS.n6433 VSS.n2422 0.04025
R10795 VSS.n6434 VSS.n6433 0.04025
R10796 VSS.n6435 VSS.n6434 0.04025
R10797 VSS.n6435 VSS.n2420 0.04025
R10798 VSS.n6439 VSS.n2420 0.04025
R10799 VSS.n6440 VSS.n6439 0.04025
R10800 VSS.n6441 VSS.n6440 0.04025
R10801 VSS.n6441 VSS.n2418 0.04025
R10802 VSS.n6445 VSS.n2418 0.04025
R10803 VSS.n6446 VSS.n6445 0.04025
R10804 VSS.n6447 VSS.n6446 0.04025
R10805 VSS.n6447 VSS.n2416 0.04025
R10806 VSS.n6451 VSS.n2416 0.04025
R10807 VSS.n6452 VSS.n6451 0.04025
R10808 VSS.n6453 VSS.n6452 0.04025
R10809 VSS.n6453 VSS.n2414 0.04025
R10810 VSS.n6457 VSS.n2414 0.04025
R10811 VSS.n6458 VSS.n6457 0.04025
R10812 VSS.n6459 VSS.n6458 0.04025
R10813 VSS.n6459 VSS.n2412 0.04025
R10814 VSS.n6463 VSS.n2412 0.04025
R10815 VSS.n6464 VSS.n6463 0.04025
R10816 VSS.n6465 VSS.n6464 0.04025
R10817 VSS.n6465 VSS.n2410 0.04025
R10818 VSS.n6469 VSS.n2410 0.04025
R10819 VSS.n6470 VSS.n6469 0.04025
R10820 VSS.n6471 VSS.n6470 0.04025
R10821 VSS.n6471 VSS.n2408 0.04025
R10822 VSS.n6475 VSS.n2408 0.04025
R10823 VSS.n6476 VSS.n6475 0.04025
R10824 VSS.n6477 VSS.n6476 0.04025
R10825 VSS.n6477 VSS.n2406 0.04025
R10826 VSS.n6481 VSS.n2406 0.04025
R10827 VSS.n6482 VSS.n6481 0.04025
R10828 VSS.n6483 VSS.n6482 0.04025
R10829 VSS.n6483 VSS.n2404 0.04025
R10830 VSS.n6487 VSS.n2404 0.04025
R10831 VSS.n6488 VSS.n6487 0.04025
R10832 VSS.n6489 VSS.n6488 0.04025
R10833 VSS.n6489 VSS.n2402 0.04025
R10834 VSS.n6493 VSS.n2402 0.04025
R10835 VSS.n6494 VSS.n6493 0.04025
R10836 VSS.n6495 VSS.n6494 0.04025
R10837 VSS.n6495 VSS.n2400 0.04025
R10838 VSS.n6499 VSS.n2400 0.04025
R10839 VSS.n6500 VSS.n6499 0.04025
R10840 VSS.n6501 VSS.n6500 0.04025
R10841 VSS.n6501 VSS.n2398 0.04025
R10842 VSS.n6505 VSS.n2398 0.04025
R10843 VSS.n6506 VSS.n6505 0.04025
R10844 VSS.n6507 VSS.n6506 0.04025
R10845 VSS.n6507 VSS.n2396 0.04025
R10846 VSS.n6511 VSS.n2396 0.04025
R10847 VSS.n6512 VSS.n6511 0.04025
R10848 VSS.n6513 VSS.n6512 0.04025
R10849 VSS.n6513 VSS.n2394 0.04025
R10850 VSS.n6517 VSS.n2394 0.04025
R10851 VSS.n6518 VSS.n6517 0.04025
R10852 VSS.n6519 VSS.n6518 0.04025
R10853 VSS.n6519 VSS.n2392 0.04025
R10854 VSS.n6523 VSS.n2392 0.04025
R10855 VSS.n6524 VSS.n6523 0.04025
R10856 VSS.n6525 VSS.n6524 0.04025
R10857 VSS.n6525 VSS.n2390 0.04025
R10858 VSS.n6529 VSS.n2390 0.04025
R10859 VSS.n6530 VSS.n6529 0.04025
R10860 VSS.n6531 VSS.n6530 0.04025
R10861 VSS.n6531 VSS.n2388 0.04025
R10862 VSS.n6535 VSS.n2388 0.04025
R10863 VSS.n6536 VSS.n6535 0.04025
R10864 VSS.n6537 VSS.n6536 0.04025
R10865 VSS.n6537 VSS.n2386 0.04025
R10866 VSS.n6541 VSS.n2386 0.04025
R10867 VSS.n6542 VSS.n6541 0.04025
R10868 VSS.n6543 VSS.n6542 0.04025
R10869 VSS.n6543 VSS.n2384 0.04025
R10870 VSS.n6547 VSS.n2384 0.04025
R10871 VSS.n6548 VSS.n6547 0.04025
R10872 VSS.n6549 VSS.n6548 0.04025
R10873 VSS.n6549 VSS.n2382 0.04025
R10874 VSS.n6553 VSS.n2382 0.04025
R10875 VSS.n6554 VSS.n6553 0.04025
R10876 VSS.n6555 VSS.n6554 0.04025
R10877 VSS.n6555 VSS.n2380 0.04025
R10878 VSS.n6559 VSS.n2380 0.04025
R10879 VSS.n6560 VSS.n6559 0.04025
R10880 VSS.n6561 VSS.n6560 0.04025
R10881 VSS.n6561 VSS.n2378 0.04025
R10882 VSS.n6565 VSS.n2378 0.04025
R10883 VSS.n6566 VSS.n6565 0.04025
R10884 VSS.n6567 VSS.n6566 0.04025
R10885 VSS.n6567 VSS.n2376 0.04025
R10886 VSS.n6571 VSS.n2376 0.04025
R10887 VSS.n6572 VSS.n6571 0.04025
R10888 VSS.n6573 VSS.n6572 0.04025
R10889 VSS.n6573 VSS.n2374 0.04025
R10890 VSS.n6577 VSS.n2374 0.04025
R10891 VSS.n6578 VSS.n6577 0.04025
R10892 VSS.n6579 VSS.n6578 0.04025
R10893 VSS.n6579 VSS.n2372 0.04025
R10894 VSS.n6583 VSS.n2372 0.04025
R10895 VSS.n6584 VSS.n6583 0.04025
R10896 VSS.n6585 VSS.n6584 0.04025
R10897 VSS.n6585 VSS.n2370 0.04025
R10898 VSS.n6589 VSS.n2370 0.04025
R10899 VSS.n6590 VSS.n6589 0.04025
R10900 VSS.n6591 VSS.n6590 0.04025
R10901 VSS.n6591 VSS.n2368 0.04025
R10902 VSS.n6595 VSS.n2368 0.04025
R10903 VSS.n6596 VSS.n6595 0.04025
R10904 VSS.n6597 VSS.n6596 0.04025
R10905 VSS.n6597 VSS.n2366 0.04025
R10906 VSS.n6601 VSS.n2366 0.04025
R10907 VSS.n6602 VSS.n6601 0.04025
R10908 VSS.n6603 VSS.n6602 0.04025
R10909 VSS.n6603 VSS.n2364 0.04025
R10910 VSS.n6607 VSS.n2364 0.04025
R10911 VSS.n6608 VSS.n6607 0.04025
R10912 VSS.n6609 VSS.n6608 0.04025
R10913 VSS.n6609 VSS.n2362 0.04025
R10914 VSS.n6613 VSS.n2362 0.04025
R10915 VSS.n6614 VSS.n6613 0.04025
R10916 VSS.n6615 VSS.n6614 0.04025
R10917 VSS.n6615 VSS.n2360 0.04025
R10918 VSS.n6619 VSS.n2360 0.04025
R10919 VSS.n6620 VSS.n6619 0.04025
R10920 VSS.n6621 VSS.n6620 0.04025
R10921 VSS.n6621 VSS.n2358 0.04025
R10922 VSS.n6625 VSS.n2358 0.04025
R10923 VSS.n6626 VSS.n6625 0.04025
R10924 VSS.n6627 VSS.n6626 0.04025
R10925 VSS.n6627 VSS.n2356 0.04025
R10926 VSS.n6631 VSS.n2356 0.04025
R10927 VSS.n6632 VSS.n6631 0.04025
R10928 VSS.n6633 VSS.n6632 0.04025
R10929 VSS.n6633 VSS.n2354 0.04025
R10930 VSS.n6637 VSS.n2354 0.04025
R10931 VSS.n6638 VSS.n6637 0.04025
R10932 VSS.n6639 VSS.n6638 0.04025
R10933 VSS.n6639 VSS.n2352 0.04025
R10934 VSS.n6643 VSS.n2352 0.04025
R10935 VSS.n6644 VSS.n6643 0.04025
R10936 VSS.n6645 VSS.n6644 0.04025
R10937 VSS.n6645 VSS.n2350 0.04025
R10938 VSS.n6649 VSS.n2350 0.04025
R10939 VSS.n6650 VSS.n6649 0.04025
R10940 VSS.n6651 VSS.n6650 0.04025
R10941 VSS.n6651 VSS.n2348 0.04025
R10942 VSS.n6655 VSS.n2348 0.04025
R10943 VSS.n6656 VSS.n6655 0.04025
R10944 VSS.n6657 VSS.n6656 0.04025
R10945 VSS.n6657 VSS.n2346 0.04025
R10946 VSS.n6661 VSS.n2346 0.04025
R10947 VSS.n6662 VSS.n6661 0.04025
R10948 VSS.n6663 VSS.n6662 0.04025
R10949 VSS.n6663 VSS.n2344 0.04025
R10950 VSS.n6667 VSS.n2344 0.04025
R10951 VSS.n6668 VSS.n6667 0.04025
R10952 VSS.n6669 VSS.n6668 0.04025
R10953 VSS.n6669 VSS.n2342 0.04025
R10954 VSS.n6673 VSS.n2342 0.04025
R10955 VSS.n6674 VSS.n6673 0.04025
R10956 VSS.n6675 VSS.n6674 0.04025
R10957 VSS.n6675 VSS.n2340 0.04025
R10958 VSS.n6679 VSS.n2340 0.04025
R10959 VSS.n6680 VSS.n6679 0.04025
R10960 VSS.n6681 VSS.n6680 0.04025
R10961 VSS.n6681 VSS.n2338 0.04025
R10962 VSS.n6685 VSS.n2338 0.04025
R10963 VSS.n6686 VSS.n6685 0.04025
R10964 VSS.n6687 VSS.n6686 0.04025
R10965 VSS.n6687 VSS.n2336 0.04025
R10966 VSS.n6691 VSS.n2336 0.04025
R10967 VSS.n6692 VSS.n6691 0.04025
R10968 VSS.n6693 VSS.n6692 0.04025
R10969 VSS.n6693 VSS.n2334 0.04025
R10970 VSS.n6697 VSS.n2334 0.04025
R10971 VSS.n6698 VSS.n6697 0.04025
R10972 VSS.n6699 VSS.n6698 0.04025
R10973 VSS.n6699 VSS.n2332 0.04025
R10974 VSS.n6703 VSS.n2332 0.04025
R10975 VSS.n6704 VSS.n6703 0.04025
R10976 VSS.n6705 VSS.n6704 0.04025
R10977 VSS.n6705 VSS.n2330 0.04025
R10978 VSS.n6709 VSS.n2330 0.04025
R10979 VSS.n6710 VSS.n6709 0.04025
R10980 VSS.n6711 VSS.n6710 0.04025
R10981 VSS.n6711 VSS.n2328 0.04025
R10982 VSS.n6715 VSS.n2328 0.04025
R10983 VSS.n6716 VSS.n6715 0.04025
R10984 VSS.n6717 VSS.n6716 0.04025
R10985 VSS.n6717 VSS.n2326 0.04025
R10986 VSS.n6721 VSS.n2326 0.04025
R10987 VSS.n6722 VSS.n6721 0.04025
R10988 VSS.n6723 VSS.n6722 0.04025
R10989 VSS.n6723 VSS.n2324 0.04025
R10990 VSS.n6727 VSS.n2324 0.04025
R10991 VSS.n6728 VSS.n6727 0.04025
R10992 VSS.n6729 VSS.n6728 0.04025
R10993 VSS.n6729 VSS.n2322 0.04025
R10994 VSS.n6733 VSS.n2322 0.04025
R10995 VSS.n6734 VSS.n6733 0.04025
R10996 VSS.n6735 VSS.n6734 0.04025
R10997 VSS.n6735 VSS.n2320 0.04025
R10998 VSS.n6739 VSS.n2320 0.04025
R10999 VSS.n6740 VSS.n6739 0.04025
R11000 VSS.n6741 VSS.n6740 0.04025
R11001 VSS.n6741 VSS.n2318 0.04025
R11002 VSS.n6745 VSS.n2318 0.04025
R11003 VSS.n6746 VSS.n6745 0.04025
R11004 VSS.n6747 VSS.n6746 0.04025
R11005 VSS.n6747 VSS.n2316 0.04025
R11006 VSS.n6751 VSS.n2316 0.04025
R11007 VSS.n6752 VSS.n6751 0.04025
R11008 VSS.n6753 VSS.n6752 0.04025
R11009 VSS.n6753 VSS.n2314 0.04025
R11010 VSS.n6757 VSS.n2314 0.04025
R11011 VSS.n6758 VSS.n6757 0.04025
R11012 VSS.n6759 VSS.n6758 0.04025
R11013 VSS.n6759 VSS.n2312 0.04025
R11014 VSS.n6763 VSS.n2312 0.04025
R11015 VSS.n6764 VSS.n6763 0.04025
R11016 VSS.n6765 VSS.n6764 0.04025
R11017 VSS.n6765 VSS.n2310 0.04025
R11018 VSS.n6769 VSS.n2310 0.04025
R11019 VSS.n6770 VSS.n6769 0.04025
R11020 VSS.n6771 VSS.n6770 0.04025
R11021 VSS.n6771 VSS.n2308 0.04025
R11022 VSS.n6775 VSS.n2308 0.04025
R11023 VSS.n6776 VSS.n6775 0.04025
R11024 VSS.n6777 VSS.n6776 0.04025
R11025 VSS.n6777 VSS.n2306 0.04025
R11026 VSS.n6781 VSS.n2306 0.04025
R11027 VSS.n6782 VSS.n6781 0.04025
R11028 VSS.n6783 VSS.n6782 0.04025
R11029 VSS.n6783 VSS.n2304 0.04025
R11030 VSS.n6787 VSS.n2304 0.04025
R11031 VSS.n6788 VSS.n6787 0.04025
R11032 VSS.n6789 VSS.n6788 0.04025
R11033 VSS.n6789 VSS.n2302 0.04025
R11034 VSS.n6793 VSS.n2302 0.04025
R11035 VSS.n6794 VSS.n6793 0.04025
R11036 VSS.n6795 VSS.n6794 0.04025
R11037 VSS.n6795 VSS.n2300 0.04025
R11038 VSS.n6799 VSS.n2300 0.04025
R11039 VSS.n6800 VSS.n6799 0.04025
R11040 VSS.n6801 VSS.n6800 0.04025
R11041 VSS.n6801 VSS.n2298 0.04025
R11042 VSS.n6805 VSS.n2298 0.04025
R11043 VSS.n6806 VSS.n6805 0.04025
R11044 VSS.n6807 VSS.n6806 0.04025
R11045 VSS.n6807 VSS.n2296 0.04025
R11046 VSS.n6811 VSS.n2296 0.04025
R11047 VSS.n6812 VSS.n6811 0.04025
R11048 VSS.n6813 VSS.n6812 0.04025
R11049 VSS.n6813 VSS.n2294 0.04025
R11050 VSS.n6817 VSS.n2294 0.04025
R11051 VSS.n6818 VSS.n6817 0.04025
R11052 VSS.n6819 VSS.n6818 0.04025
R11053 VSS.n6819 VSS.n2292 0.04025
R11054 VSS.n6823 VSS.n2292 0.04025
R11055 VSS.n6824 VSS.n6823 0.04025
R11056 VSS.n6825 VSS.n6824 0.04025
R11057 VSS.n6825 VSS.n2290 0.04025
R11058 VSS.n6829 VSS.n2290 0.04025
R11059 VSS.n6830 VSS.n6829 0.04025
R11060 VSS.n6831 VSS.n6830 0.04025
R11061 VSS.n6831 VSS.n2288 0.04025
R11062 VSS.n6835 VSS.n2288 0.04025
R11063 VSS.n6836 VSS.n6835 0.04025
R11064 VSS.n6837 VSS.n6836 0.04025
R11065 VSS.n6837 VSS.n2286 0.04025
R11066 VSS.n6841 VSS.n2286 0.04025
R11067 VSS.n6842 VSS.n6841 0.04025
R11068 VSS.n6843 VSS.n6842 0.04025
R11069 VSS.n6843 VSS.n2284 0.04025
R11070 VSS.n6847 VSS.n2284 0.04025
R11071 VSS.n6848 VSS.n6847 0.04025
R11072 VSS.n6849 VSS.n6848 0.04025
R11073 VSS.n6849 VSS.n2282 0.04025
R11074 VSS.n6853 VSS.n2282 0.04025
R11075 VSS.n6854 VSS.n6853 0.04025
R11076 VSS.n6855 VSS.n6854 0.04025
R11077 VSS.n6855 VSS.n2280 0.04025
R11078 VSS.n6859 VSS.n2280 0.04025
R11079 VSS.n6860 VSS.n6859 0.04025
R11080 VSS.n6861 VSS.n6860 0.04025
R11081 VSS.n6861 VSS.n2278 0.04025
R11082 VSS.n6865 VSS.n2278 0.04025
R11083 VSS.n6866 VSS.n6865 0.04025
R11084 VSS.n6867 VSS.n6866 0.04025
R11085 VSS.n6867 VSS.n2276 0.04025
R11086 VSS.n6871 VSS.n2276 0.04025
R11087 VSS.n6872 VSS.n6871 0.04025
R11088 VSS.n6873 VSS.n6872 0.04025
R11089 VSS.n6873 VSS.n2274 0.04025
R11090 VSS.n6877 VSS.n2274 0.04025
R11091 VSS.n6878 VSS.n6877 0.04025
R11092 VSS.n6879 VSS.n6878 0.04025
R11093 VSS.n6879 VSS.n2272 0.04025
R11094 VSS.n6883 VSS.n2272 0.04025
R11095 VSS.n6884 VSS.n6883 0.04025
R11096 VSS.n6885 VSS.n6884 0.04025
R11097 VSS.n6885 VSS.n2270 0.04025
R11098 VSS.n6889 VSS.n2270 0.04025
R11099 VSS.n6890 VSS.n6889 0.04025
R11100 VSS.n6891 VSS.n6890 0.04025
R11101 VSS.n6891 VSS.n2268 0.04025
R11102 VSS.n6895 VSS.n2268 0.04025
R11103 VSS.n6896 VSS.n6895 0.04025
R11104 VSS.n6897 VSS.n6896 0.04025
R11105 VSS.n6897 VSS.n2266 0.04025
R11106 VSS.n6901 VSS.n2266 0.04025
R11107 VSS.n6902 VSS.n6901 0.04025
R11108 VSS.n6903 VSS.n6902 0.04025
R11109 VSS.n6903 VSS.n2264 0.04025
R11110 VSS.n6907 VSS.n2264 0.04025
R11111 VSS.n8229 VSS.n1822 0.04025
R11112 VSS.n8229 VSS.n8228 0.04025
R11113 VSS.n8228 VSS.n8227 0.04025
R11114 VSS.n8227 VSS.n1824 0.04025
R11115 VSS.n8223 VSS.n1824 0.04025
R11116 VSS.n8223 VSS.n8222 0.04025
R11117 VSS.n8222 VSS.n8221 0.04025
R11118 VSS.n8221 VSS.n1826 0.04025
R11119 VSS.n8217 VSS.n1826 0.04025
R11120 VSS.n8217 VSS.n8216 0.04025
R11121 VSS.n8216 VSS.n8215 0.04025
R11122 VSS.n8215 VSS.n1828 0.04025
R11123 VSS.n8211 VSS.n1828 0.04025
R11124 VSS.n8211 VSS.n8210 0.04025
R11125 VSS.n8210 VSS.n8209 0.04025
R11126 VSS.n8209 VSS.n1830 0.04025
R11127 VSS.n8205 VSS.n1830 0.04025
R11128 VSS.n8205 VSS.n8204 0.04025
R11129 VSS.n8204 VSS.n8203 0.04025
R11130 VSS.n8203 VSS.n1832 0.04025
R11131 VSS.n8199 VSS.n1832 0.04025
R11132 VSS.n8199 VSS.n8198 0.04025
R11133 VSS.n8198 VSS.n8197 0.04025
R11134 VSS.n8197 VSS.n1834 0.04025
R11135 VSS.n8193 VSS.n1834 0.04025
R11136 VSS.n8193 VSS.n8192 0.04025
R11137 VSS.n8192 VSS.n8191 0.04025
R11138 VSS.n8191 VSS.n1836 0.04025
R11139 VSS.n8187 VSS.n1836 0.04025
R11140 VSS.n8187 VSS.n8186 0.04025
R11141 VSS.n8186 VSS.n8185 0.04025
R11142 VSS.n8185 VSS.n1838 0.04025
R11143 VSS.n8181 VSS.n1838 0.04025
R11144 VSS.n8181 VSS.n8180 0.04025
R11145 VSS.n8180 VSS.n8179 0.04025
R11146 VSS.n8179 VSS.n1840 0.04025
R11147 VSS.n8175 VSS.n1840 0.04025
R11148 VSS.n8175 VSS.n8174 0.04025
R11149 VSS.n8174 VSS.n8173 0.04025
R11150 VSS.n8173 VSS.n1842 0.04025
R11151 VSS.n8169 VSS.n1842 0.04025
R11152 VSS.n8169 VSS.n8168 0.04025
R11153 VSS.n8168 VSS.n8167 0.04025
R11154 VSS.n8167 VSS.n1844 0.04025
R11155 VSS.n8163 VSS.n1844 0.04025
R11156 VSS.n8163 VSS.n8162 0.04025
R11157 VSS.n8162 VSS.n8161 0.04025
R11158 VSS.n8161 VSS.n1846 0.04025
R11159 VSS.n8157 VSS.n1846 0.04025
R11160 VSS.n8157 VSS.n8156 0.04025
R11161 VSS.n8156 VSS.n8155 0.04025
R11162 VSS.n8155 VSS.n1848 0.04025
R11163 VSS.n8151 VSS.n1848 0.04025
R11164 VSS.n8151 VSS.n8150 0.04025
R11165 VSS.n8150 VSS.n8149 0.04025
R11166 VSS.n8149 VSS.n1850 0.04025
R11167 VSS.n8145 VSS.n1850 0.04025
R11168 VSS.n8145 VSS.n8144 0.04025
R11169 VSS.n8144 VSS.n8143 0.04025
R11170 VSS.n8143 VSS.n1852 0.04025
R11171 VSS.n8139 VSS.n1852 0.04025
R11172 VSS.n8139 VSS.n8138 0.04025
R11173 VSS.n8138 VSS.n8137 0.04025
R11174 VSS.n8137 VSS.n1854 0.04025
R11175 VSS.n8133 VSS.n1854 0.04025
R11176 VSS.n8133 VSS.n8132 0.04025
R11177 VSS.n8132 VSS.n8131 0.04025
R11178 VSS.n8131 VSS.n1856 0.04025
R11179 VSS.n8127 VSS.n1856 0.04025
R11180 VSS.n8127 VSS.n8126 0.04025
R11181 VSS.n8126 VSS.n8125 0.04025
R11182 VSS.n8125 VSS.n1858 0.04025
R11183 VSS.n8121 VSS.n1858 0.04025
R11184 VSS.n8121 VSS.n8120 0.04025
R11185 VSS.n8120 VSS.n8119 0.04025
R11186 VSS.n8119 VSS.n1860 0.04025
R11187 VSS.n8115 VSS.n1860 0.04025
R11188 VSS.n8115 VSS.n8114 0.04025
R11189 VSS.n8114 VSS.n8113 0.04025
R11190 VSS.n8113 VSS.n1862 0.04025
R11191 VSS.n8109 VSS.n1862 0.04025
R11192 VSS.n8109 VSS.n8108 0.04025
R11193 VSS.n8108 VSS.n8107 0.04025
R11194 VSS.n8107 VSS.n1864 0.04025
R11195 VSS.n8103 VSS.n1864 0.04025
R11196 VSS.n8103 VSS.n8102 0.04025
R11197 VSS.n8102 VSS.n8101 0.04025
R11198 VSS.n8101 VSS.n1866 0.04025
R11199 VSS.n8097 VSS.n1866 0.04025
R11200 VSS.n8097 VSS.n8096 0.04025
R11201 VSS.n8096 VSS.n8095 0.04025
R11202 VSS.n8095 VSS.n1868 0.04025
R11203 VSS.n8091 VSS.n1868 0.04025
R11204 VSS.n8091 VSS.n8090 0.04025
R11205 VSS.n8090 VSS.n8089 0.04025
R11206 VSS.n8089 VSS.n1870 0.04025
R11207 VSS.n8085 VSS.n1870 0.04025
R11208 VSS.n8085 VSS.n8084 0.04025
R11209 VSS.n8084 VSS.n8083 0.04025
R11210 VSS.n8083 VSS.n1872 0.04025
R11211 VSS.n8079 VSS.n1872 0.04025
R11212 VSS.n8079 VSS.n8078 0.04025
R11213 VSS.n8078 VSS.n8077 0.04025
R11214 VSS.n8077 VSS.n1874 0.04025
R11215 VSS.n8073 VSS.n1874 0.04025
R11216 VSS.n8073 VSS.n8072 0.04025
R11217 VSS.n8072 VSS.n8071 0.04025
R11218 VSS.n8071 VSS.n1876 0.04025
R11219 VSS.n8067 VSS.n1876 0.04025
R11220 VSS.n8067 VSS.n8066 0.04025
R11221 VSS.n8066 VSS.n8065 0.04025
R11222 VSS.n8065 VSS.n1878 0.04025
R11223 VSS.n8061 VSS.n1878 0.04025
R11224 VSS.n8061 VSS.n8060 0.04025
R11225 VSS.n8060 VSS.n8059 0.04025
R11226 VSS.n8059 VSS.n1880 0.04025
R11227 VSS.n8055 VSS.n1880 0.04025
R11228 VSS.n8055 VSS.n8054 0.04025
R11229 VSS.n8054 VSS.n8053 0.04025
R11230 VSS.n8053 VSS.n1882 0.04025
R11231 VSS.n8049 VSS.n1882 0.04025
R11232 VSS.n8049 VSS.n8048 0.04025
R11233 VSS.n8048 VSS.n8047 0.04025
R11234 VSS.n8047 VSS.n1884 0.04025
R11235 VSS.n8043 VSS.n1884 0.04025
R11236 VSS.n8043 VSS.n8042 0.04025
R11237 VSS.n8042 VSS.n8041 0.04025
R11238 VSS.n8041 VSS.n1886 0.04025
R11239 VSS.n8037 VSS.n1886 0.04025
R11240 VSS.n8037 VSS.n8036 0.04025
R11241 VSS.n8036 VSS.n8035 0.04025
R11242 VSS.n8035 VSS.n1888 0.04025
R11243 VSS.n8031 VSS.n1888 0.04025
R11244 VSS.n8031 VSS.n8030 0.04025
R11245 VSS.n8030 VSS.n8029 0.04025
R11246 VSS.n8029 VSS.n1890 0.04025
R11247 VSS.n8025 VSS.n1890 0.04025
R11248 VSS.n8025 VSS.n8024 0.04025
R11249 VSS.n8024 VSS.n8023 0.04025
R11250 VSS.n8023 VSS.n1892 0.04025
R11251 VSS.n8019 VSS.n1892 0.04025
R11252 VSS.n8019 VSS.n8018 0.04025
R11253 VSS.n8018 VSS.n8017 0.04025
R11254 VSS.n8017 VSS.n1894 0.04025
R11255 VSS.n8013 VSS.n1894 0.04025
R11256 VSS.n8013 VSS.n8012 0.04025
R11257 VSS.n8012 VSS.n8011 0.04025
R11258 VSS.n8011 VSS.n1896 0.04025
R11259 VSS.n8007 VSS.n1896 0.04025
R11260 VSS.n8007 VSS.n8006 0.04025
R11261 VSS.n8006 VSS.n8005 0.04025
R11262 VSS.n8005 VSS.n1898 0.04025
R11263 VSS.n8001 VSS.n1898 0.04025
R11264 VSS.n8001 VSS.n8000 0.04025
R11265 VSS.n8000 VSS.n7999 0.04025
R11266 VSS.n7999 VSS.n1900 0.04025
R11267 VSS.n7995 VSS.n1900 0.04025
R11268 VSS.n7995 VSS.n7994 0.04025
R11269 VSS.n7994 VSS.n7993 0.04025
R11270 VSS.n7993 VSS.n1902 0.04025
R11271 VSS.n7989 VSS.n1902 0.04025
R11272 VSS.n7989 VSS.n7988 0.04025
R11273 VSS.n7988 VSS.n7987 0.04025
R11274 VSS.n7987 VSS.n1904 0.04025
R11275 VSS.n7983 VSS.n1904 0.04025
R11276 VSS.n7983 VSS.n7982 0.04025
R11277 VSS.n7982 VSS.n7981 0.04025
R11278 VSS.n7981 VSS.n1906 0.04025
R11279 VSS.n7977 VSS.n1906 0.04025
R11280 VSS.n7977 VSS.n7976 0.04025
R11281 VSS.n7976 VSS.n7975 0.04025
R11282 VSS.n7975 VSS.n1908 0.04025
R11283 VSS.n7971 VSS.n1908 0.04025
R11284 VSS.n7971 VSS.n7970 0.04025
R11285 VSS.n7970 VSS.n7969 0.04025
R11286 VSS.n7969 VSS.n1910 0.04025
R11287 VSS.n7965 VSS.n1910 0.04025
R11288 VSS.n7965 VSS.n7964 0.04025
R11289 VSS.n7964 VSS.n7963 0.04025
R11290 VSS.n7963 VSS.n1912 0.04025
R11291 VSS.n7959 VSS.n1912 0.04025
R11292 VSS.n7959 VSS.n7958 0.04025
R11293 VSS.n7958 VSS.n7957 0.04025
R11294 VSS.n7957 VSS.n1914 0.04025
R11295 VSS.n7953 VSS.n1914 0.04025
R11296 VSS.n7953 VSS.n7952 0.04025
R11297 VSS.n7952 VSS.n7951 0.04025
R11298 VSS.n7951 VSS.n1916 0.04025
R11299 VSS.n7947 VSS.n1916 0.04025
R11300 VSS.n7947 VSS.n7946 0.04025
R11301 VSS.n7946 VSS.n7945 0.04025
R11302 VSS.n7945 VSS.n1918 0.04025
R11303 VSS.n7941 VSS.n1918 0.04025
R11304 VSS.n7941 VSS.n7940 0.04025
R11305 VSS.n7940 VSS.n7939 0.04025
R11306 VSS.n7939 VSS.n1920 0.04025
R11307 VSS.n7935 VSS.n1920 0.04025
R11308 VSS.n7935 VSS.n7934 0.04025
R11309 VSS.n7934 VSS.n7933 0.04025
R11310 VSS.n7933 VSS.n1922 0.04025
R11311 VSS.n7929 VSS.n1922 0.04025
R11312 VSS.n7929 VSS.n7928 0.04025
R11313 VSS.n7928 VSS.n7927 0.04025
R11314 VSS.n7927 VSS.n1924 0.04025
R11315 VSS.n7923 VSS.n1924 0.04025
R11316 VSS.n7923 VSS.n7922 0.04025
R11317 VSS.n7922 VSS.n7921 0.04025
R11318 VSS.n7921 VSS.n1926 0.04025
R11319 VSS.n7917 VSS.n1926 0.04025
R11320 VSS.n7917 VSS.n7916 0.04025
R11321 VSS.n7916 VSS.n7915 0.04025
R11322 VSS.n7915 VSS.n1928 0.04025
R11323 VSS.n7911 VSS.n1928 0.04025
R11324 VSS.n7911 VSS.n7910 0.04025
R11325 VSS.n7910 VSS.n7909 0.04025
R11326 VSS.n7909 VSS.n1930 0.04025
R11327 VSS.n7905 VSS.n1930 0.04025
R11328 VSS.n7905 VSS.n7904 0.04025
R11329 VSS.n7904 VSS.n7903 0.04025
R11330 VSS.n7903 VSS.n1932 0.04025
R11331 VSS.n7899 VSS.n1932 0.04025
R11332 VSS.n7899 VSS.n7898 0.04025
R11333 VSS.n7898 VSS.n7897 0.04025
R11334 VSS.n7897 VSS.n1934 0.04025
R11335 VSS.n7893 VSS.n1934 0.04025
R11336 VSS.n7893 VSS.n7892 0.04025
R11337 VSS.n7892 VSS.n7891 0.04025
R11338 VSS.n7891 VSS.n1936 0.04025
R11339 VSS.n7887 VSS.n1936 0.04025
R11340 VSS.n7887 VSS.n7886 0.04025
R11341 VSS.n7886 VSS.n7885 0.04025
R11342 VSS.n7885 VSS.n1938 0.04025
R11343 VSS.n7881 VSS.n1938 0.04025
R11344 VSS.n7881 VSS.n7880 0.04025
R11345 VSS.n7880 VSS.n7879 0.04025
R11346 VSS.n7879 VSS.n1940 0.04025
R11347 VSS.n7875 VSS.n1940 0.04025
R11348 VSS.n7875 VSS.n7874 0.04025
R11349 VSS.n7874 VSS.n7873 0.04025
R11350 VSS.n7873 VSS.n1942 0.04025
R11351 VSS.n7869 VSS.n1942 0.04025
R11352 VSS.n7869 VSS.n7868 0.04025
R11353 VSS.n7868 VSS.n7867 0.04025
R11354 VSS.n7867 VSS.n1944 0.04025
R11355 VSS.n7863 VSS.n1944 0.04025
R11356 VSS.n7863 VSS.n7862 0.04025
R11357 VSS.n7862 VSS.n7861 0.04025
R11358 VSS.n7861 VSS.n1946 0.04025
R11359 VSS.n7857 VSS.n1946 0.04025
R11360 VSS.n7857 VSS.n7856 0.04025
R11361 VSS.n7856 VSS.n7855 0.04025
R11362 VSS.n7855 VSS.n1948 0.04025
R11363 VSS.n7851 VSS.n1948 0.04025
R11364 VSS.n7851 VSS.n7850 0.04025
R11365 VSS.n7850 VSS.n7849 0.04025
R11366 VSS.n7849 VSS.n1950 0.04025
R11367 VSS.n7845 VSS.n1950 0.04025
R11368 VSS.n7845 VSS.n7844 0.04025
R11369 VSS.n7844 VSS.n7843 0.04025
R11370 VSS.n7843 VSS.n1952 0.04025
R11371 VSS.n7839 VSS.n1952 0.04025
R11372 VSS.n7839 VSS.n7838 0.04025
R11373 VSS.n7838 VSS.n7837 0.04025
R11374 VSS.n7837 VSS.n1954 0.04025
R11375 VSS.n7833 VSS.n1954 0.04025
R11376 VSS.n7833 VSS.n7832 0.04025
R11377 VSS.n7832 VSS.n7831 0.04025
R11378 VSS.n7831 VSS.n1956 0.04025
R11379 VSS.n7827 VSS.n1956 0.04025
R11380 VSS.n7827 VSS.n7826 0.04025
R11381 VSS.n7826 VSS.n7825 0.04025
R11382 VSS.n7825 VSS.n1958 0.04025
R11383 VSS.n7821 VSS.n1958 0.04025
R11384 VSS.n7821 VSS.n7820 0.04025
R11385 VSS.n7820 VSS.n7819 0.04025
R11386 VSS.n7819 VSS.n1960 0.04025
R11387 VSS.n7815 VSS.n1960 0.04025
R11388 VSS.n7815 VSS.n7814 0.04025
R11389 VSS.n7814 VSS.n7813 0.04025
R11390 VSS.n7813 VSS.n1962 0.04025
R11391 VSS.n7809 VSS.n1962 0.04025
R11392 VSS.n7809 VSS.n7808 0.04025
R11393 VSS.n7808 VSS.n7807 0.04025
R11394 VSS.n7807 VSS.n1964 0.04025
R11395 VSS.n7803 VSS.n1964 0.04025
R11396 VSS.n7803 VSS.n7802 0.04025
R11397 VSS.n7802 VSS.n7801 0.04025
R11398 VSS.n7801 VSS.n1966 0.04025
R11399 VSS.n7797 VSS.n1966 0.04025
R11400 VSS.n7797 VSS.n7796 0.04025
R11401 VSS.n7796 VSS.n7795 0.04025
R11402 VSS.n7795 VSS.n1968 0.04025
R11403 VSS.n7791 VSS.n1968 0.04025
R11404 VSS.n7791 VSS.n7790 0.04025
R11405 VSS.n7790 VSS.n7789 0.04025
R11406 VSS.n7789 VSS.n1970 0.04025
R11407 VSS.n7785 VSS.n1970 0.04025
R11408 VSS.n7785 VSS.n7784 0.04025
R11409 VSS.n7784 VSS.n7783 0.04025
R11410 VSS.n7783 VSS.n1972 0.04025
R11411 VSS.n7779 VSS.n1972 0.04025
R11412 VSS.n7779 VSS.n7778 0.04025
R11413 VSS.n7778 VSS.n7777 0.04025
R11414 VSS.n7777 VSS.n1974 0.04025
R11415 VSS.n7773 VSS.n1974 0.04025
R11416 VSS.n7773 VSS.n7772 0.04025
R11417 VSS.n7772 VSS.n7771 0.04025
R11418 VSS.n7771 VSS.n1976 0.04025
R11419 VSS.n7767 VSS.n1976 0.04025
R11420 VSS.n7767 VSS.n7766 0.04025
R11421 VSS.n7766 VSS.n7765 0.04025
R11422 VSS.n7765 VSS.n1978 0.04025
R11423 VSS.n7761 VSS.n1978 0.04025
R11424 VSS.n7761 VSS.n7760 0.04025
R11425 VSS.n7760 VSS.n7759 0.04025
R11426 VSS.n7759 VSS.n1980 0.04025
R11427 VSS.n7755 VSS.n1980 0.04025
R11428 VSS.n7755 VSS.n7754 0.04025
R11429 VSS.n7754 VSS.n7753 0.04025
R11430 VSS.n7753 VSS.n1982 0.04025
R11431 VSS.n7749 VSS.n1982 0.04025
R11432 VSS.n7749 VSS.n7748 0.04025
R11433 VSS.n7748 VSS.n7747 0.04025
R11434 VSS.n7747 VSS.n1984 0.04025
R11435 VSS.n7743 VSS.n1984 0.04025
R11436 VSS.n7743 VSS.n7742 0.04025
R11437 VSS.n7742 VSS.n7741 0.04025
R11438 VSS.n7741 VSS.n1986 0.04025
R11439 VSS.n7737 VSS.n1986 0.04025
R11440 VSS.n7737 VSS.n7736 0.04025
R11441 VSS.n7736 VSS.n7735 0.04025
R11442 VSS.n7735 VSS.n1988 0.04025
R11443 VSS.n7731 VSS.n1988 0.04025
R11444 VSS.n7731 VSS.n7730 0.04025
R11445 VSS.n7730 VSS.n7729 0.04025
R11446 VSS.n7729 VSS.n1990 0.04025
R11447 VSS.n7725 VSS.n1990 0.04025
R11448 VSS.n7725 VSS.n7724 0.04025
R11449 VSS.n7724 VSS.n7723 0.04025
R11450 VSS.n7723 VSS.n1992 0.04025
R11451 VSS.n7719 VSS.n1992 0.04025
R11452 VSS.n7719 VSS.n7718 0.04025
R11453 VSS.n7718 VSS.n7717 0.04025
R11454 VSS.n7717 VSS.n1994 0.04025
R11455 VSS.n7713 VSS.n1994 0.04025
R11456 VSS.n7713 VSS.n7712 0.04025
R11457 VSS.n7712 VSS.n7711 0.04025
R11458 VSS.n7711 VSS.n1996 0.04025
R11459 VSS.n7707 VSS.n1996 0.04025
R11460 VSS.n7707 VSS.n7706 0.04025
R11461 VSS.n7706 VSS.n7705 0.04025
R11462 VSS.n7705 VSS.n1998 0.04025
R11463 VSS.n7701 VSS.n1998 0.04025
R11464 VSS.n7701 VSS.n7700 0.04025
R11465 VSS.n7700 VSS.n7699 0.04025
R11466 VSS.n7699 VSS.n2000 0.04025
R11467 VSS.n7695 VSS.n2000 0.04025
R11468 VSS.n7695 VSS.n7694 0.04025
R11469 VSS.n7694 VSS.n7693 0.04025
R11470 VSS.n7693 VSS.n2002 0.04025
R11471 VSS.n7689 VSS.n2002 0.04025
R11472 VSS.n7689 VSS.n7688 0.04025
R11473 VSS.n7688 VSS.n7687 0.04025
R11474 VSS.n7687 VSS.n2004 0.04025
R11475 VSS.n7683 VSS.n2004 0.04025
R11476 VSS.n7683 VSS.n7682 0.04025
R11477 VSS.n7682 VSS.n7681 0.04025
R11478 VSS.n7681 VSS.n2006 0.04025
R11479 VSS.n7677 VSS.n2006 0.04025
R11480 VSS.n7677 VSS.n7676 0.04025
R11481 VSS.n7676 VSS.n7675 0.04025
R11482 VSS.n7675 VSS.n2008 0.04025
R11483 VSS.n7671 VSS.n2008 0.04025
R11484 VSS.n7671 VSS.n7670 0.04025
R11485 VSS.n7670 VSS.n7669 0.04025
R11486 VSS.n7669 VSS.n2010 0.04025
R11487 VSS.n7665 VSS.n2010 0.04025
R11488 VSS.n7665 VSS.n7664 0.04025
R11489 VSS.n7664 VSS.n7663 0.04025
R11490 VSS.n7663 VSS.n2012 0.04025
R11491 VSS.n7659 VSS.n2012 0.04025
R11492 VSS.n7659 VSS.n7658 0.04025
R11493 VSS.n7658 VSS.n7657 0.04025
R11494 VSS.n7657 VSS.n2014 0.04025
R11495 VSS.n7653 VSS.n2014 0.04025
R11496 VSS.n7653 VSS.n7652 0.04025
R11497 VSS.n7652 VSS.n7651 0.04025
R11498 VSS.n7651 VSS.n2016 0.04025
R11499 VSS.n7647 VSS.n2016 0.04025
R11500 VSS.n7647 VSS.n7646 0.04025
R11501 VSS.n7646 VSS.n7645 0.04025
R11502 VSS.n7645 VSS.n2018 0.04025
R11503 VSS.n7641 VSS.n2018 0.04025
R11504 VSS.n7641 VSS.n7640 0.04025
R11505 VSS.n7640 VSS.n7639 0.04025
R11506 VSS.n7639 VSS.n2020 0.04025
R11507 VSS.n7635 VSS.n2020 0.04025
R11508 VSS.n7635 VSS.n7634 0.04025
R11509 VSS.n7634 VSS.n7633 0.04025
R11510 VSS.n7633 VSS.n2022 0.04025
R11511 VSS.n7629 VSS.n2022 0.04025
R11512 VSS.n7629 VSS.n7628 0.04025
R11513 VSS.n7628 VSS.n7627 0.04025
R11514 VSS.n7627 VSS.n2024 0.04025
R11515 VSS.n7623 VSS.n2024 0.04025
R11516 VSS.n7623 VSS.n7622 0.04025
R11517 VSS.n7622 VSS.n7621 0.04025
R11518 VSS.n7621 VSS.n2026 0.04025
R11519 VSS.n7617 VSS.n2026 0.04025
R11520 VSS.n7617 VSS.n7616 0.04025
R11521 VSS.n7616 VSS.n7615 0.04025
R11522 VSS.n7615 VSS.n2028 0.04025
R11523 VSS.n7611 VSS.n2028 0.04025
R11524 VSS.n7611 VSS.n7610 0.04025
R11525 VSS.n7610 VSS.n7609 0.04025
R11526 VSS.n7609 VSS.n2030 0.04025
R11527 VSS.n7605 VSS.n2030 0.04025
R11528 VSS.n7605 VSS.n7604 0.04025
R11529 VSS.n7604 VSS.n7603 0.04025
R11530 VSS.n7603 VSS.n2032 0.04025
R11531 VSS.n7599 VSS.n2032 0.04025
R11532 VSS.n7599 VSS.n7598 0.04025
R11533 VSS.n7598 VSS.n7597 0.04025
R11534 VSS.n7597 VSS.n2034 0.04025
R11535 VSS.n7593 VSS.n2034 0.04025
R11536 VSS.n7593 VSS.n7592 0.04025
R11537 VSS.n7592 VSS.n7591 0.04025
R11538 VSS.n7591 VSS.n2036 0.04025
R11539 VSS.n7587 VSS.n2036 0.04025
R11540 VSS.n7587 VSS.n7586 0.04025
R11541 VSS.n7586 VSS.n7585 0.04025
R11542 VSS.n7585 VSS.n2038 0.04025
R11543 VSS.n7581 VSS.n2038 0.04025
R11544 VSS.n7581 VSS.n7580 0.04025
R11545 VSS.n7580 VSS.n7579 0.04025
R11546 VSS.n7579 VSS.n2040 0.04025
R11547 VSS.n7575 VSS.n2040 0.04025
R11548 VSS.n7575 VSS.n7574 0.04025
R11549 VSS.n7574 VSS.n7573 0.04025
R11550 VSS.n7573 VSS.n2042 0.04025
R11551 VSS.n7569 VSS.n2042 0.04025
R11552 VSS.n7569 VSS.n7568 0.04025
R11553 VSS.n7568 VSS.n7567 0.04025
R11554 VSS.n7567 VSS.n2044 0.04025
R11555 VSS.n7563 VSS.n2044 0.04025
R11556 VSS.n7563 VSS.n7562 0.04025
R11557 VSS.n7562 VSS.n7561 0.04025
R11558 VSS.n7561 VSS.n2046 0.04025
R11559 VSS.n7557 VSS.n2046 0.04025
R11560 VSS.n7557 VSS.n7556 0.04025
R11561 VSS.n7556 VSS.n7555 0.04025
R11562 VSS.n7555 VSS.n2048 0.04025
R11563 VSS.n7551 VSS.n2048 0.04025
R11564 VSS.n7551 VSS.n7550 0.04025
R11565 VSS.n7550 VSS.n7549 0.04025
R11566 VSS.n7549 VSS.n2050 0.04025
R11567 VSS.n7545 VSS.n2050 0.04025
R11568 VSS.n7545 VSS.n7544 0.04025
R11569 VSS.n7544 VSS.n7543 0.04025
R11570 VSS.n7543 VSS.n2052 0.04025
R11571 VSS.n7539 VSS.n2052 0.04025
R11572 VSS.n7539 VSS.n7538 0.04025
R11573 VSS.n7538 VSS.n7537 0.04025
R11574 VSS.n7537 VSS.n2054 0.04025
R11575 VSS.n7533 VSS.n2054 0.04025
R11576 VSS.n7533 VSS.n7532 0.04025
R11577 VSS.n7532 VSS.n7531 0.04025
R11578 VSS.n7531 VSS.n2056 0.04025
R11579 VSS.n7527 VSS.n2056 0.04025
R11580 VSS.n7527 VSS.n7526 0.04025
R11581 VSS.n7526 VSS.n7525 0.04025
R11582 VSS.n7525 VSS.n2058 0.04025
R11583 VSS.n7521 VSS.n2058 0.04025
R11584 VSS.n7521 VSS.n7520 0.04025
R11585 VSS.n7520 VSS.n7519 0.04025
R11586 VSS.n7519 VSS.n2060 0.04025
R11587 VSS.n7515 VSS.n2060 0.04025
R11588 VSS.n7515 VSS.n7514 0.04025
R11589 VSS.n7514 VSS.n7513 0.04025
R11590 VSS.n7513 VSS.n2062 0.04025
R11591 VSS.n7509 VSS.n2062 0.04025
R11592 VSS.n7509 VSS.n7508 0.04025
R11593 VSS.n7508 VSS.n7507 0.04025
R11594 VSS.n7507 VSS.n2064 0.04025
R11595 VSS.n7503 VSS.n2064 0.04025
R11596 VSS.n7503 VSS.n7502 0.04025
R11597 VSS.n7502 VSS.n7501 0.04025
R11598 VSS.n7501 VSS.n2066 0.04025
R11599 VSS.n7497 VSS.n2066 0.04025
R11600 VSS.n7497 VSS.n7496 0.04025
R11601 VSS.n7496 VSS.n7495 0.04025
R11602 VSS.n7495 VSS.n2068 0.04025
R11603 VSS.n7491 VSS.n2068 0.04025
R11604 VSS.n7491 VSS.n7490 0.04025
R11605 VSS.n7490 VSS.n7489 0.04025
R11606 VSS.n7489 VSS.n2070 0.04025
R11607 VSS.n7485 VSS.n2070 0.04025
R11608 VSS.n7485 VSS.n7484 0.04025
R11609 VSS.n7484 VSS.n7483 0.04025
R11610 VSS.n7483 VSS.n2072 0.04025
R11611 VSS.n7479 VSS.n2072 0.04025
R11612 VSS.n7479 VSS.n7478 0.04025
R11613 VSS.n7478 VSS.n7477 0.04025
R11614 VSS.n7477 VSS.n2074 0.04025
R11615 VSS.n7473 VSS.n2074 0.04025
R11616 VSS.n7473 VSS.n7472 0.04025
R11617 VSS.n7472 VSS.n7471 0.04025
R11618 VSS.n7471 VSS.n2076 0.04025
R11619 VSS.n7467 VSS.n2076 0.04025
R11620 VSS.n7467 VSS.n7466 0.04025
R11621 VSS.n7466 VSS.n7465 0.04025
R11622 VSS.n7465 VSS.n2078 0.04025
R11623 VSS.n7461 VSS.n2078 0.04025
R11624 VSS.n7461 VSS.n7460 0.04025
R11625 VSS.n7460 VSS.n7459 0.04025
R11626 VSS.n7459 VSS.n2080 0.04025
R11627 VSS.n7455 VSS.n2080 0.04025
R11628 VSS.n7455 VSS.n7454 0.04025
R11629 VSS.n7454 VSS.n7453 0.04025
R11630 VSS.n7453 VSS.n2082 0.04025
R11631 VSS.n7449 VSS.n2082 0.04025
R11632 VSS.n7449 VSS.n7448 0.04025
R11633 VSS.n7448 VSS.n7447 0.04025
R11634 VSS.n7447 VSS.n2084 0.04025
R11635 VSS.n7443 VSS.n2084 0.04025
R11636 VSS.n7443 VSS.n7442 0.04025
R11637 VSS.n7442 VSS.n7441 0.04025
R11638 VSS.n7441 VSS.n2086 0.04025
R11639 VSS.n7437 VSS.n2086 0.04025
R11640 VSS.n7437 VSS.n7436 0.04025
R11641 VSS.n7436 VSS.n7435 0.04025
R11642 VSS.n7435 VSS.n2088 0.04025
R11643 VSS.n7431 VSS.n2088 0.04025
R11644 VSS.n7431 VSS.n7430 0.04025
R11645 VSS.n7430 VSS.n7429 0.04025
R11646 VSS.n7429 VSS.n2090 0.04025
R11647 VSS.n7425 VSS.n2090 0.04025
R11648 VSS.n7425 VSS.n7424 0.04025
R11649 VSS.n7424 VSS.n7423 0.04025
R11650 VSS.n7423 VSS.n2092 0.04025
R11651 VSS.n7419 VSS.n2092 0.04025
R11652 VSS.n7419 VSS.n7418 0.04025
R11653 VSS.n7418 VSS.n7417 0.04025
R11654 VSS.n7417 VSS.n2094 0.04025
R11655 VSS.n7413 VSS.n2094 0.04025
R11656 VSS.n7413 VSS.n7412 0.04025
R11657 VSS.n7412 VSS.n7411 0.04025
R11658 VSS.n7411 VSS.n2096 0.04025
R11659 VSS.n7407 VSS.n2096 0.04025
R11660 VSS.n7407 VSS.n7406 0.04025
R11661 VSS.n7406 VSS.n7405 0.04025
R11662 VSS.n7405 VSS.n2098 0.04025
R11663 VSS.n7401 VSS.n2098 0.04025
R11664 VSS.n7401 VSS.n7400 0.04025
R11665 VSS.n7400 VSS.n7399 0.04025
R11666 VSS.n7399 VSS.n2100 0.04025
R11667 VSS.n7395 VSS.n2100 0.04025
R11668 VSS.n7395 VSS.n7394 0.04025
R11669 VSS.n7394 VSS.n7393 0.04025
R11670 VSS.n7393 VSS.n2102 0.04025
R11671 VSS.n7389 VSS.n2102 0.04025
R11672 VSS.n7389 VSS.n7388 0.04025
R11673 VSS.n7388 VSS.n7387 0.04025
R11674 VSS.n7387 VSS.n2104 0.04025
R11675 VSS.n7383 VSS.n2104 0.04025
R11676 VSS.n7383 VSS.n7382 0.04025
R11677 VSS.n7382 VSS.n7381 0.04025
R11678 VSS.n7381 VSS.n2106 0.04025
R11679 VSS.n7377 VSS.n2106 0.04025
R11680 VSS.n7377 VSS.n7376 0.04025
R11681 VSS.n7376 VSS.n7375 0.04025
R11682 VSS.n7375 VSS.n2108 0.04025
R11683 VSS.n7371 VSS.n2108 0.04025
R11684 VSS.n7371 VSS.n7370 0.04025
R11685 VSS.n7370 VSS.n7369 0.04025
R11686 VSS.n7369 VSS.n2110 0.04025
R11687 VSS.n7365 VSS.n2110 0.04025
R11688 VSS.n7365 VSS.n7364 0.04025
R11689 VSS.n7364 VSS.n7363 0.04025
R11690 VSS.n7363 VSS.n2112 0.04025
R11691 VSS.n7359 VSS.n2112 0.04025
R11692 VSS.n7359 VSS.n7358 0.04025
R11693 VSS.n7358 VSS.n7357 0.04025
R11694 VSS.n7357 VSS.n2114 0.04025
R11695 VSS.n7353 VSS.n2114 0.04025
R11696 VSS.n7353 VSS.n7352 0.04025
R11697 VSS.n7352 VSS.n7351 0.04025
R11698 VSS.n7351 VSS.n2116 0.04025
R11699 VSS.n7347 VSS.n2116 0.04025
R11700 VSS.n7347 VSS.n7346 0.04025
R11701 VSS.n7346 VSS.n7345 0.04025
R11702 VSS.n7345 VSS.n2118 0.04025
R11703 VSS.n7341 VSS.n2118 0.04025
R11704 VSS.n7341 VSS.n7340 0.04025
R11705 VSS.n7340 VSS.n7339 0.04025
R11706 VSS.n7339 VSS.n2120 0.04025
R11707 VSS.n7335 VSS.n2120 0.04025
R11708 VSS.n7335 VSS.n7334 0.04025
R11709 VSS.n7334 VSS.n7333 0.04025
R11710 VSS.n7333 VSS.n2122 0.04025
R11711 VSS.n7329 VSS.n2122 0.04025
R11712 VSS.n7329 VSS.n7328 0.04025
R11713 VSS.n7328 VSS.n7327 0.04025
R11714 VSS.n7327 VSS.n2124 0.04025
R11715 VSS.n7323 VSS.n2124 0.04025
R11716 VSS.n7323 VSS.n7322 0.04025
R11717 VSS.n7322 VSS.n7321 0.04025
R11718 VSS.n7321 VSS.n2126 0.04025
R11719 VSS.n7317 VSS.n2126 0.04025
R11720 VSS.n7317 VSS.n7316 0.04025
R11721 VSS.n7316 VSS.n7315 0.04025
R11722 VSS.n7315 VSS.n2128 0.04025
R11723 VSS.n7311 VSS.n2128 0.04025
R11724 VSS.n7311 VSS.n7310 0.04025
R11725 VSS.n7310 VSS.n7309 0.04025
R11726 VSS.n7309 VSS.n2130 0.04025
R11727 VSS.n7305 VSS.n2130 0.04025
R11728 VSS.n7305 VSS.n7304 0.04025
R11729 VSS.n7304 VSS.n7303 0.04025
R11730 VSS.n7303 VSS.n2132 0.04025
R11731 VSS.n7299 VSS.n2132 0.04025
R11732 VSS.n7299 VSS.n7298 0.04025
R11733 VSS.n7298 VSS.n7297 0.04025
R11734 VSS.n7297 VSS.n2134 0.04025
R11735 VSS.n7293 VSS.n2134 0.04025
R11736 VSS.n7293 VSS.n7292 0.04025
R11737 VSS.n7292 VSS.n7291 0.04025
R11738 VSS.n7291 VSS.n2136 0.04025
R11739 VSS.n7287 VSS.n2136 0.04025
R11740 VSS.n7287 VSS.n7286 0.04025
R11741 VSS.n7286 VSS.n7285 0.04025
R11742 VSS.n7285 VSS.n2138 0.04025
R11743 VSS.n7281 VSS.n2138 0.04025
R11744 VSS.n7281 VSS.n7280 0.04025
R11745 VSS.n7280 VSS.n7279 0.04025
R11746 VSS.n7279 VSS.n2140 0.04025
R11747 VSS.n7275 VSS.n2140 0.04025
R11748 VSS.n7275 VSS.n7274 0.04025
R11749 VSS.n7274 VSS.n7273 0.04025
R11750 VSS.n7273 VSS.n2142 0.04025
R11751 VSS.n7269 VSS.n2142 0.04025
R11752 VSS.n7269 VSS.n7268 0.04025
R11753 VSS.n7268 VSS.n7267 0.04025
R11754 VSS.n7267 VSS.n2144 0.04025
R11755 VSS.n7263 VSS.n2144 0.04025
R11756 VSS.n7263 VSS.n7262 0.04025
R11757 VSS.n7262 VSS.n7261 0.04025
R11758 VSS.n7261 VSS.n2146 0.04025
R11759 VSS.n7257 VSS.n2146 0.04025
R11760 VSS.n7257 VSS.n7256 0.04025
R11761 VSS.n7256 VSS.n7255 0.04025
R11762 VSS.n7255 VSS.n2148 0.04025
R11763 VSS.n7251 VSS.n2148 0.04025
R11764 VSS.n7251 VSS.n7250 0.04025
R11765 VSS.n7250 VSS.n7249 0.04025
R11766 VSS.n7249 VSS.n2150 0.04025
R11767 VSS.n7245 VSS.n2150 0.04025
R11768 VSS.n7245 VSS.n7244 0.04025
R11769 VSS.n7244 VSS.n7243 0.04025
R11770 VSS.n7243 VSS.n2152 0.04025
R11771 VSS.n7239 VSS.n2152 0.04025
R11772 VSS.n7239 VSS.n7238 0.04025
R11773 VSS.n7238 VSS.n7237 0.04025
R11774 VSS.n7237 VSS.n2154 0.04025
R11775 VSS.n7233 VSS.n2154 0.04025
R11776 VSS.n7233 VSS.n7232 0.04025
R11777 VSS.n7232 VSS.n7231 0.04025
R11778 VSS.n7231 VSS.n2156 0.04025
R11779 VSS.n7227 VSS.n2156 0.04025
R11780 VSS.n7227 VSS.n7226 0.04025
R11781 VSS.n7226 VSS.n7225 0.04025
R11782 VSS.n7225 VSS.n2158 0.04025
R11783 VSS.n7221 VSS.n2158 0.04025
R11784 VSS.n7221 VSS.n7220 0.04025
R11785 VSS.n7220 VSS.n7219 0.04025
R11786 VSS.n7219 VSS.n2160 0.04025
R11787 VSS.n7215 VSS.n2160 0.04025
R11788 VSS.n7215 VSS.n7214 0.04025
R11789 VSS.n7214 VSS.n7213 0.04025
R11790 VSS.n7213 VSS.n2162 0.04025
R11791 VSS.n7209 VSS.n2162 0.04025
R11792 VSS.n7209 VSS.n7208 0.04025
R11793 VSS.n7208 VSS.n7207 0.04025
R11794 VSS.n7207 VSS.n2164 0.04025
R11795 VSS.n7203 VSS.n2164 0.04025
R11796 VSS.n7203 VSS.n7202 0.04025
R11797 VSS.n7202 VSS.n7201 0.04025
R11798 VSS.n7201 VSS.n2166 0.04025
R11799 VSS.n7197 VSS.n2166 0.04025
R11800 VSS.n7197 VSS.n7196 0.04025
R11801 VSS.n7196 VSS.n7195 0.04025
R11802 VSS.n7195 VSS.n2168 0.04025
R11803 VSS.n7191 VSS.n2168 0.04025
R11804 VSS.n7191 VSS.n7190 0.04025
R11805 VSS.n7190 VSS.n7189 0.04025
R11806 VSS.n7189 VSS.n2170 0.04025
R11807 VSS.n7185 VSS.n2170 0.04025
R11808 VSS.n7185 VSS.n7184 0.04025
R11809 VSS.n7184 VSS.n7183 0.04025
R11810 VSS.n7183 VSS.n2172 0.04025
R11811 VSS.n7179 VSS.n2172 0.04025
R11812 VSS.n7179 VSS.n7178 0.04025
R11813 VSS.n7178 VSS.n7177 0.04025
R11814 VSS.n7177 VSS.n2174 0.04025
R11815 VSS.n7173 VSS.n2174 0.04025
R11816 VSS.n7173 VSS.n7172 0.04025
R11817 VSS.n7172 VSS.n7171 0.04025
R11818 VSS.n7171 VSS.n2176 0.04025
R11819 VSS.n7167 VSS.n2176 0.04025
R11820 VSS.n7167 VSS.n7166 0.04025
R11821 VSS.n7166 VSS.n7165 0.04025
R11822 VSS.n7165 VSS.n2178 0.04025
R11823 VSS.n7161 VSS.n2178 0.04025
R11824 VSS.n7161 VSS.n7160 0.04025
R11825 VSS.n7160 VSS.n7159 0.04025
R11826 VSS.n7159 VSS.n2180 0.04025
R11827 VSS.n7155 VSS.n2180 0.04025
R11828 VSS.n7155 VSS.n7154 0.04025
R11829 VSS.n7154 VSS.n7153 0.04025
R11830 VSS.n7153 VSS.n2182 0.04025
R11831 VSS.n7149 VSS.n2182 0.04025
R11832 VSS.n7149 VSS.n7148 0.04025
R11833 VSS.n7148 VSS.n7147 0.04025
R11834 VSS.n7147 VSS.n2184 0.04025
R11835 VSS.n7143 VSS.n2184 0.04025
R11836 VSS.n7143 VSS.n7142 0.04025
R11837 VSS.n7142 VSS.n7141 0.04025
R11838 VSS.n7141 VSS.n2186 0.04025
R11839 VSS.n7137 VSS.n2186 0.04025
R11840 VSS.n7137 VSS.n7136 0.04025
R11841 VSS.n7136 VSS.n7135 0.04025
R11842 VSS.n7135 VSS.n2188 0.04025
R11843 VSS.n7131 VSS.n2188 0.04025
R11844 VSS.n7131 VSS.n7130 0.04025
R11845 VSS.n7130 VSS.n7129 0.04025
R11846 VSS.n7129 VSS.n2190 0.04025
R11847 VSS.n7125 VSS.n2190 0.04025
R11848 VSS.n7125 VSS.n7124 0.04025
R11849 VSS.n7124 VSS.n7123 0.04025
R11850 VSS.n7123 VSS.n2192 0.04025
R11851 VSS.n7119 VSS.n2192 0.04025
R11852 VSS.n7119 VSS.n7118 0.04025
R11853 VSS.n7118 VSS.n7117 0.04025
R11854 VSS.n7117 VSS.n2194 0.04025
R11855 VSS.n7113 VSS.n2194 0.04025
R11856 VSS.n7113 VSS.n7112 0.04025
R11857 VSS.n7112 VSS.n7111 0.04025
R11858 VSS.n7111 VSS.n2196 0.04025
R11859 VSS.n7107 VSS.n2196 0.04025
R11860 VSS.n7107 VSS.n7106 0.04025
R11861 VSS.n7106 VSS.n7105 0.04025
R11862 VSS.n7105 VSS.n2198 0.04025
R11863 VSS.n7101 VSS.n2198 0.04025
R11864 VSS.n7101 VSS.n7100 0.04025
R11865 VSS.n7100 VSS.n7099 0.04025
R11866 VSS.n7099 VSS.n2200 0.04025
R11867 VSS.n7095 VSS.n2200 0.04025
R11868 VSS.n7095 VSS.n7094 0.04025
R11869 VSS.n7094 VSS.n7093 0.04025
R11870 VSS.n7093 VSS.n2202 0.04025
R11871 VSS.n7089 VSS.n2202 0.04025
R11872 VSS.n7089 VSS.n7088 0.04025
R11873 VSS.n7088 VSS.n7087 0.04025
R11874 VSS.n7087 VSS.n2204 0.04025
R11875 VSS.n7083 VSS.n2204 0.04025
R11876 VSS.n7083 VSS.n7082 0.04025
R11877 VSS.n7082 VSS.n7081 0.04025
R11878 VSS.n7081 VSS.n2206 0.04025
R11879 VSS.n7077 VSS.n2206 0.04025
R11880 VSS.n7077 VSS.n7076 0.04025
R11881 VSS.n7076 VSS.n7075 0.04025
R11882 VSS.n7075 VSS.n2208 0.04025
R11883 VSS.n7071 VSS.n2208 0.04025
R11884 VSS.n7071 VSS.n7070 0.04025
R11885 VSS.n7070 VSS.n7069 0.04025
R11886 VSS.n7069 VSS.n2210 0.04025
R11887 VSS.n7065 VSS.n2210 0.04025
R11888 VSS.n7065 VSS.n7064 0.04025
R11889 VSS.n7064 VSS.n7063 0.04025
R11890 VSS.n7063 VSS.n2212 0.04025
R11891 VSS.n7059 VSS.n2212 0.04025
R11892 VSS.n7059 VSS.n7058 0.04025
R11893 VSS.n7058 VSS.n7057 0.04025
R11894 VSS.n7057 VSS.n2214 0.04025
R11895 VSS.n7053 VSS.n2214 0.04025
R11896 VSS.n7053 VSS.n7052 0.04025
R11897 VSS.n7052 VSS.n7051 0.04025
R11898 VSS.n7051 VSS.n2216 0.04025
R11899 VSS.n7047 VSS.n2216 0.04025
R11900 VSS.n7047 VSS.n7046 0.04025
R11901 VSS.n7046 VSS.n7045 0.04025
R11902 VSS.n7045 VSS.n2218 0.04025
R11903 VSS.n7041 VSS.n2218 0.04025
R11904 VSS.n7041 VSS.n7040 0.04025
R11905 VSS.n7040 VSS.n7039 0.04025
R11906 VSS.n7039 VSS.n2220 0.04025
R11907 VSS.n7035 VSS.n2220 0.04025
R11908 VSS.n7035 VSS.n7034 0.04025
R11909 VSS.n7034 VSS.n7033 0.04025
R11910 VSS.n7033 VSS.n2222 0.04025
R11911 VSS.n7029 VSS.n2222 0.04025
R11912 VSS.n7029 VSS.n7028 0.04025
R11913 VSS.n7028 VSS.n7027 0.04025
R11914 VSS.n7027 VSS.n2224 0.04025
R11915 VSS.n7023 VSS.n2224 0.04025
R11916 VSS.n7023 VSS.n7022 0.04025
R11917 VSS.n7022 VSS.n7021 0.04025
R11918 VSS.n7021 VSS.n2226 0.04025
R11919 VSS.n7017 VSS.n2226 0.04025
R11920 VSS.n7017 VSS.n7016 0.04025
R11921 VSS.n7016 VSS.n7015 0.04025
R11922 VSS.n7015 VSS.n2228 0.04025
R11923 VSS.n7011 VSS.n2228 0.04025
R11924 VSS.n7011 VSS.n7010 0.04025
R11925 VSS.n7010 VSS.n7009 0.04025
R11926 VSS.n7009 VSS.n2230 0.04025
R11927 VSS.n7005 VSS.n2230 0.04025
R11928 VSS.n7005 VSS.n7004 0.04025
R11929 VSS.n7004 VSS.n7003 0.04025
R11930 VSS.n7003 VSS.n2232 0.04025
R11931 VSS.n6999 VSS.n2232 0.04025
R11932 VSS.n6999 VSS.n6998 0.04025
R11933 VSS.n6998 VSS.n6997 0.04025
R11934 VSS.n6997 VSS.n2234 0.04025
R11935 VSS.n6993 VSS.n2234 0.04025
R11936 VSS.n6993 VSS.n6992 0.04025
R11937 VSS.n6992 VSS.n6991 0.04025
R11938 VSS.n6991 VSS.n2236 0.04025
R11939 VSS.n6987 VSS.n2236 0.04025
R11940 VSS.n6987 VSS.n6986 0.04025
R11941 VSS.n6986 VSS.n6985 0.04025
R11942 VSS.n6985 VSS.n2238 0.04025
R11943 VSS.n6981 VSS.n2238 0.04025
R11944 VSS.n6981 VSS.n6980 0.04025
R11945 VSS.n6980 VSS.n6979 0.04025
R11946 VSS.n6979 VSS.n2240 0.04025
R11947 VSS.n6975 VSS.n2240 0.04025
R11948 VSS.n6975 VSS.n6974 0.04025
R11949 VSS.n6974 VSS.n6973 0.04025
R11950 VSS.n6973 VSS.n2242 0.04025
R11951 VSS.n6969 VSS.n2242 0.04025
R11952 VSS.n6969 VSS.n6968 0.04025
R11953 VSS.n6968 VSS.n6967 0.04025
R11954 VSS.n6967 VSS.n2244 0.04025
R11955 VSS.n6963 VSS.n2244 0.04025
R11956 VSS.n6963 VSS.n6962 0.04025
R11957 VSS.n6962 VSS.n6961 0.04025
R11958 VSS.n6961 VSS.n2246 0.04025
R11959 VSS.n6957 VSS.n2246 0.04025
R11960 VSS.n6957 VSS.n6956 0.04025
R11961 VSS.n6956 VSS.n6955 0.04025
R11962 VSS.n6955 VSS.n2248 0.04025
R11963 VSS.n6951 VSS.n2248 0.04025
R11964 VSS.n6951 VSS.n6950 0.04025
R11965 VSS.n6950 VSS.n6949 0.04025
R11966 VSS.n6949 VSS.n2250 0.04025
R11967 VSS.n6945 VSS.n2250 0.04025
R11968 VSS.n6945 VSS.n6944 0.04025
R11969 VSS.n6944 VSS.n6943 0.04025
R11970 VSS.n6943 VSS.n2252 0.04025
R11971 VSS.n6939 VSS.n2252 0.04025
R11972 VSS.n6939 VSS.n6938 0.04025
R11973 VSS.n6938 VSS.n6937 0.04025
R11974 VSS.n6937 VSS.n2254 0.04025
R11975 VSS.n6933 VSS.n2254 0.04025
R11976 VSS.n6933 VSS.n6932 0.04025
R11977 VSS.n6932 VSS.n6931 0.04025
R11978 VSS.n6931 VSS.n2256 0.04025
R11979 VSS.n6927 VSS.n2256 0.04025
R11980 VSS.n6927 VSS.n6926 0.04025
R11981 VSS.n6926 VSS.n6925 0.04025
R11982 VSS.n6925 VSS.n2258 0.04025
R11983 VSS.n6921 VSS.n2258 0.04025
R11984 VSS.n6921 VSS.n6920 0.04025
R11985 VSS.n6920 VSS.n6919 0.04025
R11986 VSS.n6919 VSS.n2260 0.04025
R11987 VSS.n6915 VSS.n2260 0.04025
R11988 VSS.n6915 VSS.n6914 0.04025
R11989 VSS.n6914 VSS.n6913 0.04025
R11990 VSS.n6913 VSS.n2262 0.04025
R11991 VSS.n6909 VSS.n2262 0.04025
R11992 VSS.n6909 VSS.n6908 0.04025
R11993 VSS.n4140 VSS.n4139 0.04025
R11994 VSS.n4139 VSS.n4138 0.04025
R11995 VSS.n4138 VSS.n3186 0.04025
R11996 VSS.n4134 VSS.n3186 0.04025
R11997 VSS.n4134 VSS.n4133 0.04025
R11998 VSS.n4133 VSS.n4132 0.04025
R11999 VSS.n4132 VSS.n3188 0.04025
R12000 VSS.n4128 VSS.n3188 0.04025
R12001 VSS.n4128 VSS.n4127 0.04025
R12002 VSS.n4127 VSS.n4126 0.04025
R12003 VSS.n4126 VSS.n3190 0.04025
R12004 VSS.n4122 VSS.n3190 0.04025
R12005 VSS.n4122 VSS.n4121 0.04025
R12006 VSS.n4121 VSS.n4120 0.04025
R12007 VSS.n4120 VSS.n3192 0.04025
R12008 VSS.n4116 VSS.n3192 0.04025
R12009 VSS.n4116 VSS.n4115 0.04025
R12010 VSS.n4115 VSS.n4114 0.04025
R12011 VSS.n4114 VSS.n3194 0.04025
R12012 VSS.n4110 VSS.n3194 0.04025
R12013 VSS.n4110 VSS.n4109 0.04025
R12014 VSS.n4109 VSS.n4108 0.04025
R12015 VSS.n4108 VSS.n3196 0.04025
R12016 VSS.n4104 VSS.n3196 0.04025
R12017 VSS.n4104 VSS.n4103 0.04025
R12018 VSS.n4103 VSS.n4102 0.04025
R12019 VSS.n4102 VSS.n3198 0.04025
R12020 VSS.n4098 VSS.n3198 0.04025
R12021 VSS.n4098 VSS.n4097 0.04025
R12022 VSS.n4097 VSS.n4096 0.04025
R12023 VSS.n4096 VSS.n3200 0.04025
R12024 VSS.n4092 VSS.n3200 0.04025
R12025 VSS.n4092 VSS.n4091 0.04025
R12026 VSS.n4091 VSS.n4090 0.04025
R12027 VSS.n4090 VSS.n3202 0.04025
R12028 VSS.n4086 VSS.n3202 0.04025
R12029 VSS.n4086 VSS.n4085 0.04025
R12030 VSS.n4085 VSS.n4084 0.04025
R12031 VSS.n4084 VSS.n3204 0.04025
R12032 VSS.n4080 VSS.n3204 0.04025
R12033 VSS.n4080 VSS.n4079 0.04025
R12034 VSS.n4079 VSS.n4078 0.04025
R12035 VSS.n4078 VSS.n3206 0.04025
R12036 VSS.n4074 VSS.n3206 0.04025
R12037 VSS.n4074 VSS.n4073 0.04025
R12038 VSS.n4073 VSS.n4072 0.04025
R12039 VSS.n4072 VSS.n3208 0.04025
R12040 VSS.n4068 VSS.n3208 0.04025
R12041 VSS.n4068 VSS.n4067 0.04025
R12042 VSS.n4067 VSS.n4066 0.04025
R12043 VSS.n4066 VSS.n3210 0.04025
R12044 VSS.n4062 VSS.n3210 0.04025
R12045 VSS.n4062 VSS.n4061 0.04025
R12046 VSS.n4061 VSS.n4060 0.04025
R12047 VSS.n4060 VSS.n3212 0.04025
R12048 VSS.n4056 VSS.n3212 0.04025
R12049 VSS.n4056 VSS.n4055 0.04025
R12050 VSS.n4055 VSS.n4054 0.04025
R12051 VSS.n4054 VSS.n3214 0.04025
R12052 VSS.n4050 VSS.n3214 0.04025
R12053 VSS.n4050 VSS.n4049 0.04025
R12054 VSS.n4049 VSS.n4048 0.04025
R12055 VSS.n4048 VSS.n3216 0.04025
R12056 VSS.n4044 VSS.n3216 0.04025
R12057 VSS.n4044 VSS.n4043 0.04025
R12058 VSS.n4043 VSS.n4042 0.04025
R12059 VSS.n4042 VSS.n3218 0.04025
R12060 VSS.n4038 VSS.n3218 0.04025
R12061 VSS.n4038 VSS.n4037 0.04025
R12062 VSS.n4037 VSS.n4036 0.04025
R12063 VSS.n4036 VSS.n3220 0.04025
R12064 VSS.n4032 VSS.n3220 0.04025
R12065 VSS.n4032 VSS.n4031 0.04025
R12066 VSS.n4031 VSS.n4030 0.04025
R12067 VSS.n4030 VSS.n3222 0.04025
R12068 VSS.n4026 VSS.n3222 0.04025
R12069 VSS.n4026 VSS.n4025 0.04025
R12070 VSS.n4025 VSS.n4024 0.04025
R12071 VSS.n4024 VSS.n3224 0.04025
R12072 VSS.n4020 VSS.n3224 0.04025
R12073 VSS.n4020 VSS.n4019 0.04025
R12074 VSS.n4019 VSS.n4018 0.04025
R12075 VSS.n4018 VSS.n3226 0.04025
R12076 VSS.n4014 VSS.n3226 0.04025
R12077 VSS.n4014 VSS.n4013 0.04025
R12078 VSS.n4013 VSS.n4012 0.04025
R12079 VSS.n4012 VSS.n3228 0.04025
R12080 VSS.n4008 VSS.n3228 0.04025
R12081 VSS.n4008 VSS.n4007 0.04025
R12082 VSS.n4007 VSS.n4006 0.04025
R12083 VSS.n4006 VSS.n3230 0.04025
R12084 VSS.n4002 VSS.n3230 0.04025
R12085 VSS.n4002 VSS.n4001 0.04025
R12086 VSS.n4001 VSS.n4000 0.04025
R12087 VSS.n4000 VSS.n3232 0.04025
R12088 VSS.n3996 VSS.n3232 0.04025
R12089 VSS.n3996 VSS.n3995 0.04025
R12090 VSS.n3995 VSS.n3994 0.04025
R12091 VSS.n3994 VSS.n3234 0.04025
R12092 VSS.n3990 VSS.n3234 0.04025
R12093 VSS.n3990 VSS.n3989 0.04025
R12094 VSS.n3989 VSS.n3988 0.04025
R12095 VSS.n3988 VSS.n3236 0.04025
R12096 VSS.n3984 VSS.n3236 0.04025
R12097 VSS.n3984 VSS.n3983 0.04025
R12098 VSS.n3983 VSS.n3982 0.04025
R12099 VSS.n3982 VSS.n3238 0.04025
R12100 VSS.n3978 VSS.n3238 0.04025
R12101 VSS.n3978 VSS.n3977 0.04025
R12102 VSS.n3977 VSS.n3976 0.04025
R12103 VSS.n3976 VSS.n3240 0.04025
R12104 VSS.n3972 VSS.n3240 0.04025
R12105 VSS.n3972 VSS.n3971 0.04025
R12106 VSS.n3971 VSS.n3970 0.04025
R12107 VSS.n3970 VSS.n3242 0.04025
R12108 VSS.n3966 VSS.n3242 0.04025
R12109 VSS.n3966 VSS.n3965 0.04025
R12110 VSS.n3965 VSS.n3964 0.04025
R12111 VSS.n3964 VSS.n3244 0.04025
R12112 VSS.n3960 VSS.n3244 0.04025
R12113 VSS.n3960 VSS.n3959 0.04025
R12114 VSS.n3959 VSS.n3958 0.04025
R12115 VSS.n3958 VSS.n3246 0.04025
R12116 VSS.n3954 VSS.n3246 0.04025
R12117 VSS.n3954 VSS.n3953 0.04025
R12118 VSS.n3953 VSS.n3952 0.04025
R12119 VSS.n3952 VSS.n3248 0.04025
R12120 VSS.n3948 VSS.n3248 0.04025
R12121 VSS.n3948 VSS.n3947 0.04025
R12122 VSS.n3947 VSS.n3946 0.04025
R12123 VSS.n3946 VSS.n3250 0.04025
R12124 VSS.n3942 VSS.n3250 0.04025
R12125 VSS.n3942 VSS.n3941 0.04025
R12126 VSS.n3941 VSS.n3940 0.04025
R12127 VSS.n3940 VSS.n3252 0.04025
R12128 VSS.n3936 VSS.n3252 0.04025
R12129 VSS.n3936 VSS.n3935 0.04025
R12130 VSS.n3935 VSS.n3934 0.04025
R12131 VSS.n3934 VSS.n3254 0.04025
R12132 VSS.n3930 VSS.n3254 0.04025
R12133 VSS.n3930 VSS.n3929 0.04025
R12134 VSS.n3929 VSS.n3928 0.04025
R12135 VSS.n3928 VSS.n3256 0.04025
R12136 VSS.n3924 VSS.n3256 0.04025
R12137 VSS.n3924 VSS.n3923 0.04025
R12138 VSS.n3923 VSS.n3922 0.04025
R12139 VSS.n3922 VSS.n3258 0.04025
R12140 VSS.n3918 VSS.n3258 0.04025
R12141 VSS.n3918 VSS.n3917 0.04025
R12142 VSS.n3917 VSS.n3916 0.04025
R12143 VSS.n3916 VSS.n3260 0.04025
R12144 VSS.n3912 VSS.n3260 0.04025
R12145 VSS.n3912 VSS.n3911 0.04025
R12146 VSS.n3911 VSS.n3910 0.04025
R12147 VSS.n3910 VSS.n3262 0.04025
R12148 VSS.n3906 VSS.n3262 0.04025
R12149 VSS.n3906 VSS.n3905 0.04025
R12150 VSS.n3905 VSS.n3904 0.04025
R12151 VSS.n3904 VSS.n3264 0.04025
R12152 VSS.n3900 VSS.n3264 0.04025
R12153 VSS.n3900 VSS.n3899 0.04025
R12154 VSS.n3899 VSS.n3898 0.04025
R12155 VSS.n3898 VSS.n3266 0.04025
R12156 VSS.n3894 VSS.n3266 0.04025
R12157 VSS.n3894 VSS.n3893 0.04025
R12158 VSS.n3893 VSS.n3892 0.04025
R12159 VSS.n3892 VSS.n3268 0.04025
R12160 VSS.n3888 VSS.n3268 0.04025
R12161 VSS.n3888 VSS.n3887 0.04025
R12162 VSS.n3887 VSS.n3886 0.04025
R12163 VSS.n3886 VSS.n3270 0.04025
R12164 VSS.n3882 VSS.n3270 0.04025
R12165 VSS.n3882 VSS.n3881 0.04025
R12166 VSS.n3881 VSS.n3880 0.04025
R12167 VSS.n3880 VSS.n3272 0.04025
R12168 VSS.n3876 VSS.n3272 0.04025
R12169 VSS.n3876 VSS.n3875 0.04025
R12170 VSS.n3875 VSS.n3874 0.04025
R12171 VSS.n3874 VSS.n3274 0.04025
R12172 VSS.n3870 VSS.n3274 0.04025
R12173 VSS.n3870 VSS.n3869 0.04025
R12174 VSS.n3869 VSS.n3868 0.04025
R12175 VSS.n3868 VSS.n3276 0.04025
R12176 VSS.n3864 VSS.n3276 0.04025
R12177 VSS.n3864 VSS.n3863 0.04025
R12178 VSS.n3863 VSS.n3862 0.04025
R12179 VSS.n3862 VSS.n3278 0.04025
R12180 VSS.n3858 VSS.n3278 0.04025
R12181 VSS.n3858 VSS.n3857 0.04025
R12182 VSS.n3857 VSS.n3856 0.04025
R12183 VSS.n3856 VSS.n3280 0.04025
R12184 VSS.n3852 VSS.n3280 0.04025
R12185 VSS.n3852 VSS.n3851 0.04025
R12186 VSS.n3851 VSS.n3850 0.04025
R12187 VSS.n3850 VSS.n3282 0.04025
R12188 VSS.n3846 VSS.n3282 0.04025
R12189 VSS.n3846 VSS.n3845 0.04025
R12190 VSS.n3845 VSS.n3844 0.04025
R12191 VSS.n3844 VSS.n3284 0.04025
R12192 VSS.n3840 VSS.n3284 0.04025
R12193 VSS.n3840 VSS.n3839 0.04025
R12194 VSS.n3839 VSS.n3838 0.04025
R12195 VSS.n3838 VSS.n3286 0.04025
R12196 VSS.n3834 VSS.n3286 0.04025
R12197 VSS.n3834 VSS.n3833 0.04025
R12198 VSS.n3833 VSS.n3832 0.04025
R12199 VSS.n3832 VSS.n3288 0.04025
R12200 VSS.n3828 VSS.n3288 0.04025
R12201 VSS.n3828 VSS.n3827 0.04025
R12202 VSS.n3827 VSS.n3826 0.04025
R12203 VSS.n3826 VSS.n3290 0.04025
R12204 VSS.n3822 VSS.n3290 0.04025
R12205 VSS.n3822 VSS.n3821 0.04025
R12206 VSS.n3821 VSS.n3820 0.04025
R12207 VSS.n3820 VSS.n3292 0.04025
R12208 VSS.n3816 VSS.n3292 0.04025
R12209 VSS.n3816 VSS.n3815 0.04025
R12210 VSS.n3815 VSS.n3814 0.04025
R12211 VSS.n3814 VSS.n3294 0.04025
R12212 VSS.n3810 VSS.n3294 0.04025
R12213 VSS.n3810 VSS.n3809 0.04025
R12214 VSS.n3809 VSS.n3808 0.04025
R12215 VSS.n3808 VSS.n3296 0.04025
R12216 VSS.n3804 VSS.n3296 0.04025
R12217 VSS.n3804 VSS.n3803 0.04025
R12218 VSS.n3803 VSS.n3802 0.04025
R12219 VSS.n3802 VSS.n3298 0.04025
R12220 VSS.n3798 VSS.n3298 0.04025
R12221 VSS.n3798 VSS.n3797 0.04025
R12222 VSS.n3797 VSS.n3796 0.04025
R12223 VSS.n3796 VSS.n3300 0.04025
R12224 VSS.n3792 VSS.n3300 0.04025
R12225 VSS.n3792 VSS.n3791 0.04025
R12226 VSS.n3791 VSS.n3790 0.04025
R12227 VSS.n3790 VSS.n3302 0.04025
R12228 VSS.n3786 VSS.n3302 0.04025
R12229 VSS.n3786 VSS.n3785 0.04025
R12230 VSS.n3785 VSS.n3784 0.04025
R12231 VSS.n3784 VSS.n3304 0.04025
R12232 VSS.n3780 VSS.n3304 0.04025
R12233 VSS.n3780 VSS.n3779 0.04025
R12234 VSS.n3779 VSS.n3778 0.04025
R12235 VSS.n3778 VSS.n3306 0.04025
R12236 VSS.n3774 VSS.n3306 0.04025
R12237 VSS.n3774 VSS.n3773 0.04025
R12238 VSS.n3773 VSS.n3772 0.04025
R12239 VSS.n3772 VSS.n3308 0.04025
R12240 VSS.n3768 VSS.n3308 0.04025
R12241 VSS.n3768 VSS.n3767 0.04025
R12242 VSS.n3767 VSS.n3766 0.04025
R12243 VSS.n3766 VSS.n3310 0.04025
R12244 VSS.n3762 VSS.n3310 0.04025
R12245 VSS.n3762 VSS.n3761 0.04025
R12246 VSS.n3761 VSS.n3760 0.04025
R12247 VSS.n3760 VSS.n3312 0.04025
R12248 VSS.n3756 VSS.n3312 0.04025
R12249 VSS.n3756 VSS.n3755 0.04025
R12250 VSS.n3755 VSS.n3754 0.04025
R12251 VSS.n3754 VSS.n3314 0.04025
R12252 VSS.n3750 VSS.n3314 0.04025
R12253 VSS.n3750 VSS.n3749 0.04025
R12254 VSS.n3749 VSS.n3748 0.04025
R12255 VSS.n3748 VSS.n3316 0.04025
R12256 VSS.n3744 VSS.n3316 0.04025
R12257 VSS.n3744 VSS.n3743 0.04025
R12258 VSS.n3743 VSS.n3742 0.04025
R12259 VSS.n3742 VSS.n3318 0.04025
R12260 VSS.n3738 VSS.n3318 0.04025
R12261 VSS.n3738 VSS.n3737 0.04025
R12262 VSS.n3737 VSS.n3736 0.04025
R12263 VSS.n3736 VSS.n3320 0.04025
R12264 VSS.n3732 VSS.n3320 0.04025
R12265 VSS.n3732 VSS.n3731 0.04025
R12266 VSS.n3731 VSS.n3730 0.04025
R12267 VSS.n3730 VSS.n3322 0.04025
R12268 VSS.n3726 VSS.n3322 0.04025
R12269 VSS.n3726 VSS.n3725 0.04025
R12270 VSS.n3725 VSS.n3724 0.04025
R12271 VSS.n3724 VSS.n3324 0.04025
R12272 VSS.n3720 VSS.n3324 0.04025
R12273 VSS.n3720 VSS.n3719 0.04025
R12274 VSS.n3719 VSS.n3718 0.04025
R12275 VSS.n3718 VSS.n3326 0.04025
R12276 VSS.n3714 VSS.n3326 0.04025
R12277 VSS.n3714 VSS.n3713 0.04025
R12278 VSS.n3713 VSS.n3712 0.04025
R12279 VSS.n3712 VSS.n3328 0.04025
R12280 VSS.n3708 VSS.n3328 0.04025
R12281 VSS.n3708 VSS.n3707 0.04025
R12282 VSS.n3707 VSS.n3706 0.04025
R12283 VSS.n3706 VSS.n3330 0.04025
R12284 VSS.n3702 VSS.n3330 0.04025
R12285 VSS.n3702 VSS.n3701 0.04025
R12286 VSS.n3701 VSS.n3700 0.04025
R12287 VSS.n3700 VSS.n3332 0.04025
R12288 VSS.n3696 VSS.n3332 0.04025
R12289 VSS.n3696 VSS.n3695 0.04025
R12290 VSS.n3695 VSS.n3694 0.04025
R12291 VSS.n3694 VSS.n3334 0.04025
R12292 VSS.n3690 VSS.n3334 0.04025
R12293 VSS.n3690 VSS.n3689 0.04025
R12294 VSS.n3689 VSS.n3688 0.04025
R12295 VSS.n3688 VSS.n3336 0.04025
R12296 VSS.n3684 VSS.n3336 0.04025
R12297 VSS.n3684 VSS.n3683 0.04025
R12298 VSS.n3683 VSS.n3682 0.04025
R12299 VSS.n3682 VSS.n3338 0.04025
R12300 VSS.n3678 VSS.n3338 0.04025
R12301 VSS.n3678 VSS.n3677 0.04025
R12302 VSS.n3677 VSS.n3676 0.04025
R12303 VSS.n3676 VSS.n3340 0.04025
R12304 VSS.n3672 VSS.n3340 0.04025
R12305 VSS.n3672 VSS.n3671 0.04025
R12306 VSS.n3671 VSS.n3670 0.04025
R12307 VSS.n3670 VSS.n3342 0.04025
R12308 VSS.n3666 VSS.n3342 0.04025
R12309 VSS.n3666 VSS.n3665 0.04025
R12310 VSS.n3665 VSS.n3664 0.04025
R12311 VSS.n3664 VSS.n3344 0.04025
R12312 VSS.n3660 VSS.n3344 0.04025
R12313 VSS.n3660 VSS.n3659 0.04025
R12314 VSS.n3659 VSS.n3658 0.04025
R12315 VSS.n3658 VSS.n3346 0.04025
R12316 VSS.n3654 VSS.n3346 0.04025
R12317 VSS.n3654 VSS.n3653 0.04025
R12318 VSS.n3653 VSS.n3652 0.04025
R12319 VSS.n3652 VSS.n3348 0.04025
R12320 VSS.n3648 VSS.n3348 0.04025
R12321 VSS.n3648 VSS.n3647 0.04025
R12322 VSS.n3647 VSS.n3646 0.04025
R12323 VSS.n3646 VSS.n3350 0.04025
R12324 VSS.n3642 VSS.n3350 0.04025
R12325 VSS.n3642 VSS.n3641 0.04025
R12326 VSS.n3641 VSS.n3640 0.04025
R12327 VSS.n3640 VSS.n3352 0.04025
R12328 VSS.n3636 VSS.n3352 0.04025
R12329 VSS.n3636 VSS.n3635 0.04025
R12330 VSS.n3635 VSS.n3634 0.04025
R12331 VSS.n3634 VSS.n3354 0.04025
R12332 VSS.n3630 VSS.n3354 0.04025
R12333 VSS.n3630 VSS.n3629 0.04025
R12334 VSS.n3629 VSS.n3628 0.04025
R12335 VSS.n3628 VSS.n3356 0.04025
R12336 VSS.n3624 VSS.n3356 0.04025
R12337 VSS.n3624 VSS.n3623 0.04025
R12338 VSS.n3623 VSS.n3622 0.04025
R12339 VSS.n3622 VSS.n3358 0.04025
R12340 VSS.n3618 VSS.n3358 0.04025
R12341 VSS.n3618 VSS.n3617 0.04025
R12342 VSS.n3617 VSS.n3616 0.04025
R12343 VSS.n3616 VSS.n3360 0.04025
R12344 VSS.n3612 VSS.n3360 0.04025
R12345 VSS.n3612 VSS.n3611 0.04025
R12346 VSS.n3611 VSS.n3610 0.04025
R12347 VSS.n3610 VSS.n3362 0.04025
R12348 VSS.n3606 VSS.n3362 0.04025
R12349 VSS.n3606 VSS.n3605 0.04025
R12350 VSS.n3605 VSS.n3604 0.04025
R12351 VSS.n3604 VSS.n3364 0.04025
R12352 VSS.n3600 VSS.n3364 0.04025
R12353 VSS.n3600 VSS.n3599 0.04025
R12354 VSS.n3599 VSS.n3598 0.04025
R12355 VSS.n3598 VSS.n3366 0.04025
R12356 VSS.n3594 VSS.n3366 0.04025
R12357 VSS.n3594 VSS.n3593 0.04025
R12358 VSS.n3593 VSS.n3592 0.04025
R12359 VSS.n3592 VSS.n3368 0.04025
R12360 VSS.n3588 VSS.n3368 0.04025
R12361 VSS.n3588 VSS.n3587 0.04025
R12362 VSS.n3587 VSS.n3586 0.04025
R12363 VSS.n3586 VSS.n3370 0.04025
R12364 VSS.n3582 VSS.n3370 0.04025
R12365 VSS.n3582 VSS.n3581 0.04025
R12366 VSS.n3581 VSS.n3580 0.04025
R12367 VSS.n3580 VSS.n3372 0.04025
R12368 VSS.n3576 VSS.n3372 0.04025
R12369 VSS.n3576 VSS.n3575 0.04025
R12370 VSS.n3575 VSS.n3574 0.04025
R12371 VSS.n3574 VSS.n3374 0.04025
R12372 VSS.n3570 VSS.n3374 0.04025
R12373 VSS.n3570 VSS.n3569 0.04025
R12374 VSS.n3569 VSS.n3568 0.04025
R12375 VSS.n3568 VSS.n3376 0.04025
R12376 VSS.n3564 VSS.n3376 0.04025
R12377 VSS.n3564 VSS.n3563 0.04025
R12378 VSS.n3563 VSS.n3562 0.04025
R12379 VSS.n3562 VSS.n3378 0.04025
R12380 VSS.n3558 VSS.n3378 0.04025
R12381 VSS.n3558 VSS.n3557 0.04025
R12382 VSS.n3557 VSS.n3556 0.04025
R12383 VSS.n3556 VSS.n3380 0.04025
R12384 VSS.n3552 VSS.n3380 0.04025
R12385 VSS.n3552 VSS.n3551 0.04025
R12386 VSS.n3551 VSS.n3550 0.04025
R12387 VSS.n3550 VSS.n3382 0.04025
R12388 VSS.n3546 VSS.n3382 0.04025
R12389 VSS.n3546 VSS.n3545 0.04025
R12390 VSS.n3545 VSS.n3544 0.04025
R12391 VSS.n3544 VSS.n3384 0.04025
R12392 VSS.n3540 VSS.n3384 0.04025
R12393 VSS.n3540 VSS.n3539 0.04025
R12394 VSS.n3539 VSS.n3538 0.04025
R12395 VSS.n3538 VSS.n3386 0.04025
R12396 VSS.n3534 VSS.n3386 0.04025
R12397 VSS.n3534 VSS.n3533 0.04025
R12398 VSS.n3533 VSS.n3532 0.04025
R12399 VSS.n3532 VSS.n3388 0.04025
R12400 VSS.n3528 VSS.n3388 0.04025
R12401 VSS.n3528 VSS.n3527 0.04025
R12402 VSS.n3527 VSS.n3526 0.04025
R12403 VSS.n3526 VSS.n3390 0.04025
R12404 VSS.n3522 VSS.n3390 0.04025
R12405 VSS.n3522 VSS.n3521 0.04025
R12406 VSS.n3521 VSS.n3520 0.04025
R12407 VSS.n3520 VSS.n3392 0.04025
R12408 VSS.n3516 VSS.n3392 0.04025
R12409 VSS.n3516 VSS.n3515 0.04025
R12410 VSS.n3515 VSS.n3514 0.04025
R12411 VSS.n3514 VSS.n3394 0.04025
R12412 VSS.n3510 VSS.n3394 0.04025
R12413 VSS.n3510 VSS.n3509 0.04025
R12414 VSS.n3509 VSS.n3508 0.04025
R12415 VSS.n3508 VSS.n3396 0.04025
R12416 VSS.n3504 VSS.n3396 0.04025
R12417 VSS.n3504 VSS.n3503 0.04025
R12418 VSS.n3503 VSS.n3502 0.04025
R12419 VSS.n3502 VSS.n3398 0.04025
R12420 VSS.n3498 VSS.n3398 0.04025
R12421 VSS.n3498 VSS.n3497 0.04025
R12422 VSS.n3497 VSS.n3496 0.04025
R12423 VSS.n3496 VSS.n3400 0.04025
R12424 VSS.n3492 VSS.n3400 0.04025
R12425 VSS.n3492 VSS.n3491 0.04025
R12426 VSS.n3491 VSS.n3490 0.04025
R12427 VSS.n3490 VSS.n3402 0.04025
R12428 VSS.n3486 VSS.n3402 0.04025
R12429 VSS.n3486 VSS.n3485 0.04025
R12430 VSS.n3485 VSS.n3484 0.04025
R12431 VSS.n3484 VSS.n3404 0.04025
R12432 VSS.n3480 VSS.n3404 0.04025
R12433 VSS.n3480 VSS.n3479 0.04025
R12434 VSS.n3479 VSS.n3478 0.04025
R12435 VSS.n3478 VSS.n3406 0.04025
R12436 VSS.n3474 VSS.n3406 0.04025
R12437 VSS.n3474 VSS.n3473 0.04025
R12438 VSS.n3473 VSS.n3472 0.04025
R12439 VSS.n3472 VSS.n3408 0.04025
R12440 VSS.n3468 VSS.n3408 0.04025
R12441 VSS.n3468 VSS.n3467 0.04025
R12442 VSS.n3467 VSS.n3466 0.04025
R12443 VSS.n3466 VSS.n3410 0.04025
R12444 VSS.n3462 VSS.n3410 0.04025
R12445 VSS.n3462 VSS.n3461 0.04025
R12446 VSS.n3461 VSS.n3460 0.04025
R12447 VSS.n3460 VSS.n3412 0.04025
R12448 VSS.n3456 VSS.n3412 0.04025
R12449 VSS.n3456 VSS.n3455 0.04025
R12450 VSS.n3455 VSS.n3454 0.04025
R12451 VSS.n3454 VSS.n3414 0.04025
R12452 VSS.n3450 VSS.n3414 0.04025
R12453 VSS.n3450 VSS.n3449 0.04025
R12454 VSS.n3449 VSS.n3448 0.04025
R12455 VSS.n3448 VSS.n3416 0.04025
R12456 VSS.n3444 VSS.n3416 0.04025
R12457 VSS.n3444 VSS.n3443 0.04025
R12458 VSS.n3443 VSS.n3442 0.04025
R12459 VSS.n3442 VSS.n3418 0.04025
R12460 VSS.n3438 VSS.n3418 0.04025
R12461 VSS.n3438 VSS.n3437 0.04025
R12462 VSS.n3437 VSS.n3436 0.04025
R12463 VSS.n3436 VSS.n3420 0.04025
R12464 VSS.n3432 VSS.n3420 0.04025
R12465 VSS.n3432 VSS.n3431 0.04025
R12466 VSS.n3431 VSS.n3430 0.04025
R12467 VSS.n3430 VSS.n3422 0.04025
R12468 VSS.n3426 VSS.n3422 0.04025
R12469 VSS.n3426 VSS.n3425 0.04025
R12470 VSS.n3425 VSS.n3424 0.04025
R12471 VSS.n3424 VSS.n1582 0.04025
R12472 VSS.n8949 VSS.n1582 0.04025
R12473 VSS.n8949 VSS.n8948 0.04025
R12474 VSS.n8948 VSS.n8947 0.04025
R12475 VSS.n8947 VSS.n1584 0.04025
R12476 VSS.n8943 VSS.n1584 0.04025
R12477 VSS.n8943 VSS.n8942 0.04025
R12478 VSS.n8942 VSS.n8941 0.04025
R12479 VSS.n8941 VSS.n1586 0.04025
R12480 VSS.n8937 VSS.n1586 0.04025
R12481 VSS.n8937 VSS.n8936 0.04025
R12482 VSS.n8936 VSS.n8935 0.04025
R12483 VSS.n8935 VSS.n1588 0.04025
R12484 VSS.n8931 VSS.n1588 0.04025
R12485 VSS.n8931 VSS.n8930 0.04025
R12486 VSS.n8930 VSS.n8929 0.04025
R12487 VSS.n8929 VSS.n1590 0.04025
R12488 VSS.n8925 VSS.n1590 0.04025
R12489 VSS.n8925 VSS.n8924 0.04025
R12490 VSS.n8924 VSS.n8923 0.04025
R12491 VSS.n8923 VSS.n1592 0.04025
R12492 VSS.n8919 VSS.n1592 0.04025
R12493 VSS.n8919 VSS.n8918 0.04025
R12494 VSS.n8918 VSS.n8917 0.04025
R12495 VSS.n8917 VSS.n1594 0.04025
R12496 VSS.n8913 VSS.n1594 0.04025
R12497 VSS.n8913 VSS.n8912 0.04025
R12498 VSS.n8912 VSS.n8911 0.04025
R12499 VSS.n8911 VSS.n1596 0.04025
R12500 VSS.n8907 VSS.n1596 0.04025
R12501 VSS.n8907 VSS.n8906 0.04025
R12502 VSS.n8906 VSS.n8905 0.04025
R12503 VSS.n8905 VSS.n1598 0.04025
R12504 VSS.n8901 VSS.n1598 0.04025
R12505 VSS.n8901 VSS.n8900 0.04025
R12506 VSS.n8900 VSS.n8899 0.04025
R12507 VSS.n8899 VSS.n1600 0.04025
R12508 VSS.n8895 VSS.n1600 0.04025
R12509 VSS.n8895 VSS.n8894 0.04025
R12510 VSS.n8894 VSS.n8893 0.04025
R12511 VSS.n8893 VSS.n1602 0.04025
R12512 VSS.n8889 VSS.n1602 0.04025
R12513 VSS.n8889 VSS.n8888 0.04025
R12514 VSS.n8888 VSS.n8887 0.04025
R12515 VSS.n8887 VSS.n1604 0.04025
R12516 VSS.n8883 VSS.n1604 0.04025
R12517 VSS.n8883 VSS.n8882 0.04025
R12518 VSS.n8882 VSS.n8881 0.04025
R12519 VSS.n8881 VSS.n1606 0.04025
R12520 VSS.n8877 VSS.n1606 0.04025
R12521 VSS.n8877 VSS.n8876 0.04025
R12522 VSS.n8876 VSS.n8875 0.04025
R12523 VSS.n8875 VSS.n1608 0.04025
R12524 VSS.n8871 VSS.n1608 0.04025
R12525 VSS.n8871 VSS.n8870 0.04025
R12526 VSS.n8870 VSS.n8869 0.04025
R12527 VSS.n8869 VSS.n1610 0.04025
R12528 VSS.n8865 VSS.n1610 0.04025
R12529 VSS.n8865 VSS.n8864 0.04025
R12530 VSS.n8864 VSS.n8863 0.04025
R12531 VSS.n8863 VSS.n1612 0.04025
R12532 VSS.n8859 VSS.n1612 0.04025
R12533 VSS.n8859 VSS.n8858 0.04025
R12534 VSS.n8858 VSS.n8857 0.04025
R12535 VSS.n8857 VSS.n1614 0.04025
R12536 VSS.n8853 VSS.n1614 0.04025
R12537 VSS.n8853 VSS.n8852 0.04025
R12538 VSS.n8852 VSS.n8851 0.04025
R12539 VSS.n8851 VSS.n1616 0.04025
R12540 VSS.n8847 VSS.n1616 0.04025
R12541 VSS.n8847 VSS.n8846 0.04025
R12542 VSS.n8846 VSS.n8845 0.04025
R12543 VSS.n8845 VSS.n1618 0.04025
R12544 VSS.n8841 VSS.n1618 0.04025
R12545 VSS.n8841 VSS.n8840 0.04025
R12546 VSS.n8840 VSS.n8839 0.04025
R12547 VSS.n8839 VSS.n1620 0.04025
R12548 VSS.n8835 VSS.n1620 0.04025
R12549 VSS.n8835 VSS.n8834 0.04025
R12550 VSS.n8834 VSS.n8833 0.04025
R12551 VSS.n8833 VSS.n1622 0.04025
R12552 VSS.n8829 VSS.n1622 0.04025
R12553 VSS.n8829 VSS.n8828 0.04025
R12554 VSS.n8828 VSS.n8827 0.04025
R12555 VSS.n8827 VSS.n1624 0.04025
R12556 VSS.n8823 VSS.n1624 0.04025
R12557 VSS.n8823 VSS.n8822 0.04025
R12558 VSS.n8822 VSS.n8821 0.04025
R12559 VSS.n8821 VSS.n1626 0.04025
R12560 VSS.n8817 VSS.n1626 0.04025
R12561 VSS.n8817 VSS.n8816 0.04025
R12562 VSS.n8816 VSS.n8815 0.04025
R12563 VSS.n8815 VSS.n1628 0.04025
R12564 VSS.n8811 VSS.n1628 0.04025
R12565 VSS.n8811 VSS.n8810 0.04025
R12566 VSS.n8810 VSS.n8809 0.04025
R12567 VSS.n8809 VSS.n1630 0.04025
R12568 VSS.n8805 VSS.n1630 0.04025
R12569 VSS.n8805 VSS.n8804 0.04025
R12570 VSS.n8804 VSS.n8803 0.04025
R12571 VSS.n8803 VSS.n1632 0.04025
R12572 VSS.n8799 VSS.n1632 0.04025
R12573 VSS.n8799 VSS.n8798 0.04025
R12574 VSS.n8798 VSS.n8797 0.04025
R12575 VSS.n8797 VSS.n1634 0.04025
R12576 VSS.n8793 VSS.n1634 0.04025
R12577 VSS.n8793 VSS.n8792 0.04025
R12578 VSS.n8792 VSS.n8791 0.04025
R12579 VSS.n8791 VSS.n1636 0.04025
R12580 VSS.n8787 VSS.n1636 0.04025
R12581 VSS.n8787 VSS.n8786 0.04025
R12582 VSS.n8786 VSS.n8785 0.04025
R12583 VSS.n8785 VSS.n1638 0.04025
R12584 VSS.n8781 VSS.n1638 0.04025
R12585 VSS.n8781 VSS.n8780 0.04025
R12586 VSS.n8780 VSS.n8779 0.04025
R12587 VSS.n8779 VSS.n1640 0.04025
R12588 VSS.n8775 VSS.n1640 0.04025
R12589 VSS.n8775 VSS.n8774 0.04025
R12590 VSS.n8774 VSS.n8773 0.04025
R12591 VSS.n8773 VSS.n1642 0.04025
R12592 VSS.n8769 VSS.n1642 0.04025
R12593 VSS.n8769 VSS.n8768 0.04025
R12594 VSS.n8768 VSS.n8767 0.04025
R12595 VSS.n8767 VSS.n1644 0.04025
R12596 VSS.n8763 VSS.n1644 0.04025
R12597 VSS.n8763 VSS.n8762 0.04025
R12598 VSS.n8762 VSS.n8761 0.04025
R12599 VSS.n8761 VSS.n1646 0.04025
R12600 VSS.n8757 VSS.n1646 0.04025
R12601 VSS.n8757 VSS.n8756 0.04025
R12602 VSS.n8756 VSS.n8755 0.04025
R12603 VSS.n8755 VSS.n1648 0.04025
R12604 VSS.n8751 VSS.n1648 0.04025
R12605 VSS.n8751 VSS.n8750 0.04025
R12606 VSS.n8750 VSS.n8749 0.04025
R12607 VSS.n8749 VSS.n1650 0.04025
R12608 VSS.n8745 VSS.n1650 0.04025
R12609 VSS.n8745 VSS.n8744 0.04025
R12610 VSS.n8744 VSS.n8743 0.04025
R12611 VSS.n8743 VSS.n1652 0.04025
R12612 VSS.n8739 VSS.n1652 0.04025
R12613 VSS.n8739 VSS.n8738 0.04025
R12614 VSS.n8738 VSS.n8737 0.04025
R12615 VSS.n8737 VSS.n1654 0.04025
R12616 VSS.n8733 VSS.n1654 0.04025
R12617 VSS.n8733 VSS.n8732 0.04025
R12618 VSS.n8732 VSS.n8731 0.04025
R12619 VSS.n8731 VSS.n1656 0.04025
R12620 VSS.n8727 VSS.n1656 0.04025
R12621 VSS.n8727 VSS.n8726 0.04025
R12622 VSS.n8726 VSS.n8725 0.04025
R12623 VSS.n8725 VSS.n1658 0.04025
R12624 VSS.n8721 VSS.n1658 0.04025
R12625 VSS.n8721 VSS.n8720 0.04025
R12626 VSS.n8720 VSS.n8719 0.04025
R12627 VSS.n8719 VSS.n1660 0.04025
R12628 VSS.n8715 VSS.n1660 0.04025
R12629 VSS.n8715 VSS.n8714 0.04025
R12630 VSS.n8714 VSS.n8713 0.04025
R12631 VSS.n8713 VSS.n1662 0.04025
R12632 VSS.n8709 VSS.n1662 0.04025
R12633 VSS.n8709 VSS.n8708 0.04025
R12634 VSS.n8708 VSS.n8707 0.04025
R12635 VSS.n8707 VSS.n1664 0.04025
R12636 VSS.n8703 VSS.n1664 0.04025
R12637 VSS.n8703 VSS.n8702 0.04025
R12638 VSS.n8702 VSS.n8701 0.04025
R12639 VSS.n8701 VSS.n1666 0.04025
R12640 VSS.n8697 VSS.n1666 0.04025
R12641 VSS.n8697 VSS.n8696 0.04025
R12642 VSS.n8696 VSS.n8695 0.04025
R12643 VSS.n8695 VSS.n1668 0.04025
R12644 VSS.n8691 VSS.n1668 0.04025
R12645 VSS.n8691 VSS.n8690 0.04025
R12646 VSS.n8690 VSS.n8689 0.04025
R12647 VSS.n8689 VSS.n1670 0.04025
R12648 VSS.n8685 VSS.n1670 0.04025
R12649 VSS.n8685 VSS.n8684 0.04025
R12650 VSS.n8684 VSS.n8683 0.04025
R12651 VSS.n8683 VSS.n1672 0.04025
R12652 VSS.n8679 VSS.n1672 0.04025
R12653 VSS.n8679 VSS.n8678 0.04025
R12654 VSS.n8678 VSS.n8677 0.04025
R12655 VSS.n8677 VSS.n1674 0.04025
R12656 VSS.n8673 VSS.n1674 0.04025
R12657 VSS.n8673 VSS.n8672 0.04025
R12658 VSS.n8672 VSS.n8671 0.04025
R12659 VSS.n8671 VSS.n1676 0.04025
R12660 VSS.n8667 VSS.n1676 0.04025
R12661 VSS.n8667 VSS.n8666 0.04025
R12662 VSS.n8666 VSS.n8665 0.04025
R12663 VSS.n8665 VSS.n1678 0.04025
R12664 VSS.n8661 VSS.n1678 0.04025
R12665 VSS.n8661 VSS.n8660 0.04025
R12666 VSS.n8660 VSS.n8659 0.04025
R12667 VSS.n8659 VSS.n1680 0.04025
R12668 VSS.n8655 VSS.n1680 0.04025
R12669 VSS.n8655 VSS.n8654 0.04025
R12670 VSS.n8654 VSS.n8653 0.04025
R12671 VSS.n8653 VSS.n1682 0.04025
R12672 VSS.n8649 VSS.n1682 0.04025
R12673 VSS.n8649 VSS.n8648 0.04025
R12674 VSS.n8648 VSS.n8647 0.04025
R12675 VSS.n8647 VSS.n1684 0.04025
R12676 VSS.n8643 VSS.n1684 0.04025
R12677 VSS.n8643 VSS.n8642 0.04025
R12678 VSS.n8642 VSS.n8641 0.04025
R12679 VSS.n8641 VSS.n1686 0.04025
R12680 VSS.n8637 VSS.n1686 0.04025
R12681 VSS.n8637 VSS.n8636 0.04025
R12682 VSS.n8636 VSS.n8635 0.04025
R12683 VSS.n8635 VSS.n1688 0.04025
R12684 VSS.n8631 VSS.n1688 0.04025
R12685 VSS.n8631 VSS.n8630 0.04025
R12686 VSS.n8630 VSS.n8629 0.04025
R12687 VSS.n8629 VSS.n1690 0.04025
R12688 VSS.n8625 VSS.n1690 0.04025
R12689 VSS.n8625 VSS.n8624 0.04025
R12690 VSS.n8624 VSS.n8623 0.04025
R12691 VSS.n8623 VSS.n1692 0.04025
R12692 VSS.n8619 VSS.n1692 0.04025
R12693 VSS.n8619 VSS.n8618 0.04025
R12694 VSS.n8618 VSS.n8617 0.04025
R12695 VSS.n8617 VSS.n1694 0.04025
R12696 VSS.n8613 VSS.n1694 0.04025
R12697 VSS.n8613 VSS.n8612 0.04025
R12698 VSS.n8612 VSS.n8611 0.04025
R12699 VSS.n8611 VSS.n1696 0.04025
R12700 VSS.n8607 VSS.n1696 0.04025
R12701 VSS.n8607 VSS.n8606 0.04025
R12702 VSS.n8606 VSS.n8605 0.04025
R12703 VSS.n8605 VSS.n1698 0.04025
R12704 VSS.n8601 VSS.n1698 0.04025
R12705 VSS.n8601 VSS.n8600 0.04025
R12706 VSS.n8600 VSS.n8599 0.04025
R12707 VSS.n8599 VSS.n1700 0.04025
R12708 VSS.n8595 VSS.n1700 0.04025
R12709 VSS.n8595 VSS.n8594 0.04025
R12710 VSS.n8594 VSS.n8593 0.04025
R12711 VSS.n8593 VSS.n1702 0.04025
R12712 VSS.n8589 VSS.n1702 0.04025
R12713 VSS.n8589 VSS.n8588 0.04025
R12714 VSS.n8588 VSS.n8587 0.04025
R12715 VSS.n8587 VSS.n1704 0.04025
R12716 VSS.n8583 VSS.n1704 0.04025
R12717 VSS.n8583 VSS.n8582 0.04025
R12718 VSS.n8582 VSS.n8581 0.04025
R12719 VSS.n8581 VSS.n1706 0.04025
R12720 VSS.n8577 VSS.n1706 0.04025
R12721 VSS.n8577 VSS.n8576 0.04025
R12722 VSS.n8576 VSS.n8575 0.04025
R12723 VSS.n8575 VSS.n1708 0.04025
R12724 VSS.n8571 VSS.n1708 0.04025
R12725 VSS.n8571 VSS.n8570 0.04025
R12726 VSS.n8570 VSS.n8569 0.04025
R12727 VSS.n8569 VSS.n1710 0.04025
R12728 VSS.n8565 VSS.n1710 0.04025
R12729 VSS.n8565 VSS.n8564 0.04025
R12730 VSS.n8564 VSS.n8563 0.04025
R12731 VSS.n8563 VSS.n1712 0.04025
R12732 VSS.n8559 VSS.n1712 0.04025
R12733 VSS.n8559 VSS.n8558 0.04025
R12734 VSS.n8558 VSS.n8557 0.04025
R12735 VSS.n8557 VSS.n1714 0.04025
R12736 VSS.n8553 VSS.n1714 0.04025
R12737 VSS.n8553 VSS.n8552 0.04025
R12738 VSS.n8552 VSS.n8551 0.04025
R12739 VSS.n8551 VSS.n1716 0.04025
R12740 VSS.n8547 VSS.n1716 0.04025
R12741 VSS.n8547 VSS.n8546 0.04025
R12742 VSS.n8546 VSS.n8545 0.04025
R12743 VSS.n8545 VSS.n1718 0.04025
R12744 VSS.n8541 VSS.n1718 0.04025
R12745 VSS.n8541 VSS.n8540 0.04025
R12746 VSS.n8540 VSS.n8539 0.04025
R12747 VSS.n8539 VSS.n1720 0.04025
R12748 VSS.n8535 VSS.n1720 0.04025
R12749 VSS.n8535 VSS.n8534 0.04025
R12750 VSS.n8534 VSS.n8533 0.04025
R12751 VSS.n8533 VSS.n1722 0.04025
R12752 VSS.n8529 VSS.n1722 0.04025
R12753 VSS.n8529 VSS.n8528 0.04025
R12754 VSS.n8528 VSS.n8527 0.04025
R12755 VSS.n8527 VSS.n1724 0.04025
R12756 VSS.n8523 VSS.n1724 0.04025
R12757 VSS.n8523 VSS.n8522 0.04025
R12758 VSS.n8522 VSS.n8521 0.04025
R12759 VSS.n8521 VSS.n1726 0.04025
R12760 VSS.n8517 VSS.n1726 0.04025
R12761 VSS.n8517 VSS.n8516 0.04025
R12762 VSS.n8516 VSS.n8515 0.04025
R12763 VSS.n8515 VSS.n1728 0.04025
R12764 VSS.n8511 VSS.n1728 0.04025
R12765 VSS.n8511 VSS.n8510 0.04025
R12766 VSS.n8510 VSS.n8509 0.04025
R12767 VSS.n8509 VSS.n1730 0.04025
R12768 VSS.n8505 VSS.n1730 0.04025
R12769 VSS.n8505 VSS.n8504 0.04025
R12770 VSS.n8504 VSS.n8503 0.04025
R12771 VSS.n8503 VSS.n1732 0.04025
R12772 VSS.n8499 VSS.n1732 0.04025
R12773 VSS.n8499 VSS.n8498 0.04025
R12774 VSS.n8498 VSS.n8497 0.04025
R12775 VSS.n8497 VSS.n1734 0.04025
R12776 VSS.n8493 VSS.n1734 0.04025
R12777 VSS.n8493 VSS.n8492 0.04025
R12778 VSS.n8492 VSS.n8491 0.04025
R12779 VSS.n8491 VSS.n1736 0.04025
R12780 VSS.n8487 VSS.n1736 0.04025
R12781 VSS.n8487 VSS.n8486 0.04025
R12782 VSS.n8486 VSS.n8485 0.04025
R12783 VSS.n8485 VSS.n1738 0.04025
R12784 VSS.n8481 VSS.n1738 0.04025
R12785 VSS.n8481 VSS.n8480 0.04025
R12786 VSS.n8480 VSS.n8479 0.04025
R12787 VSS.n8479 VSS.n1740 0.04025
R12788 VSS.n8475 VSS.n1740 0.04025
R12789 VSS.n8475 VSS.n8474 0.04025
R12790 VSS.n8474 VSS.n8473 0.04025
R12791 VSS.n8473 VSS.n1742 0.04025
R12792 VSS.n8469 VSS.n1742 0.04025
R12793 VSS.n8469 VSS.n8468 0.04025
R12794 VSS.n8468 VSS.n8467 0.04025
R12795 VSS.n8467 VSS.n1744 0.04025
R12796 VSS.n8463 VSS.n1744 0.04025
R12797 VSS.n8463 VSS.n8462 0.04025
R12798 VSS.n8462 VSS.n8461 0.04025
R12799 VSS.n8461 VSS.n1746 0.04025
R12800 VSS.n8457 VSS.n1746 0.04025
R12801 VSS.n8457 VSS.n8456 0.04025
R12802 VSS.n8456 VSS.n8455 0.04025
R12803 VSS.n8455 VSS.n1748 0.04025
R12804 VSS.n8451 VSS.n1748 0.04025
R12805 VSS.n8451 VSS.n8450 0.04025
R12806 VSS.n8450 VSS.n8449 0.04025
R12807 VSS.n8449 VSS.n1750 0.04025
R12808 VSS.n8445 VSS.n1750 0.04025
R12809 VSS.n8445 VSS.n8444 0.04025
R12810 VSS.n8444 VSS.n8443 0.04025
R12811 VSS.n8443 VSS.n1752 0.04025
R12812 VSS.n8439 VSS.n1752 0.04025
R12813 VSS.n8439 VSS.n8438 0.04025
R12814 VSS.n8438 VSS.n8437 0.04025
R12815 VSS.n8437 VSS.n1754 0.04025
R12816 VSS.n8433 VSS.n1754 0.04025
R12817 VSS.n8433 VSS.n8432 0.04025
R12818 VSS.n8432 VSS.n8431 0.04025
R12819 VSS.n8431 VSS.n1756 0.04025
R12820 VSS.n8427 VSS.n1756 0.04025
R12821 VSS.n8427 VSS.n8426 0.04025
R12822 VSS.n8426 VSS.n8425 0.04025
R12823 VSS.n8425 VSS.n1758 0.04025
R12824 VSS.n8421 VSS.n1758 0.04025
R12825 VSS.n8421 VSS.n8420 0.04025
R12826 VSS.n8420 VSS.n8419 0.04025
R12827 VSS.n8419 VSS.n1760 0.04025
R12828 VSS.n8415 VSS.n1760 0.04025
R12829 VSS.n8415 VSS.n8414 0.04025
R12830 VSS.n8414 VSS.n8413 0.04025
R12831 VSS.n8413 VSS.n1762 0.04025
R12832 VSS.n8409 VSS.n1762 0.04025
R12833 VSS.n8409 VSS.n8408 0.04025
R12834 VSS.n8408 VSS.n8407 0.04025
R12835 VSS.n8407 VSS.n1764 0.04025
R12836 VSS.n8403 VSS.n1764 0.04025
R12837 VSS.n8403 VSS.n8402 0.04025
R12838 VSS.n8402 VSS.n8401 0.04025
R12839 VSS.n8401 VSS.n1766 0.04025
R12840 VSS.n8397 VSS.n1766 0.04025
R12841 VSS.n8397 VSS.n8396 0.04025
R12842 VSS.n8396 VSS.n8395 0.04025
R12843 VSS.n8395 VSS.n1768 0.04025
R12844 VSS.n8391 VSS.n1768 0.04025
R12845 VSS.n8391 VSS.n8390 0.04025
R12846 VSS.n8390 VSS.n8389 0.04025
R12847 VSS.n8389 VSS.n1770 0.04025
R12848 VSS.n8385 VSS.n1770 0.04025
R12849 VSS.n8385 VSS.n8384 0.04025
R12850 VSS.n8384 VSS.n8383 0.04025
R12851 VSS.n8383 VSS.n1772 0.04025
R12852 VSS.n8379 VSS.n1772 0.04025
R12853 VSS.n8379 VSS.n8378 0.04025
R12854 VSS.n8378 VSS.n8377 0.04025
R12855 VSS.n8377 VSS.n1774 0.04025
R12856 VSS.n8373 VSS.n1774 0.04025
R12857 VSS.n8373 VSS.n8372 0.04025
R12858 VSS.n8372 VSS.n8371 0.04025
R12859 VSS.n8371 VSS.n1776 0.04025
R12860 VSS.n8367 VSS.n1776 0.04025
R12861 VSS.n8367 VSS.n8366 0.04025
R12862 VSS.n8366 VSS.n8365 0.04025
R12863 VSS.n8365 VSS.n1778 0.04025
R12864 VSS.n8361 VSS.n1778 0.04025
R12865 VSS.n8361 VSS.n8360 0.04025
R12866 VSS.n8360 VSS.n8359 0.04025
R12867 VSS.n8359 VSS.n1780 0.04025
R12868 VSS.n8355 VSS.n1780 0.04025
R12869 VSS.n8355 VSS.n8354 0.04025
R12870 VSS.n8354 VSS.n8353 0.04025
R12871 VSS.n8353 VSS.n1782 0.04025
R12872 VSS.n8349 VSS.n1782 0.04025
R12873 VSS.n8349 VSS.n8348 0.04025
R12874 VSS.n8348 VSS.n8347 0.04025
R12875 VSS.n8347 VSS.n1784 0.04025
R12876 VSS.n8343 VSS.n1784 0.04025
R12877 VSS.n8343 VSS.n8342 0.04025
R12878 VSS.n8342 VSS.n8341 0.04025
R12879 VSS.n8341 VSS.n1786 0.04025
R12880 VSS.n8337 VSS.n1786 0.04025
R12881 VSS.n8337 VSS.n8336 0.04025
R12882 VSS.n8336 VSS.n8335 0.04025
R12883 VSS.n8335 VSS.n1788 0.04025
R12884 VSS.n8331 VSS.n1788 0.04025
R12885 VSS.n8331 VSS.n8330 0.04025
R12886 VSS.n8330 VSS.n8329 0.04025
R12887 VSS.n8329 VSS.n1790 0.04025
R12888 VSS.n8325 VSS.n1790 0.04025
R12889 VSS.n8325 VSS.n8324 0.04025
R12890 VSS.n8324 VSS.n8323 0.04025
R12891 VSS.n8323 VSS.n1792 0.04025
R12892 VSS.n8319 VSS.n1792 0.04025
R12893 VSS.n8319 VSS.n8318 0.04025
R12894 VSS.n8318 VSS.n8317 0.04025
R12895 VSS.n8317 VSS.n1794 0.04025
R12896 VSS.n8313 VSS.n1794 0.04025
R12897 VSS.n8313 VSS.n8312 0.04025
R12898 VSS.n8312 VSS.n8311 0.04025
R12899 VSS.n8311 VSS.n1796 0.04025
R12900 VSS.n8307 VSS.n1796 0.04025
R12901 VSS.n8307 VSS.n8306 0.04025
R12902 VSS.n8306 VSS.n8305 0.04025
R12903 VSS.n8305 VSS.n1798 0.04025
R12904 VSS.n8301 VSS.n1798 0.04025
R12905 VSS.n8301 VSS.n8300 0.04025
R12906 VSS.n8300 VSS.n8299 0.04025
R12907 VSS.n8299 VSS.n1800 0.04025
R12908 VSS.n8295 VSS.n1800 0.04025
R12909 VSS.n8295 VSS.n8294 0.04025
R12910 VSS.n8294 VSS.n8293 0.04025
R12911 VSS.n8293 VSS.n1802 0.04025
R12912 VSS.n8289 VSS.n1802 0.04025
R12913 VSS.n8289 VSS.n8288 0.04025
R12914 VSS.n8288 VSS.n8287 0.04025
R12915 VSS.n8287 VSS.n1804 0.04025
R12916 VSS.n8283 VSS.n1804 0.04025
R12917 VSS.n8283 VSS.n8282 0.04025
R12918 VSS.n8282 VSS.n8281 0.04025
R12919 VSS.n8281 VSS.n1806 0.04025
R12920 VSS.n8277 VSS.n1806 0.04025
R12921 VSS.n8277 VSS.n8276 0.04025
R12922 VSS.n8276 VSS.n8275 0.04025
R12923 VSS.n8275 VSS.n1808 0.04025
R12924 VSS.n8271 VSS.n1808 0.04025
R12925 VSS.n8271 VSS.n8270 0.04025
R12926 VSS.n8270 VSS.n8269 0.04025
R12927 VSS.n8269 VSS.n1810 0.04025
R12928 VSS.n8265 VSS.n1810 0.04025
R12929 VSS.n8265 VSS.n8264 0.04025
R12930 VSS.n8264 VSS.n8263 0.04025
R12931 VSS.n8263 VSS.n1812 0.04025
R12932 VSS.n8259 VSS.n1812 0.04025
R12933 VSS.n8259 VSS.n8258 0.04025
R12934 VSS.n8258 VSS.n8257 0.04025
R12935 VSS.n8257 VSS.n1814 0.04025
R12936 VSS.n8253 VSS.n1814 0.04025
R12937 VSS.n8253 VSS.n8252 0.04025
R12938 VSS.n8252 VSS.n8251 0.04025
R12939 VSS.n8251 VSS.n1816 0.04025
R12940 VSS.n8247 VSS.n1816 0.04025
R12941 VSS.n8247 VSS.n8246 0.04025
R12942 VSS.n8246 VSS.n8245 0.04025
R12943 VSS.n8245 VSS.n1818 0.04025
R12944 VSS.n8241 VSS.n1818 0.04025
R12945 VSS.n8241 VSS.n8240 0.04025
R12946 VSS.n8240 VSS.n8239 0.04025
R12947 VSS.n8239 VSS.n1820 0.04025
R12948 VSS.n8235 VSS.n1820 0.04025
R12949 VSS.n8235 VSS.n8234 0.04025
R12950 VSS.n8234 VSS.n8233 0.04025
R12951 VSS.n4144 VSS.n3184 0.04025
R12952 VSS.n4145 VSS.n4144 0.04025
R12953 VSS.n4146 VSS.n4145 0.04025
R12954 VSS.n4146 VSS.n3182 0.04025
R12955 VSS.n4150 VSS.n3182 0.04025
R12956 VSS.n4151 VSS.n4150 0.04025
R12957 VSS.n4152 VSS.n4151 0.04025
R12958 VSS.n4152 VSS.n3180 0.04025
R12959 VSS.n4156 VSS.n3180 0.04025
R12960 VSS.n4157 VSS.n4156 0.04025
R12961 VSS.n4158 VSS.n4157 0.04025
R12962 VSS.n4158 VSS.n3178 0.04025
R12963 VSS.n4162 VSS.n3178 0.04025
R12964 VSS.n4163 VSS.n4162 0.04025
R12965 VSS.n4164 VSS.n4163 0.04025
R12966 VSS.n4164 VSS.n3176 0.04025
R12967 VSS.n4168 VSS.n3176 0.04025
R12968 VSS.n4169 VSS.n4168 0.04025
R12969 VSS.n4170 VSS.n4169 0.04025
R12970 VSS.n4170 VSS.n3174 0.04025
R12971 VSS.n4174 VSS.n3174 0.04025
R12972 VSS.n4175 VSS.n4174 0.04025
R12973 VSS.n4176 VSS.n4175 0.04025
R12974 VSS.n4176 VSS.n3172 0.04025
R12975 VSS.n4180 VSS.n3172 0.04025
R12976 VSS.n4181 VSS.n4180 0.04025
R12977 VSS.n4182 VSS.n4181 0.04025
R12978 VSS.n4182 VSS.n3170 0.04025
R12979 VSS.n4186 VSS.n3170 0.04025
R12980 VSS.n4187 VSS.n4186 0.04025
R12981 VSS.n4188 VSS.n4187 0.04025
R12982 VSS.n4188 VSS.n3168 0.04025
R12983 VSS.n4192 VSS.n3168 0.04025
R12984 VSS.n4193 VSS.n4192 0.04025
R12985 VSS.n4194 VSS.n4193 0.04025
R12986 VSS.n4194 VSS.n3166 0.04025
R12987 VSS.n4198 VSS.n3166 0.04025
R12988 VSS.n4199 VSS.n4198 0.04025
R12989 VSS.n4200 VSS.n4199 0.04025
R12990 VSS.n4200 VSS.n3164 0.04025
R12991 VSS.n4204 VSS.n3164 0.04025
R12992 VSS.n4205 VSS.n4204 0.04025
R12993 VSS.n4206 VSS.n4205 0.04025
R12994 VSS.n4206 VSS.n3162 0.04025
R12995 VSS.n4210 VSS.n3162 0.04025
R12996 VSS.n4211 VSS.n4210 0.04025
R12997 VSS.n4212 VSS.n4211 0.04025
R12998 VSS.n4212 VSS.n3160 0.04025
R12999 VSS.n4216 VSS.n3160 0.04025
R13000 VSS.n4217 VSS.n4216 0.04025
R13001 VSS.n4218 VSS.n4217 0.04025
R13002 VSS.n4218 VSS.n3158 0.04025
R13003 VSS.n4222 VSS.n3158 0.04025
R13004 VSS.n4223 VSS.n4222 0.04025
R13005 VSS.n4224 VSS.n4223 0.04025
R13006 VSS.n4224 VSS.n3156 0.04025
R13007 VSS.n4228 VSS.n3156 0.04025
R13008 VSS.n4229 VSS.n4228 0.04025
R13009 VSS.n4230 VSS.n4229 0.04025
R13010 VSS.n4230 VSS.n3154 0.04025
R13011 VSS.n4234 VSS.n3154 0.04025
R13012 VSS.n4235 VSS.n4234 0.04025
R13013 VSS.n4236 VSS.n4235 0.04025
R13014 VSS.n4236 VSS.n3152 0.04025
R13015 VSS.n4240 VSS.n3152 0.04025
R13016 VSS.n4241 VSS.n4240 0.04025
R13017 VSS.n4242 VSS.n4241 0.04025
R13018 VSS.n4242 VSS.n3150 0.04025
R13019 VSS.n4246 VSS.n3150 0.04025
R13020 VSS.n4247 VSS.n4246 0.04025
R13021 VSS.n4248 VSS.n4247 0.04025
R13022 VSS.n4248 VSS.n3148 0.04025
R13023 VSS.n4252 VSS.n3148 0.04025
R13024 VSS.n4253 VSS.n4252 0.04025
R13025 VSS.n4254 VSS.n4253 0.04025
R13026 VSS.n4254 VSS.n3146 0.04025
R13027 VSS.n4258 VSS.n3146 0.04025
R13028 VSS.n4259 VSS.n4258 0.04025
R13029 VSS.n4260 VSS.n4259 0.04025
R13030 VSS.n4260 VSS.n3144 0.04025
R13031 VSS.n4264 VSS.n3144 0.04025
R13032 VSS.n4265 VSS.n4264 0.04025
R13033 VSS.n4266 VSS.n4265 0.04025
R13034 VSS.n4266 VSS.n3142 0.04025
R13035 VSS.n4270 VSS.n3142 0.04025
R13036 VSS.n4271 VSS.n4270 0.04025
R13037 VSS.n4272 VSS.n4271 0.04025
R13038 VSS.n4272 VSS.n3140 0.04025
R13039 VSS.n4276 VSS.n3140 0.04025
R13040 VSS.n4277 VSS.n4276 0.04025
R13041 VSS.n4278 VSS.n4277 0.04025
R13042 VSS.n4278 VSS.n3138 0.04025
R13043 VSS.n4282 VSS.n3138 0.04025
R13044 VSS.n4283 VSS.n4282 0.04025
R13045 VSS.n4284 VSS.n4283 0.04025
R13046 VSS.n4284 VSS.n3136 0.04025
R13047 VSS.n4288 VSS.n3136 0.04025
R13048 VSS.n4289 VSS.n4288 0.04025
R13049 VSS.n4290 VSS.n4289 0.04025
R13050 VSS.n4290 VSS.n3134 0.04025
R13051 VSS.n4294 VSS.n3134 0.04025
R13052 VSS.n4295 VSS.n4294 0.04025
R13053 VSS.n4296 VSS.n4295 0.04025
R13054 VSS.n4296 VSS.n3132 0.04025
R13055 VSS.n4300 VSS.n3132 0.04025
R13056 VSS.n4301 VSS.n4300 0.04025
R13057 VSS.n4302 VSS.n4301 0.04025
R13058 VSS.n4302 VSS.n3130 0.04025
R13059 VSS.n4306 VSS.n3130 0.04025
R13060 VSS.n4307 VSS.n4306 0.04025
R13061 VSS.n4308 VSS.n4307 0.04025
R13062 VSS.n4308 VSS.n3128 0.04025
R13063 VSS.n4312 VSS.n3128 0.04025
R13064 VSS.n4313 VSS.n4312 0.04025
R13065 VSS.n4314 VSS.n4313 0.04025
R13066 VSS.n4314 VSS.n3126 0.04025
R13067 VSS.n4318 VSS.n3126 0.04025
R13068 VSS.n4319 VSS.n4318 0.04025
R13069 VSS.n4320 VSS.n4319 0.04025
R13070 VSS.n4320 VSS.n3124 0.04025
R13071 VSS.n4324 VSS.n3124 0.04025
R13072 VSS.n4325 VSS.n4324 0.04025
R13073 VSS.n4326 VSS.n4325 0.04025
R13074 VSS.n4326 VSS.n3122 0.04025
R13075 VSS.n4330 VSS.n3122 0.04025
R13076 VSS.n4331 VSS.n4330 0.04025
R13077 VSS.n4332 VSS.n4331 0.04025
R13078 VSS.n4332 VSS.n3120 0.04025
R13079 VSS.n4336 VSS.n3120 0.04025
R13080 VSS.n4337 VSS.n4336 0.04025
R13081 VSS.n4338 VSS.n4337 0.04025
R13082 VSS.n4338 VSS.n3118 0.04025
R13083 VSS.n4342 VSS.n3118 0.04025
R13084 VSS.n4343 VSS.n4342 0.04025
R13085 VSS.n4344 VSS.n4343 0.04025
R13086 VSS.n4344 VSS.n3116 0.04025
R13087 VSS.n4348 VSS.n3116 0.04025
R13088 VSS.n4349 VSS.n4348 0.04025
R13089 VSS.n4350 VSS.n4349 0.04025
R13090 VSS.n4350 VSS.n3114 0.04025
R13091 VSS.n4354 VSS.n3114 0.04025
R13092 VSS.n4355 VSS.n4354 0.04025
R13093 VSS.n4356 VSS.n4355 0.04025
R13094 VSS.n4356 VSS.n3112 0.04025
R13095 VSS.n4360 VSS.n3112 0.04025
R13096 VSS.n4361 VSS.n4360 0.04025
R13097 VSS.n4362 VSS.n4361 0.04025
R13098 VSS.n4362 VSS.n3110 0.04025
R13099 VSS.n4366 VSS.n3110 0.04025
R13100 VSS.n4367 VSS.n4366 0.04025
R13101 VSS.n4368 VSS.n4367 0.04025
R13102 VSS.n4368 VSS.n3108 0.04025
R13103 VSS.n4372 VSS.n3108 0.04025
R13104 VSS.n4373 VSS.n4372 0.04025
R13105 VSS.n4374 VSS.n4373 0.04025
R13106 VSS.n4374 VSS.n3106 0.04025
R13107 VSS.n4378 VSS.n3106 0.04025
R13108 VSS.n4379 VSS.n4378 0.04025
R13109 VSS.n4380 VSS.n4379 0.04025
R13110 VSS.n4380 VSS.n3104 0.04025
R13111 VSS.n4384 VSS.n3104 0.04025
R13112 VSS.n4385 VSS.n4384 0.04025
R13113 VSS.n4386 VSS.n4385 0.04025
R13114 VSS.n4386 VSS.n3102 0.04025
R13115 VSS.n4390 VSS.n3102 0.04025
R13116 VSS.n4391 VSS.n4390 0.04025
R13117 VSS.n4392 VSS.n4391 0.04025
R13118 VSS.n4392 VSS.n3100 0.04025
R13119 VSS.n4396 VSS.n3100 0.04025
R13120 VSS.n4397 VSS.n4396 0.04025
R13121 VSS.n4398 VSS.n4397 0.04025
R13122 VSS.n4398 VSS.n3098 0.04025
R13123 VSS.n4402 VSS.n3098 0.04025
R13124 VSS.n4403 VSS.n4402 0.04025
R13125 VSS.n4404 VSS.n4403 0.04025
R13126 VSS.n4404 VSS.n3096 0.04025
R13127 VSS.n4408 VSS.n3096 0.04025
R13128 VSS.n4409 VSS.n4408 0.04025
R13129 VSS.n4410 VSS.n4409 0.04025
R13130 VSS.n4410 VSS.n3094 0.04025
R13131 VSS.n4414 VSS.n3094 0.04025
R13132 VSS.n4415 VSS.n4414 0.04025
R13133 VSS.n4416 VSS.n4415 0.04025
R13134 VSS.n4416 VSS.n3092 0.04025
R13135 VSS.n4420 VSS.n3092 0.04025
R13136 VSS.n4421 VSS.n4420 0.04025
R13137 VSS.n4422 VSS.n4421 0.04025
R13138 VSS.n4422 VSS.n3090 0.04025
R13139 VSS.n4426 VSS.n3090 0.04025
R13140 VSS.n4427 VSS.n4426 0.04025
R13141 VSS.n4428 VSS.n4427 0.04025
R13142 VSS.n4428 VSS.n3088 0.04025
R13143 VSS.n4432 VSS.n3088 0.04025
R13144 VSS.n4433 VSS.n4432 0.04025
R13145 VSS.n4434 VSS.n4433 0.04025
R13146 VSS.n4434 VSS.n3086 0.04025
R13147 VSS.n4438 VSS.n3086 0.04025
R13148 VSS.n4439 VSS.n4438 0.04025
R13149 VSS.n4440 VSS.n4439 0.04025
R13150 VSS.n4440 VSS.n3084 0.04025
R13151 VSS.n4444 VSS.n3084 0.04025
R13152 VSS.n4445 VSS.n4444 0.04025
R13153 VSS.n4446 VSS.n4445 0.04025
R13154 VSS.n4446 VSS.n3082 0.04025
R13155 VSS.n4450 VSS.n3082 0.04025
R13156 VSS.n4451 VSS.n4450 0.04025
R13157 VSS.n4452 VSS.n4451 0.04025
R13158 VSS.n4452 VSS.n3080 0.04025
R13159 VSS.n4456 VSS.n3080 0.04025
R13160 VSS.n4457 VSS.n4456 0.04025
R13161 VSS.n4458 VSS.n4457 0.04025
R13162 VSS.n4458 VSS.n3078 0.04025
R13163 VSS.n4462 VSS.n3078 0.04025
R13164 VSS.n4463 VSS.n4462 0.04025
R13165 VSS.n4464 VSS.n4463 0.04025
R13166 VSS.n4464 VSS.n3076 0.04025
R13167 VSS.n4468 VSS.n3076 0.04025
R13168 VSS.n4469 VSS.n4468 0.04025
R13169 VSS.n4470 VSS.n4469 0.04025
R13170 VSS.n4470 VSS.n3074 0.04025
R13171 VSS.n4474 VSS.n3074 0.04025
R13172 VSS.n4475 VSS.n4474 0.04025
R13173 VSS.n4476 VSS.n4475 0.04025
R13174 VSS.n4476 VSS.n3072 0.04025
R13175 VSS.n4480 VSS.n3072 0.04025
R13176 VSS.n4481 VSS.n4480 0.04025
R13177 VSS.n4482 VSS.n4481 0.04025
R13178 VSS.n4482 VSS.n3070 0.04025
R13179 VSS.n4486 VSS.n3070 0.04025
R13180 VSS.n4487 VSS.n4486 0.04025
R13181 VSS.n4488 VSS.n4487 0.04025
R13182 VSS.n4488 VSS.n3068 0.04025
R13183 VSS.n4492 VSS.n3068 0.04025
R13184 VSS.n4493 VSS.n4492 0.04025
R13185 VSS.n4494 VSS.n4493 0.04025
R13186 VSS.n4494 VSS.n3066 0.04025
R13187 VSS.n4498 VSS.n3066 0.04025
R13188 VSS.n4499 VSS.n4498 0.04025
R13189 VSS.n4500 VSS.n4499 0.04025
R13190 VSS.n4500 VSS.n3064 0.04025
R13191 VSS.n4504 VSS.n3064 0.04025
R13192 VSS.n4505 VSS.n4504 0.04025
R13193 VSS.n4506 VSS.n4505 0.04025
R13194 VSS.n4506 VSS.n3062 0.04025
R13195 VSS.n4510 VSS.n3062 0.04025
R13196 VSS.n4511 VSS.n4510 0.04025
R13197 VSS.n4512 VSS.n4511 0.04025
R13198 VSS.n4512 VSS.n3060 0.04025
R13199 VSS.n4516 VSS.n3060 0.04025
R13200 VSS.n4517 VSS.n4516 0.04025
R13201 VSS.n4518 VSS.n4517 0.04025
R13202 VSS.n4518 VSS.n3058 0.04025
R13203 VSS.n4522 VSS.n3058 0.04025
R13204 VSS.n4523 VSS.n4522 0.04025
R13205 VSS.n4524 VSS.n4523 0.04025
R13206 VSS.n4524 VSS.n3056 0.04025
R13207 VSS.n4528 VSS.n3056 0.04025
R13208 VSS.n4529 VSS.n4528 0.04025
R13209 VSS.n4530 VSS.n4529 0.04025
R13210 VSS.n4530 VSS.n3054 0.04025
R13211 VSS.n4534 VSS.n3054 0.04025
R13212 VSS.n4535 VSS.n4534 0.04025
R13213 VSS.n4536 VSS.n4535 0.04025
R13214 VSS.n4536 VSS.n3052 0.04025
R13215 VSS.n4540 VSS.n3052 0.04025
R13216 VSS.n4541 VSS.n4540 0.04025
R13217 VSS.n4542 VSS.n4541 0.04025
R13218 VSS.n4542 VSS.n3050 0.04025
R13219 VSS.n4546 VSS.n3050 0.04025
R13220 VSS.n4547 VSS.n4546 0.04025
R13221 VSS.n4548 VSS.n4547 0.04025
R13222 VSS.n4548 VSS.n3048 0.04025
R13223 VSS.n4552 VSS.n3048 0.04025
R13224 VSS.n4553 VSS.n4552 0.04025
R13225 VSS.n4554 VSS.n4553 0.04025
R13226 VSS.n4554 VSS.n3046 0.04025
R13227 VSS.n4558 VSS.n3046 0.04025
R13228 VSS.n4559 VSS.n4558 0.04025
R13229 VSS.n4560 VSS.n4559 0.04025
R13230 VSS.n4560 VSS.n3044 0.04025
R13231 VSS.n4564 VSS.n3044 0.04025
R13232 VSS.n4565 VSS.n4564 0.04025
R13233 VSS.n4566 VSS.n4565 0.04025
R13234 VSS.n4566 VSS.n3042 0.04025
R13235 VSS.n4570 VSS.n3042 0.04025
R13236 VSS.n4571 VSS.n4570 0.04025
R13237 VSS.n4572 VSS.n4571 0.04025
R13238 VSS.n4572 VSS.n3040 0.04025
R13239 VSS.n4576 VSS.n3040 0.04025
R13240 VSS.n4577 VSS.n4576 0.04025
R13241 VSS.n4578 VSS.n4577 0.04025
R13242 VSS.n4578 VSS.n3038 0.04025
R13243 VSS.n4582 VSS.n3038 0.04025
R13244 VSS.n4583 VSS.n4582 0.04025
R13245 VSS.n4584 VSS.n4583 0.04025
R13246 VSS.n4584 VSS.n3036 0.04025
R13247 VSS.n4588 VSS.n3036 0.04025
R13248 VSS.n4589 VSS.n4588 0.04025
R13249 VSS.n4590 VSS.n4589 0.04025
R13250 VSS.n4590 VSS.n3034 0.04025
R13251 VSS.n4594 VSS.n3034 0.04025
R13252 VSS.n4595 VSS.n4594 0.04025
R13253 VSS.n4596 VSS.n4595 0.04025
R13254 VSS.n4596 VSS.n3032 0.04025
R13255 VSS.n4600 VSS.n3032 0.04025
R13256 VSS.n4601 VSS.n4600 0.04025
R13257 VSS.n4602 VSS.n4601 0.04025
R13258 VSS.n4602 VSS.n3030 0.04025
R13259 VSS.n4606 VSS.n3030 0.04025
R13260 VSS.n4607 VSS.n4606 0.04025
R13261 VSS.n4608 VSS.n4607 0.04025
R13262 VSS.n4608 VSS.n3028 0.04025
R13263 VSS.n4612 VSS.n3028 0.04025
R13264 VSS.n4613 VSS.n4612 0.04025
R13265 VSS.n4614 VSS.n4613 0.04025
R13266 VSS.n4614 VSS.n3026 0.04025
R13267 VSS.n4618 VSS.n3026 0.04025
R13268 VSS.n4619 VSS.n4618 0.04025
R13269 VSS.n4620 VSS.n4619 0.04025
R13270 VSS.n4620 VSS.n3024 0.04025
R13271 VSS.n4624 VSS.n3024 0.04025
R13272 VSS.n4625 VSS.n4624 0.04025
R13273 VSS.n4626 VSS.n4625 0.04025
R13274 VSS.n4626 VSS.n3022 0.04025
R13275 VSS.n4630 VSS.n3022 0.04025
R13276 VSS.n4631 VSS.n4630 0.04025
R13277 VSS.n4632 VSS.n4631 0.04025
R13278 VSS.n4632 VSS.n3020 0.04025
R13279 VSS.n4636 VSS.n3020 0.04025
R13280 VSS.n4637 VSS.n4636 0.04025
R13281 VSS.n4638 VSS.n4637 0.04025
R13282 VSS.n4638 VSS.n3018 0.04025
R13283 VSS.n4642 VSS.n3018 0.04025
R13284 VSS.n4643 VSS.n4642 0.04025
R13285 VSS.n4644 VSS.n4643 0.04025
R13286 VSS.n4644 VSS.n3016 0.04025
R13287 VSS.n4648 VSS.n3016 0.04025
R13288 VSS.n4649 VSS.n4648 0.04025
R13289 VSS.n4650 VSS.n4649 0.04025
R13290 VSS.n4650 VSS.n3014 0.04025
R13291 VSS.n4654 VSS.n3014 0.04025
R13292 VSS.n4655 VSS.n4654 0.04025
R13293 VSS.n4656 VSS.n4655 0.04025
R13294 VSS.n4656 VSS.n3012 0.04025
R13295 VSS.n4660 VSS.n3012 0.04025
R13296 VSS.n4661 VSS.n4660 0.04025
R13297 VSS.n4662 VSS.n4661 0.04025
R13298 VSS.n4662 VSS.n3010 0.04025
R13299 VSS.n4666 VSS.n3010 0.04025
R13300 VSS.n4667 VSS.n4666 0.04025
R13301 VSS.n4668 VSS.n4667 0.04025
R13302 VSS.n4668 VSS.n3008 0.04025
R13303 VSS.n4672 VSS.n3008 0.04025
R13304 VSS.n4673 VSS.n4672 0.04025
R13305 VSS.n4674 VSS.n4673 0.04025
R13306 VSS.n4674 VSS.n3006 0.04025
R13307 VSS.n4678 VSS.n3006 0.04025
R13308 VSS.n4679 VSS.n4678 0.04025
R13309 VSS.n4680 VSS.n4679 0.04025
R13310 VSS.n4680 VSS.n3004 0.04025
R13311 VSS.n4684 VSS.n3004 0.04025
R13312 VSS.n4685 VSS.n4684 0.04025
R13313 VSS.n4686 VSS.n4685 0.04025
R13314 VSS.n4686 VSS.n3002 0.04025
R13315 VSS.n4690 VSS.n3002 0.04025
R13316 VSS.n4691 VSS.n4690 0.04025
R13317 VSS.n4692 VSS.n4691 0.04025
R13318 VSS.n4692 VSS.n3000 0.04025
R13319 VSS.n4696 VSS.n3000 0.04025
R13320 VSS.n4697 VSS.n4696 0.04025
R13321 VSS.n4698 VSS.n4697 0.04025
R13322 VSS.n4698 VSS.n2998 0.04025
R13323 VSS.n4702 VSS.n2998 0.04025
R13324 VSS.n4703 VSS.n4702 0.04025
R13325 VSS.n4704 VSS.n4703 0.04025
R13326 VSS.n4704 VSS.n2996 0.04025
R13327 VSS.n4708 VSS.n2996 0.04025
R13328 VSS.n4709 VSS.n4708 0.04025
R13329 VSS.n4710 VSS.n4709 0.04025
R13330 VSS.n4710 VSS.n2994 0.04025
R13331 VSS.n4714 VSS.n2994 0.04025
R13332 VSS.n4715 VSS.n4714 0.04025
R13333 VSS.n4716 VSS.n4715 0.04025
R13334 VSS.n4716 VSS.n2992 0.04025
R13335 VSS.n4720 VSS.n2992 0.04025
R13336 VSS.n4721 VSS.n4720 0.04025
R13337 VSS.n4722 VSS.n4721 0.04025
R13338 VSS.n4722 VSS.n2990 0.04025
R13339 VSS.n4726 VSS.n2990 0.04025
R13340 VSS.n4727 VSS.n4726 0.04025
R13341 VSS.n4728 VSS.n4727 0.04025
R13342 VSS.n4728 VSS.n2988 0.04025
R13343 VSS.n4732 VSS.n2988 0.04025
R13344 VSS.n4733 VSS.n4732 0.04025
R13345 VSS.n4734 VSS.n4733 0.04025
R13346 VSS.n4734 VSS.n2986 0.04025
R13347 VSS.n4738 VSS.n2986 0.04025
R13348 VSS.n4739 VSS.n4738 0.04025
R13349 VSS.n4740 VSS.n4739 0.04025
R13350 VSS.n4740 VSS.n2984 0.04025
R13351 VSS.n4744 VSS.n2984 0.04025
R13352 VSS.n4745 VSS.n4744 0.04025
R13353 VSS.n4746 VSS.n4745 0.04025
R13354 VSS.n4746 VSS.n2982 0.04025
R13355 VSS.n4750 VSS.n2982 0.04025
R13356 VSS.n4751 VSS.n4750 0.04025
R13357 VSS.n4752 VSS.n4751 0.04025
R13358 VSS.n4752 VSS.n2980 0.04025
R13359 VSS.n4756 VSS.n2980 0.04025
R13360 VSS.n4757 VSS.n4756 0.04025
R13361 VSS.n4758 VSS.n4757 0.04025
R13362 VSS.n4758 VSS.n2978 0.04025
R13363 VSS.n4762 VSS.n2978 0.04025
R13364 VSS.n4763 VSS.n4762 0.04025
R13365 VSS.n4764 VSS.n4763 0.04025
R13366 VSS.n4764 VSS.n2976 0.04025
R13367 VSS.n4768 VSS.n2976 0.04025
R13368 VSS.n4769 VSS.n4768 0.04025
R13369 VSS.n4770 VSS.n4769 0.04025
R13370 VSS.n4770 VSS.n2974 0.04025
R13371 VSS.n4774 VSS.n2974 0.04025
R13372 VSS.n4775 VSS.n4774 0.04025
R13373 VSS.n4776 VSS.n4775 0.04025
R13374 VSS.n4776 VSS.n2972 0.04025
R13375 VSS.n4780 VSS.n2972 0.04025
R13376 VSS.n4781 VSS.n4780 0.04025
R13377 VSS.n4782 VSS.n4781 0.04025
R13378 VSS.n4782 VSS.n2970 0.04025
R13379 VSS.n4786 VSS.n2970 0.04025
R13380 VSS.n4787 VSS.n4786 0.04025
R13381 VSS.n4788 VSS.n4787 0.04025
R13382 VSS.n4788 VSS.n2968 0.04025
R13383 VSS.n4792 VSS.n2968 0.04025
R13384 VSS.n4793 VSS.n4792 0.04025
R13385 VSS.n4794 VSS.n4793 0.04025
R13386 VSS.n4794 VSS.n2966 0.04025
R13387 VSS.n4798 VSS.n2966 0.04025
R13388 VSS.n4799 VSS.n4798 0.04025
R13389 VSS.n4800 VSS.n4799 0.04025
R13390 VSS.n4800 VSS.n2964 0.04025
R13391 VSS.n4807 VSS.n2964 0.04025
R13392 VSS.n4808 VSS.n4807 0.04025
R13393 VSS.n4809 VSS.n4808 0.04025
R13394 VSS.n4809 VSS.n2962 0.04025
R13395 VSS.n4813 VSS.n2962 0.04025
R13396 VSS.n4814 VSS.n4813 0.04025
R13397 VSS.n4815 VSS.n4814 0.04025
R13398 VSS.n4815 VSS.n2960 0.04025
R13399 VSS.n4819 VSS.n2960 0.04025
R13400 VSS.n4820 VSS.n4819 0.04025
R13401 VSS.n4821 VSS.n4820 0.04025
R13402 VSS.n4821 VSS.n2958 0.04025
R13403 VSS.n4825 VSS.n2958 0.04025
R13404 VSS.n4826 VSS.n4825 0.04025
R13405 VSS.n4827 VSS.n4826 0.04025
R13406 VSS.n4827 VSS.n2956 0.04025
R13407 VSS.n4831 VSS.n2956 0.04025
R13408 VSS.n4832 VSS.n4831 0.04025
R13409 VSS.n4833 VSS.n4832 0.04025
R13410 VSS.n4833 VSS.n2954 0.04025
R13411 VSS.n4837 VSS.n2954 0.04025
R13412 VSS.n4838 VSS.n4837 0.04025
R13413 VSS.n4839 VSS.n4838 0.04025
R13414 VSS.n4839 VSS.n2952 0.04025
R13415 VSS.n4843 VSS.n2952 0.04025
R13416 VSS.n4844 VSS.n4843 0.04025
R13417 VSS.n4845 VSS.n4844 0.04025
R13418 VSS.n4845 VSS.n2950 0.04025
R13419 VSS.n4849 VSS.n2950 0.04025
R13420 VSS.n4850 VSS.n4849 0.04025
R13421 VSS.n4851 VSS.n4850 0.04025
R13422 VSS.n4851 VSS.n2948 0.04025
R13423 VSS.n4855 VSS.n2948 0.04025
R13424 VSS.n4856 VSS.n4855 0.04025
R13425 VSS.n4857 VSS.n4856 0.04025
R13426 VSS.n4857 VSS.n2946 0.04025
R13427 VSS.n4861 VSS.n2946 0.04025
R13428 VSS.n4862 VSS.n4861 0.04025
R13429 VSS.n4863 VSS.n4862 0.04025
R13430 VSS.n4863 VSS.n2944 0.04025
R13431 VSS.n4867 VSS.n2944 0.04025
R13432 VSS.n4868 VSS.n4867 0.04025
R13433 VSS.n4869 VSS.n4868 0.04025
R13434 VSS.n4869 VSS.n2942 0.04025
R13435 VSS.n4873 VSS.n2942 0.04025
R13436 VSS.n4874 VSS.n4873 0.04025
R13437 VSS.n4875 VSS.n4874 0.04025
R13438 VSS.n4875 VSS.n2940 0.04025
R13439 VSS.n4879 VSS.n2940 0.04025
R13440 VSS.n4880 VSS.n4879 0.04025
R13441 VSS.n4881 VSS.n4880 0.04025
R13442 VSS.n4881 VSS.n2938 0.04025
R13443 VSS.n4885 VSS.n2938 0.04025
R13444 VSS.n4886 VSS.n4885 0.04025
R13445 VSS.n4887 VSS.n4886 0.04025
R13446 VSS.n4887 VSS.n2936 0.04025
R13447 VSS.n4891 VSS.n2936 0.04025
R13448 VSS.n4892 VSS.n4891 0.04025
R13449 VSS.n4893 VSS.n4892 0.04025
R13450 VSS.n4893 VSS.n2934 0.04025
R13451 VSS.n4897 VSS.n2934 0.04025
R13452 VSS.n4898 VSS.n4897 0.04025
R13453 VSS.n4899 VSS.n4898 0.04025
R13454 VSS.n4899 VSS.n2932 0.04025
R13455 VSS.n4903 VSS.n2932 0.04025
R13456 VSS.n4904 VSS.n4903 0.04025
R13457 VSS.n4905 VSS.n4904 0.04025
R13458 VSS.n4905 VSS.n2930 0.04025
R13459 VSS.n4909 VSS.n2930 0.04025
R13460 VSS.n4910 VSS.n4909 0.04025
R13461 VSS.n4911 VSS.n4910 0.04025
R13462 VSS.n4911 VSS.n2928 0.04025
R13463 VSS.n4915 VSS.n2928 0.04025
R13464 VSS.n4916 VSS.n4915 0.04025
R13465 VSS.n4917 VSS.n4916 0.04025
R13466 VSS.n4917 VSS.n2926 0.04025
R13467 VSS.n4921 VSS.n2926 0.04025
R13468 VSS.n4922 VSS.n4921 0.04025
R13469 VSS.n4923 VSS.n4922 0.04025
R13470 VSS.n4923 VSS.n2924 0.04025
R13471 VSS.n4927 VSS.n2924 0.04025
R13472 VSS.n4928 VSS.n4927 0.04025
R13473 VSS.n4929 VSS.n4928 0.04025
R13474 VSS.n4929 VSS.n2922 0.04025
R13475 VSS.n4933 VSS.n2922 0.04025
R13476 VSS.n4934 VSS.n4933 0.04025
R13477 VSS.n4935 VSS.n4934 0.04025
R13478 VSS.n4935 VSS.n2920 0.04025
R13479 VSS.n4939 VSS.n2920 0.04025
R13480 VSS.n4940 VSS.n4939 0.04025
R13481 VSS.n4941 VSS.n4940 0.04025
R13482 VSS.n4941 VSS.n2918 0.04025
R13483 VSS.n4945 VSS.n2918 0.04025
R13484 VSS.n4946 VSS.n4945 0.04025
R13485 VSS.n4947 VSS.n4946 0.04025
R13486 VSS.n4947 VSS.n2916 0.04025
R13487 VSS.n4951 VSS.n2916 0.04025
R13488 VSS.n4952 VSS.n4951 0.04025
R13489 VSS.n4953 VSS.n4952 0.04025
R13490 VSS.n4953 VSS.n2914 0.04025
R13491 VSS.n4957 VSS.n2914 0.04025
R13492 VSS.n4958 VSS.n4957 0.04025
R13493 VSS.n4959 VSS.n4958 0.04025
R13494 VSS.n4959 VSS.n2912 0.04025
R13495 VSS.n4963 VSS.n2912 0.04025
R13496 VSS.n4964 VSS.n4963 0.04025
R13497 VSS.n4965 VSS.n4964 0.04025
R13498 VSS.n4965 VSS.n2910 0.04025
R13499 VSS.n4969 VSS.n2910 0.04025
R13500 VSS.n4970 VSS.n4969 0.04025
R13501 VSS.n4971 VSS.n4970 0.04025
R13502 VSS.n4971 VSS.n2908 0.04025
R13503 VSS.n4975 VSS.n2908 0.04025
R13504 VSS.n4976 VSS.n4975 0.04025
R13505 VSS.n4977 VSS.n4976 0.04025
R13506 VSS.n4977 VSS.n2906 0.04025
R13507 VSS.n4981 VSS.n2906 0.04025
R13508 VSS.n4982 VSS.n4981 0.04025
R13509 VSS.n4983 VSS.n4982 0.04025
R13510 VSS.n4983 VSS.n2904 0.04025
R13511 VSS.n4987 VSS.n2904 0.04025
R13512 VSS.n4988 VSS.n4987 0.04025
R13513 VSS.n4989 VSS.n4988 0.04025
R13514 VSS.n4989 VSS.n2902 0.04025
R13515 VSS.n4993 VSS.n2902 0.04025
R13516 VSS.n4994 VSS.n4993 0.04025
R13517 VSS.n4995 VSS.n4994 0.04025
R13518 VSS.n4995 VSS.n2900 0.04025
R13519 VSS.n4999 VSS.n2900 0.04025
R13520 VSS.n5000 VSS.n4999 0.04025
R13521 VSS.n5001 VSS.n5000 0.04025
R13522 VSS.n5001 VSS.n2898 0.04025
R13523 VSS.n5005 VSS.n2898 0.04025
R13524 VSS.n5006 VSS.n5005 0.04025
R13525 VSS.n5007 VSS.n5006 0.04025
R13526 VSS.n5007 VSS.n2896 0.04025
R13527 VSS.n5011 VSS.n2896 0.04025
R13528 VSS.n5012 VSS.n5011 0.04025
R13529 VSS.n5013 VSS.n5012 0.04025
R13530 VSS.n5013 VSS.n2894 0.04025
R13531 VSS.n5017 VSS.n2894 0.04025
R13532 VSS.n5018 VSS.n5017 0.04025
R13533 VSS.n5019 VSS.n5018 0.04025
R13534 VSS.n5019 VSS.n2892 0.04025
R13535 VSS.n5023 VSS.n2892 0.04025
R13536 VSS.n5024 VSS.n5023 0.04025
R13537 VSS.n5025 VSS.n5024 0.04025
R13538 VSS.n5025 VSS.n2890 0.04025
R13539 VSS.n5029 VSS.n2890 0.04025
R13540 VSS.n5030 VSS.n5029 0.04025
R13541 VSS.n5031 VSS.n5030 0.04025
R13542 VSS.n5031 VSS.n2888 0.04025
R13543 VSS.n5035 VSS.n2888 0.04025
R13544 VSS.n5036 VSS.n5035 0.04025
R13545 VSS.n5037 VSS.n5036 0.04025
R13546 VSS.n5037 VSS.n2886 0.04025
R13547 VSS.n5041 VSS.n2886 0.04025
R13548 VSS.n5042 VSS.n5041 0.04025
R13549 VSS.n5043 VSS.n5042 0.04025
R13550 VSS.n5043 VSS.n2884 0.04025
R13551 VSS.n5047 VSS.n2884 0.04025
R13552 VSS.n5048 VSS.n5047 0.04025
R13553 VSS.n5049 VSS.n5048 0.04025
R13554 VSS.n5049 VSS.n2882 0.04025
R13555 VSS.n5053 VSS.n2882 0.04025
R13556 VSS.n5054 VSS.n5053 0.04025
R13557 VSS.n5055 VSS.n5054 0.04025
R13558 VSS.n5055 VSS.n2880 0.04025
R13559 VSS.n5059 VSS.n2880 0.04025
R13560 VSS.n5060 VSS.n5059 0.04025
R13561 VSS.n5061 VSS.n5060 0.04025
R13562 VSS.n5061 VSS.n2878 0.04025
R13563 VSS.n5065 VSS.n2878 0.04025
R13564 VSS.n5066 VSS.n5065 0.04025
R13565 VSS.n5067 VSS.n5066 0.04025
R13566 VSS.n5067 VSS.n2876 0.04025
R13567 VSS.n5071 VSS.n2876 0.04025
R13568 VSS.n5072 VSS.n5071 0.04025
R13569 VSS.n5073 VSS.n5072 0.04025
R13570 VSS.n5073 VSS.n2874 0.04025
R13571 VSS.n5077 VSS.n2874 0.04025
R13572 VSS.n5078 VSS.n5077 0.04025
R13573 VSS.n5079 VSS.n5078 0.04025
R13574 VSS.n5079 VSS.n2872 0.04025
R13575 VSS.n5083 VSS.n2872 0.04025
R13576 VSS.n5084 VSS.n5083 0.04025
R13577 VSS.n5085 VSS.n5084 0.04025
R13578 VSS.n5085 VSS.n2870 0.04025
R13579 VSS.n5089 VSS.n2870 0.04025
R13580 VSS.n5090 VSS.n5089 0.04025
R13581 VSS.n5091 VSS.n5090 0.04025
R13582 VSS.n5091 VSS.n2868 0.04025
R13583 VSS.n5095 VSS.n2868 0.04025
R13584 VSS.n5096 VSS.n5095 0.04025
R13585 VSS.n5097 VSS.n5096 0.04025
R13586 VSS.n5097 VSS.n2866 0.04025
R13587 VSS.n5101 VSS.n2866 0.04025
R13588 VSS.n5102 VSS.n5101 0.04025
R13589 VSS.n5103 VSS.n5102 0.04025
R13590 VSS.n5103 VSS.n2864 0.04025
R13591 VSS.n5107 VSS.n2864 0.04025
R13592 VSS.n5108 VSS.n5107 0.04025
R13593 VSS.n5109 VSS.n5108 0.04025
R13594 VSS.n5109 VSS.n2862 0.04025
R13595 VSS.n5113 VSS.n2862 0.04025
R13596 VSS.n5114 VSS.n5113 0.04025
R13597 VSS.n5115 VSS.n5114 0.04025
R13598 VSS.n5115 VSS.n2860 0.04025
R13599 VSS.n5119 VSS.n2860 0.04025
R13600 VSS.n5120 VSS.n5119 0.04025
R13601 VSS.n5121 VSS.n5120 0.04025
R13602 VSS.n5121 VSS.n2858 0.04025
R13603 VSS.n5125 VSS.n2858 0.04025
R13604 VSS.n5126 VSS.n5125 0.04025
R13605 VSS.n5127 VSS.n5126 0.04025
R13606 VSS.n5127 VSS.n2856 0.04025
R13607 VSS.n5131 VSS.n2856 0.04025
R13608 VSS.n5132 VSS.n5131 0.04025
R13609 VSS.n5133 VSS.n5132 0.04025
R13610 VSS.n5133 VSS.n2854 0.04025
R13611 VSS.n5137 VSS.n2854 0.04025
R13612 VSS.n5138 VSS.n5137 0.04025
R13613 VSS.n5139 VSS.n5138 0.04025
R13614 VSS.n5139 VSS.n2852 0.04025
R13615 VSS.n5143 VSS.n2852 0.04025
R13616 VSS.n5144 VSS.n5143 0.04025
R13617 VSS.n5145 VSS.n5144 0.04025
R13618 VSS.n5145 VSS.n2850 0.04025
R13619 VSS.n5149 VSS.n2850 0.04025
R13620 VSS.n5150 VSS.n5149 0.04025
R13621 VSS.n5151 VSS.n5150 0.04025
R13622 VSS.n5151 VSS.n2848 0.04025
R13623 VSS.n5155 VSS.n2848 0.04025
R13624 VSS.n5156 VSS.n5155 0.04025
R13625 VSS.n5157 VSS.n5156 0.04025
R13626 VSS.n5157 VSS.n2846 0.04025
R13627 VSS.n5161 VSS.n2846 0.04025
R13628 VSS.n5162 VSS.n5161 0.04025
R13629 VSS.n5163 VSS.n5162 0.04025
R13630 VSS.n5163 VSS.n2844 0.04025
R13631 VSS.n5167 VSS.n2844 0.04025
R13632 VSS.n5168 VSS.n5167 0.04025
R13633 VSS.n5169 VSS.n5168 0.04025
R13634 VSS.n5169 VSS.n2842 0.04025
R13635 VSS.n5173 VSS.n2842 0.04025
R13636 VSS.n5174 VSS.n5173 0.04025
R13637 VSS.n5175 VSS.n5174 0.04025
R13638 VSS.n5175 VSS.n2840 0.04025
R13639 VSS.n5179 VSS.n2840 0.04025
R13640 VSS.n5180 VSS.n5179 0.04025
R13641 VSS.n5181 VSS.n5180 0.04025
R13642 VSS.n5181 VSS.n2838 0.04025
R13643 VSS.n5185 VSS.n2838 0.04025
R13644 VSS.n5186 VSS.n5185 0.04025
R13645 VSS.n5187 VSS.n5186 0.04025
R13646 VSS.n5187 VSS.n2836 0.04025
R13647 VSS.n5191 VSS.n2836 0.04025
R13648 VSS.n5192 VSS.n5191 0.04025
R13649 VSS.n5193 VSS.n5192 0.04025
R13650 VSS.n5193 VSS.n2834 0.04025
R13651 VSS.n5197 VSS.n2834 0.04025
R13652 VSS.n5198 VSS.n5197 0.04025
R13653 VSS.n5199 VSS.n5198 0.04025
R13654 VSS.n5199 VSS.n2832 0.04025
R13655 VSS.n5203 VSS.n2832 0.04025
R13656 VSS.n5204 VSS.n5203 0.04025
R13657 VSS.n5205 VSS.n5204 0.04025
R13658 VSS.n5205 VSS.n2830 0.04025
R13659 VSS.n5209 VSS.n2830 0.04025
R13660 VSS.n5210 VSS.n5209 0.04025
R13661 VSS.n5211 VSS.n5210 0.04025
R13662 VSS.n5211 VSS.n2828 0.04025
R13663 VSS.n5215 VSS.n2828 0.04025
R13664 VSS.n5216 VSS.n5215 0.04025
R13665 VSS.n5217 VSS.n5216 0.04025
R13666 VSS.n5217 VSS.n2826 0.04025
R13667 VSS.n5221 VSS.n2826 0.04025
R13668 VSS.n5222 VSS.n5221 0.04025
R13669 VSS.n5223 VSS.n5222 0.04025
R13670 VSS.n5223 VSS.n2824 0.04025
R13671 VSS.n5227 VSS.n2824 0.04025
R13672 VSS.n5228 VSS.n5227 0.04025
R13673 VSS.n5229 VSS.n5228 0.04025
R13674 VSS.n5229 VSS.n2822 0.04025
R13675 VSS.n5233 VSS.n2822 0.04025
R13676 VSS.n5234 VSS.n5233 0.04025
R13677 VSS.n5235 VSS.n5234 0.04025
R13678 VSS.n5235 VSS.n2820 0.04025
R13679 VSS.n5239 VSS.n2820 0.04025
R13680 VSS.n5240 VSS.n5239 0.04025
R13681 VSS.n5241 VSS.n5240 0.04025
R13682 VSS.n5241 VSS.n2818 0.04025
R13683 VSS.n5245 VSS.n2818 0.04025
R13684 VSS.n5246 VSS.n5245 0.04025
R13685 VSS.n5247 VSS.n5246 0.04025
R13686 VSS.n5247 VSS.n2816 0.04025
R13687 VSS.n5251 VSS.n2816 0.04025
R13688 VSS.n5252 VSS.n5251 0.04025
R13689 VSS.n5253 VSS.n5252 0.04025
R13690 VSS.n5253 VSS.n2814 0.04025
R13691 VSS.n5257 VSS.n2814 0.04025
R13692 VSS.n5258 VSS.n5257 0.04025
R13693 VSS.n5259 VSS.n5258 0.04025
R13694 VSS.n5259 VSS.n2812 0.04025
R13695 VSS.n5263 VSS.n2812 0.04025
R13696 VSS.n5264 VSS.n5263 0.04025
R13697 VSS.n5265 VSS.n5264 0.04025
R13698 VSS.n5265 VSS.n2810 0.04025
R13699 VSS.n5269 VSS.n2810 0.04025
R13700 VSS.n5270 VSS.n5269 0.04025
R13701 VSS.n5271 VSS.n5270 0.04025
R13702 VSS.n5271 VSS.n2808 0.04025
R13703 VSS.n5275 VSS.n2808 0.04025
R13704 VSS.n5276 VSS.n5275 0.04025
R13705 VSS.n5277 VSS.n5276 0.04025
R13706 VSS.n5277 VSS.n2806 0.04025
R13707 VSS.n5281 VSS.n2806 0.04025
R13708 VSS.n5282 VSS.n5281 0.04025
R13709 VSS.n5283 VSS.n5282 0.04025
R13710 VSS.n5283 VSS.n2804 0.04025
R13711 VSS.n5287 VSS.n2804 0.04025
R13712 VSS.n5288 VSS.n5287 0.04025
R13713 VSS.n5289 VSS.n5288 0.04025
R13714 VSS.n5289 VSS.n2802 0.04025
R13715 VSS.n5293 VSS.n2802 0.04025
R13716 VSS.n5294 VSS.n5293 0.04025
R13717 VSS.n5295 VSS.n5294 0.04025
R13718 VSS.n5295 VSS.n2800 0.04025
R13719 VSS.n5299 VSS.n2800 0.04025
R13720 VSS.n5300 VSS.n5299 0.04025
R13721 VSS.n5301 VSS.n5300 0.04025
R13722 VSS.n5301 VSS.n2798 0.04025
R13723 VSS.n5305 VSS.n2798 0.04025
R13724 VSS.n5306 VSS.n5305 0.04025
R13725 VSS.n5307 VSS.n5306 0.04025
R13726 VSS.n5307 VSS.n2796 0.04025
R13727 VSS.n5311 VSS.n2796 0.04025
R13728 VSS.n5312 VSS.n5311 0.04025
R13729 VSS.n5313 VSS.n5312 0.04025
R13730 VSS.n5313 VSS.n2794 0.04025
R13731 VSS.n5317 VSS.n2794 0.04025
R13732 VSS.n5318 VSS.n5317 0.04025
R13733 VSS.n5319 VSS.n5318 0.04025
R13734 VSS.n5319 VSS.n2792 0.04025
R13735 VSS.n5323 VSS.n2792 0.04025
R13736 VSS.n5324 VSS.n5323 0.04025
R13737 VSS.n5325 VSS.n5324 0.04025
R13738 VSS.n5325 VSS.n2790 0.04025
R13739 VSS.n5329 VSS.n2790 0.04025
R13740 VSS.n5330 VSS.n5329 0.04025
R13741 VSS.n5331 VSS.n5330 0.04025
R13742 VSS.n5331 VSS.n2788 0.04025
R13743 VSS.n5335 VSS.n2788 0.04025
R13744 VSS.n5336 VSS.n5335 0.04025
R13745 VSS.n5337 VSS.n5336 0.04025
R13746 VSS.n5337 VSS.n2786 0.04025
R13747 VSS.n5341 VSS.n2786 0.04025
R13748 VSS.n5342 VSS.n5341 0.04025
R13749 VSS.n5343 VSS.n5342 0.04025
R13750 VSS.n5343 VSS.n2784 0.04025
R13751 VSS.n5347 VSS.n2784 0.04025
R13752 VSS.n5348 VSS.n5347 0.04025
R13753 VSS.n5349 VSS.n5348 0.04025
R13754 VSS.n5349 VSS.n2782 0.04025
R13755 VSS.n5353 VSS.n2782 0.04025
R13756 VSS.n5354 VSS.n5353 0.04025
R13757 VSS.n5355 VSS.n5354 0.04025
R13758 VSS.n5355 VSS.n2780 0.04025
R13759 VSS.n5359 VSS.n2780 0.04025
R13760 VSS.n5360 VSS.n5359 0.04025
R13761 VSS.n5361 VSS.n5360 0.04025
R13762 VSS.n5361 VSS.n2778 0.04025
R13763 VSS.n5365 VSS.n2778 0.04025
R13764 VSS.n5366 VSS.n5365 0.04025
R13765 VSS.n5367 VSS.n5366 0.04025
R13766 VSS.n5367 VSS.n2776 0.04025
R13767 VSS.n5371 VSS.n2776 0.04025
R13768 VSS.n5372 VSS.n5371 0.04025
R13769 VSS.n5373 VSS.n5372 0.04025
R13770 VSS.n5373 VSS.n2774 0.04025
R13771 VSS.n5377 VSS.n2774 0.04025
R13772 VSS.n5378 VSS.n5377 0.04025
R13773 VSS.n5379 VSS.n5378 0.04025
R13774 VSS.n5379 VSS.n2772 0.04025
R13775 VSS.n5383 VSS.n2772 0.04025
R13776 VSS.n5384 VSS.n5383 0.04025
R13777 VSS.n5385 VSS.n5384 0.04025
R13778 VSS.n5385 VSS.n2770 0.04025
R13779 VSS.n5389 VSS.n2770 0.04025
R13780 VSS.n5390 VSS.n5389 0.04025
R13781 VSS.n5391 VSS.n5390 0.04025
R13782 VSS.n5391 VSS.n2768 0.04025
R13783 VSS.n5395 VSS.n2768 0.04025
R13784 VSS.n5396 VSS.n5395 0.04025
R13785 VSS.n5397 VSS.n5396 0.04025
R13786 VSS.n5397 VSS.n2766 0.04025
R13787 VSS.n5401 VSS.n2766 0.04025
R13788 VSS.n5402 VSS.n5401 0.04025
R13789 VSS.n5403 VSS.n5402 0.04025
R13790 VSS.n5403 VSS.n2764 0.04025
R13791 VSS.n5407 VSS.n2764 0.04025
R13792 VSS.n5408 VSS.n5407 0.04025
R13793 VSS.n5409 VSS.n5408 0.04025
R13794 VSS.n5409 VSS.n2762 0.04025
R13795 VSS.n5413 VSS.n2762 0.04025
R13796 VSS.n5414 VSS.n5413 0.04025
R13797 VSS.n5415 VSS.n5414 0.04025
R13798 VSS.n5415 VSS.n2760 0.04025
R13799 VSS.n5419 VSS.n2760 0.04025
R13800 VSS.n5420 VSS.n5419 0.04025
R13801 VSS.n5421 VSS.n5420 0.04025
R13802 VSS.n5421 VSS.n2758 0.04025
R13803 VSS.n5425 VSS.n2758 0.04025
R13804 VSS.n5426 VSS.n5425 0.04025
R13805 VSS.n5427 VSS.n5426 0.04025
R13806 VSS.n5427 VSS.n2756 0.04025
R13807 VSS.n5431 VSS.n2756 0.04025
R13808 VSS.n5432 VSS.n5431 0.04025
R13809 VSS.n5433 VSS.n5432 0.04025
R13810 VSS.n5433 VSS.n2754 0.04025
R13811 VSS.n5437 VSS.n2754 0.04025
R13812 VSS.n5438 VSS.n5437 0.04025
R13813 VSS.n5439 VSS.n5438 0.04025
R13814 VSS.n5439 VSS.n2752 0.04025
R13815 VSS.n5443 VSS.n2752 0.04025
R13816 VSS.n5444 VSS.n5443 0.04025
R13817 VSS.n5445 VSS.n5444 0.04025
R13818 VSS.n5445 VSS.n2750 0.04025
R13819 VSS.n5449 VSS.n2750 0.04025
R13820 VSS.n5450 VSS.n5449 0.04025
R13821 VSS.n5451 VSS.n5450 0.04025
R13822 VSS.n5451 VSS.n2748 0.04025
R13823 VSS.n5455 VSS.n2748 0.04025
R13824 VSS.n5456 VSS.n5455 0.04025
R13825 VSS.n5457 VSS.n5456 0.04025
R13826 VSS.n5457 VSS.n2746 0.04025
R13827 VSS.n5461 VSS.n2746 0.04025
R13828 VSS.n5462 VSS.n5461 0.04025
R13829 VSS.n5463 VSS.n5462 0.04025
R13830 VSS.n5463 VSS.n2744 0.04025
R13831 VSS.n5467 VSS.n2744 0.04025
R13832 VSS.n5468 VSS.n5467 0.04025
R13833 VSS.n4143 VSS.n4142 0.04025
R13834 VSS.n4143 VSS.n3183 0.04025
R13835 VSS.n4147 VSS.n3183 0.04025
R13836 VSS.n4148 VSS.n4147 0.04025
R13837 VSS.n4149 VSS.n4148 0.04025
R13838 VSS.n4149 VSS.n3181 0.04025
R13839 VSS.n4153 VSS.n3181 0.04025
R13840 VSS.n4154 VSS.n4153 0.04025
R13841 VSS.n4155 VSS.n4154 0.04025
R13842 VSS.n4155 VSS.n3179 0.04025
R13843 VSS.n4159 VSS.n3179 0.04025
R13844 VSS.n4160 VSS.n4159 0.04025
R13845 VSS.n4161 VSS.n4160 0.04025
R13846 VSS.n4161 VSS.n3177 0.04025
R13847 VSS.n4165 VSS.n3177 0.04025
R13848 VSS.n4166 VSS.n4165 0.04025
R13849 VSS.n4167 VSS.n4166 0.04025
R13850 VSS.n4167 VSS.n3175 0.04025
R13851 VSS.n4171 VSS.n3175 0.04025
R13852 VSS.n4172 VSS.n4171 0.04025
R13853 VSS.n4173 VSS.n4172 0.04025
R13854 VSS.n4173 VSS.n3173 0.04025
R13855 VSS.n4177 VSS.n3173 0.04025
R13856 VSS.n4178 VSS.n4177 0.04025
R13857 VSS.n4179 VSS.n4178 0.04025
R13858 VSS.n4179 VSS.n3171 0.04025
R13859 VSS.n4183 VSS.n3171 0.04025
R13860 VSS.n4184 VSS.n4183 0.04025
R13861 VSS.n4185 VSS.n4184 0.04025
R13862 VSS.n4185 VSS.n3169 0.04025
R13863 VSS.n4189 VSS.n3169 0.04025
R13864 VSS.n4190 VSS.n4189 0.04025
R13865 VSS.n4191 VSS.n4190 0.04025
R13866 VSS.n4191 VSS.n3167 0.04025
R13867 VSS.n4195 VSS.n3167 0.04025
R13868 VSS.n4196 VSS.n4195 0.04025
R13869 VSS.n4197 VSS.n4196 0.04025
R13870 VSS.n4197 VSS.n3165 0.04025
R13871 VSS.n4201 VSS.n3165 0.04025
R13872 VSS.n4202 VSS.n4201 0.04025
R13873 VSS.n4203 VSS.n4202 0.04025
R13874 VSS.n4203 VSS.n3163 0.04025
R13875 VSS.n4207 VSS.n3163 0.04025
R13876 VSS.n4208 VSS.n4207 0.04025
R13877 VSS.n4209 VSS.n4208 0.04025
R13878 VSS.n4209 VSS.n3161 0.04025
R13879 VSS.n4213 VSS.n3161 0.04025
R13880 VSS.n4214 VSS.n4213 0.04025
R13881 VSS.n4215 VSS.n4214 0.04025
R13882 VSS.n4215 VSS.n3159 0.04025
R13883 VSS.n4219 VSS.n3159 0.04025
R13884 VSS.n4220 VSS.n4219 0.04025
R13885 VSS.n4221 VSS.n4220 0.04025
R13886 VSS.n4221 VSS.n3157 0.04025
R13887 VSS.n4225 VSS.n3157 0.04025
R13888 VSS.n4226 VSS.n4225 0.04025
R13889 VSS.n4227 VSS.n4226 0.04025
R13890 VSS.n4227 VSS.n3155 0.04025
R13891 VSS.n4231 VSS.n3155 0.04025
R13892 VSS.n4232 VSS.n4231 0.04025
R13893 VSS.n4233 VSS.n4232 0.04025
R13894 VSS.n4233 VSS.n3153 0.04025
R13895 VSS.n4237 VSS.n3153 0.04025
R13896 VSS.n4238 VSS.n4237 0.04025
R13897 VSS.n4239 VSS.n4238 0.04025
R13898 VSS.n4239 VSS.n3151 0.04025
R13899 VSS.n4243 VSS.n3151 0.04025
R13900 VSS.n4244 VSS.n4243 0.04025
R13901 VSS.n4245 VSS.n4244 0.04025
R13902 VSS.n4245 VSS.n3149 0.04025
R13903 VSS.n4249 VSS.n3149 0.04025
R13904 VSS.n4250 VSS.n4249 0.04025
R13905 VSS.n4251 VSS.n4250 0.04025
R13906 VSS.n4251 VSS.n3147 0.04025
R13907 VSS.n4255 VSS.n3147 0.04025
R13908 VSS.n4256 VSS.n4255 0.04025
R13909 VSS.n4257 VSS.n4256 0.04025
R13910 VSS.n4257 VSS.n3145 0.04025
R13911 VSS.n4261 VSS.n3145 0.04025
R13912 VSS.n4262 VSS.n4261 0.04025
R13913 VSS.n4263 VSS.n4262 0.04025
R13914 VSS.n4263 VSS.n3143 0.04025
R13915 VSS.n4267 VSS.n3143 0.04025
R13916 VSS.n4268 VSS.n4267 0.04025
R13917 VSS.n4269 VSS.n4268 0.04025
R13918 VSS.n4269 VSS.n3141 0.04025
R13919 VSS.n4273 VSS.n3141 0.04025
R13920 VSS.n4274 VSS.n4273 0.04025
R13921 VSS.n4275 VSS.n4274 0.04025
R13922 VSS.n4275 VSS.n3139 0.04025
R13923 VSS.n4279 VSS.n3139 0.04025
R13924 VSS.n4280 VSS.n4279 0.04025
R13925 VSS.n4281 VSS.n4280 0.04025
R13926 VSS.n4281 VSS.n3137 0.04025
R13927 VSS.n4285 VSS.n3137 0.04025
R13928 VSS.n4286 VSS.n4285 0.04025
R13929 VSS.n4287 VSS.n4286 0.04025
R13930 VSS.n4287 VSS.n3135 0.04025
R13931 VSS.n4291 VSS.n3135 0.04025
R13932 VSS.n4292 VSS.n4291 0.04025
R13933 VSS.n4293 VSS.n4292 0.04025
R13934 VSS.n4293 VSS.n3133 0.04025
R13935 VSS.n4297 VSS.n3133 0.04025
R13936 VSS.n4298 VSS.n4297 0.04025
R13937 VSS.n4299 VSS.n4298 0.04025
R13938 VSS.n4299 VSS.n3131 0.04025
R13939 VSS.n4303 VSS.n3131 0.04025
R13940 VSS.n4304 VSS.n4303 0.04025
R13941 VSS.n4305 VSS.n4304 0.04025
R13942 VSS.n4305 VSS.n3129 0.04025
R13943 VSS.n4309 VSS.n3129 0.04025
R13944 VSS.n4310 VSS.n4309 0.04025
R13945 VSS.n4311 VSS.n4310 0.04025
R13946 VSS.n4311 VSS.n3127 0.04025
R13947 VSS.n4315 VSS.n3127 0.04025
R13948 VSS.n4316 VSS.n4315 0.04025
R13949 VSS.n4317 VSS.n4316 0.04025
R13950 VSS.n4317 VSS.n3125 0.04025
R13951 VSS.n4321 VSS.n3125 0.04025
R13952 VSS.n4322 VSS.n4321 0.04025
R13953 VSS.n4323 VSS.n4322 0.04025
R13954 VSS.n4323 VSS.n3123 0.04025
R13955 VSS.n4327 VSS.n3123 0.04025
R13956 VSS.n4328 VSS.n4327 0.04025
R13957 VSS.n4329 VSS.n4328 0.04025
R13958 VSS.n4329 VSS.n3121 0.04025
R13959 VSS.n4333 VSS.n3121 0.04025
R13960 VSS.n4334 VSS.n4333 0.04025
R13961 VSS.n4335 VSS.n4334 0.04025
R13962 VSS.n4335 VSS.n3119 0.04025
R13963 VSS.n4339 VSS.n3119 0.04025
R13964 VSS.n4340 VSS.n4339 0.04025
R13965 VSS.n4341 VSS.n4340 0.04025
R13966 VSS.n4341 VSS.n3117 0.04025
R13967 VSS.n4345 VSS.n3117 0.04025
R13968 VSS.n4346 VSS.n4345 0.04025
R13969 VSS.n4347 VSS.n4346 0.04025
R13970 VSS.n4347 VSS.n3115 0.04025
R13971 VSS.n4351 VSS.n3115 0.04025
R13972 VSS.n4352 VSS.n4351 0.04025
R13973 VSS.n4353 VSS.n4352 0.04025
R13974 VSS.n4353 VSS.n3113 0.04025
R13975 VSS.n4357 VSS.n3113 0.04025
R13976 VSS.n4358 VSS.n4357 0.04025
R13977 VSS.n4359 VSS.n4358 0.04025
R13978 VSS.n4359 VSS.n3111 0.04025
R13979 VSS.n4363 VSS.n3111 0.04025
R13980 VSS.n4364 VSS.n4363 0.04025
R13981 VSS.n4365 VSS.n4364 0.04025
R13982 VSS.n4365 VSS.n3109 0.04025
R13983 VSS.n4369 VSS.n3109 0.04025
R13984 VSS.n4370 VSS.n4369 0.04025
R13985 VSS.n4371 VSS.n4370 0.04025
R13986 VSS.n4371 VSS.n3107 0.04025
R13987 VSS.n4375 VSS.n3107 0.04025
R13988 VSS.n4376 VSS.n4375 0.04025
R13989 VSS.n4377 VSS.n4376 0.04025
R13990 VSS.n4377 VSS.n3105 0.04025
R13991 VSS.n4381 VSS.n3105 0.04025
R13992 VSS.n4382 VSS.n4381 0.04025
R13993 VSS.n4383 VSS.n4382 0.04025
R13994 VSS.n4383 VSS.n3103 0.04025
R13995 VSS.n4387 VSS.n3103 0.04025
R13996 VSS.n4388 VSS.n4387 0.04025
R13997 VSS.n4389 VSS.n4388 0.04025
R13998 VSS.n4389 VSS.n3101 0.04025
R13999 VSS.n4393 VSS.n3101 0.04025
R14000 VSS.n4394 VSS.n4393 0.04025
R14001 VSS.n4395 VSS.n4394 0.04025
R14002 VSS.n4395 VSS.n3099 0.04025
R14003 VSS.n4399 VSS.n3099 0.04025
R14004 VSS.n4400 VSS.n4399 0.04025
R14005 VSS.n4401 VSS.n4400 0.04025
R14006 VSS.n4401 VSS.n3097 0.04025
R14007 VSS.n4405 VSS.n3097 0.04025
R14008 VSS.n4406 VSS.n4405 0.04025
R14009 VSS.n4407 VSS.n4406 0.04025
R14010 VSS.n4407 VSS.n3095 0.04025
R14011 VSS.n4411 VSS.n3095 0.04025
R14012 VSS.n4412 VSS.n4411 0.04025
R14013 VSS.n4413 VSS.n4412 0.04025
R14014 VSS.n4413 VSS.n3093 0.04025
R14015 VSS.n4417 VSS.n3093 0.04025
R14016 VSS.n4418 VSS.n4417 0.04025
R14017 VSS.n4419 VSS.n4418 0.04025
R14018 VSS.n4419 VSS.n3091 0.04025
R14019 VSS.n4423 VSS.n3091 0.04025
R14020 VSS.n4424 VSS.n4423 0.04025
R14021 VSS.n4425 VSS.n4424 0.04025
R14022 VSS.n4425 VSS.n3089 0.04025
R14023 VSS.n4429 VSS.n3089 0.04025
R14024 VSS.n4430 VSS.n4429 0.04025
R14025 VSS.n4431 VSS.n4430 0.04025
R14026 VSS.n4431 VSS.n3087 0.04025
R14027 VSS.n4435 VSS.n3087 0.04025
R14028 VSS.n4436 VSS.n4435 0.04025
R14029 VSS.n4437 VSS.n4436 0.04025
R14030 VSS.n4437 VSS.n3085 0.04025
R14031 VSS.n4441 VSS.n3085 0.04025
R14032 VSS.n4442 VSS.n4441 0.04025
R14033 VSS.n4443 VSS.n4442 0.04025
R14034 VSS.n4443 VSS.n3083 0.04025
R14035 VSS.n4447 VSS.n3083 0.04025
R14036 VSS.n4448 VSS.n4447 0.04025
R14037 VSS.n4449 VSS.n4448 0.04025
R14038 VSS.n4449 VSS.n3081 0.04025
R14039 VSS.n4453 VSS.n3081 0.04025
R14040 VSS.n4454 VSS.n4453 0.04025
R14041 VSS.n4455 VSS.n4454 0.04025
R14042 VSS.n4455 VSS.n3079 0.04025
R14043 VSS.n4459 VSS.n3079 0.04025
R14044 VSS.n4460 VSS.n4459 0.04025
R14045 VSS.n4461 VSS.n4460 0.04025
R14046 VSS.n4461 VSS.n3077 0.04025
R14047 VSS.n4465 VSS.n3077 0.04025
R14048 VSS.n4466 VSS.n4465 0.04025
R14049 VSS.n4467 VSS.n4466 0.04025
R14050 VSS.n4467 VSS.n3075 0.04025
R14051 VSS.n4471 VSS.n3075 0.04025
R14052 VSS.n4472 VSS.n4471 0.04025
R14053 VSS.n4473 VSS.n4472 0.04025
R14054 VSS.n4473 VSS.n3073 0.04025
R14055 VSS.n4477 VSS.n3073 0.04025
R14056 VSS.n4478 VSS.n4477 0.04025
R14057 VSS.n4479 VSS.n4478 0.04025
R14058 VSS.n4479 VSS.n3071 0.04025
R14059 VSS.n4483 VSS.n3071 0.04025
R14060 VSS.n4484 VSS.n4483 0.04025
R14061 VSS.n4485 VSS.n4484 0.04025
R14062 VSS.n4485 VSS.n3069 0.04025
R14063 VSS.n4489 VSS.n3069 0.04025
R14064 VSS.n4490 VSS.n4489 0.04025
R14065 VSS.n4491 VSS.n4490 0.04025
R14066 VSS.n4491 VSS.n3067 0.04025
R14067 VSS.n4495 VSS.n3067 0.04025
R14068 VSS.n4496 VSS.n4495 0.04025
R14069 VSS.n4497 VSS.n4496 0.04025
R14070 VSS.n4497 VSS.n3065 0.04025
R14071 VSS.n4501 VSS.n3065 0.04025
R14072 VSS.n4502 VSS.n4501 0.04025
R14073 VSS.n4503 VSS.n4502 0.04025
R14074 VSS.n4503 VSS.n3063 0.04025
R14075 VSS.n4507 VSS.n3063 0.04025
R14076 VSS.n4508 VSS.n4507 0.04025
R14077 VSS.n4509 VSS.n4508 0.04025
R14078 VSS.n4509 VSS.n3061 0.04025
R14079 VSS.n4513 VSS.n3061 0.04025
R14080 VSS.n4514 VSS.n4513 0.04025
R14081 VSS.n4515 VSS.n4514 0.04025
R14082 VSS.n4515 VSS.n3059 0.04025
R14083 VSS.n4519 VSS.n3059 0.04025
R14084 VSS.n4520 VSS.n4519 0.04025
R14085 VSS.n4521 VSS.n4520 0.04025
R14086 VSS.n4521 VSS.n3057 0.04025
R14087 VSS.n4525 VSS.n3057 0.04025
R14088 VSS.n4526 VSS.n4525 0.04025
R14089 VSS.n4527 VSS.n4526 0.04025
R14090 VSS.n4527 VSS.n3055 0.04025
R14091 VSS.n4531 VSS.n3055 0.04025
R14092 VSS.n4532 VSS.n4531 0.04025
R14093 VSS.n4533 VSS.n4532 0.04025
R14094 VSS.n4533 VSS.n3053 0.04025
R14095 VSS.n4537 VSS.n3053 0.04025
R14096 VSS.n4538 VSS.n4537 0.04025
R14097 VSS.n4539 VSS.n4538 0.04025
R14098 VSS.n4539 VSS.n3051 0.04025
R14099 VSS.n4543 VSS.n3051 0.04025
R14100 VSS.n4544 VSS.n4543 0.04025
R14101 VSS.n4545 VSS.n4544 0.04025
R14102 VSS.n4545 VSS.n3049 0.04025
R14103 VSS.n4549 VSS.n3049 0.04025
R14104 VSS.n4550 VSS.n4549 0.04025
R14105 VSS.n4551 VSS.n4550 0.04025
R14106 VSS.n4551 VSS.n3047 0.04025
R14107 VSS.n4555 VSS.n3047 0.04025
R14108 VSS.n4556 VSS.n4555 0.04025
R14109 VSS.n4557 VSS.n4556 0.04025
R14110 VSS.n4557 VSS.n3045 0.04025
R14111 VSS.n4561 VSS.n3045 0.04025
R14112 VSS.n4562 VSS.n4561 0.04025
R14113 VSS.n4563 VSS.n4562 0.04025
R14114 VSS.n4563 VSS.n3043 0.04025
R14115 VSS.n4567 VSS.n3043 0.04025
R14116 VSS.n4568 VSS.n4567 0.04025
R14117 VSS.n4569 VSS.n4568 0.04025
R14118 VSS.n4569 VSS.n3041 0.04025
R14119 VSS.n4573 VSS.n3041 0.04025
R14120 VSS.n4574 VSS.n4573 0.04025
R14121 VSS.n4575 VSS.n4574 0.04025
R14122 VSS.n4575 VSS.n3039 0.04025
R14123 VSS.n4579 VSS.n3039 0.04025
R14124 VSS.n4580 VSS.n4579 0.04025
R14125 VSS.n4581 VSS.n4580 0.04025
R14126 VSS.n4581 VSS.n3037 0.04025
R14127 VSS.n4585 VSS.n3037 0.04025
R14128 VSS.n4586 VSS.n4585 0.04025
R14129 VSS.n4587 VSS.n4586 0.04025
R14130 VSS.n4587 VSS.n3035 0.04025
R14131 VSS.n4591 VSS.n3035 0.04025
R14132 VSS.n4592 VSS.n4591 0.04025
R14133 VSS.n4593 VSS.n4592 0.04025
R14134 VSS.n4593 VSS.n3033 0.04025
R14135 VSS.n4597 VSS.n3033 0.04025
R14136 VSS.n4598 VSS.n4597 0.04025
R14137 VSS.n4599 VSS.n4598 0.04025
R14138 VSS.n4599 VSS.n3031 0.04025
R14139 VSS.n4603 VSS.n3031 0.04025
R14140 VSS.n4604 VSS.n4603 0.04025
R14141 VSS.n4605 VSS.n4604 0.04025
R14142 VSS.n4605 VSS.n3029 0.04025
R14143 VSS.n4609 VSS.n3029 0.04025
R14144 VSS.n4610 VSS.n4609 0.04025
R14145 VSS.n4611 VSS.n4610 0.04025
R14146 VSS.n4611 VSS.n3027 0.04025
R14147 VSS.n4615 VSS.n3027 0.04025
R14148 VSS.n4616 VSS.n4615 0.04025
R14149 VSS.n4617 VSS.n4616 0.04025
R14150 VSS.n4617 VSS.n3025 0.04025
R14151 VSS.n4621 VSS.n3025 0.04025
R14152 VSS.n4622 VSS.n4621 0.04025
R14153 VSS.n4623 VSS.n4622 0.04025
R14154 VSS.n4623 VSS.n3023 0.04025
R14155 VSS.n4627 VSS.n3023 0.04025
R14156 VSS.n4628 VSS.n4627 0.04025
R14157 VSS.n4629 VSS.n4628 0.04025
R14158 VSS.n4629 VSS.n3021 0.04025
R14159 VSS.n4633 VSS.n3021 0.04025
R14160 VSS.n4634 VSS.n4633 0.04025
R14161 VSS.n4635 VSS.n4634 0.04025
R14162 VSS.n4635 VSS.n3019 0.04025
R14163 VSS.n4639 VSS.n3019 0.04025
R14164 VSS.n4640 VSS.n4639 0.04025
R14165 VSS.n4641 VSS.n4640 0.04025
R14166 VSS.n4641 VSS.n3017 0.04025
R14167 VSS.n4645 VSS.n3017 0.04025
R14168 VSS.n4646 VSS.n4645 0.04025
R14169 VSS.n4647 VSS.n4646 0.04025
R14170 VSS.n4647 VSS.n3015 0.04025
R14171 VSS.n4651 VSS.n3015 0.04025
R14172 VSS.n4652 VSS.n4651 0.04025
R14173 VSS.n4653 VSS.n4652 0.04025
R14174 VSS.n4653 VSS.n3013 0.04025
R14175 VSS.n4657 VSS.n3013 0.04025
R14176 VSS.n4658 VSS.n4657 0.04025
R14177 VSS.n4659 VSS.n4658 0.04025
R14178 VSS.n4659 VSS.n3011 0.04025
R14179 VSS.n4663 VSS.n3011 0.04025
R14180 VSS.n4664 VSS.n4663 0.04025
R14181 VSS.n4665 VSS.n4664 0.04025
R14182 VSS.n4665 VSS.n3009 0.04025
R14183 VSS.n4669 VSS.n3009 0.04025
R14184 VSS.n4670 VSS.n4669 0.04025
R14185 VSS.n4671 VSS.n4670 0.04025
R14186 VSS.n4671 VSS.n3007 0.04025
R14187 VSS.n4675 VSS.n3007 0.04025
R14188 VSS.n4676 VSS.n4675 0.04025
R14189 VSS.n4677 VSS.n4676 0.04025
R14190 VSS.n4677 VSS.n3005 0.04025
R14191 VSS.n4681 VSS.n3005 0.04025
R14192 VSS.n4682 VSS.n4681 0.04025
R14193 VSS.n4683 VSS.n4682 0.04025
R14194 VSS.n4683 VSS.n3003 0.04025
R14195 VSS.n4687 VSS.n3003 0.04025
R14196 VSS.n4688 VSS.n4687 0.04025
R14197 VSS.n4689 VSS.n4688 0.04025
R14198 VSS.n4689 VSS.n3001 0.04025
R14199 VSS.n4693 VSS.n3001 0.04025
R14200 VSS.n4694 VSS.n4693 0.04025
R14201 VSS.n4695 VSS.n4694 0.04025
R14202 VSS.n4695 VSS.n2999 0.04025
R14203 VSS.n4699 VSS.n2999 0.04025
R14204 VSS.n4700 VSS.n4699 0.04025
R14205 VSS.n4701 VSS.n4700 0.04025
R14206 VSS.n4701 VSS.n2997 0.04025
R14207 VSS.n4705 VSS.n2997 0.04025
R14208 VSS.n4706 VSS.n4705 0.04025
R14209 VSS.n4707 VSS.n4706 0.04025
R14210 VSS.n4707 VSS.n2995 0.04025
R14211 VSS.n4711 VSS.n2995 0.04025
R14212 VSS.n4712 VSS.n4711 0.04025
R14213 VSS.n4713 VSS.n4712 0.04025
R14214 VSS.n4713 VSS.n2993 0.04025
R14215 VSS.n4717 VSS.n2993 0.04025
R14216 VSS.n4718 VSS.n4717 0.04025
R14217 VSS.n4719 VSS.n4718 0.04025
R14218 VSS.n4719 VSS.n2991 0.04025
R14219 VSS.n4723 VSS.n2991 0.04025
R14220 VSS.n4724 VSS.n4723 0.04025
R14221 VSS.n4725 VSS.n4724 0.04025
R14222 VSS.n4725 VSS.n2989 0.04025
R14223 VSS.n4729 VSS.n2989 0.04025
R14224 VSS.n4730 VSS.n4729 0.04025
R14225 VSS.n4731 VSS.n4730 0.04025
R14226 VSS.n4731 VSS.n2987 0.04025
R14227 VSS.n4735 VSS.n2987 0.04025
R14228 VSS.n4736 VSS.n4735 0.04025
R14229 VSS.n4737 VSS.n4736 0.04025
R14230 VSS.n4737 VSS.n2985 0.04025
R14231 VSS.n4741 VSS.n2985 0.04025
R14232 VSS.n4742 VSS.n4741 0.04025
R14233 VSS.n4743 VSS.n4742 0.04025
R14234 VSS.n4743 VSS.n2983 0.04025
R14235 VSS.n4747 VSS.n2983 0.04025
R14236 VSS.n4748 VSS.n4747 0.04025
R14237 VSS.n4749 VSS.n4748 0.04025
R14238 VSS.n4749 VSS.n2981 0.04025
R14239 VSS.n4753 VSS.n2981 0.04025
R14240 VSS.n4754 VSS.n4753 0.04025
R14241 VSS.n4755 VSS.n4754 0.04025
R14242 VSS.n4755 VSS.n2979 0.04025
R14243 VSS.n4759 VSS.n2979 0.04025
R14244 VSS.n4760 VSS.n4759 0.04025
R14245 VSS.n4761 VSS.n4760 0.04025
R14246 VSS.n4761 VSS.n2977 0.04025
R14247 VSS.n4765 VSS.n2977 0.04025
R14248 VSS.n4766 VSS.n4765 0.04025
R14249 VSS.n4767 VSS.n4766 0.04025
R14250 VSS.n4767 VSS.n2975 0.04025
R14251 VSS.n4771 VSS.n2975 0.04025
R14252 VSS.n4772 VSS.n4771 0.04025
R14253 VSS.n4773 VSS.n4772 0.04025
R14254 VSS.n4773 VSS.n2973 0.04025
R14255 VSS.n4777 VSS.n2973 0.04025
R14256 VSS.n4778 VSS.n4777 0.04025
R14257 VSS.n4779 VSS.n4778 0.04025
R14258 VSS.n4779 VSS.n2971 0.04025
R14259 VSS.n4783 VSS.n2971 0.04025
R14260 VSS.n4784 VSS.n4783 0.04025
R14261 VSS.n4785 VSS.n4784 0.04025
R14262 VSS.n4785 VSS.n2969 0.04025
R14263 VSS.n4789 VSS.n2969 0.04025
R14264 VSS.n4790 VSS.n4789 0.04025
R14265 VSS.n4791 VSS.n4790 0.04025
R14266 VSS.n4791 VSS.n2967 0.04025
R14267 VSS.n4795 VSS.n2967 0.04025
R14268 VSS.n4796 VSS.n4795 0.04025
R14269 VSS.n4797 VSS.n4796 0.04025
R14270 VSS.n4797 VSS.n2965 0.04025
R14271 VSS.n4801 VSS.n2965 0.04025
R14272 VSS.n4802 VSS.n4801 0.04025
R14273 VSS.n4806 VSS.n4802 0.04025
R14274 VSS.n4806 VSS.n2963 0.04025
R14275 VSS.n4810 VSS.n2963 0.04025
R14276 VSS.n4811 VSS.n4810 0.04025
R14277 VSS.n4812 VSS.n4811 0.04025
R14278 VSS.n4812 VSS.n2961 0.04025
R14279 VSS.n4816 VSS.n2961 0.04025
R14280 VSS.n4817 VSS.n4816 0.04025
R14281 VSS.n4818 VSS.n4817 0.04025
R14282 VSS.n4818 VSS.n2959 0.04025
R14283 VSS.n4822 VSS.n2959 0.04025
R14284 VSS.n4823 VSS.n4822 0.04025
R14285 VSS.n4824 VSS.n4823 0.04025
R14286 VSS.n4824 VSS.n2957 0.04025
R14287 VSS.n4828 VSS.n2957 0.04025
R14288 VSS.n4829 VSS.n4828 0.04025
R14289 VSS.n4830 VSS.n4829 0.04025
R14290 VSS.n4830 VSS.n2955 0.04025
R14291 VSS.n4834 VSS.n2955 0.04025
R14292 VSS.n4835 VSS.n4834 0.04025
R14293 VSS.n4836 VSS.n4835 0.04025
R14294 VSS.n4836 VSS.n2953 0.04025
R14295 VSS.n4840 VSS.n2953 0.04025
R14296 VSS.n4841 VSS.n4840 0.04025
R14297 VSS.n4842 VSS.n4841 0.04025
R14298 VSS.n4842 VSS.n2951 0.04025
R14299 VSS.n4846 VSS.n2951 0.04025
R14300 VSS.n4847 VSS.n4846 0.04025
R14301 VSS.n4848 VSS.n4847 0.04025
R14302 VSS.n4848 VSS.n2949 0.04025
R14303 VSS.n4852 VSS.n2949 0.04025
R14304 VSS.n4853 VSS.n4852 0.04025
R14305 VSS.n4854 VSS.n4853 0.04025
R14306 VSS.n4854 VSS.n2947 0.04025
R14307 VSS.n4858 VSS.n2947 0.04025
R14308 VSS.n4859 VSS.n4858 0.04025
R14309 VSS.n4860 VSS.n4859 0.04025
R14310 VSS.n4860 VSS.n2945 0.04025
R14311 VSS.n4864 VSS.n2945 0.04025
R14312 VSS.n4865 VSS.n4864 0.04025
R14313 VSS.n4866 VSS.n4865 0.04025
R14314 VSS.n4866 VSS.n2943 0.04025
R14315 VSS.n4870 VSS.n2943 0.04025
R14316 VSS.n4871 VSS.n4870 0.04025
R14317 VSS.n4872 VSS.n4871 0.04025
R14318 VSS.n4872 VSS.n2941 0.04025
R14319 VSS.n4876 VSS.n2941 0.04025
R14320 VSS.n4877 VSS.n4876 0.04025
R14321 VSS.n4878 VSS.n4877 0.04025
R14322 VSS.n4878 VSS.n2939 0.04025
R14323 VSS.n4882 VSS.n2939 0.04025
R14324 VSS.n4883 VSS.n4882 0.04025
R14325 VSS.n4884 VSS.n4883 0.04025
R14326 VSS.n4884 VSS.n2937 0.04025
R14327 VSS.n4888 VSS.n2937 0.04025
R14328 VSS.n4889 VSS.n4888 0.04025
R14329 VSS.n4890 VSS.n4889 0.04025
R14330 VSS.n4890 VSS.n2935 0.04025
R14331 VSS.n4894 VSS.n2935 0.04025
R14332 VSS.n4895 VSS.n4894 0.04025
R14333 VSS.n4896 VSS.n4895 0.04025
R14334 VSS.n4896 VSS.n2933 0.04025
R14335 VSS.n4900 VSS.n2933 0.04025
R14336 VSS.n4901 VSS.n4900 0.04025
R14337 VSS.n4902 VSS.n4901 0.04025
R14338 VSS.n4902 VSS.n2931 0.04025
R14339 VSS.n4906 VSS.n2931 0.04025
R14340 VSS.n4907 VSS.n4906 0.04025
R14341 VSS.n4908 VSS.n4907 0.04025
R14342 VSS.n4908 VSS.n2929 0.04025
R14343 VSS.n4912 VSS.n2929 0.04025
R14344 VSS.n4913 VSS.n4912 0.04025
R14345 VSS.n4914 VSS.n4913 0.04025
R14346 VSS.n4914 VSS.n2927 0.04025
R14347 VSS.n4918 VSS.n2927 0.04025
R14348 VSS.n4919 VSS.n4918 0.04025
R14349 VSS.n4920 VSS.n4919 0.04025
R14350 VSS.n4920 VSS.n2925 0.04025
R14351 VSS.n4924 VSS.n2925 0.04025
R14352 VSS.n4925 VSS.n4924 0.04025
R14353 VSS.n4926 VSS.n4925 0.04025
R14354 VSS.n4926 VSS.n2923 0.04025
R14355 VSS.n4930 VSS.n2923 0.04025
R14356 VSS.n4931 VSS.n4930 0.04025
R14357 VSS.n4932 VSS.n4931 0.04025
R14358 VSS.n4932 VSS.n2921 0.04025
R14359 VSS.n4936 VSS.n2921 0.04025
R14360 VSS.n4937 VSS.n4936 0.04025
R14361 VSS.n4938 VSS.n4937 0.04025
R14362 VSS.n4938 VSS.n2919 0.04025
R14363 VSS.n4942 VSS.n2919 0.04025
R14364 VSS.n4943 VSS.n4942 0.04025
R14365 VSS.n4944 VSS.n4943 0.04025
R14366 VSS.n4944 VSS.n2917 0.04025
R14367 VSS.n4948 VSS.n2917 0.04025
R14368 VSS.n4949 VSS.n4948 0.04025
R14369 VSS.n4950 VSS.n4949 0.04025
R14370 VSS.n4950 VSS.n2915 0.04025
R14371 VSS.n4954 VSS.n2915 0.04025
R14372 VSS.n4955 VSS.n4954 0.04025
R14373 VSS.n4956 VSS.n4955 0.04025
R14374 VSS.n4956 VSS.n2913 0.04025
R14375 VSS.n4960 VSS.n2913 0.04025
R14376 VSS.n4961 VSS.n4960 0.04025
R14377 VSS.n4962 VSS.n4961 0.04025
R14378 VSS.n4962 VSS.n2911 0.04025
R14379 VSS.n4966 VSS.n2911 0.04025
R14380 VSS.n4967 VSS.n4966 0.04025
R14381 VSS.n4968 VSS.n4967 0.04025
R14382 VSS.n4968 VSS.n2909 0.04025
R14383 VSS.n4972 VSS.n2909 0.04025
R14384 VSS.n4973 VSS.n4972 0.04025
R14385 VSS.n4974 VSS.n4973 0.04025
R14386 VSS.n4974 VSS.n2907 0.04025
R14387 VSS.n4978 VSS.n2907 0.04025
R14388 VSS.n4979 VSS.n4978 0.04025
R14389 VSS.n4980 VSS.n4979 0.04025
R14390 VSS.n4980 VSS.n2905 0.04025
R14391 VSS.n4984 VSS.n2905 0.04025
R14392 VSS.n4985 VSS.n4984 0.04025
R14393 VSS.n4986 VSS.n4985 0.04025
R14394 VSS.n4986 VSS.n2903 0.04025
R14395 VSS.n4990 VSS.n2903 0.04025
R14396 VSS.n4991 VSS.n4990 0.04025
R14397 VSS.n4992 VSS.n4991 0.04025
R14398 VSS.n4992 VSS.n2901 0.04025
R14399 VSS.n4996 VSS.n2901 0.04025
R14400 VSS.n4997 VSS.n4996 0.04025
R14401 VSS.n4998 VSS.n4997 0.04025
R14402 VSS.n4998 VSS.n2899 0.04025
R14403 VSS.n5002 VSS.n2899 0.04025
R14404 VSS.n5003 VSS.n5002 0.04025
R14405 VSS.n5004 VSS.n5003 0.04025
R14406 VSS.n5004 VSS.n2897 0.04025
R14407 VSS.n5008 VSS.n2897 0.04025
R14408 VSS.n5009 VSS.n5008 0.04025
R14409 VSS.n5010 VSS.n5009 0.04025
R14410 VSS.n5010 VSS.n2895 0.04025
R14411 VSS.n5014 VSS.n2895 0.04025
R14412 VSS.n5015 VSS.n5014 0.04025
R14413 VSS.n5016 VSS.n5015 0.04025
R14414 VSS.n5016 VSS.n2893 0.04025
R14415 VSS.n5020 VSS.n2893 0.04025
R14416 VSS.n5021 VSS.n5020 0.04025
R14417 VSS.n5022 VSS.n5021 0.04025
R14418 VSS.n5022 VSS.n2891 0.04025
R14419 VSS.n5026 VSS.n2891 0.04025
R14420 VSS.n5027 VSS.n5026 0.04025
R14421 VSS.n5028 VSS.n5027 0.04025
R14422 VSS.n5028 VSS.n2889 0.04025
R14423 VSS.n5032 VSS.n2889 0.04025
R14424 VSS.n5033 VSS.n5032 0.04025
R14425 VSS.n5034 VSS.n5033 0.04025
R14426 VSS.n5034 VSS.n2887 0.04025
R14427 VSS.n5038 VSS.n2887 0.04025
R14428 VSS.n5039 VSS.n5038 0.04025
R14429 VSS.n5040 VSS.n5039 0.04025
R14430 VSS.n5040 VSS.n2885 0.04025
R14431 VSS.n5044 VSS.n2885 0.04025
R14432 VSS.n5045 VSS.n5044 0.04025
R14433 VSS.n5046 VSS.n5045 0.04025
R14434 VSS.n5046 VSS.n2883 0.04025
R14435 VSS.n5050 VSS.n2883 0.04025
R14436 VSS.n5051 VSS.n5050 0.04025
R14437 VSS.n5052 VSS.n5051 0.04025
R14438 VSS.n5052 VSS.n2881 0.04025
R14439 VSS.n5056 VSS.n2881 0.04025
R14440 VSS.n5057 VSS.n5056 0.04025
R14441 VSS.n5058 VSS.n5057 0.04025
R14442 VSS.n5058 VSS.n2879 0.04025
R14443 VSS.n5062 VSS.n2879 0.04025
R14444 VSS.n5063 VSS.n5062 0.04025
R14445 VSS.n5064 VSS.n5063 0.04025
R14446 VSS.n5064 VSS.n2877 0.04025
R14447 VSS.n5068 VSS.n2877 0.04025
R14448 VSS.n5069 VSS.n5068 0.04025
R14449 VSS.n5070 VSS.n5069 0.04025
R14450 VSS.n5070 VSS.n2875 0.04025
R14451 VSS.n5074 VSS.n2875 0.04025
R14452 VSS.n5075 VSS.n5074 0.04025
R14453 VSS.n5076 VSS.n5075 0.04025
R14454 VSS.n5076 VSS.n2873 0.04025
R14455 VSS.n5080 VSS.n2873 0.04025
R14456 VSS.n5081 VSS.n5080 0.04025
R14457 VSS.n5082 VSS.n5081 0.04025
R14458 VSS.n5082 VSS.n2871 0.04025
R14459 VSS.n5086 VSS.n2871 0.04025
R14460 VSS.n5087 VSS.n5086 0.04025
R14461 VSS.n5088 VSS.n5087 0.04025
R14462 VSS.n5088 VSS.n2869 0.04025
R14463 VSS.n5092 VSS.n2869 0.04025
R14464 VSS.n5093 VSS.n5092 0.04025
R14465 VSS.n5094 VSS.n5093 0.04025
R14466 VSS.n5094 VSS.n2867 0.04025
R14467 VSS.n5098 VSS.n2867 0.04025
R14468 VSS.n5099 VSS.n5098 0.04025
R14469 VSS.n5100 VSS.n5099 0.04025
R14470 VSS.n5100 VSS.n2865 0.04025
R14471 VSS.n5104 VSS.n2865 0.04025
R14472 VSS.n5105 VSS.n5104 0.04025
R14473 VSS.n5106 VSS.n5105 0.04025
R14474 VSS.n5106 VSS.n2863 0.04025
R14475 VSS.n5110 VSS.n2863 0.04025
R14476 VSS.n5111 VSS.n5110 0.04025
R14477 VSS.n5112 VSS.n5111 0.04025
R14478 VSS.n5112 VSS.n2861 0.04025
R14479 VSS.n5116 VSS.n2861 0.04025
R14480 VSS.n5117 VSS.n5116 0.04025
R14481 VSS.n5118 VSS.n5117 0.04025
R14482 VSS.n5118 VSS.n2859 0.04025
R14483 VSS.n5122 VSS.n2859 0.04025
R14484 VSS.n5123 VSS.n5122 0.04025
R14485 VSS.n5124 VSS.n5123 0.04025
R14486 VSS.n5124 VSS.n2857 0.04025
R14487 VSS.n5128 VSS.n2857 0.04025
R14488 VSS.n5129 VSS.n5128 0.04025
R14489 VSS.n5130 VSS.n5129 0.04025
R14490 VSS.n5130 VSS.n2855 0.04025
R14491 VSS.n5134 VSS.n2855 0.04025
R14492 VSS.n5135 VSS.n5134 0.04025
R14493 VSS.n5136 VSS.n5135 0.04025
R14494 VSS.n5136 VSS.n2853 0.04025
R14495 VSS.n5140 VSS.n2853 0.04025
R14496 VSS.n5141 VSS.n5140 0.04025
R14497 VSS.n5142 VSS.n5141 0.04025
R14498 VSS.n5142 VSS.n2851 0.04025
R14499 VSS.n5146 VSS.n2851 0.04025
R14500 VSS.n5147 VSS.n5146 0.04025
R14501 VSS.n5148 VSS.n5147 0.04025
R14502 VSS.n5148 VSS.n2849 0.04025
R14503 VSS.n5152 VSS.n2849 0.04025
R14504 VSS.n5153 VSS.n5152 0.04025
R14505 VSS.n5154 VSS.n5153 0.04025
R14506 VSS.n5154 VSS.n2847 0.04025
R14507 VSS.n5158 VSS.n2847 0.04025
R14508 VSS.n5159 VSS.n5158 0.04025
R14509 VSS.n5160 VSS.n5159 0.04025
R14510 VSS.n5160 VSS.n2845 0.04025
R14511 VSS.n5164 VSS.n2845 0.04025
R14512 VSS.n5165 VSS.n5164 0.04025
R14513 VSS.n5166 VSS.n5165 0.04025
R14514 VSS.n5166 VSS.n2843 0.04025
R14515 VSS.n5170 VSS.n2843 0.04025
R14516 VSS.n5171 VSS.n5170 0.04025
R14517 VSS.n5172 VSS.n5171 0.04025
R14518 VSS.n5172 VSS.n2841 0.04025
R14519 VSS.n5176 VSS.n2841 0.04025
R14520 VSS.n5177 VSS.n5176 0.04025
R14521 VSS.n5178 VSS.n5177 0.04025
R14522 VSS.n5178 VSS.n2839 0.04025
R14523 VSS.n5182 VSS.n2839 0.04025
R14524 VSS.n5183 VSS.n5182 0.04025
R14525 VSS.n5184 VSS.n5183 0.04025
R14526 VSS.n5184 VSS.n2837 0.04025
R14527 VSS.n5188 VSS.n2837 0.04025
R14528 VSS.n5189 VSS.n5188 0.04025
R14529 VSS.n5190 VSS.n5189 0.04025
R14530 VSS.n5190 VSS.n2835 0.04025
R14531 VSS.n5194 VSS.n2835 0.04025
R14532 VSS.n5195 VSS.n5194 0.04025
R14533 VSS.n5196 VSS.n5195 0.04025
R14534 VSS.n5196 VSS.n2833 0.04025
R14535 VSS.n5200 VSS.n2833 0.04025
R14536 VSS.n5201 VSS.n5200 0.04025
R14537 VSS.n5202 VSS.n5201 0.04025
R14538 VSS.n5202 VSS.n2831 0.04025
R14539 VSS.n5206 VSS.n2831 0.04025
R14540 VSS.n5207 VSS.n5206 0.04025
R14541 VSS.n5208 VSS.n5207 0.04025
R14542 VSS.n5208 VSS.n2829 0.04025
R14543 VSS.n5212 VSS.n2829 0.04025
R14544 VSS.n5213 VSS.n5212 0.04025
R14545 VSS.n5214 VSS.n5213 0.04025
R14546 VSS.n5214 VSS.n2827 0.04025
R14547 VSS.n5218 VSS.n2827 0.04025
R14548 VSS.n5219 VSS.n5218 0.04025
R14549 VSS.n5220 VSS.n5219 0.04025
R14550 VSS.n5220 VSS.n2825 0.04025
R14551 VSS.n5224 VSS.n2825 0.04025
R14552 VSS.n5225 VSS.n5224 0.04025
R14553 VSS.n5226 VSS.n5225 0.04025
R14554 VSS.n5226 VSS.n2823 0.04025
R14555 VSS.n5230 VSS.n2823 0.04025
R14556 VSS.n5231 VSS.n5230 0.04025
R14557 VSS.n5232 VSS.n5231 0.04025
R14558 VSS.n5232 VSS.n2821 0.04025
R14559 VSS.n5236 VSS.n2821 0.04025
R14560 VSS.n5237 VSS.n5236 0.04025
R14561 VSS.n5238 VSS.n5237 0.04025
R14562 VSS.n5238 VSS.n2819 0.04025
R14563 VSS.n5242 VSS.n2819 0.04025
R14564 VSS.n5243 VSS.n5242 0.04025
R14565 VSS.n5244 VSS.n5243 0.04025
R14566 VSS.n5244 VSS.n2817 0.04025
R14567 VSS.n5248 VSS.n2817 0.04025
R14568 VSS.n5249 VSS.n5248 0.04025
R14569 VSS.n5250 VSS.n5249 0.04025
R14570 VSS.n5250 VSS.n2815 0.04025
R14571 VSS.n5254 VSS.n2815 0.04025
R14572 VSS.n5255 VSS.n5254 0.04025
R14573 VSS.n5256 VSS.n5255 0.04025
R14574 VSS.n5256 VSS.n2813 0.04025
R14575 VSS.n5260 VSS.n2813 0.04025
R14576 VSS.n5261 VSS.n5260 0.04025
R14577 VSS.n5262 VSS.n5261 0.04025
R14578 VSS.n5262 VSS.n2811 0.04025
R14579 VSS.n5266 VSS.n2811 0.04025
R14580 VSS.n5267 VSS.n5266 0.04025
R14581 VSS.n5268 VSS.n5267 0.04025
R14582 VSS.n5268 VSS.n2809 0.04025
R14583 VSS.n5272 VSS.n2809 0.04025
R14584 VSS.n5273 VSS.n5272 0.04025
R14585 VSS.n5274 VSS.n5273 0.04025
R14586 VSS.n5274 VSS.n2807 0.04025
R14587 VSS.n5278 VSS.n2807 0.04025
R14588 VSS.n5279 VSS.n5278 0.04025
R14589 VSS.n5280 VSS.n5279 0.04025
R14590 VSS.n5280 VSS.n2805 0.04025
R14591 VSS.n5284 VSS.n2805 0.04025
R14592 VSS.n5285 VSS.n5284 0.04025
R14593 VSS.n5286 VSS.n5285 0.04025
R14594 VSS.n5286 VSS.n2803 0.04025
R14595 VSS.n5290 VSS.n2803 0.04025
R14596 VSS.n5291 VSS.n5290 0.04025
R14597 VSS.n5292 VSS.n5291 0.04025
R14598 VSS.n5292 VSS.n2801 0.04025
R14599 VSS.n5296 VSS.n2801 0.04025
R14600 VSS.n5297 VSS.n5296 0.04025
R14601 VSS.n5298 VSS.n5297 0.04025
R14602 VSS.n5298 VSS.n2799 0.04025
R14603 VSS.n5302 VSS.n2799 0.04025
R14604 VSS.n5303 VSS.n5302 0.04025
R14605 VSS.n5304 VSS.n5303 0.04025
R14606 VSS.n5304 VSS.n2797 0.04025
R14607 VSS.n5308 VSS.n2797 0.04025
R14608 VSS.n5309 VSS.n5308 0.04025
R14609 VSS.n5310 VSS.n5309 0.04025
R14610 VSS.n5310 VSS.n2795 0.04025
R14611 VSS.n5314 VSS.n2795 0.04025
R14612 VSS.n5315 VSS.n5314 0.04025
R14613 VSS.n5316 VSS.n5315 0.04025
R14614 VSS.n5316 VSS.n2793 0.04025
R14615 VSS.n5320 VSS.n2793 0.04025
R14616 VSS.n5321 VSS.n5320 0.04025
R14617 VSS.n5322 VSS.n5321 0.04025
R14618 VSS.n5322 VSS.n2791 0.04025
R14619 VSS.n5326 VSS.n2791 0.04025
R14620 VSS.n5327 VSS.n5326 0.04025
R14621 VSS.n5328 VSS.n5327 0.04025
R14622 VSS.n5328 VSS.n2789 0.04025
R14623 VSS.n5332 VSS.n2789 0.04025
R14624 VSS.n5333 VSS.n5332 0.04025
R14625 VSS.n5334 VSS.n5333 0.04025
R14626 VSS.n5334 VSS.n2787 0.04025
R14627 VSS.n5338 VSS.n2787 0.04025
R14628 VSS.n5339 VSS.n5338 0.04025
R14629 VSS.n5340 VSS.n5339 0.04025
R14630 VSS.n5340 VSS.n2785 0.04025
R14631 VSS.n5344 VSS.n2785 0.04025
R14632 VSS.n5345 VSS.n5344 0.04025
R14633 VSS.n5346 VSS.n5345 0.04025
R14634 VSS.n5346 VSS.n2783 0.04025
R14635 VSS.n5350 VSS.n2783 0.04025
R14636 VSS.n5351 VSS.n5350 0.04025
R14637 VSS.n5352 VSS.n5351 0.04025
R14638 VSS.n5352 VSS.n2781 0.04025
R14639 VSS.n5356 VSS.n2781 0.04025
R14640 VSS.n5357 VSS.n5356 0.04025
R14641 VSS.n5358 VSS.n5357 0.04025
R14642 VSS.n5358 VSS.n2779 0.04025
R14643 VSS.n5362 VSS.n2779 0.04025
R14644 VSS.n5363 VSS.n5362 0.04025
R14645 VSS.n5364 VSS.n5363 0.04025
R14646 VSS.n5364 VSS.n2777 0.04025
R14647 VSS.n5368 VSS.n2777 0.04025
R14648 VSS.n5369 VSS.n5368 0.04025
R14649 VSS.n5370 VSS.n5369 0.04025
R14650 VSS.n5370 VSS.n2775 0.04025
R14651 VSS.n5374 VSS.n2775 0.04025
R14652 VSS.n5375 VSS.n5374 0.04025
R14653 VSS.n5376 VSS.n5375 0.04025
R14654 VSS.n5376 VSS.n2773 0.04025
R14655 VSS.n5380 VSS.n2773 0.04025
R14656 VSS.n5381 VSS.n5380 0.04025
R14657 VSS.n5382 VSS.n5381 0.04025
R14658 VSS.n5382 VSS.n2771 0.04025
R14659 VSS.n5386 VSS.n2771 0.04025
R14660 VSS.n5387 VSS.n5386 0.04025
R14661 VSS.n5388 VSS.n5387 0.04025
R14662 VSS.n5388 VSS.n2769 0.04025
R14663 VSS.n5392 VSS.n2769 0.04025
R14664 VSS.n5393 VSS.n5392 0.04025
R14665 VSS.n5394 VSS.n5393 0.04025
R14666 VSS.n5394 VSS.n2767 0.04025
R14667 VSS.n5398 VSS.n2767 0.04025
R14668 VSS.n5399 VSS.n5398 0.04025
R14669 VSS.n5400 VSS.n5399 0.04025
R14670 VSS.n5400 VSS.n2765 0.04025
R14671 VSS.n5404 VSS.n2765 0.04025
R14672 VSS.n5405 VSS.n5404 0.04025
R14673 VSS.n5406 VSS.n5405 0.04025
R14674 VSS.n5406 VSS.n2763 0.04025
R14675 VSS.n5410 VSS.n2763 0.04025
R14676 VSS.n5411 VSS.n5410 0.04025
R14677 VSS.n5412 VSS.n5411 0.04025
R14678 VSS.n5412 VSS.n2761 0.04025
R14679 VSS.n5416 VSS.n2761 0.04025
R14680 VSS.n5417 VSS.n5416 0.04025
R14681 VSS.n5418 VSS.n5417 0.04025
R14682 VSS.n5418 VSS.n2759 0.04025
R14683 VSS.n5422 VSS.n2759 0.04025
R14684 VSS.n5423 VSS.n5422 0.04025
R14685 VSS.n5424 VSS.n5423 0.04025
R14686 VSS.n5424 VSS.n2757 0.04025
R14687 VSS.n5428 VSS.n2757 0.04025
R14688 VSS.n5429 VSS.n5428 0.04025
R14689 VSS.n5430 VSS.n5429 0.04025
R14690 VSS.n5430 VSS.n2755 0.04025
R14691 VSS.n5434 VSS.n2755 0.04025
R14692 VSS.n5435 VSS.n5434 0.04025
R14693 VSS.n5436 VSS.n5435 0.04025
R14694 VSS.n5436 VSS.n2753 0.04025
R14695 VSS.n5440 VSS.n2753 0.04025
R14696 VSS.n5441 VSS.n5440 0.04025
R14697 VSS.n5442 VSS.n5441 0.04025
R14698 VSS.n5442 VSS.n2751 0.04025
R14699 VSS.n5446 VSS.n2751 0.04025
R14700 VSS.n5447 VSS.n5446 0.04025
R14701 VSS.n5448 VSS.n5447 0.04025
R14702 VSS.n5448 VSS.n2749 0.04025
R14703 VSS.n5452 VSS.n2749 0.04025
R14704 VSS.n5453 VSS.n5452 0.04025
R14705 VSS.n5454 VSS.n5453 0.04025
R14706 VSS.n5454 VSS.n2747 0.04025
R14707 VSS.n5458 VSS.n2747 0.04025
R14708 VSS.n5459 VSS.n5458 0.04025
R14709 VSS.n5460 VSS.n5459 0.04025
R14710 VSS.n5460 VSS.n2745 0.04025
R14711 VSS.n5464 VSS.n2745 0.04025
R14712 VSS.n5465 VSS.n5464 0.04025
R14713 VSS.n5466 VSS.n5465 0.04025
R14714 VSS.n5466 VSS.n2743 0.04025
R14715 VSS.n5471 VSS.n5470 0.04025
R14716 VSS.n5472 VSS.n5471 0.04025
R14717 VSS.n5472 VSS.n2741 0.04025
R14718 VSS.n5476 VSS.n2741 0.04025
R14719 VSS.n5477 VSS.n5476 0.04025
R14720 VSS.n5478 VSS.n5477 0.04025
R14721 VSS.n5478 VSS.n2739 0.04025
R14722 VSS.n5482 VSS.n2739 0.04025
R14723 VSS.n5483 VSS.n5482 0.04025
R14724 VSS.n5484 VSS.n5483 0.04025
R14725 VSS.n5484 VSS.n2737 0.04025
R14726 VSS.n5488 VSS.n2737 0.04025
R14727 VSS.n5489 VSS.n5488 0.04025
R14728 VSS.n5490 VSS.n5489 0.04025
R14729 VSS.n5490 VSS.n2735 0.04025
R14730 VSS.n5494 VSS.n2735 0.04025
R14731 VSS.n5495 VSS.n5494 0.04025
R14732 VSS.n5496 VSS.n5495 0.04025
R14733 VSS.n5496 VSS.n2733 0.04025
R14734 VSS.n5500 VSS.n2733 0.04025
R14735 VSS.n5501 VSS.n5500 0.04025
R14736 VSS.n5502 VSS.n5501 0.04025
R14737 VSS.n5502 VSS.n2731 0.04025
R14738 VSS.n5506 VSS.n2731 0.04025
R14739 VSS.n5507 VSS.n5506 0.04025
R14740 VSS.n5508 VSS.n5507 0.04025
R14741 VSS.n5508 VSS.n2729 0.04025
R14742 VSS.n5512 VSS.n2729 0.04025
R14743 VSS.n5513 VSS.n5512 0.04025
R14744 VSS.n5514 VSS.n5513 0.04025
R14745 VSS.n5514 VSS.n2727 0.04025
R14746 VSS.n5518 VSS.n2727 0.04025
R14747 VSS.n5519 VSS.n5518 0.04025
R14748 VSS.n5520 VSS.n5519 0.04025
R14749 VSS.n5520 VSS.n2725 0.04025
R14750 VSS.n5524 VSS.n2725 0.04025
R14751 VSS.n5525 VSS.n5524 0.04025
R14752 VSS.n5526 VSS.n5525 0.04025
R14753 VSS.n5526 VSS.n2723 0.04025
R14754 VSS.n5530 VSS.n2723 0.04025
R14755 VSS.n5531 VSS.n5530 0.04025
R14756 VSS.n5532 VSS.n5531 0.04025
R14757 VSS.n5532 VSS.n2721 0.04025
R14758 VSS.n5536 VSS.n2721 0.04025
R14759 VSS.n5537 VSS.n5536 0.04025
R14760 VSS.n5538 VSS.n5537 0.04025
R14761 VSS.n5538 VSS.n2719 0.04025
R14762 VSS.n5542 VSS.n2719 0.04025
R14763 VSS.n5543 VSS.n5542 0.04025
R14764 VSS.n5544 VSS.n5543 0.04025
R14765 VSS.n5544 VSS.n2717 0.04025
R14766 VSS.n5548 VSS.n2717 0.04025
R14767 VSS.n5549 VSS.n5548 0.04025
R14768 VSS.n5550 VSS.n5549 0.04025
R14769 VSS.n5550 VSS.n2715 0.04025
R14770 VSS.n5554 VSS.n2715 0.04025
R14771 VSS.n5555 VSS.n5554 0.04025
R14772 VSS.n5556 VSS.n5555 0.04025
R14773 VSS.n5556 VSS.n2713 0.04025
R14774 VSS.n5560 VSS.n2713 0.04025
R14775 VSS.n5561 VSS.n5560 0.04025
R14776 VSS.n5562 VSS.n5561 0.04025
R14777 VSS.n5562 VSS.n2711 0.04025
R14778 VSS.n5566 VSS.n2711 0.04025
R14779 VSS.n5567 VSS.n5566 0.04025
R14780 VSS.n5568 VSS.n5567 0.04025
R14781 VSS.n5568 VSS.n2709 0.04025
R14782 VSS.n5572 VSS.n2709 0.04025
R14783 VSS.n5573 VSS.n5572 0.04025
R14784 VSS.n5574 VSS.n5573 0.04025
R14785 VSS.n5574 VSS.n2707 0.04025
R14786 VSS.n5578 VSS.n2707 0.04025
R14787 VSS.n5579 VSS.n5578 0.04025
R14788 VSS.n5580 VSS.n5579 0.04025
R14789 VSS.n5580 VSS.n2705 0.04025
R14790 VSS.n5584 VSS.n2705 0.04025
R14791 VSS.n5585 VSS.n5584 0.04025
R14792 VSS.n5586 VSS.n5585 0.04025
R14793 VSS.n5586 VSS.n2703 0.04025
R14794 VSS.n5590 VSS.n2703 0.04025
R14795 VSS.n5591 VSS.n5590 0.04025
R14796 VSS.n5592 VSS.n5591 0.04025
R14797 VSS.n5592 VSS.n2701 0.04025
R14798 VSS.n5596 VSS.n2701 0.04025
R14799 VSS.n5597 VSS.n5596 0.04025
R14800 VSS.n5598 VSS.n5597 0.04025
R14801 VSS.n5598 VSS.n2699 0.04025
R14802 VSS.n5602 VSS.n2699 0.04025
R14803 VSS.n5603 VSS.n5602 0.04025
R14804 VSS.n5604 VSS.n5603 0.04025
R14805 VSS.n5604 VSS.n2697 0.04025
R14806 VSS.n5608 VSS.n2697 0.04025
R14807 VSS.n5609 VSS.n5608 0.04025
R14808 VSS.n5610 VSS.n5609 0.04025
R14809 VSS.n5610 VSS.n2695 0.04025
R14810 VSS.n5614 VSS.n2695 0.04025
R14811 VSS.n5615 VSS.n5614 0.04025
R14812 VSS.n5616 VSS.n5615 0.04025
R14813 VSS.n5616 VSS.n2693 0.04025
R14814 VSS.n5620 VSS.n2693 0.04025
R14815 VSS.n5621 VSS.n5620 0.04025
R14816 VSS.n5622 VSS.n5621 0.04025
R14817 VSS.n5622 VSS.n2691 0.04025
R14818 VSS.n5626 VSS.n2691 0.04025
R14819 VSS.n5627 VSS.n5626 0.04025
R14820 VSS.n5628 VSS.n5627 0.04025
R14821 VSS.n5628 VSS.n2689 0.04025
R14822 VSS.n5632 VSS.n2689 0.04025
R14823 VSS.n5633 VSS.n5632 0.04025
R14824 VSS.n5634 VSS.n5633 0.04025
R14825 VSS.n5634 VSS.n2687 0.04025
R14826 VSS.n5638 VSS.n2687 0.04025
R14827 VSS.n5639 VSS.n5638 0.04025
R14828 VSS.n5640 VSS.n5639 0.04025
R14829 VSS.n5640 VSS.n2685 0.04025
R14830 VSS.n5644 VSS.n2685 0.04025
R14831 VSS.n5645 VSS.n5644 0.04025
R14832 VSS.n5646 VSS.n5645 0.04025
R14833 VSS.n5646 VSS.n2683 0.04025
R14834 VSS.n5650 VSS.n2683 0.04025
R14835 VSS.n5651 VSS.n5650 0.04025
R14836 VSS.n5652 VSS.n5651 0.04025
R14837 VSS.n5652 VSS.n2681 0.04025
R14838 VSS.n5656 VSS.n2681 0.04025
R14839 VSS.n5657 VSS.n5656 0.04025
R14840 VSS.n5658 VSS.n5657 0.04025
R14841 VSS.n5658 VSS.n2679 0.04025
R14842 VSS.n5662 VSS.n2679 0.04025
R14843 VSS.n5663 VSS.n5662 0.04025
R14844 VSS.n5664 VSS.n5663 0.04025
R14845 VSS.n5664 VSS.n2677 0.04025
R14846 VSS.n5668 VSS.n2677 0.04025
R14847 VSS.n5669 VSS.n5668 0.04025
R14848 VSS.n5670 VSS.n5669 0.04025
R14849 VSS.n5670 VSS.n2675 0.04025
R14850 VSS.n5674 VSS.n2675 0.04025
R14851 VSS.n5675 VSS.n5674 0.04025
R14852 VSS.n5676 VSS.n5675 0.04025
R14853 VSS.n5676 VSS.n2673 0.04025
R14854 VSS.n5680 VSS.n2673 0.04025
R14855 VSS.n5681 VSS.n5680 0.04025
R14856 VSS.n5682 VSS.n5681 0.04025
R14857 VSS.n5682 VSS.n2671 0.04025
R14858 VSS.n5686 VSS.n2671 0.04025
R14859 VSS.n5687 VSS.n5686 0.04025
R14860 VSS.n5688 VSS.n5687 0.04025
R14861 VSS.n5688 VSS.n2669 0.04025
R14862 VSS.n5692 VSS.n2669 0.04025
R14863 VSS.n5693 VSS.n5692 0.04025
R14864 VSS.n5694 VSS.n5693 0.04025
R14865 VSS.n5694 VSS.n2667 0.04025
R14866 VSS.n5698 VSS.n2667 0.04025
R14867 VSS.n5699 VSS.n5698 0.04025
R14868 VSS.n5700 VSS.n5699 0.04025
R14869 VSS.n5700 VSS.n2665 0.04025
R14870 VSS.n5704 VSS.n2665 0.04025
R14871 VSS.n5705 VSS.n5704 0.04025
R14872 VSS.n5706 VSS.n5705 0.04025
R14873 VSS.n5706 VSS.n2663 0.04025
R14874 VSS.n5710 VSS.n2663 0.04025
R14875 VSS.n5711 VSS.n5710 0.04025
R14876 VSS.n5712 VSS.n5711 0.04025
R14877 VSS.n5712 VSS.n2661 0.04025
R14878 VSS.n5716 VSS.n2661 0.04025
R14879 VSS.n5717 VSS.n5716 0.04025
R14880 VSS.n5718 VSS.n5717 0.04025
R14881 VSS.n5718 VSS.n2659 0.04025
R14882 VSS.n5722 VSS.n2659 0.04025
R14883 VSS.n5723 VSS.n5722 0.04025
R14884 VSS.n5724 VSS.n5723 0.04025
R14885 VSS.n5724 VSS.n2657 0.04025
R14886 VSS.n5728 VSS.n2657 0.04025
R14887 VSS.n5729 VSS.n5728 0.04025
R14888 VSS.n5730 VSS.n5729 0.04025
R14889 VSS.n5730 VSS.n2655 0.04025
R14890 VSS.n5734 VSS.n2655 0.04025
R14891 VSS.n5735 VSS.n5734 0.04025
R14892 VSS.n5736 VSS.n5735 0.04025
R14893 VSS.n5736 VSS.n2653 0.04025
R14894 VSS.n5740 VSS.n2653 0.04025
R14895 VSS.n5741 VSS.n5740 0.04025
R14896 VSS.n5742 VSS.n5741 0.04025
R14897 VSS.n5742 VSS.n2651 0.04025
R14898 VSS.n5746 VSS.n2651 0.04025
R14899 VSS.n5747 VSS.n5746 0.04025
R14900 VSS.n5748 VSS.n5747 0.04025
R14901 VSS.n5748 VSS.n2649 0.04025
R14902 VSS.n5752 VSS.n2649 0.04025
R14903 VSS.n5753 VSS.n5752 0.04025
R14904 VSS.n5754 VSS.n5753 0.04025
R14905 VSS.n5754 VSS.n2647 0.04025
R14906 VSS.n5758 VSS.n2647 0.04025
R14907 VSS.n5759 VSS.n5758 0.04025
R14908 VSS.n5760 VSS.n5759 0.04025
R14909 VSS.n5760 VSS.n2645 0.04025
R14910 VSS.n5764 VSS.n2645 0.04025
R14911 VSS.n5765 VSS.n5764 0.04025
R14912 VSS.n5766 VSS.n5765 0.04025
R14913 VSS.n5766 VSS.n2643 0.04025
R14914 VSS.n5770 VSS.n2643 0.04025
R14915 VSS.n5771 VSS.n5770 0.04025
R14916 VSS.n5772 VSS.n5771 0.04025
R14917 VSS.n5772 VSS.n2641 0.04025
R14918 VSS.n5776 VSS.n2641 0.04025
R14919 VSS.n5777 VSS.n5776 0.04025
R14920 VSS.n5778 VSS.n5777 0.04025
R14921 VSS.n5778 VSS.n2639 0.04025
R14922 VSS.n5782 VSS.n2639 0.04025
R14923 VSS.n5783 VSS.n5782 0.04025
R14924 VSS.n5784 VSS.n5783 0.04025
R14925 VSS.n5784 VSS.n2637 0.04025
R14926 VSS.n5788 VSS.n2637 0.04025
R14927 VSS.n5789 VSS.n5788 0.04025
R14928 VSS.n5790 VSS.n5789 0.04025
R14929 VSS.n5790 VSS.n2635 0.04025
R14930 VSS.n5794 VSS.n2635 0.04025
R14931 VSS.n5795 VSS.n5794 0.04025
R14932 VSS.n5796 VSS.n5795 0.04025
R14933 VSS.n5796 VSS.n2633 0.04025
R14934 VSS.n5800 VSS.n2633 0.04025
R14935 VSS.n5801 VSS.n5800 0.04025
R14936 VSS.n5802 VSS.n5801 0.04025
R14937 VSS.n5802 VSS.n2631 0.04025
R14938 VSS.n5806 VSS.n2631 0.04025
R14939 VSS.n5807 VSS.n5806 0.04025
R14940 VSS.n5808 VSS.n5807 0.04025
R14941 VSS.n5808 VSS.n2629 0.04025
R14942 VSS.n5812 VSS.n2629 0.04025
R14943 VSS.n5813 VSS.n5812 0.04025
R14944 VSS.n5814 VSS.n5813 0.04025
R14945 VSS.n5814 VSS.n2627 0.04025
R14946 VSS.n5818 VSS.n2627 0.04025
R14947 VSS.n5819 VSS.n5818 0.04025
R14948 VSS.n5820 VSS.n5819 0.04025
R14949 VSS.n5820 VSS.n2625 0.04025
R14950 VSS.n5824 VSS.n2625 0.04025
R14951 VSS.n5825 VSS.n5824 0.04025
R14952 VSS.n5826 VSS.n5825 0.04025
R14953 VSS.n5826 VSS.n2623 0.04025
R14954 VSS.n5830 VSS.n2623 0.04025
R14955 VSS.n5831 VSS.n5830 0.04025
R14956 VSS.n5832 VSS.n5831 0.04025
R14957 VSS.n5832 VSS.n2621 0.04025
R14958 VSS.n5836 VSS.n2621 0.04025
R14959 VSS.n5837 VSS.n5836 0.04025
R14960 VSS.n5838 VSS.n5837 0.04025
R14961 VSS.n5838 VSS.n2619 0.04025
R14962 VSS.n5842 VSS.n2619 0.04025
R14963 VSS.n5843 VSS.n5842 0.04025
R14964 VSS.n5844 VSS.n5843 0.04025
R14965 VSS.n5844 VSS.n2617 0.04025
R14966 VSS.n5848 VSS.n2617 0.04025
R14967 VSS.n5849 VSS.n5848 0.04025
R14968 VSS.n5850 VSS.n5849 0.04025
R14969 VSS.n5850 VSS.n2615 0.04025
R14970 VSS.n5854 VSS.n2615 0.04025
R14971 VSS.n5855 VSS.n5854 0.04025
R14972 VSS.n5856 VSS.n5855 0.04025
R14973 VSS.n5856 VSS.n2613 0.04025
R14974 VSS.n5860 VSS.n2613 0.04025
R14975 VSS.n5861 VSS.n5860 0.04025
R14976 VSS.n5862 VSS.n5861 0.04025
R14977 VSS.n5862 VSS.n2611 0.04025
R14978 VSS.n5866 VSS.n2611 0.04025
R14979 VSS.n5867 VSS.n5866 0.04025
R14980 VSS.n5868 VSS.n5867 0.04025
R14981 VSS.n5868 VSS.n2609 0.04025
R14982 VSS.n5872 VSS.n2609 0.04025
R14983 VSS.n5873 VSS.n5872 0.04025
R14984 VSS.n5874 VSS.n5873 0.04025
R14985 VSS.n5874 VSS.n2607 0.04025
R14986 VSS.n5878 VSS.n2607 0.04025
R14987 VSS.n5879 VSS.n5878 0.04025
R14988 VSS.n5880 VSS.n5879 0.04025
R14989 VSS.n5880 VSS.n2605 0.04025
R14990 VSS.n5884 VSS.n2605 0.04025
R14991 VSS.n5885 VSS.n5884 0.04025
R14992 VSS.n5886 VSS.n5885 0.04025
R14993 VSS.n5886 VSS.n2603 0.04025
R14994 VSS.n5890 VSS.n2603 0.04025
R14995 VSS.n5891 VSS.n5890 0.04025
R14996 VSS.n5892 VSS.n5891 0.04025
R14997 VSS.n5892 VSS.n2601 0.04025
R14998 VSS.n5896 VSS.n2601 0.04025
R14999 VSS.n5897 VSS.n5896 0.04025
R15000 VSS.n5898 VSS.n5897 0.04025
R15001 VSS.n5898 VSS.n2599 0.04025
R15002 VSS.n5902 VSS.n2599 0.04025
R15003 VSS.n5903 VSS.n5902 0.04025
R15004 VSS.n5904 VSS.n5903 0.04025
R15005 VSS.n5904 VSS.n2597 0.04025
R15006 VSS.n5908 VSS.n2597 0.04025
R15007 VSS.n5909 VSS.n5908 0.04025
R15008 VSS.n5910 VSS.n5909 0.04025
R15009 VSS.n5910 VSS.n2595 0.04025
R15010 VSS.n5914 VSS.n2595 0.04025
R15011 VSS.n5915 VSS.n5914 0.04025
R15012 VSS.n5916 VSS.n5915 0.04025
R15013 VSS.n5916 VSS.n2593 0.04025
R15014 VSS.n5920 VSS.n2593 0.04025
R15015 VSS.n5921 VSS.n5920 0.04025
R15016 VSS.n5922 VSS.n5921 0.04025
R15017 VSS.n5922 VSS.n2591 0.04025
R15018 VSS.n5926 VSS.n2591 0.04025
R15019 VSS.n5927 VSS.n5926 0.04025
R15020 VSS.n5928 VSS.n5927 0.04025
R15021 VSS.n5928 VSS.n2589 0.04025
R15022 VSS.n5932 VSS.n2589 0.04025
R15023 VSS.n5933 VSS.n5932 0.04025
R15024 VSS.n5934 VSS.n5933 0.04025
R15025 VSS.n5934 VSS.n2587 0.04025
R15026 VSS.n5938 VSS.n2587 0.04025
R15027 VSS.n5939 VSS.n5938 0.04025
R15028 VSS.n5940 VSS.n5939 0.04025
R15029 VSS.n5940 VSS.n2585 0.04025
R15030 VSS.n5944 VSS.n2585 0.04025
R15031 VSS.n5945 VSS.n5944 0.04025
R15032 VSS.n5946 VSS.n5945 0.04025
R15033 VSS.n5946 VSS.n2583 0.04025
R15034 VSS.n5950 VSS.n2583 0.04025
R15035 VSS.n5951 VSS.n5950 0.04025
R15036 VSS.n5952 VSS.n5951 0.04025
R15037 VSS.n5952 VSS.n2581 0.04025
R15038 VSS.n5956 VSS.n2581 0.04025
R15039 VSS.n5957 VSS.n5956 0.04025
R15040 VSS.n5958 VSS.n5957 0.04025
R15041 VSS.n5958 VSS.n2579 0.04025
R15042 VSS.n5962 VSS.n2579 0.04025
R15043 VSS.n5963 VSS.n5962 0.04025
R15044 VSS.n5964 VSS.n5963 0.04025
R15045 VSS.n5964 VSS.n2577 0.04025
R15046 VSS.n5968 VSS.n2577 0.04025
R15047 VSS.n5969 VSS.n5968 0.04025
R15048 VSS.n5970 VSS.n5969 0.04025
R15049 VSS.n5970 VSS.n2575 0.04025
R15050 VSS.n5974 VSS.n2575 0.04025
R15051 VSS.n5975 VSS.n5974 0.04025
R15052 VSS.n5976 VSS.n5975 0.04025
R15053 VSS.n5976 VSS.n2573 0.04025
R15054 VSS.n5980 VSS.n2573 0.04025
R15055 VSS.n5981 VSS.n5980 0.04025
R15056 VSS.n5982 VSS.n5981 0.04025
R15057 VSS.n5982 VSS.n2571 0.04025
R15058 VSS.n5986 VSS.n2571 0.04025
R15059 VSS.n5987 VSS.n5986 0.04025
R15060 VSS.n5988 VSS.n5987 0.04025
R15061 VSS.n5988 VSS.n2569 0.04025
R15062 VSS.n5992 VSS.n2569 0.04025
R15063 VSS.n5993 VSS.n5992 0.04025
R15064 VSS.n5994 VSS.n5993 0.04025
R15065 VSS.n5994 VSS.n2567 0.04025
R15066 VSS.n5998 VSS.n2567 0.04025
R15067 VSS.n5999 VSS.n5998 0.04025
R15068 VSS.n6000 VSS.n5999 0.04025
R15069 VSS.n6000 VSS.n2565 0.04025
R15070 VSS.n6004 VSS.n2565 0.04025
R15071 VSS.n6005 VSS.n6004 0.04025
R15072 VSS.n6006 VSS.n6005 0.04025
R15073 VSS.n6006 VSS.n2563 0.04025
R15074 VSS.n6010 VSS.n2563 0.04025
R15075 VSS.n6011 VSS.n6010 0.04025
R15076 VSS.n6012 VSS.n6011 0.04025
R15077 VSS.n6012 VSS.n2561 0.04025
R15078 VSS.n6016 VSS.n2561 0.04025
R15079 VSS.n6017 VSS.n6016 0.04025
R15080 VSS.n6018 VSS.n6017 0.04025
R15081 VSS.n6018 VSS.n2559 0.04025
R15082 VSS.n6022 VSS.n2559 0.04025
R15083 VSS.n6023 VSS.n6022 0.04025
R15084 VSS.n6024 VSS.n6023 0.04025
R15085 VSS.n6024 VSS.n2557 0.04025
R15086 VSS.n6028 VSS.n2557 0.04025
R15087 VSS.n6029 VSS.n6028 0.04025
R15088 VSS.n6030 VSS.n6029 0.04025
R15089 VSS.n6030 VSS.n2555 0.04025
R15090 VSS.n6034 VSS.n2555 0.04025
R15091 VSS.n6035 VSS.n6034 0.04025
R15092 VSS.n6036 VSS.n6035 0.04025
R15093 VSS.n6036 VSS.n2553 0.04025
R15094 VSS.n6040 VSS.n2553 0.04025
R15095 VSS.n6041 VSS.n6040 0.04025
R15096 VSS.n6042 VSS.n6041 0.04025
R15097 VSS.n6042 VSS.n2551 0.04025
R15098 VSS.n6046 VSS.n2551 0.04025
R15099 VSS.n6047 VSS.n6046 0.04025
R15100 VSS.n6048 VSS.n6047 0.04025
R15101 VSS.n6048 VSS.n2549 0.04025
R15102 VSS.n6052 VSS.n2549 0.04025
R15103 VSS.n6053 VSS.n6052 0.04025
R15104 VSS.n6054 VSS.n6053 0.04025
R15105 VSS.n6054 VSS.n2547 0.04025
R15106 VSS.n6058 VSS.n2547 0.04025
R15107 VSS.n6059 VSS.n6058 0.04025
R15108 VSS.n6060 VSS.n6059 0.04025
R15109 VSS.n6060 VSS.n2545 0.04025
R15110 VSS.n6064 VSS.n2545 0.04025
R15111 VSS.n6065 VSS.n6064 0.04025
R15112 VSS.n6066 VSS.n6065 0.04025
R15113 VSS.n6066 VSS.n2543 0.04025
R15114 VSS.n6070 VSS.n2543 0.04025
R15115 VSS.n6071 VSS.n6070 0.04025
R15116 VSS.n6072 VSS.n6071 0.04025
R15117 VSS.n6072 VSS.n2541 0.04025
R15118 VSS.n6076 VSS.n2541 0.04025
R15119 VSS.n6077 VSS.n6076 0.04025
R15120 VSS.n6078 VSS.n6077 0.04025
R15121 VSS.n6078 VSS.n2539 0.04025
R15122 VSS.n6082 VSS.n2539 0.04025
R15123 VSS.n6083 VSS.n6082 0.04025
R15124 VSS.n6084 VSS.n6083 0.04025
R15125 VSS.n6084 VSS.n2537 0.04025
R15126 VSS.n6088 VSS.n2537 0.04025
R15127 VSS.n6089 VSS.n6088 0.04025
R15128 VSS.n6090 VSS.n6089 0.04025
R15129 VSS.n6090 VSS.n2535 0.04025
R15130 VSS.n6094 VSS.n2535 0.04025
R15131 VSS.n6095 VSS.n6094 0.04025
R15132 VSS.n6096 VSS.n6095 0.04025
R15133 VSS.n6096 VSS.n2533 0.04025
R15134 VSS.n6100 VSS.n2533 0.04025
R15135 VSS.n6101 VSS.n6100 0.04025
R15136 VSS.n6102 VSS.n6101 0.04025
R15137 VSS.n6102 VSS.n2531 0.04025
R15138 VSS.n6106 VSS.n2531 0.04025
R15139 VSS.n6107 VSS.n6106 0.04025
R15140 VSS.n6108 VSS.n6107 0.04025
R15141 VSS.n6108 VSS.n2529 0.04025
R15142 VSS.n6112 VSS.n2529 0.04025
R15143 VSS.n6113 VSS.n6112 0.04025
R15144 VSS.n6114 VSS.n6113 0.04025
R15145 VSS.n6114 VSS.n2527 0.04025
R15146 VSS.n6118 VSS.n2527 0.04025
R15147 VSS.n6119 VSS.n6118 0.04025
R15148 VSS.n6120 VSS.n6119 0.04025
R15149 VSS.n6120 VSS.n2525 0.04025
R15150 VSS.n6124 VSS.n2525 0.04025
R15151 VSS.n6125 VSS.n6124 0.04025
R15152 VSS.n6126 VSS.n6125 0.04025
R15153 VSS.n6126 VSS.n2523 0.04025
R15154 VSS.n6130 VSS.n2523 0.04025
R15155 VSS.n6131 VSS.n6130 0.04025
R15156 VSS.n6132 VSS.n6131 0.04025
R15157 VSS.n6132 VSS.n2521 0.04025
R15158 VSS.n6136 VSS.n2521 0.04025
R15159 VSS.n6137 VSS.n6136 0.04025
R15160 VSS.n6138 VSS.n6137 0.04025
R15161 VSS.n6138 VSS.n2519 0.04025
R15162 VSS.n6142 VSS.n2519 0.04025
R15163 VSS.n6143 VSS.n6142 0.04025
R15164 VSS.n6144 VSS.n6143 0.04025
R15165 VSS.n6144 VSS.n2517 0.04025
R15166 VSS.n6148 VSS.n2517 0.04025
R15167 VSS.n6149 VSS.n6148 0.04025
R15168 VSS.n6150 VSS.n6149 0.04025
R15169 VSS.n6150 VSS.n2515 0.04025
R15170 VSS.n6154 VSS.n2515 0.04025
R15171 VSS.n6155 VSS.n6154 0.04025
R15172 VSS.n6156 VSS.n6155 0.04025
R15173 VSS.n6156 VSS.n2513 0.04025
R15174 VSS.n6160 VSS.n2513 0.04025
R15175 VSS.n6161 VSS.n6160 0.04025
R15176 VSS.n6162 VSS.n6161 0.04025
R15177 VSS.n6162 VSS.n2511 0.04025
R15178 VSS.n6166 VSS.n2511 0.04025
R15179 VSS.n6167 VSS.n6166 0.04025
R15180 VSS.n6168 VSS.n6167 0.04025
R15181 VSS.n6168 VSS.n2509 0.04025
R15182 VSS.n6172 VSS.n2509 0.04025
R15183 VSS.n6173 VSS.n6172 0.04025
R15184 VSS.n6174 VSS.n6173 0.04025
R15185 VSS.n6174 VSS.n2507 0.04025
R15186 VSS.n6178 VSS.n2507 0.04025
R15187 VSS.n6179 VSS.n6178 0.04025
R15188 VSS.n6180 VSS.n6179 0.04025
R15189 VSS.n6180 VSS.n2505 0.04025
R15190 VSS.n6184 VSS.n2505 0.04025
R15191 VSS.n6185 VSS.n6184 0.04025
R15192 VSS.n6186 VSS.n6185 0.04025
R15193 VSS.n6186 VSS.n2503 0.04025
R15194 VSS.n6190 VSS.n2503 0.04025
R15195 VSS.n6191 VSS.n6190 0.04025
R15196 VSS.n6192 VSS.n6191 0.04025
R15197 VSS.n6192 VSS.n2501 0.04025
R15198 VSS.n6196 VSS.n2501 0.04025
R15199 VSS.n6197 VSS.n6196 0.04025
R15200 VSS.n6198 VSS.n6197 0.04025
R15201 VSS.n6198 VSS.n2499 0.04025
R15202 VSS.n6202 VSS.n2499 0.04025
R15203 VSS.n6203 VSS.n6202 0.04025
R15204 VSS.n6204 VSS.n6203 0.04025
R15205 VSS.n6204 VSS.n2497 0.04025
R15206 VSS.n6208 VSS.n2497 0.04025
R15207 VSS.n6209 VSS.n6208 0.04025
R15208 VSS.n6210 VSS.n6209 0.04025
R15209 VSS.n6210 VSS.n2495 0.04025
R15210 VSS.n6214 VSS.n2495 0.04025
R15211 VSS.n6215 VSS.n6214 0.04025
R15212 VSS.n6216 VSS.n6215 0.04025
R15213 VSS.n6216 VSS.n2493 0.04025
R15214 VSS.n6220 VSS.n2493 0.04025
R15215 VSS.n6221 VSS.n6220 0.04025
R15216 VSS.n6222 VSS.n6221 0.04025
R15217 VSS.n6222 VSS.n2491 0.04025
R15218 VSS.n6226 VSS.n2491 0.04025
R15219 VSS.n6227 VSS.n6226 0.04025
R15220 VSS.n6228 VSS.n6227 0.04025
R15221 VSS.n6228 VSS.n2489 0.04025
R15222 VSS.n6232 VSS.n2489 0.04025
R15223 VSS.n6233 VSS.n6232 0.04025
R15224 VSS.n6234 VSS.n6233 0.04025
R15225 VSS.n6234 VSS.n2487 0.04025
R15226 VSS.n6238 VSS.n2487 0.04025
R15227 VSS.n6239 VSS.n6238 0.04025
R15228 VSS.n6240 VSS.n6239 0.04025
R15229 VSS.n6240 VSS.n2485 0.04025
R15230 VSS.n6244 VSS.n2485 0.04025
R15231 VSS.n6245 VSS.n6244 0.04025
R15232 VSS.n6246 VSS.n6245 0.04025
R15233 VSS.n6246 VSS.n2483 0.04025
R15234 VSS.n6250 VSS.n2483 0.04025
R15235 VSS.n6251 VSS.n6250 0.04025
R15236 VSS.n6252 VSS.n6251 0.04025
R15237 VSS.n6252 VSS.n2481 0.04025
R15238 VSS.n6256 VSS.n2481 0.04025
R15239 VSS.n6257 VSS.n6256 0.04025
R15240 VSS.n6258 VSS.n6257 0.04025
R15241 VSS.n6258 VSS.n2479 0.04025
R15242 VSS.n6262 VSS.n2479 0.04025
R15243 VSS.n6263 VSS.n6262 0.04025
R15244 VSS.n6264 VSS.n6263 0.04025
R15245 VSS.n6264 VSS.n2477 0.04025
R15246 VSS.n6268 VSS.n2477 0.04025
R15247 VSS.n6269 VSS.n6268 0.04025
R15248 VSS.n6270 VSS.n6269 0.04025
R15249 VSS.n6270 VSS.n2475 0.04025
R15250 VSS.n6274 VSS.n2475 0.04025
R15251 VSS.n6275 VSS.n6274 0.04025
R15252 VSS.n6276 VSS.n6275 0.04025
R15253 VSS.n6276 VSS.n2473 0.04025
R15254 VSS.n6280 VSS.n2473 0.04025
R15255 VSS.n6281 VSS.n6280 0.04025
R15256 VSS.n6282 VSS.n6281 0.04025
R15257 VSS.n6282 VSS.n2471 0.04025
R15258 VSS.n6286 VSS.n2471 0.04025
R15259 VSS.n6287 VSS.n6286 0.04025
R15260 VSS.n6288 VSS.n6287 0.04025
R15261 VSS.n6288 VSS.n2469 0.04025
R15262 VSS.n6292 VSS.n2469 0.04025
R15263 VSS.n6293 VSS.n6292 0.04025
R15264 VSS.n6294 VSS.n6293 0.04025
R15265 VSS.n6294 VSS.n2467 0.04025
R15266 VSS.n6298 VSS.n2467 0.04025
R15267 VSS.n6299 VSS.n6298 0.04025
R15268 VSS.n6300 VSS.n6299 0.04025
R15269 VSS.n6300 VSS.n2465 0.04025
R15270 VSS.n6304 VSS.n2465 0.04025
R15271 VSS.n6305 VSS.n6304 0.04025
R15272 VSS.n6306 VSS.n6305 0.04025
R15273 VSS.n6306 VSS.n2463 0.04025
R15274 VSS.n6310 VSS.n2463 0.04025
R15275 VSS.n6311 VSS.n6310 0.04025
R15276 VSS.n6312 VSS.n6311 0.04025
R15277 VSS.n6312 VSS.n2461 0.04025
R15278 VSS.n6316 VSS.n2461 0.04025
R15279 VSS.n6317 VSS.n6316 0.04025
R15280 VSS.n6318 VSS.n6317 0.04025
R15281 VSS.n6318 VSS.n2459 0.04025
R15282 VSS.n6322 VSS.n2459 0.04025
R15283 VSS.n6323 VSS.n6322 0.04025
R15284 VSS.n6324 VSS.n6323 0.04025
R15285 VSS.n6324 VSS.n2457 0.04025
R15286 VSS.n6328 VSS.n2457 0.04025
R15287 VSS.n6329 VSS.n6328 0.04025
R15288 VSS.n6330 VSS.n6329 0.04025
R15289 VSS.n6330 VSS.n2455 0.04025
R15290 VSS.n6334 VSS.n2455 0.04025
R15291 VSS.n6335 VSS.n6334 0.04025
R15292 VSS.n6336 VSS.n6335 0.04025
R15293 VSS.n6336 VSS.n2453 0.04025
R15294 VSS.n6340 VSS.n2453 0.04025
R15295 VSS.n6341 VSS.n6340 0.04025
R15296 VSS.n6342 VSS.n6341 0.04025
R15297 VSS.n6342 VSS.n2451 0.04025
R15298 VSS.n6346 VSS.n2451 0.04025
R15299 VSS.n6347 VSS.n6346 0.04025
R15300 VSS.n6348 VSS.n6347 0.04025
R15301 VSS.n6348 VSS.n2449 0.04025
R15302 VSS.n6352 VSS.n2449 0.04025
R15303 VSS.n6353 VSS.n6352 0.04025
R15304 VSS.n6354 VSS.n6353 0.04025
R15305 VSS.n6354 VSS.n2447 0.04025
R15306 VSS.n6358 VSS.n2447 0.04025
R15307 VSS.n6359 VSS.n6358 0.04025
R15308 VSS.n6360 VSS.n6359 0.04025
R15309 VSS.n6360 VSS.n2445 0.04025
R15310 VSS.n6364 VSS.n2445 0.04025
R15311 VSS.n6365 VSS.n6364 0.04025
R15312 VSS.n6366 VSS.n6365 0.04025
R15313 VSS.n6366 VSS.n2443 0.04025
R15314 VSS.n6370 VSS.n2443 0.04025
R15315 VSS.n6371 VSS.n6370 0.04025
R15316 VSS.n6372 VSS.n6371 0.04025
R15317 VSS.n6372 VSS.n2441 0.04025
R15318 VSS.n6376 VSS.n2441 0.04025
R15319 VSS.n6377 VSS.n6376 0.04025
R15320 VSS.n6378 VSS.n6377 0.04025
R15321 VSS.n6378 VSS.n2439 0.04025
R15322 VSS.n6382 VSS.n2439 0.04025
R15323 VSS.n6383 VSS.n6382 0.04025
R15324 VSS.n6384 VSS.n6383 0.04025
R15325 VSS.n6384 VSS.n2437 0.04025
R15326 VSS.n6388 VSS.n2437 0.04025
R15327 VSS.n6389 VSS.n6388 0.04025
R15328 VSS.n6390 VSS.n6389 0.04025
R15329 VSS.n6390 VSS.n2435 0.04025
R15330 VSS.n6394 VSS.n2435 0.04025
R15331 VSS.n6395 VSS.n6394 0.04025
R15332 VSS.n6396 VSS.n6395 0.04025
R15333 VSS.n6396 VSS.n2433 0.04025
R15334 VSS.n6400 VSS.n2433 0.04025
R15335 VSS.n6401 VSS.n6400 0.04025
R15336 VSS.n6402 VSS.n6401 0.04025
R15337 VSS.n6402 VSS.n2431 0.04025
R15338 VSS.n6406 VSS.n2431 0.04025
R15339 VSS.n6407 VSS.n6406 0.04025
R15340 VSS.n6408 VSS.n6407 0.04025
R15341 VSS.n6408 VSS.n2429 0.04025
R15342 VSS.n6412 VSS.n2429 0.04025
R15343 VSS.n6413 VSS.n6412 0.04025
R15344 VSS.n6414 VSS.n6413 0.04025
R15345 VSS.n6414 VSS.n2427 0.04025
R15346 VSS.n6418 VSS.n2427 0.04025
R15347 VSS.n6419 VSS.n6418 0.04025
R15348 VSS.n6420 VSS.n6419 0.04025
R15349 VSS.n6420 VSS.n2425 0.04025
R15350 VSS.n6424 VSS.n2425 0.04025
R15351 VSS.n6425 VSS.n6424 0.04025
R15352 VSS.n6426 VSS.n6425 0.04025
R15353 VSS.n6426 VSS.n2423 0.04025
R15354 VSS.n6430 VSS.n2423 0.04025
R15355 VSS.n6431 VSS.n6430 0.04025
R15356 VSS.n6432 VSS.n6431 0.04025
R15357 VSS.n6432 VSS.n2421 0.04025
R15358 VSS.n6436 VSS.n2421 0.04025
R15359 VSS.n6437 VSS.n6436 0.04025
R15360 VSS.n6438 VSS.n6437 0.04025
R15361 VSS.n6438 VSS.n2419 0.04025
R15362 VSS.n6442 VSS.n2419 0.04025
R15363 VSS.n6443 VSS.n6442 0.04025
R15364 VSS.n6444 VSS.n6443 0.04025
R15365 VSS.n6444 VSS.n2417 0.04025
R15366 VSS.n6448 VSS.n2417 0.04025
R15367 VSS.n6449 VSS.n6448 0.04025
R15368 VSS.n6450 VSS.n6449 0.04025
R15369 VSS.n6450 VSS.n2415 0.04025
R15370 VSS.n6454 VSS.n2415 0.04025
R15371 VSS.n6455 VSS.n6454 0.04025
R15372 VSS.n6456 VSS.n6455 0.04025
R15373 VSS.n6456 VSS.n2413 0.04025
R15374 VSS.n6460 VSS.n2413 0.04025
R15375 VSS.n6461 VSS.n6460 0.04025
R15376 VSS.n6462 VSS.n6461 0.04025
R15377 VSS.n6462 VSS.n2411 0.04025
R15378 VSS.n6466 VSS.n2411 0.04025
R15379 VSS.n6467 VSS.n6466 0.04025
R15380 VSS.n6468 VSS.n6467 0.04025
R15381 VSS.n6468 VSS.n2409 0.04025
R15382 VSS.n6472 VSS.n2409 0.04025
R15383 VSS.n6473 VSS.n6472 0.04025
R15384 VSS.n6474 VSS.n6473 0.04025
R15385 VSS.n6474 VSS.n2407 0.04025
R15386 VSS.n6478 VSS.n2407 0.04025
R15387 VSS.n6479 VSS.n6478 0.04025
R15388 VSS.n6480 VSS.n6479 0.04025
R15389 VSS.n6480 VSS.n2405 0.04025
R15390 VSS.n6484 VSS.n2405 0.04025
R15391 VSS.n6485 VSS.n6484 0.04025
R15392 VSS.n6486 VSS.n6485 0.04025
R15393 VSS.n6486 VSS.n2403 0.04025
R15394 VSS.n6490 VSS.n2403 0.04025
R15395 VSS.n6491 VSS.n6490 0.04025
R15396 VSS.n6492 VSS.n6491 0.04025
R15397 VSS.n6492 VSS.n2401 0.04025
R15398 VSS.n6496 VSS.n2401 0.04025
R15399 VSS.n6497 VSS.n6496 0.04025
R15400 VSS.n6498 VSS.n6497 0.04025
R15401 VSS.n6498 VSS.n2399 0.04025
R15402 VSS.n6502 VSS.n2399 0.04025
R15403 VSS.n6503 VSS.n6502 0.04025
R15404 VSS.n6504 VSS.n6503 0.04025
R15405 VSS.n6504 VSS.n2397 0.04025
R15406 VSS.n6508 VSS.n2397 0.04025
R15407 VSS.n6509 VSS.n6508 0.04025
R15408 VSS.n6510 VSS.n6509 0.04025
R15409 VSS.n6510 VSS.n2395 0.04025
R15410 VSS.n6514 VSS.n2395 0.04025
R15411 VSS.n6515 VSS.n6514 0.04025
R15412 VSS.n6516 VSS.n6515 0.04025
R15413 VSS.n6516 VSS.n2393 0.04025
R15414 VSS.n6520 VSS.n2393 0.04025
R15415 VSS.n6521 VSS.n6520 0.04025
R15416 VSS.n6522 VSS.n6521 0.04025
R15417 VSS.n6522 VSS.n2391 0.04025
R15418 VSS.n6526 VSS.n2391 0.04025
R15419 VSS.n6527 VSS.n6526 0.04025
R15420 VSS.n6528 VSS.n6527 0.04025
R15421 VSS.n6528 VSS.n2389 0.04025
R15422 VSS.n6532 VSS.n2389 0.04025
R15423 VSS.n6533 VSS.n6532 0.04025
R15424 VSS.n6534 VSS.n6533 0.04025
R15425 VSS.n6534 VSS.n2387 0.04025
R15426 VSS.n6538 VSS.n2387 0.04025
R15427 VSS.n6539 VSS.n6538 0.04025
R15428 VSS.n6540 VSS.n6539 0.04025
R15429 VSS.n6540 VSS.n2385 0.04025
R15430 VSS.n6544 VSS.n2385 0.04025
R15431 VSS.n6545 VSS.n6544 0.04025
R15432 VSS.n6546 VSS.n6545 0.04025
R15433 VSS.n6546 VSS.n2383 0.04025
R15434 VSS.n6550 VSS.n2383 0.04025
R15435 VSS.n6551 VSS.n6550 0.04025
R15436 VSS.n6552 VSS.n6551 0.04025
R15437 VSS.n6552 VSS.n2381 0.04025
R15438 VSS.n6556 VSS.n2381 0.04025
R15439 VSS.n6557 VSS.n6556 0.04025
R15440 VSS.n6558 VSS.n6557 0.04025
R15441 VSS.n6558 VSS.n2379 0.04025
R15442 VSS.n6562 VSS.n2379 0.04025
R15443 VSS.n6563 VSS.n6562 0.04025
R15444 VSS.n6564 VSS.n6563 0.04025
R15445 VSS.n6564 VSS.n2377 0.04025
R15446 VSS.n6568 VSS.n2377 0.04025
R15447 VSS.n6569 VSS.n6568 0.04025
R15448 VSS.n6570 VSS.n6569 0.04025
R15449 VSS.n6570 VSS.n2375 0.04025
R15450 VSS.n6574 VSS.n2375 0.04025
R15451 VSS.n6575 VSS.n6574 0.04025
R15452 VSS.n6576 VSS.n6575 0.04025
R15453 VSS.n6576 VSS.n2373 0.04025
R15454 VSS.n6580 VSS.n2373 0.04025
R15455 VSS.n6581 VSS.n6580 0.04025
R15456 VSS.n6582 VSS.n6581 0.04025
R15457 VSS.n6582 VSS.n2371 0.04025
R15458 VSS.n6586 VSS.n2371 0.04025
R15459 VSS.n6587 VSS.n6586 0.04025
R15460 VSS.n6588 VSS.n6587 0.04025
R15461 VSS.n6588 VSS.n2369 0.04025
R15462 VSS.n6592 VSS.n2369 0.04025
R15463 VSS.n6593 VSS.n6592 0.04025
R15464 VSS.n6594 VSS.n6593 0.04025
R15465 VSS.n6594 VSS.n2367 0.04025
R15466 VSS.n6598 VSS.n2367 0.04025
R15467 VSS.n6599 VSS.n6598 0.04025
R15468 VSS.n6600 VSS.n6599 0.04025
R15469 VSS.n6600 VSS.n2365 0.04025
R15470 VSS.n6604 VSS.n2365 0.04025
R15471 VSS.n6605 VSS.n6604 0.04025
R15472 VSS.n6606 VSS.n6605 0.04025
R15473 VSS.n6606 VSS.n2363 0.04025
R15474 VSS.n6610 VSS.n2363 0.04025
R15475 VSS.n6611 VSS.n6610 0.04025
R15476 VSS.n6612 VSS.n6611 0.04025
R15477 VSS.n6612 VSS.n2361 0.04025
R15478 VSS.n6616 VSS.n2361 0.04025
R15479 VSS.n6617 VSS.n6616 0.04025
R15480 VSS.n6618 VSS.n6617 0.04025
R15481 VSS.n6618 VSS.n2359 0.04025
R15482 VSS.n6622 VSS.n2359 0.04025
R15483 VSS.n6623 VSS.n6622 0.04025
R15484 VSS.n6624 VSS.n6623 0.04025
R15485 VSS.n6624 VSS.n2357 0.04025
R15486 VSS.n6628 VSS.n2357 0.04025
R15487 VSS.n6629 VSS.n6628 0.04025
R15488 VSS.n6630 VSS.n6629 0.04025
R15489 VSS.n6630 VSS.n2355 0.04025
R15490 VSS.n6634 VSS.n2355 0.04025
R15491 VSS.n6635 VSS.n6634 0.04025
R15492 VSS.n6636 VSS.n6635 0.04025
R15493 VSS.n6636 VSS.n2353 0.04025
R15494 VSS.n6640 VSS.n2353 0.04025
R15495 VSS.n6641 VSS.n6640 0.04025
R15496 VSS.n6642 VSS.n6641 0.04025
R15497 VSS.n6642 VSS.n2351 0.04025
R15498 VSS.n6646 VSS.n2351 0.04025
R15499 VSS.n6647 VSS.n6646 0.04025
R15500 VSS.n6648 VSS.n6647 0.04025
R15501 VSS.n6648 VSS.n2349 0.04025
R15502 VSS.n6652 VSS.n2349 0.04025
R15503 VSS.n6653 VSS.n6652 0.04025
R15504 VSS.n6654 VSS.n6653 0.04025
R15505 VSS.n6654 VSS.n2347 0.04025
R15506 VSS.n6658 VSS.n2347 0.04025
R15507 VSS.n6659 VSS.n6658 0.04025
R15508 VSS.n6660 VSS.n6659 0.04025
R15509 VSS.n6660 VSS.n2345 0.04025
R15510 VSS.n6664 VSS.n2345 0.04025
R15511 VSS.n6665 VSS.n6664 0.04025
R15512 VSS.n6666 VSS.n6665 0.04025
R15513 VSS.n6666 VSS.n2343 0.04025
R15514 VSS.n6670 VSS.n2343 0.04025
R15515 VSS.n6671 VSS.n6670 0.04025
R15516 VSS.n6672 VSS.n6671 0.04025
R15517 VSS.n6672 VSS.n2341 0.04025
R15518 VSS.n6676 VSS.n2341 0.04025
R15519 VSS.n6677 VSS.n6676 0.04025
R15520 VSS.n6678 VSS.n6677 0.04025
R15521 VSS.n6678 VSS.n2339 0.04025
R15522 VSS.n6682 VSS.n2339 0.04025
R15523 VSS.n6683 VSS.n6682 0.04025
R15524 VSS.n6684 VSS.n6683 0.04025
R15525 VSS.n6684 VSS.n2337 0.04025
R15526 VSS.n6688 VSS.n2337 0.04025
R15527 VSS.n6689 VSS.n6688 0.04025
R15528 VSS.n6690 VSS.n6689 0.04025
R15529 VSS.n6690 VSS.n2335 0.04025
R15530 VSS.n6694 VSS.n2335 0.04025
R15531 VSS.n6695 VSS.n6694 0.04025
R15532 VSS.n6696 VSS.n6695 0.04025
R15533 VSS.n6696 VSS.n2333 0.04025
R15534 VSS.n6700 VSS.n2333 0.04025
R15535 VSS.n6701 VSS.n6700 0.04025
R15536 VSS.n6702 VSS.n6701 0.04025
R15537 VSS.n6702 VSS.n2331 0.04025
R15538 VSS.n6706 VSS.n2331 0.04025
R15539 VSS.n6707 VSS.n6706 0.04025
R15540 VSS.n6708 VSS.n6707 0.04025
R15541 VSS.n6708 VSS.n2329 0.04025
R15542 VSS.n6712 VSS.n2329 0.04025
R15543 VSS.n6713 VSS.n6712 0.04025
R15544 VSS.n6714 VSS.n6713 0.04025
R15545 VSS.n6714 VSS.n2327 0.04025
R15546 VSS.n6718 VSS.n2327 0.04025
R15547 VSS.n6719 VSS.n6718 0.04025
R15548 VSS.n6720 VSS.n6719 0.04025
R15549 VSS.n6720 VSS.n2325 0.04025
R15550 VSS.n6724 VSS.n2325 0.04025
R15551 VSS.n6725 VSS.n6724 0.04025
R15552 VSS.n6726 VSS.n6725 0.04025
R15553 VSS.n6726 VSS.n2323 0.04025
R15554 VSS.n6730 VSS.n2323 0.04025
R15555 VSS.n6731 VSS.n6730 0.04025
R15556 VSS.n6732 VSS.n6731 0.04025
R15557 VSS.n6732 VSS.n2321 0.04025
R15558 VSS.n6736 VSS.n2321 0.04025
R15559 VSS.n6737 VSS.n6736 0.04025
R15560 VSS.n6738 VSS.n6737 0.04025
R15561 VSS.n6738 VSS.n2319 0.04025
R15562 VSS.n6742 VSS.n2319 0.04025
R15563 VSS.n6743 VSS.n6742 0.04025
R15564 VSS.n6744 VSS.n6743 0.04025
R15565 VSS.n6744 VSS.n2317 0.04025
R15566 VSS.n6748 VSS.n2317 0.04025
R15567 VSS.n6749 VSS.n6748 0.04025
R15568 VSS.n6750 VSS.n6749 0.04025
R15569 VSS.n6750 VSS.n2315 0.04025
R15570 VSS.n6754 VSS.n2315 0.04025
R15571 VSS.n6755 VSS.n6754 0.04025
R15572 VSS.n6756 VSS.n6755 0.04025
R15573 VSS.n6756 VSS.n2313 0.04025
R15574 VSS.n6760 VSS.n2313 0.04025
R15575 VSS.n6761 VSS.n6760 0.04025
R15576 VSS.n6762 VSS.n6761 0.04025
R15577 VSS.n6762 VSS.n2311 0.04025
R15578 VSS.n6766 VSS.n2311 0.04025
R15579 VSS.n6767 VSS.n6766 0.04025
R15580 VSS.n6768 VSS.n6767 0.04025
R15581 VSS.n6768 VSS.n2309 0.04025
R15582 VSS.n6772 VSS.n2309 0.04025
R15583 VSS.n6773 VSS.n6772 0.04025
R15584 VSS.n6774 VSS.n6773 0.04025
R15585 VSS.n6774 VSS.n2307 0.04025
R15586 VSS.n6778 VSS.n2307 0.04025
R15587 VSS.n6779 VSS.n6778 0.04025
R15588 VSS.n6780 VSS.n6779 0.04025
R15589 VSS.n6780 VSS.n2305 0.04025
R15590 VSS.n6784 VSS.n2305 0.04025
R15591 VSS.n6785 VSS.n6784 0.04025
R15592 VSS.n6786 VSS.n6785 0.04025
R15593 VSS.n6786 VSS.n2303 0.04025
R15594 VSS.n6790 VSS.n2303 0.04025
R15595 VSS.n6791 VSS.n6790 0.04025
R15596 VSS.n6792 VSS.n6791 0.04025
R15597 VSS.n6792 VSS.n2301 0.04025
R15598 VSS.n6796 VSS.n2301 0.04025
R15599 VSS.n6797 VSS.n6796 0.04025
R15600 VSS.n6798 VSS.n6797 0.04025
R15601 VSS.n6798 VSS.n2299 0.04025
R15602 VSS.n6802 VSS.n2299 0.04025
R15603 VSS.n6803 VSS.n6802 0.04025
R15604 VSS.n6804 VSS.n6803 0.04025
R15605 VSS.n6804 VSS.n2297 0.04025
R15606 VSS.n6808 VSS.n2297 0.04025
R15607 VSS.n6809 VSS.n6808 0.04025
R15608 VSS.n6810 VSS.n6809 0.04025
R15609 VSS.n6810 VSS.n2295 0.04025
R15610 VSS.n6814 VSS.n2295 0.04025
R15611 VSS.n6815 VSS.n6814 0.04025
R15612 VSS.n6816 VSS.n6815 0.04025
R15613 VSS.n6816 VSS.n2293 0.04025
R15614 VSS.n6820 VSS.n2293 0.04025
R15615 VSS.n6821 VSS.n6820 0.04025
R15616 VSS.n6822 VSS.n6821 0.04025
R15617 VSS.n6822 VSS.n2291 0.04025
R15618 VSS.n6826 VSS.n2291 0.04025
R15619 VSS.n6827 VSS.n6826 0.04025
R15620 VSS.n6828 VSS.n6827 0.04025
R15621 VSS.n6828 VSS.n2289 0.04025
R15622 VSS.n6832 VSS.n2289 0.04025
R15623 VSS.n6833 VSS.n6832 0.04025
R15624 VSS.n6834 VSS.n6833 0.04025
R15625 VSS.n6834 VSS.n2287 0.04025
R15626 VSS.n6838 VSS.n2287 0.04025
R15627 VSS.n6839 VSS.n6838 0.04025
R15628 VSS.n6840 VSS.n6839 0.04025
R15629 VSS.n6840 VSS.n2285 0.04025
R15630 VSS.n6844 VSS.n2285 0.04025
R15631 VSS.n6845 VSS.n6844 0.04025
R15632 VSS.n6846 VSS.n6845 0.04025
R15633 VSS.n6846 VSS.n2283 0.04025
R15634 VSS.n6850 VSS.n2283 0.04025
R15635 VSS.n6851 VSS.n6850 0.04025
R15636 VSS.n6852 VSS.n6851 0.04025
R15637 VSS.n6852 VSS.n2281 0.04025
R15638 VSS.n6856 VSS.n2281 0.04025
R15639 VSS.n6857 VSS.n6856 0.04025
R15640 VSS.n6858 VSS.n6857 0.04025
R15641 VSS.n6858 VSS.n2279 0.04025
R15642 VSS.n6862 VSS.n2279 0.04025
R15643 VSS.n6863 VSS.n6862 0.04025
R15644 VSS.n6864 VSS.n6863 0.04025
R15645 VSS.n6864 VSS.n2277 0.04025
R15646 VSS.n6868 VSS.n2277 0.04025
R15647 VSS.n6869 VSS.n6868 0.04025
R15648 VSS.n6870 VSS.n6869 0.04025
R15649 VSS.n6870 VSS.n2275 0.04025
R15650 VSS.n6874 VSS.n2275 0.04025
R15651 VSS.n6875 VSS.n6874 0.04025
R15652 VSS.n6876 VSS.n6875 0.04025
R15653 VSS.n6876 VSS.n2273 0.04025
R15654 VSS.n6880 VSS.n2273 0.04025
R15655 VSS.n6881 VSS.n6880 0.04025
R15656 VSS.n6882 VSS.n6881 0.04025
R15657 VSS.n6882 VSS.n2271 0.04025
R15658 VSS.n6886 VSS.n2271 0.04025
R15659 VSS.n6887 VSS.n6886 0.04025
R15660 VSS.n6888 VSS.n6887 0.04025
R15661 VSS.n6888 VSS.n2269 0.04025
R15662 VSS.n6892 VSS.n2269 0.04025
R15663 VSS.n6893 VSS.n6892 0.04025
R15664 VSS.n6894 VSS.n6893 0.04025
R15665 VSS.n6894 VSS.n2267 0.04025
R15666 VSS.n6898 VSS.n2267 0.04025
R15667 VSS.n6899 VSS.n6898 0.04025
R15668 VSS.n6900 VSS.n6899 0.04025
R15669 VSS.n6900 VSS.n2265 0.04025
R15670 VSS.n6904 VSS.n2265 0.04025
R15671 VSS.n6905 VSS.n6904 0.04025
R15672 VSS.n6906 VSS.n6905 0.04025
R15673 VSS.n8231 VSS.n8230 0.04025
R15674 VSS.n8230 VSS.n1823 0.04025
R15675 VSS.n8226 VSS.n1823 0.04025
R15676 VSS.n8226 VSS.n8225 0.04025
R15677 VSS.n8225 VSS.n8224 0.04025
R15678 VSS.n8224 VSS.n1825 0.04025
R15679 VSS.n8220 VSS.n1825 0.04025
R15680 VSS.n8220 VSS.n8219 0.04025
R15681 VSS.n8219 VSS.n8218 0.04025
R15682 VSS.n8218 VSS.n1827 0.04025
R15683 VSS.n8214 VSS.n1827 0.04025
R15684 VSS.n8214 VSS.n8213 0.04025
R15685 VSS.n8213 VSS.n8212 0.04025
R15686 VSS.n8212 VSS.n1829 0.04025
R15687 VSS.n8208 VSS.n1829 0.04025
R15688 VSS.n8208 VSS.n8207 0.04025
R15689 VSS.n8207 VSS.n8206 0.04025
R15690 VSS.n8206 VSS.n1831 0.04025
R15691 VSS.n8202 VSS.n1831 0.04025
R15692 VSS.n8202 VSS.n8201 0.04025
R15693 VSS.n8201 VSS.n8200 0.04025
R15694 VSS.n8200 VSS.n1833 0.04025
R15695 VSS.n8196 VSS.n1833 0.04025
R15696 VSS.n8196 VSS.n8195 0.04025
R15697 VSS.n8195 VSS.n8194 0.04025
R15698 VSS.n8194 VSS.n1835 0.04025
R15699 VSS.n8190 VSS.n1835 0.04025
R15700 VSS.n8190 VSS.n8189 0.04025
R15701 VSS.n8189 VSS.n8188 0.04025
R15702 VSS.n8188 VSS.n1837 0.04025
R15703 VSS.n8184 VSS.n1837 0.04025
R15704 VSS.n8184 VSS.n8183 0.04025
R15705 VSS.n8183 VSS.n8182 0.04025
R15706 VSS.n8182 VSS.n1839 0.04025
R15707 VSS.n8178 VSS.n1839 0.04025
R15708 VSS.n8178 VSS.n8177 0.04025
R15709 VSS.n8177 VSS.n8176 0.04025
R15710 VSS.n8176 VSS.n1841 0.04025
R15711 VSS.n8172 VSS.n1841 0.04025
R15712 VSS.n8172 VSS.n8171 0.04025
R15713 VSS.n8171 VSS.n8170 0.04025
R15714 VSS.n8170 VSS.n1843 0.04025
R15715 VSS.n8166 VSS.n1843 0.04025
R15716 VSS.n8166 VSS.n8165 0.04025
R15717 VSS.n8165 VSS.n8164 0.04025
R15718 VSS.n8164 VSS.n1845 0.04025
R15719 VSS.n8160 VSS.n1845 0.04025
R15720 VSS.n8160 VSS.n8159 0.04025
R15721 VSS.n8159 VSS.n8158 0.04025
R15722 VSS.n8158 VSS.n1847 0.04025
R15723 VSS.n8154 VSS.n1847 0.04025
R15724 VSS.n8154 VSS.n8153 0.04025
R15725 VSS.n8153 VSS.n8152 0.04025
R15726 VSS.n8152 VSS.n1849 0.04025
R15727 VSS.n8148 VSS.n1849 0.04025
R15728 VSS.n8148 VSS.n8147 0.04025
R15729 VSS.n8147 VSS.n8146 0.04025
R15730 VSS.n8146 VSS.n1851 0.04025
R15731 VSS.n8142 VSS.n1851 0.04025
R15732 VSS.n8142 VSS.n8141 0.04025
R15733 VSS.n8141 VSS.n8140 0.04025
R15734 VSS.n8140 VSS.n1853 0.04025
R15735 VSS.n8136 VSS.n1853 0.04025
R15736 VSS.n8136 VSS.n8135 0.04025
R15737 VSS.n8135 VSS.n8134 0.04025
R15738 VSS.n8134 VSS.n1855 0.04025
R15739 VSS.n8130 VSS.n1855 0.04025
R15740 VSS.n8130 VSS.n8129 0.04025
R15741 VSS.n8129 VSS.n8128 0.04025
R15742 VSS.n8128 VSS.n1857 0.04025
R15743 VSS.n8124 VSS.n1857 0.04025
R15744 VSS.n8124 VSS.n8123 0.04025
R15745 VSS.n8123 VSS.n8122 0.04025
R15746 VSS.n8122 VSS.n1859 0.04025
R15747 VSS.n8118 VSS.n1859 0.04025
R15748 VSS.n8118 VSS.n8117 0.04025
R15749 VSS.n8117 VSS.n8116 0.04025
R15750 VSS.n8116 VSS.n1861 0.04025
R15751 VSS.n8112 VSS.n1861 0.04025
R15752 VSS.n8112 VSS.n8111 0.04025
R15753 VSS.n8111 VSS.n8110 0.04025
R15754 VSS.n8110 VSS.n1863 0.04025
R15755 VSS.n8106 VSS.n1863 0.04025
R15756 VSS.n8106 VSS.n8105 0.04025
R15757 VSS.n8105 VSS.n8104 0.04025
R15758 VSS.n8104 VSS.n1865 0.04025
R15759 VSS.n8100 VSS.n1865 0.04025
R15760 VSS.n8100 VSS.n8099 0.04025
R15761 VSS.n8099 VSS.n8098 0.04025
R15762 VSS.n8098 VSS.n1867 0.04025
R15763 VSS.n8094 VSS.n1867 0.04025
R15764 VSS.n8094 VSS.n8093 0.04025
R15765 VSS.n8093 VSS.n8092 0.04025
R15766 VSS.n8092 VSS.n1869 0.04025
R15767 VSS.n8088 VSS.n1869 0.04025
R15768 VSS.n8088 VSS.n8087 0.04025
R15769 VSS.n8087 VSS.n8086 0.04025
R15770 VSS.n8086 VSS.n1871 0.04025
R15771 VSS.n8082 VSS.n1871 0.04025
R15772 VSS.n8082 VSS.n8081 0.04025
R15773 VSS.n8081 VSS.n8080 0.04025
R15774 VSS.n8080 VSS.n1873 0.04025
R15775 VSS.n8076 VSS.n1873 0.04025
R15776 VSS.n8076 VSS.n8075 0.04025
R15777 VSS.n8075 VSS.n8074 0.04025
R15778 VSS.n8074 VSS.n1875 0.04025
R15779 VSS.n8070 VSS.n1875 0.04025
R15780 VSS.n8070 VSS.n8069 0.04025
R15781 VSS.n8069 VSS.n8068 0.04025
R15782 VSS.n8068 VSS.n1877 0.04025
R15783 VSS.n8064 VSS.n1877 0.04025
R15784 VSS.n8064 VSS.n8063 0.04025
R15785 VSS.n8063 VSS.n8062 0.04025
R15786 VSS.n8062 VSS.n1879 0.04025
R15787 VSS.n8058 VSS.n1879 0.04025
R15788 VSS.n8058 VSS.n8057 0.04025
R15789 VSS.n8057 VSS.n8056 0.04025
R15790 VSS.n8056 VSS.n1881 0.04025
R15791 VSS.n8052 VSS.n1881 0.04025
R15792 VSS.n8052 VSS.n8051 0.04025
R15793 VSS.n8051 VSS.n8050 0.04025
R15794 VSS.n8050 VSS.n1883 0.04025
R15795 VSS.n8046 VSS.n1883 0.04025
R15796 VSS.n8046 VSS.n8045 0.04025
R15797 VSS.n8045 VSS.n8044 0.04025
R15798 VSS.n8044 VSS.n1885 0.04025
R15799 VSS.n8040 VSS.n1885 0.04025
R15800 VSS.n8040 VSS.n8039 0.04025
R15801 VSS.n8039 VSS.n8038 0.04025
R15802 VSS.n8038 VSS.n1887 0.04025
R15803 VSS.n8034 VSS.n1887 0.04025
R15804 VSS.n8034 VSS.n8033 0.04025
R15805 VSS.n8033 VSS.n8032 0.04025
R15806 VSS.n8032 VSS.n1889 0.04025
R15807 VSS.n8028 VSS.n1889 0.04025
R15808 VSS.n8028 VSS.n8027 0.04025
R15809 VSS.n8027 VSS.n8026 0.04025
R15810 VSS.n8026 VSS.n1891 0.04025
R15811 VSS.n8022 VSS.n1891 0.04025
R15812 VSS.n8022 VSS.n8021 0.04025
R15813 VSS.n8021 VSS.n8020 0.04025
R15814 VSS.n8020 VSS.n1893 0.04025
R15815 VSS.n8016 VSS.n1893 0.04025
R15816 VSS.n8016 VSS.n8015 0.04025
R15817 VSS.n8015 VSS.n8014 0.04025
R15818 VSS.n8014 VSS.n1895 0.04025
R15819 VSS.n8010 VSS.n1895 0.04025
R15820 VSS.n8010 VSS.n8009 0.04025
R15821 VSS.n8009 VSS.n8008 0.04025
R15822 VSS.n8008 VSS.n1897 0.04025
R15823 VSS.n8004 VSS.n1897 0.04025
R15824 VSS.n8004 VSS.n8003 0.04025
R15825 VSS.n8003 VSS.n8002 0.04025
R15826 VSS.n8002 VSS.n1899 0.04025
R15827 VSS.n7998 VSS.n1899 0.04025
R15828 VSS.n7998 VSS.n7997 0.04025
R15829 VSS.n7997 VSS.n7996 0.04025
R15830 VSS.n7996 VSS.n1901 0.04025
R15831 VSS.n7992 VSS.n1901 0.04025
R15832 VSS.n7992 VSS.n7991 0.04025
R15833 VSS.n7991 VSS.n7990 0.04025
R15834 VSS.n7990 VSS.n1903 0.04025
R15835 VSS.n7986 VSS.n1903 0.04025
R15836 VSS.n7986 VSS.n7985 0.04025
R15837 VSS.n7985 VSS.n7984 0.04025
R15838 VSS.n7984 VSS.n1905 0.04025
R15839 VSS.n7980 VSS.n1905 0.04025
R15840 VSS.n7980 VSS.n7979 0.04025
R15841 VSS.n7979 VSS.n7978 0.04025
R15842 VSS.n7978 VSS.n1907 0.04025
R15843 VSS.n7974 VSS.n1907 0.04025
R15844 VSS.n7974 VSS.n7973 0.04025
R15845 VSS.n7973 VSS.n7972 0.04025
R15846 VSS.n7972 VSS.n1909 0.04025
R15847 VSS.n7968 VSS.n1909 0.04025
R15848 VSS.n7968 VSS.n7967 0.04025
R15849 VSS.n7967 VSS.n7966 0.04025
R15850 VSS.n7966 VSS.n1911 0.04025
R15851 VSS.n7962 VSS.n1911 0.04025
R15852 VSS.n7962 VSS.n7961 0.04025
R15853 VSS.n7961 VSS.n7960 0.04025
R15854 VSS.n7960 VSS.n1913 0.04025
R15855 VSS.n7956 VSS.n1913 0.04025
R15856 VSS.n7956 VSS.n7955 0.04025
R15857 VSS.n7955 VSS.n7954 0.04025
R15858 VSS.n7954 VSS.n1915 0.04025
R15859 VSS.n7950 VSS.n1915 0.04025
R15860 VSS.n7950 VSS.n7949 0.04025
R15861 VSS.n7949 VSS.n7948 0.04025
R15862 VSS.n7948 VSS.n1917 0.04025
R15863 VSS.n7944 VSS.n1917 0.04025
R15864 VSS.n7944 VSS.n7943 0.04025
R15865 VSS.n7943 VSS.n7942 0.04025
R15866 VSS.n7942 VSS.n1919 0.04025
R15867 VSS.n7938 VSS.n1919 0.04025
R15868 VSS.n7938 VSS.n7937 0.04025
R15869 VSS.n7937 VSS.n7936 0.04025
R15870 VSS.n7936 VSS.n1921 0.04025
R15871 VSS.n7932 VSS.n1921 0.04025
R15872 VSS.n7932 VSS.n7931 0.04025
R15873 VSS.n7931 VSS.n7930 0.04025
R15874 VSS.n7930 VSS.n1923 0.04025
R15875 VSS.n7926 VSS.n1923 0.04025
R15876 VSS.n7926 VSS.n7925 0.04025
R15877 VSS.n7925 VSS.n7924 0.04025
R15878 VSS.n7924 VSS.n1925 0.04025
R15879 VSS.n7920 VSS.n1925 0.04025
R15880 VSS.n7920 VSS.n7919 0.04025
R15881 VSS.n7919 VSS.n7918 0.04025
R15882 VSS.n7918 VSS.n1927 0.04025
R15883 VSS.n7914 VSS.n1927 0.04025
R15884 VSS.n7914 VSS.n7913 0.04025
R15885 VSS.n7913 VSS.n7912 0.04025
R15886 VSS.n7912 VSS.n1929 0.04025
R15887 VSS.n7908 VSS.n1929 0.04025
R15888 VSS.n7908 VSS.n7907 0.04025
R15889 VSS.n7907 VSS.n7906 0.04025
R15890 VSS.n7906 VSS.n1931 0.04025
R15891 VSS.n7902 VSS.n1931 0.04025
R15892 VSS.n7902 VSS.n7901 0.04025
R15893 VSS.n7901 VSS.n7900 0.04025
R15894 VSS.n7900 VSS.n1933 0.04025
R15895 VSS.n7896 VSS.n1933 0.04025
R15896 VSS.n7896 VSS.n7895 0.04025
R15897 VSS.n7895 VSS.n7894 0.04025
R15898 VSS.n7894 VSS.n1935 0.04025
R15899 VSS.n7890 VSS.n1935 0.04025
R15900 VSS.n7890 VSS.n7889 0.04025
R15901 VSS.n7889 VSS.n7888 0.04025
R15902 VSS.n7888 VSS.n1937 0.04025
R15903 VSS.n7884 VSS.n1937 0.04025
R15904 VSS.n7884 VSS.n7883 0.04025
R15905 VSS.n7883 VSS.n7882 0.04025
R15906 VSS.n7882 VSS.n1939 0.04025
R15907 VSS.n7878 VSS.n1939 0.04025
R15908 VSS.n7878 VSS.n7877 0.04025
R15909 VSS.n7877 VSS.n7876 0.04025
R15910 VSS.n7876 VSS.n1941 0.04025
R15911 VSS.n7872 VSS.n1941 0.04025
R15912 VSS.n7872 VSS.n7871 0.04025
R15913 VSS.n7871 VSS.n7870 0.04025
R15914 VSS.n7870 VSS.n1943 0.04025
R15915 VSS.n7866 VSS.n1943 0.04025
R15916 VSS.n7866 VSS.n7865 0.04025
R15917 VSS.n7865 VSS.n7864 0.04025
R15918 VSS.n7864 VSS.n1945 0.04025
R15919 VSS.n7860 VSS.n1945 0.04025
R15920 VSS.n7860 VSS.n7859 0.04025
R15921 VSS.n7859 VSS.n7858 0.04025
R15922 VSS.n7858 VSS.n1947 0.04025
R15923 VSS.n7854 VSS.n1947 0.04025
R15924 VSS.n7854 VSS.n7853 0.04025
R15925 VSS.n7853 VSS.n7852 0.04025
R15926 VSS.n7852 VSS.n1949 0.04025
R15927 VSS.n7848 VSS.n1949 0.04025
R15928 VSS.n7848 VSS.n7847 0.04025
R15929 VSS.n7847 VSS.n7846 0.04025
R15930 VSS.n7846 VSS.n1951 0.04025
R15931 VSS.n7842 VSS.n1951 0.04025
R15932 VSS.n7842 VSS.n7841 0.04025
R15933 VSS.n7841 VSS.n7840 0.04025
R15934 VSS.n7840 VSS.n1953 0.04025
R15935 VSS.n7836 VSS.n1953 0.04025
R15936 VSS.n7836 VSS.n7835 0.04025
R15937 VSS.n7835 VSS.n7834 0.04025
R15938 VSS.n7834 VSS.n1955 0.04025
R15939 VSS.n7830 VSS.n1955 0.04025
R15940 VSS.n7830 VSS.n7829 0.04025
R15941 VSS.n7829 VSS.n7828 0.04025
R15942 VSS.n7828 VSS.n1957 0.04025
R15943 VSS.n7824 VSS.n1957 0.04025
R15944 VSS.n7824 VSS.n7823 0.04025
R15945 VSS.n7823 VSS.n7822 0.04025
R15946 VSS.n7822 VSS.n1959 0.04025
R15947 VSS.n7818 VSS.n1959 0.04025
R15948 VSS.n7818 VSS.n7817 0.04025
R15949 VSS.n7817 VSS.n7816 0.04025
R15950 VSS.n7816 VSS.n1961 0.04025
R15951 VSS.n7812 VSS.n1961 0.04025
R15952 VSS.n7812 VSS.n7811 0.04025
R15953 VSS.n7811 VSS.n7810 0.04025
R15954 VSS.n7810 VSS.n1963 0.04025
R15955 VSS.n7806 VSS.n1963 0.04025
R15956 VSS.n7806 VSS.n7805 0.04025
R15957 VSS.n7805 VSS.n7804 0.04025
R15958 VSS.n7804 VSS.n1965 0.04025
R15959 VSS.n7800 VSS.n1965 0.04025
R15960 VSS.n7800 VSS.n7799 0.04025
R15961 VSS.n7799 VSS.n7798 0.04025
R15962 VSS.n7798 VSS.n1967 0.04025
R15963 VSS.n7794 VSS.n1967 0.04025
R15964 VSS.n7794 VSS.n7793 0.04025
R15965 VSS.n7793 VSS.n7792 0.04025
R15966 VSS.n7792 VSS.n1969 0.04025
R15967 VSS.n7788 VSS.n1969 0.04025
R15968 VSS.n7788 VSS.n7787 0.04025
R15969 VSS.n7787 VSS.n7786 0.04025
R15970 VSS.n7786 VSS.n1971 0.04025
R15971 VSS.n7782 VSS.n1971 0.04025
R15972 VSS.n7782 VSS.n7781 0.04025
R15973 VSS.n7781 VSS.n7780 0.04025
R15974 VSS.n7780 VSS.n1973 0.04025
R15975 VSS.n7776 VSS.n1973 0.04025
R15976 VSS.n7776 VSS.n7775 0.04025
R15977 VSS.n7775 VSS.n7774 0.04025
R15978 VSS.n7774 VSS.n1975 0.04025
R15979 VSS.n7770 VSS.n1975 0.04025
R15980 VSS.n7770 VSS.n7769 0.04025
R15981 VSS.n7769 VSS.n7768 0.04025
R15982 VSS.n7768 VSS.n1977 0.04025
R15983 VSS.n7764 VSS.n1977 0.04025
R15984 VSS.n7764 VSS.n7763 0.04025
R15985 VSS.n7763 VSS.n7762 0.04025
R15986 VSS.n7762 VSS.n1979 0.04025
R15987 VSS.n7758 VSS.n1979 0.04025
R15988 VSS.n7758 VSS.n7757 0.04025
R15989 VSS.n7757 VSS.n7756 0.04025
R15990 VSS.n7756 VSS.n1981 0.04025
R15991 VSS.n7752 VSS.n1981 0.04025
R15992 VSS.n7752 VSS.n7751 0.04025
R15993 VSS.n7751 VSS.n7750 0.04025
R15994 VSS.n7750 VSS.n1983 0.04025
R15995 VSS.n7746 VSS.n1983 0.04025
R15996 VSS.n7746 VSS.n7745 0.04025
R15997 VSS.n7745 VSS.n7744 0.04025
R15998 VSS.n7744 VSS.n1985 0.04025
R15999 VSS.n7740 VSS.n1985 0.04025
R16000 VSS.n7740 VSS.n7739 0.04025
R16001 VSS.n7739 VSS.n7738 0.04025
R16002 VSS.n7738 VSS.n1987 0.04025
R16003 VSS.n7734 VSS.n1987 0.04025
R16004 VSS.n7734 VSS.n7733 0.04025
R16005 VSS.n7733 VSS.n7732 0.04025
R16006 VSS.n7732 VSS.n1989 0.04025
R16007 VSS.n7728 VSS.n1989 0.04025
R16008 VSS.n7728 VSS.n7727 0.04025
R16009 VSS.n7727 VSS.n7726 0.04025
R16010 VSS.n7726 VSS.n1991 0.04025
R16011 VSS.n7722 VSS.n1991 0.04025
R16012 VSS.n7722 VSS.n7721 0.04025
R16013 VSS.n7721 VSS.n7720 0.04025
R16014 VSS.n7720 VSS.n1993 0.04025
R16015 VSS.n7716 VSS.n1993 0.04025
R16016 VSS.n7716 VSS.n7715 0.04025
R16017 VSS.n7715 VSS.n7714 0.04025
R16018 VSS.n7714 VSS.n1995 0.04025
R16019 VSS.n7710 VSS.n1995 0.04025
R16020 VSS.n7710 VSS.n7709 0.04025
R16021 VSS.n7709 VSS.n7708 0.04025
R16022 VSS.n7708 VSS.n1997 0.04025
R16023 VSS.n7704 VSS.n1997 0.04025
R16024 VSS.n7704 VSS.n7703 0.04025
R16025 VSS.n7703 VSS.n7702 0.04025
R16026 VSS.n7702 VSS.n1999 0.04025
R16027 VSS.n7698 VSS.n1999 0.04025
R16028 VSS.n7698 VSS.n7697 0.04025
R16029 VSS.n7697 VSS.n7696 0.04025
R16030 VSS.n7696 VSS.n2001 0.04025
R16031 VSS.n7692 VSS.n2001 0.04025
R16032 VSS.n7692 VSS.n7691 0.04025
R16033 VSS.n7691 VSS.n7690 0.04025
R16034 VSS.n7690 VSS.n2003 0.04025
R16035 VSS.n7686 VSS.n2003 0.04025
R16036 VSS.n7686 VSS.n7685 0.04025
R16037 VSS.n7685 VSS.n7684 0.04025
R16038 VSS.n7684 VSS.n2005 0.04025
R16039 VSS.n7680 VSS.n2005 0.04025
R16040 VSS.n7680 VSS.n7679 0.04025
R16041 VSS.n7679 VSS.n7678 0.04025
R16042 VSS.n7678 VSS.n2007 0.04025
R16043 VSS.n7674 VSS.n2007 0.04025
R16044 VSS.n7674 VSS.n7673 0.04025
R16045 VSS.n7673 VSS.n7672 0.04025
R16046 VSS.n7672 VSS.n2009 0.04025
R16047 VSS.n7668 VSS.n2009 0.04025
R16048 VSS.n7668 VSS.n7667 0.04025
R16049 VSS.n7667 VSS.n7666 0.04025
R16050 VSS.n7666 VSS.n2011 0.04025
R16051 VSS.n7662 VSS.n2011 0.04025
R16052 VSS.n7662 VSS.n7661 0.04025
R16053 VSS.n7661 VSS.n7660 0.04025
R16054 VSS.n7660 VSS.n2013 0.04025
R16055 VSS.n7656 VSS.n2013 0.04025
R16056 VSS.n7656 VSS.n7655 0.04025
R16057 VSS.n7655 VSS.n7654 0.04025
R16058 VSS.n7654 VSS.n2015 0.04025
R16059 VSS.n7650 VSS.n2015 0.04025
R16060 VSS.n7650 VSS.n7649 0.04025
R16061 VSS.n7649 VSS.n7648 0.04025
R16062 VSS.n7648 VSS.n2017 0.04025
R16063 VSS.n7644 VSS.n2017 0.04025
R16064 VSS.n7644 VSS.n7643 0.04025
R16065 VSS.n7643 VSS.n7642 0.04025
R16066 VSS.n7642 VSS.n2019 0.04025
R16067 VSS.n7638 VSS.n2019 0.04025
R16068 VSS.n7638 VSS.n7637 0.04025
R16069 VSS.n7637 VSS.n7636 0.04025
R16070 VSS.n7636 VSS.n2021 0.04025
R16071 VSS.n7632 VSS.n2021 0.04025
R16072 VSS.n7632 VSS.n7631 0.04025
R16073 VSS.n7631 VSS.n7630 0.04025
R16074 VSS.n7630 VSS.n2023 0.04025
R16075 VSS.n7626 VSS.n2023 0.04025
R16076 VSS.n7626 VSS.n7625 0.04025
R16077 VSS.n7625 VSS.n7624 0.04025
R16078 VSS.n7624 VSS.n2025 0.04025
R16079 VSS.n7620 VSS.n2025 0.04025
R16080 VSS.n7620 VSS.n7619 0.04025
R16081 VSS.n7619 VSS.n7618 0.04025
R16082 VSS.n7618 VSS.n2027 0.04025
R16083 VSS.n7614 VSS.n2027 0.04025
R16084 VSS.n7614 VSS.n7613 0.04025
R16085 VSS.n7613 VSS.n7612 0.04025
R16086 VSS.n7612 VSS.n2029 0.04025
R16087 VSS.n7608 VSS.n2029 0.04025
R16088 VSS.n7608 VSS.n7607 0.04025
R16089 VSS.n7607 VSS.n7606 0.04025
R16090 VSS.n7606 VSS.n2031 0.04025
R16091 VSS.n7602 VSS.n2031 0.04025
R16092 VSS.n7602 VSS.n7601 0.04025
R16093 VSS.n7601 VSS.n7600 0.04025
R16094 VSS.n7600 VSS.n2033 0.04025
R16095 VSS.n7596 VSS.n2033 0.04025
R16096 VSS.n7596 VSS.n7595 0.04025
R16097 VSS.n7595 VSS.n7594 0.04025
R16098 VSS.n7594 VSS.n2035 0.04025
R16099 VSS.n7590 VSS.n2035 0.04025
R16100 VSS.n7590 VSS.n7589 0.04025
R16101 VSS.n7589 VSS.n7588 0.04025
R16102 VSS.n7588 VSS.n2037 0.04025
R16103 VSS.n7584 VSS.n2037 0.04025
R16104 VSS.n7584 VSS.n7583 0.04025
R16105 VSS.n7583 VSS.n7582 0.04025
R16106 VSS.n7582 VSS.n2039 0.04025
R16107 VSS.n7578 VSS.n2039 0.04025
R16108 VSS.n7578 VSS.n7577 0.04025
R16109 VSS.n7577 VSS.n7576 0.04025
R16110 VSS.n7576 VSS.n2041 0.04025
R16111 VSS.n7572 VSS.n2041 0.04025
R16112 VSS.n7572 VSS.n7571 0.04025
R16113 VSS.n7571 VSS.n7570 0.04025
R16114 VSS.n7570 VSS.n2043 0.04025
R16115 VSS.n7566 VSS.n2043 0.04025
R16116 VSS.n7566 VSS.n7565 0.04025
R16117 VSS.n7565 VSS.n7564 0.04025
R16118 VSS.n7564 VSS.n2045 0.04025
R16119 VSS.n7560 VSS.n2045 0.04025
R16120 VSS.n7560 VSS.n7559 0.04025
R16121 VSS.n7559 VSS.n7558 0.04025
R16122 VSS.n7558 VSS.n2047 0.04025
R16123 VSS.n7554 VSS.n2047 0.04025
R16124 VSS.n7554 VSS.n7553 0.04025
R16125 VSS.n7553 VSS.n7552 0.04025
R16126 VSS.n7552 VSS.n2049 0.04025
R16127 VSS.n7548 VSS.n2049 0.04025
R16128 VSS.n7548 VSS.n7547 0.04025
R16129 VSS.n7547 VSS.n7546 0.04025
R16130 VSS.n7546 VSS.n2051 0.04025
R16131 VSS.n7542 VSS.n2051 0.04025
R16132 VSS.n7542 VSS.n7541 0.04025
R16133 VSS.n7541 VSS.n7540 0.04025
R16134 VSS.n7540 VSS.n2053 0.04025
R16135 VSS.n7536 VSS.n2053 0.04025
R16136 VSS.n7536 VSS.n7535 0.04025
R16137 VSS.n7535 VSS.n7534 0.04025
R16138 VSS.n7534 VSS.n2055 0.04025
R16139 VSS.n7530 VSS.n2055 0.04025
R16140 VSS.n7530 VSS.n7529 0.04025
R16141 VSS.n7529 VSS.n7528 0.04025
R16142 VSS.n7528 VSS.n2057 0.04025
R16143 VSS.n7524 VSS.n2057 0.04025
R16144 VSS.n7524 VSS.n7523 0.04025
R16145 VSS.n7523 VSS.n7522 0.04025
R16146 VSS.n7522 VSS.n2059 0.04025
R16147 VSS.n7518 VSS.n2059 0.04025
R16148 VSS.n7518 VSS.n7517 0.04025
R16149 VSS.n7517 VSS.n7516 0.04025
R16150 VSS.n7516 VSS.n2061 0.04025
R16151 VSS.n7512 VSS.n2061 0.04025
R16152 VSS.n7512 VSS.n7511 0.04025
R16153 VSS.n7511 VSS.n7510 0.04025
R16154 VSS.n7510 VSS.n2063 0.04025
R16155 VSS.n7506 VSS.n2063 0.04025
R16156 VSS.n7506 VSS.n7505 0.04025
R16157 VSS.n7505 VSS.n7504 0.04025
R16158 VSS.n7504 VSS.n2065 0.04025
R16159 VSS.n7500 VSS.n2065 0.04025
R16160 VSS.n7500 VSS.n7499 0.04025
R16161 VSS.n7499 VSS.n7498 0.04025
R16162 VSS.n7498 VSS.n2067 0.04025
R16163 VSS.n7494 VSS.n2067 0.04025
R16164 VSS.n7494 VSS.n7493 0.04025
R16165 VSS.n7493 VSS.n7492 0.04025
R16166 VSS.n7492 VSS.n2069 0.04025
R16167 VSS.n7488 VSS.n2069 0.04025
R16168 VSS.n7488 VSS.n7487 0.04025
R16169 VSS.n7487 VSS.n7486 0.04025
R16170 VSS.n7486 VSS.n2071 0.04025
R16171 VSS.n7482 VSS.n2071 0.04025
R16172 VSS.n7482 VSS.n7481 0.04025
R16173 VSS.n7481 VSS.n7480 0.04025
R16174 VSS.n7480 VSS.n2073 0.04025
R16175 VSS.n7476 VSS.n2073 0.04025
R16176 VSS.n7476 VSS.n7475 0.04025
R16177 VSS.n7475 VSS.n7474 0.04025
R16178 VSS.n7474 VSS.n2075 0.04025
R16179 VSS.n7470 VSS.n2075 0.04025
R16180 VSS.n7470 VSS.n7469 0.04025
R16181 VSS.n7469 VSS.n7468 0.04025
R16182 VSS.n7468 VSS.n2077 0.04025
R16183 VSS.n7464 VSS.n2077 0.04025
R16184 VSS.n7464 VSS.n7463 0.04025
R16185 VSS.n7463 VSS.n7462 0.04025
R16186 VSS.n7462 VSS.n2079 0.04025
R16187 VSS.n7458 VSS.n2079 0.04025
R16188 VSS.n7458 VSS.n7457 0.04025
R16189 VSS.n7457 VSS.n7456 0.04025
R16190 VSS.n7456 VSS.n2081 0.04025
R16191 VSS.n7452 VSS.n2081 0.04025
R16192 VSS.n7452 VSS.n7451 0.04025
R16193 VSS.n7451 VSS.n7450 0.04025
R16194 VSS.n7450 VSS.n2083 0.04025
R16195 VSS.n7446 VSS.n2083 0.04025
R16196 VSS.n7446 VSS.n7445 0.04025
R16197 VSS.n7445 VSS.n7444 0.04025
R16198 VSS.n7444 VSS.n2085 0.04025
R16199 VSS.n7440 VSS.n2085 0.04025
R16200 VSS.n7440 VSS.n7439 0.04025
R16201 VSS.n7439 VSS.n7438 0.04025
R16202 VSS.n7438 VSS.n2087 0.04025
R16203 VSS.n7434 VSS.n2087 0.04025
R16204 VSS.n7434 VSS.n7433 0.04025
R16205 VSS.n7433 VSS.n7432 0.04025
R16206 VSS.n7432 VSS.n2089 0.04025
R16207 VSS.n7428 VSS.n2089 0.04025
R16208 VSS.n7428 VSS.n7427 0.04025
R16209 VSS.n7427 VSS.n7426 0.04025
R16210 VSS.n7426 VSS.n2091 0.04025
R16211 VSS.n7422 VSS.n2091 0.04025
R16212 VSS.n7422 VSS.n7421 0.04025
R16213 VSS.n7421 VSS.n7420 0.04025
R16214 VSS.n7420 VSS.n2093 0.04025
R16215 VSS.n7416 VSS.n2093 0.04025
R16216 VSS.n7416 VSS.n7415 0.04025
R16217 VSS.n7415 VSS.n7414 0.04025
R16218 VSS.n7414 VSS.n2095 0.04025
R16219 VSS.n7410 VSS.n2095 0.04025
R16220 VSS.n7410 VSS.n7409 0.04025
R16221 VSS.n7409 VSS.n7408 0.04025
R16222 VSS.n7408 VSS.n2097 0.04025
R16223 VSS.n7404 VSS.n2097 0.04025
R16224 VSS.n7404 VSS.n7403 0.04025
R16225 VSS.n7403 VSS.n7402 0.04025
R16226 VSS.n7402 VSS.n2099 0.04025
R16227 VSS.n7398 VSS.n2099 0.04025
R16228 VSS.n7398 VSS.n7397 0.04025
R16229 VSS.n7397 VSS.n7396 0.04025
R16230 VSS.n7396 VSS.n2101 0.04025
R16231 VSS.n7392 VSS.n2101 0.04025
R16232 VSS.n7392 VSS.n7391 0.04025
R16233 VSS.n7391 VSS.n7390 0.04025
R16234 VSS.n7390 VSS.n2103 0.04025
R16235 VSS.n7386 VSS.n2103 0.04025
R16236 VSS.n7386 VSS.n7385 0.04025
R16237 VSS.n7385 VSS.n7384 0.04025
R16238 VSS.n7384 VSS.n2105 0.04025
R16239 VSS.n7380 VSS.n2105 0.04025
R16240 VSS.n7380 VSS.n7379 0.04025
R16241 VSS.n7379 VSS.n7378 0.04025
R16242 VSS.n7378 VSS.n2107 0.04025
R16243 VSS.n7374 VSS.n2107 0.04025
R16244 VSS.n7374 VSS.n7373 0.04025
R16245 VSS.n7373 VSS.n7372 0.04025
R16246 VSS.n7372 VSS.n2109 0.04025
R16247 VSS.n7368 VSS.n2109 0.04025
R16248 VSS.n7368 VSS.n7367 0.04025
R16249 VSS.n7367 VSS.n7366 0.04025
R16250 VSS.n7366 VSS.n2111 0.04025
R16251 VSS.n7362 VSS.n2111 0.04025
R16252 VSS.n7362 VSS.n7361 0.04025
R16253 VSS.n7361 VSS.n7360 0.04025
R16254 VSS.n7360 VSS.n2113 0.04025
R16255 VSS.n7356 VSS.n2113 0.04025
R16256 VSS.n7356 VSS.n7355 0.04025
R16257 VSS.n7355 VSS.n7354 0.04025
R16258 VSS.n7354 VSS.n2115 0.04025
R16259 VSS.n7350 VSS.n2115 0.04025
R16260 VSS.n7350 VSS.n7349 0.04025
R16261 VSS.n7349 VSS.n7348 0.04025
R16262 VSS.n7348 VSS.n2117 0.04025
R16263 VSS.n7344 VSS.n2117 0.04025
R16264 VSS.n7344 VSS.n7343 0.04025
R16265 VSS.n7343 VSS.n7342 0.04025
R16266 VSS.n7342 VSS.n2119 0.04025
R16267 VSS.n7338 VSS.n2119 0.04025
R16268 VSS.n7338 VSS.n7337 0.04025
R16269 VSS.n7337 VSS.n7336 0.04025
R16270 VSS.n7336 VSS.n2121 0.04025
R16271 VSS.n7332 VSS.n2121 0.04025
R16272 VSS.n7332 VSS.n7331 0.04025
R16273 VSS.n7331 VSS.n7330 0.04025
R16274 VSS.n7330 VSS.n2123 0.04025
R16275 VSS.n7326 VSS.n2123 0.04025
R16276 VSS.n7326 VSS.n7325 0.04025
R16277 VSS.n7325 VSS.n7324 0.04025
R16278 VSS.n7324 VSS.n2125 0.04025
R16279 VSS.n7320 VSS.n2125 0.04025
R16280 VSS.n7320 VSS.n7319 0.04025
R16281 VSS.n7319 VSS.n7318 0.04025
R16282 VSS.n7318 VSS.n2127 0.04025
R16283 VSS.n7314 VSS.n2127 0.04025
R16284 VSS.n7314 VSS.n7313 0.04025
R16285 VSS.n7313 VSS.n7312 0.04025
R16286 VSS.n7312 VSS.n2129 0.04025
R16287 VSS.n7308 VSS.n2129 0.04025
R16288 VSS.n7308 VSS.n7307 0.04025
R16289 VSS.n7307 VSS.n7306 0.04025
R16290 VSS.n7306 VSS.n2131 0.04025
R16291 VSS.n7302 VSS.n2131 0.04025
R16292 VSS.n7302 VSS.n7301 0.04025
R16293 VSS.n7301 VSS.n7300 0.04025
R16294 VSS.n7300 VSS.n2133 0.04025
R16295 VSS.n7296 VSS.n2133 0.04025
R16296 VSS.n7296 VSS.n7295 0.04025
R16297 VSS.n7295 VSS.n7294 0.04025
R16298 VSS.n7294 VSS.n2135 0.04025
R16299 VSS.n7290 VSS.n2135 0.04025
R16300 VSS.n7290 VSS.n7289 0.04025
R16301 VSS.n7289 VSS.n7288 0.04025
R16302 VSS.n7288 VSS.n2137 0.04025
R16303 VSS.n7284 VSS.n2137 0.04025
R16304 VSS.n7284 VSS.n7283 0.04025
R16305 VSS.n7283 VSS.n7282 0.04025
R16306 VSS.n7282 VSS.n2139 0.04025
R16307 VSS.n7278 VSS.n2139 0.04025
R16308 VSS.n7278 VSS.n7277 0.04025
R16309 VSS.n7277 VSS.n7276 0.04025
R16310 VSS.n7276 VSS.n2141 0.04025
R16311 VSS.n7272 VSS.n2141 0.04025
R16312 VSS.n7272 VSS.n7271 0.04025
R16313 VSS.n7271 VSS.n7270 0.04025
R16314 VSS.n7270 VSS.n2143 0.04025
R16315 VSS.n7266 VSS.n2143 0.04025
R16316 VSS.n7266 VSS.n7265 0.04025
R16317 VSS.n7265 VSS.n7264 0.04025
R16318 VSS.n7264 VSS.n2145 0.04025
R16319 VSS.n7260 VSS.n2145 0.04025
R16320 VSS.n7260 VSS.n7259 0.04025
R16321 VSS.n7259 VSS.n7258 0.04025
R16322 VSS.n7258 VSS.n2147 0.04025
R16323 VSS.n7254 VSS.n2147 0.04025
R16324 VSS.n7254 VSS.n7253 0.04025
R16325 VSS.n7253 VSS.n7252 0.04025
R16326 VSS.n7252 VSS.n2149 0.04025
R16327 VSS.n7248 VSS.n2149 0.04025
R16328 VSS.n7248 VSS.n7247 0.04025
R16329 VSS.n7247 VSS.n7246 0.04025
R16330 VSS.n7246 VSS.n2151 0.04025
R16331 VSS.n7242 VSS.n2151 0.04025
R16332 VSS.n7242 VSS.n7241 0.04025
R16333 VSS.n7241 VSS.n7240 0.04025
R16334 VSS.n7240 VSS.n2153 0.04025
R16335 VSS.n7236 VSS.n2153 0.04025
R16336 VSS.n7236 VSS.n7235 0.04025
R16337 VSS.n7235 VSS.n7234 0.04025
R16338 VSS.n7234 VSS.n2155 0.04025
R16339 VSS.n7230 VSS.n2155 0.04025
R16340 VSS.n7230 VSS.n7229 0.04025
R16341 VSS.n7229 VSS.n7228 0.04025
R16342 VSS.n7228 VSS.n2157 0.04025
R16343 VSS.n7224 VSS.n2157 0.04025
R16344 VSS.n7224 VSS.n7223 0.04025
R16345 VSS.n7223 VSS.n7222 0.04025
R16346 VSS.n7222 VSS.n2159 0.04025
R16347 VSS.n7218 VSS.n2159 0.04025
R16348 VSS.n7218 VSS.n7217 0.04025
R16349 VSS.n7217 VSS.n7216 0.04025
R16350 VSS.n7216 VSS.n2161 0.04025
R16351 VSS.n7212 VSS.n2161 0.04025
R16352 VSS.n7212 VSS.n7211 0.04025
R16353 VSS.n7211 VSS.n7210 0.04025
R16354 VSS.n7210 VSS.n2163 0.04025
R16355 VSS.n7206 VSS.n2163 0.04025
R16356 VSS.n7206 VSS.n7205 0.04025
R16357 VSS.n7205 VSS.n7204 0.04025
R16358 VSS.n7204 VSS.n2165 0.04025
R16359 VSS.n7200 VSS.n2165 0.04025
R16360 VSS.n7200 VSS.n7199 0.04025
R16361 VSS.n7199 VSS.n7198 0.04025
R16362 VSS.n7198 VSS.n2167 0.04025
R16363 VSS.n7194 VSS.n2167 0.04025
R16364 VSS.n7194 VSS.n7193 0.04025
R16365 VSS.n7193 VSS.n7192 0.04025
R16366 VSS.n7192 VSS.n2169 0.04025
R16367 VSS.n7188 VSS.n2169 0.04025
R16368 VSS.n7188 VSS.n7187 0.04025
R16369 VSS.n7187 VSS.n7186 0.04025
R16370 VSS.n7186 VSS.n2171 0.04025
R16371 VSS.n7182 VSS.n2171 0.04025
R16372 VSS.n7182 VSS.n7181 0.04025
R16373 VSS.n7181 VSS.n7180 0.04025
R16374 VSS.n7180 VSS.n2173 0.04025
R16375 VSS.n7176 VSS.n2173 0.04025
R16376 VSS.n7176 VSS.n7175 0.04025
R16377 VSS.n7175 VSS.n7174 0.04025
R16378 VSS.n7174 VSS.n2175 0.04025
R16379 VSS.n7170 VSS.n2175 0.04025
R16380 VSS.n7170 VSS.n7169 0.04025
R16381 VSS.n7169 VSS.n7168 0.04025
R16382 VSS.n7168 VSS.n2177 0.04025
R16383 VSS.n7164 VSS.n2177 0.04025
R16384 VSS.n7164 VSS.n7163 0.04025
R16385 VSS.n7163 VSS.n7162 0.04025
R16386 VSS.n7162 VSS.n2179 0.04025
R16387 VSS.n7158 VSS.n2179 0.04025
R16388 VSS.n7158 VSS.n7157 0.04025
R16389 VSS.n7157 VSS.n7156 0.04025
R16390 VSS.n7156 VSS.n2181 0.04025
R16391 VSS.n7152 VSS.n2181 0.04025
R16392 VSS.n7152 VSS.n7151 0.04025
R16393 VSS.n7151 VSS.n7150 0.04025
R16394 VSS.n7150 VSS.n2183 0.04025
R16395 VSS.n7146 VSS.n2183 0.04025
R16396 VSS.n7146 VSS.n7145 0.04025
R16397 VSS.n7145 VSS.n7144 0.04025
R16398 VSS.n7144 VSS.n2185 0.04025
R16399 VSS.n7140 VSS.n2185 0.04025
R16400 VSS.n7140 VSS.n7139 0.04025
R16401 VSS.n7139 VSS.n7138 0.04025
R16402 VSS.n7138 VSS.n2187 0.04025
R16403 VSS.n7134 VSS.n2187 0.04025
R16404 VSS.n7134 VSS.n7133 0.04025
R16405 VSS.n7133 VSS.n7132 0.04025
R16406 VSS.n7132 VSS.n2189 0.04025
R16407 VSS.n7128 VSS.n2189 0.04025
R16408 VSS.n7128 VSS.n7127 0.04025
R16409 VSS.n7127 VSS.n7126 0.04025
R16410 VSS.n7126 VSS.n2191 0.04025
R16411 VSS.n7122 VSS.n2191 0.04025
R16412 VSS.n7122 VSS.n7121 0.04025
R16413 VSS.n7121 VSS.n7120 0.04025
R16414 VSS.n7120 VSS.n2193 0.04025
R16415 VSS.n7116 VSS.n2193 0.04025
R16416 VSS.n7116 VSS.n7115 0.04025
R16417 VSS.n7115 VSS.n7114 0.04025
R16418 VSS.n7114 VSS.n2195 0.04025
R16419 VSS.n7110 VSS.n2195 0.04025
R16420 VSS.n7110 VSS.n7109 0.04025
R16421 VSS.n7109 VSS.n7108 0.04025
R16422 VSS.n7108 VSS.n2197 0.04025
R16423 VSS.n7104 VSS.n2197 0.04025
R16424 VSS.n7104 VSS.n7103 0.04025
R16425 VSS.n7103 VSS.n7102 0.04025
R16426 VSS.n7102 VSS.n2199 0.04025
R16427 VSS.n7098 VSS.n2199 0.04025
R16428 VSS.n7098 VSS.n7097 0.04025
R16429 VSS.n7097 VSS.n7096 0.04025
R16430 VSS.n7096 VSS.n2201 0.04025
R16431 VSS.n7092 VSS.n2201 0.04025
R16432 VSS.n7092 VSS.n7091 0.04025
R16433 VSS.n7091 VSS.n7090 0.04025
R16434 VSS.n7090 VSS.n2203 0.04025
R16435 VSS.n7086 VSS.n2203 0.04025
R16436 VSS.n7086 VSS.n7085 0.04025
R16437 VSS.n7085 VSS.n7084 0.04025
R16438 VSS.n7084 VSS.n2205 0.04025
R16439 VSS.n7080 VSS.n2205 0.04025
R16440 VSS.n7080 VSS.n7079 0.04025
R16441 VSS.n7079 VSS.n7078 0.04025
R16442 VSS.n7078 VSS.n2207 0.04025
R16443 VSS.n7074 VSS.n2207 0.04025
R16444 VSS.n7074 VSS.n7073 0.04025
R16445 VSS.n7073 VSS.n7072 0.04025
R16446 VSS.n7072 VSS.n2209 0.04025
R16447 VSS.n7068 VSS.n2209 0.04025
R16448 VSS.n7068 VSS.n7067 0.04025
R16449 VSS.n7067 VSS.n7066 0.04025
R16450 VSS.n7066 VSS.n2211 0.04025
R16451 VSS.n7062 VSS.n2211 0.04025
R16452 VSS.n7062 VSS.n7061 0.04025
R16453 VSS.n7061 VSS.n7060 0.04025
R16454 VSS.n7060 VSS.n2213 0.04025
R16455 VSS.n7056 VSS.n2213 0.04025
R16456 VSS.n7056 VSS.n7055 0.04025
R16457 VSS.n7055 VSS.n7054 0.04025
R16458 VSS.n7054 VSS.n2215 0.04025
R16459 VSS.n7050 VSS.n2215 0.04025
R16460 VSS.n7050 VSS.n7049 0.04025
R16461 VSS.n7049 VSS.n7048 0.04025
R16462 VSS.n7048 VSS.n2217 0.04025
R16463 VSS.n7044 VSS.n2217 0.04025
R16464 VSS.n7044 VSS.n7043 0.04025
R16465 VSS.n7043 VSS.n7042 0.04025
R16466 VSS.n7042 VSS.n2219 0.04025
R16467 VSS.n7038 VSS.n2219 0.04025
R16468 VSS.n7038 VSS.n7037 0.04025
R16469 VSS.n7037 VSS.n7036 0.04025
R16470 VSS.n7036 VSS.n2221 0.04025
R16471 VSS.n7032 VSS.n2221 0.04025
R16472 VSS.n7032 VSS.n7031 0.04025
R16473 VSS.n7031 VSS.n7030 0.04025
R16474 VSS.n7030 VSS.n2223 0.04025
R16475 VSS.n7026 VSS.n2223 0.04025
R16476 VSS.n7026 VSS.n7025 0.04025
R16477 VSS.n7025 VSS.n7024 0.04025
R16478 VSS.n7024 VSS.n2225 0.04025
R16479 VSS.n7020 VSS.n2225 0.04025
R16480 VSS.n7020 VSS.n7019 0.04025
R16481 VSS.n7019 VSS.n7018 0.04025
R16482 VSS.n7018 VSS.n2227 0.04025
R16483 VSS.n7014 VSS.n2227 0.04025
R16484 VSS.n7014 VSS.n7013 0.04025
R16485 VSS.n7013 VSS.n7012 0.04025
R16486 VSS.n7012 VSS.n2229 0.04025
R16487 VSS.n7008 VSS.n2229 0.04025
R16488 VSS.n7008 VSS.n7007 0.04025
R16489 VSS.n7007 VSS.n7006 0.04025
R16490 VSS.n7006 VSS.n2231 0.04025
R16491 VSS.n7002 VSS.n2231 0.04025
R16492 VSS.n7002 VSS.n7001 0.04025
R16493 VSS.n7001 VSS.n7000 0.04025
R16494 VSS.n7000 VSS.n2233 0.04025
R16495 VSS.n6996 VSS.n2233 0.04025
R16496 VSS.n6996 VSS.n6995 0.04025
R16497 VSS.n6995 VSS.n6994 0.04025
R16498 VSS.n6994 VSS.n2235 0.04025
R16499 VSS.n6990 VSS.n2235 0.04025
R16500 VSS.n6990 VSS.n6989 0.04025
R16501 VSS.n6989 VSS.n6988 0.04025
R16502 VSS.n6988 VSS.n2237 0.04025
R16503 VSS.n6984 VSS.n2237 0.04025
R16504 VSS.n6984 VSS.n6983 0.04025
R16505 VSS.n6983 VSS.n6982 0.04025
R16506 VSS.n6982 VSS.n2239 0.04025
R16507 VSS.n6978 VSS.n2239 0.04025
R16508 VSS.n6978 VSS.n6977 0.04025
R16509 VSS.n6977 VSS.n6976 0.04025
R16510 VSS.n6976 VSS.n2241 0.04025
R16511 VSS.n6972 VSS.n2241 0.04025
R16512 VSS.n6972 VSS.n6971 0.04025
R16513 VSS.n6971 VSS.n6970 0.04025
R16514 VSS.n6970 VSS.n2243 0.04025
R16515 VSS.n6966 VSS.n2243 0.04025
R16516 VSS.n6966 VSS.n6965 0.04025
R16517 VSS.n6965 VSS.n6964 0.04025
R16518 VSS.n6964 VSS.n2245 0.04025
R16519 VSS.n6960 VSS.n2245 0.04025
R16520 VSS.n6960 VSS.n6959 0.04025
R16521 VSS.n6959 VSS.n6958 0.04025
R16522 VSS.n6958 VSS.n2247 0.04025
R16523 VSS.n6954 VSS.n2247 0.04025
R16524 VSS.n6954 VSS.n6953 0.04025
R16525 VSS.n6953 VSS.n6952 0.04025
R16526 VSS.n6952 VSS.n2249 0.04025
R16527 VSS.n6948 VSS.n2249 0.04025
R16528 VSS.n6948 VSS.n6947 0.04025
R16529 VSS.n6947 VSS.n6946 0.04025
R16530 VSS.n6946 VSS.n2251 0.04025
R16531 VSS.n6942 VSS.n2251 0.04025
R16532 VSS.n6942 VSS.n6941 0.04025
R16533 VSS.n6941 VSS.n6940 0.04025
R16534 VSS.n6940 VSS.n2253 0.04025
R16535 VSS.n6936 VSS.n6935 0.04025
R16536 VSS.n6935 VSS.n6934 0.04025
R16537 VSS.n6934 VSS.n2255 0.04025
R16538 VSS.n6930 VSS.n2255 0.04025
R16539 VSS.n6930 VSS.n6929 0.04025
R16540 VSS.n6929 VSS.n6928 0.04025
R16541 VSS.n6928 VSS.n2257 0.04025
R16542 VSS.n6924 VSS.n2257 0.04025
R16543 VSS.n6924 VSS.n6923 0.04025
R16544 VSS.n6923 VSS.n6922 0.04025
R16545 VSS.n6922 VSS.n2259 0.04025
R16546 VSS.n6918 VSS.n2259 0.04025
R16547 VSS.n6918 VSS.n6917 0.04025
R16548 VSS.n6917 VSS.n6916 0.04025
R16549 VSS.n6916 VSS.n2261 0.04025
R16550 VSS.n6912 VSS.n2261 0.04025
R16551 VSS.n6912 VSS.n6911 0.04025
R16552 VSS.n6911 VSS.n6910 0.04025
R16553 VSS.n6910 VSS.n2263 0.04025
R16554 VSS.n4141 VSS.n3185 0.04025
R16555 VSS.n4137 VSS.n3185 0.04025
R16556 VSS.n4137 VSS.n4136 0.04025
R16557 VSS.n4136 VSS.n4135 0.04025
R16558 VSS.n4135 VSS.n3187 0.04025
R16559 VSS.n4131 VSS.n3187 0.04025
R16560 VSS.n4131 VSS.n4130 0.04025
R16561 VSS.n4130 VSS.n4129 0.04025
R16562 VSS.n4129 VSS.n3189 0.04025
R16563 VSS.n4125 VSS.n3189 0.04025
R16564 VSS.n4125 VSS.n4124 0.04025
R16565 VSS.n4124 VSS.n4123 0.04025
R16566 VSS.n4123 VSS.n3191 0.04025
R16567 VSS.n4119 VSS.n3191 0.04025
R16568 VSS.n4119 VSS.n4118 0.04025
R16569 VSS.n4118 VSS.n4117 0.04025
R16570 VSS.n4117 VSS.n3193 0.04025
R16571 VSS.n4113 VSS.n3193 0.04025
R16572 VSS.n4113 VSS.n4112 0.04025
R16573 VSS.n4112 VSS.n4111 0.04025
R16574 VSS.n4111 VSS.n3195 0.04025
R16575 VSS.n4107 VSS.n3195 0.04025
R16576 VSS.n4107 VSS.n4106 0.04025
R16577 VSS.n4106 VSS.n4105 0.04025
R16578 VSS.n4105 VSS.n3197 0.04025
R16579 VSS.n4101 VSS.n3197 0.04025
R16580 VSS.n4101 VSS.n4100 0.04025
R16581 VSS.n4100 VSS.n4099 0.04025
R16582 VSS.n4099 VSS.n3199 0.04025
R16583 VSS.n4095 VSS.n3199 0.04025
R16584 VSS.n4095 VSS.n4094 0.04025
R16585 VSS.n4094 VSS.n4093 0.04025
R16586 VSS.n4093 VSS.n3201 0.04025
R16587 VSS.n4089 VSS.n3201 0.04025
R16588 VSS.n4089 VSS.n4088 0.04025
R16589 VSS.n4088 VSS.n4087 0.04025
R16590 VSS.n4087 VSS.n3203 0.04025
R16591 VSS.n4083 VSS.n3203 0.04025
R16592 VSS.n4083 VSS.n4082 0.04025
R16593 VSS.n4082 VSS.n4081 0.04025
R16594 VSS.n4081 VSS.n3205 0.04025
R16595 VSS.n4077 VSS.n3205 0.04025
R16596 VSS.n4077 VSS.n4076 0.04025
R16597 VSS.n4076 VSS.n4075 0.04025
R16598 VSS.n4075 VSS.n3207 0.04025
R16599 VSS.n4071 VSS.n3207 0.04025
R16600 VSS.n4071 VSS.n4070 0.04025
R16601 VSS.n4070 VSS.n4069 0.04025
R16602 VSS.n4069 VSS.n3209 0.04025
R16603 VSS.n4065 VSS.n3209 0.04025
R16604 VSS.n4065 VSS.n4064 0.04025
R16605 VSS.n4064 VSS.n4063 0.04025
R16606 VSS.n4063 VSS.n3211 0.04025
R16607 VSS.n4059 VSS.n3211 0.04025
R16608 VSS.n4059 VSS.n4058 0.04025
R16609 VSS.n4058 VSS.n4057 0.04025
R16610 VSS.n4057 VSS.n3213 0.04025
R16611 VSS.n4053 VSS.n3213 0.04025
R16612 VSS.n4053 VSS.n4052 0.04025
R16613 VSS.n4052 VSS.n4051 0.04025
R16614 VSS.n4051 VSS.n3215 0.04025
R16615 VSS.n4047 VSS.n3215 0.04025
R16616 VSS.n4047 VSS.n4046 0.04025
R16617 VSS.n4046 VSS.n4045 0.04025
R16618 VSS.n4045 VSS.n3217 0.04025
R16619 VSS.n4041 VSS.n3217 0.04025
R16620 VSS.n4041 VSS.n4040 0.04025
R16621 VSS.n4040 VSS.n4039 0.04025
R16622 VSS.n4039 VSS.n3219 0.04025
R16623 VSS.n4035 VSS.n3219 0.04025
R16624 VSS.n4035 VSS.n4034 0.04025
R16625 VSS.n4034 VSS.n4033 0.04025
R16626 VSS.n4033 VSS.n3221 0.04025
R16627 VSS.n4029 VSS.n3221 0.04025
R16628 VSS.n4029 VSS.n4028 0.04025
R16629 VSS.n4028 VSS.n4027 0.04025
R16630 VSS.n4027 VSS.n3223 0.04025
R16631 VSS.n4023 VSS.n3223 0.04025
R16632 VSS.n4023 VSS.n4022 0.04025
R16633 VSS.n4022 VSS.n4021 0.04025
R16634 VSS.n4021 VSS.n3225 0.04025
R16635 VSS.n4017 VSS.n3225 0.04025
R16636 VSS.n4017 VSS.n4016 0.04025
R16637 VSS.n4016 VSS.n4015 0.04025
R16638 VSS.n4015 VSS.n3227 0.04025
R16639 VSS.n4011 VSS.n3227 0.04025
R16640 VSS.n4011 VSS.n4010 0.04025
R16641 VSS.n4010 VSS.n4009 0.04025
R16642 VSS.n4009 VSS.n3229 0.04025
R16643 VSS.n4005 VSS.n3229 0.04025
R16644 VSS.n4005 VSS.n4004 0.04025
R16645 VSS.n4004 VSS.n4003 0.04025
R16646 VSS.n4003 VSS.n3231 0.04025
R16647 VSS.n3999 VSS.n3231 0.04025
R16648 VSS.n3999 VSS.n3998 0.04025
R16649 VSS.n3998 VSS.n3997 0.04025
R16650 VSS.n3997 VSS.n3233 0.04025
R16651 VSS.n3993 VSS.n3233 0.04025
R16652 VSS.n3993 VSS.n3992 0.04025
R16653 VSS.n3992 VSS.n3991 0.04025
R16654 VSS.n3991 VSS.n3235 0.04025
R16655 VSS.n3987 VSS.n3235 0.04025
R16656 VSS.n3987 VSS.n3986 0.04025
R16657 VSS.n3986 VSS.n3985 0.04025
R16658 VSS.n3985 VSS.n3237 0.04025
R16659 VSS.n3981 VSS.n3237 0.04025
R16660 VSS.n3981 VSS.n3980 0.04025
R16661 VSS.n3980 VSS.n3979 0.04025
R16662 VSS.n3979 VSS.n3239 0.04025
R16663 VSS.n3975 VSS.n3239 0.04025
R16664 VSS.n3975 VSS.n3974 0.04025
R16665 VSS.n3974 VSS.n3973 0.04025
R16666 VSS.n3973 VSS.n3241 0.04025
R16667 VSS.n3969 VSS.n3241 0.04025
R16668 VSS.n3969 VSS.n3968 0.04025
R16669 VSS.n3968 VSS.n3967 0.04025
R16670 VSS.n3967 VSS.n3243 0.04025
R16671 VSS.n3963 VSS.n3243 0.04025
R16672 VSS.n3963 VSS.n3962 0.04025
R16673 VSS.n3962 VSS.n3961 0.04025
R16674 VSS.n3961 VSS.n3245 0.04025
R16675 VSS.n3957 VSS.n3245 0.04025
R16676 VSS.n3957 VSS.n3956 0.04025
R16677 VSS.n3956 VSS.n3955 0.04025
R16678 VSS.n3955 VSS.n3247 0.04025
R16679 VSS.n3951 VSS.n3247 0.04025
R16680 VSS.n3951 VSS.n3950 0.04025
R16681 VSS.n3950 VSS.n3949 0.04025
R16682 VSS.n3949 VSS.n3249 0.04025
R16683 VSS.n3945 VSS.n3249 0.04025
R16684 VSS.n3945 VSS.n3944 0.04025
R16685 VSS.n3944 VSS.n3943 0.04025
R16686 VSS.n3943 VSS.n3251 0.04025
R16687 VSS.n3939 VSS.n3251 0.04025
R16688 VSS.n3939 VSS.n3938 0.04025
R16689 VSS.n3938 VSS.n3937 0.04025
R16690 VSS.n3937 VSS.n3253 0.04025
R16691 VSS.n3933 VSS.n3253 0.04025
R16692 VSS.n3933 VSS.n3932 0.04025
R16693 VSS.n3932 VSS.n3931 0.04025
R16694 VSS.n3931 VSS.n3255 0.04025
R16695 VSS.n3927 VSS.n3255 0.04025
R16696 VSS.n3927 VSS.n3926 0.04025
R16697 VSS.n3926 VSS.n3925 0.04025
R16698 VSS.n3925 VSS.n3257 0.04025
R16699 VSS.n3921 VSS.n3257 0.04025
R16700 VSS.n3921 VSS.n3920 0.04025
R16701 VSS.n3920 VSS.n3919 0.04025
R16702 VSS.n3919 VSS.n3259 0.04025
R16703 VSS.n3915 VSS.n3259 0.04025
R16704 VSS.n3915 VSS.n3914 0.04025
R16705 VSS.n3914 VSS.n3913 0.04025
R16706 VSS.n3913 VSS.n3261 0.04025
R16707 VSS.n3909 VSS.n3261 0.04025
R16708 VSS.n3909 VSS.n3908 0.04025
R16709 VSS.n3908 VSS.n3907 0.04025
R16710 VSS.n3907 VSS.n3263 0.04025
R16711 VSS.n3903 VSS.n3263 0.04025
R16712 VSS.n3903 VSS.n3902 0.04025
R16713 VSS.n3902 VSS.n3901 0.04025
R16714 VSS.n3901 VSS.n3265 0.04025
R16715 VSS.n3897 VSS.n3265 0.04025
R16716 VSS.n3897 VSS.n3896 0.04025
R16717 VSS.n3896 VSS.n3895 0.04025
R16718 VSS.n3895 VSS.n3267 0.04025
R16719 VSS.n3891 VSS.n3267 0.04025
R16720 VSS.n3891 VSS.n3890 0.04025
R16721 VSS.n3890 VSS.n3889 0.04025
R16722 VSS.n3889 VSS.n3269 0.04025
R16723 VSS.n3885 VSS.n3269 0.04025
R16724 VSS.n3885 VSS.n3884 0.04025
R16725 VSS.n3884 VSS.n3883 0.04025
R16726 VSS.n3883 VSS.n3271 0.04025
R16727 VSS.n3879 VSS.n3271 0.04025
R16728 VSS.n3879 VSS.n3878 0.04025
R16729 VSS.n3878 VSS.n3877 0.04025
R16730 VSS.n3877 VSS.n3273 0.04025
R16731 VSS.n3873 VSS.n3273 0.04025
R16732 VSS.n3873 VSS.n3872 0.04025
R16733 VSS.n3872 VSS.n3871 0.04025
R16734 VSS.n3871 VSS.n3275 0.04025
R16735 VSS.n3867 VSS.n3275 0.04025
R16736 VSS.n3867 VSS.n3866 0.04025
R16737 VSS.n3866 VSS.n3865 0.04025
R16738 VSS.n3865 VSS.n3277 0.04025
R16739 VSS.n3861 VSS.n3277 0.04025
R16740 VSS.n3861 VSS.n3860 0.04025
R16741 VSS.n3860 VSS.n3859 0.04025
R16742 VSS.n3859 VSS.n3279 0.04025
R16743 VSS.n3855 VSS.n3279 0.04025
R16744 VSS.n3855 VSS.n3854 0.04025
R16745 VSS.n3854 VSS.n3853 0.04025
R16746 VSS.n3853 VSS.n3281 0.04025
R16747 VSS.n3849 VSS.n3281 0.04025
R16748 VSS.n3849 VSS.n3848 0.04025
R16749 VSS.n3848 VSS.n3847 0.04025
R16750 VSS.n3847 VSS.n3283 0.04025
R16751 VSS.n3843 VSS.n3283 0.04025
R16752 VSS.n3843 VSS.n3842 0.04025
R16753 VSS.n3842 VSS.n3841 0.04025
R16754 VSS.n3841 VSS.n3285 0.04025
R16755 VSS.n3837 VSS.n3285 0.04025
R16756 VSS.n3837 VSS.n3836 0.04025
R16757 VSS.n3836 VSS.n3835 0.04025
R16758 VSS.n3835 VSS.n3287 0.04025
R16759 VSS.n3831 VSS.n3287 0.04025
R16760 VSS.n3831 VSS.n3830 0.04025
R16761 VSS.n3830 VSS.n3829 0.04025
R16762 VSS.n3829 VSS.n3289 0.04025
R16763 VSS.n3825 VSS.n3289 0.04025
R16764 VSS.n3825 VSS.n3824 0.04025
R16765 VSS.n3824 VSS.n3823 0.04025
R16766 VSS.n3823 VSS.n3291 0.04025
R16767 VSS.n3819 VSS.n3291 0.04025
R16768 VSS.n3819 VSS.n3818 0.04025
R16769 VSS.n3818 VSS.n3817 0.04025
R16770 VSS.n3817 VSS.n3293 0.04025
R16771 VSS.n3813 VSS.n3293 0.04025
R16772 VSS.n3813 VSS.n3812 0.04025
R16773 VSS.n3812 VSS.n3811 0.04025
R16774 VSS.n3811 VSS.n3295 0.04025
R16775 VSS.n3807 VSS.n3295 0.04025
R16776 VSS.n3807 VSS.n3806 0.04025
R16777 VSS.n3806 VSS.n3805 0.04025
R16778 VSS.n3805 VSS.n3297 0.04025
R16779 VSS.n3801 VSS.n3297 0.04025
R16780 VSS.n3801 VSS.n3800 0.04025
R16781 VSS.n3800 VSS.n3799 0.04025
R16782 VSS.n3799 VSS.n3299 0.04025
R16783 VSS.n3795 VSS.n3299 0.04025
R16784 VSS.n3795 VSS.n3794 0.04025
R16785 VSS.n3794 VSS.n3793 0.04025
R16786 VSS.n3793 VSS.n3301 0.04025
R16787 VSS.n3789 VSS.n3301 0.04025
R16788 VSS.n3789 VSS.n3788 0.04025
R16789 VSS.n3788 VSS.n3787 0.04025
R16790 VSS.n3787 VSS.n3303 0.04025
R16791 VSS.n3783 VSS.n3303 0.04025
R16792 VSS.n3783 VSS.n3782 0.04025
R16793 VSS.n3782 VSS.n3781 0.04025
R16794 VSS.n3781 VSS.n3305 0.04025
R16795 VSS.n3777 VSS.n3305 0.04025
R16796 VSS.n3777 VSS.n3776 0.04025
R16797 VSS.n3776 VSS.n3775 0.04025
R16798 VSS.n3775 VSS.n3307 0.04025
R16799 VSS.n3771 VSS.n3307 0.04025
R16800 VSS.n3771 VSS.n3770 0.04025
R16801 VSS.n3770 VSS.n3769 0.04025
R16802 VSS.n3769 VSS.n3309 0.04025
R16803 VSS.n3765 VSS.n3309 0.04025
R16804 VSS.n3765 VSS.n3764 0.04025
R16805 VSS.n3764 VSS.n3763 0.04025
R16806 VSS.n3763 VSS.n3311 0.04025
R16807 VSS.n3759 VSS.n3311 0.04025
R16808 VSS.n3759 VSS.n3758 0.04025
R16809 VSS.n3758 VSS.n3757 0.04025
R16810 VSS.n3757 VSS.n3313 0.04025
R16811 VSS.n3753 VSS.n3313 0.04025
R16812 VSS.n3753 VSS.n3752 0.04025
R16813 VSS.n3752 VSS.n3751 0.04025
R16814 VSS.n3751 VSS.n3315 0.04025
R16815 VSS.n3747 VSS.n3315 0.04025
R16816 VSS.n3747 VSS.n3746 0.04025
R16817 VSS.n3746 VSS.n3745 0.04025
R16818 VSS.n3745 VSS.n3317 0.04025
R16819 VSS.n3741 VSS.n3317 0.04025
R16820 VSS.n3741 VSS.n3740 0.04025
R16821 VSS.n3740 VSS.n3739 0.04025
R16822 VSS.n3739 VSS.n3319 0.04025
R16823 VSS.n3735 VSS.n3319 0.04025
R16824 VSS.n3735 VSS.n3734 0.04025
R16825 VSS.n3734 VSS.n3733 0.04025
R16826 VSS.n3733 VSS.n3321 0.04025
R16827 VSS.n3729 VSS.n3321 0.04025
R16828 VSS.n3729 VSS.n3728 0.04025
R16829 VSS.n3728 VSS.n3727 0.04025
R16830 VSS.n3727 VSS.n3323 0.04025
R16831 VSS.n3723 VSS.n3323 0.04025
R16832 VSS.n3723 VSS.n3722 0.04025
R16833 VSS.n3722 VSS.n3721 0.04025
R16834 VSS.n3721 VSS.n3325 0.04025
R16835 VSS.n3717 VSS.n3325 0.04025
R16836 VSS.n3717 VSS.n3716 0.04025
R16837 VSS.n3716 VSS.n3715 0.04025
R16838 VSS.n3715 VSS.n3327 0.04025
R16839 VSS.n3711 VSS.n3327 0.04025
R16840 VSS.n3711 VSS.n3710 0.04025
R16841 VSS.n3710 VSS.n3709 0.04025
R16842 VSS.n3709 VSS.n3329 0.04025
R16843 VSS.n3705 VSS.n3329 0.04025
R16844 VSS.n3705 VSS.n3704 0.04025
R16845 VSS.n3704 VSS.n3703 0.04025
R16846 VSS.n3703 VSS.n3331 0.04025
R16847 VSS.n3699 VSS.n3331 0.04025
R16848 VSS.n3699 VSS.n3698 0.04025
R16849 VSS.n3698 VSS.n3697 0.04025
R16850 VSS.n3697 VSS.n3333 0.04025
R16851 VSS.n3693 VSS.n3333 0.04025
R16852 VSS.n3693 VSS.n3692 0.04025
R16853 VSS.n3692 VSS.n3691 0.04025
R16854 VSS.n3691 VSS.n3335 0.04025
R16855 VSS.n3687 VSS.n3335 0.04025
R16856 VSS.n3687 VSS.n3686 0.04025
R16857 VSS.n3686 VSS.n3685 0.04025
R16858 VSS.n3685 VSS.n3337 0.04025
R16859 VSS.n3681 VSS.n3337 0.04025
R16860 VSS.n3681 VSS.n3680 0.04025
R16861 VSS.n3680 VSS.n3679 0.04025
R16862 VSS.n3679 VSS.n3339 0.04025
R16863 VSS.n3675 VSS.n3339 0.04025
R16864 VSS.n3675 VSS.n3674 0.04025
R16865 VSS.n3674 VSS.n3673 0.04025
R16866 VSS.n3673 VSS.n3341 0.04025
R16867 VSS.n3669 VSS.n3341 0.04025
R16868 VSS.n3669 VSS.n3668 0.04025
R16869 VSS.n3668 VSS.n3667 0.04025
R16870 VSS.n3667 VSS.n3343 0.04025
R16871 VSS.n3663 VSS.n3343 0.04025
R16872 VSS.n3663 VSS.n3662 0.04025
R16873 VSS.n3662 VSS.n3661 0.04025
R16874 VSS.n3661 VSS.n3345 0.04025
R16875 VSS.n3657 VSS.n3345 0.04025
R16876 VSS.n3657 VSS.n3656 0.04025
R16877 VSS.n3656 VSS.n3655 0.04025
R16878 VSS.n3655 VSS.n3347 0.04025
R16879 VSS.n3651 VSS.n3347 0.04025
R16880 VSS.n3651 VSS.n3650 0.04025
R16881 VSS.n3650 VSS.n3649 0.04025
R16882 VSS.n3649 VSS.n3349 0.04025
R16883 VSS.n3645 VSS.n3349 0.04025
R16884 VSS.n3645 VSS.n3644 0.04025
R16885 VSS.n3644 VSS.n3643 0.04025
R16886 VSS.n3643 VSS.n3351 0.04025
R16887 VSS.n3639 VSS.n3351 0.04025
R16888 VSS.n3639 VSS.n3638 0.04025
R16889 VSS.n3638 VSS.n3637 0.04025
R16890 VSS.n3637 VSS.n3353 0.04025
R16891 VSS.n3633 VSS.n3353 0.04025
R16892 VSS.n3633 VSS.n3632 0.04025
R16893 VSS.n3632 VSS.n3631 0.04025
R16894 VSS.n3631 VSS.n3355 0.04025
R16895 VSS.n3627 VSS.n3355 0.04025
R16896 VSS.n3627 VSS.n3626 0.04025
R16897 VSS.n3626 VSS.n3625 0.04025
R16898 VSS.n3625 VSS.n3357 0.04025
R16899 VSS.n3621 VSS.n3357 0.04025
R16900 VSS.n3621 VSS.n3620 0.04025
R16901 VSS.n3620 VSS.n3619 0.04025
R16902 VSS.n3619 VSS.n3359 0.04025
R16903 VSS.n3615 VSS.n3359 0.04025
R16904 VSS.n3615 VSS.n3614 0.04025
R16905 VSS.n3614 VSS.n3613 0.04025
R16906 VSS.n3613 VSS.n3361 0.04025
R16907 VSS.n3609 VSS.n3361 0.04025
R16908 VSS.n3609 VSS.n3608 0.04025
R16909 VSS.n3608 VSS.n3607 0.04025
R16910 VSS.n3607 VSS.n3363 0.04025
R16911 VSS.n3603 VSS.n3363 0.04025
R16912 VSS.n3603 VSS.n3602 0.04025
R16913 VSS.n3602 VSS.n3601 0.04025
R16914 VSS.n3601 VSS.n3365 0.04025
R16915 VSS.n3597 VSS.n3365 0.04025
R16916 VSS.n3597 VSS.n3596 0.04025
R16917 VSS.n3596 VSS.n3595 0.04025
R16918 VSS.n3595 VSS.n3367 0.04025
R16919 VSS.n3591 VSS.n3367 0.04025
R16920 VSS.n3591 VSS.n3590 0.04025
R16921 VSS.n3590 VSS.n3589 0.04025
R16922 VSS.n3589 VSS.n3369 0.04025
R16923 VSS.n3585 VSS.n3369 0.04025
R16924 VSS.n3585 VSS.n3584 0.04025
R16925 VSS.n3584 VSS.n3583 0.04025
R16926 VSS.n3583 VSS.n3371 0.04025
R16927 VSS.n3579 VSS.n3371 0.04025
R16928 VSS.n3579 VSS.n3578 0.04025
R16929 VSS.n3578 VSS.n3577 0.04025
R16930 VSS.n3577 VSS.n3373 0.04025
R16931 VSS.n3573 VSS.n3373 0.04025
R16932 VSS.n3573 VSS.n3572 0.04025
R16933 VSS.n3572 VSS.n3571 0.04025
R16934 VSS.n3571 VSS.n3375 0.04025
R16935 VSS.n3567 VSS.n3375 0.04025
R16936 VSS.n3567 VSS.n3566 0.04025
R16937 VSS.n3566 VSS.n3565 0.04025
R16938 VSS.n3565 VSS.n3377 0.04025
R16939 VSS.n3561 VSS.n3377 0.04025
R16940 VSS.n3561 VSS.n3560 0.04025
R16941 VSS.n3560 VSS.n3559 0.04025
R16942 VSS.n3559 VSS.n3379 0.04025
R16943 VSS.n3555 VSS.n3379 0.04025
R16944 VSS.n3555 VSS.n3554 0.04025
R16945 VSS.n3554 VSS.n3553 0.04025
R16946 VSS.n3553 VSS.n3381 0.04025
R16947 VSS.n3549 VSS.n3381 0.04025
R16948 VSS.n3549 VSS.n3548 0.04025
R16949 VSS.n3548 VSS.n3547 0.04025
R16950 VSS.n3547 VSS.n3383 0.04025
R16951 VSS.n3543 VSS.n3383 0.04025
R16952 VSS.n3543 VSS.n3542 0.04025
R16953 VSS.n3542 VSS.n3541 0.04025
R16954 VSS.n3541 VSS.n3385 0.04025
R16955 VSS.n3537 VSS.n3385 0.04025
R16956 VSS.n3537 VSS.n3536 0.04025
R16957 VSS.n3536 VSS.n3535 0.04025
R16958 VSS.n3535 VSS.n3387 0.04025
R16959 VSS.n3531 VSS.n3387 0.04025
R16960 VSS.n3531 VSS.n3530 0.04025
R16961 VSS.n3530 VSS.n3529 0.04025
R16962 VSS.n3529 VSS.n3389 0.04025
R16963 VSS.n3525 VSS.n3389 0.04025
R16964 VSS.n3525 VSS.n3524 0.04025
R16965 VSS.n3524 VSS.n3523 0.04025
R16966 VSS.n3523 VSS.n3391 0.04025
R16967 VSS.n3519 VSS.n3391 0.04025
R16968 VSS.n3519 VSS.n3518 0.04025
R16969 VSS.n3518 VSS.n3517 0.04025
R16970 VSS.n3517 VSS.n3393 0.04025
R16971 VSS.n3513 VSS.n3393 0.04025
R16972 VSS.n3513 VSS.n3512 0.04025
R16973 VSS.n3512 VSS.n3511 0.04025
R16974 VSS.n3511 VSS.n3395 0.04025
R16975 VSS.n3507 VSS.n3395 0.04025
R16976 VSS.n3507 VSS.n3506 0.04025
R16977 VSS.n3506 VSS.n3505 0.04025
R16978 VSS.n3505 VSS.n3397 0.04025
R16979 VSS.n3501 VSS.n3397 0.04025
R16980 VSS.n3501 VSS.n3500 0.04025
R16981 VSS.n3500 VSS.n3499 0.04025
R16982 VSS.n3499 VSS.n3399 0.04025
R16983 VSS.n3495 VSS.n3399 0.04025
R16984 VSS.n3495 VSS.n3494 0.04025
R16985 VSS.n3494 VSS.n3493 0.04025
R16986 VSS.n3493 VSS.n3401 0.04025
R16987 VSS.n3489 VSS.n3401 0.04025
R16988 VSS.n3489 VSS.n3488 0.04025
R16989 VSS.n3488 VSS.n3487 0.04025
R16990 VSS.n3487 VSS.n3403 0.04025
R16991 VSS.n3483 VSS.n3403 0.04025
R16992 VSS.n3483 VSS.n3482 0.04025
R16993 VSS.n3482 VSS.n3481 0.04025
R16994 VSS.n3481 VSS.n3405 0.04025
R16995 VSS.n3477 VSS.n3405 0.04025
R16996 VSS.n3477 VSS.n3476 0.04025
R16997 VSS.n3476 VSS.n3475 0.04025
R16998 VSS.n3475 VSS.n3407 0.04025
R16999 VSS.n3471 VSS.n3407 0.04025
R17000 VSS.n3471 VSS.n3470 0.04025
R17001 VSS.n3470 VSS.n3469 0.04025
R17002 VSS.n3469 VSS.n3409 0.04025
R17003 VSS.n3465 VSS.n3409 0.04025
R17004 VSS.n3465 VSS.n3464 0.04025
R17005 VSS.n3464 VSS.n3463 0.04025
R17006 VSS.n3463 VSS.n3411 0.04025
R17007 VSS.n3459 VSS.n3411 0.04025
R17008 VSS.n3459 VSS.n3458 0.04025
R17009 VSS.n3458 VSS.n3457 0.04025
R17010 VSS.n3457 VSS.n3413 0.04025
R17011 VSS.n3453 VSS.n3413 0.04025
R17012 VSS.n3453 VSS.n3452 0.04025
R17013 VSS.n3452 VSS.n3451 0.04025
R17014 VSS.n3451 VSS.n3415 0.04025
R17015 VSS.n3447 VSS.n3415 0.04025
R17016 VSS.n3447 VSS.n3446 0.04025
R17017 VSS.n3446 VSS.n3445 0.04025
R17018 VSS.n3445 VSS.n3417 0.04025
R17019 VSS.n3441 VSS.n3417 0.04025
R17020 VSS.n3441 VSS.n3440 0.04025
R17021 VSS.n3440 VSS.n3439 0.04025
R17022 VSS.n3439 VSS.n3419 0.04025
R17023 VSS.n3435 VSS.n3419 0.04025
R17024 VSS.n3435 VSS.n3434 0.04025
R17025 VSS.n3434 VSS.n3433 0.04025
R17026 VSS.n3433 VSS.n3421 0.04025
R17027 VSS.n3429 VSS.n3421 0.04025
R17028 VSS.n3429 VSS.n3428 0.04025
R17029 VSS.n3428 VSS.n3427 0.04025
R17030 VSS.n3427 VSS.n3423 0.04025
R17031 VSS.n3423 VSS.n1581 0.04025
R17032 VSS.n8951 VSS.n1581 0.04025
R17033 VSS.n8951 VSS.n8950 0.04025
R17034 VSS.n8950 VSS.n1583 0.04025
R17035 VSS.n8946 VSS.n1583 0.04025
R17036 VSS.n8946 VSS.n8945 0.04025
R17037 VSS.n8945 VSS.n8944 0.04025
R17038 VSS.n8944 VSS.n1585 0.04025
R17039 VSS.n8940 VSS.n1585 0.04025
R17040 VSS.n8940 VSS.n8939 0.04025
R17041 VSS.n8939 VSS.n8938 0.04025
R17042 VSS.n8938 VSS.n1587 0.04025
R17043 VSS.n8934 VSS.n1587 0.04025
R17044 VSS.n8934 VSS.n8933 0.04025
R17045 VSS.n8933 VSS.n8932 0.04025
R17046 VSS.n8932 VSS.n1589 0.04025
R17047 VSS.n8928 VSS.n1589 0.04025
R17048 VSS.n8928 VSS.n8927 0.04025
R17049 VSS.n8927 VSS.n8926 0.04025
R17050 VSS.n8926 VSS.n1591 0.04025
R17051 VSS.n8922 VSS.n1591 0.04025
R17052 VSS.n8922 VSS.n8921 0.04025
R17053 VSS.n8921 VSS.n8920 0.04025
R17054 VSS.n8920 VSS.n1593 0.04025
R17055 VSS.n8916 VSS.n1593 0.04025
R17056 VSS.n8916 VSS.n8915 0.04025
R17057 VSS.n8915 VSS.n8914 0.04025
R17058 VSS.n8914 VSS.n1595 0.04025
R17059 VSS.n8910 VSS.n1595 0.04025
R17060 VSS.n8910 VSS.n8909 0.04025
R17061 VSS.n8909 VSS.n8908 0.04025
R17062 VSS.n8908 VSS.n1597 0.04025
R17063 VSS.n8904 VSS.n1597 0.04025
R17064 VSS.n8904 VSS.n8903 0.04025
R17065 VSS.n8903 VSS.n8902 0.04025
R17066 VSS.n8902 VSS.n1599 0.04025
R17067 VSS.n8898 VSS.n1599 0.04025
R17068 VSS.n8898 VSS.n8897 0.04025
R17069 VSS.n8897 VSS.n8896 0.04025
R17070 VSS.n8896 VSS.n1601 0.04025
R17071 VSS.n8892 VSS.n1601 0.04025
R17072 VSS.n8892 VSS.n8891 0.04025
R17073 VSS.n8891 VSS.n8890 0.04025
R17074 VSS.n8890 VSS.n1603 0.04025
R17075 VSS.n8886 VSS.n1603 0.04025
R17076 VSS.n8886 VSS.n8885 0.04025
R17077 VSS.n8885 VSS.n8884 0.04025
R17078 VSS.n8884 VSS.n1605 0.04025
R17079 VSS.n8880 VSS.n1605 0.04025
R17080 VSS.n8880 VSS.n8879 0.04025
R17081 VSS.n8879 VSS.n8878 0.04025
R17082 VSS.n8878 VSS.n1607 0.04025
R17083 VSS.n8874 VSS.n1607 0.04025
R17084 VSS.n8874 VSS.n8873 0.04025
R17085 VSS.n8873 VSS.n8872 0.04025
R17086 VSS.n8872 VSS.n1609 0.04025
R17087 VSS.n8868 VSS.n1609 0.04025
R17088 VSS.n8868 VSS.n8867 0.04025
R17089 VSS.n8867 VSS.n8866 0.04025
R17090 VSS.n8866 VSS.n1611 0.04025
R17091 VSS.n8862 VSS.n1611 0.04025
R17092 VSS.n8862 VSS.n8861 0.04025
R17093 VSS.n8861 VSS.n8860 0.04025
R17094 VSS.n8860 VSS.n1613 0.04025
R17095 VSS.n8856 VSS.n1613 0.04025
R17096 VSS.n8856 VSS.n8855 0.04025
R17097 VSS.n8855 VSS.n8854 0.04025
R17098 VSS.n8854 VSS.n1615 0.04025
R17099 VSS.n8850 VSS.n1615 0.04025
R17100 VSS.n8850 VSS.n8849 0.04025
R17101 VSS.n8849 VSS.n8848 0.04025
R17102 VSS.n8848 VSS.n1617 0.04025
R17103 VSS.n8844 VSS.n1617 0.04025
R17104 VSS.n8844 VSS.n8843 0.04025
R17105 VSS.n8843 VSS.n8842 0.04025
R17106 VSS.n8842 VSS.n1619 0.04025
R17107 VSS.n8838 VSS.n1619 0.04025
R17108 VSS.n8838 VSS.n8837 0.04025
R17109 VSS.n8837 VSS.n8836 0.04025
R17110 VSS.n8836 VSS.n1621 0.04025
R17111 VSS.n8832 VSS.n1621 0.04025
R17112 VSS.n8832 VSS.n8831 0.04025
R17113 VSS.n8831 VSS.n8830 0.04025
R17114 VSS.n8830 VSS.n1623 0.04025
R17115 VSS.n8826 VSS.n1623 0.04025
R17116 VSS.n8826 VSS.n8825 0.04025
R17117 VSS.n8825 VSS.n8824 0.04025
R17118 VSS.n8824 VSS.n1625 0.04025
R17119 VSS.n8820 VSS.n1625 0.04025
R17120 VSS.n8820 VSS.n8819 0.04025
R17121 VSS.n8819 VSS.n8818 0.04025
R17122 VSS.n8818 VSS.n1627 0.04025
R17123 VSS.n8814 VSS.n1627 0.04025
R17124 VSS.n8814 VSS.n8813 0.04025
R17125 VSS.n8813 VSS.n8812 0.04025
R17126 VSS.n8812 VSS.n1629 0.04025
R17127 VSS.n8808 VSS.n1629 0.04025
R17128 VSS.n8808 VSS.n8807 0.04025
R17129 VSS.n8807 VSS.n8806 0.04025
R17130 VSS.n8806 VSS.n1631 0.04025
R17131 VSS.n8802 VSS.n1631 0.04025
R17132 VSS.n8802 VSS.n8801 0.04025
R17133 VSS.n8801 VSS.n8800 0.04025
R17134 VSS.n8800 VSS.n1633 0.04025
R17135 VSS.n8796 VSS.n1633 0.04025
R17136 VSS.n8796 VSS.n8795 0.04025
R17137 VSS.n8795 VSS.n8794 0.04025
R17138 VSS.n8794 VSS.n1635 0.04025
R17139 VSS.n8790 VSS.n1635 0.04025
R17140 VSS.n8790 VSS.n8789 0.04025
R17141 VSS.n8789 VSS.n8788 0.04025
R17142 VSS.n8788 VSS.n1637 0.04025
R17143 VSS.n8784 VSS.n1637 0.04025
R17144 VSS.n8784 VSS.n8783 0.04025
R17145 VSS.n8783 VSS.n8782 0.04025
R17146 VSS.n8782 VSS.n1639 0.04025
R17147 VSS.n8778 VSS.n1639 0.04025
R17148 VSS.n8778 VSS.n8777 0.04025
R17149 VSS.n8777 VSS.n8776 0.04025
R17150 VSS.n8776 VSS.n1641 0.04025
R17151 VSS.n8772 VSS.n1641 0.04025
R17152 VSS.n8772 VSS.n8771 0.04025
R17153 VSS.n8771 VSS.n8770 0.04025
R17154 VSS.n8770 VSS.n1643 0.04025
R17155 VSS.n8766 VSS.n1643 0.04025
R17156 VSS.n8766 VSS.n8765 0.04025
R17157 VSS.n8765 VSS.n8764 0.04025
R17158 VSS.n8764 VSS.n1645 0.04025
R17159 VSS.n8760 VSS.n1645 0.04025
R17160 VSS.n8760 VSS.n8759 0.04025
R17161 VSS.n8759 VSS.n8758 0.04025
R17162 VSS.n8758 VSS.n1647 0.04025
R17163 VSS.n8754 VSS.n1647 0.04025
R17164 VSS.n8754 VSS.n8753 0.04025
R17165 VSS.n8753 VSS.n8752 0.04025
R17166 VSS.n8752 VSS.n1649 0.04025
R17167 VSS.n8748 VSS.n1649 0.04025
R17168 VSS.n8748 VSS.n8747 0.04025
R17169 VSS.n8747 VSS.n8746 0.04025
R17170 VSS.n8746 VSS.n1651 0.04025
R17171 VSS.n8742 VSS.n1651 0.04025
R17172 VSS.n8742 VSS.n8741 0.04025
R17173 VSS.n8741 VSS.n8740 0.04025
R17174 VSS.n8740 VSS.n1653 0.04025
R17175 VSS.n8736 VSS.n1653 0.04025
R17176 VSS.n8736 VSS.n8735 0.04025
R17177 VSS.n8735 VSS.n8734 0.04025
R17178 VSS.n8734 VSS.n1655 0.04025
R17179 VSS.n8730 VSS.n1655 0.04025
R17180 VSS.n8730 VSS.n8729 0.04025
R17181 VSS.n8729 VSS.n8728 0.04025
R17182 VSS.n8728 VSS.n1657 0.04025
R17183 VSS.n8724 VSS.n1657 0.04025
R17184 VSS.n8724 VSS.n8723 0.04025
R17185 VSS.n8723 VSS.n8722 0.04025
R17186 VSS.n8722 VSS.n1659 0.04025
R17187 VSS.n8718 VSS.n1659 0.04025
R17188 VSS.n8718 VSS.n8717 0.04025
R17189 VSS.n8717 VSS.n8716 0.04025
R17190 VSS.n8716 VSS.n1661 0.04025
R17191 VSS.n8712 VSS.n1661 0.04025
R17192 VSS.n8712 VSS.n8711 0.04025
R17193 VSS.n8711 VSS.n8710 0.04025
R17194 VSS.n8710 VSS.n1663 0.04025
R17195 VSS.n8706 VSS.n1663 0.04025
R17196 VSS.n8706 VSS.n8705 0.04025
R17197 VSS.n8705 VSS.n8704 0.04025
R17198 VSS.n8704 VSS.n1665 0.04025
R17199 VSS.n8700 VSS.n1665 0.04025
R17200 VSS.n8700 VSS.n8699 0.04025
R17201 VSS.n8699 VSS.n8698 0.04025
R17202 VSS.n8698 VSS.n1667 0.04025
R17203 VSS.n8694 VSS.n1667 0.04025
R17204 VSS.n8694 VSS.n8693 0.04025
R17205 VSS.n8693 VSS.n8692 0.04025
R17206 VSS.n8692 VSS.n1669 0.04025
R17207 VSS.n8688 VSS.n1669 0.04025
R17208 VSS.n8688 VSS.n8687 0.04025
R17209 VSS.n8687 VSS.n8686 0.04025
R17210 VSS.n8686 VSS.n1671 0.04025
R17211 VSS.n8682 VSS.n1671 0.04025
R17212 VSS.n8682 VSS.n8681 0.04025
R17213 VSS.n8681 VSS.n8680 0.04025
R17214 VSS.n8680 VSS.n1673 0.04025
R17215 VSS.n8676 VSS.n1673 0.04025
R17216 VSS.n8676 VSS.n8675 0.04025
R17217 VSS.n8675 VSS.n8674 0.04025
R17218 VSS.n8674 VSS.n1675 0.04025
R17219 VSS.n8670 VSS.n1675 0.04025
R17220 VSS.n8670 VSS.n8669 0.04025
R17221 VSS.n8669 VSS.n8668 0.04025
R17222 VSS.n8668 VSS.n1677 0.04025
R17223 VSS.n8664 VSS.n1677 0.04025
R17224 VSS.n8664 VSS.n8663 0.04025
R17225 VSS.n8663 VSS.n8662 0.04025
R17226 VSS.n8662 VSS.n1679 0.04025
R17227 VSS.n8658 VSS.n1679 0.04025
R17228 VSS.n8658 VSS.n8657 0.04025
R17229 VSS.n8657 VSS.n8656 0.04025
R17230 VSS.n8656 VSS.n1681 0.04025
R17231 VSS.n8652 VSS.n1681 0.04025
R17232 VSS.n8652 VSS.n8651 0.04025
R17233 VSS.n8651 VSS.n8650 0.04025
R17234 VSS.n8650 VSS.n1683 0.04025
R17235 VSS.n8646 VSS.n1683 0.04025
R17236 VSS.n8646 VSS.n8645 0.04025
R17237 VSS.n8645 VSS.n8644 0.04025
R17238 VSS.n8644 VSS.n1685 0.04025
R17239 VSS.n8640 VSS.n1685 0.04025
R17240 VSS.n8640 VSS.n8639 0.04025
R17241 VSS.n8639 VSS.n8638 0.04025
R17242 VSS.n8638 VSS.n1687 0.04025
R17243 VSS.n8634 VSS.n1687 0.04025
R17244 VSS.n8634 VSS.n8633 0.04025
R17245 VSS.n8633 VSS.n8632 0.04025
R17246 VSS.n8632 VSS.n1689 0.04025
R17247 VSS.n8628 VSS.n1689 0.04025
R17248 VSS.n8628 VSS.n8627 0.04025
R17249 VSS.n8627 VSS.n8626 0.04025
R17250 VSS.n8626 VSS.n1691 0.04025
R17251 VSS.n8622 VSS.n1691 0.04025
R17252 VSS.n8622 VSS.n8621 0.04025
R17253 VSS.n8621 VSS.n8620 0.04025
R17254 VSS.n8620 VSS.n1693 0.04025
R17255 VSS.n8616 VSS.n1693 0.04025
R17256 VSS.n8616 VSS.n8615 0.04025
R17257 VSS.n8615 VSS.n8614 0.04025
R17258 VSS.n8614 VSS.n1695 0.04025
R17259 VSS.n8610 VSS.n1695 0.04025
R17260 VSS.n8610 VSS.n8609 0.04025
R17261 VSS.n8609 VSS.n8608 0.04025
R17262 VSS.n8608 VSS.n1697 0.04025
R17263 VSS.n8604 VSS.n1697 0.04025
R17264 VSS.n8604 VSS.n8603 0.04025
R17265 VSS.n8603 VSS.n8602 0.04025
R17266 VSS.n8602 VSS.n1699 0.04025
R17267 VSS.n8598 VSS.n1699 0.04025
R17268 VSS.n8598 VSS.n8597 0.04025
R17269 VSS.n8597 VSS.n8596 0.04025
R17270 VSS.n8596 VSS.n1701 0.04025
R17271 VSS.n8592 VSS.n1701 0.04025
R17272 VSS.n8592 VSS.n8591 0.04025
R17273 VSS.n8591 VSS.n8590 0.04025
R17274 VSS.n8590 VSS.n1703 0.04025
R17275 VSS.n8586 VSS.n1703 0.04025
R17276 VSS.n8586 VSS.n8585 0.04025
R17277 VSS.n8585 VSS.n8584 0.04025
R17278 VSS.n8584 VSS.n1705 0.04025
R17279 VSS.n8580 VSS.n1705 0.04025
R17280 VSS.n8580 VSS.n8579 0.04025
R17281 VSS.n8579 VSS.n8578 0.04025
R17282 VSS.n8578 VSS.n1707 0.04025
R17283 VSS.n8574 VSS.n1707 0.04025
R17284 VSS.n8574 VSS.n8573 0.04025
R17285 VSS.n8573 VSS.n8572 0.04025
R17286 VSS.n8572 VSS.n1709 0.04025
R17287 VSS.n8568 VSS.n1709 0.04025
R17288 VSS.n8568 VSS.n8567 0.04025
R17289 VSS.n8567 VSS.n8566 0.04025
R17290 VSS.n8566 VSS.n1711 0.04025
R17291 VSS.n8562 VSS.n1711 0.04025
R17292 VSS.n8562 VSS.n8561 0.04025
R17293 VSS.n8561 VSS.n8560 0.04025
R17294 VSS.n8560 VSS.n1713 0.04025
R17295 VSS.n8556 VSS.n1713 0.04025
R17296 VSS.n8556 VSS.n8555 0.04025
R17297 VSS.n8555 VSS.n8554 0.04025
R17298 VSS.n8554 VSS.n1715 0.04025
R17299 VSS.n8550 VSS.n1715 0.04025
R17300 VSS.n8550 VSS.n8549 0.04025
R17301 VSS.n8549 VSS.n8548 0.04025
R17302 VSS.n8548 VSS.n1717 0.04025
R17303 VSS.n8544 VSS.n1717 0.04025
R17304 VSS.n8544 VSS.n8543 0.04025
R17305 VSS.n8543 VSS.n8542 0.04025
R17306 VSS.n8542 VSS.n1719 0.04025
R17307 VSS.n8538 VSS.n1719 0.04025
R17308 VSS.n8538 VSS.n8537 0.04025
R17309 VSS.n8537 VSS.n8536 0.04025
R17310 VSS.n8536 VSS.n1721 0.04025
R17311 VSS.n8532 VSS.n1721 0.04025
R17312 VSS.n8532 VSS.n8531 0.04025
R17313 VSS.n8531 VSS.n8530 0.04025
R17314 VSS.n8530 VSS.n1723 0.04025
R17315 VSS.n8526 VSS.n1723 0.04025
R17316 VSS.n8526 VSS.n8525 0.04025
R17317 VSS.n8525 VSS.n8524 0.04025
R17318 VSS.n8524 VSS.n1725 0.04025
R17319 VSS.n8520 VSS.n1725 0.04025
R17320 VSS.n8520 VSS.n8519 0.04025
R17321 VSS.n8519 VSS.n8518 0.04025
R17322 VSS.n8518 VSS.n1727 0.04025
R17323 VSS.n8514 VSS.n1727 0.04025
R17324 VSS.n8514 VSS.n8513 0.04025
R17325 VSS.n8513 VSS.n8512 0.04025
R17326 VSS.n8512 VSS.n1729 0.04025
R17327 VSS.n8508 VSS.n1729 0.04025
R17328 VSS.n8508 VSS.n8507 0.04025
R17329 VSS.n8507 VSS.n8506 0.04025
R17330 VSS.n8506 VSS.n1731 0.04025
R17331 VSS.n8502 VSS.n1731 0.04025
R17332 VSS.n8502 VSS.n8501 0.04025
R17333 VSS.n8501 VSS.n8500 0.04025
R17334 VSS.n8500 VSS.n1733 0.04025
R17335 VSS.n8496 VSS.n1733 0.04025
R17336 VSS.n8496 VSS.n8495 0.04025
R17337 VSS.n8495 VSS.n8494 0.04025
R17338 VSS.n8494 VSS.n1735 0.04025
R17339 VSS.n8490 VSS.n1735 0.04025
R17340 VSS.n8490 VSS.n8489 0.04025
R17341 VSS.n8489 VSS.n8488 0.04025
R17342 VSS.n8488 VSS.n1737 0.04025
R17343 VSS.n8484 VSS.n1737 0.04025
R17344 VSS.n8484 VSS.n8483 0.04025
R17345 VSS.n8483 VSS.n8482 0.04025
R17346 VSS.n8482 VSS.n1739 0.04025
R17347 VSS.n8478 VSS.n1739 0.04025
R17348 VSS.n8478 VSS.n8477 0.04025
R17349 VSS.n8477 VSS.n8476 0.04025
R17350 VSS.n8476 VSS.n1741 0.04025
R17351 VSS.n8472 VSS.n1741 0.04025
R17352 VSS.n8472 VSS.n8471 0.04025
R17353 VSS.n8471 VSS.n8470 0.04025
R17354 VSS.n8470 VSS.n1743 0.04025
R17355 VSS.n8466 VSS.n1743 0.04025
R17356 VSS.n8466 VSS.n8465 0.04025
R17357 VSS.n8465 VSS.n8464 0.04025
R17358 VSS.n8464 VSS.n1745 0.04025
R17359 VSS.n8460 VSS.n1745 0.04025
R17360 VSS.n8460 VSS.n8459 0.04025
R17361 VSS.n8459 VSS.n8458 0.04025
R17362 VSS.n8458 VSS.n1747 0.04025
R17363 VSS.n8454 VSS.n1747 0.04025
R17364 VSS.n8454 VSS.n8453 0.04025
R17365 VSS.n8453 VSS.n8452 0.04025
R17366 VSS.n8452 VSS.n1749 0.04025
R17367 VSS.n8448 VSS.n1749 0.04025
R17368 VSS.n8448 VSS.n8447 0.04025
R17369 VSS.n8447 VSS.n8446 0.04025
R17370 VSS.n8446 VSS.n1751 0.04025
R17371 VSS.n8442 VSS.n1751 0.04025
R17372 VSS.n8442 VSS.n8441 0.04025
R17373 VSS.n8441 VSS.n8440 0.04025
R17374 VSS.n8440 VSS.n1753 0.04025
R17375 VSS.n8436 VSS.n1753 0.04025
R17376 VSS.n8436 VSS.n8435 0.04025
R17377 VSS.n8435 VSS.n8434 0.04025
R17378 VSS.n8434 VSS.n1755 0.04025
R17379 VSS.n8430 VSS.n1755 0.04025
R17380 VSS.n8430 VSS.n8429 0.04025
R17381 VSS.n8429 VSS.n8428 0.04025
R17382 VSS.n8428 VSS.n1757 0.04025
R17383 VSS.n8424 VSS.n1757 0.04025
R17384 VSS.n8424 VSS.n8423 0.04025
R17385 VSS.n8423 VSS.n8422 0.04025
R17386 VSS.n8422 VSS.n1759 0.04025
R17387 VSS.n8418 VSS.n1759 0.04025
R17388 VSS.n8418 VSS.n8417 0.04025
R17389 VSS.n8417 VSS.n8416 0.04025
R17390 VSS.n8416 VSS.n1761 0.04025
R17391 VSS.n8412 VSS.n1761 0.04025
R17392 VSS.n8412 VSS.n8411 0.04025
R17393 VSS.n8411 VSS.n8410 0.04025
R17394 VSS.n8410 VSS.n1763 0.04025
R17395 VSS.n8406 VSS.n1763 0.04025
R17396 VSS.n8406 VSS.n8405 0.04025
R17397 VSS.n8405 VSS.n8404 0.04025
R17398 VSS.n8404 VSS.n1765 0.04025
R17399 VSS.n8400 VSS.n1765 0.04025
R17400 VSS.n8400 VSS.n8399 0.04025
R17401 VSS.n8399 VSS.n8398 0.04025
R17402 VSS.n8398 VSS.n1767 0.04025
R17403 VSS.n8394 VSS.n1767 0.04025
R17404 VSS.n8394 VSS.n8393 0.04025
R17405 VSS.n8393 VSS.n8392 0.04025
R17406 VSS.n8392 VSS.n1769 0.04025
R17407 VSS.n8388 VSS.n1769 0.04025
R17408 VSS.n8388 VSS.n8387 0.04025
R17409 VSS.n8387 VSS.n8386 0.04025
R17410 VSS.n8386 VSS.n1771 0.04025
R17411 VSS.n8382 VSS.n1771 0.04025
R17412 VSS.n8382 VSS.n8381 0.04025
R17413 VSS.n8381 VSS.n8380 0.04025
R17414 VSS.n8380 VSS.n1773 0.04025
R17415 VSS.n8376 VSS.n1773 0.04025
R17416 VSS.n8376 VSS.n8375 0.04025
R17417 VSS.n8375 VSS.n8374 0.04025
R17418 VSS.n8374 VSS.n1775 0.04025
R17419 VSS.n8370 VSS.n1775 0.04025
R17420 VSS.n8370 VSS.n8369 0.04025
R17421 VSS.n8369 VSS.n8368 0.04025
R17422 VSS.n8368 VSS.n1777 0.04025
R17423 VSS.n8364 VSS.n1777 0.04025
R17424 VSS.n8364 VSS.n8363 0.04025
R17425 VSS.n8363 VSS.n8362 0.04025
R17426 VSS.n8362 VSS.n1779 0.04025
R17427 VSS.n8358 VSS.n1779 0.04025
R17428 VSS.n8358 VSS.n8357 0.04025
R17429 VSS.n8357 VSS.n8356 0.04025
R17430 VSS.n8356 VSS.n1781 0.04025
R17431 VSS.n8352 VSS.n1781 0.04025
R17432 VSS.n8352 VSS.n8351 0.04025
R17433 VSS.n8351 VSS.n8350 0.04025
R17434 VSS.n8350 VSS.n1783 0.04025
R17435 VSS.n8346 VSS.n1783 0.04025
R17436 VSS.n8346 VSS.n8345 0.04025
R17437 VSS.n8345 VSS.n8344 0.04025
R17438 VSS.n8344 VSS.n1785 0.04025
R17439 VSS.n8340 VSS.n1785 0.04025
R17440 VSS.n8340 VSS.n8339 0.04025
R17441 VSS.n8339 VSS.n8338 0.04025
R17442 VSS.n8338 VSS.n1787 0.04025
R17443 VSS.n8334 VSS.n1787 0.04025
R17444 VSS.n8334 VSS.n8333 0.04025
R17445 VSS.n8333 VSS.n8332 0.04025
R17446 VSS.n8332 VSS.n1789 0.04025
R17447 VSS.n8328 VSS.n1789 0.04025
R17448 VSS.n8328 VSS.n8327 0.04025
R17449 VSS.n8327 VSS.n8326 0.04025
R17450 VSS.n8326 VSS.n1791 0.04025
R17451 VSS.n8322 VSS.n1791 0.04025
R17452 VSS.n8322 VSS.n8321 0.04025
R17453 VSS.n8321 VSS.n8320 0.04025
R17454 VSS.n8320 VSS.n1793 0.04025
R17455 VSS.n8316 VSS.n1793 0.04025
R17456 VSS.n8316 VSS.n8315 0.04025
R17457 VSS.n8315 VSS.n8314 0.04025
R17458 VSS.n8314 VSS.n1795 0.04025
R17459 VSS.n8310 VSS.n1795 0.04025
R17460 VSS.n8310 VSS.n8309 0.04025
R17461 VSS.n8309 VSS.n8308 0.04025
R17462 VSS.n8308 VSS.n1797 0.04025
R17463 VSS.n8304 VSS.n1797 0.04025
R17464 VSS.n8304 VSS.n8303 0.04025
R17465 VSS.n8303 VSS.n8302 0.04025
R17466 VSS.n8302 VSS.n1799 0.04025
R17467 VSS.n8298 VSS.n1799 0.04025
R17468 VSS.n8298 VSS.n8297 0.04025
R17469 VSS.n8297 VSS.n8296 0.04025
R17470 VSS.n8296 VSS.n1801 0.04025
R17471 VSS.n8292 VSS.n1801 0.04025
R17472 VSS.n8292 VSS.n8291 0.04025
R17473 VSS.n8291 VSS.n8290 0.04025
R17474 VSS.n8290 VSS.n1803 0.04025
R17475 VSS.n8286 VSS.n1803 0.04025
R17476 VSS.n8286 VSS.n8285 0.04025
R17477 VSS.n8285 VSS.n8284 0.04025
R17478 VSS.n8284 VSS.n1805 0.04025
R17479 VSS.n8280 VSS.n1805 0.04025
R17480 VSS.n8280 VSS.n8279 0.04025
R17481 VSS.n8279 VSS.n8278 0.04025
R17482 VSS.n8278 VSS.n1807 0.04025
R17483 VSS.n8274 VSS.n1807 0.04025
R17484 VSS.n8274 VSS.n8273 0.04025
R17485 VSS.n8273 VSS.n8272 0.04025
R17486 VSS.n8272 VSS.n1809 0.04025
R17487 VSS.n8268 VSS.n1809 0.04025
R17488 VSS.n8268 VSS.n8267 0.04025
R17489 VSS.n8267 VSS.n8266 0.04025
R17490 VSS.n8266 VSS.n1811 0.04025
R17491 VSS.n8262 VSS.n1811 0.04025
R17492 VSS.n8262 VSS.n8261 0.04025
R17493 VSS.n8261 VSS.n8260 0.04025
R17494 VSS.n8260 VSS.n1813 0.04025
R17495 VSS.n8256 VSS.n1813 0.04025
R17496 VSS.n8256 VSS.n8255 0.04025
R17497 VSS.n8255 VSS.n8254 0.04025
R17498 VSS.n8254 VSS.n1815 0.04025
R17499 VSS.n8250 VSS.n1815 0.04025
R17500 VSS.n8250 VSS.n8249 0.04025
R17501 VSS.n8249 VSS.n8248 0.04025
R17502 VSS.n8248 VSS.n1817 0.04025
R17503 VSS.n8244 VSS.n1817 0.04025
R17504 VSS.n8244 VSS.n8243 0.04025
R17505 VSS.n8243 VSS.n8242 0.04025
R17506 VSS.n8242 VSS.n1819 0.04025
R17507 VSS.n8238 VSS.n1819 0.04025
R17508 VSS.n8238 VSS.n8237 0.04025
R17509 VSS.n8237 VSS.n8236 0.04025
R17510 VSS.n8236 VSS.n1821 0.04025
R17511 VSS.n8232 VSS.n1821 0.04025
R17512 VSS.n10642 VSS.n10641 0.039811
R17513 VSS.n11335 VSS.n11334 0.0390622
R17514 VSS.n77 VSS.n76 0.0390622
R17515 VSS.n11398 VSS.n0 0.0389239
R17516 VSS.n1575 VSS.n1573 0.0385696
R17517 VSS.n8962 VSS.n8961 0.0385696
R17518 VSS.n962 VSS.n961 0.0385696
R17519 VSS.n10280 VSS.n10279 0.0385696
R17520 VSS.n10454 VSS.n10453 0.0385295
R17521 VSS.n10476 VSS.n10475 0.0385295
R17522 VSS VSS.n0 0.0379215
R17523 VSS.n65 VSS.n63 0.0377578
R17524 VSS.n11333 VSS.n11332 0.0371211
R17525 VSS.n11328 VSS.n11327 0.0371211
R17526 VSS.n67 VSS.n66 0.0371211
R17527 VSS.n74 VSS.n73 0.0371211
R17528 VSS.n1577 VSS.n1576 0.0366533
R17529 VSS.n8959 VSS.n8958 0.0366533
R17530 VSS.n960 VSS.n959 0.0366533
R17531 VSS.n10282 VSS.n10281 0.0366533
R17532 VSS.n11326 VSS.n11325 0.0366035
R17533 VSS.n9434 VSS.n9433 0.0359944
R17534 VSS.n10868 VSS.n238 0.0359286
R17535 VSS.n11337 VSS.n111 0.0359286
R17536 VSS.n11399 VSS.n58 0.0359286
R17537 VSS.n10536 VSS.n10493 0.0359286
R17538 VSS VSS.n11470 0.0357042
R17539 VSS.n9448 VSS.n9447 0.035639
R17540 VSS.n10670 VSS.n10669 0.0354077
R17541 VSS.n10358 VSS.n10357 0.0354077
R17542 VSS.n10424 VSS.n10423 0.0354077
R17543 VSS.n10432 VSS.n10431 0.0354077
R17544 VSS.n10469 VSS.n10468 0.0353617
R17545 VSS.n10461 VSS.n10460 0.0353617
R17546 VSS.n10867 VSS.n239 0.0345
R17547 VSS.n11315 VSS.n106 0.0345
R17548 VSS.n11389 VSS.n11388 0.0345
R17549 VSS.n11394 VSS.n11393 0.0345
R17550 VSS.n11320 VSS.n11319 0.0345
R17551 VSS.n35 VSS.n34 0.0345
R17552 VSS.n10706 VSS.n10705 0.0345
R17553 VSS.n10529 VSS.n10499 0.0345
R17554 VSS.n11313 VSS.n11312 0.0345
R17555 VSS.n10566 VSS.n10565 0.0345
R17556 VSS.n10865 VSS.n225 0.0345
R17557 VSS.n10605 VSS.n10604 0.0342762
R17558 VSS.n10753 VSS.n10752 0.0342758
R17559 VSS.n8979 VSS.n8971 0.0341
R17560 VSS.n8977 VSS.n8971 0.0341
R17561 VSS.n8972 VSS.n1554 0.0341
R17562 VSS.n9096 VSS.n9095 0.0341
R17563 VSS.n9097 VSS.n9096 0.0341
R17564 VSS.n9097 VSS.n1553 0.0341
R17565 VSS.n9099 VSS.n1553 0.0341
R17566 VSS.n8966 VSS.n8965 0.0341
R17567 VSS.n8967 VSS.n8966 0.0341
R17568 VSS.n8967 VSS.n1565 0.0341
R17569 VSS.n8969 VSS.n1565 0.0341
R17570 VSS.n9007 VSS.n8970 0.0341
R17571 VSS.n9005 VSS.n8970 0.0341
R17572 VSS.n9005 VSS.n9004 0.0341
R17573 VSS.n9004 VSS.n9003 0.0341
R17574 VSS.n842 VSS.n838 0.0341
R17575 VSS.n840 VSS.n838 0.0341
R17576 VSS.n840 VSS.n839 0.0341
R17577 VSS.n839 VSS.n221 0.0341
R17578 VSS.n10926 VSS.n222 0.0341
R17579 VSS.n10924 VSS.n222 0.0341
R17580 VSS.n10924 VSS.n10923 0.0341
R17581 VSS.n10923 VSS.n10922 0.0341
R17582 VSS.n877 VSS.n836 0.0341
R17583 VSS.n875 VSS.n836 0.0341
R17584 VSS.n870 VSS.n869 0.0341
R17585 VSS.n866 VSS.n837 0.0341
R17586 VSS.n864 VSS.n837 0.0341
R17587 VSS.n864 VSS.n863 0.0341
R17588 VSS.n863 VSS.n862 0.0341
R17589 VSS.n1121 VSS.n1120 0.0341
R17590 VSS.n1122 VSS.n1121 0.0341
R17591 VSS.n1122 VSS.n879 0.0341
R17592 VSS.n1124 VSS.n879 0.0341
R17593 VSS.n1127 VSS.n1126 0.0341
R17594 VSS.n1128 VSS.n1127 0.0341
R17595 VSS.n1128 VSS.n878 0.0341
R17596 VSS.n1130 VSS.n878 0.0341
R17597 VSS.n1109 VSS.n1108 0.0341
R17598 VSS.n1110 VSS.n1109 0.0341
R17599 VSS.n1110 VSS.n902 0.0341
R17600 VSS.n1112 VSS.n902 0.0341
R17601 VSS.n1115 VSS.n1114 0.0341
R17602 VSS.n1116 VSS.n1115 0.0341
R17603 VSS.n1116 VSS.n901 0.0341
R17604 VSS.n1118 VSS.n901 0.0341
R17605 VSS.n1084 VSS.n1083 0.0341
R17606 VSS.n1089 VSS.n1084 0.0341
R17607 VSS.n1091 VSS.n904 0.0341
R17608 VSS.n1094 VSS.n1093 0.0341
R17609 VSS.n1095 VSS.n1094 0.0341
R17610 VSS.n1095 VSS.n903 0.0341
R17611 VSS.n1097 VSS.n903 0.0341
R17612 VSS.n1072 VSS.n1071 0.0341
R17613 VSS.n1073 VSS.n1072 0.0341
R17614 VSS.n1073 VSS.n915 0.0341
R17615 VSS.n1075 VSS.n915 0.0341
R17616 VSS.n1078 VSS.n1077 0.0341
R17617 VSS.n1079 VSS.n1078 0.0341
R17618 VSS.n1079 VSS.n914 0.0341
R17619 VSS.n1081 VSS.n914 0.0341
R17620 VSS.n1051 VSS.n1050 0.0341
R17621 VSS.n1052 VSS.n1051 0.0341
R17622 VSS.n1052 VSS.n917 0.0341
R17623 VSS.n1054 VSS.n917 0.0341
R17624 VSS.n1057 VSS.n1056 0.0341
R17625 VSS.n1058 VSS.n1057 0.0341
R17626 VSS.n1058 VSS.n916 0.0341
R17627 VSS.n1060 VSS.n916 0.0341
R17628 VSS.n1035 VSS.n1034 0.0341
R17629 VSS.n1040 VSS.n1035 0.0341
R17630 VSS.n1042 VSS.n928 0.0341
R17631 VSS.n1045 VSS.n1044 0.0341
R17632 VSS.n1046 VSS.n1045 0.0341
R17633 VSS.n1046 VSS.n927 0.0341
R17634 VSS.n1048 VSS.n927 0.0341
R17635 VSS.n1014 VSS.n1013 0.0341
R17636 VSS.n1015 VSS.n1014 0.0341
R17637 VSS.n1015 VSS.n930 0.0341
R17638 VSS.n1017 VSS.n930 0.0341
R17639 VSS.n1020 VSS.n1019 0.0341
R17640 VSS.n1021 VSS.n1020 0.0341
R17641 VSS.n1021 VSS.n929 0.0341
R17642 VSS.n1023 VSS.n929 0.0341
R17643 VSS.n1002 VSS.n1001 0.0341
R17644 VSS.n1003 VSS.n1002 0.0341
R17645 VSS.n1003 VSS.n941 0.0341
R17646 VSS.n1005 VSS.n941 0.0341
R17647 VSS.n1008 VSS.n1007 0.0341
R17648 VSS.n1009 VSS.n1008 0.0341
R17649 VSS.n1009 VSS.n940 0.0341
R17650 VSS.n1011 VSS.n940 0.0341
R17651 VSS.n977 VSS.n976 0.0341
R17652 VSS.n982 VSS.n977 0.0341
R17653 VSS.n984 VSS.n943 0.0341
R17654 VSS.n987 VSS.n986 0.0341
R17655 VSS.n988 VSS.n987 0.0341
R17656 VSS.n988 VSS.n942 0.0341
R17657 VSS.n990 VSS.n942 0.0341
R17658 VSS.n965 VSS.n964 0.0341
R17659 VSS.n966 VSS.n965 0.0341
R17660 VSS.n966 VSS.n954 0.0341
R17661 VSS.n968 VSS.n954 0.0341
R17662 VSS.n971 VSS.n970 0.0341
R17663 VSS.n972 VSS.n971 0.0341
R17664 VSS.n972 VSS.n953 0.0341
R17665 VSS.n974 VSS.n953 0.0341
R17666 VSS.n10920 VSS.n10916 0.0341
R17667 VSS.n10918 VSS.n10916 0.0341
R17668 VSS.n10918 VSS.n10917 0.0341
R17669 VSS.n10917 VSS.n207 0.0341
R17670 VSS.n10986 VSS.n10985 0.0341
R17671 VSS.n10987 VSS.n10986 0.0341
R17672 VSS.n10987 VSS.n206 0.0341
R17673 VSS.n10989 VSS.n206 0.0341
R17674 VSS.n10998 VSS.n10990 0.0341
R17675 VSS.n10996 VSS.n10990 0.0341
R17676 VSS.n10991 VSS.n96 0.0341
R17677 VSS.n11358 VSS.n97 0.0341
R17678 VSS.n11356 VSS.n97 0.0341
R17679 VSS.n11356 VSS.n11355 0.0341
R17680 VSS.n11355 VSS.n11354 0.0341
R17681 VSS.n11352 VSS.n101 0.0341
R17682 VSS.n11350 VSS.n101 0.0341
R17683 VSS.n11350 VSS.n11349 0.0341
R17684 VSS.n11349 VSS.n11348 0.0341
R17685 VSS.n11345 VSS.n102 0.0341
R17686 VSS.n11343 VSS.n102 0.0341
R17687 VSS.n11343 VSS.n11342 0.0341
R17688 VSS.n11342 VSS.n11341 0.0341
R17689 VSS.n11371 VSS.n11370 0.0341
R17690 VSS.n11372 VSS.n11371 0.0341
R17691 VSS.n11372 VSS.n85 0.0341
R17692 VSS.n11374 VSS.n85 0.0341
R17693 VSS.n11378 VSS.n11377 0.0341
R17694 VSS.n11379 VSS.n11378 0.0341
R17695 VSS.n11379 VSS.n84 0.0341
R17696 VSS.n11381 VSS.n84 0.0341
R17697 VSS.n10952 VSS.n10944 0.0341
R17698 VSS.n10950 VSS.n10944 0.0341
R17699 VSS.n10945 VSS.n90 0.0341
R17700 VSS.n11365 VSS.n11364 0.0341
R17701 VSS.n11366 VSS.n11365 0.0341
R17702 VSS.n11366 VSS.n89 0.0341
R17703 VSS.n11368 VSS.n89 0.0341
R17704 VSS.n10939 VSS.n10938 0.0341
R17705 VSS.n10940 VSS.n10939 0.0341
R17706 VSS.n10940 VSS.n209 0.0341
R17707 VSS.n10942 VSS.n209 0.0341
R17708 VSS.n10979 VSS.n10943 0.0341
R17709 VSS.n10977 VSS.n10943 0.0341
R17710 VSS.n10977 VSS.n10976 0.0341
R17711 VSS.n10976 VSS.n10975 0.0341
R17712 VSS.n1168 VSS.n1164 0.0341
R17713 VSS.n1166 VSS.n1164 0.0341
R17714 VSS.n1166 VSS.n1165 0.0341
R17715 VSS.n1165 VSS.n214 0.0341
R17716 VSS.n10933 VSS.n10932 0.0341
R17717 VSS.n10934 VSS.n10933 0.0341
R17718 VSS.n10934 VSS.n213 0.0341
R17719 VSS.n10936 VSS.n213 0.0341
R17720 VSS.n1214 VSS.n1162 0.0341
R17721 VSS.n1212 VSS.n1162 0.0341
R17722 VSS.n1207 VSS.n1206 0.0341
R17723 VSS.n1204 VSS.n1163 0.0341
R17724 VSS.n1202 VSS.n1163 0.0341
R17725 VSS.n1202 VSS.n1201 0.0341
R17726 VSS.n1201 VSS.n1200 0.0341
R17727 VSS.n9537 VSS.n9536 0.0341
R17728 VSS.n9538 VSS.n9537 0.0341
R17729 VSS.n9538 VSS.n1216 0.0341
R17730 VSS.n9540 VSS.n1216 0.0341
R17731 VSS.n9544 VSS.n9543 0.0341
R17732 VSS.n9545 VSS.n9544 0.0341
R17733 VSS.n9545 VSS.n1215 0.0341
R17734 VSS.n9547 VSS.n1215 0.0341
R17735 VSS.n1402 VSS.n1398 0.0341
R17736 VSS.n1400 VSS.n1398 0.0341
R17737 VSS.n1400 VSS.n1399 0.0341
R17738 VSS.n1399 VSS.n1221 0.0341
R17739 VSS.n9531 VSS.n9530 0.0341
R17740 VSS.n9532 VSS.n9531 0.0341
R17741 VSS.n9532 VSS.n1220 0.0341
R17742 VSS.n9534 VSS.n1220 0.0341
R17743 VSS.n1494 VSS.n1486 0.0341
R17744 VSS.n1492 VSS.n1486 0.0341
R17745 VSS.n1487 VSS.n1396 0.0341
R17746 VSS.n9419 VSS.n1397 0.0341
R17747 VSS.n9417 VSS.n1397 0.0341
R17748 VSS.n9417 VSS.n9416 0.0341
R17749 VSS.n9416 VSS.n9415 0.0341
R17750 VSS.n9268 VSS.n9264 0.0341
R17751 VSS.n9266 VSS.n9264 0.0341
R17752 VSS.n9266 VSS.n9265 0.0341
R17753 VSS.n9265 VSS.n1496 0.0341
R17754 VSS.n9351 VSS.n9350 0.0341
R17755 VSS.n9352 VSS.n9351 0.0341
R17756 VSS.n9352 VSS.n1495 0.0341
R17757 VSS.n9354 VSS.n1495 0.0341
R17758 VSS.n9259 VSS.n9258 0.0341
R17759 VSS.n9260 VSS.n9259 0.0341
R17760 VSS.n9260 VSS.n1508 0.0341
R17761 VSS.n9262 VSS.n1508 0.0341
R17762 VSS.n9296 VSS.n9263 0.0341
R17763 VSS.n9294 VSS.n9263 0.0341
R17764 VSS.n9294 VSS.n9293 0.0341
R17765 VSS.n9293 VSS.n9292 0.0341
R17766 VSS.n9146 VSS.n9138 0.0341
R17767 VSS.n9144 VSS.n9138 0.0341
R17768 VSS.n9139 VSS.n1513 0.0341
R17769 VSS.n9253 VSS.n9252 0.0341
R17770 VSS.n9254 VSS.n9253 0.0341
R17771 VSS.n9254 VSS.n1512 0.0341
R17772 VSS.n9256 VSS.n1512 0.0341
R17773 VSS.n9133 VSS.n9132 0.0341
R17774 VSS.n9134 VSS.n9133 0.0341
R17775 VSS.n9134 VSS.n1526 0.0341
R17776 VSS.n9136 VSS.n1526 0.0341
R17777 VSS.n9174 VSS.n9137 0.0341
R17778 VSS.n9172 VSS.n9137 0.0341
R17779 VSS.n9172 VSS.n9171 0.0341
R17780 VSS.n9171 VSS.n9170 0.0341
R17781 VSS.n1552 VSS.n1541 0.0341
R17782 VSS.n1550 VSS.n1541 0.0341
R17783 VSS.n1550 VSS.n1549 0.0341
R17784 VSS.n1549 VSS.n1548 0.0341
R17785 VSS.n1546 VSS.n1542 0.0341
R17786 VSS.n1544 VSS.n1542 0.0341
R17787 VSS.n1544 VSS.n1543 0.0341
R17788 VSS.n1543 VSS.n1527 0.0341
R17789 VSS.n11401 VSS.n11400 0.033821
R17790 VSS.n10676 VSS.n10336 0.0337454
R17791 VSS.n10674 VSS.n10336 0.0337454
R17792 VSS.n10674 VSS.n10673 0.0337454
R17793 VSS.n10673 VSS.n10672 0.0337454
R17794 VSS.n10672 VSS.n10337 0.0337454
R17795 VSS.n10670 VSS.n10337 0.0337454
R17796 VSS.n10669 VSS.n10338 0.0337454
R17797 VSS.n10667 VSS.n10338 0.0337454
R17798 VSS.n10667 VSS.n10666 0.0337454
R17799 VSS.n10355 VSS.n10339 0.0337454
R17800 VSS.n10357 VSS.n10355 0.0337454
R17801 VSS.n10358 VSS.n10354 0.0337454
R17802 VSS.n10360 VSS.n10354 0.0337454
R17803 VSS.n10361 VSS.n10360 0.0337454
R17804 VSS.n10362 VSS.n10361 0.0337454
R17805 VSS.n10362 VSS.n10353 0.0337454
R17806 VSS.n10364 VSS.n10353 0.0337454
R17807 VSS.n10417 VSS.n10291 0.0337454
R17808 VSS.n10419 VSS.n10417 0.0337454
R17809 VSS.n10420 VSS.n10419 0.0337454
R17810 VSS.n10421 VSS.n10420 0.0337454
R17811 VSS.n10421 VSS.n10416 0.0337454
R17812 VSS.n10423 VSS.n10416 0.0337454
R17813 VSS.n10424 VSS.n10415 0.0337454
R17814 VSS.n10426 VSS.n10415 0.0337454
R17815 VSS.n10427 VSS.n10426 0.0337454
R17816 VSS.n10429 VSS.n10414 0.0337454
R17817 VSS.n10431 VSS.n10414 0.0337454
R17818 VSS.n10432 VSS.n10413 0.0337454
R17819 VSS.n10434 VSS.n10413 0.0337454
R17820 VSS.n10435 VSS.n10434 0.0337454
R17821 VSS.n10436 VSS.n10435 0.0337454
R17822 VSS.n10436 VSS.n10412 0.0337454
R17823 VSS.n10438 VSS.n10412 0.0337454
R17824 VSS.n10475 VSS.n10443 0.0337016
R17825 VSS.n10473 VSS.n10443 0.0337016
R17826 VSS.n10473 VSS.n10472 0.0337016
R17827 VSS.n10472 VSS.n10471 0.0337016
R17828 VSS.n10471 VSS.n10444 0.0337016
R17829 VSS.n10469 VSS.n10444 0.0337016
R17830 VSS.n10468 VSS.n10445 0.0337016
R17831 VSS.n10466 VSS.n10445 0.0337016
R17832 VSS.n10466 VSS.n10465 0.0337016
R17833 VSS.n10463 VSS.n10446 0.0337016
R17834 VSS.n10461 VSS.n10446 0.0337016
R17835 VSS.n10460 VSS.n10447 0.0337016
R17836 VSS.n10458 VSS.n10447 0.0337016
R17837 VSS.n10458 VSS.n10457 0.0337016
R17838 VSS.n10457 VSS.n10456 0.0337016
R17839 VSS.n10456 VSS.n10448 0.0337016
R17840 VSS.n10454 VSS.n10448 0.0337016
R17841 VSS.n10665 VSS.n10339 0.033033
R17842 VSS.n10429 VSS.n10428 0.033033
R17843 VSS.n10464 VSS.n10463 0.0329901
R17844 VSS.n9486 VSS.n9485 0.0329468
R17845 VSS.n9484 VSS.n9483 0.0329468
R17846 VSS.n9482 VSS.n9481 0.0329468
R17847 VSS.n1410 VSS.n1409 0.0329468
R17848 VSS.n1412 VSS.n1411 0.0329468
R17849 VSS.n1414 VSS.n1413 0.0329468
R17850 VSS.n1321 VSS.n1320 0.0329468
R17851 VSS.n1323 VSS.n1322 0.0329468
R17852 VSS.n1325 VSS.n1324 0.0329468
R17853 VSS.n9509 VSS.n9508 0.0329468
R17854 VSS.n10819 VSS.n10818 0.032073
R17855 VSS.n10777 VSS.n10776 0.032073
R17856 VSS.n10788 VSS.n10787 0.032073
R17857 VSS.n9485 VSS.n9477 0.0319894
R17858 VSS.n9484 VSS.n9477 0.0319894
R17859 VSS.n9483 VSS.n9478 0.0319894
R17860 VSS.n9482 VSS.n9478 0.0319894
R17861 VSS.n9481 VSS.n9479 0.0319894
R17862 VSS.n9480 VSS.n9479 0.0319894
R17863 VSS.n1386 VSS.n1385 0.0319894
R17864 VSS.n1408 VSS.n1407 0.0319894
R17865 VSS.n1409 VSS.n1407 0.0319894
R17866 VSS.n1410 VSS.n1406 0.0319894
R17867 VSS.n1411 VSS.n1406 0.0319894
R17868 VSS.n1412 VSS.n1405 0.0319894
R17869 VSS.n1413 VSS.n1405 0.0319894
R17870 VSS.n1414 VSS.n1404 0.0319894
R17871 VSS.n1415 VSS.n1404 0.0319894
R17872 VSS.n1319 VSS.n1271 0.0319894
R17873 VSS.n1320 VSS.n1271 0.0319894
R17874 VSS.n1321 VSS.n1270 0.0319894
R17875 VSS.n1322 VSS.n1270 0.0319894
R17876 VSS.n1323 VSS.n1269 0.0319894
R17877 VSS.n1324 VSS.n1269 0.0319894
R17878 VSS.n1325 VSS.n1268 0.0319894
R17879 VSS.n1326 VSS.n1268 0.0319894
R17880 VSS.n1332 VSS.n1331 0.0319894
R17881 VSS.n9510 VSS.n1334 0.0319894
R17882 VSS.n9509 VSS.n1334 0.0319894
R17883 VSS.n10752 VSS.n10747 0.0319607
R17884 VSS.n10750 VSS.n10747 0.0319607
R17885 VSS.n10750 VSS.n10749 0.0319607
R17886 VSS.n10749 VSS.n10748 0.0319607
R17887 VSS.n10815 VSS.n10814 0.0319607
R17888 VSS.n10816 VSS.n10815 0.0319607
R17889 VSS.n10816 VSS.n10813 0.0319607
R17890 VSS.n10818 VSS.n10813 0.0319607
R17891 VSS.n10778 VSS.n10777 0.0319607
R17892 VSS.n10779 VSS.n10778 0.0319607
R17893 VSS.n10779 VSS.n10737 0.0319607
R17894 VSS.n10781 VSS.n10737 0.0319607
R17895 VSS.n10784 VSS.n10783 0.0319607
R17896 VSS.n10785 VSS.n10784 0.0319607
R17897 VSS.n10785 VSS.n10736 0.0319607
R17898 VSS.n10787 VSS.n10736 0.0319607
R17899 VSS.n10494 VSS.n10441 0.0319161
R17900 VSS.n10582 VSS.n10581 0.0315563
R17901 VSS.n10649 VSS.n10648 0.0315563
R17902 VSS.n10453 VSS.n10452 0.0314767
R17903 VSS.n10451 VSS.n10450 0.0314767
R17904 VSS.n10449 VSS.n10345 0.0314767
R17905 VSS.n10659 VSS.n10658 0.0314767
R17906 VSS.n10657 VSS.n10656 0.0314767
R17907 VSS.n10477 VSS.n10476 0.0314767
R17908 VSS.n10479 VSS.n10478 0.0314767
R17909 VSS.n10481 VSS.n10480 0.0314767
R17910 VSS.n10596 VSS.n10595 0.0314767
R17911 VSS.n10594 VSS.n10593 0.0314767
R17912 VSS.n10560 VSS.n10559 0.0314767
R17913 VSS.n10558 VSS.n10290 0.0314767
R17914 VSS.n10693 VSS.n10692 0.0314767
R17915 VSS.n10691 VSS.n10690 0.0314767
R17916 VSS.n10689 VSS.n10688 0.0314767
R17917 VSS.n10641 VSS.n10640 0.0314767
R17918 VSS.n10572 VSS.n10561 0.0313721
R17919 VSS.n1388 VSS.n1387 0.0311383
R17920 VSS.n1333 VSS.n1330 0.0311383
R17921 VSS.n11331 VSS.n11330 0.0301981
R17922 VSS.n72 VSS.n70 0.0301981
R17923 VSS.n10575 VSS.n10574 0.0301831
R17924 VSS.n10278 VSS.n10277 0.0301505
R17925 VSS.n1572 VSS.n1570 0.0300866
R17926 VSS.n10575 VSS.n10555 0.0300775
R17927 VSS.n10577 VSS.n10555 0.0300775
R17928 VSS.n10578 VSS.n10577 0.0300775
R17929 VSS.n10579 VSS.n10578 0.0300775
R17930 VSS.n10579 VSS.n10554 0.0300775
R17931 VSS.n10581 VSS.n10554 0.0300775
R17932 VSS.n10582 VSS.n10553 0.0300775
R17933 VSS.n10584 VSS.n10553 0.0300775
R17934 VSS.n10585 VSS.n10584 0.0300775
R17935 VSS.n10651 VSS.n10650 0.0300775
R17936 VSS.n10650 VSS.n10649 0.0300775
R17937 VSS.n10648 VSS.n10350 0.0300775
R17938 VSS.n10646 VSS.n10350 0.0300775
R17939 VSS.n10646 VSS.n10645 0.0300775
R17940 VSS.n10645 VSS.n10644 0.0300775
R17941 VSS.n10644 VSS.n10351 0.0300775
R17942 VSS.n10642 VSS.n10351 0.0300775
R17943 VSS.n8965 VSS.n8964 0.0299989
R17944 VSS.n964 VSS.n963 0.0299989
R17945 VSS.n8957 VSS.n8955 0.0298187
R17946 VSS.n9073 VSS.n9046 0.0294988
R17947 VSS.n9071 VSS.n9046 0.0294988
R17948 VSS.n9071 VSS.n9070 0.0294988
R17949 VSS.n9070 VSS.n9069 0.0294988
R17950 VSS.n9067 VSS.n9047 0.0294988
R17951 VSS.n9065 VSS.n9047 0.0294988
R17952 VSS.n9065 VSS.n9064 0.0294988
R17953 VSS.n9064 VSS.n9063 0.0294988
R17954 VSS.n9041 VSS.n9040 0.0294988
R17955 VSS.n9042 VSS.n9041 0.0294988
R17956 VSS.n9042 VSS.n1556 0.0294988
R17957 VSS.n9044 VSS.n1556 0.0294988
R17958 VSS.n9088 VSS.n9045 0.0294988
R17959 VSS.n9086 VSS.n9045 0.0294988
R17960 VSS.n9086 VSS.n9085 0.0294988
R17961 VSS.n9085 VSS.n9084 0.0294988
R17962 VSS.n1570 VSS.n1566 0.0294988
R17963 VSS.n1568 VSS.n1566 0.0294988
R17964 VSS.n1568 VSS.n1567 0.0294988
R17965 VSS.n1567 VSS.n1561 0.0294988
R17966 VSS.n9017 VSS.n9016 0.0294988
R17967 VSS.n9036 VSS.n9017 0.0294988
R17968 VSS.n9036 VSS.n9035 0.0294988
R17969 VSS.n1285 VSS.n416 0.0294988
R17970 VSS.n1286 VSS.n1285 0.0294988
R17971 VSS.n1286 VSS.n1284 0.0294988
R17972 VSS.n1288 VSS.n1284 0.0294988
R17973 VSS.n1291 VSS.n1290 0.0294988
R17974 VSS.n1292 VSS.n1291 0.0294988
R17975 VSS.n1292 VSS.n1283 0.0294988
R17976 VSS.n1294 VSS.n1283 0.0294988
R17977 VSS.n10157 VSS.n401 0.0294988
R17978 VSS.n10155 VSS.n401 0.0294988
R17979 VSS.n10155 VSS.n10154 0.0294988
R17980 VSS.n10154 VSS.n10153 0.0294988
R17981 VSS.n10151 VSS.n402 0.0294988
R17982 VSS.n10149 VSS.n402 0.0294988
R17983 VSS.n10149 VSS.n10148 0.0294988
R17984 VSS.n387 VSS.n386 0.0294988
R17985 VSS.n388 VSS.n387 0.0294988
R17986 VSS.n388 VSS.n363 0.0294988
R17987 VSS.n390 VSS.n363 0.0294988
R17988 VSS.n10160 VSS.n10159 0.0294988
R17989 VSS.n10161 VSS.n10160 0.0294988
R17990 VSS.n10161 VSS.n10158 0.0294988
R17991 VSS.n10163 VSS.n10158 0.0294988
R17992 VSS.n366 VSS.n344 0.0294988
R17993 VSS.n367 VSS.n366 0.0294988
R17994 VSS.n367 VSS.n365 0.0294988
R17995 VSS.n369 VSS.n365 0.0294988
R17996 VSS.n372 VSS.n371 0.0294988
R17997 VSS.n373 VSS.n372 0.0294988
R17998 VSS.n373 VSS.n364 0.0294988
R17999 VSS.n375 VSS.n364 0.0294988
R18000 VSS.n10217 VSS.n329 0.0294988
R18001 VSS.n10215 VSS.n329 0.0294988
R18002 VSS.n10215 VSS.n10214 0.0294988
R18003 VSS.n10214 VSS.n10213 0.0294988
R18004 VSS.n10211 VSS.n330 0.0294988
R18005 VSS.n10209 VSS.n330 0.0294988
R18006 VSS.n10209 VSS.n10208 0.0294988
R18007 VSS.n315 VSS.n314 0.0294988
R18008 VSS.n316 VSS.n315 0.0294988
R18009 VSS.n316 VSS.n291 0.0294988
R18010 VSS.n318 VSS.n291 0.0294988
R18011 VSS.n10220 VSS.n10219 0.0294988
R18012 VSS.n10221 VSS.n10220 0.0294988
R18013 VSS.n10221 VSS.n10218 0.0294988
R18014 VSS.n10223 VSS.n10218 0.0294988
R18015 VSS.n303 VSS.n272 0.0294988
R18016 VSS.n304 VSS.n303 0.0294988
R18017 VSS.n304 VSS.n302 0.0294988
R18018 VSS.n306 VSS.n302 0.0294988
R18019 VSS.n309 VSS.n308 0.0294988
R18020 VSS.n310 VSS.n309 0.0294988
R18021 VSS.n310 VSS.n301 0.0294988
R18022 VSS.n312 VSS.n301 0.0294988
R18023 VSS.n10277 VSS.n257 0.0294988
R18024 VSS.n10275 VSS.n257 0.0294988
R18025 VSS.n10275 VSS.n10274 0.0294988
R18026 VSS.n10274 VSS.n10273 0.0294988
R18027 VSS.n10271 VSS.n258 0.0294988
R18028 VSS.n10269 VSS.n258 0.0294988
R18029 VSS.n10269 VSS.n10268 0.0294988
R18030 VSS.n9377 VSS.n9376 0.0294988
R18031 VSS.n9378 VSS.n9377 0.0294988
R18032 VSS.n9378 VSS.n1477 0.0294988
R18033 VSS.n9380 VSS.n1477 0.0294988
R18034 VSS.n9384 VSS.n9383 0.0294988
R18035 VSS.n9385 VSS.n9384 0.0294988
R18036 VSS.n9385 VSS.n1476 0.0294988
R18037 VSS.n9387 VSS.n1476 0.0294988
R18038 VSS.n9317 VSS.n9316 0.0294988
R18039 VSS.n9318 VSS.n9317 0.0294988
R18040 VSS.n9318 VSS.n1500 0.0294988
R18041 VSS.n9320 VSS.n1500 0.0294988
R18042 VSS.n9343 VSS.n9321 0.0294988
R18043 VSS.n9341 VSS.n9321 0.0294988
R18044 VSS.n9341 VSS.n9340 0.0294988
R18045 VSS.n9217 VSS.n9213 0.0294988
R18046 VSS.n9215 VSS.n9213 0.0294988
R18047 VSS.n9215 VSS.n9214 0.0294988
R18048 VSS.n9214 VSS.n1505 0.0294988
R18049 VSS.n9311 VSS.n9310 0.0294988
R18050 VSS.n9312 VSS.n9311 0.0294988
R18051 VSS.n9312 VSS.n1504 0.0294988
R18052 VSS.n9314 VSS.n1504 0.0294988
R18053 VSS.n9208 VSS.n9207 0.0294988
R18054 VSS.n9209 VSS.n9208 0.0294988
R18055 VSS.n9209 VSS.n1518 0.0294988
R18056 VSS.n9211 VSS.n1518 0.0294988
R18057 VSS.n9245 VSS.n9212 0.0294988
R18058 VSS.n9243 VSS.n9212 0.0294988
R18059 VSS.n9243 VSS.n9242 0.0294988
R18060 VSS.n9242 VSS.n9241 0.0294988
R18061 VSS.n9061 VSS.n9057 0.0294988
R18062 VSS.n9059 VSS.n9057 0.0294988
R18063 VSS.n9059 VSS.n9058 0.0294988
R18064 VSS.n9058 VSS.n1523 0.0294988
R18065 VSS.n9184 VSS.n9183 0.0294988
R18066 VSS.n9203 VSS.n9184 0.0294988
R18067 VSS.n9203 VSS.n9202 0.0294988
R18068 VSS.n10825 VSS.n10821 0.029033
R18069 VSS.n9487 VSS.n9486 0.0286128
R18070 VSS.n10769 VSS.n10768 0.0280818
R18071 VSS.n10634 VSS.n10352 0.0277138
R18072 VSS.n9002 VSS.n8979 0.02738
R18073 VSS.n9100 VSS.n9099 0.02738
R18074 VSS.n9003 VSS.n9002 0.02738
R18075 VSS.n861 VSS.n842 0.02738
R18076 VSS.n10922 VSS.n10921 0.02738
R18077 VSS.n1131 VSS.n877 0.02738
R18078 VSS.n862 VSS.n861 0.02738
R18079 VSS.n1120 VSS.n1119 0.02738
R18080 VSS.n1131 VSS.n1130 0.02738
R18081 VSS.n1108 VSS.n1107 0.02738
R18082 VSS.n1119 VSS.n1118 0.02738
R18083 VSS.n1083 VSS.n1082 0.02738
R18084 VSS.n1107 VSS.n1097 0.02738
R18085 VSS.n1071 VSS.n1070 0.02738
R18086 VSS.n1082 VSS.n1081 0.02738
R18087 VSS.n1050 VSS.n1049 0.02738
R18088 VSS.n1070 VSS.n1060 0.02738
R18089 VSS.n1034 VSS.n1033 0.02738
R18090 VSS.n1049 VSS.n1048 0.02738
R18091 VSS.n1013 VSS.n1012 0.02738
R18092 VSS.n1033 VSS.n1023 0.02738
R18093 VSS.n1001 VSS.n1000 0.02738
R18094 VSS.n1012 VSS.n1011 0.02738
R18095 VSS.n976 VSS.n975 0.02738
R18096 VSS.n1000 VSS.n990 0.02738
R18097 VSS.n975 VSS.n974 0.02738
R18098 VSS.n10921 VSS.n10920 0.02738
R18099 VSS.n10999 VSS.n10989 0.02738
R18100 VSS.n10999 VSS.n10998 0.02738
R18101 VSS.n11354 VSS.n11353 0.02738
R18102 VSS.n11353 VSS.n11352 0.02738
R18103 VSS.n11341 VSS.n11340 0.02738
R18104 VSS.n11370 VSS.n11369 0.02738
R18105 VSS.n11382 VSS.n11381 0.02738
R18106 VSS.n10974 VSS.n10952 0.02738
R18107 VSS.n11369 VSS.n11368 0.02738
R18108 VSS.n10938 VSS.n10937 0.02738
R18109 VSS.n10975 VSS.n10974 0.02738
R18110 VSS.n1199 VSS.n1168 0.02738
R18111 VSS.n10937 VSS.n10936 0.02738
R18112 VSS.n9548 VSS.n1214 0.02738
R18113 VSS.n1200 VSS.n1199 0.02738
R18114 VSS.n9536 VSS.n9535 0.02738
R18115 VSS.n9548 VSS.n9547 0.02738
R18116 VSS.n9414 VSS.n1402 0.02738
R18117 VSS.n9535 VSS.n9534 0.02738
R18118 VSS.n9355 VSS.n1494 0.02738
R18119 VSS.n9415 VSS.n9414 0.02738
R18120 VSS.n9291 VSS.n9268 0.02738
R18121 VSS.n9355 VSS.n9354 0.02738
R18122 VSS.n9258 VSS.n9257 0.02738
R18123 VSS.n9292 VSS.n9291 0.02738
R18124 VSS.n9169 VSS.n9146 0.02738
R18125 VSS.n9257 VSS.n9256 0.02738
R18126 VSS.n9132 VSS.n9131 0.02738
R18127 VSS.n9170 VSS.n9169 0.02738
R18128 VSS.n9100 VSS.n1552 0.02738
R18129 VSS.n9131 VSS.n1527 0.02738
R18130 VSS.n10633 VSS.n10364 0.0271502
R18131 VSS.n10842 VSS.n10841 0.0261855
R18132 VSS.n10763 VSS.n10762 0.0259315
R18133 VSS.n10746 VSS.n10745 0.0255699
R18134 VSS.n9198 VSS.n9186 0.0255051
R18135 VSS.n9335 VSS.n9334 0.0255051
R18136 VSS.n172 VSS.n160 0.0255051
R18137 VSS.n9582 VSS.n9580 0.0255051
R18138 VSS.n11140 VSS.n200 0.0255051
R18139 VSS.n482 VSS.n481 0.0255051
R18140 VSS.n9031 VSS.n9019 0.0255051
R18141 VSS.n10263 VSS.n271 0.0255051
R18142 VSS.n10203 VSS.n343 0.0255051
R18143 VSS.n10143 VSS.n415 0.0255051
R18144 VSS.n10823 VSS.n10822 0.024829
R18145 VSS.n9083 VSS.n9073 0.0236991
R18146 VSS.n9063 VSS.n9062 0.0236991
R18147 VSS.n9040 VSS.n9039 0.0236991
R18148 VSS.n9084 VSS.n9083 0.0236991
R18149 VSS.n9039 VSS.n9038 0.0236991
R18150 VSS.n10141 VSS.n416 0.0236991
R18151 VSS.n1295 VSS.n1294 0.0236991
R18152 VSS.n10164 VSS.n10157 0.0236991
R18153 VSS.n10142 VSS.n10141 0.0236991
R18154 VSS.n386 VSS.n385 0.0236991
R18155 VSS.n10164 VSS.n10163 0.0236991
R18156 VSS.n10201 VSS.n344 0.0236991
R18157 VSS.n385 VSS.n375 0.0236991
R18158 VSS.n10224 VSS.n10217 0.0236991
R18159 VSS.n10202 VSS.n10201 0.0236991
R18160 VSS.n314 VSS.n313 0.0236991
R18161 VSS.n10224 VSS.n10223 0.0236991
R18162 VSS.n10261 VSS.n272 0.0236991
R18163 VSS.n313 VSS.n312 0.0236991
R18164 VSS.n10262 VSS.n10261 0.0236991
R18165 VSS.n9376 VSS.n9375 0.0236991
R18166 VSS.n9388 VSS.n9387 0.0236991
R18167 VSS.n9316 VSS.n9315 0.0236991
R18168 VSS.n9375 VSS.n1478 0.0236991
R18169 VSS.n9240 VSS.n9217 0.0236991
R18170 VSS.n9315 VSS.n9314 0.0236991
R18171 VSS.n9207 VSS.n9206 0.0236991
R18172 VSS.n9241 VSS.n9240 0.0236991
R18173 VSS.n9062 VSS.n9061 0.0236991
R18174 VSS.n9206 VSS.n9205 0.0236991
R18175 VSS.n10651 VSS.n10349 0.0231186
R18176 VSS.n6936 VSS.n61 0.023
R18177 VSS.n10843 VSS.n10733 0.0229499
R18178 VSS.n8977 VSS.n8976 0.022805
R18179 VSS.n875 VSS.n874 0.022805
R18180 VSS.n1089 VSS.n1088 0.022805
R18181 VSS.n1040 VSS.n1039 0.022805
R18182 VSS.n982 VSS.n981 0.022805
R18183 VSS.n10996 VSS.n10995 0.022805
R18184 VSS.n10950 VSS.n10949 0.022805
R18185 VSS.n1212 VSS.n1211 0.022805
R18186 VSS.n1492 VSS.n1491 0.022805
R18187 VSS.n9144 VSS.n9143 0.022805
R18188 VSS.n10639 VSS.n10638 0.0217442
R18189 VSS.n9200 VSS.n9198 0.0215309
R18190 VSS.n9338 VSS.n9334 0.0215309
R18191 VSS.n175 VSS.n172 0.0215309
R18192 VSS.n9585 VSS.n9580 0.0215309
R18193 VSS.n11143 VSS.n200 0.0215309
R18194 VSS.n481 VSS.n480 0.0215309
R18195 VSS.n9033 VSS.n9031 0.0215309
R18196 VSS.n10266 VSS.n271 0.0215309
R18197 VSS.n10206 VSS.n343 0.0215309
R18198 VSS.n10146 VSS.n415 0.0215309
R18199 VSS.n10688 VSS.n10687 0.0213083
R18200 VSS.n10496 VSS.n10495 0.0209545
R18201 VSS.n10607 VSS.n10606 0.0208496
R18202 VSS.n9752 VSS.n9649 0.0206923
R18203 VSS.n9864 VSS.n178 0.0206923
R18204 VSS.n1260 VSS.n455 0.0206923
R18205 VSS.n634 VSS.n499 0.0206923
R18206 VSS.n10015 VSS.n9934 0.0206923
R18207 VSS.n9993 VSS.n9954 0.0206923
R18208 VSS.n11195 VSS.n11194 0.0206923
R18209 VSS.n9626 VSS.n9625 0.0206923
R18210 VSS.n10677 VSS.n10676 0.0206172
R18211 VSS.n10687 VSS.n10291 0.0206172
R18212 VSS.n786 VSS.n785 0.0205874
R18213 VSS.n9730 VSS.n9693 0.0205874
R18214 VSS.n9842 VSS.n9841 0.0205874
R18215 VSS.n10015 VSS.n578 0.0205874
R18216 VSS.n9626 VSS.n804 0.0205874
R18217 VSS.n9752 VSS.n9661 0.0205874
R18218 VSS.n10048 VSS.n546 0.0205874
R18219 VSS.n9730 VSS.n9717 0.0205874
R18220 VSS.n590 VSS.n184 0.0205874
R18221 VSS.n11051 VSS.n11050 0.0205874
R18222 VSS.n9993 VSS.n9966 0.0205874
R18223 VSS.n9602 VSS.n9601 0.0205874
R18224 VSS.n10439 VSS.n10438 0.0204409
R18225 VSS.n11330 VSS.n11329 0.0203634
R18226 VSS.n70 VSS.n69 0.0203634
R18227 VSS.n10284 VSS.n10283 0.0201097
R18228 VSS.n9095 VSS.n9094 0.01994
R18229 VSS.n9008 VSS.n9007 0.01994
R18230 VSS.n10927 VSS.n10926 0.01994
R18231 VSS.n868 VSS.n866 0.01994
R18232 VSS.n1126 VSS.n1125 0.01994
R18233 VSS.n1114 VSS.n1113 0.01994
R18234 VSS.n1093 VSS.n1092 0.01994
R18235 VSS.n1077 VSS.n1076 0.01994
R18236 VSS.n1056 VSS.n1055 0.01994
R18237 VSS.n1044 VSS.n1043 0.01994
R18238 VSS.n1019 VSS.n1018 0.01994
R18239 VSS.n1007 VSS.n1006 0.01994
R18240 VSS.n986 VSS.n985 0.01994
R18241 VSS.n970 VSS.n969 0.01994
R18242 VSS.n10985 VSS.n10984 0.01994
R18243 VSS.n11359 VSS.n11358 0.01994
R18244 VSS.n11347 VSS.n11345 0.01994
R18245 VSS.n11377 VSS.n11376 0.01994
R18246 VSS.n11364 VSS.n11363 0.01994
R18247 VSS.n10980 VSS.n10979 0.01994
R18248 VSS.n10932 VSS.n10931 0.01994
R18249 VSS.n1205 VSS.n1204 0.01994
R18250 VSS.n9543 VSS.n9542 0.01994
R18251 VSS.n9530 VSS.n9529 0.01994
R18252 VSS.n9420 VSS.n9419 0.01994
R18253 VSS.n9350 VSS.n9349 0.01994
R18254 VSS.n9297 VSS.n9296 0.01994
R18255 VSS.n9252 VSS.n9251 0.01994
R18256 VSS.n9175 VSS.n9174 0.01994
R18257 VSS.n1547 VSS.n1546 0.01994
R18258 VSS.n11334 VSS.n11333 0.0196517
R18259 VSS.n11332 VSS.n11331 0.0196517
R18260 VSS.n11329 VSS.n11328 0.0196517
R18261 VSS.n11327 VSS.n11326 0.0196517
R18262 VSS.n66 VSS.n65 0.0196517
R18263 VSS.n69 VSS.n67 0.0196517
R18264 VSS.n73 VSS.n72 0.0196517
R18265 VSS.n76 VSS.n74 0.0196517
R18266 VSS.n9080 VSS.n9079 0.0194273
R18267 VSS.n9105 VSS.n9103 0.0194273
R18268 VSS.n858 VSS.n857 0.0194273
R18269 VSS.n1104 VSS.n1103 0.0194273
R18270 VSS.n1279 VSS.n1278 0.0194273
R18271 VSS.n924 VSS.n923 0.0194273
R18272 VSS.n381 VSS.n380 0.0194273
R18273 VSS.n997 VSS.n996 0.0194273
R18274 VSS.n297 VSS.n296 0.0194273
R18275 VSS.n11063 VSS.n11060 0.0194273
R18276 VSS.n11211 VSS.n11209 0.0194273
R18277 VSS.n1195 VSS.n1194 0.0194273
R18278 VSS.n9395 VSS.n9392 0.0194273
R18279 VSS.n9410 VSS.n9409 0.0194273
R18280 VSS.n9237 VSS.n9236 0.0194273
R18281 VSS.n9225 VSS.n9223 0.0194273
R18282 VSS.n1573 VSS.n1572 0.019407
R18283 VSS.n1576 VSS.n1575 0.019407
R18284 VSS.n1579 VSS.n1577 0.019407
R18285 VSS.n8958 VSS.n8957 0.019407
R18286 VSS.n8961 VSS.n8959 0.019407
R18287 VSS.n8964 VSS.n8962 0.019407
R18288 VSS.n963 VSS.n962 0.019407
R18289 VSS.n961 VSS.n960 0.019407
R18290 VSS.n959 VSS.n958 0.019407
R18291 VSS.n10283 VSS.n10282 0.019407
R18292 VSS.n10281 VSS.n10280 0.019407
R18293 VSS.n10279 VSS.n10278 0.019407
R18294 VSS.n9445 VSS.n9444 0.0192683
R18295 VSS.n9436 VSS.n9435 0.0192683
R18296 VSS.n8983 VSS.n8980 0.0189267
R18297 VSS.n8998 VSS.n8997 0.0189267
R18298 VSS.n1138 VSS.n1135 0.0189267
R18299 VSS.n911 VSS.n910 0.0189267
R18300 VSS.n10137 VSS.n10136 0.0189267
R18301 VSS.n1030 VSS.n1029 0.0189267
R18302 VSS.n10197 VSS.n10196 0.0189267
R18303 VSS.n950 VSS.n949 0.0189267
R18304 VSS.n10257 VSS.n10256 0.0189267
R18305 VSS.n11006 VSS.n11003 0.0189267
R18306 VSS.n10970 VSS.n10969 0.0189267
R18307 VSS.n9553 VSS.n9551 0.0189267
R18308 VSS.n9372 VSS.n9371 0.0189267
R18309 VSS.n9360 VSS.n9358 0.0189267
R18310 VSS.n9150 VSS.n9147 0.0189267
R18311 VSS.n9165 VSS.n9164 0.0189267
R18312 VSS VSS.n10823 0.0186978
R18313 VSS.n111 VSS.n110 0.0186448
R18314 VSS.n107 VSS.n106 0.0186448
R18315 VSS.n11385 VSS.n83 0.0186448
R18316 VSS.n83 VSS.n82 0.0186448
R18317 VSS.n11388 VSS.n79 0.0186448
R18318 VSS.n11397 VSS.n56 0.0186448
R18319 VSS.n11394 VSS.n55 0.0186448
R18320 VSS.n37 VSS.n30 0.0186448
R18321 VSS.n33 VSS.n30 0.0186448
R18322 VSS.n35 VSS.n29 0.0186448
R18323 VSS.n10704 VSS.n10702 0.0186448
R18324 VSS.n10704 VSS.n10699 0.0186448
R18325 VSS.n10705 VSS.n10700 0.0186448
R18326 VSS.n11307 VSS.n11306 0.0186448
R18327 VSS.n11307 VSS.n126 0.0186448
R18328 VSS.n11312 VSS.n11311 0.0186448
R18329 VSS.n10564 VSS.n10557 0.0186448
R18330 VSS.n10568 VSS.n10557 0.0186448
R18331 VSS.n10569 VSS.n10562 0.0186448
R18332 VSS.n10568 VSS.n10563 0.0186448
R18333 VSS.n10566 VSS.n10562 0.0186448
R18334 VSS.n10571 VSS.n10564 0.0186448
R18335 VSS.n230 VSS.n226 0.0186448
R18336 VSS.n10911 VSS.n225 0.0186448
R18337 VSS.n230 VSS.n229 0.0186448
R18338 VSS.n10912 VSS.n10911 0.0186448
R18339 VSS.n227 VSS.n226 0.0186448
R18340 VSS.n108 VSS.n107 0.0186448
R18341 VSS.n110 VSS.n109 0.0186448
R18342 VSS.n37 VSS.n32 0.0186448
R18343 VSS.n11432 VSS.n33 0.0186448
R18344 VSS.n11430 VSS.n29 0.0186448
R18345 VSS.n11396 VSS.n55 0.0186448
R18346 VSS.n11397 VSS.n58 0.0186448
R18347 VSS.n11386 VSS.n11385 0.0186448
R18348 VSS.n11383 VSS.n79 0.0186448
R18349 VSS.n82 VSS.n62 0.0186448
R18350 VSS.n11311 VSS.n124 0.0186448
R18351 VSS.n126 VSS.n122 0.0186448
R18352 VSS.n11309 VSS.n11306 0.0186448
R18353 VSS.n10729 VSS.n10700 0.0186448
R18354 VSS.n10707 VSS.n10699 0.0186448
R18355 VSS.n10731 VSS.n10702 0.0186448
R18356 VSS.n9077 VSS.n9076 0.0184746
R18357 VSS.n9107 VSS.n9106 0.0184746
R18358 VSS.n855 VSS.n854 0.0184746
R18359 VSS.n848 VSS.n847 0.0184746
R18360 VSS.n1101 VSS.n1100 0.0184746
R18361 VSS.n1275 VSS.n1274 0.0184746
R18362 VSS.n921 VSS.n920 0.0184746
R18363 VSS.n377 VSS.n376 0.0184746
R18364 VSS.n994 VSS.n993 0.0184746
R18365 VSS.n293 VSS.n292 0.0184746
R18366 VSS.n11065 VSS.n11064 0.0184746
R18367 VSS.n11074 VSS.n11073 0.0184746
R18368 VSS.n11220 VSS.n11219 0.0184746
R18369 VSS.n11213 VSS.n11212 0.0184746
R18370 VSS.n1170 VSS.n1169 0.0184746
R18371 VSS.n1191 VSS.n1190 0.0184746
R18372 VSS.n9397 VSS.n9396 0.0184746
R18373 VSS.n9406 VSS.n9405 0.0184746
R18374 VSS.n9234 VSS.n9233 0.0184746
R18375 VSS.n9227 VSS.n9226 0.0184746
R18376 VSS.n898 VSS.n897 0.0183443
R18377 VSS.n1067 VSS.n1066 0.0183443
R18378 VSS.n10169 VSS.n10167 0.0183443
R18379 VSS.n937 VSS.n936 0.0183443
R18380 VSS.n10229 VSS.n10227 0.0183443
R18381 VSS.n10909 VSS.n10908 0.0183443
R18382 VSS.n713 VSS.n711 0.0183443
R18383 VSS.n1227 VSS.n1225 0.0183443
R18384 VSS.n9272 VSS.n9269 0.0183443
R18385 VSS.n9287 VSS.n9286 0.0183443
R18386 VSS.n9054 VSS.n9053 0.0183443
R18387 VSS.n9127 VSS.n9126 0.0183443
R18388 VSS.n9069 VSS.n9068 0.0183136
R18389 VSS.n9089 VSS.n9044 0.0183136
R18390 VSS.n9015 VSS.n1561 0.0183136
R18391 VSS.n1289 VSS.n1288 0.0183136
R18392 VSS.n10153 VSS.n10152 0.0183136
R18393 VSS.n391 VSS.n390 0.0183136
R18394 VSS.n370 VSS.n369 0.0183136
R18395 VSS.n10213 VSS.n10212 0.0183136
R18396 VSS.n319 VSS.n318 0.0183136
R18397 VSS.n307 VSS.n306 0.0183136
R18398 VSS.n10273 VSS.n10272 0.0183136
R18399 VSS.n9382 VSS.n9380 0.0183136
R18400 VSS.n9344 VSS.n9320 0.0183136
R18401 VSS.n9309 VSS.n1505 0.0183136
R18402 VSS.n9246 VSS.n9211 0.0183136
R18403 VSS.n9182 VSS.n1523 0.0183136
R18404 VSS.n10060 VSS.n536 0.0182205
R18405 VSS.n11078 VSS.n11077 0.0182205
R18406 VSS.n11223 VSS.n11222 0.0182205
R18407 VSS.n9823 VSS.n768 0.0182205
R18408 VSS.n9467 VSS.n1380 0.0181966
R18409 VSS.n10771 VSS.n10770 0.0181748
R18410 VSS.n9463 VSS.n9452 0.0180195
R18411 VSS.n958 VSS.n253 0.0180018
R18412 VSS.n8985 VSS.n8984 0.0179991
R18413 VSS.n8994 VSS.n8993 0.0179991
R18414 VSS.n1140 VSS.n1139 0.0179991
R18415 VSS.n1149 VSS.n1148 0.0179991
R18416 VSS.n908 VSS.n907 0.0179991
R18417 VSS.n10133 VSS.n10132 0.0179991
R18418 VSS.n1027 VSS.n1026 0.0179991
R18419 VSS.n10193 VSS.n10192 0.0179991
R18420 VSS.n947 VSS.n946 0.0179991
R18421 VSS.n10253 VSS.n10252 0.0179991
R18422 VSS.n11008 VSS.n11007 0.0179991
R18423 VSS.n11017 VSS.n11016 0.0179991
R18424 VSS.n10957 VSS.n10956 0.0179991
R18425 VSS.n10966 VSS.n10965 0.0179991
R18426 VSS.n1155 VSS.n1154 0.0179991
R18427 VSS.n9555 VSS.n9554 0.0179991
R18428 VSS.n9369 VSS.n9368 0.0179991
R18429 VSS.n9362 VSS.n9361 0.0179991
R18430 VSS.n9152 VSS.n9151 0.0179991
R18431 VSS.n9161 VSS.n9160 0.0179991
R18432 VSS.n1147 VSS.n491 0.0177518
R18433 VSS.n11022 VSS.n11020 0.0177518
R18434 VSS.n10955 VSS.n151 0.0177518
R18435 VSS.n9781 VSS.n793 0.0177518
R18436 VSS.n2253 VSS.n61 0.01775
R18437 VSS.n895 VSS.n894 0.0174461
R18438 VSS.n888 VSS.n887 0.0174461
R18439 VSS.n1064 VSS.n1063 0.0174461
R18440 VSS.n10171 VSS.n10170 0.0174461
R18441 VSS.n934 VSS.n933 0.0174461
R18442 VSS.n10231 VSS.n10230 0.0174461
R18443 VSS.n10906 VSS.n10905 0.0174461
R18444 VSS.n10899 VSS.n10898 0.0174461
R18445 VSS.n722 VSS.n721 0.0174461
R18446 VSS.n715 VSS.n714 0.0174461
R18447 VSS.n1435 VSS.n1434 0.0174461
R18448 VSS.n1229 VSS.n1228 0.0174461
R18449 VSS.n9274 VSS.n9273 0.0174461
R18450 VSS.n9283 VSS.n9282 0.0174461
R18451 VSS.n9051 VSS.n9050 0.0174461
R18452 VSS.n9123 VSS.n9122 0.0174461
R18453 VSS.n9443 VSS.n9442 0.0174024
R18454 VSS.n9438 VSS.n9437 0.0174024
R18455 VSS.n10757 VSS.n10740 0.0173337
R18456 VSS.n10755 VSS.n10740 0.0173337
R18457 VSS.n886 VSS.n448 0.0172066
R18458 VSS.n10897 VSS.n10895 0.0172066
R18459 VSS.n725 VSS.n724 0.0172066
R18460 VSS.n1438 VSS.n1437 0.0172066
R18461 VSS.n1386 VSS.n811 0.0169894
R18462 VSS.n1332 VSS.n1327 0.0169894
R18463 VSS.n10759 VSS.n10758 0.0169128
R18464 VSS.n1408 VSS.n814 0.0167766
R18465 VSS.n9511 VSS.n9510 0.0167766
R18466 VSS.n9446 VSS.n9445 0.0167439
R18467 VSS.n9444 VSS.n9424 0.0167439
R18468 VSS.n9443 VSS.n9424 0.0167439
R18469 VSS.n9442 VSS.n9425 0.0167439
R18470 VSS.n9441 VSS.n9425 0.0167439
R18471 VSS.n9439 VSS.n9426 0.0167439
R18472 VSS.n9438 VSS.n9426 0.0167439
R18473 VSS.n9437 VSS.n9427 0.0167439
R18474 VSS.n9436 VSS.n9427 0.0167439
R18475 VSS.n9435 VSS.n9428 0.0167439
R18476 VSS.n10726 VSS.n10708 0.0167142
R18477 VSS.n10725 VSS.n10708 0.0167142
R18478 VSS.n10724 VSS.n10709 0.0167142
R18479 VSS.n10723 VSS.n10709 0.0167142
R18480 VSS.n10722 VSS.n10710 0.0167142
R18481 VSS.n10721 VSS.n10710 0.0167142
R18482 VSS.n10719 VSS.n10711 0.0167142
R18483 VSS.n10718 VSS.n10711 0.0167142
R18484 VSS.n1387 VSS.n814 0.0166702
R18485 VSS.n9511 VSS.n1333 0.0166702
R18486 VSS.n10677 VSS.n10335 0.016599
R18487 VSS.n9648 VSS.n9647 0.0164965
R18488 VSS.n9646 VSS.n9645 0.0164965
R18489 VSS.n9644 VSS.n9643 0.0164965
R18490 VSS.n780 VSS.n779 0.0164965
R18491 VSS.n782 VSS.n781 0.0164965
R18492 VSS.n784 VSS.n783 0.0164965
R18493 VSS.n662 VSS.n661 0.0164965
R18494 VSS.n664 VSS.n663 0.0164965
R18495 VSS.n666 VSS.n665 0.0164965
R18496 VSS.n9870 VSS.n9869 0.0164965
R18497 VSS.n9868 VSS.n9867 0.0164965
R18498 VSS.n9866 VSS.n9865 0.0164965
R18499 VSS.n1262 VSS.n1261 0.0164965
R18500 VSS.n1264 VSS.n1263 0.0164965
R18501 VSS.n1266 VSS.n1265 0.0164965
R18502 VSS.n1246 VSS.n1245 0.0164965
R18503 VSS.n1244 VSS.n1243 0.0164965
R18504 VSS.n1242 VSS.n1241 0.0164965
R18505 VSS.n636 VSS.n635 0.0164965
R18506 VSS.n638 VSS.n637 0.0164965
R18507 VSS.n640 VSS.n639 0.0164965
R18508 VSS.n9656 VSS.n9655 0.0164965
R18509 VSS.n9658 VSS.n9657 0.0164965
R18510 VSS.n9660 VSS.n9659 0.0164965
R18511 VSS.n592 VSS.n591 0.0164965
R18512 VSS.n594 VSS.n593 0.0164965
R18513 VSS.n596 VSS.n595 0.0164965
R18514 VSS.n9929 VSS.n9928 0.0164965
R18515 VSS.n9931 VSS.n9930 0.0164965
R18516 VSS.n9933 VSS.n9932 0.0164965
R18517 VSS.n11049 VSS.n11048 0.0164965
R18518 VSS.n11047 VSS.n11046 0.0164965
R18519 VSS.n11045 VSS.n11044 0.0164965
R18520 VSS.n9949 VSS.n9948 0.0164965
R18521 VSS.n9951 VSS.n9950 0.0164965
R18522 VSS.n9953 VSS.n9952 0.0164965
R18523 VSS.n9965 VSS.n9964 0.0164965
R18524 VSS.n9963 VSS.n9962 0.0164965
R18525 VSS.n9961 VSS.n9960 0.0164965
R18526 VSS.n11189 VSS.n11188 0.0164965
R18527 VSS.n11191 VSS.n11190 0.0164965
R18528 VSS.n11193 VSS.n11192 0.0164965
R18529 VSS.n9624 VSS.n9623 0.0164965
R18530 VSS.n9622 VSS.n9621 0.0164965
R18531 VSS.n9620 VSS.n9619 0.0164965
R18532 VSS.n9608 VSS.n9607 0.0164965
R18533 VSS.n9606 VSS.n9605 0.0164965
R18534 VSS.n9604 VSS.n9603 0.0164965
R18535 VSS.n9480 VSS.n811 0.0164574
R18536 VSS.n1327 VSS.n1326 0.0164574
R18537 VSS.n10754 VSS.n10753 0.0164441
R18538 VSS.n9691 VSS.n9690 0.0163916
R18539 VSS.n9688 VSS.n9687 0.0163916
R18540 VSS.n9685 VSS.n9684 0.0163916
R18541 VSS.n9851 VSS.n9850 0.0163916
R18542 VSS.n9848 VSS.n9847 0.0163916
R18543 VSS.n9845 VSS.n9844 0.0163916
R18544 VSS.n606 VSS.n605 0.0163916
R18545 VSS.n611 VSS.n610 0.0163916
R18546 VSS.n616 VSS.n615 0.0163916
R18547 VSS.n9703 VSS.n9702 0.0163916
R18548 VSS.n9708 VSS.n9707 0.0163916
R18549 VSS.n9713 VSS.n9712 0.0163916
R18550 VSS.n10743 VSS.n10742 0.0160769
R18551 VSS.n10497 VSS.n10496 0.0160245
R18552 VSS.n10495 VSS.n10494 0.0160245
R18553 VSS.n10606 VSS.n10605 0.0160245
R18554 VSS.n10608 VSS.n10607 0.0160245
R18555 VSS.n9649 VSS.n9639 0.0160245
R18556 VSS.n9648 VSS.n9639 0.0160245
R18557 VSS.n9647 VSS.n9640 0.0160245
R18558 VSS.n9646 VSS.n9640 0.0160245
R18559 VSS.n9645 VSS.n9641 0.0160245
R18560 VSS.n9644 VSS.n9641 0.0160245
R18561 VSS.n9643 VSS.n9642 0.0160245
R18562 VSS.n9642 VSS.n649 0.0160245
R18563 VSS.n9885 VSS.n647 0.0160245
R18564 VSS.n778 VSS.n777 0.0160245
R18565 VSS.n779 VSS.n777 0.0160245
R18566 VSS.n780 VSS.n776 0.0160245
R18567 VSS.n781 VSS.n776 0.0160245
R18568 VSS.n782 VSS.n775 0.0160245
R18569 VSS.n783 VSS.n775 0.0160245
R18570 VSS.n784 VSS.n774 0.0160245
R18571 VSS.n785 VSS.n774 0.0160245
R18572 VSS.n660 VSS.n578 0.0160245
R18573 VSS.n661 VSS.n660 0.0160245
R18574 VSS.n662 VSS.n659 0.0160245
R18575 VSS.n663 VSS.n659 0.0160245
R18576 VSS.n664 VSS.n658 0.0160245
R18577 VSS.n665 VSS.n658 0.0160245
R18578 VSS.n666 VSS.n657 0.0160245
R18579 VSS.n667 VSS.n657 0.0160245
R18580 VSS.n673 VSS.n672 0.0160245
R18581 VSS.n9871 VSS.n9860 0.0160245
R18582 VSS.n9870 VSS.n9860 0.0160245
R18583 VSS.n9869 VSS.n9861 0.0160245
R18584 VSS.n9868 VSS.n9861 0.0160245
R18585 VSS.n9867 VSS.n9862 0.0160245
R18586 VSS.n9866 VSS.n9862 0.0160245
R18587 VSS.n9865 VSS.n9863 0.0160245
R18588 VSS.n9864 VSS.n9863 0.0160245
R18589 VSS.n1260 VSS.n1259 0.0160245
R18590 VSS.n1261 VSS.n1259 0.0160245
R18591 VSS.n1262 VSS.n1258 0.0160245
R18592 VSS.n1263 VSS.n1258 0.0160245
R18593 VSS.n1264 VSS.n1257 0.0160245
R18594 VSS.n1265 VSS.n1257 0.0160245
R18595 VSS.n1266 VSS.n1256 0.0160245
R18596 VSS.n1267 VSS.n1256 0.0160245
R18597 VSS.n9519 VSS.n1236 0.0160245
R18598 VSS.n1247 VSS.n1237 0.0160245
R18599 VSS.n1246 VSS.n1237 0.0160245
R18600 VSS.n1245 VSS.n1238 0.0160245
R18601 VSS.n1244 VSS.n1238 0.0160245
R18602 VSS.n1243 VSS.n1239 0.0160245
R18603 VSS.n1242 VSS.n1239 0.0160245
R18604 VSS.n1241 VSS.n1240 0.0160245
R18605 VSS.n1240 VSS.n804 0.0160245
R18606 VSS.n634 VSS.n633 0.0160245
R18607 VSS.n635 VSS.n633 0.0160245
R18608 VSS.n636 VSS.n632 0.0160245
R18609 VSS.n637 VSS.n632 0.0160245
R18610 VSS.n638 VSS.n631 0.0160245
R18611 VSS.n639 VSS.n631 0.0160245
R18612 VSS.n640 VSS.n630 0.0160245
R18613 VSS.n641 VSS.n630 0.0160245
R18614 VSS.n9894 VSS.n643 0.0160245
R18615 VSS.n9654 VSS.n9653 0.0160245
R18616 VSS.n9655 VSS.n9653 0.0160245
R18617 VSS.n9656 VSS.n9652 0.0160245
R18618 VSS.n9657 VSS.n9652 0.0160245
R18619 VSS.n9658 VSS.n9651 0.0160245
R18620 VSS.n9659 VSS.n9651 0.0160245
R18621 VSS.n9660 VSS.n9650 0.0160245
R18622 VSS.n9661 VSS.n9650 0.0160245
R18623 VSS.n590 VSS.n589 0.0160245
R18624 VSS.n591 VSS.n589 0.0160245
R18625 VSS.n592 VSS.n588 0.0160245
R18626 VSS.n593 VSS.n588 0.0160245
R18627 VSS.n594 VSS.n587 0.0160245
R18628 VSS.n595 VSS.n587 0.0160245
R18629 VSS.n596 VSS.n586 0.0160245
R18630 VSS.n597 VSS.n586 0.0160245
R18631 VSS.n9915 VSS.n583 0.0160245
R18632 VSS.n9927 VSS.n582 0.0160245
R18633 VSS.n9928 VSS.n582 0.0160245
R18634 VSS.n9929 VSS.n581 0.0160245
R18635 VSS.n9930 VSS.n581 0.0160245
R18636 VSS.n9931 VSS.n580 0.0160245
R18637 VSS.n9932 VSS.n580 0.0160245
R18638 VSS.n9933 VSS.n579 0.0160245
R18639 VSS.n9934 VSS.n579 0.0160245
R18640 VSS.n11050 VSS.n11039 0.0160245
R18641 VSS.n11049 VSS.n11039 0.0160245
R18642 VSS.n11048 VSS.n11040 0.0160245
R18643 VSS.n11047 VSS.n11040 0.0160245
R18644 VSS.n11046 VSS.n11041 0.0160245
R18645 VSS.n11045 VSS.n11041 0.0160245
R18646 VSS.n11044 VSS.n11042 0.0160245
R18647 VSS.n11043 VSS.n11042 0.0160245
R18648 VSS.n11283 VSS.n11282 0.0160245
R18649 VSS.n9947 VSS.n9946 0.0160245
R18650 VSS.n9948 VSS.n9946 0.0160245
R18651 VSS.n9949 VSS.n9945 0.0160245
R18652 VSS.n9950 VSS.n9945 0.0160245
R18653 VSS.n9951 VSS.n9944 0.0160245
R18654 VSS.n9952 VSS.n9944 0.0160245
R18655 VSS.n9953 VSS.n9943 0.0160245
R18656 VSS.n9954 VSS.n9943 0.0160245
R18657 VSS.n9966 VSS.n9955 0.0160245
R18658 VSS.n9965 VSS.n9955 0.0160245
R18659 VSS.n9964 VSS.n9956 0.0160245
R18660 VSS.n9963 VSS.n9956 0.0160245
R18661 VSS.n9962 VSS.n9957 0.0160245
R18662 VSS.n9961 VSS.n9957 0.0160245
R18663 VSS.n9960 VSS.n9958 0.0160245
R18664 VSS.n9959 VSS.n9958 0.0160245
R18665 VSS.n142 VSS.n141 0.0160245
R18666 VSS.n11187 VSS.n11186 0.0160245
R18667 VSS.n11188 VSS.n11186 0.0160245
R18668 VSS.n11189 VSS.n11185 0.0160245
R18669 VSS.n11190 VSS.n11185 0.0160245
R18670 VSS.n11191 VSS.n11184 0.0160245
R18671 VSS.n11192 VSS.n11184 0.0160245
R18672 VSS.n11193 VSS.n11183 0.0160245
R18673 VSS.n11194 VSS.n11183 0.0160245
R18674 VSS.n9625 VSS.n806 0.0160245
R18675 VSS.n9624 VSS.n806 0.0160245
R18676 VSS.n9623 VSS.n807 0.0160245
R18677 VSS.n9622 VSS.n807 0.0160245
R18678 VSS.n9621 VSS.n808 0.0160245
R18679 VSS.n9620 VSS.n808 0.0160245
R18680 VSS.n9619 VSS.n809 0.0160245
R18681 VSS.n9618 VSS.n809 0.0160245
R18682 VSS.n1233 VSS.n810 0.0160245
R18683 VSS.n9609 VSS.n823 0.0160245
R18684 VSS.n9608 VSS.n823 0.0160245
R18685 VSS.n9607 VSS.n824 0.0160245
R18686 VSS.n9606 VSS.n824 0.0160245
R18687 VSS.n9605 VSS.n825 0.0160245
R18688 VSS.n9604 VSS.n825 0.0160245
R18689 VSS.n9603 VSS.n826 0.0160245
R18690 VSS.n9602 VSS.n826 0.0160245
R18691 VSS.n10824 VSS 0.0159286
R18692 VSS.n9672 VSS.n9671 0.0159196
R18693 VSS.n9692 VSS.n9673 0.0159196
R18694 VSS.n9675 VSS.n9674 0.0159196
R18695 VSS.n9689 VSS.n9676 0.0159196
R18696 VSS.n9678 VSS.n9677 0.0159196
R18697 VSS.n9686 VSS.n9679 0.0159196
R18698 VSS.n9681 VSS.n9680 0.0159196
R18699 VSS.n9683 VSS.n9682 0.0159196
R18700 VSS.n681 VSS.n680 0.0159196
R18701 VSS.n9852 VSS.n682 0.0159196
R18702 VSS.n684 VSS.n683 0.0159196
R18703 VSS.n9849 VSS.n685 0.0159196
R18704 VSS.n687 VSS.n686 0.0159196
R18705 VSS.n9846 VSS.n688 0.0159196
R18706 VSS.n690 VSS.n689 0.0159196
R18707 VSS.n9843 VSS.n691 0.0159196
R18708 VSS.n604 VSS.n603 0.0159196
R18709 VSS.n602 VSS.n601 0.0159196
R18710 VSS.n609 VSS.n608 0.0159196
R18711 VSS.n607 VSS.n600 0.0159196
R18712 VSS.n614 VSS.n613 0.0159196
R18713 VSS.n612 VSS.n599 0.0159196
R18714 VSS.n619 VSS.n618 0.0159196
R18715 VSS.n617 VSS.n598 0.0159196
R18716 VSS.n9701 VSS.n9700 0.0159196
R18717 VSS.n9699 VSS.n9697 0.0159196
R18718 VSS.n9706 VSS.n9705 0.0159196
R18719 VSS.n9704 VSS.n9696 0.0159196
R18720 VSS.n9711 VSS.n9710 0.0159196
R18721 VSS.n9709 VSS.n9695 0.0159196
R18722 VSS.n9716 VSS.n9715 0.0159196
R18723 VSS.n9714 VSS.n9694 0.0159196
R18724 VSS.n10439 VSS.n10335 0.0158871
R18725 VSS.n10587 VSS.n10586 0.0157873
R18726 VSS.n10814 VSS.n250 0.0156685
R18727 VSS.n10783 VSS.n10782 0.0156685
R18728 VSS.n10717 VSS.n10712 0.0156595
R18729 VSS.n9887 VSS.n9886 0.0156049
R18730 VSS.n671 VSS.n668 0.0156049
R18731 VSS.n9521 VSS.n9520 0.0156049
R18732 VSS.n9893 VSS.n9892 0.0156049
R18733 VSS.n9917 VSS.n9916 0.0156049
R18734 VSS.n11284 VSS.n11281 0.0156049
R18735 VSS.n143 VSS.n140 0.0156049
R18736 VSS.n1234 VSS.n815 0.0156049
R18737 VSS.n1177 VSS.n1176 0.0155
R18738 VSS.n1180 VSS.n1179 0.0155
R18739 VSS.n623 VSS.n622 0.0155
R18740 VSS.n9905 VSS.n626 0.0155
R18741 VSS.n11470 VSS.n3 0.0152621
R18742 VSS.n8955 VSS.n8954 0.0152551
R18743 VSS.n9094 VSS.n1554 0.01514
R18744 VSS.n9008 VSS.n8969 0.01514
R18745 VSS.n10927 VSS.n221 0.01514
R18746 VSS.n869 VSS.n868 0.01514
R18747 VSS.n1125 VSS.n1124 0.01514
R18748 VSS.n1113 VSS.n1112 0.01514
R18749 VSS.n1092 VSS.n1091 0.01514
R18750 VSS.n1076 VSS.n1075 0.01514
R18751 VSS.n1055 VSS.n1054 0.01514
R18752 VSS.n1043 VSS.n1042 0.01514
R18753 VSS.n1018 VSS.n1017 0.01514
R18754 VSS.n1006 VSS.n1005 0.01514
R18755 VSS.n985 VSS.n984 0.01514
R18756 VSS.n969 VSS.n968 0.01514
R18757 VSS.n10984 VSS.n207 0.01514
R18758 VSS.n11359 VSS.n96 0.01514
R18759 VSS.n11348 VSS.n11347 0.01514
R18760 VSS.n11376 VSS.n11374 0.01514
R18761 VSS.n11363 VSS.n90 0.01514
R18762 VSS.n10980 VSS.n10942 0.01514
R18763 VSS.n10931 VSS.n214 0.01514
R18764 VSS.n1206 VSS.n1205 0.01514
R18765 VSS.n9542 VSS.n9540 0.01514
R18766 VSS.n9529 VSS.n1221 0.01514
R18767 VSS.n9420 VSS.n1396 0.01514
R18768 VSS.n9349 VSS.n1496 0.01514
R18769 VSS.n9297 VSS.n9262 0.01514
R18770 VSS.n9251 VSS.n1513 0.01514
R18771 VSS.n9175 VSS.n9136 0.01514
R18772 VSS.n1548 VSS.n1547 0.01514
R18773 VSS.n9110 VSS.n9109 0.0150766
R18774 VSS.n853 VSS.n851 0.0150766
R18775 VSS.n10121 VSS.n427 0.0150766
R18776 VSS.n10181 VSS.n357 0.0150766
R18777 VSS.n10241 VSS.n285 0.0150766
R18778 VSS.n11069 VSS.n11068 0.0150766
R18779 VSS.n11216 VSS.n11215 0.0150766
R18780 VSS.n1189 VSS.n1186 0.0150766
R18781 VSS.n9404 VSS.n9401 0.0150766
R18782 VSS.n9230 VSS.n9229 0.0150766
R18783 VSS.n8992 VSS.n8989 0.014691
R18784 VSS.n1152 VSS.n1143 0.014691
R18785 VSS.n10128 VSS.n419 0.014691
R18786 VSS.n10188 VSS.n347 0.014691
R18787 VSS.n10248 VSS.n275 0.014691
R18788 VSS.n11012 VSS.n11011 0.014691
R18789 VSS.n10964 VSS.n10961 0.014691
R18790 VSS.n9558 VSS.n9557 0.014691
R18791 VSS.n9365 VSS.n9364 0.014691
R18792 VSS.n9159 VSS.n9156 0.014691
R18793 VSS.n78 VSS.n77 0.014605
R18794 VSS.n10716 VSS.n10712 0.0144843
R18795 VSS.n10715 VSS.n10713 0.0144843
R18796 VSS.n10714 VSS.n10713 0.0144843
R18797 VSS.n893 VSS.n891 0.0142425
R18798 VSS.n10174 VSS.n397 0.0142425
R18799 VSS.n10234 VSS.n325 0.0142425
R18800 VSS.n10904 VSS.n10902 0.0142425
R18801 VSS.n718 VSS.n717 0.0142425
R18802 VSS.n1232 VSS.n1231 0.0142425
R18803 VSS.n9281 VSS.n9278 0.0142425
R18804 VSS.n9121 VSS.n9118 0.0142425
R18805 VSS.n9038 VSS.n1560 0.0141709
R18806 VSS.n10144 VSS.n10142 0.0141709
R18807 VSS.n10204 VSS.n10202 0.0141709
R18808 VSS.n10264 VSS.n10262 0.0141709
R18809 VSS.n9336 VSS.n1478 0.0141709
R18810 VSS.n9205 VSS.n1522 0.0141709
R18811 VSS.n9629 VSS.n9628 0.0139852
R18812 VSS.n9755 VSS.n9754 0.0139852
R18813 VSS.n9750 VSS.n9749 0.0139852
R18814 VSS.n9733 VSS.n9732 0.0139852
R18815 VSS.n9728 VSS.n9727 0.0139852
R18816 VSS.n10013 VSS.n10012 0.0139852
R18817 VSS.n9996 VSS.n9995 0.0139852
R18818 VSS.n9991 VSS.n9990 0.0139852
R18819 VSS.n10634 VSS.n10633 0.0137679
R18820 VSS.n10748 VSS.n250 0.0136461
R18821 VSS.n10782 VSS.n10781 0.0136461
R18822 VSS.n11436 VSS.n11435 0.0133485
R18823 VSS.n11403 VSS.n11402 0.0133485
R18824 VSS.n11427 VSS.n11426 0.0132877
R18825 VSS.n9032 VSS.n9018 0.0132388
R18826 VSS.n10145 VSS.n403 0.0132388
R18827 VSS.n10205 VSS.n331 0.0132388
R18828 VSS.n10265 VSS.n259 0.0132388
R18829 VSS.n9337 VSS.n9322 0.0132388
R18830 VSS.n9199 VSS.n9185 0.0132388
R18831 VSS.n1363 VSS.n1362 0.013182
R18832 VSS.n9760 VSS.n9759 0.013182
R18833 VSS.n9738 VSS.n9737 0.013182
R18834 VSS.n10001 VSS.n10000 0.013182
R18835 VSS.n9979 VSS.n9978 0.013182
R18836 VSS.n8976 VSS.n8972 0.0127708
R18837 VSS.n874 VSS.n870 0.0127708
R18838 VSS.n1088 VSS.n904 0.0127708
R18839 VSS.n1039 VSS.n928 0.0127708
R18840 VSS.n981 VSS.n943 0.0127708
R18841 VSS.n10995 VSS.n10991 0.0127708
R18842 VSS.n10949 VSS.n10945 0.0127708
R18843 VSS.n1211 VSS.n1207 0.0127708
R18844 VSS.n1491 VSS.n1487 0.0127708
R18845 VSS.n9143 VSS.n9139 0.0127708
R18846 VSS.n9508 VSS.n1335 0.012534
R18847 VSS.n9493 VSS.n1374 0.0123788
R18848 VSS.n9974 VSS.n31 0.0123788
R18849 VSS.n1374 VSS.n1346 0.0123365
R18850 VSS.n1372 VSS.n1346 0.0123365
R18851 VSS.n1372 VSS.n1371 0.0123365
R18852 VSS.n1371 VSS.n1370 0.0123365
R18853 VSS.n1369 VSS.n1368 0.0123365
R18854 VSS.n1368 VSS.n1348 0.0123365
R18855 VSS.n1366 VSS.n1365 0.0123365
R18856 VSS.n1365 VSS.n1364 0.0123365
R18857 VSS.n1362 VSS.n1351 0.0123365
R18858 VSS.n1360 VSS.n1351 0.0123365
R18859 VSS.n1360 VSS.n1359 0.0123365
R18860 VSS.n1355 VSS.n1354 0.0123365
R18861 VSS.n1354 VSS.n805 0.0123365
R18862 VSS.n9627 VSS.n803 0.0123365
R18863 VSS.n9628 VSS.n803 0.0123365
R18864 VSS.n9629 VSS.n802 0.0123365
R18865 VSS.n9631 VSS.n802 0.0123365
R18866 VSS.n9631 VSS.n801 0.0123365
R18867 VSS.n9633 VSS.n801 0.0123365
R18868 VSS.n9635 VSS.n9634 0.0123365
R18869 VSS.n9635 VSS.n798 0.0123365
R18870 VSS.n9763 VSS.n800 0.0123365
R18871 VSS.n9761 VSS.n800 0.0123365
R18872 VSS.n9759 VSS.n9636 0.0123365
R18873 VSS.n9757 VSS.n9636 0.0123365
R18874 VSS.n9757 VSS.n9756 0.0123365
R18875 VSS.n9756 VSS.n9755 0.0123365
R18876 VSS.n9754 VSS.n9638 0.0123365
R18877 VSS.n9753 VSS.n9638 0.0123365
R18878 VSS.n9751 VSS.n9662 0.0123365
R18879 VSS.n9750 VSS.n9662 0.0123365
R18880 VSS.n9749 VSS.n9663 0.0123365
R18881 VSS.n9747 VSS.n9663 0.0123365
R18882 VSS.n9747 VSS.n9746 0.0123365
R18883 VSS.n9746 VSS.n9745 0.0123365
R18884 VSS.n9744 VSS.n9743 0.0123365
R18885 VSS.n9743 VSS.n9665 0.0123365
R18886 VSS.n9741 VSS.n9740 0.0123365
R18887 VSS.n9740 VSS.n9739 0.0123365
R18888 VSS.n9737 VSS.n9668 0.0123365
R18889 VSS.n9735 VSS.n9668 0.0123365
R18890 VSS.n9735 VSS.n9734 0.0123365
R18891 VSS.n9734 VSS.n9733 0.0123365
R18892 VSS.n9732 VSS.n9670 0.0123365
R18893 VSS.n9731 VSS.n9670 0.0123365
R18894 VSS.n9729 VSS.n9718 0.0123365
R18895 VSS.n9728 VSS.n9718 0.0123365
R18896 VSS.n9727 VSS.n9719 0.0123365
R18897 VSS.n9725 VSS.n9719 0.0123365
R18898 VSS.n9725 VSS.n9724 0.0123365
R18899 VSS.n9724 VSS.n9723 0.0123365
R18900 VSS.n9722 VSS.n9721 0.0123365
R18901 VSS.n9721 VSS.n569 0.0123365
R18902 VSS.n10029 VSS.n571 0.0123365
R18903 VSS.n10027 VSS.n571 0.0123365
R18904 VSS.n10022 VSS.n574 0.0123365
R18905 VSS.n10022 VSS.n10021 0.0123365
R18906 VSS.n10017 VSS.n577 0.0123365
R18907 VSS.n10016 VSS.n577 0.0123365
R18908 VSS.n10014 VSS.n9935 0.0123365
R18909 VSS.n10013 VSS.n9935 0.0123365
R18910 VSS.n10012 VSS.n9936 0.0123365
R18911 VSS.n10010 VSS.n9936 0.0123365
R18912 VSS.n10010 VSS.n10009 0.0123365
R18913 VSS.n10009 VSS.n10008 0.0123365
R18914 VSS.n10007 VSS.n10006 0.0123365
R18915 VSS.n10006 VSS.n9938 0.0123365
R18916 VSS.n10004 VSS.n10003 0.0123365
R18917 VSS.n10003 VSS.n10002 0.0123365
R18918 VSS.n10000 VSS.n9940 0.0123365
R18919 VSS.n9998 VSS.n9940 0.0123365
R18920 VSS.n9998 VSS.n9997 0.0123365
R18921 VSS.n9997 VSS.n9996 0.0123365
R18922 VSS.n9995 VSS.n9942 0.0123365
R18923 VSS.n9994 VSS.n9942 0.0123365
R18924 VSS.n9992 VSS.n9967 0.0123365
R18925 VSS.n9991 VSS.n9967 0.0123365
R18926 VSS.n9990 VSS.n9968 0.0123365
R18927 VSS.n9988 VSS.n9968 0.0123365
R18928 VSS.n9988 VSS.n9987 0.0123365
R18929 VSS.n9987 VSS.n9986 0.0123365
R18930 VSS.n9985 VSS.n9984 0.0123365
R18931 VSS.n9984 VSS.n9970 0.0123365
R18932 VSS.n9982 VSS.n9981 0.0123365
R18933 VSS.n9981 VSS.n9980 0.0123365
R18934 VSS.n9978 VSS.n9972 0.0123365
R18935 VSS.n9976 VSS.n9972 0.0123365
R18936 VSS.n9976 VSS.n9975 0.0123365
R18937 VSS.n9975 VSS.n9974 0.0123365
R18938 VSS.n10284 VSS.n253 0.0123169
R18939 VSS.n11460 VSS.n11459 0.0121335
R18940 VSS.n9068 VSS.n9067 0.0120995
R18941 VSS.n9089 VSS.n9088 0.0120995
R18942 VSS.n9016 VSS.n9015 0.0120995
R18943 VSS.n1290 VSS.n1289 0.0120995
R18944 VSS.n10152 VSS.n10151 0.0120995
R18945 VSS.n10159 VSS.n391 0.0120995
R18946 VSS.n371 VSS.n370 0.0120995
R18947 VSS.n10212 VSS.n10211 0.0120995
R18948 VSS.n10219 VSS.n319 0.0120995
R18949 VSS.n308 VSS.n307 0.0120995
R18950 VSS.n10272 VSS.n10271 0.0120995
R18951 VSS.n9383 VSS.n9382 0.0120995
R18952 VSS.n9344 VSS.n9343 0.0120995
R18953 VSS.n9310 VSS.n9309 0.0120995
R18954 VSS.n9246 VSS.n9245 0.0120995
R18955 VSS.n9183 VSS.n9182 0.0120995
R18956 VSS.n1349 VSS.n1348 0.0119138
R18957 VSS.n9764 VSS.n798 0.0119138
R18958 VSS.n9666 VSS.n9665 0.0119138
R18959 VSS.n10030 VSS.n569 0.0119138
R18960 VSS.n9938 VSS.n147 0.0119138
R18961 VSS.n9970 VSS.n138 0.0119138
R18962 VSS.n10727 VSS.n10726 0.0118938
R18963 VSS.n10725 VSS.n10724 0.0118938
R18964 VSS.n10723 VSS.n10722 0.0118938
R18965 VSS.n10718 VSS.n10717 0.0118938
R18966 VSS.n10772 VSS.n10771 0.0118287
R18967 VSS.n10774 VSS.n10773 0.011514
R18968 VSS.n9626 VSS.n805 0.0114911
R18969 VSS.n9627 VSS.n9626 0.0114911
R18970 VSS.n9753 VSS.n9752 0.0114911
R18971 VSS.n9752 VSS.n9751 0.0114911
R18972 VSS.n9731 VSS.n9730 0.0114911
R18973 VSS.n9730 VSS.n9729 0.0114911
R18974 VSS.n10016 VSS.n10015 0.0114911
R18975 VSS.n10015 VSS.n10014 0.0114911
R18976 VSS.n9994 VSS.n9993 0.0114911
R18977 VSS.n9993 VSS.n9992 0.0114911
R18978 VSS.n10638 VSS.n10352 0.0113855
R18979 VSS.n10610 VSS.n10440 0.0113305
R18980 VSS.n11336 VSS.n11335 0.0112405
R18981 VSS.n1356 VSS.n1355 0.0111529
R18982 VSS.n10018 VSS.n10017 0.0111529
R18983 VSS.n11434 VSS.n11433 0.0111311
R18984 VSS.n10745 VSS.n10744 0.0105699
R18985 VSS.n10755 VSS.n10754 0.0105401
R18986 VSS.n10026 VSS.n10025 0.0105188
R18987 VSS.n10728 VSS.n10727 0.0104148
R18988 VSS.n10716 VSS.n10715 0.0103268
R18989 VSS.n10714 VSS.n125 0.0103268
R18990 VSS.n9110 VSS.n1536 0.0102495
R18991 VSS.n851 VSS.n850 0.0102495
R18992 VSS.n10121 VSS.n430 0.0102495
R18993 VSS.n10181 VSS.n360 0.0102495
R18994 VSS.n10241 VSS.n288 0.0102495
R18995 VSS.n11072 VSS.n11069 0.0102495
R18996 VSS.n11218 VSS.n11216 0.0102495
R18997 VSS.n1186 VSS.n1173 0.0102495
R18998 VSS.n9401 VSS.n9400 0.0102495
R18999 VSS.n9232 VSS.n9230 0.0102495
R19000 VSS.n10574 VSS.n10573 0.0101279
R19001 VSS.n10857 VSS.n10856 0.00999301
R19002 VSS.n8989 VSS.n8988 0.00999158
R19003 VSS.n1152 VSS.n1151 0.00999158
R19004 VSS.n10131 VSS.n10128 0.00999158
R19005 VSS.n10191 VSS.n10188 0.00999158
R19006 VSS.n10251 VSS.n10248 0.00999158
R19007 VSS.n11015 VSS.n11012 0.00999158
R19008 VSS.n10961 VSS.n10960 0.00999158
R19009 VSS.n9558 VSS.n1158 0.00999158
R19010 VSS.n9367 VSS.n9365 0.00999158
R19011 VSS.n9156 VSS.n9155 0.00999158
R19012 VSS.n1359 VSS.n1358 0.00992696
R19013 VSS.n10021 VSS.n10020 0.00992696
R19014 VSS.n9082 VSS.n9080 0.00990014
R19015 VSS.n9079 VSS.n9077 0.00990014
R19016 VSS.n9076 VSS.n1536 0.00990014
R19017 VSS.n9109 VSS.n9107 0.00990014
R19018 VSS.n9106 VSS.n9105 0.00990014
R19019 VSS.n9103 VSS.n9102 0.00990014
R19020 VSS.n860 VSS.n858 0.00990014
R19021 VSS.n857 VSS.n855 0.00990014
R19022 VSS.n854 VSS.n853 0.00990014
R19023 VSS.n850 VSS.n848 0.00990014
R19024 VSS.n847 VSS.n536 0.00990014
R19025 VSS.n1106 VSS.n1104 0.00990014
R19026 VSS.n1103 VSS.n1101 0.00990014
R19027 VSS.n1100 VSS.n427 0.00990014
R19028 VSS.n1274 VSS.n430 0.00990014
R19029 VSS.n1278 VSS.n1275 0.00990014
R19030 VSS.n1282 VSS.n1279 0.00990014
R19031 VSS.n926 VSS.n924 0.00990014
R19032 VSS.n923 VSS.n921 0.00990014
R19033 VSS.n920 VSS.n357 0.00990014
R19034 VSS.n376 VSS.n360 0.00990014
R19035 VSS.n380 VSS.n377 0.00990014
R19036 VSS.n384 VSS.n381 0.00990014
R19037 VSS.n999 VSS.n997 0.00990014
R19038 VSS.n996 VSS.n994 0.00990014
R19039 VSS.n993 VSS.n285 0.00990014
R19040 VSS.n292 VSS.n288 0.00990014
R19041 VSS.n296 VSS.n293 0.00990014
R19042 VSS.n300 VSS.n297 0.00990014
R19043 VSS.n11060 VSS.n100 0.00990014
R19044 VSS.n11064 VSS.n11063 0.00990014
R19045 VSS.n11068 VSS.n11065 0.00990014
R19046 VSS.n11073 VSS.n11072 0.00990014
R19047 VSS.n11077 VSS.n11074 0.00990014
R19048 VSS.n11222 VSS.n11220 0.00990014
R19049 VSS.n11219 VSS.n11218 0.00990014
R19050 VSS.n11215 VSS.n11213 0.00990014
R19051 VSS.n11212 VSS.n11211 0.00990014
R19052 VSS.n11209 VSS.n88 0.00990014
R19053 VSS.n1169 VSS.n768 0.00990014
R19054 VSS.n1173 VSS.n1170 0.00990014
R19055 VSS.n1190 VSS.n1189 0.00990014
R19056 VSS.n1194 VSS.n1191 0.00990014
R19057 VSS.n1198 VSS.n1195 0.00990014
R19058 VSS.n9392 VSS.n9391 0.00990014
R19059 VSS.n9396 VSS.n9395 0.00990014
R19060 VSS.n9400 VSS.n9397 0.00990014
R19061 VSS.n9405 VSS.n9404 0.00990014
R19062 VSS.n9409 VSS.n9406 0.00990014
R19063 VSS.n9413 VSS.n9410 0.00990014
R19064 VSS.n9239 VSS.n9237 0.00990014
R19065 VSS.n9236 VSS.n9234 0.00990014
R19066 VSS.n9233 VSS.n9232 0.00990014
R19067 VSS.n9229 VSS.n9227 0.00990014
R19068 VSS.n9226 VSS.n9225 0.00990014
R19069 VSS.n9223 VSS.n1511 0.00990014
R19070 VSS.n11458 VSS.n11457 0.00976426
R19071 VSS.n11456 VSS.n11455 0.00976426
R19072 VSS.n11454 VSS.n11453 0.00976426
R19073 VSS.n11442 VSS.n11441 0.00976426
R19074 VSS.n11440 VSS.n11439 0.00976426
R19075 VSS.n11438 VSS.n11437 0.00976426
R19076 VSS.n11425 VSS.n11424 0.00976426
R19077 VSS.n11423 VSS.n11422 0.00976426
R19078 VSS.n11421 VSS.n11420 0.00976426
R19079 VSS.n11409 VSS.n11408 0.00976426
R19080 VSS.n11407 VSS.n11406 0.00976426
R19081 VSS.n11405 VSS.n11404 0.00976426
R19082 VSS.n574 VSS.n573 0.00975787
R19083 VSS.n891 VSS.n890 0.00969162
R19084 VSS.n10174 VSS.n10173 0.00969162
R19085 VSS.n10234 VSS.n10233 0.00969162
R19086 VSS.n10902 VSS.n10901 0.00969162
R19087 VSS.n720 VSS.n718 0.00969162
R19088 VSS.n1433 VSS.n1232 0.00969162
R19089 VSS.n9278 VSS.n9277 0.00969162
R19090 VSS.n9118 VSS.n1530 0.00969162
R19091 VSS.n8980 VSS.n1559 0.00965149
R19092 VSS.n8984 VSS.n8983 0.00965149
R19093 VSS.n8988 VSS.n8985 0.00965149
R19094 VSS.n8993 VSS.n8992 0.00965149
R19095 VSS.n8997 VSS.n8994 0.00965149
R19096 VSS.n9001 VSS.n8998 0.00965149
R19097 VSS.n1135 VSS.n1134 0.00965149
R19098 VSS.n1139 VSS.n1138 0.00965149
R19099 VSS.n1143 VSS.n1140 0.00965149
R19100 VSS.n1151 VSS.n1149 0.00965149
R19101 VSS.n1148 VSS.n1147 0.00965149
R19102 VSS.n913 VSS.n911 0.00965149
R19103 VSS.n910 VSS.n908 0.00965149
R19104 VSS.n907 VSS.n419 0.00965149
R19105 VSS.n10132 VSS.n10131 0.00965149
R19106 VSS.n10136 VSS.n10133 0.00965149
R19107 VSS.n10140 VSS.n10137 0.00965149
R19108 VSS.n1032 VSS.n1030 0.00965149
R19109 VSS.n1029 VSS.n1027 0.00965149
R19110 VSS.n1026 VSS.n347 0.00965149
R19111 VSS.n10192 VSS.n10191 0.00965149
R19112 VSS.n10196 VSS.n10193 0.00965149
R19113 VSS.n10200 VSS.n10197 0.00965149
R19114 VSS.n952 VSS.n950 0.00965149
R19115 VSS.n949 VSS.n947 0.00965149
R19116 VSS.n946 VSS.n275 0.00965149
R19117 VSS.n10252 VSS.n10251 0.00965149
R19118 VSS.n10256 VSS.n10253 0.00965149
R19119 VSS.n10260 VSS.n10257 0.00965149
R19120 VSS.n11003 VSS.n11002 0.00965149
R19121 VSS.n11007 VSS.n11006 0.00965149
R19122 VSS.n11011 VSS.n11008 0.00965149
R19123 VSS.n11016 VSS.n11015 0.00965149
R19124 VSS.n11020 VSS.n11017 0.00965149
R19125 VSS.n10956 VSS.n10955 0.00965149
R19126 VSS.n10960 VSS.n10957 0.00965149
R19127 VSS.n10965 VSS.n10964 0.00965149
R19128 VSS.n10969 VSS.n10966 0.00965149
R19129 VSS.n10973 VSS.n10970 0.00965149
R19130 VSS.n1154 VSS.n793 0.00965149
R19131 VSS.n1158 VSS.n1155 0.00965149
R19132 VSS.n9557 VSS.n9555 0.00965149
R19133 VSS.n9554 VSS.n9553 0.00965149
R19134 VSS.n9551 VSS.n9550 0.00965149
R19135 VSS.n9374 VSS.n9372 0.00965149
R19136 VSS.n9371 VSS.n9369 0.00965149
R19137 VSS.n9368 VSS.n9367 0.00965149
R19138 VSS.n9364 VSS.n9362 0.00965149
R19139 VSS.n9361 VSS.n9360 0.00965149
R19140 VSS.n9358 VSS.n9357 0.00965149
R19141 VSS.n9147 VSS.n1521 0.00965149
R19142 VSS.n9151 VSS.n9150 0.00965149
R19143 VSS.n9155 VSS.n9152 0.00965149
R19144 VSS.n9160 VSS.n9159 0.00965149
R19145 VSS.n9164 VSS.n9161 0.00965149
R19146 VSS.n9168 VSS.n9165 0.00965149
R19147 VSS.n11431 VSS.n11428 0.00958201
R19148 VSS.n11459 VSS.n14 0.00949089
R19149 VSS.n11458 VSS.n14 0.00949089
R19150 VSS.n11457 VSS.n15 0.00949089
R19151 VSS.n11456 VSS.n15 0.00949089
R19152 VSS.n11455 VSS.n16 0.00949089
R19153 VSS.n11454 VSS.n16 0.00949089
R19154 VSS.n11453 VSS.n17 0.00949089
R19155 VSS.n11452 VSS.n17 0.00949089
R19156 VSS.n11294 VSS.n23 0.00949089
R19157 VSS.n11443 VSS.n24 0.00949089
R19158 VSS.n11442 VSS.n24 0.00949089
R19159 VSS.n11441 VSS.n25 0.00949089
R19160 VSS.n11440 VSS.n25 0.00949089
R19161 VSS.n11439 VSS.n26 0.00949089
R19162 VSS.n11438 VSS.n26 0.00949089
R19163 VSS.n11437 VSS.n27 0.00949089
R19164 VSS.n11436 VSS.n27 0.00949089
R19165 VSS.n11435 VSS.n28 0.00949089
R19166 VSS.n11434 VSS.n28 0.00949089
R19167 VSS.n11428 VSS.n38 0.00949089
R19168 VSS.n11427 VSS.n38 0.00949089
R19169 VSS.n11426 VSS.n39 0.00949089
R19170 VSS.n11425 VSS.n39 0.00949089
R19171 VSS.n11424 VSS.n40 0.00949089
R19172 VSS.n11423 VSS.n40 0.00949089
R19173 VSS.n11422 VSS.n41 0.00949089
R19174 VSS.n11421 VSS.n41 0.00949089
R19175 VSS.n11420 VSS.n42 0.00949089
R19176 VSS.n11419 VSS.n42 0.00949089
R19177 VSS.n133 VSS.n48 0.00949089
R19178 VSS.n11410 VSS.n49 0.00949089
R19179 VSS.n11409 VSS.n49 0.00949089
R19180 VSS.n11408 VSS.n50 0.00949089
R19181 VSS.n11407 VSS.n50 0.00949089
R19182 VSS.n11406 VSS.n51 0.00949089
R19183 VSS.n11405 VSS.n51 0.00949089
R19184 VSS.n11404 VSS.n52 0.00949089
R19185 VSS.n11403 VSS.n52 0.00949089
R19186 VSS.n11402 VSS.n53 0.00949089
R19187 VSS.n11401 VSS.n53 0.00949089
R19188 VSS.n63 VSS.n3 0.00949089
R19189 VSS.n11310 VSS.n125 0.00947638
R19190 VSS.n900 VSS.n898 0.00936227
R19191 VSS.n897 VSS.n895 0.00936227
R19192 VSS.n894 VSS.n893 0.00936227
R19193 VSS.n890 VSS.n888 0.00936227
R19194 VSS.n887 VSS.n886 0.00936227
R19195 VSS.n1069 VSS.n1067 0.00936227
R19196 VSS.n1066 VSS.n1064 0.00936227
R19197 VSS.n1063 VSS.n397 0.00936227
R19198 VSS.n10173 VSS.n10171 0.00936227
R19199 VSS.n10170 VSS.n10169 0.00936227
R19200 VSS.n10167 VSS.n10166 0.00936227
R19201 VSS.n939 VSS.n937 0.00936227
R19202 VSS.n936 VSS.n934 0.00936227
R19203 VSS.n933 VSS.n325 0.00936227
R19204 VSS.n10233 VSS.n10231 0.00936227
R19205 VSS.n10230 VSS.n10229 0.00936227
R19206 VSS.n10227 VSS.n10226 0.00936227
R19207 VSS.n10908 VSS.n10906 0.00936227
R19208 VSS.n10905 VSS.n10904 0.00936227
R19209 VSS.n10901 VSS.n10899 0.00936227
R19210 VSS.n10898 VSS.n10897 0.00936227
R19211 VSS.n724 VSS.n722 0.00936227
R19212 VSS.n721 VSS.n720 0.00936227
R19213 VSS.n717 VSS.n715 0.00936227
R19214 VSS.n714 VSS.n713 0.00936227
R19215 VSS.n711 VSS.n212 0.00936227
R19216 VSS.n1437 VSS.n1435 0.00936227
R19217 VSS.n1434 VSS.n1433 0.00936227
R19218 VSS.n1231 VSS.n1229 0.00936227
R19219 VSS.n1228 VSS.n1227 0.00936227
R19220 VSS.n1225 VSS.n1219 0.00936227
R19221 VSS.n9269 VSS.n1503 0.00936227
R19222 VSS.n9273 VSS.n9272 0.00936227
R19223 VSS.n9277 VSS.n9274 0.00936227
R19224 VSS.n9282 VSS.n9281 0.00936227
R19225 VSS.n9286 VSS.n9283 0.00936227
R19226 VSS.n9290 VSS.n9287 0.00936227
R19227 VSS.n9056 VSS.n9054 0.00936227
R19228 VSS.n9053 VSS.n9051 0.00936227
R19229 VSS.n9050 VSS.n1530 0.00936227
R19230 VSS.n9122 VSS.n9121 0.00936227
R19231 VSS.n9126 VSS.n9123 0.00936227
R19232 VSS.n9130 VSS.n9127 0.00936227
R19233 VSS.n10840 VSS.n10734 0.0092701
R19234 VSS.n11295 VSS.n18 0.00924789
R19235 VSS.n134 VSS.n43 0.00924789
R19236 VSS.n9885 VSS.n9884 0.00862937
R19237 VSS.n9872 VSS.n673 0.00862937
R19238 VSS.n9519 VSS.n9518 0.00862937
R19239 VSS.n9895 VSS.n9894 0.00862937
R19240 VSS.n9926 VSS.n583 0.00862937
R19241 VSS.n11282 VSS.n22 0.00862937
R19242 VSS.n141 VSS.n47 0.00862937
R19243 VSS.n9617 VSS.n810 0.00862937
R19244 VSS.n778 VSS.n648 0.00852448
R19245 VSS.n9879 VSS.n667 0.00852448
R19246 VSS.n1255 VSS.n1247 0.00852448
R19247 VSS.n9654 VSS.n628 0.00852448
R19248 VSS.n9918 VSS.n597 0.00852448
R19249 VSS.n11043 VSS.n19 0.00852448
R19250 VSS.n9959 VSS.n44 0.00852448
R19251 VSS.n9610 VSS.n9609 0.00852448
R19252 VSS.n9496 VSS.n9493 0.00847863
R19253 VSS.n9886 VSS.n648 0.00847203
R19254 VSS.n9881 VSS.n654 0.00847203
R19255 VSS.n1178 VSS.n679 0.00847203
R19256 VSS.n9879 VSS.n668 0.00847203
R19257 VSS.n9520 VSS.n1255 0.00847203
R19258 VSS.n9893 VSS.n628 0.00847203
R19259 VSS.n9907 VSS.n9906 0.00847203
R19260 VSS.n9904 VSS.n9903 0.00847203
R19261 VSS.n9918 VSS.n9917 0.00847203
R19262 VSS.n11281 VSS.n19 0.00847203
R19263 VSS.n140 VSS.n44 0.00847203
R19264 VSS.n9610 VSS.n815 0.00847203
R19265 VSS.n9884 VSS.n649 0.00836713
R19266 VSS.n9882 VSS.n653 0.00836713
R19267 VSS.n9854 VSS.n9853 0.00836713
R19268 VSS.n9872 VSS.n9871 0.00836713
R19269 VSS.n9518 VSS.n1267 0.00836713
R19270 VSS.n9895 VSS.n641 0.00836713
R19271 VSS.n621 VSS.n620 0.00836713
R19272 VSS.n9698 VSS.n627 0.00836713
R19273 VSS.n9927 VSS.n9926 0.00836713
R19274 VSS.n9947 VSS.n22 0.00836713
R19275 VSS.n11187 VSS.n47 0.00836713
R19276 VSS.n9618 VSS.n9617 0.00836713
R19277 VSS.n9500 VSS.n9499 0.00819275
R19278 VSS.n9492 VSS.n1375 0.00819275
R19279 VSS.n10552 VSS.n10551 0.00799437
R19280 VSS.n10540 VSS.n10539 0.00799437
R19281 VSS.n9469 VSS.n9468 0.00788202
R19282 VSS.n9462 VSS.n9458 0.00780812
R19283 VSS.n9441 VSS.n9440 0.00779878
R19284 VSS.n10839 VSS.n10735 0.00773913
R19285 VSS.n10836 VSS.n10790 0.00773913
R19286 VSS.n10835 VSS.n10790 0.00773913
R19287 VSS.n10829 VSS.n10811 0.00773913
R19288 VSS.n10826 VSS.n10820 0.00773913
R19289 VSS.n9506 VSS.n9505 0.00767297
R19290 VSS.n1339 VSS.n1338 0.00767297
R19291 VSS.n10811 VSS.n10810 0.00761685
R19292 VSS.n10590 VSS.n10589 0.00752176
R19293 VSS.n10490 VSS.n10489 0.00752176
R19294 VSS.n10538 VSS.n10491 0.00752176
R19295 VSS.n10525 VSS.n10524 0.007488
R19296 VSS.n10513 VSS.n10512 0.007488
R19297 VSS.n10741 VSS.n247 0.00721329
R19298 VSS.n10636 VSS.n10635 0.00704376
R19299 VSS.n10760 VSS.n241 0.00704376
R19300 VSS.n10761 VSS.n10760 0.00704376
R19301 VSS.n11384 VSS.n11382 0.00703487
R19302 VSS.n10505 VSS.n10504 0.00701538
R19303 VSS.n10522 VSS.n10506 0.00701538
R19304 VSS.n10521 VSS.n10507 0.00701538
R19305 VSS.n10509 VSS.n10508 0.00701538
R19306 VSS.n10518 VSS.n10517 0.00701538
R19307 VSS.n10516 VSS.n10515 0.00701538
R19308 VSS.n9447 VSS.n9446 0.00681098
R19309 VSS.n10567 VSS.n10556 0.00674846
R19310 VSS.n10570 VSS.n10567 0.00674846
R19311 VSS.n9503 VSS.n9502 0.00671138
R19312 VSS.n1342 VSS.n1341 0.00671138
R19313 VSS.n10484 VSS.n10483 0.00667779
R19314 VSS.n10549 VSS.n10485 0.00667779
R19315 VSS.n10548 VSS.n10486 0.00667779
R19316 VSS.n10488 VSS.n10487 0.00667779
R19317 VSS.n10545 VSS.n10544 0.00667779
R19318 VSS.n10543 VSS.n10542 0.00667779
R19319 VSS.n9434 VSS.n9428 0.00659146
R19320 VSS.n10720 VSS.n10719 0.00658034
R19321 VSS.n10773 VSS.n10772 0.00653147
R19322 VSS.n9504 VSS.n1340 0.00647748
R19323 VSS.n9501 VSS.n1343 0.00639951
R19324 VSS.n10775 VSS.n10774 0.00632168
R19325 VSS.n10732 VSS.n10701 0.00625167
R19326 VSS.n10610 VSS.n10609 0.00619059
R19327 VSS.n10592 VSS.n10482 0.00617142
R19328 VSS.n10527 VSS.n10500 0.00617142
R19329 VSS.n10503 VSS.n10502 0.00617142
R19330 VSS.n10511 VSS.n10510 0.00617142
R19331 VSS.n10348 VSS.n10347 0.00617142
R19332 VSS.n9488 VSS.n9487 0.00616561
R19333 VSS.n10856 VSS.n10855 0.00611189
R19334 VSS.n9490 VSS.n9489 0.00582775
R19335 VSS.n9474 VSS.n1377 0.00582775
R19336 VSS.n10721 VSS.n10720 0.00581345
R19337 VSS.n10825 VSS.n10824 0.00559341
R19338 VSS.n81 VSS.n78 0.00554673
R19339 VSS.n10894 VSS.n10893 0.00554202
R19340 VSS.n11463 VSS.n11462 0.00554202
R19341 VSS.n11462 VSS.n11461 0.00554202
R19342 VSS.n11310 VSS.n127 0.00550787
R19343 VSS.n11102 VSS.n11101 0.005488
R19344 VSS.n11084 VSS.n11080 0.005488
R19345 VSS.n10910 VSS.n10909 0.00547006
R19346 VSS.n11082 VSS.n11081 0.00536194
R19347 VSS.n8954 VSS.n1579 0.00535451
R19348 VSS.n10827 VSS.n10812 0.00529348
R19349 VSS.n10873 VSS.n10872 0.00528992
R19350 VSS.n192 VSS.n191 0.00523684
R19351 VSS.n197 VSS.n196 0.00523684
R19352 VSS.n470 VSS.n469 0.00523684
R19353 VSS.n475 VSS.n474 0.00523684
R19354 VSS.n263 VSS.n262 0.00523684
R19355 VSS.n268 VSS.n267 0.00523684
R19356 VSS.n335 VSS.n334 0.00523684
R19357 VSS.n340 VSS.n339 0.00523684
R19358 VSS.n407 VSS.n406 0.00523684
R19359 VSS.n412 VSS.n411 0.00523684
R19360 VSS.n11099 VSS.n11086 0.00523589
R19361 VSS.n11444 VSS.n23 0.00520807
R19362 VSS.n11411 VSS.n48 0.00520807
R19363 VSS.n1337 VSS.n1336 0.00520401
R19364 VSS.n10060 VSS.n10059 0.00516387
R19365 VSS.n11083 VSS.n11078 0.00516387
R19366 VSS.n11452 VSS.n11451 0.00514732
R19367 VSS.n11419 VSS.n11418 0.00514732
R19368 VSS.n10108 VSS.n10107 0.00512785
R19369 VSS.n450 VSS.n449 0.00512785
R19370 VSS.n10105 VSS.n451 0.00512785
R19371 VSS.n11451 VSS.n18 0.00511694
R19372 VSS.n11418 VSS.n43 0.00511694
R19373 VSS.n538 VSS.n537 0.00507383
R19374 VSS.n10057 VSS.n539 0.00507383
R19375 VSS.n10056 VSS.n540 0.00507383
R19376 VSS.n542 VSS.n541 0.00507383
R19377 VSS.n11444 VSS.n11443 0.00505619
R19378 VSS.n11411 VSS.n11410 0.00505619
R19379 VSS.n1316 VSS.n1315 0.00496579
R19380 VSS.n1297 VSS.n1273 0.00496579
R19381 VSS.n10891 VSS.n10874 0.00492977
R19382 VSS.n10890 VSS.n10889 0.00492977
R19383 VSS.n10888 VSS.n10875 0.00492977
R19384 VSS.n10855 VSS.n10854 0.00490559
R19385 VSS.n10637 VSS.n240 0.00489366
R19386 VSS.n10863 VSS.n241 0.00489366
R19387 VSS.n1296 VSS.n1295 0.00487585
R19388 VSS.n9495 VSS.n9494 0.00486616
R19389 VSS.n9497 VSS.n1345 0.00486616
R19390 VSS.n10834 VSS.n10833 0.00485326
R19391 VSS.n551 VSS.n549 0.00483974
R19392 VSS.n10045 VSS.n10044 0.00483974
R19393 VSS.n11105 VSS.n11104 0.00483974
R19394 VSS.n10100 VSS.n457 0.00482173
R19395 VSS.n10099 VSS.n10098 0.00482173
R19396 VSS.n10097 VSS.n10096 0.00482173
R19397 VSS.n10054 VSS.n10053 0.0047497
R19398 VSS.n186 VSS.n185 0.00469568
R19399 VSS.n11147 VSS.n187 0.00469568
R19400 VSS.n11146 VSS.n11145 0.00469568
R19401 VSS.n10530 VSS.n10498 0.00465229
R19402 VSS.n531 VSS.n530 0.00464166
R19403 VSS.n529 VSS.n528 0.00464166
R19404 VSS.n515 VSS.n514 0.00464166
R19405 VSS.n10061 VSS.n533 0.00464166
R19406 VSS.n10809 VSS.n10808 0.00463315
R19407 VSS.n9491 VSS.n1376 0.00463225
R19408 VSS.n10877 VSS.n10876 0.00460564
R19409 VSS.n10886 VSS.n10885 0.00460564
R19410 VSS.n11336 VSS.n105 0.00455578
R19411 VSS.n11338 VSS.n105 0.00455578
R19412 VSS.n11098 VSS.n11087 0.00455162
R19413 VSS.n11089 VSS.n11088 0.00455162
R19414 VSS.n11096 VSS.n11095 0.00455162
R19415 VSS.n11091 VSS.n11090 0.00455162
R19416 VSS.n11093 VSS.n11092 0.00455162
R19417 VSS.n456 VSS.n455 0.00446158
R19418 VSS.n10064 VSS.n513 0.00446158
R19419 VSS.n10838 VSS.n10789 0.0044375
R19420 VSS.n10638 VSS.n10637 0.00442625
R19421 VSS.n10104 VSS.n452 0.00442557
R19422 VSS.n454 VSS.n453 0.00442557
R19423 VSS.n747 VSS.n726 0.0044234
R19424 VSS.n747 VSS.n746 0.0044234
R19425 VSS.n10838 VSS.n10837 0.00441304
R19426 VSS.n10048 VSS.n10047 0.00440756
R19427 VSS.n11246 VSS.n11245 0.00438136
R19428 VSS.n11229 VSS.n11225 0.00438136
R19429 VSS.n11243 VSS.n11230 0.00438136
R19430 VSS.n10895 VSS.n235 0.00437155
R19431 VSS.n119 VSS.n13 0.00436387
R19432 VSS.n1309 VSS.n1308 0.00433553
R19433 VSS.n1307 VSS.n1306 0.00433553
R19434 VSS.n10854 VSS.n10853 0.00432867
R19435 VSS.n11227 VSS.n11226 0.00428328
R19436 VSS.n10502 VSS.n10500 0.00428095
R19437 VSS.n10525 VSS.n10503 0.00428095
R19438 VSS.n10512 VSS.n10511 0.00428095
R19439 VSS.n10510 VSS.n10346 0.00428095
R19440 VSS.n10655 VSS.n10346 0.00428095
R19441 VSS.n10654 VSS.n10347 0.00428095
R19442 VSS.n1313 VSS.n1311 0.00426351
R19443 VSS.n10535 VSS.n10534 0.00424719
R19444 VSS.n10528 VSS.n10527 0.00424719
R19445 VSS.n10792 VSS.n10791 0.00424185
R19446 VSS.n11055 VSS.n11054 0.00422749
R19447 VSS.n11108 VSS.n11056 0.00422749
R19448 VSS.n11107 VSS.n11057 0.00422749
R19449 VSS.n11059 VSS.n11058 0.00422749
R19450 VSS.n461 VSS.n459 0.00419148
R19451 VSS.n10093 VSS.n10092 0.00419148
R19452 VSS.n478 VSS.n460 0.00419148
R19453 VSS.n553 VSS.n550 0.00413745
R19454 VSS.n10042 VSS.n554 0.00413745
R19455 VSS.n9826 VSS.n9823 0.00412915
R19456 VSS.n11228 VSS.n11223 0.00412915
R19457 VSS.n10103 VSS.n10102 0.00410144
R19458 VSS.n1450 VSS.n1449 0.00410112
R19459 VSS.n1440 VSS.n1439 0.00410112
R19460 VSS.n1447 VSS.n1441 0.00410112
R19461 VSS.n1376 VSS.n1375 0.0040605
R19462 VSS.n9491 VSS.n9490 0.0040605
R19463 VSS.n9825 VSS.n9824 0.00405908
R19464 VSS.n9828 VSS.n765 0.00405908
R19465 VSS.n9831 VSS.n9830 0.00405908
R19466 VSS.n9829 VSS.n764 0.00405908
R19467 VSS.n9195 VSS.n9194 0.00405263
R19468 VSS.n9190 VSS.n9189 0.00405263
R19469 VSS.n9331 VSS.n9330 0.00405263
R19470 VSS.n9326 VSS.n9325 0.00405263
R19471 VSS.n169 VSS.n168 0.00405263
R19472 VSS.n164 VSS.n163 0.00405263
R19473 VSS.n9577 VSS.n9576 0.00405263
R19474 VSS.n9572 VSS.n9571 0.00405263
R19475 VSS.n9028 VSS.n9027 0.00405263
R19476 VSS.n9023 VSS.n9022 0.00405263
R19477 VSS.n544 VSS.n543 0.00404742
R19478 VSS.n10051 VSS.n545 0.00404742
R19479 VSS.n10050 VSS.n10049 0.00404742
R19480 VSS.n10728 VSS.n10703 0.00401077
R19481 VSS.n10730 VSS.n10703 0.00401077
R19482 VSS.n4805 VSS.n1580 0.00400211
R19483 VSS.n10833 VSS.n10791 0.00399728
R19484 VSS.n9388 VSS.n1475 0.00399694
R19485 VSS.n11120 VSS.n11119 0.0039934
R19486 VSS.n11035 VSS.n11034 0.0039934
R19487 VSS.n1473 VSS.n1418 0.00397501
R19488 VSS.n1472 VSS.n1471 0.00397501
R19489 VSS.n448 VSS.n447 0.00395738
R19490 VSS.n745 VSS.n727 0.00394699
R19491 VSS.n729 VSS.n728 0.00394699
R19492 VSS.n743 VSS.n742 0.00394699
R19493 VSS.n11 VSS.n10 0.00392137
R19494 VSS.n11463 VSS.n12 0.00392137
R19495 VSS.n10884 VSS.n10878 0.00390336
R19496 VSS.n10880 VSS.n10879 0.00390336
R19497 VSS.n10883 VSS.n10882 0.00390336
R19498 VSS.n11111 VSS.n11110 0.00390336
R19499 VSS.n697 VSS.n695 0.00387693
R19500 VSS.n761 VSS.n760 0.00387693
R19501 VSS.n11249 VSS.n11248 0.00387693
R19502 VSS.n9599 VSS.n828 0.00386291
R19503 VSS.n830 VSS.n829 0.00386291
R19504 VSS.n9598 VSS.n9597 0.00386291
R19505 VSS.n10776 VSS.n10769 0.00385664
R19506 VSS.n9494 VSS.n1345 0.0038266
R19507 VSS.n9497 VSS.n9496 0.0038266
R19508 VSS.n10041 VSS.n555 0.00381333
R19509 VSS.n557 VSS.n556 0.00381333
R19510 VSS.n9834 VSS.n9833 0.00380687
R19511 VSS.n10074 VSS.n497 0.00379532
R19512 VSS.n11325 VSS.n11324 0.00377731
R19513 VSS.n10551 VSS.n10483 0.00377457
R19514 VSS.n10485 VSS.n10484 0.00377457
R19515 VSS.n10549 VSS.n10548 0.00377457
R19516 VSS.n10487 VSS.n10486 0.00377457
R19517 VSS.n10545 VSS.n10488 0.00377457
R19518 VSS.n10544 VSS.n10543 0.00377457
R19519 VSS.n10542 VSS.n10540 0.00377457
R19520 VSS.n11157 VSS.n11156 0.00376483
R19521 VSS.n11159 VSS.n158 0.00376483
R19522 VSS.n11158 VSS.n177 0.00376483
R19523 VSS.n1301 VSS.n1300 0.00372329
R19524 VSS.n1304 VSS.n1302 0.00372329
R19525 VSS.n9813 VSS.n9812 0.00372279
R19526 VSS.n9811 VSS.n770 0.00372279
R19527 VSS.n9818 VSS.n9817 0.00372279
R19528 VSS.n9821 VSS.n769 0.00372279
R19529 VSS.n1295 VSS.n1282 0.00370748
R19530 VSS.n385 VSS.n384 0.00370748
R19531 VSS.n313 VSS.n300 0.00370748
R19532 VSS.n517 VSS.n503 0.00370528
R19533 VSS.n519 VSS.n518 0.00370528
R19534 VSS.n524 VSS.n521 0.00370528
R19535 VSS.n523 VSS.n522 0.00370528
R19536 VSS.n526 VSS.n516 0.00370528
R19537 VSS.n740 VSS.n739 0.00369477
R19538 VSS.n731 VSS.n730 0.00369477
R19539 VSS.n11129 VSS.n11128 0.00368728
R19540 VSS.n11025 VSS.n11024 0.00368728
R19541 VSS.n119 VSS.n118 0.00367595
R19542 VSS.n9083 VSS.n9082 0.00367572
R19543 VSS.n9391 VSS.n9388 0.00367572
R19544 VSS.n9240 VSS.n9239 0.00367572
R19545 VSS.n11340 VSS.n103 0.00367038
R19546 VSS.n11138 VSS.n11137 0.00366927
R19547 VSS.n203 VSS.n202 0.00366927
R19548 VSS.n11135 VSS.n204 0.00366927
R19549 VSS.n11134 VSS.n11132 0.00366927
R19550 VSS.n11242 VSS.n11231 0.00365273
R19551 VSS.n11233 VSS.n11232 0.00365273
R19552 VSS.n11240 VSS.n11239 0.00365273
R19553 VSS.n11235 VSS.n11234 0.00365273
R19554 VSS.n11237 VSS.n11236 0.00365273
R19555 VSS.n1318 VSS.n1272 0.00365126
R19556 VSS.n10141 VSS.n10140 0.00362264
R19557 VSS.n10201 VSS.n10200 0.00362264
R19558 VSS.n10261 VSS.n10260 0.00362264
R19559 VSS.n11038 VSS.n11036 0.00359724
R19560 VSS.n11305 VSS.n123 0.00359693
R19561 VSS.n11308 VSS.n123 0.00359693
R19562 VSS.n9039 VSS.n1559 0.00359172
R19563 VSS.n9375 VSS.n9374 0.00359172
R19564 VSS.n9206 VSS.n1521 0.00359172
R19565 VSS.n9601 VSS.n9600 0.00358267
R19566 VSS.n9816 VSS.n9815 0.00358267
R19567 VSS.n11117 VSS.n11051 0.00356122
R19568 VSS.n10828 VSS.n10827 0.00355707
R19569 VSS.n1446 VSS.n1442 0.00355465
R19570 VSS.n1444 VSS.n1443 0.00355465
R19571 VSS.n9841 VSS.n9840 0.00354064
R19572 VSS.n10166 VSS.n10164 0.00352395
R19573 VSS.n10226 VSS.n10224 0.00352395
R19574 VSS.n749 VSS.n725 0.00351261
R19575 VSS.n9315 VSS.n1503 0.00349401
R19576 VSS.n9062 VSS.n9056 0.00349401
R19577 VSS.n1468 VSS.n1467 0.00348459
R19578 VSS.n1466 VSS.n1465 0.00348459
R19579 VSS.n1424 VSS.n1423 0.00348459
R19580 VSS.n496 VSS.n495 0.00347119
R19581 VSS.n10076 VSS.n10075 0.00347119
R19582 VSS.n10524 VSS.n10504 0.00343698
R19583 VSS.n10506 VSS.n10505 0.00343698
R19584 VSS.n10522 VSS.n10521 0.00343698
R19585 VSS.n10508 VSS.n10507 0.00343698
R19586 VSS.n10518 VSS.n10509 0.00343698
R19587 VSS.n10517 VSS.n10516 0.00343698
R19588 VSS.n10515 VSS.n10513 0.00343698
R19589 VSS.n499 VSS.n498 0.00343517
R19590 VSS.n11126 VSS.n11027 0.00343517
R19591 VSS.n1470 VSS.n1419 0.00342854
R19592 VSS.n11199 VSS.n11198 0.00340051
R19593 VSS.n11252 VSS.n11200 0.00340051
R19594 VSS.n11251 VSS.n11201 0.00340051
R19595 VSS.n11203 VSS.n11202 0.00340051
R19596 VSS.n1303 VSS.n441 0.00339916
R19597 VSS.n10114 VSS.n442 0.00339916
R19598 VSS.n444 VSS.n443 0.00339916
R19599 VSS.n10112 VSS.n10111 0.00339916
R19600 VSS.n10084 VSS.n10083 0.00339916
R19601 VSS.n9475 VSS.n9474 0.00338478
R19602 VSS.n11022 VSS.n11021 0.00338115
R19603 VSS.n9589 VSS.n9567 0.00337249
R19604 VSS.n9593 VSS.n9592 0.00337249
R19605 VSS.n9588 VSS.n9587 0.00337249
R19606 VSS.n10039 VSS.n10038 0.00334514
R19607 VSS.n1357 VSS.n1356 0.00333232
R19608 VSS.n10019 VSS.n10018 0.00333232
R19609 VSS.n699 VSS.n696 0.00333045
R19610 VSS.n758 VSS.n700 0.00333045
R19611 VSS.n1445 VSS.n827 0.00330243
R19612 VSS.n9440 VSS.n9439 0.00329878
R19613 VSS.n11122 VSS.n11031 0.00329112
R19614 VSS.n11033 VSS.n11032 0.00329112
R19615 VSS.n9476 VSS.n9475 0.00328083
R19616 VSS.n493 VSS.n492 0.00327311
R19617 VSS.n10081 VSS.n10080 0.00327311
R19618 VSS.n10079 VSS.n10078 0.00327311
R19619 VSS.n495 VSS.n494 0.00327311
R19620 VSS.n9836 VSS.n9835 0.00326039
R19621 VSS.n9838 VSS.n763 0.00326039
R19622 VSS.n9837 VSS.n692 0.00326039
R19623 VSS.n10111 VSS.n10110 0.0032551
R19624 VSS.n447 VSS.n446 0.0032551
R19625 VSS.n10089 VSS.n484 0.0032551
R19626 VSS.n486 VSS.n485 0.0032551
R19627 VSS.n10087 VSS.n10086 0.0032551
R19628 VSS.n489 VSS.n488 0.0032551
R19629 VSS.n10084 VSS.n490 0.0032551
R19630 VSS.n11267 VSS.n11180 0.00321836
R19631 VSS.n11182 VSS.n11181 0.00321836
R19632 VSS.n10831 VSS.n10830 0.00321467
R19633 VSS.n11053 VSS.n11052 0.00320108
R19634 VSS.n11115 VSS.n11114 0.00320108
R19635 VSS.n11113 VSS.n11112 0.00320108
R19636 VSS.n1438 VSS.n1429 0.00319033
R19637 VSS.n10533 VSS.n10532 0.00316692
R19638 VSS.n10025 VSS.n10024 0.00316322
R19639 VSS.n11340 VSS.n11339 0.00315277
R19640 VSS.n737 VSS.n732 0.0031483
R19641 VSS.n736 VSS.n735 0.0031483
R19642 VSS.n734 VSS.n733 0.0031483
R19643 VSS.n11255 VSS.n11254 0.0031483
R19644 VSS.n10832 VSS.n10809 0.0031413
R19645 VSS.n10638 VSS.n10635 0.0031175
R19646 VSS.n10535 VSS.n10492 0.0030994
R19647 VSS.n11433 VSS.n31 0.00308184
R19648 VSS.n10024 VSS.n573 0.00307868
R19649 VSS.n757 VSS.n701 0.00307823
R19650 VSS.n703 VSS.n702 0.00307823
R19651 VSS.n492 VSS.n491 0.00307503
R19652 VSS.n10072 VSS.n10071 0.00307503
R19653 VSS.n501 VSS.n500 0.00307503
R19654 VSS.n10070 VSS.n502 0.00307503
R19655 VSS.n11125 VSS.n11028 0.00307503
R19656 VSS.n11030 VSS.n11029 0.00307503
R19657 VSS.n9495 VSS.n1344 0.00307291
R19658 VSS.n9793 VSS.n9792 0.00306422
R19659 VSS.n11131 VSS.n205 0.00305702
R19660 VSS.n1463 VSS.n1425 0.00300817
R19661 VSS.n4806 VSS.n4805 0.00300278
R19662 VSS.n9803 VSS.n9802 0.00299416
R19663 VSS.n9801 VSS.n772 0.00299416
R19664 VSS.n9808 VSS.n9805 0.00299416
R19665 VSS.n9807 VSS.n9806 0.00299416
R19666 VSS.n9810 VSS.n771 0.00299416
R19667 VSS.n11132 VSS.n11131 0.00298499
R19668 VSS.n11021 VSS.n205 0.00298499
R19669 VSS.n11276 VSS.n152 0.00298015
R19670 VSS.n11173 VSS.n11172 0.00298015
R19671 VSS.n11274 VSS.n11273 0.00298015
R19672 VSS.n10083 VSS.n491 0.00296699
R19673 VSS.n10071 VSS.n500 0.00296699
R19674 VSS.n502 VSS.n501 0.00296699
R19675 VSS.n11126 VSS.n11125 0.00296699
R19676 VSS.n11029 VSS.n11028 0.00296699
R19677 VSS.n11123 VSS.n11030 0.00296699
R19678 VSS.n11163 VSS.n11162 0.00296614
R19679 VSS.n11165 VSS.n11164 0.00296614
R19680 VSS.n11168 VSS.n155 0.00296614
R19681 VSS.n10604 VSS.n10441 0.00296504
R19682 VSS.n1416 VSS.n1403 0.00295213
R19683 VSS.n10587 VSS.n10482 0.00293061
R19684 VSS.n10591 VSS.n10590 0.00293061
R19685 VSS.n10589 VSS.n10552 0.00293061
R19686 VSS.n10539 VSS.n10489 0.00293061
R19687 VSS.n10491 VSS.n10490 0.00293061
R19688 VSS.n11461 VSS.n11460 0.00291297
R19689 VSS.n11265 VSS.n11264 0.00291009
R19690 VSS.n1358 VSS.n1357 0.00290958
R19691 VSS.n10020 VSS.n10019 0.00290958
R19692 VSS.n11261 VSS.n11195 0.00288206
R19693 VSS.n9035 VSS.n9034 0.00288205
R19694 VSS.n10148 VSS.n10147 0.00288205
R19695 VSS.n10208 VSS.n10207 0.00288205
R19696 VSS.n10268 VSS.n10267 0.00288205
R19697 VSS.n9340 VSS.n9339 0.00288205
R19698 VSS.n9202 VSS.n9201 0.00288205
R19699 VSS.n10090 VSS.n483 0.00287695
R19700 VSS.n11141 VSS.n11139 0.00287695
R19701 VSS.n10832 VSS.n10831 0.00287228
R19702 VSS.n9489 VSS.n1377 0.002865
R19703 VSS.n10440 VSS.n10335 0.00286014
R19704 VSS.n11115 VSS.n11053 0.00284094
R19705 VSS.n11114 VSS.n11113 0.00284094
R19706 VSS.n11112 VSS.n11111 0.00284094
R19707 VSS.n10046 VSS.n548 0.00282293
R19708 VSS.n9791 VSS.n789 0.002812
R19709 VSS.n9790 VSS.n787 0.002812
R19710 VSS.n11460 VSS.n13 0.00280492
R19711 VSS.n8952 VSS.n8951 0.00280297
R19712 VSS.n4803 VSS.n2503 0.00280297
R19713 VSS.n10788 VSS.n10735 0.00279891
R19714 VSS.n10110 VSS.n446 0.00278691
R19715 VSS.n485 VSS.n484 0.00278691
R19716 VSS.n10086 VSS.n488 0.00278691
R19717 VSS.n490 VSS.n489 0.00278691
R19718 VSS.n788 VSS.n786 0.00278398
R19719 VSS.n10081 VSS.n493 0.00276891
R19720 VSS.n10080 VSS.n10079 0.00276891
R19721 VSS.n10078 VSS.n494 0.00276891
R19722 VSS.n1462 VSS.n1461 0.00275596
R19723 VSS.n1456 VSS.n1455 0.00275596
R19724 VSS.n1459 VSS.n1427 0.00275596
R19725 VSS.n9780 VSS.n9779 0.00275596
R19726 VSS.n11123 VSS.n11122 0.0027509
R19727 VSS.n11032 VSS.n11031 0.0027509
R19728 VSS.n11120 VSS.n11033 0.0027509
R19729 VSS.n154 VSS.n151 0.00274194
R19730 VSS.n9507 VSS.n1336 0.00273506
R19731 VSS.n11321 VSS.n117 0.00273289
R19732 VSS.n11178 VSS.n11177 0.00267188
R19733 VSS.n11268 VSS.n11179 0.00267188
R19734 VSS.n11431 VSS.n36 0.00266998
R19735 VSS.n57 VSS.n54 0.00266998
R19736 VSS.n11398 VSS.n11395 0.00266998
R19737 VSS.n11429 VSS.n36 0.00266998
R19738 VSS.n11400 VSS.n54 0.00266998
R19739 VSS.n11395 VSS.n57 0.00266998
R19740 VSS.n10035 VSS.n10034 0.00266086
R19741 VSS.n9783 VSS.n9782 0.00265787
R19742 VSS.n9785 VSS.n9784 0.00265787
R19743 VSS.n9788 VSS.n790 0.00265787
R19744 VSS.n9787 VSS.n789 0.00265787
R19745 VSS.n10776 VSS.n10775 0.00265035
R19746 VSS.n10742 VSS.n10741 0.00265035
R19747 VSS.n10910 VSS.n228 0.0026461
R19748 VSS.n10913 VSS.n228 0.0026461
R19749 VSS.n1453 VSS.n1452 0.00264386
R19750 VSS.n1429 VSS.n1428 0.00264386
R19751 VSS.n9772 VSS.n9771 0.00264386
R19752 VSS.n9770 VSS.n9769 0.00264386
R19753 VSS.n9777 VSS.n795 0.00264386
R19754 VSS.n9776 VSS.n9775 0.00264386
R19755 VSS.n443 VSS.n442 0.00264286
R19756 VSS.n10112 VSS.n444 0.00264286
R19757 VSS.n487 VSS.n486 0.00260684
R19758 VSS.n10072 VSS.n499 0.00260684
R19759 VSS.n754 VSS.n753 0.00260182
R19760 VSS.n705 VSS.n704 0.00260182
R19761 VSS.n751 VSS.n706 0.00260182
R19762 VSS.n11197 VSS.n11196 0.00260182
R19763 VSS.n11259 VSS.n11258 0.00260182
R19764 VSS.n11257 VSS.n11256 0.00260182
R19765 VSS.n10076 VSS.n496 0.00257083
R19766 VSS.n11387 VSS.n81 0.00257045
R19767 VSS.n1454 VSS.n1453 0.00255979
R19768 VSS.n10829 VSS.n10828 0.00252989
R19769 VSS.n9488 VSS.n9476 0.00252714
R19770 VSS.n1298 VSS.n433 0.00251681
R19771 VSS.n462 VSS.n458 0.00251681
R19772 VSS.n10069 VSS.n503 0.00251681
R19773 VSS.n552 VSS.n548 0.00251681
R19774 VSS.n11150 VSS.n11149 0.00251681
R19775 VSS.n11466 VSS.n11465 0.00251681
R19776 VSS.n9782 VSS.n9781 0.00250374
R19777 VSS.n9798 VSS.n9795 0.00250374
R19778 VSS.n9797 VSS.n9796 0.00250374
R19779 VSS.n9799 VSS.n773 0.00250374
R19780 VSS.n11175 VSS.n11174 0.00250374
R19781 VSS.n11271 VSS.n11176 0.00250374
R19782 VSS.n156 VSS.n153 0.00248972
R19783 VSS.n11171 VSS.n11170 0.00248972
R19784 VSS.n11023 VSS.n11022 0.00248079
R19785 VSS.n11052 VSS.n11051 0.00248079
R19786 VSS.n10115 VSS.n441 0.00246279
R19787 VSS.n10090 VSS.n10089 0.00246279
R19788 VSS.n9779 VSS.n794 0.00244769
R19789 VSS.n11171 VSS.n153 0.00243368
R19790 VSS.n11170 VSS.n154 0.00243368
R19791 VSS.n9781 VSS.n9780 0.00241966
R19792 VSS.n9798 VSS.n9797 0.00241966
R19793 VSS.n9796 VSS.n773 0.00241966
R19794 VSS.n11273 VSS.n11174 0.00241966
R19795 VSS.n11176 VSS.n11175 0.00241966
R19796 VSS.n11271 VSS.n11270 0.00241966
R19797 VSS.n10655 VSS.n10654 0.00239047
R19798 VSS.n11137 VSS.n202 0.00237275
R19799 VSS.n204 VSS.n203 0.00237275
R19800 VSS.n11135 VSS.n11134 0.00237275
R19801 VSS.n11128 VSS.n11024 0.00235474
R19802 VSS.n11026 VSS.n11025 0.00235474
R19803 VSS.n9583 VSS.n796 0.0023496
R19804 VSS.n11161 VSS.n157 0.0023496
R19805 VSS.n518 VSS.n517 0.00233673
R19806 VSS.n521 VSS.n519 0.00233673
R19807 VSS.n524 VSS.n523 0.00233673
R19808 VSS.n522 VSS.n516 0.00233673
R19809 VSS.n753 VSS.n704 0.00232158
R19810 VSS.n706 VSS.n705 0.00232158
R19811 VSS.n11259 VSS.n11197 0.00232158
R19812 VSS.n11258 VSS.n11257 0.00232158
R19813 VSS.n11256 VSS.n11255 0.00232158
R19814 VSS.n1312 VSS.n433 0.00231873
R19815 VSS.n1302 VSS.n1301 0.00231873
R19816 VSS.n1304 VSS.n1303 0.00231873
R19817 VSS.n11150 VSS.n184 0.00231873
R19818 VSS.n11322 VSS.n11321 0.00231873
R19819 VSS.n762 VSS.n694 0.00230757
R19820 VSS.n1343 VSS.n1342 0.00229324
R19821 VSS.n9501 VSS.n9500 0.00229324
R19822 VSS.n1452 VSS.n1428 0.00227954
R19823 VSS.n9771 VSS.n9770 0.00227954
R19824 VSS.n9777 VSS.n9776 0.00227954
R19825 VSS.n9775 VSS.n9774 0.00227954
R19826 VSS.n10574 VSS.n10556 0.00227907
R19827 VSS.n9785 VSS.n9783 0.00226553
R19828 VSS.n9784 VSS.n790 0.00226553
R19829 VSS.n9788 VSS.n9787 0.00226553
R19830 VSS.n10037 VSS.n236 0.00226471
R19831 VSS.n11270 VSS.n11177 0.00225152
R19832 VSS.n11179 VSS.n11178 0.00225152
R19833 VSS.n11268 VSS.n11267 0.00225152
R19834 VSS.n10075 VSS.n10074 0.0022467
R19835 VSS.n498 VSS.n497 0.0022467
R19836 VSS.n10857 VSS.n246 0.00223077
R19837 VSS.n556 VSS.n555 0.00222869
R19838 VSS.n10039 VSS.n557 0.00222869
R19839 VSS.n1340 VSS.n1339 0.00221528
R19840 VSS.n9504 VSS.n9503 0.00221528
R19841 VSS.n11093 VSS.n9 0.00219268
R19842 VSS.n751 VSS.n750 0.00218146
R19843 VSS.n10095 VSS.n458 0.00217467
R19844 VSS.n1455 VSS.n1427 0.00216745
R19845 VSS.n1459 VSS.n1458 0.00216745
R19846 VSS.n10870 VSS.n10869 0.00215666
R19847 VSS.n9769 VSS.n9768 0.00213942
R19848 VSS.n9795 VSS.n786 0.00213942
R19849 VSS.n10885 VSS.n10884 0.00213866
R19850 VSS.n10879 VSS.n10878 0.00213866
R19851 VSS.n10883 VSS.n10880 0.00213866
R19852 VSS.n10035 VSS.n560 0.00212065
R19853 VSS.n11118 VSS.n11117 0.00212065
R19854 VSS.n11465 VSS.n10 0.00212065
R19855 VSS.n12 VSS.n11 0.00212065
R19856 VSS.n9791 VSS.n9790 0.0021114
R19857 VSS.n10537 VSS.n10492 0.00208665
R19858 VSS.n10108 VSS.n448 0.00208463
R19859 VSS.n1422 VSS.n1421 0.00206936
R19860 VSS.n9590 VSS.n9566 0.00206936
R19861 VSS.n9803 VSS.n9800 0.00206936
R19862 VSS.n698 VSS.n694 0.00206936
R19863 VSS.n11155 VSS.n11154 0.00206936
R19864 VSS.n11139 VSS.n11138 0.00204862
R19865 VSS.n11119 VSS.n11034 0.00204862
R19866 VSS.n11036 VSS.n11035 0.00204862
R19867 VSS.n11277 VSS.n151 0.00204134
R19868 VSS.n11196 VSS.n11195 0.00204134
R19869 VSS.n1461 VSS.n1426 0.00202732
R19870 VSS.n9772 VSS.n796 0.00202732
R19871 VSS.n10053 VSS.n543 0.0019946
R19872 VSS.n545 VSS.n544 0.0019946
R19873 VSS.n10051 VSS.n10050 0.0019946
R19874 VSS.n9502 VSS.n1341 0.00198137
R19875 VSS.n10921 VSS.n223 0.00196707
R19876 VSS.n11165 VSS.n11163 0.00195726
R19877 VSS.n11164 VSS.n155 0.00195726
R19878 VSS.n11168 VSS.n11167 0.00195726
R19879 VSS.n9499 VSS.n9498 0.00195539
R19880 VSS.n11172 VSS.n152 0.00194325
R19881 VSS.n11274 VSS.n11173 0.00194325
R19882 VSS.n1370 VSS.n1369 0.00193729
R19883 VSS.n9634 VSS.n9633 0.00193729
R19884 VSS.n9745 VSS.n9744 0.00193729
R19885 VSS.n9723 VSS.n9722 0.00193729
R19886 VSS.n10008 VSS.n10007 0.00193729
R19887 VSS.n9986 VSS.n9985 0.00193729
R19888 VSS.n9802 VSS.n9801 0.00192924
R19889 VSS.n9805 VSS.n772 0.00192924
R19890 VSS.n9808 VSS.n9807 0.00192924
R19891 VSS.n9806 VSS.n771 0.00192924
R19892 VSS.n10868 VSS.n10867 0.00192857
R19893 VSS.n11315 VSS.n109 0.00192857
R19894 VSS.n11389 VSS.n62 0.00192857
R19895 VSS.n11393 VSS.n56 0.00192857
R19896 VSS.n11319 VSS.n120 0.00192857
R19897 VSS.n11432 VSS.n34 0.00192857
R19898 VSS.n10707 VSS.n10706 0.00192857
R19899 VSS.n10499 VSS.n10493 0.00192857
R19900 VSS.n11313 VSS.n122 0.00192857
R19901 VSS.n10565 VSS.n10563 0.00192857
R19902 VSS.n10865 VSS.n229 0.00192857
R19903 VSS.n10096 VSS.n10095 0.00192257
R19904 VSS.n10820 VSS.n10819 0.00191848
R19905 VSS.n9468 VSS.n9467 0.00191573
R19906 VSS.n1421 VSS.n1420 0.00191523
R19907 VSS.n1425 VSS.n1424 0.00191523
R19908 VSS.n1463 VSS.n1462 0.00191523
R19909 VSS.n11154 VSS.n178 0.00191523
R19910 VSS.n10044 VSS.n550 0.00190456
R19911 VSS.n554 VSS.n553 0.00190456
R19912 VSS.n10042 VSS.n10041 0.00190456
R19913 VSS.n11466 VSS.n9 0.00190456
R19914 VSS.n9463 VSS.n9462 0.00190156
R19915 VSS.n9793 VSS.n787 0.00185918
R19916 VSS.n9792 VSS.n788 0.00185918
R19917 VSS.n462 VSS.n461 0.00185054
R19918 VSS.n10093 VSS.n459 0.00185054
R19919 VSS.n10092 VSS.n460 0.00185054
R19920 VSS.n11325 VSS.n116 0.00185054
R19921 VSS.n10592 VSS.n10591 0.00185034
R19922 VSS.n702 VSS.n701 0.00184517
R19923 VSS.n755 VSS.n703 0.00184517
R19924 VSS.n10531 VSS.n10530 0.00181658
R19925 VSS.n1318 VSS.n1317 0.00181453
R19926 VSS.n11110 VSS.n11054 0.00181453
R19927 VSS.n11056 VSS.n11055 0.00181453
R19928 VSS.n11108 VSS.n11107 0.00181453
R19929 VSS.n11058 VSS.n11057 0.00181453
R19930 VSS.n11105 VSS.n11059 0.00181453
R19931 VSS.n9595 VSS.n9566 0.00180313
R19932 VSS.n9102 VSS.n9100 0.00180205
R19933 VSS.n861 VSS.n860 0.00180205
R19934 VSS.n1107 VSS.n1106 0.00180205
R19935 VSS.n1049 VSS.n926 0.00180205
R19936 VSS.n1000 VSS.n999 0.00180205
R19937 VSS.n11353 VSS.n100 0.00180205
R19938 VSS.n11369 VSS.n88 0.00180205
R19939 VSS.n1199 VSS.n1198 0.00180205
R19940 VSS.n9414 VSS.n9413 0.00180205
R19941 VSS.n9257 VSS.n1511 0.00180205
R19942 VSS.n11339 VSS.n11338 0.00179403
R19943 VSS.n1311 VSS.n1297 0.00177851
R19944 VSS.n1313 VSS.n1312 0.00177851
R19945 VSS.n10882 VSS.n184 0.00177851
R19946 VSS.n732 VSS.n731 0.00177511
R19947 VSS.n737 VSS.n736 0.00177511
R19948 VSS.n735 VSS.n734 0.00177511
R19949 VSS.n9002 VSS.n9001 0.00176761
R19950 VSS.n1134 VSS.n1131 0.00176761
R19951 VSS.n1082 VSS.n913 0.00176761
R19952 VSS.n1033 VSS.n1032 0.00176761
R19953 VSS.n975 VSS.n952 0.00176761
R19954 VSS.n11002 VSS.n10999 0.00176761
R19955 VSS.n10974 VSS.n10973 0.00176761
R19956 VSS.n9550 VSS.n9548 0.00176761
R19957 VSS.n9357 VSS.n9355 0.00176761
R19958 VSS.n9169 VSS.n9168 0.00176761
R19959 VSS.n11262 VSS.n11261 0.00176109
R19960 VSS.n10744 VSS.n10743 0.00175874
R19961 VSS.n1450 VSS.n1438 0.00173307
R19962 VSS.n1119 VSS.n900 0.00172754
R19963 VSS.n1070 VSS.n1069 0.00172754
R19964 VSS.n1012 VSS.n939 0.00172754
R19965 VSS.n10921 VSS.n10915 0.00172754
R19966 VSS.n10937 VSS.n212 0.00172754
R19967 VSS.n9535 VSS.n1219 0.00172754
R19968 VSS.n9291 VSS.n9290 0.00172754
R19969 VSS.n9131 VSS.n9130 0.00172754
R19970 VSS.n1309 VSS.n1298 0.00170648
R19971 VSS.n1308 VSS.n1307 0.00170648
R19972 VSS.n1306 VSS.n1299 0.00170648
R19973 VSS.n11162 VSS.n11161 0.00170504
R19974 VSS.n11181 VSS.n11180 0.00170504
R19975 VSS.n11265 VSS.n11182 0.00170504
R19976 VSS.n558 VSS.n237 0.00168848
R19977 VSS.n10806 VSS.n10804 0.00168421
R19978 VSS.n10800 VSS.n10798 0.00168421
R19979 VSS.n10630 VSS.n10629 0.00168421
R19980 VSS.n10626 VSS.n10625 0.00168421
R19981 VSS.n10621 VSS.n10620 0.00168421
R19982 VSS.n10617 VSS.n10616 0.00168421
R19983 VSS.n10385 VSS.n10384 0.00168421
R19984 VSS.n10381 VSS.n10380 0.00168421
R19985 VSS.n10376 VSS.n10375 0.00168421
R19986 VSS.n10302 VSS.n10299 0.00168421
R19987 VSS.n10681 VSS.n10297 0.00168421
R19988 VSS.n10684 VSS.n10294 0.00168421
R19989 VSS.n9813 VSS.n9810 0.00167702
R19990 VSS.n10837 VSS.n10836 0.00167391
R19991 VSS.n10826 VSS.n10825 0.00167391
R19992 VSS.n10895 VSS.n10894 0.00167047
R19993 VSS.n9836 VSS.n9834 0.00166301
R19994 VSS.n9835 VSS.n763 0.00166301
R19995 VSS.n9838 VSS.n9837 0.00166301
R19996 VSS.n559 VSS.n558 0.00165246
R19997 VSS.n10049 VSS.n10048 0.00163445
R19998 VSS.n10105 VSS.n10104 0.00161645
R19999 VSS.n453 VSS.n452 0.00161645
R20000 VSS.n10103 VSS.n454 0.00161645
R20001 VSS.n201 VSS.n188 0.00161645
R20002 VSS.n9597 VSS.n9595 0.00160696
R20003 VSS.n11142 VSS.n201 0.00159844
R20004 VSS.n760 VSS.n696 0.00159295
R20005 VSS.n700 VSS.n699 0.00159295
R20006 VSS.n758 VSS.n757 0.00159295
R20007 VSS.n10102 VSS.n455 0.00158043
R20008 VSS.n560 VSS.n559 0.00158043
R20009 VSS.n10766 VSS.n10765 0.00156599
R20010 VSS.n10762 VSS.n10761 0.00155167
R20011 VSS.n9590 VSS.n9589 0.00155091
R20012 VSS.n9593 VSS.n9567 0.00155091
R20013 VSS.n9592 VSS.n9588 0.00155091
R20014 VSS.n10869 VSS.n237 0.00154442
R20015 VSS.n10819 VSS.n10812 0.00152717
R20016 VSS.n1417 VSS.n1416 0.00152289
R20017 VSS.n11254 VSS.n11198 0.00152289
R20018 VSS.n11200 VSS.n11199 0.00152289
R20019 VSS.n11252 VSS.n11251 0.00152289
R20020 VSS.n11202 VSS.n11201 0.00152289
R20021 VSS.n9584 VSS.n9581 0.00150887
R20022 VSS.n10789 VSS.n10788 0.00150272
R20023 VSS.n1471 VSS.n1470 0.00149486
R20024 VSS.n1420 VSS.n1419 0.00149486
R20025 VSS.n733 VSS.n178 0.00149486
R20026 VSS.n11088 VSS.n11087 0.0014904
R20027 VSS.n11096 VSS.n11089 0.0014904
R20028 VSS.n11095 VSS.n11090 0.0014904
R20029 VSS.n11092 VSS.n11091 0.0014904
R20030 VSS.n118 VSS.n117 0.0014904
R20031 VSS.n1468 VSS.n1422 0.00143881
R20032 VSS.n1467 VSS.n1466 0.00143881
R20033 VSS.n1465 VSS.n1423 0.00143881
R20034 VSS.n10886 VSS.n10877 0.00143638
R20035 VSS.n466 VSS.n465 0.00141837
R20036 VSS.n726 VSS.n725 0.00141079
R20037 VSS.n531 VSS.n527 0.00140036
R20038 VSS.n530 VSS.n529 0.00140036
R20039 VSS.n528 VSS.n513 0.00140036
R20040 VSS.n10063 VSS.n514 0.00140036
R20041 VSS.n533 VSS.n515 0.00140036
R20042 VSS.n10754 VSS.n10746 0.00139161
R20043 VSS.n9841 VSS.n692 0.00138277
R20044 VSS.n1447 VSS.n1446 0.00136875
R20045 VSS.n1443 VSS.n1442 0.00136875
R20046 VSS.n1445 VSS.n1444 0.00136875
R20047 VSS.n173 VSS.n159 0.00136875
R20048 VSS.n174 VSS.n173 0.00135474
R20049 VSS.n1388 VSS.n1385 0.00135106
R20050 VSS.n1331 VSS.n1330 0.00135106
R20051 VSS.n11149 VSS.n185 0.00134634
R20052 VSS.n187 VSS.n186 0.00134634
R20053 VSS.n11147 VSS.n11146 0.00134634
R20054 VSS.n10538 VSS.n10537 0.00134396
R20055 VSS.n9601 VSS.n827 0.00134073
R20056 VSS.n11303 VSS.n129 0.00130178
R20057 VSS.n10844 VSS.n10698 0.00130178
R20058 VSS.n10853 VSS.n247 0.00128671
R20059 VSS.n11237 VSS.n0 0.00128468
R20060 VSS.n10047 VSS.n10046 0.00127431
R20061 VSS.n11232 VSS.n11231 0.00127067
R20062 VSS.n11240 VSS.n11233 0.00127067
R20063 VSS.n11239 VSS.n11234 0.00127067
R20064 VSS.n11236 VSS.n11235 0.00127067
R20065 VSS.n11429 VSS.n31 0.00125937
R20066 VSS.n1337 VSS.n1335 0.00125368
R20067 VSS.n9507 VSS.n9506 0.00125368
R20068 VSS.n9498 VSS.n1344 0.00125368
R20069 VSS.n10835 VSS.n10834 0.0012337
R20070 VSS.n739 VSS.n730 0.00122863
R20071 VSS.n457 VSS.n456 0.00122029
R20072 VSS.n10100 VSS.n10099 0.00122029
R20073 VSS.n10098 VSS.n10097 0.00122029
R20074 VSS.n9581 VSS.n9568 0.00121462
R20075 VSS.n10666 VSS.n10665 0.0012124
R20076 VSS.n10428 VSS.n10427 0.0012124
R20077 VSS.n10465 VSS.n10464 0.00121146
R20078 VSS.n552 VSS.n551 0.00120228
R20079 VSS.n10045 VSS.n549 0.00120228
R20080 VSS.n9812 VSS.n9811 0.00120061
R20081 VSS.n9815 VSS.n770 0.00120061
R20082 VSS.n9819 VSS.n9818 0.00120061
R20083 VSS.n9817 VSS.n769 0.00120061
R20084 VSS.n464 VSS.n463 0.00118427
R20085 VSS.n11099 VSS.n11098 0.00116627
R20086 VSS.n11157 VSS.n11155 0.00115857
R20087 VSS.n11156 VSS.n158 0.00115857
R20088 VSS.n11159 VSS.n11158 0.00115857
R20089 VSS.n10586 VSS.n10585 0.0011338
R20090 VSS.n1300 VSS.n1299 0.00111224
R20091 VSS.n465 VSS.n464 0.00111224
R20092 VSS.n527 VSS.n526 0.00111224
R20093 VSS.n10874 VSS.n10873 0.00111224
R20094 VSS.n10891 VSS.n10890 0.00111224
R20095 VSS.n10889 VSS.n10888 0.00111224
R20096 VSS.n10876 VSS.n10875 0.00111224
R20097 VSS.n9840 VSS.n762 0.00110252
R20098 VSS.n10915 VSS.n10913 0.0010988
R20099 VSS.n1364 VSS.n1363 0.00109183
R20100 VSS.n9761 VSS.n9760 0.00109183
R20101 VSS.n9739 VSS.n9738 0.00109183
R20102 VSS.n10027 VSS.n10026 0.00109183
R20103 VSS.n10002 VSS.n10001 0.00109183
R20104 VSS.n9980 VSS.n9979 0.00109183
R20105 VSS.n11387 VSS.n11382 0.00108231
R20106 VSS.n1296 VSS.n1272 0.00107623
R20107 VSS.n1317 VSS.n1316 0.00107623
R20108 VSS.n1315 VSS.n1273 0.00107623
R20109 VSS.n10870 VSS.n236 0.00107623
R20110 VSS.n9600 VSS.n9599 0.00106049
R20111 VSS.n829 VSS.n828 0.00106049
R20112 VSS.n9598 VSS.n830 0.00106049
R20113 VSS.n11317 VSS.n59 0.00104767
R20114 VSS.n698 VSS.n697 0.00104647
R20115 VSS.n761 VSS.n695 0.00104647
R20116 VSS.n11249 VSS.n11204 0.00104647
R20117 VSS.n10070 VSS.n10069 0.00102221
R20118 VSS.n10061 VSS.n10060 0.00102221
R20119 VSS.n9505 VSS.n1338 0.00101978
R20120 VSS.n11243 VSS.n11242 0.00101845
R20121 VSS.n10733 VSS.n10732 0.000993001
R20122 VSS.n755 VSS.n754 0.000976413
R20123 VSS.n746 VSS.n745 0.000976413
R20124 VSS.n728 VSS.n727 0.000976413
R20125 VSS.n743 VSS.n729 0.000976413
R20126 VSS.n742 VSS.n740 0.000976413
R20127 VSS.n11167 VSS.n156 0.000976413
R20128 VSS.n11204 VSS.n11203 0.000976413
R20129 VSS.n10059 VSS.n537 0.000968187
R20130 VSS.n539 VSS.n538 0.000968187
R20131 VSS.n10057 VSS.n10056 0.000968187
R20132 VSS.n541 VSS.n540 0.000968187
R20133 VSS.n10054 VSS.n542 0.000968187
R20134 VSS.n10038 VSS.n10037 0.000968187
R20135 VSS.n1475 VSS.n1403 0.000948389
R20136 VSS.n1418 VSS.n1417 0.000948389
R20137 VSS.n1473 VSS.n1472 0.000948389
R20138 VSS.n10534 VSS.n10533 0.00093886
R20139 VSS.n1366 VSS.n1349 0.000922734
R20140 VSS.n9764 VSS.n9763 0.000922734
R20141 VSS.n9741 VSS.n9666 0.000922734
R20142 VSS.n10030 VSS.n10029 0.000922734
R20143 VSS.n10004 VSS.n147 0.000922734
R20144 VSS.n9982 VSS.n138 0.000922734
R20145 VSS.n10758 VSS.n10757 0.000920842
R20146 VSS.n9887 VSS.n647 0.00091958
R20147 VSS.n1176 VSS.n1175 0.00091958
R20148 VSS.n1180 VSS.n1174 0.00091958
R20149 VSS.n672 VSS.n671 0.00091958
R20150 VSS.n9521 VSS.n1236 0.00091958
R20151 VSS.n9892 VSS.n643 0.00091958
R20152 VSS.n624 VSS.n623 0.00091958
R20153 VSS.n626 VSS.n625 0.00091958
R20154 VSS.n9916 VSS.n9915 0.00091958
R20155 VSS.n11284 VSS.n11283 0.00091958
R20156 VSS.n143 VSS.n142 0.00091958
R20157 VSS.n1234 VSS.n1233 0.00091958
R20158 VSS.n10107 VSS.n449 0.000914166
R20159 VSS.n451 VSS.n450 0.000914166
R20160 VSS.n479 VSS.n478 0.000914166
R20161 VSS.n11145 VSS.n11144 0.000914166
R20162 VSS.n11322 VSS.n116 0.000914166
R20163 VSS.n9800 VSS.n9799 0.000906352
R20164 VSS.n11118 VSS.n11038 0.000896158
R20165 VSS.n10808 VSS.n10793 0.000866848
R20166 VSS.n9826 VSS.n9825 0.000864316
R20167 VSS.n9824 VSS.n765 0.000864316
R20168 VSS.n9831 VSS.n9828 0.000864316
R20169 VSS.n9830 VSS.n9829 0.000864316
R20170 VSS.n9833 VSS.n764 0.000864316
R20171 VSS.n11104 VSS.n11078 0.00082413
R20172 VSS.n1449 VSS.n1439 0.000822279
R20173 VSS.n1441 VSS.n1440 0.000822279
R20174 VSS.n9587 VSS.n9586 0.000822279
R20175 VSS.n177 VSS.n176 0.000822279
R20176 VSS.n11264 VSS.n11262 0.000808267
R20177 VSS.n10730 VSS.n10701 0.000773889
R20178 VSS.n10840 VSS.n10839 0.000769022
R20179 VSS.n11248 VSS.n11223 0.000752219
R20180 VSS.n10893 VSS.n10872 0.000752101
R20181 VSS.n11027 VSS.n11026 0.000752101
R20182 VSS.n11086 VSS.n11085 0.000752101
R20183 VSS.n11295 VSS.n11294 0.000742997
R20184 VSS.n134 VSS.n133 0.000742997
R20185 VSS.n9823 VSS.n9822 0.000710182
R20186 VSS.n10532 VSS.n10531 0.000702551
R20187 VSS.n10349 VSS.n10348 0.000702551
R20188 VSS.n1458 VSS.n1454 0.00069617
R20189 VSS.n9774 VSS.n794 0.00069617
R20190 VSS.n9822 VSS.n9821 0.00069617
R20191 VSS.n11308 VSS.n127 0.000688976
R20192 VSS.n10115 VSS.n10114 0.000680072
R20193 VSS.n10087 VSS.n487 0.000680072
R20194 VSS.n10064 VSS.n10063 0.000680072
R20195 VSS.n10034 VSS.n235 0.000680072
R20196 VSS.n11129 VSS.n11023 0.000680072
R20197 VSS.n1456 VSS.n1426 0.000640121
R20198 VSS.n9768 VSS.n795 0.000640121
R20199 VSS.n9819 VSS.n9816 0.000640121
R20200 VSS.n750 VSS.n749 0.000640121
R20201 VSS.n11277 VSS.n11276 0.000640121
R20202 VSS.n11081 VSS.n11079 0.00062605
R20203 VSS.n10830 VSS.n10810 0.000622283
R20204 VSS.n10770 VSS.n246 0.000604895
R20205 VSS.n9693 VSS.n9671 0.000604895
R20206 VSS.n9673 VSS.n9672 0.000604895
R20207 VSS.n9692 VSS.n9691 0.000604895
R20208 VSS.n9690 VSS.n9674 0.000604895
R20209 VSS.n9676 VSS.n9675 0.000604895
R20210 VSS.n9689 VSS.n9688 0.000604895
R20211 VSS.n9687 VSS.n9677 0.000604895
R20212 VSS.n9679 VSS.n9678 0.000604895
R20213 VSS.n9686 VSS.n9685 0.000604895
R20214 VSS.n9684 VSS.n9680 0.000604895
R20215 VSS.n9682 VSS.n9681 0.000604895
R20216 VSS.n9683 VSS.n653 0.000604895
R20217 VSS.n1177 VSS.n654 0.000604895
R20218 VSS.n1175 VSS.n1174 0.000604895
R20219 VSS.n1179 VSS.n1178 0.000604895
R20220 VSS.n9853 VSS.n680 0.000604895
R20221 VSS.n682 VSS.n681 0.000604895
R20222 VSS.n9852 VSS.n9851 0.000604895
R20223 VSS.n9850 VSS.n683 0.000604895
R20224 VSS.n685 VSS.n684 0.000604895
R20225 VSS.n9849 VSS.n9848 0.000604895
R20226 VSS.n9847 VSS.n686 0.000604895
R20227 VSS.n688 VSS.n687 0.000604895
R20228 VSS.n9846 VSS.n9845 0.000604895
R20229 VSS.n9844 VSS.n689 0.000604895
R20230 VSS.n691 VSS.n690 0.000604895
R20231 VSS.n9843 VSS.n9842 0.000604895
R20232 VSS.n604 VSS.n546 0.000604895
R20233 VSS.n603 VSS.n602 0.000604895
R20234 VSS.n605 VSS.n601 0.000604895
R20235 VSS.n609 VSS.n606 0.000604895
R20236 VSS.n608 VSS.n607 0.000604895
R20237 VSS.n610 VSS.n600 0.000604895
R20238 VSS.n614 VSS.n611 0.000604895
R20239 VSS.n613 VSS.n612 0.000604895
R20240 VSS.n615 VSS.n599 0.000604895
R20241 VSS.n619 VSS.n616 0.000604895
R20242 VSS.n618 VSS.n617 0.000604895
R20243 VSS.n620 VSS.n598 0.000604895
R20244 VSS.n9906 VSS.n622 0.000604895
R20245 VSS.n625 VSS.n624 0.000604895
R20246 VSS.n9905 VSS.n9904 0.000604895
R20247 VSS.n9701 VSS.n9698 0.000604895
R20248 VSS.n9700 VSS.n9699 0.000604895
R20249 VSS.n9702 VSS.n9697 0.000604895
R20250 VSS.n9706 VSS.n9703 0.000604895
R20251 VSS.n9705 VSS.n9704 0.000604895
R20252 VSS.n9707 VSS.n9696 0.000604895
R20253 VSS.n9711 VSS.n9708 0.000604895
R20254 VSS.n9710 VSS.n9709 0.000604895
R20255 VSS.n9712 VSS.n9695 0.000604895
R20256 VSS.n9716 VSS.n9713 0.000604895
R20257 VSS.n9715 VSS.n9714 0.000604895
R20258 VSS.n9717 VSS.n9694 0.000604895
R20259 VSS.n10573 VSS.n10572 0.000604651
R20260 VSS.n9034 VSS.n9018 0.000603567
R20261 VSS.n9032 VSS.n1560 0.000603567
R20262 VSS.n10147 VSS.n403 0.000603567
R20263 VSS.n10145 VSS.n10144 0.000603567
R20264 VSS.n10207 VSS.n331 0.000603567
R20265 VSS.n10205 VSS.n10204 0.000603567
R20266 VSS.n10267 VSS.n259 0.000603567
R20267 VSS.n10265 VSS.n10264 0.000603567
R20268 VSS.n9339 VSS.n9322 0.000603567
R20269 VSS.n9337 VSS.n9336 0.000603567
R20270 VSS.n9201 VSS.n9185 0.000603567
R20271 VSS.n9199 VSS.n1522 0.000603567
R20272 VSS.n11226 VSS.n11224 0.000598085
R20273 VSS.n10793 VSS.n10792 0.000597826
R20274 VSS.n11083 VSS.n11082 0.000554022
R20275 VSS.n11102 VSS.n11079 0.000554022
R20276 VSS.n11101 VSS.n11080 0.000554022
R20277 VSS.n11085 VSS.n11084 0.000554022
R20278 VSS.n9882 VSS.n9881 0.000552448
R20279 VSS.n9854 VSS.n679 0.000552448
R20280 VSS.n9907 VSS.n621 0.000552448
R20281 VSS.n9903 VSS.n627 0.000552448
R20282 VSS.n11305 VSS.n11304 0.000547244
R20283 VSS.n11228 VSS.n11227 0.000542036
R20284 VSS.n11246 VSS.n11224 0.000542036
R20285 VSS.n11245 VSS.n11225 0.000542036
R20286 VSS.n11230 VSS.n11229 0.000542036
R20287 VSS.n10528 VSS.n10498 0.000533758
R20288 VSS.n9493 VSS.n9492 0.000525989
R20289 VSS.n479 VSS.n466 0.000518007
R20290 VSS.n483 VSS.n463 0.000518007
R20291 VSS.n11144 VSS.n188 0.000518007
R20292 VSS.n11142 VSS.n11141 0.000518007
R20293 VSS.n9586 VSS.n9568 0.000514012
R20294 VSS.n9584 VSS.n9583 0.000514012
R20295 VSS.n176 VSS.n159 0.000514012
R20296 VSS.n174 VSS.n157 0.000514012
R20297 a_52635_34067.t1 a_52635_34067.t61 9.46371
R20298 a_52635_34067.t17 a_52635_34067.t40 8.7152
R20299 a_52635_34067.t27 a_52635_34067.t44 8.7152
R20300 a_52635_34067.n7 a_52635_34067.t133 9.1601
R20301 a_52635_34067.n9 a_52635_34067.t234 9.1601
R20302 a_52635_34067.n13 a_52635_34067.t176 9.17607
R20303 a_52635_34067.n24 a_52635_34067.t121 9.17607
R20304 a_52635_34067.n109 a_52635_34067.t228 8.10567
R20305 a_52635_34067.n92 a_52635_34067.t159 8.10567
R20306 a_52635_34067.n92 a_52635_34067.t98 8.10567
R20307 a_52635_34067.n92 a_52635_34067.t233 8.10567
R20308 a_52635_34067.n92 a_52635_34067.t163 8.10567
R20309 a_52635_34067.n55 a_52635_34067.t169 8.10567
R20310 a_52635_34067.n55 a_52635_34067.t175 8.10567
R20311 a_52635_34067.n55 a_52635_34067.t114 8.10567
R20312 a_52635_34067.n55 a_52635_34067.t201 8.10567
R20313 a_52635_34067.n60 a_52635_34067.t177 8.10567
R20314 a_52635_34067.n60 a_52635_34067.t160 8.10567
R20315 a_52635_34067.n60 a_52635_34067.t99 8.10567
R20316 a_52635_34067.n60 a_52635_34067.t183 8.10567
R20317 a_52635_34067.n90 a_52635_34067.t209 8.10567
R20318 a_52635_34067.n90 a_52635_34067.t100 8.10567
R20319 a_52635_34067.n90 a_52635_34067.t223 8.10567
R20320 a_52635_34067.n58 a_52635_34067.t222 8.10567
R20321 a_52635_34067.n58 a_52635_34067.t118 8.10567
R20322 a_52635_34067.n58 a_52635_34067.t102 8.10567
R20323 a_52635_34067.n109 a_52635_34067.t198 8.10567
R20324 a_52635_34067.n109 a_52635_34067.t129 8.10567
R20325 a_52635_34067.n109 a_52635_34067.t197 8.10567
R20326 a_52635_34067.n116 a_52635_34067.t224 8.10567
R20327 a_52635_34067.n107 a_52635_34067.t149 8.10567
R20328 a_52635_34067.n107 a_52635_34067.t88 8.10567
R20329 a_52635_34067.n107 a_52635_34067.t232 8.10567
R20330 a_52635_34067.n107 a_52635_34067.t155 8.10567
R20331 a_52635_34067.n74 a_52635_34067.t161 8.10567
R20332 a_52635_34067.n74 a_52635_34067.t165 8.10567
R20333 a_52635_34067.n74 a_52635_34067.t106 8.10567
R20334 a_52635_34067.n74 a_52635_34067.t194 8.10567
R20335 a_52635_34067.n75 a_52635_34067.t168 8.10567
R20336 a_52635_34067.n75 a_52635_34067.t151 8.10567
R20337 a_52635_34067.n75 a_52635_34067.t93 8.10567
R20338 a_52635_34067.n75 a_52635_34067.t174 8.10567
R20339 a_52635_34067.n102 a_52635_34067.t162 8.10567
R20340 a_52635_34067.n102 a_52635_34067.t238 8.10567
R20341 a_52635_34067.n102 a_52635_34067.t189 8.10567
R20342 a_52635_34067.n100 a_52635_34067.t182 8.10567
R20343 a_52635_34067.n100 a_52635_34067.t79 8.10567
R20344 a_52635_34067.n100 a_52635_34067.t65 8.10567
R20345 a_52635_34067.n116 a_52635_34067.t187 8.10567
R20346 a_52635_34067.n116 a_52635_34067.t123 8.10567
R20347 a_52635_34067.n116 a_52635_34067.t185 8.10567
R20348 a_52635_34067.n111 a_52635_34067.t179 8.10567
R20349 a_52635_34067.n95 a_52635_34067.t105 8.10567
R20350 a_52635_34067.n95 a_52635_34067.t225 8.10567
R20351 a_52635_34067.n95 a_52635_34067.t195 8.10567
R20352 a_52635_34067.n95 a_52635_34067.t112 8.10567
R20353 a_52635_34067.n64 a_52635_34067.t116 8.10567
R20354 a_52635_34067.n64 a_52635_34067.t120 8.10567
R20355 a_52635_34067.n64 a_52635_34067.t235 8.10567
R20356 a_52635_34067.n64 a_52635_34067.t140 8.10567
R20357 a_52635_34067.n68 a_52635_34067.t122 8.10567
R20358 a_52635_34067.n68 a_52635_34067.t109 8.10567
R20359 a_52635_34067.n68 a_52635_34067.t226 8.10567
R20360 a_52635_34067.n68 a_52635_34067.t127 8.10567
R20361 a_52635_34067.n88 a_52635_34067.t146 8.10567
R20362 a_52635_34067.n88 a_52635_34067.t229 8.10567
R20363 a_52635_34067.n88 a_52635_34067.t171 8.10567
R20364 a_52635_34067.n86 a_52635_34067.t164 8.10567
R20365 a_52635_34067.n86 a_52635_34067.t66 8.10567
R20366 a_52635_34067.n86 a_52635_34067.t231 8.10567
R20367 a_52635_34067.n111 a_52635_34067.t137 8.10567
R20368 a_52635_34067.n111 a_52635_34067.t77 8.10567
R20369 a_52635_34067.n111 a_52635_34067.t136 8.10567
R20370 a_52635_34067.n112 a_52635_34067.t145 8.10567
R20371 a_52635_34067.n104 a_52635_34067.t72 8.10567
R20372 a_52635_34067.n104 a_52635_34067.t205 8.10567
R20373 a_52635_34067.n104 a_52635_34067.t158 8.10567
R20374 a_52635_34067.n104 a_52635_34067.t81 8.10567
R20375 a_52635_34067.n82 a_52635_34067.t83 8.10567
R20376 a_52635_34067.n82 a_52635_34067.t89 8.10567
R20377 a_52635_34067.n82 a_52635_34067.t217 8.10567
R20378 a_52635_34067.n82 a_52635_34067.t113 8.10567
R20379 a_52635_34067.n79 a_52635_34067.t92 8.10567
R20380 a_52635_34067.n79 a_52635_34067.t76 8.10567
R20381 a_52635_34067.n79 a_52635_34067.t206 8.10567
R20382 a_52635_34067.n79 a_52635_34067.t97 8.10567
R20383 a_52635_34067.n98 a_52635_34067.t86 8.10567
R20384 a_52635_34067.n98 a_52635_34067.t170 8.10567
R20385 a_52635_34067.n98 a_52635_34067.t111 8.10567
R20386 a_52635_34067.n96 a_52635_34067.t104 8.10567
R20387 a_52635_34067.n96 a_52635_34067.t191 8.10567
R20388 a_52635_34067.n96 a_52635_34067.t172 8.10567
R20389 a_52635_34067.n112 a_52635_34067.t110 8.10567
R20390 a_52635_34067.n112 a_52635_34067.t227 8.10567
R20391 a_52635_34067.n112 a_52635_34067.t108 8.10567
R20392 a_52635_34067.n19 a_52635_34067.t188 8.10567
R20393 a_52635_34067.n19 a_52635_34067.t196 8.10567
R20394 a_52635_34067.n19 a_52635_34067.t128 8.10567
R20395 a_52635_34067.n19 a_52635_34067.t216 8.10567
R20396 a_52635_34067.n11 a_52635_34067.t193 8.10567
R20397 a_52635_34067.n177 a_52635_34067.t84 8.10567
R20398 a_52635_34067.n176 a_52635_34067.t214 8.10567
R20399 a_52635_34067.n12 a_52635_34067.t115 8.10567
R20400 a_52635_34067.n12 a_52635_34067.t69 8.10567
R20401 a_52635_34067.n12 a_52635_34067.t181 8.10567
R20402 a_52635_34067.n1 a_52635_34067.t240 8.10567
R20403 a_52635_34067.n1 a_52635_34067.t213 8.10567
R20404 a_52635_34067.n1 a_52635_34067.t144 8.10567
R20405 a_52635_34067.n41 a_52635_34067.t210 8.10567
R20406 a_52635_34067.n175 a_52635_34067.t101 8.10567
R20407 a_52635_34067.n174 a_52635_34067.t85 8.10567
R20408 a_52635_34067.n16 a_52635_34067.t199 8.10567
R20409 a_52635_34067.n16 a_52635_34067.t178 8.10567
R20410 a_52635_34067.n42 a_52635_34067.t117 8.10567
R20411 a_52635_34067.n42 a_52635_34067.t203 8.10567
R20412 a_52635_34067.n36 a_52635_34067.t143 8.10567
R20413 a_52635_34067.n36 a_52635_34067.t148 8.10567
R20414 a_52635_34067.n36 a_52635_34067.t87 8.10567
R20415 a_52635_34067.n36 a_52635_34067.t173 8.10567
R20416 a_52635_34067.n5 a_52635_34067.t180 8.10567
R20417 a_52635_34067.n155 a_52635_34067.t78 8.10567
R20418 a_52635_34067.n154 a_52635_34067.t207 8.10567
R20419 a_52635_34067.n6 a_52635_34067.t70 8.10567
R20420 a_52635_34067.n6 a_52635_34067.t221 8.10567
R20421 a_52635_34067.n6 a_52635_34067.t139 8.10567
R20422 a_52635_34067.n27 a_52635_34067.t215 8.10567
R20423 a_52635_34067.n27 a_52635_34067.t167 8.10567
R20424 a_52635_34067.n27 a_52635_34067.t107 8.10567
R20425 a_52635_34067.n51 a_52635_34067.t202 8.10567
R20426 a_52635_34067.n153 a_52635_34067.t95 8.10567
R20427 a_52635_34067.n152 a_52635_34067.t80 8.10567
R20428 a_52635_34067.n43 a_52635_34067.t150 8.10567
R20429 a_52635_34067.n43 a_52635_34067.t134 8.10567
R20430 a_52635_34067.n47 a_52635_34067.t74 8.10567
R20431 a_52635_34067.n47 a_52635_34067.t156 8.10567
R20432 a_52635_34067.n21 a_52635_34067.t130 8.10567
R20433 a_52635_34067.n21 a_52635_34067.t135 8.10567
R20434 a_52635_34067.n21 a_52635_34067.t75 8.10567
R20435 a_52635_34067.n21 a_52635_34067.t157 8.10567
R20436 a_52635_34067.n157 a_52635_34067.t132 8.10567
R20437 a_52635_34067.n158 a_52635_34067.t219 8.10567
R20438 a_52635_34067.n20 a_52635_34067.t154 8.10567
R20439 a_52635_34067.n25 a_52635_34067.t236 8.10567
R20440 a_52635_34067.n25 a_52635_34067.t211 8.10567
R20441 a_52635_34067.n25 a_52635_34067.t126 8.10567
R20442 a_52635_34067.n4 a_52635_34067.t200 8.10567
R20443 a_52635_34067.n4 a_52635_34067.t153 8.10567
R20444 a_52635_34067.n4 a_52635_34067.t94 8.10567
R20445 a_52635_34067.n37 a_52635_34067.t147 8.10567
R20446 a_52635_34067.n151 a_52635_34067.t230 8.10567
R20447 a_52635_34067.n150 a_52635_34067.t220 8.10567
R20448 a_52635_34067.n38 a_52635_34067.t138 8.10567
R20449 a_52635_34067.n38 a_52635_34067.t124 8.10567
R20450 a_52635_34067.n39 a_52635_34067.t239 8.10567
R20451 a_52635_34067.n39 a_52635_34067.t142 8.10567
R20452 a_52635_34067.n33 a_52635_34067.t68 8.10567
R20453 a_52635_34067.n33 a_52635_34067.t71 8.10567
R20454 a_52635_34067.n33 a_52635_34067.t204 8.10567
R20455 a_52635_34067.n33 a_52635_34067.t96 8.10567
R20456 a_52635_34067.n162 a_52635_34067.t103 8.10567
R20457 a_52635_34067.n163 a_52635_34067.t190 8.10567
R20458 a_52635_34067.n31 a_52635_34067.t125 8.10567
R20459 a_52635_34067.n10 a_52635_34067.t184 8.10567
R20460 a_52635_34067.n10 a_52635_34067.t141 8.10567
R20461 a_52635_34067.n10 a_52635_34067.t67 8.10567
R20462 a_52635_34067.n30 a_52635_34067.t131 8.10567
R20463 a_52635_34067.n30 a_52635_34067.t91 8.10567
R20464 a_52635_34067.n30 a_52635_34067.t218 8.10567
R20465 a_52635_34067.n48 a_52635_34067.t119 8.10567
R20466 a_52635_34067.n161 a_52635_34067.t208 8.10567
R20467 a_52635_34067.n160 a_52635_34067.t192 8.10567
R20468 a_52635_34067.n45 a_52635_34067.t73 8.10567
R20469 a_52635_34067.n45 a_52635_34067.t237 8.10567
R20470 a_52635_34067.n49 a_52635_34067.t186 8.10567
R20471 a_52635_34067.n49 a_52635_34067.t82 8.10567
R20472 a_52635_34067.t17 a_52635_34067.n212 7.22198
R20473 a_52635_34067.t27 a_52635_34067.n195 7.22198
R20474 a_52635_34067.t4 a_52635_34067.t0 7.12006
R20475 a_52635_34067.n182 a_52635_34067.t10 6.77653
R20476 a_52635_34067.n142 a_52635_34067.t60 6.77653
R20477 a_52635_34067.n141 a_52635_34067.t49 6.7761
R20478 a_52635_34067.n205 a_52635_34067.t50 6.7761
R20479 a_52635_34067.n138 a_52635_34067.t2 6.86989
R20480 a_52635_34067.n127 a_52635_34067.t19 6.77231
R20481 a_52635_34067.n137 a_52635_34067.t28 6.77231
R20482 a_52635_34067.n188 a_52635_34067.t3 6.14835
R20483 a_52635_34067.n186 a_52635_34067.t62 6.14517
R20484 a_52635_34067.n140 a_52635_34067.t45 5.85898
R20485 a_52635_34067.t21 a_52635_34067.t18 5.70489
R20486 a_52635_34067.n195 a_52635_34067.t30 5.70489
R20487 a_52635_34067.t13 a_52635_34067.t39 5.70489
R20488 a_52635_34067.n212 a_52635_34067.t22 5.70489
R20489 a_52635_34067.n185 a_52635_34067.t64 5.61877
R20490 a_52635_34067.n143 a_52635_34067.t31 5.50607
R20491 a_52635_34067.n203 a_52635_34067.t53 5.50607
R20492 a_52635_34067.n183 a_52635_34067.t33 5.50607
R20493 a_52635_34067.n142 a_52635_34067.t48 5.50475
R20494 a_52635_34067.n141 a_52635_34067.t34 5.50475
R20495 a_52635_34067.n182 a_52635_34067.t11 5.50475
R20496 a_52635_34067.n199 a_52635_34067.t43 5.50475
R20497 a_52635_34067.n202 a_52635_34067.t47 5.50475
R20498 a_52635_34067.n205 a_52635_34067.t35 5.50475
R20499 a_52635_34067.n216 a_52635_34067.t42 5.50475
R20500 a_52635_34067.n139 a_52635_34067.t52 5.50475
R20501 a_52635_34067.n144 a_52635_34067.t55 5.50475
R20502 a_52635_34067.n204 a_52635_34067.t51 5.50475
R20503 a_52635_34067.n201 a_52635_34067.t15 5.50475
R20504 a_52635_34067.n200 a_52635_34067.t56 5.50475
R20505 a_52635_34067.n184 a_52635_34067.t59 5.50475
R20506 a_52635_34067.t5 a_52635_34067.n140 5.50475
R20507 a_52635_34067.n17 a_52635_34067.n16 0.595624
R20508 a_52635_34067.n85 a_52635_34067.n38 0.595624
R20509 a_52635_34067.n34 a_52635_34067.n43 0.607617
R20510 a_52635_34067.n46 a_52635_34067.n45 0.607617
R20511 a_52635_34067.n118 a_52635_34067.t37 5.5012
R20512 a_52635_34067.t57 a_52635_34067.n119 5.5012
R20513 a_52635_34067.t58 a_52635_34067.n120 5.5012
R20514 a_52635_34067.t6 a_52635_34067.n121 5.5012
R20515 a_52635_34067.t25 a_52635_34067.n122 5.5012
R20516 a_52635_34067.t7 a_52635_34067.n123 5.5012
R20517 a_52635_34067.t46 a_52635_34067.n124 5.5012
R20518 a_52635_34067.t12 a_52635_34067.n125 5.5012
R20519 a_52635_34067.t36 a_52635_34067.n126 5.5012
R20520 a_52635_34067.t20 a_52635_34067.n127 5.5012
R20521 a_52635_34067.n128 a_52635_34067.t41 5.5012
R20522 a_52635_34067.n129 a_52635_34067.t14 5.5012
R20523 a_52635_34067.n130 a_52635_34067.t16 5.5012
R20524 a_52635_34067.n131 a_52635_34067.t23 5.5012
R20525 a_52635_34067.n132 a_52635_34067.t32 5.5012
R20526 a_52635_34067.n133 a_52635_34067.t24 5.5012
R20527 a_52635_34067.n134 a_52635_34067.t9 5.5012
R20528 a_52635_34067.t26 a_52635_34067.n135 5.5012
R20529 a_52635_34067.t38 a_52635_34067.n136 5.5012
R20530 a_52635_34067.t29 a_52635_34067.n137 5.5012
R20531 a_52635_34067.t63 a_52635_34067.n138 5.66099
R20532 a_52635_34067.n107 a_52635_34067.n106 0.020246
R20533 a_52635_34067.n105 a_52635_34067.n104 0.020246
R20534 a_52635_34067.n74 a_52635_34067.n72 0.150783
R20535 a_52635_34067.n75 a_52635_34067.n71 0.150803
R20536 a_52635_34067.n116 a_52635_34067.n115 0.0676355
R20537 a_52635_34067.n82 a_52635_34067.n81 0.150803
R20538 a_52635_34067.n80 a_52635_34067.n79 0.150806
R20539 a_52635_34067.n113 a_52635_34067.n112 0.0676255
R20540 a_52635_34067.n60 a_52635_34067.n53 0.153625
R20541 a_52635_34067.n55 a_52635_34067.n54 0.153625
R20542 a_52635_34067.n93 a_52635_34067.n92 0.020088
R20543 a_52635_34067.n76 a_52635_34067.n75 0.246907
R20544 a_52635_34067.n74 a_52635_34067.n73 0.246877
R20545 a_52635_34067.n69 a_52635_34067.n68 0.153625
R20546 a_52635_34067.n65 a_52635_34067.n64 0.153625
R20547 a_52635_34067.n95 a_52635_34067.n94 0.020088
R20548 a_52635_34067.n111 a_52635_34067.n110 0.0201939
R20549 a_52635_34067.n68 a_52635_34067.n67 0.246907
R20550 a_52635_34067.n64 a_52635_34067.n63 0.246907
R20551 a_52635_34067.n79 a_52635_34067.n84 0.246907
R20552 a_52635_34067.n83 a_52635_34067.n82 0.246907
R20553 a_52635_34067.n109 a_52635_34067.n57 0.0201939
R20554 a_52635_34067.n61 a_52635_34067.n60 0.246907
R20555 a_52635_34067.n56 a_52635_34067.n55 0.246907
R20556 a_52635_34067.n27 a_52635_34067.n26 0.260442
R20557 a_52635_34067.n52 a_52635_34067.n47 0.591264
R20558 a_52635_34067.n36 a_52635_34067.n35 0.310971
R20559 a_52635_34067.n7 a_52635_34067.n6 0.258567
R20560 a_52635_34067.n4 a_52635_34067.n3 0.208479
R20561 a_52635_34067.n40 a_52635_34067.n39 0.591642
R20562 a_52635_34067.n22 a_52635_34067.n21 0.623337
R20563 a_52635_34067.n25 a_52635_34067.n24 0.259585
R20564 a_52635_34067.n30 a_52635_34067.n29 0.260442
R20565 a_52635_34067.n50 a_52635_34067.n49 0.591264
R20566 a_52635_34067.n33 a_52635_34067.n32 0.310971
R20567 a_52635_34067.n10 a_52635_34067.n9 0.258567
R20568 a_52635_34067.n1 a_52635_34067.n0 0.208479
R20569 a_52635_34067.n42 a_52635_34067.n15 0.591642
R20570 a_52635_34067.n19 a_52635_34067.n18 0.623337
R20571 a_52635_34067.n13 a_52635_34067.n12 0.259585
R20572 a_52635_34067.n191 a_52635_34067.n190 3.48654
R20573 a_52635_34067.n194 a_52635_34067.n190 3.42822
R20574 a_52635_34067.n147 a_52635_34067.n145 3.37173
R20575 a_52635_34067.t13 a_52635_34067.n211 3.23904
R20576 a_52635_34067.t21 a_52635_34067.n181 3.23904
R20577 a_52635_34067.n187 a_52635_34067.t4 3.23004
R20578 a_52635_34067.n201 a_52635_34067.n200 2.60203
R20579 a_52635_34067.n140 a_52635_34067.n139 2.60203
R20580 a_52635_34067.n184 a_52635_34067.n183 2.52436
R20581 a_52635_34067.n204 a_52635_34067.n203 2.52436
R20582 a_52635_34067.n144 a_52635_34067.n143 2.52436
R20583 a_52635_34067.n171 a_52635_34067.n170 2.40699
R20584 a_52635_34067.n159 a_52635_34067.n149 2.30989
R20585 a_52635_34067.n156 a_52635_34067.n44 2.30989
R20586 a_52635_34067.n187 a_52635_34067.n186 2.2807
R20587 a_52635_34067.n91 a_52635_34067.n90 0.427602
R20588 a_52635_34067.n59 a_52635_34067.n58 0.427602
R20589 a_52635_34067.n89 a_52635_34067.n88 0.427602
R20590 a_52635_34067.n87 a_52635_34067.n86 0.427602
R20591 a_52635_34067.n103 a_52635_34067.n102 0.420727
R20592 a_52635_34067.n101 a_52635_34067.n100 0.420727
R20593 a_52635_34067.n99 a_52635_34067.n98 0.420727
R20594 a_52635_34067.n97 a_52635_34067.n96 0.420727
R20595 a_52635_34067.n67 a_52635_34067.n66 2.96488
R20596 a_52635_34067.n62 a_52635_34067.n94 2.94096
R20597 a_52635_34067.n108 a_52635_34067.n61 2.96488
R20598 a_52635_34067.n93 a_52635_34067.n117 2.94096
R20599 a_52635_34067.n166 a_52635_34067.n114 2.07182
R20600 a_52635_34067.n167 a_52635_34067.n70 2.07182
R20601 a_52635_34067.n114 a_52635_34067.n71 2.75706
R20602 a_52635_34067.n106 a_52635_34067.n70 2.90773
R20603 a_52635_34067.n80 a_52635_34067.n78 2.75704
R20604 a_52635_34067.n77 a_52635_34067.n105 2.90773
R20605 a_52635_34067.n169 a_52635_34067.n147 1.80314
R20606 a_52635_34067.n180 a_52635_34067.n179 1.70908
R20607 a_52635_34067.n172 a_52635_34067.n171 1.68395
R20608 a_52635_34067.n179 a_52635_34067.n178 1.68395
R20609 a_52635_34067.n78 a_52635_34067.n165 1.5005
R20610 a_52635_34067.n66 a_52635_34067.n166 1.5005
R20611 a_52635_34067.n170 a_52635_34067.n108 1.5005
R20612 a_52635_34067.n117 a_52635_34067.n169 1.5005
R20613 a_52635_34067.n168 a_52635_34067.n77 1.5005
R20614 a_52635_34067.n167 a_52635_34067.n62 1.5005
R20615 a_52635_34067.n164 a_52635_34067.n28 1.5005
R20616 a_52635_34067.n159 a_52635_34067.n2 1.5005
R20617 a_52635_34067.n173 a_52635_34067.n172 1.5005
R20618 a_52635_34067.n178 a_52635_34067.n14 1.5005
R20619 a_52635_34067.n8 a_52635_34067.n148 1.5005
R20620 a_52635_34067.n23 a_52635_34067.n156 1.5005
R20621 a_52635_34067.n194 a_52635_34067.n193 1.5005
R20622 a_52635_34067.n196 a_52635_34067.t27 1.5005
R20623 a_52635_34067.n198 a_52635_34067.n197 1.5005
R20624 a_52635_34067.n208 a_52635_34067.n146 1.5005
R20625 a_52635_34067.n213 a_52635_34067.t17 1.5005
R20626 a_52635_34067.n189 a_52635_34067.n188 1.5005
R20627 a_52635_34067.n192 a_52635_34067.n191 1.5005
R20628 a_52635_34067.n207 a_52635_34067.n206 1.5005
R20629 a_52635_34067.n210 a_52635_34067.n209 1.5005
R20630 a_52635_34067.n180 a_52635_34067.t45 1.5005
R20631 a_52635_34067.n215 a_52635_34067.n214 1.5005
R20632 a_52635_34067.n166 a_52635_34067.n165 1.47516
R20633 a_52635_34067.n168 a_52635_34067.n167 1.47516
R20634 a_52635_34067.n190 a_52635_34067.n189 1.41182
R20635 a_52635_34067.n26 a_52635_34067.t166 9.17619
R20636 a_52635_34067.n29 a_52635_34067.t90 9.17619
R20637 a_52635_34067.n212 a_52635_34067.t13 1.27228
R20638 a_52635_34067.n200 a_52635_34067.n199 1.27228
R20639 a_52635_34067.n202 a_52635_34067.n201 1.27228
R20640 a_52635_34067.n195 a_52635_34067.t21 1.27228
R20641 a_52635_34067.n139 a_52635_34067.n216 1.27228
R20642 a_52635_34067.n183 a_52635_34067.n182 1.26756
R20643 a_52635_34067.n203 a_52635_34067.n202 1.26756
R20644 a_52635_34067.n143 a_52635_34067.n142 1.26756
R20645 a_52635_34067.n6 a_52635_34067.n5 1.24866
R20646 a_52635_34067.n47 a_52635_34067.n51 1.24866
R20647 a_52635_34067.n162 a_52635_34067.n10 1.24866
R20648 a_52635_34067.n49 a_52635_34067.n48 1.24866
R20649 a_52635_34067.n152 a_52635_34067.n27 1.24629
R20650 a_52635_34067.n160 a_52635_34067.n30 1.24629
R20651 a_52635_34067.n164 a_52635_34067.n159 1.23709
R20652 a_52635_34067.n156 a_52635_34067.n148 1.23709
R20653 a_52635_34067.n176 a_52635_34067.n19 1.22261
R20654 a_52635_34067.n174 a_52635_34067.n1 1.22261
R20655 a_52635_34067.n21 a_52635_34067.n20 1.22261
R20656 a_52635_34067.n150 a_52635_34067.n4 1.22261
R20657 a_52635_34067.n12 a_52635_34067.n11 1.21313
R20658 a_52635_34067.n42 a_52635_34067.n41 1.21313
R20659 a_52635_34067.n157 a_52635_34067.n25 1.21313
R20660 a_52635_34067.n39 a_52635_34067.n37 1.21313
R20661 a_52635_34067.n214 a_52635_34067.n145 1.10472
R20662 a_52635_34067.n172 a_52635_34067.n164 0.809892
R20663 a_52635_34067.n178 a_52635_34067.n148 0.809892
R20664 a_52635_34067.n198 a_52635_34067.n184 0.796291
R20665 a_52635_34067.n206 a_52635_34067.n204 0.796291
R20666 a_52635_34067.n215 a_52635_34067.n144 0.796291
R20667 a_52635_34067.n213 a_52635_34067.n146 0.780703
R20668 a_52635_34067.n196 a_52635_34067.n194 0.780703
R20669 a_52635_34067.n211 a_52635_34067.n210 0.780703
R20670 a_52635_34067.n191 a_52635_34067.n181 0.780703
R20671 a_52635_34067.n188 a_52635_34067.t1 0.769291
R20672 a_52635_34067.n186 a_52635_34067.n185 0.767125
R20673 a_52635_34067.n52 a_52635_34067.n149 1.14908
R20674 a_52635_34067.n44 a_52635_34067.n7 1.39299
R20675 a_52635_34067.n28 a_52635_34067.n50 1.14908
R20676 a_52635_34067.n9 a_52635_34067.n8 1.39299
R20677 a_52635_34067.n2 a_52635_34067.n40 1.11421
R20678 a_52635_34067.n24 a_52635_34067.n23 1.35707
R20679 a_52635_34067.n173 a_52635_34067.n15 1.11421
R20680 a_52635_34067.n14 a_52635_34067.n13 1.35707
R20681 a_52635_34067.n177 a_52635_34067.n176 0.673132
R20682 a_52635_34067.n11 a_52635_34067.n177 0.673132
R20683 a_52635_34067.n175 a_52635_34067.n174 0.673132
R20684 a_52635_34067.n41 a_52635_34067.n175 0.673132
R20685 a_52635_34067.n155 a_52635_34067.n154 0.673132
R20686 a_52635_34067.n5 a_52635_34067.n155 0.673132
R20687 a_52635_34067.n153 a_52635_34067.n152 0.673132
R20688 a_52635_34067.n51 a_52635_34067.n153 0.673132
R20689 a_52635_34067.n20 a_52635_34067.n158 0.673132
R20690 a_52635_34067.n158 a_52635_34067.n157 0.673132
R20691 a_52635_34067.n151 a_52635_34067.n150 0.673132
R20692 a_52635_34067.n37 a_52635_34067.n151 0.673132
R20693 a_52635_34067.n31 a_52635_34067.n163 0.673132
R20694 a_52635_34067.n163 a_52635_34067.n162 0.673132
R20695 a_52635_34067.n161 a_52635_34067.n160 0.673132
R20696 a_52635_34067.n48 a_52635_34067.n161 0.673132
R20697 a_52635_34067.n214 a_52635_34067.n213 0.638405
R20698 a_52635_34067.n197 a_52635_34067.n196 0.638405
R20699 a_52635_34067.n189 a_52635_34067.n187 0.638405
R20700 a_52635_34067.n211 a_52635_34067.n180 0.638405
R20701 a_52635_34067.n207 a_52635_34067.n181 0.638405
R20702 a_52635_34067.n197 a_52635_34067.n146 0.628372
R20703 a_52635_34067.n210 a_52635_34067.n207 0.628372
R20704 a_52635_34067.n179 a_52635_34067.n147 0.604355
R20705 a_52635_34067.n171 a_52635_34067.n145 0.603852
R20706 a_52635_34067.n170 a_52635_34067.n165 0.571818
R20707 a_52635_34067.n169 a_52635_34067.n168 0.571818
R20708 a_52635_34067.n199 a_52635_34067.n198 0.476484
R20709 a_52635_34067.n206 a_52635_34067.n205 0.476484
R20710 a_52635_34067.n216 a_52635_34067.n215 0.476484
R20711 a_52635_34067.t45 a_52635_34067.n141 0.476484
R20712 a_52635_34067.n52 a_52635_34067.n34 1.14166
R20713 a_52635_34067.n44 a_52635_34067.n35 2.75347
R20714 a_52635_34067.n46 a_52635_34067.n50 1.14166
R20715 a_52635_34067.n8 a_52635_34067.n32 2.75347
R20716 a_52635_34067.n124 a_52635_34067.n208 0.478684
R20717 a_52635_34067.n209 a_52635_34067.n118 0.478684
R20718 a_52635_34067.n193 a_52635_34067.n134 0.478684
R20719 a_52635_34067.n192 a_52635_34067.n128 0.478684
R20720 a_52635_34067.n59 a_52635_34067.n57 2.03311
R20721 a_52635_34067.n53 a_52635_34067.n59 2.04491
R20722 a_52635_34067.n54 a_52635_34067.n53 4.37762
R20723 a_52635_34067.n91 a_52635_34067.n54 1.87961
R20724 a_52635_34067.n91 a_52635_34067.n93 2.19836
R20725 a_52635_34067.n101 a_52635_34067.n115 2.03667
R20726 a_52635_34067.n76 a_52635_34067.n101 2.2172
R20727 a_52635_34067.n76 a_52635_34067.n73 4.49278
R20728 a_52635_34067.n103 a_52635_34067.n73 1.82125
R20729 a_52635_34067.n103 a_52635_34067.n106 2.19319
R20730 a_52635_34067.n115 a_52635_34067.n114 1.65342
R20731 a_52635_34067.n72 a_52635_34067.n71 4.34534
R20732 a_52635_34067.n72 a_52635_34067.n70 1.50598
R20733 a_52635_34067.n87 a_52635_34067.n110 2.03311
R20734 a_52635_34067.n69 a_52635_34067.n87 2.04491
R20735 a_52635_34067.n65 a_52635_34067.n69 4.37762
R20736 a_52635_34067.n89 a_52635_34067.n65 1.87961
R20737 a_52635_34067.n94 a_52635_34067.n89 2.19836
R20738 a_52635_34067.n66 a_52635_34067.n110 1.65903
R20739 a_52635_34067.n67 a_52635_34067.n63 4.49309
R20740 a_52635_34067.n63 a_52635_34067.n62 1.44546
R20741 a_52635_34067.n97 a_52635_34067.n113 2.03657
R20742 a_52635_34067.n97 a_52635_34067.n84 2.21715
R20743 a_52635_34067.n83 a_52635_34067.n84 4.49317
R20744 a_52635_34067.n99 a_52635_34067.n83 1.82113
R20745 a_52635_34067.n105 a_52635_34067.n99 2.19319
R20746 a_52635_34067.n78 a_52635_34067.n113 1.65366
R20747 a_52635_34067.n81 a_52635_34067.n80 4.34574
R20748 a_52635_34067.n81 a_52635_34067.n77 1.50586
R20749 a_52635_34067.n57 a_52635_34067.n108 1.65903
R20750 a_52635_34067.n61 a_52635_34067.n56 4.49309
R20751 a_52635_34067.n56 a_52635_34067.n117 1.44546
R20752 a_52635_34067.n149 a_52635_34067.n26 2.8103
R20753 a_52635_34067.n35 a_52635_34067.n34 4.38327
R20754 a_52635_34067.n3 a_52635_34067.n2 2.83621
R20755 a_52635_34067.n40 a_52635_34067.n85 1.15119
R20756 a_52635_34067.n85 a_52635_34067.n22 4.37089
R20757 a_52635_34067.n22 a_52635_34067.n23 2.6764
R20758 a_52635_34067.n29 a_52635_34067.n28 2.8103
R20759 a_52635_34067.n46 a_52635_34067.n32 4.38327
R20760 a_52635_34067.n173 a_52635_34067.n0 2.83621
R20761 a_52635_34067.n17 a_52635_34067.n15 1.15119
R20762 a_52635_34067.n18 a_52635_34067.n17 4.37089
R20763 a_52635_34067.n18 a_52635_34067.n14 2.6764
R20764 a_52635_34067.n126 a_52635_34067.n127 1.27228
R20765 a_52635_34067.n125 a_52635_34067.n126 2.51878
R20766 a_52635_34067.n208 a_52635_34067.n125 0.794091
R20767 a_52635_34067.n123 a_52635_34067.n124 1.27228
R20768 a_52635_34067.n122 a_52635_34067.n123 2.60203
R20769 a_52635_34067.n121 a_52635_34067.n122 1.27228
R20770 a_52635_34067.n120 a_52635_34067.n121 1.27228
R20771 a_52635_34067.n119 a_52635_34067.n120 2.51878
R20772 a_52635_34067.n209 a_52635_34067.n119 0.794091
R20773 a_52635_34067.t54 a_52635_34067.n118 6.77266
R20774 a_52635_34067.n136 a_52635_34067.n137 1.27228
R20775 a_52635_34067.n135 a_52635_34067.n136 2.51878
R20776 a_52635_34067.n193 a_52635_34067.n135 0.794091
R20777 a_52635_34067.n133 a_52635_34067.n134 1.27228
R20778 a_52635_34067.n132 a_52635_34067.n133 2.60203
R20779 a_52635_34067.n131 a_52635_34067.n132 1.27228
R20780 a_52635_34067.n130 a_52635_34067.n131 1.27228
R20781 a_52635_34067.n129 a_52635_34067.n130 2.51878
R20782 a_52635_34067.n192 a_52635_34067.n129 0.794091
R20783 a_52635_34067.t8 a_52635_34067.n128 6.77266
R20784 a_52635_34067.n185 a_52635_34067.n138 3.17898
R20785 a_52635_34067.n16 a_52635_34067.n42 2.16997
R20786 a_52635_34067.n39 a_52635_34067.n38 2.16997
R20787 a_52635_34067.n154 a_52635_34067.n36 2.13563
R20788 a_52635_34067.n33 a_52635_34067.n31 2.13563
R20789 a_52635_34067.n43 a_52635_34067.n47 2.13445
R20790 a_52635_34067.n49 a_52635_34067.n45 2.13445
R20791 a_52635_34067.t152 a_52635_34067.n3 9.16748
R20792 a_52635_34067.t212 a_52635_34067.n0 9.16748
R20793 VDD.n7996 VDD.n2188 714.056
R20794 VDD.n7994 VDD.n2188 712.232
R20795 VDD.n7996 VDD.n2187 707.59
R20796 VDD.n7994 VDD.n2187 705.766
R20797 VDD.n1743 VDD.n686 694.492
R20798 VDD.n1717 VDD.n710 694.492
R20799 VDD.n1351 VDD.n1350 694.492
R20800 VDD.n1427 VDD.n850 694.492
R20801 VDD.n1416 VDD.n845 694.492
R20802 VDD.n1720 VDD.n707 694.492
R20803 VDD.n1653 VDD.n758 694.492
R20804 VDD.n1344 VDD.n1343 694.492
R20805 VDD.n1357 VDD.n848 694.492
R20806 VDD.n1413 VDD.n875 694.492
R20807 VDD.n762 VDD.n760 694.492
R20808 VDD.n1741 VDD.n691 694.492
R20809 VDD.n688 VDD.n686 694.078
R20810 VDD.n711 VDD.n710 694.078
R20811 VDD.n1351 VDD.n1276 694.078
R20812 VDD.n1427 VDD.n849 694.078
R20813 VDD.n1416 VDD.n846 694.078
R20814 VDD.n1720 VDD.n708 694.078
R20815 VDD.n761 VDD.n758 694.078
R20816 VDD.n1348 VDD.n1344 694.078
R20817 VDD.n1355 VDD.n848 694.078
R20818 VDD.n1390 VDD.n875 694.078
R20819 VDD.n1651 VDD.n762 694.078
R20820 VDD.n691 VDD.n689 694.078
R20821 VDD.n1743 VDD.n687 692.172
R20822 VDD.n1717 VDD.n712 692.172
R20823 VDD.n1350 VDD.n1277 692.172
R20824 VDD.n1353 VDD.n850 692.172
R20825 VDD.n1430 VDD.n845 692.172
R20826 VDD.n859 VDD.n707 692.172
R20827 VDD.n1653 VDD.n759 692.172
R20828 VDD.n1347 VDD.n1343 692.172
R20829 VDD.n1357 VDD.n1083 692.172
R20830 VDD.n1413 VDD.n847 692.172
R20831 VDD.n764 VDD.n760 692.172
R20832 VDD.n1741 VDD.n692 692.172
R20833 VDD.n688 VDD.n687 691.758
R20834 VDD.n712 VDD.n711 691.758
R20835 VDD.n1277 VDD.n1276 691.758
R20836 VDD.n1353 VDD.n849 691.758
R20837 VDD.n1430 VDD.n846 691.758
R20838 VDD.n859 VDD.n708 691.758
R20839 VDD.n761 VDD.n759 691.758
R20840 VDD.n1348 VDD.n1347 691.758
R20841 VDD.n1355 VDD.n1083 691.758
R20842 VDD.n1390 VDD.n847 691.758
R20843 VDD.n1651 VDD.n764 691.758
R20844 VDD.n692 VDD.n689 691.758
R20845 VDD.n2331 VDD.n2235 647.574
R20846 VDD.n2351 VDD.n2321 647.574
R20847 VDD.n5276 VDD.n5221 647.574
R20848 VDD.n5305 VDD.n5304 647.574
R20849 VDD.n7042 VDD.n7041 647.574
R20850 VDD.n5277 VDD.n5264 647.574
R20851 VDD.n5312 VDD.n5306 647.574
R20852 VDD.n2332 VDD.n2236 647.574
R20853 VDD.n2367 VDD.n2352 647.574
R20854 VDD.n5278 VDD.n5266 647.574
R20855 VDD.n5378 VDD.n5307 647.574
R20856 VDD.n7835 VDD.n2234 647.574
R20857 VDD.n2353 VDD.n2312 647.574
R20858 VDD.n6578 VDD.n5270 647.574
R20859 VDD.n5942 VDD.n5308 647.574
R20860 VDD.n7833 VDD.n2238 647.574
R20861 VDD.n2331 VDD.n2318 642.269
R20862 VDD.n2369 VDD.n2351 642.269
R20863 VDD.n5282 VDD.n5276 642.269
R20864 VDD.n5305 VDD.n5303 642.269
R20865 VDD.n7041 VDD.n2349 642.269
R20866 VDD.n6371 VDD.n5277 642.269
R20867 VDD.n5311 VDD.n5306 642.269
R20868 VDD.n2332 VDD.n2319 642.269
R20869 VDD.n6634 VDD.n2352 642.269
R20870 VDD.n6369 VDD.n5278 642.269
R20871 VDD.n6310 VDD.n5307 642.269
R20872 VDD.n7134 VDD.n2234 642.269
R20873 VDD.n6632 VDD.n2353 642.269
R20874 VDD.n6578 VDD.n5275 642.269
R20875 VDD.n6312 VDD.n5308 642.269
R20876 VDD.n7132 VDD.n2238 642.269
R20877 VDD.n7087 VDD.n2235 640.197
R20878 VDD.n7039 VDD.n2321 640.197
R20879 VDD.n6576 VDD.n5221 640.197
R20880 VDD.n6397 VDD.n5304 640.197
R20881 VDD.n7042 VDD.n2348 640.197
R20882 VDD.n5281 VDD.n5264 640.197
R20883 VDD.n6395 VDD.n5312 640.197
R20884 VDD.n7085 VDD.n2236 640.197
R20885 VDD.n2368 VDD.n2367 640.197
R20886 VDD.n5280 VDD.n5266 640.197
R20887 VDD.n5378 VDD.n5310 640.197
R20888 VDD.n7835 VDD.n2210 640.197
R20889 VDD.n2357 VDD.n2312 640.197
R20890 VDD.n5279 VDD.n5270 640.197
R20891 VDD.n5942 VDD.n5309 640.197
R20892 VDD.n7833 VDD.n2237 640.197
R20893 VDD.n7087 VDD.n2318 634.891
R20894 VDD.n7039 VDD.n2369 634.891
R20895 VDD.n6576 VDD.n5282 634.891
R20896 VDD.n6397 VDD.n5303 634.891
R20897 VDD.n2349 VDD.n2348 634.891
R20898 VDD.n6371 VDD.n5281 634.891
R20899 VDD.n6395 VDD.n5311 634.891
R20900 VDD.n7085 VDD.n2319 634.891
R20901 VDD.n6634 VDD.n2368 634.891
R20902 VDD.n6369 VDD.n5280 634.891
R20903 VDD.n6310 VDD.n5310 634.891
R20904 VDD.n7134 VDD.n2210 634.891
R20905 VDD.n6632 VDD.n2357 634.891
R20906 VDD.n5279 VDD.n5275 634.891
R20907 VDD.n6312 VDD.n5309 634.891
R20908 VDD.n7132 VDD.n2237 634.891
R20909 VDD.n1550 VDD.n1521 614.001
R20910 VDD.n1550 VDD.n1549 613.338
R20911 VDD.n1552 VDD.n1521 607.537
R20912 VDD.n1552 VDD.n1549 606.872
R20913 VDD.n12614 VDD.n13 477.971
R20914 VDD.n12610 VDD.n16 477.971
R20915 VDD.n12529 VDD.n31 477.971
R20916 VDD.n12522 VDD.n43 477.971
R20917 VDD.n12516 VDD.n96 477.971
R20918 VDD.n12473 VDD.n111 477.971
R20919 VDD.n11027 VDD.n1771 477.971
R20920 VDD.n11006 VDD.n1785 477.971
R20921 VDD.n10999 VDD.n10998 477.971
R20922 VDD.n10994 VDD.n1833 477.971
R20923 VDD.n10951 VDD.n1848 477.971
R20924 VDD.n10944 VDD.n10943 477.971
R20925 VDD.n10939 VDD.n1898 477.971
R20926 VDD.n10896 VDD.n1913 477.971
R20927 VDD.n10889 VDD.n10888 477.971
R20928 VDD.n10884 VDD.n1925 477.971
R20929 VDD.n10841 VDD.n1940 477.971
R20930 VDD.n10834 VDD.n10833 477.971
R20931 VDD.n10829 VDD.n1990 477.971
R20932 VDD.n10783 VDD.n2013 477.971
R20933 VDD.n10776 VDD.n10775 477.971
R20934 VDD.n9157 VDD.n8473 477.971
R20935 VDD.n9033 VDD.n8491 477.971
R20936 VDD.n9014 VDD.n8500 477.971
R20937 VDD.n8936 VDD.n8508 477.971
R20938 VDD.n8883 VDD.n8519 477.971
R20939 VDD.n8805 VDD.n8527 477.971
R20940 VDD.n12460 VDD.n176 477.971
R20941 VDD.n12466 VDD.n123 477.971
R20942 VDD.n9178 VDD.n8460 477.971
R20943 VDD.n12592 VDD.n14 470.842
R20944 VDD.n30 VDD.n17 470.842
R20945 VDD.n12524 VDD.n32 470.842
R20946 VDD.n12521 VDD.n44 470.842
R20947 VDD.n110 VDD.n97 470.842
R20948 VDD.n12468 VDD.n112 470.842
R20949 VDD.n11030 VDD.n1772 470.842
R20950 VDD.n11001 VDD.n1784 470.842
R20951 VDD.n1795 VDD.n1794 470.842
R20952 VDD.n1846 VDD.n1832 470.842
R20953 VDD.n10946 VDD.n1847 470.842
R20954 VDD.n1860 VDD.n1859 470.842
R20955 VDD.n1911 VDD.n1897 470.842
R20956 VDD.n10891 VDD.n1912 470.842
R20957 VDD.n1921 VDD.n1920 470.842
R20958 VDD.n1938 VDD.n1924 470.842
R20959 VDD.n10836 VDD.n1939 470.842
R20960 VDD.n1952 VDD.n1951 470.842
R20961 VDD.n2011 VDD.n1989 470.842
R20962 VDD.n10778 VDD.n2012 470.842
R20963 VDD.n2025 VDD.n2024 470.842
R20964 VDD.n9160 VDD.n8466 470.842
R20965 VDD.n9036 VDD.n8480 470.842
R20966 VDD.n9009 VDD.n8501 470.842
R20967 VDD.n8939 VDD.n8509 470.842
R20968 VDD.n8878 VDD.n8520 470.842
R20969 VDD.n8808 VDD.n8528 470.842
R20970 VDD.n8539 VDD.n177 470.842
R20971 VDD.n12465 VDD.n124 470.842
R20972 VDD.n9182 VDD.n8461 470.842
R20973 VDD.n12614 VDD.n14 470.842
R20974 VDD.n30 VDD.n16 470.842
R20975 VDD.n12524 VDD.n31 470.842
R20976 VDD.n44 VDD.n43 470.842
R20977 VDD.n110 VDD.n96 470.842
R20978 VDD.n12468 VDD.n111 470.842
R20979 VDD.n11027 VDD.n1772 470.842
R20980 VDD.n11001 VDD.n1785 470.842
R20981 VDD.n10998 VDD.n1795 470.842
R20982 VDD.n1846 VDD.n1833 470.842
R20983 VDD.n10946 VDD.n1848 470.842
R20984 VDD.n10943 VDD.n1860 470.842
R20985 VDD.n1911 VDD.n1898 470.842
R20986 VDD.n10891 VDD.n1913 470.842
R20987 VDD.n10888 VDD.n1921 470.842
R20988 VDD.n1938 VDD.n1925 470.842
R20989 VDD.n10836 VDD.n1940 470.842
R20990 VDD.n10833 VDD.n1952 470.842
R20991 VDD.n2011 VDD.n1990 470.842
R20992 VDD.n10778 VDD.n2013 470.842
R20993 VDD.n10775 VDD.n2025 470.842
R20994 VDD.n9157 VDD.n8466 470.842
R20995 VDD.n9033 VDD.n8480 470.842
R20996 VDD.n9014 VDD.n8501 470.842
R20997 VDD.n8936 VDD.n8509 470.842
R20998 VDD.n8883 VDD.n8520 470.842
R20999 VDD.n8805 VDD.n8528 470.842
R21000 VDD.n8539 VDD.n176 470.842
R21001 VDD.n124 VDD.n123 470.842
R21002 VDD.n9182 VDD.n8460 470.842
R21003 VDD.n12592 VDD.n13 469.683
R21004 VDD.n12610 VDD.n17 469.683
R21005 VDD.n12529 VDD.n32 469.683
R21006 VDD.n12522 VDD.n12521 469.683
R21007 VDD.n12516 VDD.n97 469.683
R21008 VDD.n12473 VDD.n112 469.683
R21009 VDD.n11030 VDD.n1771 469.683
R21010 VDD.n11006 VDD.n1784 469.683
R21011 VDD.n10999 VDD.n1794 469.683
R21012 VDD.n10994 VDD.n1832 469.683
R21013 VDD.n10951 VDD.n1847 469.683
R21014 VDD.n10944 VDD.n1859 469.683
R21015 VDD.n10939 VDD.n1897 469.683
R21016 VDD.n10896 VDD.n1912 469.683
R21017 VDD.n10889 VDD.n1920 469.683
R21018 VDD.n10884 VDD.n1924 469.683
R21019 VDD.n10841 VDD.n1939 469.683
R21020 VDD.n10834 VDD.n1951 469.683
R21021 VDD.n10829 VDD.n1989 469.683
R21022 VDD.n10783 VDD.n2012 469.683
R21023 VDD.n10776 VDD.n2024 469.683
R21024 VDD.n9160 VDD.n8473 469.683
R21025 VDD.n9036 VDD.n8491 469.683
R21026 VDD.n9009 VDD.n8500 469.683
R21027 VDD.n8939 VDD.n8508 469.683
R21028 VDD.n8878 VDD.n8519 469.683
R21029 VDD.n8808 VDD.n8527 469.683
R21030 VDD.n12460 VDD.n177 469.683
R21031 VDD.n12466 VDD.n12465 469.683
R21032 VDD.n9178 VDD.n8461 469.683
R21033 VDD.n8078 VDD.n2123 351.805
R21034 VDD.n8078 VDD.n2124 351.639
R21035 VDD.n8076 VDD.n2123 350.479
R21036 VDD.n8076 VDD.n2124 350.313
R21037 VDD.t1667 VDD.t923 338.731
R21038 VDD.t997 VDD.t2302 338.731
R21039 VDD.t695 VDD.t1667 260.622
R21040 VDD.t1191 VDD.t997 260.622
R21041 VDD.t923 VDD.n1521 167.008
R21042 VDD.t2302 VDD.n1549 167.008
R21043 VDD.n1551 VDD.t695 156.792
R21044 VDD.n1551 VDD.t1191 155.268
R21045 VDD.t376 VDD.t1102 142.93
R21046 VDD.t1422 VDD.t375 142.93
R21047 VDD.t1749 VDD.t526 142.93
R21048 VDD.t527 VDD.t2234 142.93
R21049 VDD.t324 VDD.t2488 142.93
R21050 VDD.t323 VDD.t947 142.93
R21051 VDD.t503 VDD.t920 142.93
R21052 VDD.t2779 VDD.t500 142.93
R21053 VDD.t896 VDD.t557 142.93
R21054 VDD.t556 VDD.t700 142.93
R21055 VDD.t647 VDD.t804 142.93
R21056 VDD.t2776 VDD.t1052 142.93
R21057 VDD.t1843 VDD.t2122 142.93
R21058 VDD.t1186 VDD.t2926 142.93
R21059 VDD.t1368 VDD.t490 142.93
R21060 VDD.t488 VDD.t1801 142.93
R21061 VDD.t1381 VDD.t878 142.93
R21062 VDD.t2264 VDD.t1265 142.93
R21063 VDD.t493 VDD.t642 142.93
R21064 VDD.t2575 VDD.t492 142.93
R21065 VDD.t958 VDD.t3748 142.93
R21066 VDD.t3679 VDD.t1373 142.93
R21067 VDD.t496 VDD.t1551 142.93
R21068 VDD.t497 VDD.t652 142.93
R21069 VDD.t290 VDD.t1716 142.93
R21070 VDD.t1209 VDD.t291 142.93
R21071 VDD.t1180 VDD.t1497 142.93
R21072 VDD.t3424 VDD.t680 142.93
R21073 VDD.t12 VDD.t2352 142.93
R21074 VDD.t351 VDD.t1352 142.93
R21075 VDD.t331 VDD.t1484 142.93
R21076 VDD.t328 VDD.t1089 142.93
R21077 VDD.t1293 VDD.t1572 142.93
R21078 VDD.t1158 VDD.t1906 142.93
R21079 VDD.t1517 VDD.t528 142.93
R21080 VDD.t529 VDD.t1613 142.93
R21081 VDD.t1998 VDD.t629 142.93
R21082 VDD.t798 VDD.t751 142.93
R21083 VDD.t551 VDD.t1655 142.93
R21084 VDD.t831 VDD.t549 142.93
R21085 VDD.t728 VDD.t1489 142.93
R21086 VDD.t2731 VDD.t1823 142.93
R21087 VDD.t2100 VDD.t1789 142.93
R21088 VDD.t2347 VDD.t614 142.93
R21089 VDD.t2061 VDD.t795 142.93
R21090 VDD.t1411 VDD.t2254 142.93
R21091 VDD.t901 VDD.t3 142.93
R21092 VDD.t0 VDD.t1492 142.93
R21093 VDD.t2467 VDD.t547 142.93
R21094 VDD.t544 VDD.t2103 142.93
R21095 VDD.t634 VDD.t334 142.93
R21096 VDD.t322 VDD.t670 142.93
R21097 VDD.t845 VDD.t2328 142.93
R21098 VDD.t2561 VDD.t839 142.93
R21099 VDD.t2082 VDD.t1798 142.93
R21100 VDD.t564 VDD.t2164 142.93
R21101 VDD.t2159 VDD.t1895 142.93
R21102 VDD.t683 VDD.t2257 142.93
R21103 VDD.t554 VDD.t2146 142.93
R21104 VDD.t2402 VDD.t626 142.93
R21105 VDD.t1102 VDD.t968 96.8792
R21106 VDD.t373 VDD.t376 96.8792
R21107 VDD.t375 VDD.t374 96.8792
R21108 VDD.t1644 VDD.t1422 96.8792
R21109 VDD.t1357 VDD.t1749 96.8792
R21110 VDD.t526 VDD.t525 96.8792
R21111 VDD.t524 VDD.t527 96.8792
R21112 VDD.t2234 VDD.t1115 96.8792
R21113 VDD.t2488 VDD.t855 96.8792
R21114 VDD.t325 VDD.t324 96.8792
R21115 VDD.t301 VDD.t323 96.8792
R21116 VDD.t947 VDD.t748 96.8792
R21117 VDD.t920 VDD.t792 96.8792
R21118 VDD.t502 VDD.t503 96.8792
R21119 VDD.t500 VDD.t501 96.8792
R21120 VDD.t1145 VDD.t2779 96.8792
R21121 VDD.t938 VDD.t896 96.8792
R21122 VDD.t557 VDD.t559 96.8792
R21123 VDD.t558 VDD.t556 96.8792
R21124 VDD.t700 VDD.t783 96.8792
R21125 VDD.t804 VDD.t1660 96.8792
R21126 VDD.t1445 VDD.t647 96.8792
R21127 VDD.t3355 VDD.t2776 96.8792
R21128 VDD.t1052 VDD.t2682 96.8792
R21129 VDD.t2122 VDD.t858 96.8792
R21130 VDD.t575 VDD.t1843 96.8792
R21131 VDD.t2926 VDD.t3571 96.8792
R21132 VDD.t908 VDD.t1186 96.8792
R21133 VDD.t2572 VDD.t1368 96.8792
R21134 VDD.t490 VDD.t491 96.8792
R21135 VDD.t489 VDD.t488 96.8792
R21136 VDD.t1801 VDD.t1959 96.8792
R21137 VDD.t878 VDD.t1938 96.8792
R21138 VDD.t869 VDD.t1381 96.8792
R21139 VDD.t1341 VDD.t2264 96.8792
R21140 VDD.t1265 VDD.t1212 96.8792
R21141 VDD.t642 VDD.t801 96.8792
R21142 VDD.t495 VDD.t493 96.8792
R21143 VDD.t492 VDD.t494 96.8792
R21144 VDD.t1376 VDD.t2575 96.8792
R21145 VDD.t816 VDD.t958 96.8792
R21146 VDD.t3748 VDD.t2923 96.8792
R21147 VDD.t1408 VDD.t3679 96.8792
R21148 VDD.t1373 VDD.t1183 96.8792
R21149 VDD.t1551 VDD.t677 96.8792
R21150 VDD.t498 VDD.t496 96.8792
R21151 VDD.t512 VDD.t497 96.8792
R21152 VDD.t652 VDD.t1442 96.8792
R21153 VDD.t1716 VDD.t1167 96.8792
R21154 VDD.t293 VDD.t290 96.8792
R21155 VDD.t291 VDD.t292 96.8792
R21156 VDD.t1084 VDD.t1209 96.8792
R21157 VDD.t1325 VDD.t1180 96.8792
R21158 VDD.t1497 VDD.t1713 96.8792
R21159 VDD.t3614 VDD.t3424 96.8792
R21160 VDD.t680 VDD.t933 96.8792
R21161 VDD.t2352 VDD.t602 96.8792
R21162 VDD.t304 VDD.t12 96.8792
R21163 VDD.t13 VDD.t351 96.8792
R21164 VDD.t1352 VDD.t758 96.8792
R21165 VDD.t1484 VDD.t836 96.8792
R21166 VDD.t329 VDD.t331 96.8792
R21167 VDD.t330 VDD.t328 96.8792
R21168 VDD.t1089 VDD.t1782 96.8792
R21169 VDD.t1572 VDD.t1221 96.8792
R21170 VDD.t1542 VDD.t1293 96.8792
R21171 VDD.t1906 VDD.t848 96.8792
R21172 VDD.t1886 VDD.t1158 96.8792
R21173 VDD.t1302 VDD.t1517 96.8792
R21174 VDD.t528 VDD.t530 96.8792
R21175 VDD.t535 VDD.t529 96.8792
R21176 VDD.t1613 VDD.t689 96.8792
R21177 VDD.t629 VDD.t639 96.8792
R21178 VDD.t2243 VDD.t1998 96.8792
R21179 VDD.t2425 VDD.t798 96.8792
R21180 VDD.t751 VDD.t979 96.8792
R21181 VDD.t1655 VDD.t1427 96.8792
R21182 VDD.t550 VDD.t551 96.8792
R21183 VDD.t549 VDD.t548 96.8792
R21184 VDD.t623 VDD.t831 96.8792
R21185 VDD.t1508 VDD.t728 96.8792
R21186 VDD.t1489 VDD.t1710 96.8792
R21187 VDD.t1852 VDD.t2731 96.8792
R21188 VDD.t1823 VDD.t2079 96.8792
R21189 VDD.t1789 VDD.t1055 96.8792
R21190 VDD.t2385 VDD.t2100 96.8792
R21191 VDD.t2046 VDD.t2347 96.8792
R21192 VDD.t614 VDD.t826 96.8792
R21193 VDD.t795 VDD.t1130 96.8792
R21194 VDD.t2814 VDD.t2061 96.8792
R21195 VDD.t2254 VDD.t2023 96.8792
R21196 VDD.t813 VDD.t1411 96.8792
R21197 VDD.t1198 VDD.t901 96.8792
R21198 VDD.t3 VDD.t6 96.8792
R21199 VDD.t1 VDD.t0 96.8792
R21200 VDD.t1492 VDD.t1336 96.8792
R21201 VDD.t1268 VDD.t2467 96.8792
R21202 VDD.t547 VDD.t545 96.8792
R21203 VDD.t546 VDD.t544 96.8792
R21204 VDD.t2103 VDD.t1018 96.8792
R21205 VDD.t1820 VDD.t634 96.8792
R21206 VDD.t334 VDD.t296 96.8792
R21207 VDD.t420 VDD.t322 96.8792
R21208 VDD.t670 VDD.t982 96.8792
R21209 VDD.t1254 VDD.t845 96.8792
R21210 VDD.t2328 VDD.t710 96.8792
R21211 VDD.t2291 VDD.t2561 96.8792
R21212 VDD.t839 VDD.t1045 96.8792
R21213 VDD.t1826 VDD.t2082 96.8792
R21214 VDD.t1798 VDD.t2064 96.8792
R21215 VDD.t2193 VDD.t564 96.8792
R21216 VDD.t2164 VDD.t2450 96.8792
R21217 VDD.t1919 VDD.t2159 96.8792
R21218 VDD.t1895 VDD.t2131 96.8792
R21219 VDD.t2305 VDD.t683 96.8792
R21220 VDD.t2257 VDD.t607 96.8792
R21221 VDD.t2146 VDD.t1869 96.8792
R21222 VDD.t2091 VDD.t554 96.8792
R21223 VDD.t626 VDD.t552 96.8792
R21224 VDD.t723 VDD.t2402 96.8792
R21225 VDD.t572 VDD.t404 85.1494
R21226 VDD.t15 VDD.t913 85.1494
R21227 VDD.t37 VDD.t928 85.1494
R21228 VDD.t389 VDD.t965 81.7244
R21229 VDD.t968 VDD.n1771 81.1238
R21230 VDD.t758 VDD.n2025 81.1238
R21231 VDD.t836 VDD.n13 81.1238
R21232 VDD.n9182 VDD.t723 81.1238
R21233 VDD.n1786 VDD.t1644 81.017
R21234 VDD.n11005 VDD.t1357 81.017
R21235 VDD.t1115 VDD.n11002 81.017
R21236 VDD.t855 VDD.n1787 81.017
R21237 VDD.t748 VDD.n10996 81.017
R21238 VDD.n10995 VDD.t792 81.017
R21239 VDD.n1851 VDD.t1145 81.017
R21240 VDD.n10950 VDD.t938 81.017
R21241 VDD.t783 VDD.n10947 81.017
R21242 VDD.t1660 VDD.n1852 81.017
R21243 VDD.t2682 VDD.n10941 81.017
R21244 VDD.n10940 VDD.t858 81.017
R21245 VDD.n1916 VDD.t908 81.017
R21246 VDD.n10895 VDD.t2572 81.017
R21247 VDD.t1959 VDD.n10892 81.017
R21248 VDD.t1938 VDD.n1917 81.017
R21249 VDD.t1212 VDD.n10886 81.017
R21250 VDD.n10885 VDD.t801 81.017
R21251 VDD.n1943 VDD.t1376 81.017
R21252 VDD.n10840 VDD.t816 81.017
R21253 VDD.t1183 VDD.n10837 81.017
R21254 VDD.t677 VDD.n1944 81.017
R21255 VDD.t1442 VDD.n10831 81.017
R21256 VDD.n10830 VDD.t1167 81.017
R21257 VDD.n2016 VDD.t1084 81.017
R21258 VDD.n10782 VDD.t1325 81.017
R21259 VDD.t933 VDD.n10779 81.017
R21260 VDD.t602 VDD.n2017 81.017
R21261 VDD.t1782 VDD.n12612 81.017
R21262 VDD.n12611 VDD.t1221 81.017
R21263 VDD.n35 VDD.t1886 81.017
R21264 VDD.n12528 VDD.t1302 81.017
R21265 VDD.t689 VDD.n12525 81.017
R21266 VDD.t639 VDD.n36 81.017
R21267 VDD.t979 VDD.n12518 81.017
R21268 VDD.n12517 VDD.t1427 81.017
R21269 VDD.n115 VDD.t623 81.017
R21270 VDD.n12472 VDD.t1508 81.017
R21271 VDD.t2079 VDD.n12469 81.017
R21272 VDD.t1055 VDD.n116 81.017
R21273 VDD.t826 VDD.n12462 81.017
R21274 VDD.n12461 VDD.t1130 81.017
R21275 VDD.n8538 VDD.t813 81.017
R21276 VDD.n8537 VDD.t1198 81.017
R21277 VDD.t1336 VDD.n8530 81.017
R21278 VDD.n8529 VDD.t1268 81.017
R21279 VDD.t1018 VDD.n8881 81.017
R21280 VDD.n8880 VDD.t1820 81.017
R21281 VDD.t982 VDD.n8511 81.017
R21282 VDD.n8510 VDD.t1254 81.017
R21283 VDD.t1045 VDD.n9012 81.017
R21284 VDD.n9011 VDD.t1826 81.017
R21285 VDD.t2450 VDD.n8493 81.017
R21286 VDD.n8492 VDD.t1919 81.017
R21287 VDD.t607 VDD.n8462 81.017
R21288 VDD.t1869 VDD.n9179 81.017
R21289 VDD.t19 VDD.t30 79.7265
R21290 VDD.t17 VDD.t35 79.7265
R21291 VDD.t406 VDD.t389 79.5362
R21292 VDD.n11029 VDD.t373 70.2717
R21293 VDD.t525 VDD.n11004 70.2717
R21294 VDD.n1831 VDD.t325 70.2717
R21295 VDD.n1849 VDD.t502 70.2717
R21296 VDD.t559 VDD.n10949 70.2717
R21297 VDD.n1896 VDD.t1445 70.2717
R21298 VDD.n1914 VDD.t575 70.2717
R21299 VDD.t491 VDD.n10894 70.2717
R21300 VDD.n1923 VDD.t869 70.2717
R21301 VDD.n1941 VDD.t495 70.2717
R21302 VDD.t2923 VDD.n10839 70.2717
R21303 VDD.n1988 VDD.t498 70.2717
R21304 VDD.n2014 VDD.t293 70.2717
R21305 VDD.t1713 VDD.n10781 70.2717
R21306 VDD.n10773 VDD.t304 70.2717
R21307 VDD.n15 VDD.t329 70.2717
R21308 VDD.n33 VDD.t1542 70.2717
R21309 VDD.t530 VDD.n12527 70.2717
R21310 VDD.n12520 VDD.t2243 70.2717
R21311 VDD.n113 VDD.t550 70.2717
R21312 VDD.t1710 VDD.n12471 70.2717
R21313 VDD.n12464 VDD.t2385 70.2717
R21314 VDD.n8535 VDD.t2814 70.2717
R21315 VDD.n8807 VDD.t6 70.2717
R21316 VDD.n8879 VDD.t545 70.2717
R21317 VDD.n8938 VDD.t296 70.2717
R21318 VDD.n9010 VDD.t710 70.2717
R21319 VDD.n9035 VDD.t2064 70.2717
R21320 VDD.n9159 VDD.t2131 70.2717
R21321 VDD.n9180 VDD.t2091 70.2717
R21322 VDD.n11028 VDD.t374 64.1315
R21323 VDD.n11003 VDD.t524 64.1315
R21324 VDD.n10997 VDD.t301 64.1315
R21325 VDD.t501 VDD.n1850 64.1315
R21326 VDD.n10948 VDD.t558 64.1315
R21327 VDD.n10942 VDD.t3355 64.1315
R21328 VDD.t3571 VDD.n1915 64.1315
R21329 VDD.n10893 VDD.t489 64.1315
R21330 VDD.n10887 VDD.t1341 64.1315
R21331 VDD.t494 VDD.n1942 64.1315
R21332 VDD.n10838 VDD.t1408 64.1315
R21333 VDD.n10832 VDD.t512 64.1315
R21334 VDD.t292 VDD.n2015 64.1315
R21335 VDD.n10780 VDD.t3614 64.1315
R21336 VDD.n10774 VDD.t13 64.1315
R21337 VDD.n12613 VDD.t330 64.1315
R21338 VDD.t848 VDD.n34 64.1315
R21339 VDD.n12526 VDD.t535 64.1315
R21340 VDD.n12519 VDD.t2425 64.1315
R21341 VDD.t548 VDD.n114 64.1315
R21342 VDD.n12470 VDD.t1852 64.1315
R21343 VDD.n12463 VDD.t2046 64.1315
R21344 VDD.t2023 VDD.n8536 64.1315
R21345 VDD.n8806 VDD.t1 64.1315
R21346 VDD.n8882 VDD.t546 64.1315
R21347 VDD.n8937 VDD.t420 64.1315
R21348 VDD.n9013 VDD.t2291 64.1315
R21349 VDD.n9034 VDD.t2193 64.1315
R21350 VDD.n9158 VDD.t2305 64.1315
R21351 VDD.t552 VDD.n9181 64.1315
R21352 VDD.t404 VDD.t401 54.0391
R21353 VDD.t41 VDD.t15 54.0391
R21354 VDD.t21 VDD.t19 54.0391
R21355 VDD.t26 VDD.t17 54.0391
R21356 VDD.t35 VDD.t28 54.0391
R21357 VDD.t28 VDD.t23 54.0391
R21358 VDD.t23 VDD.t37 54.0391
R21359 VDD.n7995 VDD.t30 50.3287
R21360 VDD.n6633 VDD.n5268 46.8594
R21361 VDD.t965 VDD.n2123 45.4522
R21362 VDD.t928 VDD.n2188 45.3596
R21363 VDD.n2354 VDD.t572 45.2864
R21364 VDD.t913 VDD.n2355 45.2864
R21365 VDD.n2356 VDD.t21 42.0517
R21366 VDD.t686 VDD.t471 38.7904
R21367 VDD.t745 VDD.t469 38.7904
R21368 VDD.t692 VDD.t467 38.7904
R21369 VDD.t660 VDD.t470 38.7904
R21370 VDD.t881 VDD.t473 38.7904
R21371 VDD.t468 VDD.t561 38.7904
R21372 VDD.t317 VDD.t567 38.7904
R21373 VDD.t309 VDD.t821 38.7904
R21374 VDD.t316 VDD.t703 38.7904
R21375 VDD.t657 VDD.t308 38.7904
R21376 VDD.t665 VDD.t312 38.7904
R21377 VDD.t578 VDD.t306 38.7904
R21378 VDD.n8077 VDD.t401 37.9607
R21379 VDD.t471 VDD.t426 36.32
R21380 VDD.t469 VDD.t422 36.32
R21381 VDD.t467 VDD.t424 36.32
R21382 VDD.t470 VDD.t428 36.32
R21383 VDD.t473 VDD.t438 36.32
R21384 VDD.t433 VDD.t468 36.32
R21385 VDD.t315 VDD.t317 36.32
R21386 VDD.t318 VDD.t309 36.32
R21387 VDD.t332 VDD.t316 36.32
R21388 VDD.t308 VDD.t313 36.32
R21389 VDD.t312 VDD.t311 36.32
R21390 VDD.t306 VDD.t321 36.32
R21391 VDD.t590 VDD.t392 31.8205
R21392 VDD.t842 VDD.t394 31.8205
R21393 VDD.t620 VDD.t390 31.8205
R21394 VDD.t397 VDD.t617 31.8205
R21395 VDD.t889 VDD.t85 31.8205
R21396 VDD.t73 VDD.t587 31.8205
R21397 VDD.t52 VDD.t886 31.8205
R21398 VDD.t58 VDD.t597 31.8205
R21399 VDD.t405 VDD.t409 29.7939
R21400 VDD.t396 VDD.t400 29.7939
R21401 VDD.t402 VDD.t403 29.7939
R21402 VDD.t395 VDD.t399 29.7939
R21403 VDD.t63 VDD.t81 29.7939
R21404 VDD.t67 VDD.t50 29.7939
R21405 VDD.t79 VDD.t65 29.7939
R21406 VDD.t61 VDD.t123 29.7939
R21407 VDD.n10996 VDD.n10995 29.1665
R21408 VDD.n10941 VDD.n10940 29.1665
R21409 VDD.n10886 VDD.n10885 29.1665
R21410 VDD.n10831 VDD.n10830 29.1665
R21411 VDD.n12525 VDD.n36 29.1665
R21412 VDD.n12469 VDD.n116 29.1665
R21413 VDD.n8530 VDD.n8529 29.1665
R21414 VDD.n9012 VDD.n9011 29.1665
R21415 VDD.t426 VDD.t431 24.618
R21416 VDD.t424 VDD.t441 24.618
R21417 VDD.t438 VDD.t443 24.618
R21418 VDD.t319 VDD.t315 24.618
R21419 VDD.t320 VDD.t332 24.618
R21420 VDD.t311 VDD.t314 24.618
R21421 VDD.n11005 VDD.n1786 24.5613
R21422 VDD.n11002 VDD.n1787 24.5613
R21423 VDD.n10950 VDD.n1851 24.5613
R21424 VDD.n10947 VDD.n1852 24.5613
R21425 VDD.n10895 VDD.n1916 24.5613
R21426 VDD.n10892 VDD.n1917 24.5613
R21427 VDD.n10840 VDD.n1943 24.5613
R21428 VDD.n10837 VDD.n1944 24.5613
R21429 VDD.n10782 VDD.n2016 24.5613
R21430 VDD.n10779 VDD.n2017 24.5613
R21431 VDD.n12612 VDD.n12611 24.5613
R21432 VDD.n12528 VDD.n35 24.5613
R21433 VDD.n12518 VDD.n12517 24.5613
R21434 VDD.n12472 VDD.n115 24.5613
R21435 VDD.n12462 VDD.n12461 24.5613
R21436 VDD.n8538 VDD.n8537 24.5613
R21437 VDD.n8881 VDD.n8880 24.5613
R21438 VDD.n8511 VDD.n8510 24.5613
R21439 VDD.n8493 VDD.n8492 24.5613
R21440 VDD.n9179 VDD.n8462 24.5613
R21441 VDD.n1742 VDD.t422 24.0112
R21442 VDD.n1718 VDD.t428 24.0112
R21443 VDD.n1414 VDD.t433 24.0112
R21444 VDD.n1356 VDD.t318 24.0112
R21445 VDD.n1349 VDD.t313 24.0112
R21446 VDD.n1652 VDD.t321 24.0112
R21447 VDD.n690 VDD.t686 20.6307
R21448 VDD.n709 VDD.t745 20.6307
R21449 VDD.n1719 VDD.t692 20.6307
R21450 VDD.n874 VDD.t660 20.6307
R21451 VDD.n1415 VDD.t881 20.6307
R21452 VDD.n1429 VDD.t561 20.6307
R21453 VDD.n1428 VDD.t567 20.6307
R21454 VDD.t821 VDD.n1354 20.6307
R21455 VDD.t703 VDD.n1084 20.6307
R21456 VDD.n1346 VDD.t657 20.6307
R21457 VDD.n1345 VDD.t665 20.6307
R21458 VDD.n763 VDD.t578 20.6307
R21459 VDD.t392 VDD.t415 20.1946
R21460 VDD.t415 VDD.t393 20.1946
R21461 VDD.t393 VDD.t405 20.1946
R21462 VDD.t400 VDD.t412 20.1946
R21463 VDD.t411 VDD.t396 20.1946
R21464 VDD.t398 VDD.t411 20.1946
R21465 VDD.t394 VDD.t398 20.1946
R21466 VDD.t390 VDD.t414 20.1946
R21467 VDD.t414 VDD.t391 20.1946
R21468 VDD.t391 VDD.t402 20.1946
R21469 VDD.t408 VDD.t395 20.1946
R21470 VDD.t399 VDD.t407 20.1946
R21471 VDD.t407 VDD.t410 20.1946
R21472 VDD.t410 VDD.t397 20.1946
R21473 VDD.t85 VDD.t140 20.1946
R21474 VDD.t140 VDD.t71 20.1946
R21475 VDD.t71 VDD.t63 20.1946
R21476 VDD.t99 VDD.t67 20.1946
R21477 VDD.t50 VDD.t56 20.1946
R21478 VDD.t56 VDD.t118 20.1946
R21479 VDD.t118 VDD.t73 20.1946
R21480 VDD.t69 VDD.t52 20.1946
R21481 VDD.t137 VDD.t69 20.1946
R21482 VDD.t65 VDD.t137 20.1946
R21483 VDD.t76 VDD.t61 20.1946
R21484 VDD.t123 VDD.t54 20.1946
R21485 VDD.t54 VDD.t125 20.1946
R21486 VDD.t125 VDD.t58 20.1946
R21487 VDD.n6396 VDD.t409 19.0569
R21488 VDD.n6577 VDD.t403 19.0569
R21489 VDD.n7040 VDD.t81 19.0569
R21490 VDD.n7086 VDD.t79 19.0569
R21491 VDD.n6311 VDD.t590 16.9237
R21492 VDD.n5376 VDD.t842 16.9237
R21493 VDD.n6370 VDD.t620 16.9237
R21494 VDD.t617 VDD.n5268 16.9237
R21495 VDD.n6633 VDD.t889 16.9237
R21496 VDD.n7133 VDD.t886 16.9237
R21497 VDD.n7834 VDD.t597 16.9237
R21498 VDD.n8077 VDD.t406 16.0789
R21499 VDD.t587 VDD.n2356 15.3594
R21500 VDD.n2355 VDD.n2354 13.7004
R21501 VDD.n2356 VDD.t41 11.9879
R21502 VDD.n696 VDD.t486 10.8219
R21503 VDD.n949 VDD.t475 10.378
R21504 VDD.n1448 VDD.t387 9.30374
R21505 VDD.n11029 VDD.n11028 8.52856
R21506 VDD.n11004 VDD.n11003 8.52856
R21507 VDD.n10997 VDD.n1831 8.52856
R21508 VDD.n1850 VDD.n1849 8.52856
R21509 VDD.n10949 VDD.n10948 8.52856
R21510 VDD.n10942 VDD.n1896 8.52856
R21511 VDD.n1915 VDD.n1914 8.52856
R21512 VDD.n10894 VDD.n10893 8.52856
R21513 VDD.n10887 VDD.n1923 8.52856
R21514 VDD.n1942 VDD.n1941 8.52856
R21515 VDD.n10839 VDD.n10838 8.52856
R21516 VDD.n10832 VDD.n1988 8.52856
R21517 VDD.n2015 VDD.n2014 8.52856
R21518 VDD.n10781 VDD.n10780 8.52856
R21519 VDD.n10774 VDD.n10773 8.52856
R21520 VDD.n12613 VDD.n15 8.52856
R21521 VDD.n34 VDD.n33 8.52856
R21522 VDD.n12527 VDD.n12526 8.52856
R21523 VDD.n12520 VDD.n12519 8.52856
R21524 VDD.n114 VDD.n113 8.52856
R21525 VDD.n12471 VDD.n12470 8.52856
R21526 VDD.n12464 VDD.n12463 8.52856
R21527 VDD.n8536 VDD.n8535 8.52856
R21528 VDD.n8807 VDD.n8806 8.52856
R21529 VDD.n8882 VDD.n8879 8.52856
R21530 VDD.n8938 VDD.n8937 8.52856
R21531 VDD.n9013 VDD.n9010 8.52856
R21532 VDD.n9035 VDD.n9034 8.52856
R21533 VDD.n9159 VDD.n9158 8.52856
R21534 VDD.n9181 VDD.n9180 8.52856
R21535 VDD.n1442 VDD.t3074 8.19583
R21536 VDD.n1478 VDD.t2765 8.14522
R21537 VDD.t1069 VDD.n1611 8.14522
R21538 VDD.n1609 VDD.t3836 8.14522
R21539 VDD.n1477 VDD.t4070 8.14522
R21540 VDD.t1171 VDD.n1751 8.11081
R21541 VDD VDD.t4000 8.10685
R21542 VDD.n1752 VDD.t1171 8.10567
R21543 VDD.n969 VDD.t3581 8.10567
R21544 VDD.t3581 VDD.n682 8.10567
R21545 VDD.n971 VDD.t2546 8.10567
R21546 VDD.t2546 VDD.n970 8.10567
R21547 VDD.n973 VDD.t2669 8.10567
R21548 VDD.t2669 VDD.n972 8.10567
R21549 VDD.n975 VDD.t1433 8.10567
R21550 VDD.t1433 VDD.n974 8.10567
R21551 VDD.n977 VDD.t1561 8.10567
R21552 VDD.t1561 VDD.n976 8.10567
R21553 VDD.n987 VDD.t4610 8.10567
R21554 VDD.t4610 VDD.n986 8.10567
R21555 VDD.n989 VDD.t808 8.10567
R21556 VDD.t808 VDD.n988 8.10567
R21557 VDD.n991 VDD.t3846 8.10567
R21558 VDD.t3846 VDD.n990 8.10567
R21559 VDD.n993 VDD.t3978 8.10567
R21560 VDD.t3978 VDD.n992 8.10567
R21561 VDD.n995 VDD.t2932 8.10567
R21562 VDD.t2932 VDD.n994 8.10567
R21563 VDD.n997 VDD.t940 8.10567
R21564 VDD.t940 VDD.n996 8.10567
R21565 VDD.n1006 VDD.t685 8.10567
R21566 VDD.t685 VDD.n1005 8.10567
R21567 VDD.n1008 VDD.t3330 8.10567
R21568 VDD.t3330 VDD.n1007 8.10567
R21569 VDD.n1010 VDD.t2227 8.10567
R21570 VDD.t2227 VDD.n1009 8.10567
R21571 VDD.n1012 VDD.t2623 8.10567
R21572 VDD.t2623 VDD.n1011 8.10567
R21573 VDD.n1014 VDD.t2500 8.10567
R21574 VDD.t2500 VDD.n1013 8.10567
R21575 VDD.n1016 VDD.t2629 8.10567
R21576 VDD.t2629 VDD.n1015 8.10567
R21577 VDD.t1399 VDD.n1030 8.10567
R21578 VDD.n1031 VDD.t1399 8.10567
R21579 VDD.t1512 VDD.n1028 8.10567
R21580 VDD.n1029 VDD.t1512 8.10567
R21581 VDD.t4544 VDD.n1026 8.10567
R21582 VDD.n1027 VDD.t4544 8.10567
R21583 VDD.t2567 VDD.n1024 8.10567
R21584 VDD.n1025 VDD.t2567 8.10567
R21585 VDD.t1343 VDD.n1022 8.10567
R21586 VDD.n1023 VDD.t1343 8.10567
R21587 VDD.t4000 VDD.n12643 8.10567
R21588 VDD.n12563 VDD.t1483 8.10567
R21589 VDD.n12563 VDD.t835 8.10567
R21590 VDD.n12566 VDD.t1849 8.10567
R21591 VDD.n12566 VDD.t1164 8.10567
R21592 VDD.n12567 VDD.t2563 8.10567
R21593 VDD.n12567 VDD.t1767 8.10567
R21594 VDD.n12573 VDD.t1862 8.10567
R21595 VDD.n12573 VDD.t1175 8.10567
R21596 VDD.n12574 VDD.t2297 8.10567
R21597 VDD.n12574 VDD.t1537 8.10567
R21598 VDD.n12577 VDD.t3852 8.10567
R21599 VDD.n12577 VDD.t3218 8.10567
R21600 VDD.n8633 VDD.t1809 8.10567
R21601 VDD.n8634 VDD.t2641 8.10567
R21602 VDD.n12617 VDD.t1467 8.10567
R21603 VDD.n11 VDD.t2665 8.10567
R21604 VDD.n8630 VDD.t1571 8.10567
R21605 VDD.n8630 VDD.t3124 8.10567
R21606 VDD.n8627 VDD.t1940 8.10567
R21607 VDD.n8627 VDD.t3438 8.10567
R21608 VDD.n8626 VDD.t2653 8.10567
R21609 VDD.n8626 VDD.t4044 8.10567
R21610 VDD.n12606 VDD.t1967 8.10567
R21611 VDD.n12606 VDD.t3448 8.10567
R21612 VDD.n12605 VDD.t2416 8.10567
R21613 VDD.n12605 VDD.t3806 8.10567
R21614 VDD.n12602 VDD.t3944 8.10567
R21615 VDD.n12602 VDD.t1220 8.10567
R21616 VDD.n8630 VDD.t1781 8.10567
R21617 VDD.n8630 VDD.t2996 8.10567
R21618 VDD.n8627 VDD.t2184 8.10567
R21619 VDD.n8627 VDD.t3298 8.10567
R21620 VDD.n8626 VDD.t2864 8.10567
R21621 VDD.n8626 VDD.t3872 8.10567
R21622 VDD.n12606 VDD.t2207 8.10567
R21623 VDD.n12606 VDD.t3308 8.10567
R21624 VDD.n12605 VDD.t2645 8.10567
R21625 VDD.n12605 VDD.t3638 8.10567
R21626 VDD.n12602 VDD.t4172 8.10567
R21627 VDD.n12602 VDD.t1088 8.10567
R21628 VDD.n12555 VDD.t4188 8.10567
R21629 VDD.n12595 VDD.t755 8.10567
R21630 VDD.n12556 VDD.t3828 8.10567
R21631 VDD.n12588 VDD.t780 8.10567
R21632 VDD.n12545 VDD.t4266 8.10567
R21633 VDD.n25 VDD.t847 8.10567
R21634 VDD.n12551 VDD.t3916 8.10567
R21635 VDD.n24 VDD.t1292 8.10567
R21636 VDD.n8661 VDD.t3371 8.10567
R21637 VDD.n8661 VDD.t3208 8.10567
R21638 VDD.n8658 VDD.t3719 8.10567
R21639 VDD.n8658 VDD.t3508 8.10567
R21640 VDD.n8657 VDD.t4328 8.10567
R21641 VDD.n8657 VDD.t4134 8.10567
R21642 VDD.n12534 VDD.t3735 8.10567
R21643 VDD.n12534 VDD.t3528 8.10567
R21644 VDD.n12535 VDD.t4128 8.10567
R21645 VDD.n12535 VDD.t3892 8.10567
R21646 VDD.n12539 VDD.t1516 8.10567
R21647 VDD.n12539 VDD.t1301 8.10567
R21648 VDD.n8661 VDD.t1885 8.10567
R21649 VDD.n8661 VDD.t3064 8.10567
R21650 VDD.n8658 VDD.t2288 8.10567
R21651 VDD.n8658 VDD.t3357 8.10567
R21652 VDD.n8657 VDD.t2960 8.10567
R21653 VDD.n8657 VDD.t3974 8.10567
R21654 VDD.n12534 VDD.t2321 8.10567
R21655 VDD.n12534 VDD.t3373 8.10567
R21656 VDD.n12535 VDD.t2739 8.10567
R21657 VDD.n12535 VDD.t3741 8.10567
R21658 VDD.n12539 VDD.t4252 8.10567
R21659 VDD.n12539 VDD.t1157 8.10567
R21660 VDD.n8621 VDD.t1905 8.10567
R21661 VDD.n8651 VDD.t2735 8.10567
R21662 VDD.n8622 VDD.t1541 8.10567
R21663 VDD.n8645 VDD.t3190 8.10567
R21664 VDD.n8619 VDD.t3681 8.10567
R21665 VDD.n8672 VDD.t730 8.10567
R21666 VDD.n8620 VDD.t3346 8.10567
R21667 VDD.n8666 VDD.t766 8.10567
R21668 VDD.n8616 VDD.t4064 8.10567
R21669 VDD.n8616 VDD.t3842 8.10567
R21670 VDD.n8613 VDD.t4390 8.10567
R21671 VDD.n8613 VDD.t4212 8.10567
R21672 VDD.n8612 VDD.t893 8.10567
R21673 VDD.n8612 VDD.t638 8.10567
R21674 VDD.n80 VDD.t4404 8.10567
R21675 VDD.n80 VDD.t4230 8.10567
R21676 VDD.n81 VDD.t628 8.10567
R21677 VDD.n81 VDD.t4550 8.10567
R21678 VDD.n85 VDD.t2266 8.10567
R21679 VDD.n85 VDD.t2033 8.10567
R21680 VDD.n8616 VDD.t688 8.10567
R21681 VDD.n8616 VDD.t3468 8.10567
R21682 VDD.n8613 VDD.t1059 8.10567
R21683 VDD.n8613 VDD.t3800 8.10567
R21684 VDD.n8612 VDD.t1650 8.10567
R21685 VDD.n8612 VDD.t4400 8.10567
R21686 VDD.n80 VDD.t1077 8.10567
R21687 VDD.n80 VDD.t3820 8.10567
R21688 VDD.n81 VDD.t1417 8.10567
R21689 VDD.n81 VDD.t4220 8.10567
R21690 VDD.n85 VDD.t3104 8.10567
R21691 VDD.n85 VDD.t1612 8.10567
R21692 VDD.n73 VDD.t1854 8.10567
R21693 VDD.n54 VDD.t3128 8.10567
R21694 VDD.n47 VDD.t1494 8.10567
R21695 VDD.n48 VDD.t3152 8.10567
R21696 VDD.n12499 VDD.t797 8.10567
R21697 VDD.n12501 VDD.t2424 8.10567
R21698 VDD.n45 VDD.t2242 8.10567
R21699 VDD.n91 VDD.t1997 8.10567
R21700 VDD.n8694 VDD.t1654 8.10567
R21701 VDD.n8694 VDD.t1426 8.10567
R21702 VDD.n8691 VDD.t2035 8.10567
R21703 VDD.n8691 VDD.t1777 8.10567
R21704 VDD.n8690 VDD.t2724 8.10567
R21705 VDD.n8690 VDD.t2512 8.10567
R21706 VDD.n12512 VDD.t2056 8.10567
R21707 VDD.n12512 VDD.t1791 8.10567
R21708 VDD.n12511 VDD.t2502 8.10567
R21709 VDD.n12511 VDD.t2223 8.10567
R21710 VDD.n12508 VDD.t4016 8.10567
R21711 VDD.n12508 VDD.t3794 8.10567
R21712 VDD.n8694 VDD.t4354 8.10567
R21713 VDD.n8694 VDD.t4166 8.10567
R21714 VDD.n8691 VDD.t4704 8.10567
R21715 VDD.n8691 VDD.t4482 8.10567
R21716 VDD.n8690 VDD.t1155 8.10567
R21717 VDD.n8690 VDD.t986 8.10567
R21718 VDD.n12512 VDD.t4722 8.10567
R21719 VDD.n12512 VDD.t4490 8.10567
R21720 VDD.n12511 VDD.t978 8.10567
R21721 VDD.n12511 VDD.t750 8.10567
R21722 VDD.n12508 VDD.t2635 8.10567
R21723 VDD.n12508 VDD.t2410 8.10567
R21724 VDD.n8608 VDD.t2684 8.10567
R21725 VDD.n8684 VDD.t4182 8.10567
R21726 VDD.n8609 VDD.t4048 8.10567
R21727 VDD.n8678 VDD.t3818 8.10567
R21728 VDD.n8605 VDD.t2789 8.10567
R21729 VDD.n8710 VDD.t4260 8.10567
R21730 VDD.n8606 VDD.t1633 8.10567
R21731 VDD.n8704 VDD.t1405 8.10567
R21732 VDD.n8602 VDD.t4148 8.10567
R21733 VDD.n8602 VDD.t1507 8.10567
R21734 VDD.n8599 VDD.t4470 8.10567
R21735 VDD.n8599 VDD.t1875 8.10567
R21736 VDD.n8598 VDD.t970 8.10567
R21737 VDD.n8598 VDD.t2599 8.10567
R21738 VDD.n12478 VDD.t4484 8.10567
R21739 VDD.n12478 VDD.t1892 8.10567
R21740 VDD.n12479 VDD.t727 8.10567
R21741 VDD.n12479 VDD.t2349 8.10567
R21742 VDD.n12483 VDD.t2387 8.10567
R21743 VDD.n12483 VDD.t3878 8.10567
R21744 VDD.n8602 VDD.t4440 8.10567
R21745 VDD.n8602 VDD.t4246 8.10567
R21746 VDD.n8599 VDD.t622 8.10567
R21747 VDD.n8599 VDD.t4548 8.10567
R21748 VDD.n8598 VDD.t1235 8.10567
R21749 VDD.n8598 VDD.t1049 8.10567
R21750 VDD.n12478 VDD.t654 8.10567
R21751 VDD.n12478 VDD.t4574 8.10567
R21752 VDD.n12479 VDD.t1038 8.10567
R21753 VDD.n12479 VDD.t830 8.10567
R21754 VDD.n12483 VDD.t2714 8.10567
R21755 VDD.n12483 VDD.t2498 8.10567
R21756 VDD.n12489 VDD.t905 8.10567
R21757 VDD.n105 VDD.t2524 8.10567
R21758 VDD.n12495 VDD.t3996 8.10567
R21759 VDD.n104 VDD.t3772 8.10567
R21760 VDD.n162 VDD.t2730 8.10567
R21761 VDD.n143 VDD.t4228 8.10567
R21762 VDD.n136 VDD.t4078 8.10567
R21763 VDD.n137 VDD.t3858 8.10567
R21764 VDD.n8732 VDD.t3630 8.10567
R21765 VDD.n8732 VDD.t1054 8.10567
R21766 VDD.n8729 VDD.t4008 8.10567
R21767 VDD.n8729 VDD.t1385 8.10567
R21768 VDD.n8728 VDD.t4586 8.10567
R21769 VDD.n8728 VDD.t2014 8.10567
R21770 VDD.n126 VDD.t4030 8.10567
R21771 VDD.n126 VDD.t1395 8.10567
R21772 VDD.n127 VDD.t4376 8.10567
R21773 VDD.n127 VDD.t1765 8.10567
R21774 VDD.n131 VDD.t1788 8.10567
R21775 VDD.n131 VDD.t3393 8.10567
R21776 VDD.n8732 VDD.t2078 8.10567
R21777 VDD.n8732 VDD.t1822 8.10567
R21778 VDD.n8729 VDD.t2496 8.10567
R21779 VDD.n8729 VDD.t2221 8.10567
R21780 VDD.n8728 VDD.t3096 8.10567
R21781 VDD.n8728 VDD.t2892 8.10567
R21782 VDD.n126 VDD.t2516 8.10567
R21783 VDD.n126 VDD.t2238 8.10567
R21784 VDD.n127 VDD.t2880 8.10567
R21785 VDD.n127 VDD.t2673 8.10567
R21786 VDD.n131 VDD.t4382 8.10567
R21787 VDD.n131 VDD.t4196 8.10567
R21788 VDD.n8594 VDD.t4454 8.10567
R21789 VDD.n8722 VDD.t1851 8.10567
R21790 VDD.n8595 VDD.t1709 8.10567
R21791 VDD.n8716 VDD.t1488 8.10567
R21792 VDD.n8592 VDD.t2346 8.10567
R21793 VDD.n8743 VDD.t3850 8.10567
R21794 VDD.n8593 VDD.t2384 8.10567
R21795 VDD.n8737 VDD.t2099 8.10567
R21796 VDD.n8589 VDD.t4218 8.10567
R21797 VDD.n8589 VDD.t1129 8.10567
R21798 VDD.n8586 VDD.t4524 8.10567
R21799 VDD.n8586 VDD.t1461 8.10567
R21800 VDD.n8585 VDD.t1022 8.10567
R21801 VDD.n8585 VDD.t2109 8.10567
R21802 VDD.n12456 VDD.t4532 8.10567
R21803 VDD.n12456 VDD.t1477 8.10567
R21804 VDD.n12455 VDD.t794 8.10567
R21805 VDD.n12455 VDD.t1860 8.10567
R21806 VDD.n12452 VDD.t2456 8.10567
R21807 VDD.n12452 VDD.t3486 8.10567
R21808 VDD.n8589 VDD.t2716 8.10567
R21809 VDD.n8589 VDD.t3826 8.10567
R21810 VDD.n8586 VDD.t3058 8.10567
R21811 VDD.n8586 VDD.t4194 8.10567
R21812 VDD.n8585 VDD.t3601 8.10567
R21813 VDD.n8585 VDD.t613 8.10567
R21814 VDD.n12456 VDD.t3076 8.10567
R21815 VDD.n12456 VDD.t4216 8.10567
R21816 VDD.n12455 VDD.t3385 8.10567
R21817 VDD.n12455 VDD.t4534 8.10567
R21818 VDD.n12452 VDD.t825 8.10567
R21819 VDD.n12452 VDD.t2004 8.10567
R21820 VDD.n669 VDD.t3126 8.10567
R21821 VDD.n669 VDD.t1671 8.10567
R21822 VDD.n11063 VDD.t2799 8.10567
R21823 VDD.n11063 VDD.t1312 8.10567
R21824 VDD.n661 VDD.t1101 8.10567
R21825 VDD.n661 VDD.t3882 8.10567
R21826 VDD.n11097 VDD.t2791 8.10567
R21827 VDD.n11097 VDD.t1295 8.10567
R21828 VDD.n651 VDD.t2393 8.10567
R21829 VDD.n651 VDD.t967 8.10567
R21830 VDD.n11119 VDD.t2043 8.10567
R21831 VDD.n11119 VDD.t3942 8.10567
R21832 VDD.n5717 VDD.t4222 8.10567
R21833 VDD.n5718 VDD.t1755 8.10567
R21834 VDD.n11033 VDD.t1243 8.10567
R21835 VDD.n1769 VDD.t3591 8.10567
R21836 VDD.n5714 VDD.t2613 8.10567
R21837 VDD.n5714 VDD.t2128 8.10567
R21838 VDD.n5711 VDD.t2186 8.10567
R21839 VDD.n5711 VDD.t1740 8.10567
R21840 VDD.n5710 VDD.t4702 8.10567
R21841 VDD.n5710 VDD.t4306 8.10567
R21842 VDD.n11011 VDD.t2170 8.10567
R21843 VDD.n11011 VDD.t1730 8.10567
R21844 VDD.n11012 VDD.t1748 8.10567
R21845 VDD.n11012 VDD.t1356 8.10567
R21846 VDD.n11016 VDD.t2868 8.10567
R21847 VDD.n11016 VDD.t2070 8.10567
R21848 VDD.n5714 VDD.t2490 8.10567
R21849 VDD.n5714 VDD.t4706 8.10567
R21850 VDD.n5711 VDD.t2068 8.10567
R21851 VDD.n5711 VDD.t4358 8.10567
R21852 VDD.n5710 VDD.t4560 8.10567
R21853 VDD.n5710 VDD.t2836 8.10567
R21854 VDD.n11011 VDD.t2048 8.10567
R21855 VDD.n11011 VDD.t4348 8.10567
R21856 VDD.n11012 VDD.t1643 8.10567
R21857 VDD.n11012 VDD.t3982 8.10567
R21858 VDD.n11016 VDD.t2364 8.10567
R21859 VDD.n11016 VDD.t1421 8.10567
R21860 VDD.n11022 VDD.t3693 8.10567
R21861 VDD.n1779 VDD.t2615 8.10567
R21862 VDD.n1773 VDD.t584 8.10567
R21863 VDD.n1775 VDD.t3946 8.10567
R21864 VDD.n1806 VDD.t4452 8.10567
R21865 VDD.n1820 VDD.t3316 8.10567
R21866 VDD.n1807 VDD.t1359 8.10567
R21867 VDD.n1814 VDD.t1555 8.10567
R21868 VDD.n5740 VDD.t4356 8.10567
R21869 VDD.n5740 VDD.t1559 8.10567
R21870 VDD.n5737 VDD.t4020 8.10567
R21871 VDD.n5737 VDD.t1202 8.10567
R21872 VDD.n5736 VDD.t2487 8.10567
R21873 VDD.n5736 VDD.t3778 8.10567
R21874 VDD.n1797 VDD.t4002 8.10567
R21875 VDD.n1797 VDD.t1193 8.10567
R21876 VDD.n1798 VDD.t3620 8.10567
R21877 VDD.n1798 VDD.t854 8.10567
R21878 VDD.n1802 VDD.t4034 8.10567
R21879 VDD.n1802 VDD.t2886 8.10567
R21880 VDD.n5740 VDD.t1847 8.10567
R21881 VDD.n5740 VDD.t4190 8.10567
R21882 VDD.n5737 VDD.t1481 8.10567
R21883 VDD.n5737 VDD.t3824 8.10567
R21884 VDD.n5736 VDD.t4056 8.10567
R21885 VDD.n5736 VDD.t2236 8.10567
R21886 VDD.n1797 VDD.t1473 8.10567
R21887 VDD.n1797 VDD.t3810 8.10567
R21888 VDD.n1798 VDD.t1114 8.10567
R21889 VDD.n1798 VDD.t3450 8.10567
R21890 VDD.n1802 VDD.t3114 8.10567
R21891 VDD.n1802 VDD.t2233 8.10567
R21892 VDD.n5706 VDD.t3648 8.10567
R21893 VDD.n5730 VDD.t1227 8.10567
R21894 VDD.n5707 VDD.t732 8.10567
R21895 VDD.n5724 VDD.t1617 8.10567
R21896 VDD.n5753 VDD.t1318 8.10567
R21897 VDD.n5751 VDD.t1662 8.10567
R21898 VDD.n5705 VDD.t2657 8.10567
R21899 VDD.n5745 VDD.t3490 8.10567
R21900 VDD.n5701 VDD.t3948 8.10567
R21901 VDD.n5701 VDD.t1140 8.10567
R21902 VDD.n5698 VDD.t3585 8.10567
R21903 VDD.n5698 VDD.t806 8.10567
R21904 VDD.n5697 VDD.t1969 8.10567
R21905 VDD.n5697 VDD.t3352 8.10567
R21906 VDD.n10990 VDD.t3566 8.10567
R21907 VDD.n10990 VDD.t791 8.10567
R21908 VDD.n10989 VDD.t3246 8.10567
R21909 VDD.n10989 VDD.t4530 8.10567
R21910 VDD.n10986 VDD.t919 8.10567
R21911 VDD.n10986 VDD.t3844 8.10567
R21912 VDD.n5701 VDD.t747 8.10567
R21913 VDD.n5701 VDD.t946 8.10567
R21914 VDD.n5698 VDD.t4508 8.10567
R21915 VDD.n5698 VDD.t4712 8.10567
R21916 VDD.n5697 VDD.t3012 8.10567
R21917 VDD.n5697 VDD.t3168 8.10567
R21918 VDD.n10990 VDD.t4496 8.10567
R21919 VDD.n10990 VDD.t4698 8.10567
R21920 VDD.n10989 VDD.t4162 8.10567
R21921 VDD.n10989 VDD.t4326 8.10567
R21922 VDD.n10986 VDD.t4606 8.10567
R21923 VDD.n10986 VDD.t3140 8.10567
R21924 VDD.n10977 VDD.t1503 8.10567
R21925 VDD.n10979 VDD.t1387 8.10567
R21926 VDD.n1796 VDD.t2692 8.10567
R21927 VDD.n1826 VDD.t2888 8.10567
R21928 VDD.n10967 VDD.t1138 8.10567
R21929 VDD.n1841 VDD.t1331 8.10567
R21930 VDD.n10973 VDD.t3628 8.10567
R21931 VDD.n1840 VDD.t2520 8.10567
R21932 VDD.n5795 VDD.t1598 8.10567
R21933 VDD.n5795 VDD.t3068 8.10567
R21934 VDD.n5792 VDD.t1237 8.10567
R21935 VDD.n5792 VDD.t2728 8.10567
R21936 VDD.n5791 VDD.t3804 8.10567
R21937 VDD.n5791 VDD.t1032 8.10567
R21938 VDD.n10956 VDD.t1229 8.10567
R21939 VDD.n10956 VDD.t2706 8.10567
R21940 VDD.n10957 VDD.t895 8.10567
R21941 VDD.n10957 VDD.t2282 8.10567
R21942 VDD.n10961 VDD.t2126 8.10567
R21943 VDD.n10961 VDD.t937 8.10567
R21944 VDD.n5795 VDD.t3306 8.10567
R21945 VDD.n5795 VDD.t4642 8.10567
R21946 VDD.n5792 VDD.t3008 8.10567
R21947 VDD.n5792 VDD.t4292 8.10567
R21948 VDD.n5791 VDD.t1284 8.10567
R21949 VDD.n5791 VDD.t2778 8.10567
R21950 VDD.n10956 VDD.t2992 8.10567
R21951 VDD.n10956 VDD.t4280 8.10567
R21952 VDD.n10957 VDD.t2619 8.10567
R21953 VDD.n10957 VDD.t3910 8.10567
R21954 VDD.n10961 VDD.t1144 8.10567
R21955 VDD.n10961 VDD.t4126 8.10567
R21956 VDD.n5693 VDD.t1363 8.10567
R21957 VDD.n5785 VDD.t2366 8.10567
R21958 VDD.n5694 VDD.t2143 8.10567
R21959 VDD.n5779 VDD.t3524 8.10567
R21960 VDD.n5691 VDD.t871 8.10567
R21961 VDD.n5806 VDD.t1728 8.10567
R21962 VDD.n5692 VDD.t3984 8.10567
R21963 VDD.n5800 VDD.t1177 8.10567
R21964 VDD.n5688 VDD.t1519 8.10567
R21965 VDD.n5688 VDD.t2542 8.10567
R21966 VDD.n5685 VDD.t1173 8.10567
R21967 VDD.n5685 VDD.t2107 8.10567
R21968 VDD.n5684 VDD.t3737 8.10567
R21969 VDD.n5684 VDD.t4628 8.10567
R21970 VDD.n1880 VDD.t1160 8.10567
R21971 VDD.n1880 VDD.t2095 8.10567
R21972 VDD.n1881 VDD.t803 8.10567
R21973 VDD.n1881 VDD.t1687 8.10567
R21974 VDD.n1885 VDD.t1439 8.10567
R21975 VDD.n1885 VDD.t1659 8.10567
R21976 VDD.n5688 VDD.t2816 8.10567
R21977 VDD.n5688 VDD.t4130 8.10567
R21978 VDD.n5685 VDD.t2458 8.10567
R21979 VDD.n5685 VDD.t3760 8.10567
R21980 VDD.n5684 VDD.t782 8.10567
R21981 VDD.n5684 VDD.t2156 8.10567
R21982 VDD.n1880 VDD.t2445 8.10567
R21983 VDD.n1880 VDD.t3743 8.10567
R21984 VDD.n1881 VDD.t1983 8.10567
R21985 VDD.n1881 VDD.t3375 8.10567
R21986 VDD.n1885 VDD.t1903 8.10567
R21987 VDD.n1885 VDD.t699 8.10567
R21988 VDD.n1862 VDD.t1901 8.10567
R21989 VDD.n1876 VDD.t2119 8.10567
R21990 VDD.n1863 VDD.t705 8.10567
R21991 VDD.n1870 VDD.t3654 8.10567
R21992 VDD.n10922 VDD.t3200 8.10567
R21993 VDD.n10924 VDD.t3354 8.10567
R21994 VDD.n1861 VDD.t1444 8.10567
R21995 VDD.n1891 VDD.t4402 8.10567
R21996 VDD.n5850 VDD.t4104 8.10567
R21997 VDD.n5850 VDD.t857 8.10567
R21998 VDD.n5847 VDD.t3729 8.10567
R21999 VDD.n5847 VDD.t4622 8.10567
R22000 VDD.n5846 VDD.t2121 8.10567
R22001 VDD.n5846 VDD.t3094 8.10567
R22002 VDD.n10935 VDD.t3717 8.10567
R22003 VDD.n10935 VDD.t4602 8.10567
R22004 VDD.n10934 VDD.t3340 8.10567
R22005 VDD.n10934 VDD.t4254 8.10567
R22006 VDD.n10931 VDD.t2178 8.10567
R22007 VDD.n10931 VDD.t2443 8.10567
R22008 VDD.n5850 VDD.t4538 8.10567
R22009 VDD.n5850 VDD.t1769 8.10567
R22010 VDD.n5847 VDD.t4234 8.10567
R22011 VDD.n5847 VDD.t1413 8.10567
R22012 VDD.n5846 VDD.t2681 8.10567
R22013 VDD.n5846 VDD.t3992 8.10567
R22014 VDD.n10935 VDD.t4224 8.10567
R22015 VDD.n10935 VDD.t1401 8.10567
R22016 VDD.n10934 VDD.t3830 8.10567
R22017 VDD.n10934 VDD.t1051 8.10567
R22018 VDD.n10931 VDD.t3202 8.10567
R22019 VDD.n10931 VDD.t1925 8.10567
R22020 VDD.n5820 VDD.t2775 8.10567
R22021 VDD.n5818 VDD.t3593 8.10567
R22022 VDD.n5681 VDD.t3458 8.10567
R22023 VDD.n5812 VDD.t646 8.10567
R22024 VDD.n5678 VDD.t2925 8.10567
R22025 VDD.n5861 VDD.t3750 8.10567
R22026 VDD.n5679 VDD.t4626 8.10567
R22027 VDD.n5855 VDD.t1842 8.10567
R22028 VDD.n5675 VDD.t2141 8.10567
R22029 VDD.n5675 VDD.t4444 8.10567
R22030 VDD.n5672 VDD.t1753 8.10567
R22031 VDD.n5672 VDD.t4118 8.10567
R22032 VDD.n5671 VDD.t4320 8.10567
R22033 VDD.n5671 VDD.t2571 8.10567
R22034 VDD.n10901 VDD.t1738 8.10567
R22035 VDD.n10901 VDD.t4098 8.10567
R22036 VDD.n10902 VDD.t1367 8.10567
R22037 VDD.n10902 VDD.t3703 8.10567
R22038 VDD.n10906 VDD.t3976 8.10567
R22039 VDD.n10906 VDD.t3182 8.10567
R22040 VDD.n5675 VDD.t1602 8.10567
R22041 VDD.n5675 VDD.t1946 8.10567
R22042 VDD.n5672 VDD.t1241 8.10567
R22043 VDD.n5672 VDD.t1582 8.10567
R22044 VDD.n5671 VDD.t3814 8.10567
R22045 VDD.n5671 VDD.t4160 8.10567
R22046 VDD.n10901 VDD.t1231 8.10567
R22047 VDD.n10901 VDD.t1557 8.10567
R22048 VDD.n10902 VDD.t907 8.10567
R22049 VDD.n10902 VDD.t1185 8.10567
R22050 VDD.n10906 VDD.t2358 8.10567
R22051 VDD.n10906 VDD.t2176 8.10567
R22052 VDD.n10912 VDD.t3369 8.10567
R22053 VDD.n1906 VDD.t3570 8.10567
R22054 VDD.n10918 VDD.t574 8.10567
R22055 VDD.n1905 VDD.t3568 8.10567
R22056 VDD.n5510 VDD.t4562 8.10567
R22057 VDD.n5524 VDD.t3399 8.10567
R22058 VDD.n5511 VDD.t2974 8.10567
R22059 VDD.n5518 VDD.t611 8.10567
R22060 VDD.n5897 VDD.t1578 8.10567
R22061 VDD.n5897 VDD.t3922 8.10567
R22062 VDD.n5894 VDD.t1225 8.10567
R22063 VDD.n5894 VDD.t3564 8.10567
R22064 VDD.n5893 VDD.t3790 8.10567
R22065 VDD.n5893 VDD.t1937 8.10567
R22066 VDD.n5494 VDD.t1200 8.10567
R22067 VDD.n5494 VDD.t3546 8.10567
R22068 VDD.n5495 VDD.t877 8.10567
R22069 VDD.n5495 VDD.t3224 8.10567
R22070 VDD.n5499 VDD.t4710 8.10567
R22071 VDD.n5499 VDD.t3884 8.10567
R22072 VDD.n5897 VDD.t3940 8.10567
R22073 VDD.n5897 VDD.t3796 8.10567
R22074 VDD.n5894 VDD.t3579 8.10567
R22075 VDD.n5894 VDD.t3462 8.10567
R22076 VDD.n5893 VDD.t1958 8.10567
R22077 VDD.n5893 VDD.t1800 8.10567
R22078 VDD.n5494 VDD.t3556 8.10567
R22079 VDD.n5494 VDD.t3442 8.10567
R22080 VDD.n5495 VDD.t3240 8.10567
R22081 VDD.n5495 VDD.t3112 8.10567
R22082 VDD.n5499 VDD.t2115 8.10567
R22083 VDD.n5499 VDD.t3403 8.10567
R22084 VDD.n5667 VDD.t4676 8.10567
R22085 VDD.n5873 VDD.t1888 8.10567
R22086 VDD.n5668 VDD.t935 8.10567
R22087 VDD.n5867 VDD.t3697 8.10567
R22088 VDD.n5545 VDD.t2818 8.10567
R22089 VDD.n5543 VDD.t1340 8.10567
R22090 VDD.n5663 VDD.t868 8.10567
R22091 VDD.n5542 VDD.t3214 8.10567
R22092 VDD.n5633 VDD.t1030 8.10567
R22093 VDD.n5633 VDD.t2850 8.10567
R22094 VDD.n5630 VDD.t662 8.10567
R22095 VDD.n5630 VDD.t2494 8.10567
R22096 VDD.n5629 VDD.t3274 8.10567
R22097 VDD.n5629 VDD.t800 8.10567
R22098 VDD.n10880 VDD.t641 8.10567
R22099 VDD.n10880 VDD.t2485 8.10567
R22100 VDD.n10879 VDD.t4412 8.10567
R22101 VDD.n10879 VDD.t2025 8.10567
R22102 VDD.n10876 VDD.t4332 8.10567
R22103 VDD.n10876 VDD.t3216 8.10567
R22104 VDD.n5633 VDD.t1975 8.10567
R22105 VDD.n5633 VDD.t3294 8.10567
R22106 VDD.n5630 VDD.t1606 8.10567
R22107 VDD.n5630 VDD.t2988 8.10567
R22108 VDD.n5629 VDD.t4186 8.10567
R22109 VDD.n5629 VDD.t1264 8.10567
R22110 VDD.n10880 VDD.t1590 8.10567
R22111 VDD.n10880 VDD.t2966 8.10567
R22112 VDD.n10879 VDD.t1211 8.10567
R22113 VDD.n10879 VDD.t2597 8.10567
R22114 VDD.n10876 VDD.t3912 8.10567
R22115 VDD.n10876 VDD.t4168 8.10567
R22116 VDD.n10867 VDD.t2263 8.10567
R22117 VDD.n10869 VDD.t4164 8.10567
R22118 VDD.n5506 VDD.t2261 8.10567
R22119 VDD.n5504 VDD.t1380 8.10567
R22120 VDD.n10857 VDD.t2544 8.10567
R22121 VDD.n1933 VDD.t667 8.10567
R22122 VDD.n10863 VDD.t3014 8.10567
R22123 VDD.n1932 VDD.t2097 8.10567
R22124 VDD.n5612 VDD.t4624 8.10567
R22125 VDD.n5612 VDD.t828 8.10567
R22126 VDD.n5609 VDD.t4288 8.10567
R22127 VDD.n5609 VDD.t4600 8.10567
R22128 VDD.n5608 VDD.t2759 8.10567
R22129 VDD.n5608 VDD.t3080 8.10567
R22130 VDD.n10846 VDD.t4272 8.10567
R22131 VDD.n10846 VDD.t4576 8.10567
R22132 VDD.n10847 VDD.t3896 8.10567
R22133 VDD.n10847 VDD.t4240 8.10567
R22134 VDD.n10851 VDD.t957 8.10567
R22135 VDD.n10851 VDD.t815 8.10567
R22136 VDD.n5612 VDD.t2154 8.10567
R22137 VDD.n5612 VDD.t4448 8.10567
R22138 VDD.n5609 VDD.t1759 8.10567
R22139 VDD.n5609 VDD.t4122 8.10567
R22140 VDD.n5608 VDD.t4324 8.10567
R22141 VDD.n5608 VDD.t2574 8.10567
R22142 VDD.n10846 VDD.t1744 8.10567
R22143 VDD.n10846 VDD.t4100 8.10567
R22144 VDD.n10847 VDD.t1375 8.10567
R22145 VDD.n10847 VDD.t3709 8.10567
R22146 VDD.n10851 VDD.t4144 8.10567
R22147 VDD.n10851 VDD.t3320 8.10567
R22148 VDD.n5617 VDD.t2984 8.10567
R22149 VDD.n5548 VDD.t3906 8.10567
R22150 VDD.n5623 VDD.t3391 8.10567
R22151 VDD.n5547 VDD.t1514 8.10567
R22152 VDD.n5596 VDD.t4724 8.10567
R22153 VDD.n5550 VDD.t3365 8.10567
R22154 VDD.n5602 VDD.t2922 8.10567
R22155 VDD.n5549 VDD.t3747 8.10567
R22156 VDD.n5591 VDD.t2404 8.10567
R22157 VDD.n5591 VDD.t2749 8.10567
R22158 VDD.n5588 VDD.t1971 8.10567
R22159 VDD.n5588 VDD.t2376 8.10567
R22160 VDD.n5587 VDD.t4488 8.10567
R22161 VDD.n5587 VDD.t676 8.10567
R22162 VDD.n1972 VDD.t1944 8.10567
R22163 VDD.n1972 VDD.t2356 8.10567
R22164 VDD.n1973 VDD.t1550 8.10567
R22165 VDD.n1973 VDD.t1897 8.10567
R22166 VDD.n1977 VDD.t2182 8.10567
R22167 VDD.n1977 VDD.t2052 8.10567
R22168 VDD.n5591 VDD.t3988 8.10567
R22169 VDD.n5591 VDD.t2152 8.10567
R22170 VDD.n5588 VDD.t3624 8.10567
R22171 VDD.n5588 VDD.t1757 8.10567
R22172 VDD.n5587 VDD.t2012 8.10567
R22173 VDD.n5587 VDD.t4322 8.10567
R22174 VDD.n1972 VDD.t3609 8.10567
R22175 VDD.n1972 VDD.t1742 8.10567
R22176 VDD.n1973 VDD.t3284 8.10567
R22177 VDD.n1973 VDD.t1372 8.10567
R22178 VDD.n1977 VDD.t1182 8.10567
R22179 VDD.n1977 VDD.t4494 8.10567
R22180 VDD.n1954 VDD.t3678 8.10567
R22181 VDD.n1968 VDD.t1407 8.10567
R22182 VDD.n1955 VDD.t3676 8.10567
R22183 VDD.n1962 VDD.t3888 8.10567
R22184 VDD.n10809 VDD.t4436 8.10567
R22185 VDD.n10811 VDD.t3290 8.10567
R22186 VDD.n1953 VDD.t4432 8.10567
R22187 VDD.n1983 VDD.t4634 8.10567
R22188 VDD.n2116 VDD.t2569 8.10567
R22189 VDD.n2116 VDD.t3864 8.10567
R22190 VDD.n2113 VDD.t2137 8.10567
R22191 VDD.n2113 VDD.t3516 8.10567
R22192 VDD.n2112 VDD.t4666 8.10567
R22193 VDD.n2112 VDD.t1877 8.10567
R22194 VDD.n10825 VDD.t2117 8.10567
R22195 VDD.n10825 VDD.t3504 8.10567
R22196 VDD.n10824 VDD.t1715 8.10567
R22197 VDD.n10824 VDD.t3174 8.10567
R22198 VDD.n10821 VDD.t2471 8.10567
R22199 VDD.n10821 VDD.t1166 8.10567
R22200 VDD.n2116 VDD.t3464 8.10567
R22201 VDD.n2116 VDD.t651 8.10567
R22202 VDD.n2113 VDD.t3154 8.10567
R22203 VDD.n2113 VDD.t4456 8.10567
R22204 VDD.n2112 VDD.t1441 8.10567
R22205 VDD.n2112 VDD.t2934 8.10567
R22206 VDD.n10825 VDD.t3132 8.10567
R22207 VDD.n10825 VDD.t4430 8.10567
R22208 VDD.n10824 VDD.t2793 8.10567
R22209 VDD.n10824 VDD.t4074 8.10567
R22210 VDD.n10821 VDD.t1956 8.10567
R22211 VDD.n10821 VDD.t772 8.10567
R22212 VDD.n5554 VDD.t4210 8.10567
R22213 VDD.n5552 VDD.t1393 8.10567
R22214 VDD.n5581 VDD.t2380 8.10567
R22215 VDD.n5551 VDD.t3266 8.10567
R22216 VDD.n2102 VDD.t4106 8.10567
R22217 VDD.n8106 VDD.t864 8.10567
R22218 VDD.n2103 VDD.t674 8.10567
R22219 VDD.n8100 VDD.t2084 8.10567
R22220 VDD.n2099 VDD.t1931 8.10567
R22221 VDD.n2099 VDD.t3334 8.10567
R22222 VDD.n2096 VDD.t1565 8.10567
R22223 VDD.n2096 VDD.t3042 8.10567
R22224 VDD.n2095 VDD.t4152 8.10567
R22225 VDD.n2095 VDD.t1324 8.10567
R22226 VDD.n10788 VDD.t1544 8.10567
R22227 VDD.n10788 VDD.t3028 8.10567
R22228 VDD.n10789 VDD.t1179 8.10567
R22229 VDD.n10789 VDD.t2663 8.10567
R22230 VDD.n10793 VDD.t3204 8.10567
R22231 VDD.n10793 VDD.t1927 8.10567
R22232 VDD.n2099 VDD.t1795 8.10567
R22233 VDD.n2099 VDD.t3256 8.10567
R22234 VDD.n2096 VDD.t1435 8.10567
R22235 VDD.n2096 VDD.t2928 8.10567
R22236 VDD.n2095 VDD.t4028 8.10567
R22237 VDD.n2095 VDD.t1208 8.10567
R22238 VDD.n10788 VDD.t1424 8.10567
R22239 VDD.n10788 VDD.t2908 8.10567
R22240 VDD.n10789 VDD.t1083 8.10567
R22241 VDD.n10789 VDD.t2540 8.10567
R22242 VDD.n10793 VDD.t2743 8.10567
R22243 VDD.n10793 VDD.t1415 8.10567
R22244 VDD.n10799 VDD.t2741 8.10567
R22245 VDD.n2006 VDD.t2938 8.10567
R22246 VDD.n10805 VDD.t1003 8.10567
R22247 VDD.n2005 VDD.t3938 8.10567
R22248 VDD.n2036 VDD.t3423 8.10567
R22249 VDD.n2050 VDD.t3613 8.10567
R22250 VDD.n2037 VDD.t1712 8.10567
R22251 VDD.n2044 VDD.t4682 8.10567
R22252 VDD.n8128 VDD.t4258 8.10567
R22253 VDD.n8128 VDD.t1015 8.10567
R22254 VDD.n8125 VDD.t3902 8.10567
R22255 VDD.n8125 VDD.t636 8.10567
R22256 VDD.n8124 VDD.t2351 8.10567
R22257 VDD.n8124 VDD.t3250 8.10567
R22258 VDD.n2027 VDD.t3880 8.10567
R22259 VDD.n2027 VDD.t601 8.10567
R22260 VDD.n2028 VDD.t3512 8.10567
R22261 VDD.n2028 VDD.t4394 8.10567
R22262 VDD.n2032 VDD.t3038 8.10567
R22263 VDD.n2032 VDD.t3222 8.10567
R22264 VDD.n8128 VDD.t1262 8.10567
R22265 VDD.n8128 VDD.t2753 8.10567
R22266 VDD.n8125 VDD.t955 8.10567
R22267 VDD.n8125 VDD.t2382 8.10567
R22268 VDD.n8124 VDD.t3488 8.10567
R22269 VDD.n8124 VDD.t679 8.10567
R22270 VDD.n2027 VDD.t932 8.10567
R22271 VDD.n2027 VDD.t2362 8.10567
R22272 VDD.n2028 VDD.t4684 8.10567
R22273 VDD.n2028 VDD.t1899 8.10567
R22274 VDD.n2032 VDD.t3426 8.10567
R22275 VDD.n2032 VDD.t2229 8.10567
R22276 VDD.n2091 VDD.t3550 8.10567
R22277 VDD.n8118 VDD.t4450 8.10567
R22278 VDD.n2092 VDD.t4298 8.10567
R22279 VDD.n8112 VDD.t1496 8.10567
R22280 VDD.n8141 VDD.t1206 8.10567
R22281 VDD.n8139 VDD.t2150 8.10567
R22282 VDD.n2090 VDD.t1981 8.10567
R22283 VDD.n8133 VDD.t3367 8.10567
R22284 VDD.n8173 VDD.t757 8.10567
R22285 VDD.n8173 VDD.t2124 8.10567
R22286 VDD.n8188 VDD.t4518 8.10567
R22287 VDD.n8188 VDD.t1734 8.10567
R22288 VDD.n2078 VDD.t3020 8.10567
R22289 VDD.n2078 VDD.t4304 8.10567
R22290 VDD.n8222 VDD.t4504 8.10567
R22291 VDD.n8222 VDD.t1720 8.10567
R22292 VDD.n8229 VDD.t4174 8.10567
R22293 VDD.n8229 VDD.t1351 8.10567
R22294 VDD.n2064 VDD.t4184 8.10567
R22295 VDD.n2064 VDD.t3036 8.10567
R22296 VDD.n10768 VDD.t4616 8.10567
R22297 VDD.n2060 VDD.t672 8.10567
R22298 VDD.n2026 VDD.t3040 8.10567
R22299 VDD.n2056 VDD.t1732 8.10567
R22300 VDD.n2248 VDD.t3954 8.10567
R22301 VDD.n2250 VDD.t3587 8.10567
R22302 VDD.n7780 VDD.t1081 8.10567
R22303 VDD.n2272 VDD.t1093 8.10567
R22304 VDD.n7719 VDD.t2828 8.10567
R22305 VDD.n2282 VDD.t2454 8.10567
R22306 VDD.n2292 VDD.t2712 8.10567
R22307 VDD.n7825 VDD.t2054 8.10567
R22308 VDD.n7824 VDD.t1664 8.10567
R22309 VDD.n2240 VDD.t2332 8.10567
R22310 VDD.n7097 VDD.t3108 8.10567
R22311 VDD.n7093 VDD.t3964 8.10567
R22312 VDD.n7102 VDD.t1149 8.10567
R22313 VDD.n7090 VDD.t3970 8.10567
R22314 VDD.n7089 VDD.t3046 8.10567
R22315 VDD.n7109 VDD.t4700 8.10567
R22316 VDD.n2329 VDD.t1921 8.10567
R22317 VDD.n7115 VDD.t2427 8.10567
R22318 VDD.n2327 VDD.t3725 8.10567
R22319 VDD.n7120 VDD.t974 8.10567
R22320 VDD.n2324 VDD.t2249 8.10567
R22321 VDD.n2240 VDD.t4336 8.10567
R22322 VDD.n7097 VDD.t972 8.10567
R22323 VDD.n7093 VDD.t1832 8.10567
R22324 VDD.n7102 VDD.t3282 8.10567
R22325 VDD.n7090 VDD.t1840 8.10567
R22326 VDD.n7089 VDD.t903 8.10567
R22327 VDD.n7109 VDD.t2702 8.10567
R22328 VDD.n2329 VDD.t4004 8.10567
R22329 VDD.n7115 VDD.t4392 8.10567
R22330 VDD.n2327 VDD.t1615 8.10567
R22331 VDD.n7120 VDD.t3082 8.10567
R22332 VDD.n2324 VDD.t4284 8.10567
R22333 VDD.n2400 VDD.t2874 8.10567
R22334 VDD.n2398 VDD.t4426 8.10567
R22335 VDD.n2397 VDD.t4092 8.10567
R22336 VDD.n7129 VDD.t994 8.10567
R22337 VDD.n7128 VDD.t4742 8.10567
R22338 VDD.n7126 VDD.t2295 8.10567
R22339 VDD.n2400 VDD.t2528 8.10567
R22340 VDD.n2398 VDD.t4114 8.10567
R22341 VDD.n2397 VDD.t3733 8.10567
R22342 VDD.n7129 VDD.t586 8.10567
R22343 VDD.n7128 VDD.t4396 8.10567
R22344 VDD.n7126 VDD.t1890 8.10567
R22345 VDD.n2343 VDD.t4310 8.10567
R22346 VDD.n2345 VDD.t2018 8.10567
R22347 VDD.n2346 VDD.t1641 8.10567
R22348 VDD.n7045 VDD.t3930 8.10567
R22349 VDD.n7046 VDD.t3562 8.10567
R22350 VDD.n2343 VDD.t3980 8.10567
R22351 VDD.n2345 VDD.t1657 8.10567
R22352 VDD.n2346 VDD.t1286 8.10567
R22353 VDD.n7045 VDD.t3577 8.10567
R22354 VDD.n7046 VDD.t3268 8.10567
R22355 VDD.n7071 VDD.t1815 8.10567
R22356 VDD.n7069 VDD.t2832 8.10567
R22357 VDD.n7076 VDD.t4142 8.10567
R22358 VDD.n7066 VDD.t2840 8.10567
R22359 VDD.n2335 VDD.t1736 8.10567
R22360 VDD.n7083 VDD.t3520 8.10567
R22361 VDD.n7063 VDD.t734 8.10567
R22362 VDD.n2336 VDD.t1134 8.10567
R22363 VDD.n2337 VDD.t2617 8.10567
R22364 VDD.n2338 VDD.t3908 8.10567
R22365 VDD.n2339 VDD.t1024 8.10567
R22366 VDD.n2340 VDD.t1063 8.10567
R22367 VDD.n6655 VDD.t697 8.10567
R22368 VDD.n6658 VDD.t1437 8.10567
R22369 VDD.n6653 VDD.t2930 8.10567
R22370 VDD.n6663 VDD.t3756 8.10567
R22371 VDD.n6650 VDD.t1316 8.10567
R22372 VDD.n6649 VDD.t833 8.10567
R22373 VDD.n6648 VDD.t3192 8.10567
R22374 VDD.n6647 VDD.t4492 8.10567
R22375 VDD.n6676 VDD.t4012 8.10567
R22376 VDD.n6645 VDD.t1112 8.10567
R22377 VDD.n6681 VDD.t2577 8.10567
R22378 VDD.n6642 VDD.t3415 8.10567
R22379 VDD.n7071 VDD.t1834 8.10567
R22380 VDD.n7069 VDD.t2848 8.10567
R22381 VDD.n7076 VDD.t4158 8.10567
R22382 VDD.n7066 VDD.t2854 8.10567
R22383 VDD.n2335 VDD.t1751 8.10567
R22384 VDD.n7083 VDD.t3532 8.10567
R22385 VDD.n7063 VDD.t760 8.10567
R22386 VDD.n2336 VDD.t1147 8.10567
R22387 VDD.n2337 VDD.t2633 8.10567
R22388 VDD.n2338 VDD.t3926 8.10567
R22389 VDD.n2339 VDD.t1036 8.10567
R22390 VDD.n2340 VDD.t1073 8.10567
R22391 VDD.n6655 VDD.t718 8.10567
R22392 VDD.n6658 VDD.t1469 8.10567
R22393 VDD.n6653 VDD.t2958 8.10567
R22394 VDD.n6663 VDD.t3776 8.10567
R22395 VDD.n6650 VDD.t1329 8.10567
R22396 VDD.n6649 VDD.t860 8.10567
R22397 VDD.n6648 VDD.t3212 8.10567
R22398 VDD.n6647 VDD.t4506 8.10567
R22399 VDD.n6676 VDD.t4026 8.10567
R22400 VDD.n6645 VDD.t1123 8.10567
R22401 VDD.n6681 VDD.t2595 8.10567
R22402 VDD.n6642 VDD.t3430 8.10567
R22403 VDD.n6711 VDD.t2872 8.10567
R22404 VDD.n6709 VDD.t4424 8.10567
R22405 VDD.n6708 VDD.t4090 8.10567
R22406 VDD.n6704 VDD.t992 8.10567
R22407 VDD.n6703 VDD.t4740 8.10567
R22408 VDD.n6701 VDD.t2293 8.10567
R22409 VDD.n6711 VDD.t707 8.10567
R22410 VDD.n6709 VDD.t2447 8.10567
R22411 VDD.n6708 VDD.t2000 8.10567
R22412 VDD.n6704 VDD.t3110 8.10567
R22413 VDD.n6703 VDD.t2781 8.10567
R22414 VDD.n6701 VDD.t4330 8.10567
R22415 VDD.n6697 VDD.t4308 8.10567
R22416 VDD.n6695 VDD.t2016 8.10567
R22417 VDD.n6694 VDD.t1639 8.10567
R22418 VDD.n6690 VDD.t3928 8.10567
R22419 VDD.n6689 VDD.t3560 8.10567
R22420 VDD.n6687 VDD.t1061 8.10567
R22421 VDD.n6697 VDD.t2259 8.10567
R22422 VDD.n6695 VDD.t4112 8.10567
R22423 VDD.n6694 VDD.t3731 8.10567
R22424 VDD.n6690 VDD.t1817 8.10567
R22425 VDD.n6689 VDD.t1451 8.10567
R22426 VDD.n6687 VDD.t3188 8.10567
R22427 VDD.n6640 VDD.t1075 8.10567
R22428 VDD.n6638 VDD.t2807 8.10567
R22429 VDD.n6637 VDD.t2437 8.10567
R22430 VDD.n5434 VDD.t2690 8.10567
R22431 VDD.n5435 VDD.t2276 8.10567
R22432 VDD.n5437 VDD.t1954 8.10567
R22433 VDD.n6640 VDD.t3206 8.10567
R22434 VDD.n6638 VDD.t616 8.10567
R22435 VDD.n6637 VDD.t4410 8.10567
R22436 VDD.n5434 VDD.t4678 8.10567
R22437 VDD.n5435 VDD.t4316 8.10567
R22438 VDD.n5437 VDD.t4050 8.10567
R22439 VDD.n5442 VDD.t888 8.10567
R22440 VDD.n5440 VDD.t2605 8.10567
R22441 VDD.n5439 VDD.t2168 8.10567
R22442 VDD.n6629 VDD.t2219 8.10567
R22443 VDD.n6628 VDD.t1807 8.10567
R22444 VDD.n6626 VDD.t3685 8.10567
R22445 VDD.n5442 VDD.t3022 8.10567
R22446 VDD.n5440 VDD.t4558 8.10567
R22447 VDD.n5439 VDD.t4242 8.10567
R22448 VDD.n6629 VDD.t4274 8.10567
R22449 VDD.n6628 VDD.t3920 8.10567
R22450 VDD.n6626 VDD.t1594 8.10567
R22451 VDD.n2374 VDD.t3270 8.10567
R22452 VDD.n2373 VDD.t4554 8.10567
R22453 VDD.n7030 VDD.t1314 8.10567
R22454 VDD.n2372 VDD.t3150 8.10567
R22455 VDD.n2371 VDD.t2651 8.10567
R22456 VDD.n7037 VDD.t725 8.10567
R22457 VDD.n6716 VDD.t2105 8.10567
R22458 VDD.n6715 VDD.t1553 8.10567
R22459 VDD.n6722 VDD.t2946 8.10567
R22460 VDD.n2407 VDD.t4244 8.10567
R22461 VDD.n2406 VDD.t1007 8.10567
R22462 VDD.n2385 VDD.t3589 8.10567
R22463 VDD.n6872 VDD.t4474 8.10567
R22464 VDD.n2391 VDD.t1689 8.10567
R22465 VDD.n6867 VDD.t4478 8.10567
R22466 VDD.n2392 VDD.t3514 8.10567
R22467 VDD.n6862 VDD.t1095 8.10567
R22468 VDD.n2393 VDD.t2556 8.10567
R22469 VDD.n2394 VDD.t2976 8.10567
R22470 VDD.n6854 VDD.t4268 8.10567
R22471 VDD.n2395 VDD.t1463 8.10567
R22472 VDD.n2404 VDD.t2844 8.10567
R22473 VDD.n5236 VDD.t2763 8.10567
R22474 VDD.n5234 VDD.t4058 8.10567
R22475 VDD.n5241 VDD.t810 8.10567
R22476 VDD.n5231 VDD.t2637 8.10567
R22477 VDD.n5230 VDD.t2041 8.10567
R22478 VDD.n5248 VDD.t4340 8.10567
R22479 VDD.n5227 VDD.t1533 8.10567
R22480 VDD.n5254 VDD.t1047 8.10567
R22481 VDD.n5225 VDD.t2391 8.10567
R22482 VDD.n5259 VDD.t3691 8.10567
R22483 VDD.n5222 VDD.t4572 8.10567
R22484 VDD.n5236 VDD.t4726 8.10567
R22485 VDD.n5234 VDD.t1948 8.10567
R22486 VDD.n5241 VDD.t2956 8.10567
R22487 VDD.n5231 VDD.t4578 8.10567
R22488 VDD.n5230 VDD.t4102 8.10567
R22489 VDD.n5248 VDD.t2280 8.10567
R22490 VDD.n5227 VDD.t3622 8.10567
R22491 VDD.n5254 VDD.t3162 8.10567
R22492 VDD.n5225 VDD.t4364 8.10567
R22493 VDD.n5259 VDD.t1576 8.10567
R22494 VDD.n5222 VDD.t2593 8.10567
R22495 VDD.n5474 VDD.t4418 8.10567
R22496 VDD.n5475 VDD.t569 8.10567
R22497 VDD.n5476 VDD.t1987 8.10567
R22498 VDD.n5477 VDD.t4300 8.10567
R22499 VDD.n5478 VDD.t3788 8.10567
R22500 VDD.n5479 VDD.t1935 8.10567
R22501 VDD.n5480 VDD.t2336 8.10567
R22502 VDD.n5482 VDD.t3230 8.10567
R22503 VDD.n5483 VDD.t4088 8.10567
R22504 VDD.n5484 VDD.t1274 8.10567
R22505 VDD.n5485 VDD.t4096 8.10567
R22506 VDD.n5486 VDD.t4372 8.10567
R22507 VDD.n5474 VDD.t3338 8.10567
R22508 VDD.n5475 VDD.t3660 8.10567
R22509 VDD.n5476 VDD.t917 8.10567
R22510 VDD.n5477 VDD.t3264 8.10567
R22511 VDD.n5478 VDD.t2787 8.10567
R22512 VDD.n5479 VDD.t875 8.10567
R22513 VDD.n5480 VDD.t1169 8.10567
R22514 VDD.n5482 VDD.t2088 8.10567
R22515 VDD.n5483 VDD.t3052 8.10567
R22516 VDD.n5484 VDD.t4350 8.10567
R22517 VDD.n5485 VDD.t3056 8.10567
R22518 VDD.n5486 VDD.t3310 8.10567
R22519 VDD.n5446 VDD.t631 8.10567
R22520 VDD.n5391 VDD.t2039 8.10567
R22521 VDD.n5451 VDD.t3018 8.10567
R22522 VDD.n5388 VDD.t4668 8.10567
R22523 VDD.n5387 VDD.t4176 8.10567
R22524 VDD.n5458 VDD.t2389 8.10567
R22525 VDD.n5384 VDD.t3689 8.10567
R22526 VDD.n5464 VDD.t4542 8.10567
R22527 VDD.n5382 VDD.t4438 8.10567
R22528 VDD.n5469 VDD.t1652 8.10567
R22529 VDD.n5379 VDD.t3994 8.10567
R22530 VDD.n5446 VDD.t3701 8.10567
R22531 VDD.n5391 VDD.t951 8.10567
R22532 VDD.n5451 VDD.t1811 8.10567
R22533 VDD.n5388 VDD.t3583 8.10567
R22534 VDD.n5387 VDD.t3122 8.10567
R22535 VDD.n5458 VDD.t1195 8.10567
R22536 VDD.n5384 VDD.t2679 8.10567
R22537 VDD.n5464 VDD.t3500 8.10567
R22538 VDD.n5382 VDD.t3359 8.10567
R22539 VDD.n5469 VDD.t4714 8.10567
R22540 VDD.n5379 VDD.t2972 8.10567
R22541 VDD.n6264 VDD.t2481 8.10567
R22542 VDD.n6263 VDD.t2050 8.10567
R22543 VDD.n6366 VDD.t2344 8.10567
R22544 VDD.n6365 VDD.t1910 8.10567
R22545 VDD.n6363 VDD.t1623 8.10567
R22546 VDD.n6264 VDD.t3389 8.10567
R22547 VDD.n6263 VDD.t3090 8.10567
R22548 VDD.n6366 VDD.t3304 8.10567
R22549 VDD.n6365 VDD.t3002 8.10567
R22550 VDD.n6363 VDD.t2708 8.10567
R22551 VDD.n5937 VDD.t4690 8.10567
R22552 VDD.n5939 VDD.t2215 8.10567
R22553 VDD.n5940 VDD.t1803 8.10567
R22554 VDD.n5945 VDD.t1856 8.10567
R22555 VDD.n5946 VDD.t1486 8.10567
R22556 VDD.n5948 VDD.t3381 8.10567
R22557 VDD.n5937 VDD.t1501 8.10567
R22558 VDD.n5939 VDD.t3238 8.10567
R22559 VDD.n5940 VDD.t2898 8.10567
R22560 VDD.n5945 VDD.t2952 8.10567
R22561 VDD.n5946 VDD.t2585 8.10567
R22562 VDD.n5948 VDD.t4352 8.10567
R22563 VDD.n5271 VDD.t2460 8.10567
R22564 VDD.n6590 VDD.t3758 8.10567
R22565 VDD.n5272 VDD.t4648 8.10567
R22566 VDD.n6585 VDD.t2284 8.10567
R22567 VDD.n5273 VDD.t1701 8.10567
R22568 VDD.n6580 VDD.t4052 8.10567
R22569 VDD.n5924 VDD.t1245 8.10567
R22570 VDD.n5928 VDD.t2174 8.10567
R22571 VDD.n5923 VDD.t2029 8.10567
R22572 VDD.n5933 VDD.t3413 8.10567
R22573 VDD.n5922 VDD.t1529 8.10567
R22574 VDD.n6234 VDD.t3900 8.10567
R22575 VDD.n6232 VDD.t1117 8.10567
R22576 VDD.n6239 VDD.t2037 8.10567
R22577 VDD.n6229 VDD.t3770 8.10567
R22578 VDD.n6228 VDD.t3292 8.10567
R22579 VDD.n6246 VDD.t1391 8.10567
R22580 VDD.n6225 VDD.t2866 8.10567
R22581 VDD.n6252 VDD.t3664 8.10567
R22582 VDD.n6223 VDD.t3540 8.10567
R22583 VDD.n6257 VDD.t776 8.10567
R22584 VDD.n6220 VDD.t3142 8.10567
R22585 VDD.n6219 VDD.t736 8.10567
R22586 VDD.n6215 VDD.t1691 8.10567
R22587 VDD.n6270 VDD.t3534 8.10567
R22588 VDD.n6213 VDD.t3862 8.10567
R22589 VDD.n6275 VDD.t1086 8.10567
R22590 VDD.n6210 VDD.t3411 8.10567
R22591 VDD.n6209 VDD.t2964 8.10567
R22592 VDD.n6282 VDD.t1040 8.10567
R22593 VDD.n6206 VDD.t1349 8.10567
R22594 VDD.n6288 VDD.t2311 8.10567
R22595 VDD.n6204 VDD.t3228 8.10567
R22596 VDD.n6293 VDD.t4520 8.10567
R22597 VDD.n6201 VDD.t3234 8.10567
R22598 VDD.n6200 VDD.t3492 8.10567
R22599 VDD.n6234 VDD.t3918 8.10567
R22600 VDD.n6232 VDD.t1127 8.10567
R22601 VDD.n6239 VDD.t2058 8.10567
R22602 VDD.n6229 VDD.t3786 8.10567
R22603 VDD.n6228 VDD.t3300 8.10567
R22604 VDD.n6246 VDD.t1403 8.10567
R22605 VDD.n6225 VDD.t2878 8.10567
R22606 VDD.n6252 VDD.t3683 8.10567
R22607 VDD.n6223 VDD.t3552 8.10567
R22608 VDD.n6257 VDD.t787 8.10567
R22609 VDD.n6220 VDD.t3156 8.10567
R22610 VDD.n6219 VDD.t762 8.10567
R22611 VDD.n6215 VDD.t1707 8.10567
R22612 VDD.n6270 VDD.t3544 8.10567
R22613 VDD.n6213 VDD.t3876 8.10567
R22614 VDD.n6275 VDD.t1104 8.10567
R22615 VDD.n6210 VDD.t3432 8.10567
R22616 VDD.n6209 VDD.t2980 8.10567
R22617 VDD.n6282 VDD.t1065 8.10567
R22618 VDD.n6206 VDD.t1365 8.10567
R22619 VDD.n6288 VDD.t2334 8.10567
R22620 VDD.n6204 VDD.t3242 8.10567
R22621 VDD.n6293 VDD.t4526 8.10567
R22622 VDD.n6201 VDD.t3248 8.10567
R22623 VDD.n6200 VDD.t3502 8.10567
R22624 VDD.n6302 VDD.t1009 8.10567
R22625 VDD.n6303 VDD.t589 8.10567
R22626 VDD.n6307 VDD.t898 8.10567
R22627 VDD.n6306 VDD.t4652 8.10567
R22628 VDD.n5985 VDD.t789 8.10567
R22629 VDD.n5986 VDD.t4536 8.10567
R22630 VDD.n6315 VDD.t4594 8.10567
R22631 VDD.n6316 VDD.t4262 8.10567
R22632 VDD.n6318 VDD.t1950 8.10567
R22633 VDD.n5952 VDD.t2010 8.10567
R22634 VDD.n5921 VDD.t2418 8.10567
R22635 VDD.n5957 VDD.t3721 8.10567
R22636 VDD.n5920 VDD.t1864 8.10567
R22637 VDD.n5919 VDD.t1338 8.10567
R22638 VDD.n5964 VDD.t3674 8.10567
R22639 VDD.n5918 VDD.t4024 8.10567
R22640 VDD.n5970 VDD.t764 8.10567
R22641 VDD.n5917 VDD.t1637 8.10567
R22642 VDD.n5975 VDD.t3098 8.10567
R22643 VDD.n5916 VDD.t1646 8.10567
R22644 VDD.n6180 VDD.t1067 8.10567
R22645 VDD.n6182 VDD.t2797 8.10567
R22646 VDD.n6183 VDD.t2420 8.10567
R22647 VDD.n6187 VDD.t3405 8.10567
R22648 VDD.n6188 VDD.t3092 8.10567
R22649 VDD.n6192 VDD.t4420 8.10567
R22650 VDD.n6193 VDD.t4086 8.10567
R22651 VDD.n6197 VDD.t2209 8.10567
R22652 VDD.n6198 VDD.t1793 8.10567
R22653 VDD.n6381 VDD.t4720 8.10567
R22654 VDD.n5319 VDD.t930 8.10567
R22655 VDD.n6386 VDD.t2342 8.10567
R22656 VDD.n5316 VDD.t4570 8.10567
R22657 VDD.n5315 VDD.t4094 8.10567
R22658 VDD.n6393 VDD.t2272 8.10567
R22659 VDD.n5995 VDD.t2661 8.10567
R22660 VDD.n5999 VDD.t3482 8.10567
R22661 VDD.n5992 VDD.t4362 8.10567
R22662 VDD.n6004 VDD.t1567 8.10567
R22663 VDD.n5989 VDD.t4368 8.10567
R22664 VDD.n6010 VDD.t4672 8.10567
R22665 VDD.n6381 VDD.t2718 8.10567
R22666 VDD.n5319 VDD.t3044 8.10567
R22667 VDD.n6386 VDD.t4342 8.10567
R22668 VDD.n5316 VDD.t2591 8.10567
R22669 VDD.n5315 VDD.t1979 8.10567
R22670 VDD.n6393 VDD.t4296 8.10567
R22671 VDD.n5995 VDD.t4614 8.10567
R22672 VDD.n5999 VDD.t1345 8.10567
R22673 VDD.n5992 VDD.t2330 8.10567
R22674 VDD.n6004 VDD.t3640 8.10567
R22675 VDD.n5989 VDD.t2340 8.10567
R22676 VDD.n6010 VDD.t2667 8.10567
R22677 VDD.n5335 VDD.t962 8.10567
R22678 VDD.n5333 VDD.t2395 8.10567
R22679 VDD.n5340 VDD.t3278 8.10567
R22680 VDD.n5330 VDD.t823 8.10567
R22681 VDD.n5329 VDD.t4442 8.10567
R22682 VDD.n5347 VDD.t2696 8.10567
R22683 VDD.n5326 VDD.t3998 8.10567
R22684 VDD.n5353 VDD.t716 8.10567
R22685 VDD.n5324 VDD.t4732 8.10567
R22686 VDD.n5358 VDD.t1961 8.10567
R22687 VDD.n5321 VDD.t4278 8.10567
R22688 VDD.n5335 VDD.t3078 8.10567
R22689 VDD.n5333 VDD.t4370 8.10567
R22690 VDD.n5340 VDD.t1125 8.10567
R22691 VDD.n5330 VDD.t2962 8.10567
R22692 VDD.n5329 VDD.t2433 8.10567
R22693 VDD.n5347 VDD.t4662 8.10567
R22694 VDD.n5326 VDD.t1873 8.10567
R22695 VDD.n5353 VDD.t2862 8.10567
R22696 VDD.n5324 VDD.t2737 8.10567
R22697 VDD.n5358 VDD.t4040 8.10567
R22698 VDD.n5321 VDD.t2203 8.10567
R22699 VDD.n5363 VDD.t2558 8.10567
R22700 VDD.n5365 VDD.t4138 8.10567
R22701 VDD.n5366 VDD.t3764 8.10567
R22702 VDD.n5370 VDD.t619 8.10567
R22703 VDD.n5371 VDD.t4422 8.10567
R22704 VDD.n5373 VDD.t1923 8.10567
R22705 VDD.n5363 VDD.t3472 8.10567
R22706 VDD.n5365 VDD.t976 8.10567
R22707 VDD.n5366 VDD.t4734 8.10567
R22708 VDD.n5370 VDD.t1610 8.10567
R22709 VDD.n5371 VDD.t1251 8.10567
R22710 VDD.n5373 VDD.t3010 8.10567
R22711 VDD.n6377 VDD.t4006 8.10567
R22712 VDD.n6375 VDD.t1673 8.10567
R22713 VDD.n6374 VDD.t1308 8.10567
R22714 VDD.n6216 VDD.t3597 8.10567
R22715 VDD.n6217 VDD.t3288 8.10567
R22716 VDD.n6377 VDD.t841 8.10567
R22717 VDD.n6375 VDD.t2773 8.10567
R22718 VDD.n6374 VDD.t2397 8.10567
R22719 VDD.n6216 VDD.t4546 8.10567
R22720 VDD.n6217 VDD.t4238 8.10567
R22721 VDD.n5298 VDD.t1110 8.10567
R22722 VDD.n6409 VDD.t1419 8.10567
R22723 VDD.n5300 VDD.t2900 8.10567
R22724 VDD.n6404 VDD.t1005 8.10567
R22725 VDD.n5301 VDD.t4596 8.10567
R22726 VDD.n6399 VDD.t2860 8.10567
R22727 VDD.n6159 VDD.t3170 8.10567
R22728 VDD.n6163 VDD.t4014 8.10567
R22729 VDD.n6158 VDD.t770 8.10567
R22730 VDD.n6168 VDD.t2135 8.10567
R22731 VDD.n6018 VDD.t778 8.10567
R22732 VDD.n5287 VDD.t1453 8.10567
R22733 VDD.n5286 VDD.t2948 8.10567
R22734 VDD.n6567 VDD.t3768 8.10567
R22735 VDD.n5285 VDD.t1320 8.10567
R22736 VDD.n5284 VDD.t852 8.10567
R22737 VDD.n6574 VDD.t3210 8.10567
R22738 VDD.n6026 VDD.t4500 8.10567
R22739 VDD.n6025 VDD.t1233 8.10567
R22740 VDD.n6032 VDD.t1121 8.10567
R22741 VDD.n6023 VDD.t2583 8.10567
R22742 VDD.n6022 VDD.t649 8.10567
R22743 VDD.n8065 VDD.t1099 8.10567
R22744 VDD.n2159 VDD.t3752 8.10567
R22745 VDD.n2161 VDD.t2172 8.10567
R22746 VDD.n8014 VDD.t912 8.10567
R22747 VDD.n7861 VDD.t1383 8.10567
R22748 VDD.n7862 VDD.t3966 8.10567
R22749 VDD.n7911 VDD.t2307 8.10567
R22750 VDD.n7852 VDD.t2694 8.10567
R22751 VDD.n2207 VDD.t1216 8.10567
R22752 VDD.n2214 VDD.t4386 8.10567
R22753 VDD.n2232 VDD.t1993 8.10567
R22754 VDD.n2221 VDD.t3379 8.10567
R22755 VDD.n7987 VDD.t3792 8.10567
R22756 VDD.n2191 VDD.t1020 8.10567
R22757 VDD.n2195 VDD.t2473 8.10567
R22758 VDD.n2194 VDD.t3646 8.10567
R22759 VDD.n2198 VDD.t3687 8.10567
R22760 VDD.n2200 VDD.t3350 8.10567
R22761 VDD.n7961 VDD.t4132 8.10567
R22762 VDD.n6599 VDD.t1306 8.10567
R22763 VDD.n2205 VDD.t2785 8.10567
R22764 VDD.n2217 VDD.t4480 8.10567
R22765 VDD.n2213 VDD.t1693 8.10567
R22766 VDD.n2211 VDD.t3062 8.10567
R22767 VDD.n2220 VDD.t4360 8.10567
R22768 VDD.n7988 VDD.t1108 8.10567
R22769 VDD.n2190 VDD.t2008 8.10567
R22770 VDD.n2196 VDD.t3401 8.10567
R22771 VDD.n2197 VDD.t1431 8.10567
R22772 VDD.n7974 VDD.t2441 8.10567
R22773 VDD.n2201 VDD.t1013 8.10567
R22774 VDD.n7967 VDD.t1883 8.10567
R22775 VDD.n7962 VDD.t2757 8.10567
R22776 VDD.n6602 VDD.t2268 8.10567
R22777 VDD.n6598 VDD.t3990 8.10567
R22778 VDD.n6597 VDD.t3480 8.10567
R22779 VDD.n6609 VDD.t1604 8.10567
R22780 VDD.n6596 VDD.t3072 8.10567
R22781 VDD.n6615 VDD.t2565 8.10567
R22782 VDD.n6595 VDD.t3754 8.10567
R22783 VDD.n6620 VDD.t1001 8.10567
R22784 VDD.n6594 VDD.t1866 8.10567
R22785 VDD.n2358 VDD.t2805 8.10567
R22786 VDD.n2359 VDD.t2435 8.10567
R22787 VDD.n2364 VDD.t2688 8.10567
R22788 VDD.n2363 VDD.t2274 8.10567
R22789 VDD.n2361 VDD.t1952 8.10567
R22790 VDD.n2358 VDD.t2452 8.10567
R22791 VDD.n2359 VDD.t2006 8.10567
R22792 VDD.n2364 VDD.t2309 8.10567
R22793 VDD.n2363 VDD.t1881 8.10567
R22794 VDD.n2361 VDD.t1596 8.10567
R22795 VDD.n7140 VDD.t885 8.10567
R22796 VDD.n7138 VDD.t2603 8.10567
R22797 VDD.n7137 VDD.t2166 8.10567
R22798 VDD.n2315 VDD.t2217 8.10567
R22799 VDD.n2314 VDD.t1805 8.10567
R22800 VDD.n7140 VDD.t4664 8.10567
R22801 VDD.n7138 VDD.t2180 8.10567
R22802 VDD.n7137 VDD.t1775 8.10567
R22803 VDD.n2315 VDD.t1828 8.10567
R22804 VDD.n2314 VDD.t1465 8.10567
R22805 VDD.n5407 VDD.t2462 8.10567
R22806 VDD.n5405 VDD.t3762 8.10567
R22807 VDD.n5412 VDD.t4650 8.10567
R22808 VDD.n5402 VDD.t2286 8.10567
R22809 VDD.n5401 VDD.t1703 8.10567
R22810 VDD.n5419 VDD.t4054 8.10567
R22811 VDD.n5398 VDD.t1247 8.10567
R22812 VDD.n5425 VDD.t768 8.10567
R22813 VDD.n5396 VDD.t2031 8.10567
R22814 VDD.n5430 VDD.t3417 8.10567
R22815 VDD.n5393 VDD.t4302 8.10567
R22816 VDD.n5407 VDD.t1260 8.10567
R22817 VDD.n5405 VDD.t2751 8.10567
R22818 VDD.n5412 VDD.t3575 8.10567
R22819 VDD.n5402 VDD.t1136 8.10567
R22820 VDD.n5401 VDD.t604 8.10567
R22821 VDD.n5419 VDD.t3026 8.10567
R22822 VDD.n5398 VDD.t4318 8.10567
R22823 VDD.n5425 VDD.t3808 8.10567
R22824 VDD.n5396 VDD.t949 8.10567
R22825 VDD.n5430 VDD.t2372 8.10567
R22826 VDD.n5393 VDD.t3262 8.10567
R22827 VDD.n2297 VDD.t1977 8.10567
R22828 VDD.n2298 VDD.t2834 8.10567
R22829 VDD.n2299 VDD.t3644 8.10567
R22830 VDD.n2300 VDD.t910 8.10567
R22831 VDD.n2301 VDD.t3652 8.10567
R22832 VDD.n2302 VDD.t2761 8.10567
R22833 VDD.n2303 VDD.t4398 8.10567
R22834 VDD.n2304 VDD.t1621 8.10567
R22835 VDD.n2306 VDD.t2076 8.10567
R22836 VDD.n2307 VDD.t3454 8.10567
R22837 VDD.n2308 VDD.t644 8.10567
R22838 VDD.n2309 VDD.t1916 8.10567
R22839 VDD.n2297 VDD.t915 8.10567
R22840 VDD.n2298 VDD.t1635 8.10567
R22841 VDD.n2299 VDD.t2643 8.10567
R22842 VDD.n2300 VDD.t3950 8.10567
R22843 VDD.n2301 VDD.t2655 8.10567
R22844 VDD.n2302 VDD.t1548 8.10567
R22845 VDD.n2303 VDD.t3332 8.10567
R22846 VDD.n2304 VDD.t4688 8.10567
R22847 VDD.n2306 VDD.t988 8.10567
R22848 VDD.n2307 VDD.t2414 8.10567
R22849 VDD.n2308 VDD.t3713 8.10567
R22850 VDD.n2309 VDD.t850 8.10567
R22851 VDD.n2295 VDD.t2627 8.10567
R22852 VDD.n2294 VDD.t2195 8.10567
R22853 VDD.n7838 VDD.t2245 8.10567
R22854 VDD.n7839 VDD.t1836 8.10567
R22855 VDD.n7841 VDD.t3711 8.10567
R22856 VDD.n7844 VDD.t4466 8.10567
R22857 VDD.n2208 VDD.t1204 8.10567
R22858 VDD.n7177 VDD.t2315 8.10567
R22859 VDD.n7945 VDD.t1397 8.10567
R22860 VDD.n7944 VDD.t3986 8.10567
R22861 VDD.n7854 VDD.t2338 8.10567
R22862 VDD.n2148 VDD.t1119 8.10567
R22863 VDD.n8050 VDD.t3780 8.10567
R22864 VDD.n8049 VDD.t2199 8.10567
R22865 VDD.n2149 VDD.t927 8.10567
R22866 VDD.n2174 VDD.t2803 8.10567
R22867 VDD.n2171 VDD.t4108 8.10567
R22868 VDD.n2179 VDD.t1188 8.10567
R22869 VDD.n2170 VDD.t2671 8.10567
R22870 VDD.n2169 VDD.t3494 8.10567
R22871 VDD.n2186 VDD.t4374 8.10567
R22872 VDD.n2168 VDD.t1586 8.10567
R22873 VDD.n8002 VDD.t3834 8.10567
R22874 VDD.n2167 VDD.t4728 8.10567
R22875 VDD.n8007 VDD.t3377 8.10567
R22876 VDD.n2166 VDD.t4276 8.10567
R22877 VDD.n2389 VDD.t2896 8.10567
R22878 VDD.n2387 VDD.t4458 8.10567
R22879 VDD.n2386 VDD.t4120 8.10567
R22880 VDD.n7830 VDD.t1011 8.10567
R22881 VDD.n7829 VDD.t596 8.10567
R22882 VDD.n9133 VDD.t3518 8.10567
R22883 VDD.n9128 VDD.t3322 8.10567
R22884 VDD.n9133 VDD.t3000 8.10567
R22885 VDD.n9128 VDD.t2795 8.10567
R22886 VDD.n9127 VDD.t3314 8.10567
R22887 VDD.n9127 VDD.t3134 8.10567
R22888 VDD.n9125 VDD.t722 8.10567
R22889 VDD.n9125 VDD.t4646 8.10567
R22890 VDD.n9137 VDD.t2631 8.10567
R22891 VDD.n9137 VDD.t2401 8.10567
R22892 VDD.n9135 VDD.t2978 8.10567
R22893 VDD.n9135 VDD.t2767 8.10567
R22894 VDD.n9140 VDD.t2548 8.10567
R22895 VDD.n9085 VDD.t4042 8.10567
R22896 VDD.n9146 VDD.t3898 8.10567
R22897 VDD.n9084 VDD.t3672 8.10567
R22898 VDD.n9081 VDD.t2145 8.10567
R22899 VDD.n9081 VDD.t3695 8.10567
R22900 VDD.n9078 VDD.t2581 8.10567
R22901 VDD.n9078 VDD.t4062 8.10567
R22902 VDD.n9077 VDD.t3166 8.10567
R22903 VDD.n9077 VDD.t4656 8.10567
R22904 VDD.n9174 VDD.t2601 8.10567
R22905 VDD.n9174 VDD.t4076 8.10567
R22906 VDD.n9173 VDD.t2970 8.10567
R22907 VDD.n9173 VDD.t4434 8.10567
R22908 VDD.n9170 VDD.t4464 8.10567
R22909 VDD.n9170 VDD.t1868 8.10567
R22910 VDD.n9081 VDD.t2538 8.10567
R22911 VDD.n9081 VDD.t2256 8.10567
R22912 VDD.n9078 VDD.t2882 8.10567
R22913 VDD.n9078 VDD.t2675 8.10567
R22914 VDD.n9077 VDD.t3440 8.10567
R22915 VDD.n9077 VDD.t3260 8.10567
R22916 VDD.n9174 VDD.t2904 8.10567
R22917 VDD.n9174 VDD.t2686 8.10567
R22918 VDD.n9173 VDD.t3254 8.10567
R22919 VDD.n9173 VDD.t3054 8.10567
R22920 VDD.n9170 VDD.t606 8.10567
R22921 VDD.n9170 VDD.t4540 8.10567
R22922 VDD.n8471 VDD.t3102 8.10567
R22923 VDD.n9163 VDD.t4568 8.10567
R22924 VDD.n8485 VDD.t4460 8.10567
R22925 VDD.n8484 VDD.t4256 8.10567
R22926 VDD.n8580 VDD.t4060 8.10567
R22927 VDD.n8760 VDD.t3840 8.10567
R22928 VDD.n8581 VDD.t4516 8.10567
R22929 VDD.n8754 VDD.t3860 8.10567
R22930 VDD.n8577 VDD.t4282 8.10567
R22931 VDD.n8577 VDD.t1197 8.10567
R22932 VDD.n8574 VDD.t4618 8.10567
R22933 VDD.n8574 VDD.t1539 8.10567
R22934 VDD.n8573 VDD.t1097 8.10567
R22935 VDD.n8573 VDD.t2211 8.10567
R22936 VDD.n8567 VDD.t4644 8.10567
R22937 VDD.n8567 VDD.t1563 8.10567
R22938 VDD.n8566 VDD.t900 8.10567
R22939 VDD.n8566 VDD.t1965 8.10567
R22940 VDD.n8563 VDD.t2550 8.10567
R22941 VDD.n8563 VDD.t3558 8.10567
R22942 VDD.n8577 VDD.t2704 8.10567
R22943 VDD.n8577 VDD.t1410 8.10567
R22944 VDD.n8574 VDD.t3048 8.10567
R22945 VDD.n8574 VDD.t1763 8.10567
R22946 VDD.n8573 VDD.t3595 8.10567
R22947 VDD.n8573 VDD.t2492 8.10567
R22948 VDD.n8567 VDD.t3066 8.10567
R22949 VDD.n8567 VDD.t1779 8.10567
R22950 VDD.n8566 VDD.t3383 8.10567
R22951 VDD.n8566 VDD.t2205 8.10567
R22952 VDD.n8563 VDD.t812 8.10567
R22953 VDD.n8563 VDD.t3782 8.10567
R22954 VDD.n8548 VDD.t2253 8.10567
R22955 VDD.n8556 VDD.t2022 8.10567
R22956 VDD.n8549 VDD.t2813 8.10567
R22957 VDD.n8550 VDD.t2060 8.10567
R22958 VDD.n8830 VDD.t2870 8.10567
R22959 VDD.n8811 VDD.t2111 8.10567
R22960 VDD.n8544 VDD.t1034 8.10567
R22961 VDD.n8543 VDD.t2133 8.10567
R22962 VDD.n8795 VDD.t2466 8.10567
R22963 VDD.n8795 VDD.t3164 8.10567
R22964 VDD.n8792 VDD.t2822 8.10567
R22965 VDD.n8792 VDD.t3476 8.10567
R22966 VDD.n8791 VDD.t3361 8.10567
R22967 VDD.n8791 VDD.t4084 8.10567
R22968 VDD.n8785 VDD.t2838 8.10567
R22969 VDD.n8785 VDD.t3496 8.10567
R22970 VDD.n8784 VDD.t3186 8.10567
R22971 VDD.n8784 VDD.t3854 8.10567
R22972 VDD.n8781 VDD.t4708 8.10567
R22973 VDD.n8781 VDD.t1267 8.10567
R22974 VDD.n8795 VDD.t3236 8.10567
R22975 VDD.n8795 VDD.t1491 8.10567
R22976 VDD.n8792 VDD.t3538 8.10567
R22977 VDD.n8792 VDD.t1858 8.10567
R22978 VDD.n8791 VDD.t4170 8.10567
R22979 VDD.n8791 VDD.t2579 8.10567
R22980 VDD.n8785 VDD.t3548 8.10567
R22981 VDD.n8785 VDD.t1879 8.10567
R22982 VDD.n8784 VDD.t3936 8.10567
R22983 VDD.n8784 VDD.t2319 8.10567
R22984 VDD.n8781 VDD.t1335 8.10567
R22985 VDD.n8781 VDD.t3866 8.10567
R22986 VDD.n8800 VDD.t4584 8.10567
R22987 VDD.n8770 VDD.t3934 8.10567
R22988 VDD.n8531 VDD.t2942 8.10567
R22989 VDD.n8766 VDD.t3958 8.10567
R22990 VDD.n8517 VDD.t2522 8.10567
R22991 VDD.n8886 VDD.t3446 8.10567
R22992 VDD.n8772 VDD.t2439 8.10567
R22993 VDD.n8771 VDD.t3470 8.10567
R22994 VDD.n8849 VDD.t2554 8.10567
R22995 VDD.n8849 VDD.t3650 8.10567
R22996 VDD.n8853 VDD.t2902 8.10567
R22997 VDD.n8853 VDD.t4032 8.10567
R22998 VDD.n8854 VDD.t3460 8.10567
R22999 VDD.n8854 VDD.t4612 8.10567
R23000 VDD.n8862 VDD.t2914 8.10567
R23001 VDD.n8862 VDD.t4046 8.10567
R23002 VDD.n8863 VDD.t3276 8.10567
R23003 VDD.n8863 VDD.t4388 8.10567
R23004 VDD.n8867 VDD.t633 8.10567
R23005 VDD.n8867 VDD.t1819 8.10567
R23006 VDD.n8849 VDD.t1017 8.10567
R23007 VDD.n8849 VDD.t2102 8.10567
R23008 VDD.n8853 VDD.t1333 8.10567
R23009 VDD.n8853 VDD.t2534 8.10567
R23010 VDD.n8854 VDD.t1973 8.10567
R23011 VDD.n8854 VDD.t3130 8.10567
R23012 VDD.n8862 VDD.t1354 8.10567
R23013 VDD.n8862 VDD.t2552 8.10567
R23014 VDD.n8863 VDD.t1726 8.10567
R23015 VDD.n8863 VDD.t2920 8.10567
R23016 VDD.n8867 VDD.t3348 8.10567
R23017 VDD.n8867 VDD.t4416 8.10567
R23018 VDD.n8873 VDD.t580 8.10567
R23019 VDD.n8843 VDD.t1592 8.10567
R23020 VDD.n8521 VDD.t4692 8.10567
R23021 VDD.n8839 VDD.t1619 8.10567
R23022 VDD.n8506 VDD.t2469 8.10567
R23023 VDD.n8942 VDD.t1677 8.10567
R23024 VDD.n8845 VDD.t599 8.10567
R23025 VDD.n8844 VDD.t2213 8.10567
R23026 VDD.n8926 VDD.t4250 8.10567
R23027 VDD.n8926 VDD.t1253 8.10567
R23028 VDD.n8923 VDD.t4556 8.10567
R23029 VDD.n8923 VDD.t1608 8.10567
R23030 VDD.n8922 VDD.t1057 8.10567
R23031 VDD.n8922 VDD.t2270 8.10567
R23032 VDD.n8916 VDD.t4580 8.10567
R23033 VDD.n8916 VDD.t1627 8.10567
R23034 VDD.n8915 VDD.t844 8.10567
R23035 VDD.n8915 VDD.t2020 8.10567
R23036 VDD.n8912 VDD.t2506 8.10567
R23037 VDD.n8912 VDD.t3611 8.10567
R23038 VDD.n8926 VDD.t2856 8.10567
R23039 VDD.n8926 VDD.t3868 8.10567
R23040 VDD.n8923 VDD.t3184 8.10567
R23041 VDD.n8923 VDD.t4236 8.10567
R23042 VDD.n8922 VDD.t3745 8.10567
R23043 VDD.n8922 VDD.t669 8.10567
R23044 VDD.n8916 VDD.t3198 8.10567
R23045 VDD.n8916 VDD.t4248 8.10567
R23046 VDD.n8915 VDD.t3530 8.10567
R23047 VDD.n8915 VDD.t4590 8.10567
R23048 VDD.n8912 VDD.t981 8.10567
R23049 VDD.n8912 VDD.t2066 8.10567
R23050 VDD.n8931 VDD.t4226 8.10567
R23051 VDD.n8901 VDD.t3526 8.10567
R23052 VDD.n8512 VDD.t2530 8.10567
R23053 VDD.n8897 VDD.t4018 8.10567
R23054 VDD.n8498 VDD.t4290 8.10567
R23055 VDD.n9017 VDD.t4082 8.10567
R23056 VDD.n8903 VDD.t2625 8.10567
R23057 VDD.n8902 VDD.t4110 8.10567
R23058 VDD.n8976 VDD.t2081 8.10567
R23059 VDD.n8976 VDD.t1825 8.10567
R23060 VDD.n8980 VDD.t2504 8.10567
R23061 VDD.n8980 VDD.t2225 8.10567
R23062 VDD.n8981 VDD.t3100 8.10567
R23063 VDD.n8981 VDD.t2894 8.10567
R23064 VDD.n8989 VDD.t2518 8.10567
R23065 VDD.n8989 VDD.t2240 8.10567
R23066 VDD.n8990 VDD.t2884 8.10567
R23067 VDD.n8990 VDD.t2677 8.10567
R23068 VDD.n8994 VDD.t4384 8.10567
R23069 VDD.n8994 VDD.t4202 8.10567
R23070 VDD.n8976 VDD.t2950 8.10567
R23071 VDD.n8976 VDD.t2733 8.10567
R23072 VDD.n8980 VDD.t3272 8.10567
R23073 VDD.n8980 VDD.t3070 8.10567
R23074 VDD.n8981 VDD.t3832 8.10567
R23075 VDD.n8981 VDD.t3616 8.10567
R23076 VDD.n8989 VDD.t3280 8.10567
R23077 VDD.n8989 VDD.t3084 8.10567
R23078 VDD.n8990 VDD.t3605 8.10567
R23079 VDD.n8990 VDD.t3407 8.10567
R23080 VDD.n8994 VDD.t1044 8.10567
R23081 VDD.n8994 VDD.t838 8.10567
R23082 VDD.n8970 VDD.t2560 8.10567
R23083 VDD.n8952 VDD.t2290 8.10567
R23084 VDD.n8502 VDD.t709 8.10567
R23085 VDD.n8948 VDD.t2327 8.10567
R23086 VDD.n8489 VDD.t3024 8.10567
R23087 VDD.n9039 VDD.t4486 8.10567
R23088 VDD.n8972 VDD.t4366 8.10567
R23089 VDD.n8971 VDD.t4178 8.10567
R23090 VDD.n9060 VDD.t2158 8.10567
R23091 VDD.n9060 VDD.t1918 8.10567
R23092 VDD.n9057 VDD.t2587 8.10567
R23093 VDD.n9057 VDD.t2354 8.10567
R23094 VDD.n9056 VDD.t3176 8.10567
R23095 VDD.n9056 VDD.t2990 8.10567
R23096 VDD.n9050 VDD.t2609 8.10567
R23097 VDD.n9050 VDD.t2374 8.10567
R23098 VDD.n9049 VDD.t2982 8.10567
R23099 VDD.n9049 VDD.t2769 8.10567
R23100 VDD.n9046 VDD.t4468 8.10567
R23101 VDD.n9046 VDD.t4270 8.10567
R23102 VDD.n9060 VDD.t2449 8.10567
R23103 VDD.n9060 VDD.t2163 8.10567
R23104 VDD.n9057 VDD.t2809 8.10567
R23105 VDD.n9057 VDD.t2589 8.10567
R23106 VDD.n9056 VDD.t3336 8.10567
R23107 VDD.n9056 VDD.t3178 8.10567
R23108 VDD.n9050 VDD.t2824 8.10567
R23109 VDD.n9050 VDD.t2611 8.10567
R23110 VDD.n9049 VDD.t3172 8.10567
R23111 VDD.n9049 VDD.t2986 8.10567
R23112 VDD.n9046 VDD.t4694 8.10567
R23113 VDD.n9046 VDD.t4472 8.10567
R23114 VDD.n9028 VDD.t563 8.10567
R23115 VDD.n9027 VDD.t2192 8.10567
R23116 VDD.n8494 VDD.t2063 8.10567
R23117 VDD.n9023 VDD.t1797 8.10567
R23118 VDD.n9152 VDD.t682 8.10567
R23119 VDD.n9074 VDD.t2304 8.10567
R23120 VDD.n8474 VDD.t2130 8.10567
R23121 VDD.n9070 VDD.t1894 8.10567
R23122 VDD.n185 VDD.t4604 8.10567
R23123 VDD.n187 VDD.t2045 8.10567
R23124 VDD.n125 VDD.t4630 8.10567
R23125 VDD.n171 VDD.t4406 8.10567
R23126 VDD.n9117 VDD.t625 8.10567
R23127 VDD.n9098 VDD.t2231 8.10567
R23128 VDD.n9091 VDD.t2090 8.10567
R23129 VDD.n9092 VDD.t1838 8.10567
R23130 VDD.n1155 VDD.t3607 8.10567
R23131 VDD.t3607 VDD.n1139 8.10567
R23132 VDD.t4264 VDD.n1153 8.10567
R23133 VDD.n1154 VDD.t4264 8.10567
R23134 VDD.t3196 VDD.n1151 8.10567
R23135 VDD.n1152 VDD.t3196 8.10567
R23136 VDD.t3302 VDD.n1149 8.10567
R23137 VDD.n1150 VDD.t3302 8.10567
R23138 VDD.t2161 VDD.n1147 8.10567
R23139 VDD.n1148 VDD.t2161 8.10567
R23140 VDD.t2323 VDD.n1145 8.10567
R23141 VDD.n1146 VDD.t2323 8.10567
R23142 VDD.n1723 VDD.t1142 8.10567
R23143 VDD.t1142 VDD.n1722 8.10567
R23144 VDD.n1725 VDD.t1459 8.10567
R23145 VDD.t1459 VDD.n1724 8.10567
R23146 VDD.n1727 VDD.t4502 8.10567
R23147 VDD.t4502 VDD.n1726 8.10567
R23148 VDD.n1729 VDD.t4636 8.10567
R23149 VDD.t4636 VDD.n1728 8.10567
R23150 VDD.n1731 VDD.t3536 8.10567
R23151 VDD.t3536 VDD.n1730 8.10567
R23152 VDD.n1155 VDD.t753 8.10567
R23153 VDD.t753 VDD.n1139 8.10567
R23154 VDD.n1153 VDD.t3914 8.10567
R23155 VDD.n1154 VDD.t3914 8.10567
R23156 VDD.n1151 VDD.t2876 8.10567
R23157 VDD.n1152 VDD.t2876 8.10567
R23158 VDD.n1149 VDD.t3006 8.10567
R23159 VDD.n1150 VDD.t3006 8.10567
R23160 VDD.n1147 VDD.t1773 8.10567
R23161 VDD.n1148 VDD.t1773 8.10567
R23162 VDD.n1145 VDD.t1914 8.10567
R23163 VDD.n1146 VDD.t1914 8.10567
R23164 VDD.n1723 VDD.t818 8.10567
R23165 VDD.n1722 VDD.t818 8.10567
R23166 VDD.n1725 VDD.t1132 8.10567
R23167 VDD.n1724 VDD.t1132 8.10567
R23168 VDD.n1727 VDD.t4192 8.10567
R23169 VDD.n1726 VDD.t4192 8.10567
R23170 VDD.n1729 VDD.t4294 8.10567
R23171 VDD.n1728 VDD.t4294 8.10567
R23172 VDD.n1731 VDD.t3244 8.10567
R23173 VDD.n1730 VDD.t3244 8.10567
R23174 VDD.n928 VDD.t691 8.10567
R23175 VDD.t691 VDD.n699 8.10567
R23176 VDD.n930 VDD.t3739 8.10567
R23177 VDD.t3739 VDD.n929 8.10567
R23178 VDD.n932 VDD.t4072 8.10567
R23179 VDD.t4072 VDD.n931 8.10567
R23180 VDD.n934 VDD.t3962 8.10567
R23181 VDD.t3962 VDD.n933 8.10567
R23182 VDD.n936 VDD.t4080 8.10567
R23183 VDD.t4080 VDD.n935 8.10567
R23184 VDD.n1048 VDD.t3034 8.10567
R23185 VDD.t3034 VDD.n1047 8.10567
R23186 VDD.n1050 VDD.t3144 8.10567
R23187 VDD.t3144 VDD.n1049 8.10567
R23188 VDD.n1052 VDD.t1963 8.10567
R23189 VDD.t1963 VDD.n1051 8.10567
R23190 VDD.n1054 VDD.t4036 8.10567
R23191 VDD.t4036 VDD.n1053 8.10567
R23192 VDD.n1056 VDD.t2994 8.10567
R23193 VDD.t2994 VDD.n1055 8.10567
R23194 VDD.n1058 VDD.t1347 8.10567
R23195 VDD.t1347 VDD.n1057 8.10567
R23196 VDD.n928 VDD.t4232 8.10567
R23197 VDD.t4232 VDD.n699 8.10567
R23198 VDD.n930 VDD.t3160 8.10567
R23199 VDD.n929 VDD.t3160 8.10567
R23200 VDD.n932 VDD.t3452 8.10567
R23201 VDD.n931 VDD.t3452 8.10567
R23202 VDD.n934 VDD.t3328 8.10567
R23203 VDD.n933 VDD.t3328 8.10567
R23204 VDD.n936 VDD.t3456 8.10567
R23205 VDD.n935 VDD.t3456 8.10567
R23206 VDD.n1048 VDD.t2399 8.10567
R23207 VDD.n1047 VDD.t2399 8.10567
R23208 VDD.n1050 VDD.t2526 8.10567
R23209 VDD.n1049 VDD.t2526 8.10567
R23210 VDD.n1052 VDD.t1299 8.10567
R23211 VDD.n1051 VDD.t1299 8.10567
R23212 VDD.n1054 VDD.t3397 8.10567
R23213 VDD.n1053 VDD.t3397 8.10567
R23214 VDD.n1056 VDD.t2317 8.10567
R23215 VDD.n1055 VDD.t2317 8.10567
R23216 VDD.n1058 VDD.t744 8.10567
R23217 VDD.n1057 VDD.t744 8.10567
R23218 VDD.t2148 VDD.n1706 8.10567
R23219 VDD.n1707 VDD.t2148 8.10567
R23220 VDD.t1028 VDD.n1704 8.10567
R23221 VDD.n1705 VDD.t1028 8.10567
R23222 VDD.t1322 VDD.n1702 8.10567
R23223 VDD.n1703 VDD.t1322 8.10567
R23224 VDD.t1214 VDD.n1700 8.10567
R23225 VDD.n1701 VDD.t1214 8.10567
R23226 VDD.t1327 VDD.n1698 8.10567
R23227 VDD.n1699 VDD.t1327 8.10567
R23228 VDD.n886 VDD.t4380 8.10567
R23229 VDD.t4380 VDD.n885 8.10567
R23230 VDD.n888 VDD.t4498 8.10567
R23231 VDD.t4498 VDD.n887 8.10567
R23232 VDD.n890 VDD.t3421 8.10567
R23233 VDD.t3421 VDD.n889 8.10567
R23234 VDD.n892 VDD.t1282 8.10567
R23235 VDD.t1282 VDD.n891 8.10567
R23236 VDD.n894 VDD.t4346 8.10567
R23237 VDD.t4346 VDD.n893 8.10567
R23238 VDD.n896 VDD.t2890 8.10567
R23239 VDD.t2890 VDD.n895 8.10567
R23240 VDD.n1706 VDD.t1475 8.10567
R23241 VDD.n1707 VDD.t1475 8.10567
R23242 VDD.n1704 VDD.t4514 8.10567
R23243 VDD.n1705 VDD.t4514 8.10567
R23244 VDD.n1702 VDD.t712 8.10567
R23245 VDD.n1703 VDD.t712 8.10567
R23246 VDD.n1700 VDD.t4736 8.10567
R23247 VDD.n1701 VDD.t4736 8.10567
R23248 VDD.n1698 VDD.t714 8.10567
R23249 VDD.n1699 VDD.t714 8.10567
R23250 VDD.n886 VDD.t3766 8.10567
R23251 VDD.n885 VDD.t3766 8.10567
R23252 VDD.n888 VDD.t3886 8.10567
R23253 VDD.n887 VDD.t3886 8.10567
R23254 VDD.n890 VDD.t2852 8.10567
R23255 VDD.n889 VDD.t2852 8.10567
R23256 VDD.n892 VDD.t659 8.10567
R23257 VDD.n891 VDD.t659 8.10567
R23258 VDD.n894 VDD.t3705 8.10567
R23259 VDD.n893 VDD.t3705 8.10567
R23260 VDD.n896 VDD.t2197 8.10567
R23261 VDD.n895 VDD.t2197 8.10567
R23262 VDD.t4214 VDD.n1475 8.10567
R23263 VDD.n1476 VDD.t4214 8.10567
R23264 VDD.t3148 VDD.n1473 8.10567
R23265 VDD.n1474 VDD.t3148 8.10567
R23266 VDD.t3428 VDD.n1471 8.10567
R23267 VDD.n1472 VDD.t3428 8.10567
R23268 VDD.t3324 VDD.n1469 8.10567
R23269 VDD.n1470 VDD.t3324 8.10567
R23270 VDD.t3436 VDD.n1467 8.10567
R23271 VDD.n1468 VDD.t3436 8.10567
R23272 VDD.n1293 VDD.t2370 8.10567
R23273 VDD.t2370 VDD.n742 8.10567
R23274 VDD.n1295 VDD.t2510 8.10567
R23275 VDD.t2510 VDD.n1294 8.10567
R23276 VDD.n1297 VDD.t1280 8.10567
R23277 VDD.t1280 VDD.n1296 8.10567
R23278 VDD.n1299 VDD.t3363 8.10567
R23279 VDD.t3363 VDD.n1298 8.10567
R23280 VDD.n1301 VDD.t2278 8.10567
R23281 VDD.t2278 VDD.n1300 8.10567
R23282 VDD.n1303 VDD.t702 8.10567
R23283 VDD.t702 VDD.n1302 8.10567
R23284 VDD.n1475 VDD.t820 8.10567
R23285 VDD.n1476 VDD.t820 8.10567
R23286 VDD.n1473 VDD.t3856 8.10567
R23287 VDD.n1474 VDD.t3856 8.10567
R23288 VDD.n1471 VDD.t4200 8.10567
R23289 VDD.n1472 VDD.t4200 8.10567
R23290 VDD.n1469 VDD.t4066 8.10567
R23291 VDD.n1470 VDD.t4066 8.10567
R23292 VDD.n1467 VDD.t4208 8.10567
R23293 VDD.n1468 VDD.t4208 8.10567
R23294 VDD.n1293 VDD.t3138 8.10567
R23295 VDD.t3138 VDD.n742 8.10567
R23296 VDD.n1295 VDD.t3252 8.10567
R23297 VDD.n1294 VDD.t3252 8.10567
R23298 VDD.n1297 VDD.t2093 8.10567
R23299 VDD.n1296 VDD.t2093 8.10567
R23300 VDD.n1299 VDD.t4154 8.10567
R23301 VDD.n1298 VDD.t4154 8.10567
R23302 VDD.n1301 VDD.t3088 8.10567
R23303 VDD.n1300 VDD.t3088 8.10567
R23304 VDD.n1303 VDD.t1457 8.10567
R23305 VDD.n1302 VDD.t1457 8.10567
R23306 VDD.n1234 VDD.t1786 8.10567
R23307 VDD.t1786 VDD.n1219 8.10567
R23308 VDD.t3670 VDD.n1232 8.10567
R23309 VDD.n1233 VDD.t3670 8.10567
R23310 VDD.t2649 VDD.n1230 8.10567
R23311 VDD.n1231 VDD.t2649 8.10567
R23312 VDD.t2783 VDD.n1228 8.10567
R23313 VDD.n1229 VDD.t2783 8.10567
R23314 VDD.t1535 VDD.n1226 8.10567
R23315 VDD.n1227 VDD.t1535 8.10567
R23316 VDD.t1669 VDD.n1085 8.10567
R23317 VDD.n1225 VDD.t1669 8.10567
R23318 VDD.t4718 VDD.n1099 8.10567
R23319 VDD.n1100 VDD.t4718 8.10567
R23320 VDD.t925 VDD.n1097 8.10567
R23321 VDD.n1098 VDD.t925 8.10567
R23322 VDD.t3956 VDD.n1095 8.10567
R23323 VDD.n1096 VDD.t3956 8.10567
R23324 VDD.t4070 VDD.n813 8.10567
R23325 VDD.n1234 VDD.t4204 8.10567
R23326 VDD.t4204 VDD.n1219 8.10567
R23327 VDD.n1232 VDD.t2360 8.10567
R23328 VDD.n1233 VDD.t2360 8.10567
R23329 VDD.n1230 VDD.t1151 8.10567
R23330 VDD.n1231 VDD.t1151 8.10567
R23331 VDD.n1228 VDD.t1270 8.10567
R23332 VDD.n1229 VDD.t1270 8.10567
R23333 VDD.n1226 VDD.t4334 8.10567
R23334 VDD.n1227 VDD.t4334 8.10567
R23335 VDD.t4446 VDD.n1085 8.10567
R23336 VDD.n1225 VDD.t4446 8.10567
R23337 VDD.n1099 VDD.t3344 8.10567
R23338 VDD.n1100 VDD.t3344 8.10567
R23339 VDD.n1097 VDD.t3656 8.10567
R23340 VDD.n1098 VDD.t3656 8.10567
R23341 VDD.n1095 VDD.t2639 8.10567
R23342 VDD.n1096 VDD.t2639 8.10567
R23343 VDD.t2765 VDD.n813 8.10567
R23344 VDD.n1267 VDD.t2906 8.10567
R23345 VDD.t2906 VDD.n1251 8.10567
R23346 VDD.t664 VDD.n1265 8.10567
R23347 VDD.n1266 VDD.t664 8.10567
R23348 VDD.t3715 VDD.n1263 8.10567
R23349 VDD.n1264 VDD.t3715 8.10567
R23350 VDD.t3838 VDD.n1261 8.10567
R23351 VDD.n1262 VDD.t3838 8.10567
R23352 VDD.t2811 VDD.n1259 8.10567
R23353 VDD.n1260 VDD.t2811 8.10567
R23354 VDD.t2918 VDD.n1257 8.10567
R23355 VDD.n1258 VDD.t2918 8.10567
R23356 VDD.t1697 VDD.n1617 8.10567
R23357 VDD.n1618 VDD.t1697 8.10567
R23358 VDD.t2072 VDD.n1615 8.10567
R23359 VDD.n1616 VDD.t2072 8.10567
R23360 VDD.t960 VDD.n1613 8.10567
R23361 VDD.n1614 VDD.t960 8.10567
R23362 VDD.n1267 VDD.t1042 8.10567
R23363 VDD.t1042 VDD.n1251 8.10567
R23364 VDD.n1265 VDD.t3466 8.10567
R23365 VDD.n1266 VDD.t3466 8.10567
R23366 VDD.n1263 VDD.t2406 8.10567
R23367 VDD.n1264 VDD.t2406 8.10567
R23368 VDD.n1261 VDD.t2532 8.10567
R23369 VDD.n1262 VDD.t2532 8.10567
R23370 VDD.n1259 VDD.t1304 8.10567
R23371 VDD.n1260 VDD.t1304 8.10567
R23372 VDD.n1257 VDD.t1429 8.10567
R23373 VDD.n1258 VDD.t1429 8.10567
R23374 VDD.n1617 VDD.t4476 8.10567
R23375 VDD.n1618 VDD.t4476 8.10567
R23376 VDD.n1615 VDD.t656 8.10567
R23377 VDD.n1616 VDD.t656 8.10567
R23378 VDD.n1613 VDD.t3699 8.10567
R23379 VDD.n1614 VDD.t3699 8.10567
R23380 VDD.n1612 VDD.t1069 8.10567
R23381 VDD.n1612 VDD.t3836 8.10567
R23382 VDD.t2464 VDD.n1590 8.10567
R23383 VDD.n1591 VDD.t2464 8.10567
R23384 VDD.t1239 VDD.n1588 8.10567
R23385 VDD.n1589 VDD.t1239 8.10567
R23386 VDD.t1569 VDD.n1586 8.10567
R23387 VDD.n1587 VDD.t1569 8.10567
R23388 VDD.t1447 VDD.n1584 8.10567
R23389 VDD.n1585 VDD.t1447 8.10567
R23390 VDD.t1580 VDD.n1582 8.10567
R23391 VDD.n1583 VDD.t1580 8.10567
R23392 VDD.t4620 VDD.n1670 8.10567
R23393 VDD.n1671 VDD.t4620 8.10567
R23394 VDD.t4744 VDD.n1668 8.10567
R23395 VDD.n1669 VDD.t4744 8.10567
R23396 VDD.t3632 VDD.n1666 8.10567
R23397 VDD.n1667 VDD.t3632 8.10567
R23398 VDD.n1576 VDD.t2755 8.10567
R23399 VDD.t2755 VDD.n1575 8.10567
R23400 VDD.n1570 VDD.t577 8.10567
R23401 VDD.t577 VDD.n1569 8.10567
R23402 VDD.n1572 VDD.t3642 8.10567
R23403 VDD.t3642 VDD.n1571 8.10567
R23404 VDD.n1574 VDD.t3784 8.10567
R23405 VDD.t3784 VDD.n1573 8.10567
R23406 VDD.t2325 VDD.n1637 8.10567
R23407 VDD.n1638 VDD.t2325 8.10567
R23408 VDD.n1634 VDD.t2483 8.10567
R23409 VDD.t2483 VDD.n774 8.10567
R23410 VDD.n1631 VDD.t1258 8.10567
R23411 VDD.t1258 VDD.n777 8.10567
R23412 VDD.n1628 VDD.t1389 8.10567
R23413 VDD.t1389 VDD.n779 8.10567
R23414 VDD.n1568 VDD.t4428 8.10567
R23415 VDD.t4428 VDD.n1567 8.10567
R23416 VDD.t3409 VDD.n1641 8.10567
R23417 VDD.n1642 VDD.t3409 8.10567
R23418 VDD.n1133 VDD.t953 8.10567
R23419 VDD.t953 VDD.n1118 8.10567
R23420 VDD.t3626 VDD.n1131 8.10567
R23421 VDD.n1132 VDD.t3626 8.10567
R23422 VDD.t2607 VDD.n1129 8.10567
R23423 VDD.n1130 VDD.t2607 8.10567
R23424 VDD.t2726 VDD.n1127 8.10567
R23425 VDD.n1128 VDD.t2726 8.10567
R23426 VDD.t1499 VDD.n1125 8.10567
R23427 VDD.n1126 VDD.t1499 8.10567
R23428 VDD.t1631 VDD.n852 8.10567
R23429 VDD.n1124 VDD.t1631 8.10567
R23430 VDD.t4680 VDD.n872 8.10567
R23431 VDD.n873 VDD.t4680 8.10567
R23432 VDD.t880 VDD.n870 8.10567
R23433 VDD.n871 VDD.t880 8.10567
R23434 VDD.t3904 VDD.n868 8.10567
R23435 VDD.n869 VDD.t3904 8.10567
R23436 VDD.t4038 VDD.n866 8.10567
R23437 VDD.n867 VDD.t4038 8.10567
R23438 VDD.t2998 VDD.n728 8.10567
R23439 VDD.n865 VDD.t2998 8.10567
R23440 VDD.n1133 VDD.t2247 8.10567
R23441 VDD.t2247 VDD.n1118 8.10567
R23442 VDD.n1131 VDD.t3318 8.10567
R23443 VDD.n1132 VDD.t3318 8.10567
R23444 VDD.n1129 VDD.t2190 8.10567
R23445 VDD.n1130 VDD.t2190 8.10567
R23446 VDD.n1127 VDD.t2368 8.10567
R23447 VDD.n1128 VDD.t2368 8.10567
R23448 VDD.n1125 VDD.t1162 8.10567
R23449 VDD.n1126 VDD.t1162 8.10567
R23450 VDD.t1276 VDD.n852 8.10567
R23451 VDD.n1124 VDD.t1276 8.10567
R23452 VDD.n872 VDD.t4338 8.10567
R23453 VDD.n873 VDD.t4338 8.10567
R23454 VDD.n870 VDD.t4658 8.10567
R23455 VDD.n871 VDD.t4658 8.10567
R23456 VDD.n868 VDD.t3554 8.10567
R23457 VDD.n869 VDD.t3554 8.10567
R23458 VDD.n866 VDD.t3666 8.10567
R23459 VDD.n867 VDD.t3666 8.10567
R23460 VDD.t2647 VDD.n728 8.10567
R23461 VDD.n865 VDD.t2647 8.10567
R23462 VDD.n1204 VDD.t4180 8.10567
R23463 VDD.t4180 VDD.n1189 8.10567
R23464 VDD.t3723 VDD.n1202 8.10567
R23465 VDD.n1203 VDD.t3723 8.10567
R23466 VDD.t2698 VDD.n1200 8.10567
R23467 VDD.n1201 VDD.t2698 8.10567
R23468 VDD.t2820 VDD.n1198 8.10567
R23469 VDD.n1199 VDD.t2820 8.10567
R23470 VDD.t1600 VDD.n1196 8.10567
R23471 VDD.n1197 VDD.t1600 8.10567
R23472 VDD.t1718 VDD.n851 8.10567
R23473 VDD.n1195 VDD.t1718 8.10567
R23474 VDD.n1433 VDD.t594 8.10567
R23475 VDD.t594 VDD.n1432 8.10567
R23476 VDD.n1435 VDD.t984 8.10567
R23477 VDD.t984 VDD.n1434 8.10567
R23478 VDD.n1437 VDD.t4010 8.10567
R23479 VDD.t4010 VDD.n1436 8.10567
R23480 VDD.n1439 VDD.t4136 8.10567
R23481 VDD.t4136 VDD.n1438 8.10567
R23482 VDD.n1204 VDD.t1272 8.10567
R23483 VDD.t1272 VDD.n1189 8.10567
R23484 VDD.n1202 VDD.t3387 8.10567
R23485 VDD.n1203 VDD.t3387 8.10567
R23486 VDD.n1200 VDD.t2313 8.10567
R23487 VDD.n1201 VDD.t2313 8.10567
R23488 VDD.n1198 VDD.t2477 8.10567
R23489 VDD.n1199 VDD.t2477 8.10567
R23490 VDD.n1196 VDD.t1256 8.10567
R23491 VDD.n1197 VDD.t1256 8.10567
R23492 VDD.t1378 VDD.n851 8.10567
R23493 VDD.n1195 VDD.t1378 8.10567
R23494 VDD.n1433 VDD.t4414 8.10567
R23495 VDD.n1432 VDD.t4414 8.10567
R23496 VDD.n1435 VDD.t560 8.10567
R23497 VDD.n1434 VDD.t560 8.10567
R23498 VDD.n1437 VDD.t3634 8.10567
R23499 VDD.n1436 VDD.t3634 8.10567
R23500 VDD.n1439 VDD.t3774 8.10567
R23501 VDD.n1438 VDD.t3774 8.10567
R23502 VDD.t3074 VDD.n1440 8.10567
R23503 VDD.t3968 VDD.n801 8.10567
R23504 VDD.n802 VDD.t3968 8.10567
R23505 VDD.t2916 VDD.n799 8.10567
R23506 VDD.n800 VDD.t2916 8.10567
R23507 VDD.t3226 VDD.n797 8.10567
R23508 VDD.n798 VDD.t3226 8.10567
R23509 VDD.t3116 VDD.n795 8.10567
R23510 VDD.n796 VDD.t3116 8.10567
R23511 VDD.t3232 VDD.n793 8.10567
R23512 VDD.n794 VDD.t3232 8.10567
R23513 VDD.n1325 VDD.t2074 8.10567
R23514 VDD.t2074 VDD.n745 8.10567
R23515 VDD.n1327 VDD.t2201 8.10567
R23516 VDD.t2201 VDD.n1326 8.10567
R23517 VDD.n1329 VDD.t1071 8.10567
R23518 VDD.t1071 VDD.n1328 8.10567
R23519 VDD.n1331 VDD.t3180 8.10567
R23520 VDD.t3180 VDD.n1330 8.10567
R23521 VDD.n1333 VDD.t2002 8.10567
R23522 VDD.t2002 VDD.n1332 8.10567
R23523 VDD.n1335 VDD.t4608 8.10567
R23524 VDD.t4608 VDD.n1334 8.10567
R23525 VDD.n801 VDD.t4716 8.10567
R23526 VDD.n802 VDD.t4716 8.10567
R23527 VDD.n799 VDD.t3618 8.10567
R23528 VDD.n800 VDD.t3618 8.10567
R23529 VDD.n797 VDD.t3952 8.10567
R23530 VDD.n798 VDD.t3952 8.10567
R23531 VDD.n795 VDD.t3822 8.10567
R23532 VDD.n796 VDD.t3822 8.10567
R23533 VDD.n793 VDD.t3960 8.10567
R23534 VDD.n794 VDD.t3960 8.10567
R23535 VDD.n1325 VDD.t2910 8.10567
R23536 VDD.t2910 VDD.n745 8.10567
R23537 VDD.n1327 VDD.t3032 8.10567
R23538 VDD.n1326 VDD.t3032 8.10567
R23539 VDD.n1329 VDD.t1813 8.10567
R23540 VDD.n1328 VDD.t1813 8.10567
R23541 VDD.n1331 VDD.t3894 8.10567
R23542 VDD.n1330 VDD.t3894 8.10567
R23543 VDD.n1333 VDD.t2858 8.10567
R23544 VDD.n1332 VDD.t2858 8.10567
R23545 VDD.n1335 VDD.t1223 8.10567
R23546 VDD.n1334 VDD.t1223 8.10567
R23547 VDD.n1665 VDD.t1521 8.10567
R23548 VDD.t1521 VDD.n1664 8.10567
R23549 VDD.t4552 VDD.n1662 8.10567
R23550 VDD.n1663 VDD.t4552 8.10567
R23551 VDD.t2475 VDD.n838 8.10567
R23552 VDD.n839 VDD.t2475 8.10567
R23553 VDD.t1249 VDD.n836 8.10567
R23554 VDD.n837 VDD.t1249 8.10567
R23555 VDD.t1584 VDD.n834 8.10567
R23556 VDD.n835 VDD.t1584 8.10567
R23557 VDD.t1455 VDD.n832 8.10567
R23558 VDD.n833 VDD.t1455 8.10567
R23559 VDD.t1588 VDD.n830 8.10567
R23560 VDD.n831 VDD.t1588 8.10567
R23561 VDD.n1372 VDD.t4632 8.10567
R23562 VDD.t4632 VDD.n1371 8.10567
R23563 VDD.n1374 VDD.t566 8.10567
R23564 VDD.t566 VDD.n1373 8.10567
R23565 VDD.n1376 VDD.t3636 8.10567
R23566 VDD.t3636 VDD.n1375 8.10567
R23567 VDD.n1378 VDD.t1525 8.10567
R23568 VDD.t1525 VDD.n1377 8.10567
R23569 VDD.n1380 VDD.t4564 8.10567
R23570 VDD.t4564 VDD.n1379 8.10567
R23571 VDD.n1382 VDD.t3120 8.10567
R23572 VDD.t3120 VDD.n1381 8.10567
R23573 VDD.n838 VDD.t1722 8.10567
R23574 VDD.n839 VDD.t1722 8.10567
R23575 VDD.n836 VDD.t609 8.10567
R23576 VDD.n837 VDD.t609 8.10567
R23577 VDD.n834 VDD.t990 8.10567
R23578 VDD.n835 VDD.t990 8.10567
R23579 VDD.n832 VDD.t873 8.10567
R23580 VDD.n833 VDD.t873 8.10567
R23581 VDD.n830 VDD.t999 8.10567
R23582 VDD.n831 VDD.t999 8.10567
R23583 VDD.n1372 VDD.t4022 8.10567
R23584 VDD.n1371 VDD.t4022 8.10567
R23585 VDD.n1374 VDD.t4146 8.10567
R23586 VDD.n1373 VDD.t4146 8.10567
R23587 VDD.n1376 VDD.t3086 8.10567
R23588 VDD.n1375 VDD.t3086 8.10567
R23589 VDD.n1378 VDD.t942 8.10567
R23590 VDD.n1377 VDD.t942 8.10567
R23591 VDD.n1380 VDD.t3972 8.10567
R23592 VDD.n1379 VDD.t3972 8.10567
R23593 VDD.n1382 VDD.t2514 8.10567
R23594 VDD.n1381 VDD.t2514 8.10567
R23595 VDD.n8070 VDD.t1361 6.64567
R23596 VDD.n2126 VDD.t2842 6.64567
R23597 VDD.n2125 VDD.t944 6.64567
R23598 VDD.n2127 VDD.t2086 6.64567
R23599 VDD.n2141 VDD.t1026 6.64567
R23600 VDD.n2139 VDD.t2412 6.64567
R23601 VDD.n2138 VDD.t3326 6.64567
R23602 VDD.n2138 VDD.t2299 6.64567
R23603 VDD.n2134 VDD.t774 6.64567
R23604 VDD.n2134 VDD.t3870 6.64567
R23605 VDD.n2133 VDD.t3802 6.64567
R23606 VDD.n2133 VDD.t2846 6.64567
R23607 VDD.n2131 VDD.t1991 6.64567
R23608 VDD.n2131 VDD.t964 6.64567
R23609 VDD.n8085 VDD.t1278 6.64567
R23610 VDD.n8080 VDD.t2771 6.64567
R23611 VDD.n2122 VDD.t862 6.64567
R23612 VDD.n8066 VDD.t571 6.64567
R23613 VDD.n2156 VDD.t1912 6.64567
R23614 VDD.n2158 VDD.t1830 6.64567
R23615 VDD.n2165 VDD.t3474 6.64567
R23616 VDD.n8016 VDD.t2429 6.64567
R23617 VDD.n8013 VDD.t4686 6.64567
R23618 VDD.n6021 VDD.t4886 6.58663
R23619 VDD.n6094 VDD.t4962 6.58663
R23620 VDD.n6846 VDD.t272 6.58663
R23621 VDD.n6796 VDD.t180 6.58663
R23622 VDD.n7009 VDD.n7005 6.50088
R23623 VDD.n6958 VDD.n6957 6.50088
R23624 VDD.n6548 VDD.n6547 6.50088
R23625 VDD.n6501 VDD.n6497 6.50088
R23626 VDD.n6116 VDD.n6109 6.45575
R23627 VDD.n6073 VDD.n6066 6.45575
R23628 VDD.n6801 VDD.n6800 6.45575
R23629 VDD.n6752 VDD.n6746 6.45575
R23630 VDD.n1719 VDD.n709 6.24156
R23631 VDD.n1415 VDD.n874 6.24156
R23632 VDD.n1429 VDD.n1428 6.24156
R23633 VDD.n1354 VDD.n1084 6.24156
R23634 VDD.n1346 VDD.n1345 6.24156
R23635 VDD.n6153 VDD.n6152 5.95439
R23636 VDD.n6096 VDD.n6095 5.95439
R23637 VDD.n6847 VDD.n6844 5.95439
R23638 VDD.n6797 VDD.n6794 5.95439
R23639 VDD.n8643 VDD.n8642 5.76894
R23640 VDD.n8702 VDD.n8701 5.76894
R23641 VDD.n1812 VDD.n1811 5.76894
R23642 VDD.n1868 VDD.n1867 5.76894
R23643 VDD.n5516 VDD.n5515 5.76894
R23644 VDD.n1960 VDD.n1959 5.76894
R23645 VDD.n2042 VDD.n2041 5.76894
R23646 VDD.n8752 VDD.n8751 5.76894
R23647 VDD.n8895 VDD.n8894 5.76894
R23648 VDD.n9068 VDD.n9067 5.76894
R23649 VDD.n8642 VDD.n8641 5.33948
R23650 VDD.n8701 VDD.n8700 5.33948
R23651 VDD.n1811 VDD.n1810 5.33948
R23652 VDD.n1867 VDD.n1866 5.33948
R23653 VDD.n5515 VDD.n5514 5.33948
R23654 VDD.n1959 VDD.n1958 5.33948
R23655 VDD.n2041 VDD.n2040 5.33948
R23656 VDD.n8751 VDD.n8750 5.33948
R23657 VDD.n8894 VDD.n8893 5.33948
R23658 VDD.n9067 VDD.n9066 5.33948
R23659 VDD.n6153 VDD.t4866 5.31528
R23660 VDD.n6096 VDD.t4944 5.31528
R23661 VDD.n6844 VDD.t93 5.31528
R23662 VDD.n6794 VDD.t228 5.31528
R23663 VDD.n2130 VDD.t413 5.19255
R23664 VDD.n983 VDD.t453 5.17005
R23665 VDD.n1034 VDD.t462 5.17005
R23666 VDD.n1044 VDD.t448 5.17005
R23667 VDD.n1105 VDD.t352 5.17005
R23668 VDD.n1620 VDD.t360 5.17005
R23669 VDD.n1086 VDD.t371 5.17005
R23670 VDD.n1419 VDD.t446 5.17005
R23671 VDD.n853 VDD.t459 5.17005
R23672 VDD.n1677 VDD.t343 5.17005
R23673 VDD.n1683 VDD.t333 5.17005
R23674 VDD.n1689 VDD.t363 5.17005
R23675 VDD.n1696 VDD.t439 5.17005
R23676 VDD.n979 VDD.t430 5.1669
R23677 VDD.n1039 VDD.t449 5.1669
R23678 VDD.n735 VDD.t465 5.1669
R23679 VDD.n784 VDD.t350 5.1669
R23680 VDD.n1625 VDD.t327 5.1669
R23681 VDD.n1091 VDD.t487 5.1669
R23682 VDD.n1424 VDD.t447 5.1669
R23683 VDD.n858 VDD.t440 5.1669
R23684 VDD.n1673 VDD.t348 5.1669
R23685 VDD.n1679 VDD.t364 5.1669
R23686 VDD.n1685 VDD.t359 5.1669
R23687 VDD.n1692 VDD.t450 5.1669
R23688 VDD.n7952 VDD.t109 5.12594
R23689 VDD.n6370 VDD.n5376 5.12014
R23690 VDD.n7133 VDD.n2317 5.12014
R23691 VDD.n8057 VDD.t209 5.09041
R23692 VDD.n8069 VDD.t1362 5.0505
R23693 VDD.t945 VDD.n2145 5.0505
R23694 VDD.n2144 VDD.t2087 5.0505
R23695 VDD.t2087 VDD.n2143 5.0505
R23696 VDD.n2128 VDD.t863 5.0505
R23697 VDD.n8084 VDD.t1279 5.0505
R23698 VDD.n6743 VDD.n6742 4.96877
R23699 VDD.n6070 VDD.n6069 4.96877
R23700 VDD.n6113 VDD.n6112 4.96877
R23701 VDD.n6737 VDD.n6736 4.96877
R23702 VDD.n2379 VDD.n2377 4.92758
R23703 VDD.n6962 VDD.n6960 4.92758
R23704 VDD.n5292 VDD.n5290 4.92758
R23705 VDD.n6507 VDD.n6505 4.92758
R23706 VDD.n6887 VDD.n6886 4.78594
R23707 VDD.n6906 VDD.n6905 4.78594
R23708 VDD.n6420 VDD.n6419 4.78594
R23709 VDD.n6457 VDD.n6456 4.78594
R23710 VDD.n6744 VDD.n6743 4.61712
R23711 VDD.n6756 VDD.n6755 4.61712
R23712 VDD.n6071 VDD.n6070 4.61712
R23713 VDD.n6061 VDD.n6060 4.61712
R23714 VDD.n6114 VDD.n6113 4.61712
R23715 VDD.n6104 VDD.n6103 4.61712
R23716 VDD.n6738 VDD.n6737 4.61712
R23717 VDD.n6805 VDD.n6804 4.61712
R23718 VDD.n61 VDD.n60 4.61205
R23719 VDD.n70 VDD.n69 4.61205
R23720 VDD.n150 VDD.n149 4.61205
R23721 VDD.n159 VDD.n158 4.61205
R23722 VDD.n5769 VDD.n5768 4.61205
R23723 VDD.n5760 VDD.n5759 4.61205
R23724 VDD.n5836 VDD.n5835 4.61205
R23725 VDD.n5827 VDD.n5826 4.61205
R23726 VDD.n5653 VDD.n5652 4.61205
R23727 VDD.n5644 VDD.n5643 4.61205
R23728 VDD.n5571 VDD.n5570 4.61205
R23729 VDD.n5562 VDD.n5561 4.61205
R23730 VDD.n8157 VDD.n8156 4.61205
R23731 VDD.n8148 VDD.n8147 4.61205
R23732 VDD.n9105 VDD.n9104 4.61205
R23733 VDD.n9114 VDD.n9113 4.61205
R23734 VDD.n8818 VDD.n8817 4.61205
R23735 VDD.n8827 VDD.n8826 4.61205
R23736 VDD.n8958 VDD.n8957 4.61205
R23737 VDD.n8967 VDD.n8966 4.61205
R23738 VDD.n6754 VDD.n6753 4.61078
R23739 VDD.n6997 VDD.n6994 4.61078
R23740 VDD.n6992 VDD.n6989 4.61078
R23741 VDD.n6987 VDD.n6984 4.61078
R23742 VDD.n6982 VDD.n6979 4.61078
R23743 VDD.n6900 VDD.n6897 4.61078
R23744 VDD.n6895 VDD.n6892 4.61078
R23745 VDD.n6890 VDD.n6887 4.61078
R23746 VDD.n6949 VDD.n6946 4.61078
R23747 VDD.n6944 VDD.n6941 4.61078
R23748 VDD.n6939 VDD.n6936 4.61078
R23749 VDD.n6934 VDD.n6931 4.61078
R23750 VDD.n6919 VDD.n6916 4.61078
R23751 VDD.n6914 VDD.n6911 4.61078
R23752 VDD.n6909 VDD.n6906 4.61078
R23753 VDD.n6525 VDD.n6524 4.61078
R23754 VDD.n6528 VDD.n6527 4.61078
R23755 VDD.n6531 VDD.n6530 4.61078
R23756 VDD.n6534 VDD.n6533 4.61078
R23757 VDD.n6433 VDD.n6430 4.61078
R23758 VDD.n6428 VDD.n6425 4.61078
R23759 VDD.n6423 VDD.n6420 4.61078
R23760 VDD.n6485 VDD.n6484 4.61078
R23761 VDD.n6488 VDD.n6487 4.61078
R23762 VDD.n6491 VDD.n6490 4.61078
R23763 VDD.n6494 VDD.n6493 4.61078
R23764 VDD.n6470 VDD.n6467 4.61078
R23765 VDD.n6465 VDD.n6462 4.61078
R23766 VDD.n6460 VDD.n6457 4.61078
R23767 VDD.n6065 VDD.n6062 4.61078
R23768 VDD.n6108 VDD.n6105 4.61078
R23769 VDD.n7893 VDD.n7892 4.61078
R23770 VDD.n7896 VDD.n7895 4.61078
R23771 VDD.n7899 VDD.n7898 4.61078
R23772 VDD.n7902 VDD.n7901 4.61078
R23773 VDD.n7905 VDD.n7904 4.61078
R23774 VDD.n7908 VDD.n7907 4.61078
R23775 VDD.n8045 VDD.n8042 4.61078
R23776 VDD.n8040 VDD.n8037 4.61078
R23777 VDD.n8035 VDD.n8032 4.61078
R23778 VDD.n8030 VDD.n8028 4.61078
R23779 VDD.n8026 VDD.n8023 4.61078
R23780 VDD.n8021 VDD.n8018 4.61078
R23781 VDD.n6803 VDD.n6802 4.61078
R23782 VDD.n7940 VDD.n7937 4.60951
R23783 VDD.n7941 VDD.n7940 4.60951
R23784 VDD.n7935 VDD.n7932 4.60951
R23785 VDD.n7936 VDD.n7935 4.60951
R23786 VDD.n7930 VDD.n7927 4.60951
R23787 VDD.n7931 VDD.n7930 4.60951
R23788 VDD.n7925 VDD.n7923 4.60951
R23789 VDD.n7926 VDD.n7925 4.60951
R23790 VDD.n7921 VDD.n7918 4.60951
R23791 VDD.n7922 VDD.n7921 4.60951
R23792 VDD.n7916 VDD.n7913 4.60951
R23793 VDD.n7917 VDD.n7916 4.60951
R23794 VDD.n6753 VDD.n6752 4.60825
R23795 VDD.n6998 VDD.n6997 4.60825
R23796 VDD.n6993 VDD.n6992 4.60825
R23797 VDD.n6988 VDD.n6987 4.60825
R23798 VDD.n6983 VDD.n6982 4.60825
R23799 VDD.n6901 VDD.n6900 4.60825
R23800 VDD.n6896 VDD.n6895 4.60825
R23801 VDD.n6891 VDD.n6890 4.60825
R23802 VDD.n6950 VDD.n6949 4.60825
R23803 VDD.n6945 VDD.n6944 4.60825
R23804 VDD.n6940 VDD.n6939 4.60825
R23805 VDD.n6935 VDD.n6934 4.60825
R23806 VDD.n6920 VDD.n6919 4.60825
R23807 VDD.n6915 VDD.n6914 4.60825
R23808 VDD.n6910 VDD.n6909 4.60825
R23809 VDD.n6524 VDD.n6523 4.60825
R23810 VDD.n6527 VDD.n6526 4.60825
R23811 VDD.n6530 VDD.n6529 4.60825
R23812 VDD.n6533 VDD.n6532 4.60825
R23813 VDD.n6434 VDD.n6433 4.60825
R23814 VDD.n6429 VDD.n6428 4.60825
R23815 VDD.n6424 VDD.n6423 4.60825
R23816 VDD.n6484 VDD.n6447 4.60825
R23817 VDD.n6487 VDD.n6486 4.60825
R23818 VDD.n6490 VDD.n6489 4.60825
R23819 VDD.n6493 VDD.n6492 4.60825
R23820 VDD.n6471 VDD.n6470 4.60825
R23821 VDD.n6466 VDD.n6465 4.60825
R23822 VDD.n6461 VDD.n6460 4.60825
R23823 VDD.n6066 VDD.n6065 4.60825
R23824 VDD.n6109 VDD.n6108 4.60825
R23825 VDD.n7892 VDD.n7891 4.60825
R23826 VDD.n7895 VDD.n7894 4.60825
R23827 VDD.n7898 VDD.n7897 4.60825
R23828 VDD.n7901 VDD.n7900 4.60825
R23829 VDD.n7904 VDD.n7903 4.60825
R23830 VDD.n7907 VDD.n7906 4.60825
R23831 VDD.n8046 VDD.n8045 4.60825
R23832 VDD.n8041 VDD.n8040 4.60825
R23833 VDD.n8036 VDD.n8035 4.60825
R23834 VDD.n8031 VDD.n8030 4.60825
R23835 VDD.n8027 VDD.n8026 4.60825
R23836 VDD.n8022 VDD.n8021 4.60825
R23837 VDD.n6802 VDD.n6801 4.60825
R23838 VDD.n6745 VDD.n6744 4.60191
R23839 VDD.n6757 VDD.n6756 4.60191
R23840 VDD.n6072 VDD.n6071 4.60191
R23841 VDD.n6060 VDD.n6041 4.60191
R23842 VDD.n6115 VDD.n6114 4.60191
R23843 VDD.n6103 VDD.n6101 4.60191
R23844 VDD.n6739 VDD.n6738 4.60191
R23845 VDD.n6806 VDD.n6805 4.60191
R23846 VDD.n8644 VDD.n8643 4.57315
R23847 VDD.n8703 VDD.n8702 4.57315
R23848 VDD.n1813 VDD.n1812 4.57315
R23849 VDD.n1869 VDD.n1868 4.57315
R23850 VDD.n5517 VDD.n5516 4.57315
R23851 VDD.n1961 VDD.n1960 4.57315
R23852 VDD.n2043 VDD.n2042 4.57315
R23853 VDD.n8753 VDD.n8752 4.57315
R23854 VDD.n8896 VDD.n8895 4.57315
R23855 VDD.n9069 VDD.n9068 4.57315
R23856 VDD.n8643 VDD.n8639 4.56231
R23857 VDD.n8702 VDD.n8698 4.56231
R23858 VDD.n1812 VDD.n1780 4.56231
R23859 VDD.n1868 VDD.n1842 4.56231
R23860 VDD.n5516 VDD.n1907 4.56231
R23861 VDD.n1960 VDD.n1934 4.56231
R23862 VDD.n2042 VDD.n2007 4.56231
R23863 VDD.n8752 VDD.n8748 4.56231
R23864 VDD.n8895 VDD.n8891 4.56231
R23865 VDD.n9068 VDD.n9064 4.56231
R23866 VDD.n6156 VDD.n6155 4.50663
R23867 VDD.n6099 VDD.n6098 4.50663
R23868 VDD.n6843 VDD.n6841 4.50663
R23869 VDD.n6793 VDD.n6728 4.50663
R23870 VDD.n59 VDD.n58 4.5005
R23871 VDD.n68 VDD.n63 4.5005
R23872 VDD.n148 VDD.n147 4.5005
R23873 VDD.n157 VDD.n152 4.5005
R23874 VDD.n5763 VDD.n5762 4.5005
R23875 VDD.n5758 VDD.n5757 4.5005
R23876 VDD.n5830 VDD.n5829 4.5005
R23877 VDD.n5825 VDD.n5824 4.5005
R23878 VDD.n5647 VDD.n5646 4.5005
R23879 VDD.n5642 VDD.n5641 4.5005
R23880 VDD.n5565 VDD.n5564 4.5005
R23881 VDD.n5560 VDD.n5559 4.5005
R23882 VDD.n8151 VDD.n8150 4.5005
R23883 VDD.n8146 VDD.n8145 4.5005
R23884 VDD.n6889 VDD.n6885 4.5005
R23885 VDD.n6894 VDD.n6884 4.5005
R23886 VDD.n6899 VDD.n6883 4.5005
R23887 VDD.n6981 VDD.n6882 4.5005
R23888 VDD.n6986 VDD.n6881 4.5005
R23889 VDD.n6991 VDD.n6880 4.5005
R23890 VDD.n6996 VDD.n6879 4.5005
R23891 VDD.n6908 VDD.n6904 4.5005
R23892 VDD.n6913 VDD.n6903 4.5005
R23893 VDD.n6918 VDD.n6902 4.5005
R23894 VDD.n6933 VDD.n6930 4.5005
R23895 VDD.n6938 VDD.n6929 4.5005
R23896 VDD.n6943 VDD.n6928 4.5005
R23897 VDD.n6948 VDD.n6927 4.5005
R23898 VDD.n5983 VDD.n5914 4.5005
R23899 VDD.n6322 VDD.n5914 4.5005
R23900 VDD.n6323 VDD.n6322 4.5005
R23901 VDD.n6324 VDD.n5914 4.5005
R23902 VDD.n5981 VDD.n5914 4.5005
R23903 VDD.n6323 VDD.n5981 4.5005
R23904 VDD.n6324 VDD.n6323 4.5005
R23905 VDD.n6422 VDD.n6418 4.5005
R23906 VDD.n6427 VDD.n6417 4.5005
R23907 VDD.n6432 VDD.n6416 4.5005
R23908 VDD.n6437 VDD.n6435 4.5005
R23909 VDD.n6440 VDD.n6438 4.5005
R23910 VDD.n6443 VDD.n6441 4.5005
R23911 VDD.n6446 VDD.n6444 4.5005
R23912 VDD.n6459 VDD.n6455 4.5005
R23913 VDD.n6464 VDD.n6454 4.5005
R23914 VDD.n6469 VDD.n6453 4.5005
R23915 VDD.n6474 VDD.n6472 4.5005
R23916 VDD.n6477 VDD.n6475 4.5005
R23917 VDD.n6480 VDD.n6478 4.5005
R23918 VDD.n6483 VDD.n6481 4.5005
R23919 VDD.n6102 VDD.n6040 4.5005
R23920 VDD.n6107 VDD.n6039 4.5005
R23921 VDD.n6111 VDD.n6110 4.5005
R23922 VDD.n6059 VDD.n6058 4.5005
R23923 VDD.n6064 VDD.n6057 4.5005
R23924 VDD.n6068 VDD.n6067 4.5005
R23925 VDD.n6173 VDD.n6015 4.5005
R23926 VDD.n6179 VDD.n6015 4.5005
R23927 VDD.n6179 VDD.n6012 4.5005
R23928 VDD.n6179 VDD.n6011 4.5005
R23929 VDD.n6179 VDD.n6178 4.5005
R23930 VDD.n6178 VDD.n6177 4.5005
R23931 VDD.n6177 VDD.n6011 4.5005
R23932 VDD.n7915 VDD.n7860 4.5005
R23933 VDD.n7920 VDD.n7859 4.5005
R23934 VDD.n7924 VDD.n7858 4.5005
R23935 VDD.n7929 VDD.n7857 4.5005
R23936 VDD.n7934 VDD.n7856 4.5005
R23937 VDD.n7939 VDD.n7855 4.5005
R23938 VDD.n7867 VDD.n7865 4.5005
R23939 VDD.n7871 VDD.n7869 4.5005
R23940 VDD.n7874 VDD.n7873 4.5005
R23941 VDD.n7877 VDD.n7875 4.5005
R23942 VDD.n7881 VDD.n7879 4.5005
R23943 VDD.n7885 VDD.n7883 4.5005
R23944 VDD.n8020 VDD.n2155 4.5005
R23945 VDD.n8025 VDD.n2154 4.5005
R23946 VDD.n8029 VDD.n2153 4.5005
R23947 VDD.n8034 VDD.n2152 4.5005
R23948 VDD.n8039 VDD.n2151 4.5005
R23949 VDD.n8044 VDD.n2150 4.5005
R23950 VDD.n6730 VDD.n6729 4.5005
R23951 VDD.n6733 VDD.n6731 4.5005
R23952 VDD.n6735 VDD.n6734 4.5005
R23953 VDD.n6748 VDD.n6747 4.5005
R23954 VDD.n6751 VDD.n6749 4.5005
R23955 VDD.n6741 VDD.n6740 4.5005
R23956 VDD.n8161 VDD.n8160 4.5005
R23957 VDD.n8160 VDD.n8142 4.5005
R23958 VDD.n8143 VDD.n8140 4.5005
R23959 VDD.n8143 VDD.n2089 4.5005
R23960 VDD.n5575 VDD.n5574 4.5005
R23961 VDD.n5574 VDD.n5555 4.5005
R23962 VDD.n5557 VDD.n5553 4.5005
R23963 VDD.n5557 VDD.n5556 4.5005
R23964 VDD.n10817 VDD.n2002 4.5005
R23965 VDD.n8092 VDD.n8091 4.5005
R23966 VDD.n8092 VDD.n2109 4.5005
R23967 VDD.n8095 VDD.n2109 4.5005
R23968 VDD.n8095 VDD.n8094 4.5005
R23969 VDD.n8094 VDD.n2105 4.5005
R23970 VDD.n2110 VDD.n2105 4.5005
R23971 VDD.n8091 VDD.n2105 4.5005
R23972 VDD.n10819 VDD.n2004 4.5005
R23973 VDD.n2004 VDD.n1996 4.5005
R23974 VDD.n2004 VDD.n2001 4.5005
R23975 VDD.n10820 VDD.n2001 4.5005
R23976 VDD.n10820 VDD.n1997 4.5005
R23977 VDD.n10820 VDD.n2002 4.5005
R23978 VDD.n10820 VDD.n1996 4.5005
R23979 VDD.n10820 VDD.n10819 4.5005
R23980 VDD.n5657 VDD.n5656 4.5005
R23981 VDD.n5656 VDD.n5546 4.5005
R23982 VDD.n5639 VDD.n5638 4.5005
R23983 VDD.n5639 VDD.n5544 4.5005
R23984 VDD.n5907 VDD.n5540 4.5005
R23985 VDD.n5908 VDD.n5907 4.5005
R23986 VDD.n5534 VDD.n5533 4.5005
R23987 VDD.n5533 VDD.n5503 4.5005
R23988 VDD.n5883 VDD.n1919 4.5005
R23989 VDD.n5890 VDD.n5883 4.5005
R23990 VDD.n5531 VDD.n5503 4.5005
R23991 VDD.n5890 VDD.n5881 4.5005
R23992 VDD.n5904 VDD.n5902 4.5005
R23993 VDD.n5535 VDD.n5534 4.5005
R23994 VDD.n5529 VDD.n5489 4.5005
R23995 VDD.n5535 VDD.n5529 4.5005
R23996 VDD.n5902 VDD.n5540 4.5005
R23997 VDD.n5908 VDD.n5902 4.5005
R23998 VDD.n5890 VDD.n5885 4.5005
R23999 VDD.n5890 VDD.n5880 4.5005
R24000 VDD.n5885 VDD.n1919 4.5005
R24001 VDD.n5880 VDD.n1919 4.5005
R24002 VDD.n5503 VDD.n5489 4.5005
R24003 VDD.n5840 VDD.n5839 4.5005
R24004 VDD.n5839 VDD.n5821 4.5005
R24005 VDD.n5822 VDD.n5819 4.5005
R24006 VDD.n5822 VDD.n5680 4.5005
R24007 VDD.n5773 VDD.n5772 4.5005
R24008 VDD.n5772 VDD.n5754 4.5005
R24009 VDD.n5755 VDD.n5752 4.5005
R24010 VDD.n5755 VDD.n5704 4.5005
R24011 VDD.n11048 VDD.n11047 4.5005
R24012 VDD.n11047 VDD.n11046 4.5005
R24013 VDD.n11046 VDD.n675 4.5005
R24014 VDD.n11046 VDD.n1764 4.5005
R24015 VDD.n11046 VDD.n674 4.5005
R24016 VDD.n11046 VDD.n11045 4.5005
R24017 VDD.n11045 VDD.n11044 4.5005
R24018 VDD.n11044 VDD.n674 4.5005
R24019 VDD.n11044 VDD.n1764 4.5005
R24020 VDD.n11130 VDD.n636 4.5005
R24021 VDD.n640 VDD.n636 4.5005
R24022 VDD.n11129 VDD.n640 4.5005
R24023 VDD.n640 VDD.n635 4.5005
R24024 VDD.n11127 VDD.n634 4.5005
R24025 VDD.n11130 VDD.n635 4.5005
R24026 VDD.n11130 VDD.n637 4.5005
R24027 VDD.n11130 VDD.n634 4.5005
R24028 VDD.n11130 VDD.n11129 4.5005
R24029 VDD.n5220 VDD.n4593 4.5005
R24030 VDD.n5220 VDD.n4594 4.5005
R24031 VDD.n5220 VDD.n5219 4.5005
R24032 VDD.n5204 VDD.n2408 4.5005
R24033 VDD.n4599 VDD.n2408 4.5005
R24034 VDD.n4591 VDD.n2425 4.5005
R24035 VDD.n4592 VDD.n4591 4.5005
R24036 VDD.n5219 VDD.n5218 4.5005
R24037 VDD.n9103 VDD.n9102 4.5005
R24038 VDD.n9112 VDD.n9107 4.5005
R24039 VDD.n8816 VDD.n8815 4.5005
R24040 VDD.n8825 VDD.n8820 4.5005
R24041 VDD.n8956 VDD.n8955 4.5005
R24042 VDD.n8965 VDD.n8960 4.5005
R24043 VDD.n9003 VDD.n9002 4.5005
R24044 VDD.n9004 VDD.n9003 4.5005
R24045 VDD.n9001 VDD.n9000 4.5005
R24046 VDD.n9000 VDD.n8953 4.5005
R24047 VDD.n8832 VDD.n8831 4.5005
R24048 VDD.n8833 VDD.n8832 4.5005
R24049 VDD.n8813 VDD.n8525 4.5005
R24050 VDD.n8813 VDD.n8812 4.5005
R24051 VDD.n9100 VDD.n9090 4.5005
R24052 VDD.n9100 VDD.n9099 4.5005
R24053 VDD.n9120 VDD.n9119 4.5005
R24054 VDD.n9119 VDD.n9118 4.5005
R24055 VDD.n9200 VDD.n9184 4.5005
R24056 VDD.n9184 VDD.n8458 4.5005
R24057 VDD.n12448 VDD.n194 4.5005
R24058 VDD.n12448 VDD.n12447 4.5005
R24059 VDD.n164 VDD.n163 4.5005
R24060 VDD.n165 VDD.n164 4.5005
R24061 VDD.n145 VDD.n135 4.5005
R24062 VDD.n145 VDD.n144 4.5005
R24063 VDD.n75 VDD.n74 4.5005
R24064 VDD.n76 VDD.n75 4.5005
R24065 VDD.n56 VDD.n46 4.5005
R24066 VDD.n56 VDD.n55 4.5005
R24067 VDD.n12583 VDD.n12580 4.5005
R24068 VDD.n12584 VDD.n12583 4.5005
R24069 VDD.n12581 VDD.n12580 4.5005
R24070 VDD.n12581 VDD.n12561 4.5005
R24071 VDD.n12585 VDD.n12561 4.5005
R24072 VDD.n12585 VDD.n12559 4.5005
R24073 VDD.n12585 VDD.n12584 4.5005
R24074 VDD.n12626 VDD.n8 4.5005
R24075 VDD.n12628 VDD.n9 4.5005
R24076 VDD.n12630 VDD.n12628 4.5005
R24077 VDD.n12630 VDD.n12623 4.5005
R24078 VDD.n12630 VDD.n8 4.5005
R24079 VDD.n12631 VDD.n9 4.5005
R24080 VDD.n12629 VDD.n9 4.5005
R24081 VDD.n12631 VDD.n12630 4.5005
R24082 VDD.n12630 VDD.n12629 4.5005
R24083 VDD.n1757 VDD.n680 4.5005
R24084 VDD.n1759 VDD.n680 4.5005
R24085 VDD.n1755 VDD.n680 4.5005
R24086 VDD.n1757 VDD.n678 4.5005
R24087 VDD.n1759 VDD.n678 4.5005
R24088 VDD.n678 VDD.n677 4.5005
R24089 VDD.n1755 VDD.n678 4.5005
R24090 VDD.n1756 VDD.n677 4.5005
R24091 VDD.n1756 VDD.n1755 4.5005
R24092 VDD.n1002 VDD.n1001 4.5005
R24093 VDD.n1003 VDD.n1002 4.5005
R24094 VDD.n956 VDD.n954 4.5005
R24095 VDD.n956 VDD.n953 4.5005
R24096 VDD.n1001 VDD.n956 4.5005
R24097 VDD.n1003 VDD.n956 4.5005
R24098 VDD.n1004 VDD.n954 4.5005
R24099 VDD.n1004 VDD.n953 4.5005
R24100 VDD.n1004 VDD.n1003 4.5005
R24101 VDD.n12641 VDD.n1 4.5005
R24102 VDD.n12642 VDD.n5 4.5005
R24103 VDD.n12642 VDD.n3 4.5005
R24104 VDD.n12642 VDD.n12636 4.5005
R24105 VDD.n12642 VDD.n12641 4.5005
R24106 VDD.n12640 VDD.n5 4.5005
R24107 VDD.n12640 VDD.n3 4.5005
R24108 VDD.n12640 VDD.n12636 4.5005
R24109 VDD.n12641 VDD.n12640 4.5005
R24110 VDD.n6092 VDD.n6041 4.32507
R24111 VDD.n6758 VDD.n6757 4.32507
R24112 VDD.n823 VDD.t2747 4.07396
R24113 VDD.n6952 VDD.t200 4.06712
R24114 VDD.n6925 VDD.t250 4.06712
R24115 VDD.n7010 VDD.t289 4.06712
R24116 VDD.n7003 VDD.t115 4.06712
R24117 VDD.n6502 VDD.t4945 4.06712
R24118 VDD.n6451 VDD.t4929 4.06712
R24119 VDD.n6542 VDD.t4868 4.06712
R24120 VDD.n6540 VDD.t4846 4.06712
R24121 VDD.n1477 VDD.t3030 4.05637
R24122 VDD.n1611 VDD.t4124 4.05637
R24123 VDD.n1609 VDD.t2801 4.05637
R24124 VDD.n1478 VDD.t1531 4.05637
R24125 VDD.n1117 VDD.t1629 4.05408
R24126 VDD.n1116 VDD.t4566 4.05408
R24127 VDD.n1182 VDD.t1989 4.05408
R24128 VDD.n1115 VDD.t1761 4.05408
R24129 VDD.n1114 VDD.t4730 4.05408
R24130 VDD.n1138 VDD.t1218 4.05408
R24131 VDD.n1137 VDD.t1685 4.05408
R24132 VDD.n1169 VDD.t3004 4.05408
R24133 VDD.n1136 VDD.t4140 4.05408
R24134 VDD.n1135 VDD.t1479 4.05408
R24135 VDD.n1312 VDD.t2378 4.05408
R24136 VDD.n1313 VDD.t3848 4.05408
R24137 VDD.n757 VDD.t2745 4.05408
R24138 VDD.n756 VDD.t1091 4.05408
R24139 VDD.n755 VDD.t2710 4.05408
R24140 VDD.n754 VDD.t3118 4.05408
R24141 VDD.n1280 VDD.t883 4.05408
R24142 VDD.n1308 VDD.t592 4.05408
R24143 VDD.n1278 VDD.t866 4.05408
R24144 VDD.n1279 VDD.t3798 4.05408
R24145 VDD.n1311 VDD.t3573 4.05408
R24146 VDD.n1080 VDD.t3498 4.05408
R24147 VDD.n1081 VDD.t891 4.05408
R24148 VDD.n1359 VDD.t3478 4.05408
R24149 VDD.n1282 VDD.t3668 4.05408
R24150 VDD.n1281 VDD.t3812 4.05408
R24151 VDD.n878 VDD.t3286 4.05408
R24152 VDD.n1076 VDD.t582 4.05408
R24153 VDD.n876 VDD.t2027 4.05408
R24154 VDD.n877 VDD.t4592 4.05408
R24155 VDD.n1079 VDD.t1995 4.05408
R24156 VDD.n1244 VDD.t4598 4.05408
R24157 VDD.n1245 VDD.t3434 4.05408
R24158 VDD.n765 VDD.t3542 4.05408
R24159 VDD.n766 VDD.t3342 4.05408
R24160 VDD.n767 VDD.t2139 4.05408
R24161 VDD.n768 VDD.t2936 4.05408
R24162 VDD.n805 VDD.t2113 4.05408
R24163 VDD.n1497 VDD.t1310 4.05408
R24164 VDD.n1498 VDD.t3220 4.05408
R24165 VDD.n1499 VDD.t4696 4.05408
R24166 VDD.n1601 VDD.t3522 4.05408
R24167 VDD.n1502 VDD.t1942 4.05408
R24168 VDD.n1503 VDD.t3506 4.05408
R24169 VDD.n1504 VDD.t3924 4.05408
R24170 VDD.n805 VDD.t2408 4.05408
R24171 VDD.n1497 VDD.t1523 4.05408
R24172 VDD.n1498 VDD.t3395 4.05408
R24173 VDD.n1499 VDD.t785 4.05408
R24174 VDD.n1601 VDD.t3727 4.05408
R24175 VDD.n1502 VDD.t2188 4.05408
R24176 VDD.n1503 VDD.t3707 4.05408
R24177 VDD.n1504 VDD.t4150 4.05408
R24178 VDD.n1109 VDD.t3194 4.05408
R24179 VDD.n1240 VDD.t4674 4.05408
R24180 VDD.n1107 VDD.t1705 4.05408
R24181 VDD.n1108 VDD.t1845 4.05408
R24182 VDD.n1243 VDD.t3419 4.05408
R24183 VDD.n1113 VDD.t720 4.05408
R24184 VDD.n1112 VDD.t3658 4.05408
R24185 VDD.n1212 VDD.t3484 4.05408
R24186 VDD.n1111 VDD.t4670 4.05408
R24187 VDD.n1110 VDD.t2479 4.05408
R24188 VDD.n727 VDD.t3106 4.05408
R24189 VDD.n1396 VDD.t3662 4.05408
R24190 VDD.n1395 VDD.t4116 4.05408
R24191 VDD.n1394 VDD.t1449 4.05408
R24192 VDD.n1391 VDD.t2968 4.05408
R24193 VDD.n1393 VDD.t1297 4.05408
R24194 VDD.n1404 VDD.t2954 4.05408
R24195 VDD.n1405 VDD.t3312 4.05408
R24196 VDD.n822 VDD.t3932 4.05408
R24197 VDD.n1446 VDD.t4344 4.05408
R24198 VDD.n819 VDD.t1699 4.05408
R24199 VDD.n820 VDD.t4314 4.05408
R24200 VDD.n817 VDD.t4510 4.05408
R24201 VDD.n816 VDD.t4660 4.05408
R24202 VDD.n815 VDD.t2422 4.05408
R24203 VDD.n812 VDD.t1546 4.05408
R24204 VDD.n811 VDD.t1695 4.05408
R24205 VDD.n809 VDD.t1471 4.05408
R24206 VDD.n810 VDD.t1681 4.05408
R24207 VDD.n807 VDD.t4654 4.05408
R24208 VDD.n806 VDD.t4408 4.05408
R24209 VDD.n727 VDD.t3296 4.05408
R24210 VDD.n1396 VDD.t3890 4.05408
R24211 VDD.n1395 VDD.t4312 4.05408
R24212 VDD.n1394 VDD.t1675 4.05408
R24213 VDD.n1391 VDD.t3158 4.05408
R24214 VDD.n1393 VDD.t1510 4.05408
R24215 VDD.n1404 VDD.t3146 4.05408
R24216 VDD.n1405 VDD.t3510 4.05408
R24217 VDD.n822 VDD.t4156 4.05408
R24218 VDD.n1446 VDD.t4528 4.05408
R24219 VDD.n819 VDD.t1933 4.05408
R24220 VDD.n820 VDD.t4512 4.05408
R24221 VDD.n817 VDD.t4738 4.05408
R24222 VDD.n816 VDD.t742 4.05408
R24223 VDD.n815 VDD.t2659 4.05408
R24224 VDD.n812 VDD.t1771 4.05408
R24225 VDD.n811 VDD.t1929 4.05408
R24226 VDD.n809 VDD.t1683 4.05408
R24227 VDD.n810 VDD.t1908 4.05408
R24228 VDD.n807 VDD.t738 4.05408
R24229 VDD.n806 VDD.t4638 4.05408
R24230 VDD.n900 VDD.t3258 4.05408
R24231 VDD.n899 VDD.t1527 4.05408
R24232 VDD.n1065 VDD.t1746 4.05408
R24233 VDD.n898 VDD.t1985 4.05408
R24234 VDD.n897 VDD.t1724 4.05408
R24235 VDD.n904 VDD.t1648 4.05408
R24236 VDD.n903 VDD.t2826 4.05408
R24237 VDD.n910 VDD.t4378 4.05408
R24238 VDD.n902 VDD.t4582 4.05408
R24239 VDD.n901 VDD.t4462 4.05408
R24240 VDD.n943 VDD.t2621 4.05408
R24241 VDD.n944 VDD.t3599 4.05408
R24242 VDD.n693 VDD.t1106 4.05408
R24243 VDD.n695 VDD.t1288 4.05408
R24244 VDD.n697 VDD.t1153 4.05408
R24245 VDD.n943 VDD.t2830 4.05408
R24246 VDD.n944 VDD.t3816 4.05408
R24247 VDD.n693 VDD.t1290 4.05408
R24248 VDD.n695 VDD.t1505 4.05408
R24249 VDD.n697 VDD.t1370 4.05408
R24250 VDD.n698 VDD.t1574 4.05408
R24251 VDD.n718 VDD.t2251 4.05408
R24252 VDD.n717 VDD.t4068 4.05408
R24253 VDD.n716 VDD.t2508 4.05408
R24254 VDD.n713 VDD.t2720 4.05408
R24255 VDD.n715 VDD.t2940 4.05408
R24256 VDD.n726 VDD.t2700 4.05408
R24257 VDD.n698 VDD.t1784 4.05408
R24258 VDD.n718 VDD.t2536 4.05408
R24259 VDD.n717 VDD.t4286 4.05408
R24260 VDD.n716 VDD.t2722 4.05408
R24261 VDD.n713 VDD.t2944 4.05408
R24262 VDD.n715 VDD.t3136 4.05408
R24263 VDD.n726 VDD.t2912 4.05408
R24264 VDD.n683 VDD.t3050 4.05408
R24265 VDD.n684 VDD.t740 4.05408
R24266 VDD.n1745 VDD.t4640 4.05408
R24267 VDD.n1158 VDD.t1679 4.05408
R24268 VDD.n1157 VDD.t4198 4.05408
R24269 VDD.n57 VDD.t534 4.00905
R24270 VDD.n146 VDD.t4765 4.00905
R24271 VDD.n9101 VDD.t4747 4.00905
R24272 VDD.n8814 VDD.t10 4.00905
R24273 VDD.n8954 VDD.t4805 4.00905
R24274 VDD.n5756 VDD.t367 4.00848
R24275 VDD.n5823 VDD.t4797 4.00848
R24276 VDD.n5640 VDD.t4750 4.00848
R24277 VDD.n5558 VDD.t516 4.00848
R24278 VDD.n8144 VDD.t305 4.00848
R24279 VDD.n60 VDD.t539 4.00673
R24280 VDD.n149 VDD.t4763 4.00673
R24281 VDD.n9104 VDD.t4757 4.00673
R24282 VDD.n8817 VDD.t5 4.00673
R24283 VDD.n8957 VDD.t4801 4.00673
R24284 VDD.n5759 VDD.t302 4.00554
R24285 VDD.n5826 VDD.t4796 4.00554
R24286 VDD.n5643 VDD.t4755 4.00554
R24287 VDD.n5561 VDD.t519 4.00554
R24288 VDD.n8147 VDD.t303 4.00554
R24289 VDD.n7012 VDD.n7011 3.96014
R24290 VDD.n6953 VDD.n6951 3.96014
R24291 VDD.n6543 VDD.n5289 3.96014
R24292 VDD.n6504 VDD.n6503 3.96014
R24293 VDD.n6952 VDD.t62 3.86107
R24294 VDD.n6925 VDD.t127 3.86107
R24295 VDD.n7010 VDD.t237 3.86107
R24296 VDD.n7003 VDD.t282 3.86107
R24297 VDD.n6502 VDD.t4855 3.86107
R24298 VDD.n6451 VDD.t4838 3.86107
R24299 VDD.n6542 VDD.t4916 3.86107
R24300 VDD.n6540 VDD.t4901 3.86107
R24301 VDD.n8641 VDD.t540 3.8555
R24302 VDD.n8700 VDD.t4786 3.8555
R24303 VDD.n1810 VDD.t416 3.8555
R24304 VDD.n1866 VDD.t4769 3.8555
R24305 VDD.n5514 VDD.t4785 3.8555
R24306 VDD.n1958 VDD.t510 3.8555
R24307 VDD.n2040 VDD.t505 3.8555
R24308 VDD.n8750 VDD.t299 3.8555
R24309 VDD.n8893 VDD.t523 3.8555
R24310 VDD.n9066 VDD.t4775 3.8555
R24311 VDD.n8640 VDD.t541 3.85313
R24312 VDD.n8699 VDD.t4788 3.85313
R24313 VDD.n1809 VDD.t417 3.85313
R24314 VDD.n1865 VDD.t4770 3.85313
R24315 VDD.n5513 VDD.t4784 3.85313
R24316 VDD.n1957 VDD.t508 3.85313
R24317 VDD.n2039 VDD.t507 3.85313
R24318 VDD.n8749 VDD.t298 3.85313
R24319 VDD.n8892 VDD.t520 3.85313
R24320 VDD.n9065 VDD.t4774 3.85313
R24321 VDD.n6741 VDD.t153 3.84568
R24322 VDD.n6748 VDD.t171 3.84568
R24323 VDD.n6068 VDD.t4825 3.84568
R24324 VDD.n6059 VDD.t4946 3.84568
R24325 VDD.n6111 VDD.t4877 3.84568
R24326 VDD.n6102 VDD.t4817 3.84568
R24327 VDD.n6735 VDD.t80 3.84568
R24328 VDD.n6730 VDD.t103 3.84568
R24329 VDD.n6021 VDD.n6020 3.84528
R24330 VDD.n6155 VDD.n6154 3.84528
R24331 VDD.n6094 VDD.n6093 3.84528
R24332 VDD.n6098 VDD.n6097 3.84528
R24333 VDD.n6846 VDD.n6845 3.84528
R24334 VDD.n6843 VDD.n6842 3.84528
R24335 VDD.n6796 VDD.n6795 3.84528
R24336 VDD.n6793 VDD.n6792 3.84528
R24337 VDD.n7901 VDD.t31 3.84449
R24338 VDD.n2381 VDD.n2379 3.79678
R24339 VDD.n7019 VDD.n7017 3.79678
R24340 VDD.n6964 VDD.n6962 3.79678
R24341 VDD.n6972 VDD.n6970 3.79678
R24342 VDD.n5294 VDD.n5292 3.79678
R24343 VDD.n6557 VDD.n6555 3.79678
R24344 VDD.n6509 VDD.n6507 3.79678
R24345 VDD.n6518 VDD.n6516 3.79678
R24346 VDD.n6129 VDD.n6125 3.79678
R24347 VDD.n6144 VDD.n6140 3.79678
R24348 VDD.n6087 VDD.n6083 3.79678
R24349 VDD.n6052 VDD.n6048 3.79678
R24350 VDD.n6835 VDD.n6831 3.79678
R24351 VDD.n6818 VDD.n6814 3.79678
R24352 VDD.n6770 VDD.n6766 3.79678
R24353 VDD.n6785 VDD.n6781 3.79678
R24354 VDD.n5756 VDD.t326 3.78097
R24355 VDD.n5823 VDD.t4795 3.78097
R24356 VDD.n5640 VDD.t4749 3.78097
R24357 VDD.n5558 VDD.t515 3.78097
R24358 VDD.n8144 VDD.t339 3.78097
R24359 VDD.n5764 VDD.t368 3.78097
R24360 VDD.n5831 VDD.t4794 3.78097
R24361 VDD.n5648 VDD.t4748 3.78097
R24362 VDD.n5566 VDD.t514 3.78097
R24363 VDD.n8152 VDD.t366 3.78097
R24364 VDD.n57 VDD.t531 3.7804
R24365 VDD.n64 VDD.t532 3.7804
R24366 VDD.n146 VDD.t4759 3.7804
R24367 VDD.n153 VDD.t4761 3.7804
R24368 VDD.n9101 VDD.t4756 3.7804
R24369 VDD.n9108 VDD.t4746 3.7804
R24370 VDD.n8814 VDD.t7 3.7804
R24371 VDD.n8821 VDD.t8 3.7804
R24372 VDD.n8954 VDD.t4802 3.7804
R24373 VDD.n8961 VDD.t4803 3.7804
R24374 VDD.n59 VDD.t536 3.77818
R24375 VDD.n68 VDD.t537 3.77818
R24376 VDD.n148 VDD.t4758 3.77818
R24377 VDD.n157 VDD.t4760 3.77818
R24378 VDD.n5763 VDD.t419 3.77818
R24379 VDD.n5758 VDD.t418 3.77818
R24380 VDD.n5830 VDD.t4792 3.77818
R24381 VDD.n5825 VDD.t4793 3.77818
R24382 VDD.n5647 VDD.t4753 3.77818
R24383 VDD.n5642 VDD.t4754 3.77818
R24384 VDD.n5565 VDD.t517 3.77818
R24385 VDD.n5560 VDD.t518 3.77818
R24386 VDD.n8151 VDD.t14 3.77818
R24387 VDD.n8146 VDD.t365 3.77818
R24388 VDD.n9103 VDD.t555 3.77818
R24389 VDD.n9112 VDD.t553 3.77818
R24390 VDD.n8816 VDD.t11 3.77818
R24391 VDD.n8825 VDD.t2 3.77818
R24392 VDD.n8956 VDD.t4806 3.77818
R24393 VDD.n8965 VDD.t4807 3.77818
R24394 VDD.n6101 VDD.n6100 3.74038
R24395 VDD.n6807 VDD.n6806 3.74038
R24396 VDD.n6149 VDD.n6133 3.73034
R24397 VDD.n6079 VDD.n6075 3.73034
R24398 VDD.n6827 VDD.n6823 3.73034
R24399 VDD.n6790 VDD.n6774 3.73034
R24400 VDD.n7995 VDD.t26 3.7109
R24401 VDD.n980 VDD.n978 3.70005
R24402 VDD.n1038 VDD.n1037 3.70005
R24403 VDD.n1041 VDD.n1040 3.70005
R24404 VDD.n1102 VDD.n1101 3.70005
R24405 VDD.n1624 VDD.n1623 3.70005
R24406 VDD.n1090 VDD.n1089 3.70005
R24407 VDD.n1423 VDD.n1422 3.70005
R24408 VDD.n857 VDD.n856 3.70005
R24409 VDD.n1674 VDD.n746 3.70005
R24410 VDD.n1680 VDD.n743 3.70005
R24411 VDD.n1686 VDD.n740 3.70005
R24412 VDD.n1693 VDD.n737 3.70005
R24413 VDD.n982 VDD.n981 3.6965
R24414 VDD.n1036 VDD.n1035 3.6965
R24415 VDD.n1043 VDD.n1042 3.6965
R24416 VDD.n1104 VDD.n1103 3.6965
R24417 VDD.n1622 VDD.n1621 3.6965
R24418 VDD.n1088 VDD.n1087 3.6965
R24419 VDD.n1421 VDD.n1420 3.6965
R24420 VDD.n855 VDD.n854 3.6965
R24421 VDD.n1676 VDD.n1675 3.6965
R24422 VDD.n1682 VDD.n1681 3.6965
R24423 VDD.n1688 VDD.n1687 3.6965
R24424 VDD.n1695 VDD.n1694 3.6965
R24425 VDD.n8640 VDD.t543 3.68497
R24426 VDD.n8699 VDD.t4787 3.68497
R24427 VDD.n1809 VDD.t295 3.68497
R24428 VDD.n1865 VDD.t4768 3.68497
R24429 VDD.n5513 VDD.t4782 3.68497
R24430 VDD.n1957 VDD.t511 3.68497
R24431 VDD.n2039 VDD.t506 3.68497
R24432 VDD.n8749 VDD.t300 3.68497
R24433 VDD.n8892 VDD.t522 3.68497
R24434 VDD.n9065 VDD.t4772 3.68497
R24435 VDD.n7874 VDD.t34 3.68344
R24436 VDD.n8641 VDD.t542 3.68261
R24437 VDD.n8700 VDD.t4789 3.68261
R24438 VDD.n1810 VDD.t294 3.68261
R24439 VDD.n1866 VDD.t4771 3.68261
R24440 VDD.n5514 VDD.t4783 3.68261
R24441 VDD.n1958 VDD.t509 3.68261
R24442 VDD.n2040 VDD.t504 3.68261
R24443 VDD.n8750 VDD.t297 3.68261
R24444 VDD.n8893 VDD.t521 3.68261
R24445 VDD.n9066 VDD.t4773 3.68261
R24446 VDD.n7954 VDD.n7953 3.65594
R24447 VDD.n7015 VDD.n7014 3.65581
R24448 VDD.n7017 VDD.n7016 3.65581
R24449 VDD.n7019 VDD.n7018 3.65581
R24450 VDD.n7021 VDD.n7020 3.65581
R24451 VDD.n2383 VDD.n2382 3.65581
R24452 VDD.n2381 VDD.n2380 3.65581
R24453 VDD.n2379 VDD.n2378 3.65581
R24454 VDD.n6968 VDD.n6967 3.65581
R24455 VDD.n6970 VDD.n6969 3.65581
R24456 VDD.n6972 VDD.n6971 3.65581
R24457 VDD.n6974 VDD.n6973 3.65581
R24458 VDD.n6966 VDD.n6965 3.65581
R24459 VDD.n6964 VDD.n6963 3.65581
R24460 VDD.n6962 VDD.n6961 3.65581
R24461 VDD.n6559 VDD.n6558 3.65581
R24462 VDD.n6557 VDD.n6556 3.65581
R24463 VDD.n6555 VDD.n6554 3.65581
R24464 VDD.n6553 VDD.n6552 3.65581
R24465 VDD.n5296 VDD.n5295 3.65581
R24466 VDD.n5294 VDD.n5293 3.65581
R24467 VDD.n5292 VDD.n5291 3.65581
R24468 VDD.n6520 VDD.n6519 3.65581
R24469 VDD.n6518 VDD.n6517 3.65581
R24470 VDD.n6516 VDD.n6515 3.65581
R24471 VDD.n6514 VDD.n6513 3.65581
R24472 VDD.n6511 VDD.n6510 3.65581
R24473 VDD.n6509 VDD.n6508 3.65581
R24474 VDD.n6507 VDD.n6506 3.65581
R24475 VDD.n7949 VDD.n7948 3.6512
R24476 VDD.n7958 VDD.n7957 3.6512
R24477 VDD.n7951 VDD.n7950 3.6512
R24478 VDD.n7956 VDD.n7955 3.6512
R24479 VDD.n7022 VDD.n7021 3.64443
R24480 VDD.n6975 VDD.n6974 3.64443
R24481 VDD.n6553 VDD.n6551 3.64443
R24482 VDD.n6514 VDD.n6512 3.64443
R24483 VDD.n8029 VDD.t169 3.6266
R24484 VDD.n8054 VDD.n8053 3.62041
R24485 VDD.n8056 VDD.n8055 3.62041
R24486 VDD.n8059 VDD.n8058 3.62041
R24487 VDD.n8061 VDD.n8060 3.62041
R24488 VDD.n8063 VDD.n8062 3.62041
R24489 VDD.n7924 VDD.t60 3.61594
R24490 VDD.n62 VDD.n61 3.54958
R24491 VDD.n151 VDD.n150 3.54958
R24492 VDD.n5761 VDD.n5760 3.54958
R24493 VDD.n5828 VDD.n5827 3.54958
R24494 VDD.n5645 VDD.n5644 3.54958
R24495 VDD.n5563 VDD.n5562 3.54958
R24496 VDD.n8149 VDD.n8148 3.54958
R24497 VDD.n9106 VDD.n9105 3.54958
R24498 VDD.n8819 VDD.n8818 3.54958
R24499 VDD.n8959 VDD.n8958 3.54958
R24500 VDD.n6892 VDD.n6891 3.524
R24501 VDD.n6989 VDD.n6988 3.524
R24502 VDD.n6911 VDD.n6910 3.524
R24503 VDD.n6941 VDD.n6940 3.524
R24504 VDD.n6425 VDD.n6424 3.524
R24505 VDD.n6529 VDD.n6528 3.524
R24506 VDD.n6462 VDD.n6461 3.524
R24507 VDD.n6489 VDD.n6488 3.524
R24508 VDD.n6979 VDD.n6978 3.506
R24509 VDD.n6931 VDD.n6921 3.506
R24510 VDD.n6535 VDD.n6534 3.506
R24511 VDD.n6495 VDD.n6494 3.506
R24512 VDD.n1441 VDD.t383 3.3982
R24513 VDD.n804 VDD.t382 3.3982
R24514 VDD.n803 VDD.t385 3.3982
R24515 VDD.n1479 VDD.t379 3.3982
R24516 VDD.n814 VDD.t310 3.3982
R24517 VDD.n751 VDD.t386 3.37007
R24518 VDD.n1506 VDD.t307 3.37007
R24519 VDD.n6326 VDD.n5912 3.31078
R24520 VDD.n968 VDD.t484 3.29673
R24521 VDD.n941 VDD.t485 3.29673
R24522 VDD.n1140 VDD.t483 3.29673
R24523 VDD.n1141 VDD.t476 3.29673
R24524 VDD.n927 VDD.t482 3.29673
R24525 VDD.n926 VDD.t480 3.29673
R24526 VDD.n730 VDD.t481 3.29673
R24527 VDD.n731 VDD.t474 3.29673
R24528 VDD.n1289 VDD.t381 3.29673
R24529 VDD.n1288 VDD.t380 3.29673
R24530 VDD.n1119 VDD.t479 3.29673
R24531 VDD.n1120 VDD.t478 3.29673
R24532 VDD.n1191 VDD.t477 3.29673
R24533 VDD.n1321 VDD.t384 3.29673
R24534 VDD.n1320 VDD.t378 3.29673
R24535 VDD.n826 VDD.t472 3.29673
R24536 VDD.n1366 VDD.t388 3.29673
R24537 VDD.n5766 VDD.n5761 3.27995
R24538 VDD.n5833 VDD.n5828 3.27995
R24539 VDD.n5650 VDD.n5645 3.27995
R24540 VDD.n5568 VDD.n5563 3.27995
R24541 VDD.n8154 VDD.n8149 3.27995
R24542 VDD.n66 VDD.n62 3.27994
R24543 VDD.n155 VDD.n151 3.27994
R24544 VDD.n9110 VDD.n9106 3.27994
R24545 VDD.n8823 VDD.n8819 3.27994
R24546 VDD.n8963 VDD.n8959 3.27994
R24547 VDD.n1661 VDD.t3119 3.22144
R24548 VDD.t2937 VDD.n1643 3.22144
R24549 VDD.t1008 VDD.n6714 3.21228
R24550 VDD.n8637 VDD.t1810 3.20383
R24551 VDD.t2642 VDD.n12 3.20383
R24552 VDD.n12616 VDD.t1468 3.20383
R24553 VDD.n12620 VDD.t2666 3.20383
R24554 VDD.n12598 VDD.t4189 3.20383
R24555 VDD.n12594 VDD.t756 3.20383
R24556 VDD.n12591 VDD.t3829 3.20383
R24557 VDD.n12587 VDD.t781 3.20383
R24558 VDD.n12544 VDD.t4267 3.20383
R24559 VDD.n12548 VDD.t849 3.20383
R24560 VDD.n12550 VDD.t3917 3.20383
R24561 VDD.n12554 VDD.t1294 3.20383
R24562 VDD.n8654 VDD.t1907 3.20383
R24563 VDD.n8650 VDD.t2736 3.20383
R24564 VDD.n8648 VDD.t1543 3.20383
R24565 VDD.n8623 VDD.t3191 3.20383
R24566 VDD.n8675 VDD.t3682 3.20383
R24567 VDD.n8671 VDD.t731 3.20383
R24568 VDD.n8669 VDD.t3347 3.20383
R24569 VDD.n8665 VDD.t767 3.20383
R24570 VDD.n65 VDD.t533 3.20383
R24571 VDD.n67 VDD.t538 3.20383
R24572 VDD.n79 VDD.t1855 3.20383
R24573 VDD.n53 VDD.t3129 3.20383
R24574 VDD.n51 VDD.t1495 3.20383
R24575 VDD.t3153 VDD.n26 3.20383
R24576 VDD.n12504 VDD.t799 3.20383
R24577 VDD.n12500 VDD.t2426 3.20383
R24578 VDD.n94 VDD.t2244 3.20383
R24579 VDD.n90 VDD.t1999 3.20383
R24580 VDD.n8687 VDD.t2685 3.20383
R24581 VDD.n8683 VDD.t4183 3.20383
R24582 VDD.n8681 VDD.t4049 3.20383
R24583 VDD.n8677 VDD.t3819 3.20383
R24584 VDD.n8713 VDD.t2790 3.20383
R24585 VDD.n8709 VDD.t4261 3.20383
R24586 VDD.n8707 VDD.t1634 3.20383
R24587 VDD.n8607 VDD.t1406 3.20383
R24588 VDD.n12488 VDD.t906 3.20383
R24589 VDD.n12492 VDD.t2525 3.20383
R24590 VDD.n12494 VDD.t3997 3.20383
R24591 VDD.n12498 VDD.t3773 3.20383
R24592 VDD.n154 VDD.t4764 3.20383
R24593 VDD.n156 VDD.t4762 3.20383
R24594 VDD.n168 VDD.t2732 3.20383
R24595 VDD.n142 VDD.t4229 3.20383
R24596 VDD.n140 VDD.t4079 3.20383
R24597 VDD.t3859 VDD.n106 3.20383
R24598 VDD.n8725 VDD.t4455 3.20383
R24599 VDD.n8721 VDD.t1853 3.20383
R24600 VDD.n8719 VDD.t1711 3.20383
R24601 VDD.n8715 VDD.t1490 3.20383
R24602 VDD.n8746 VDD.t2348 3.20383
R24603 VDD.n8742 VDD.t3851 3.20383
R24604 VDD.n8740 VDD.t2386 3.20383
R24605 VDD.n8736 VDD.t2101 3.20383
R24606 VDD.n5721 VDD.t4223 3.20383
R24607 VDD.t1756 VDD.n1770 3.20383
R24608 VDD.n11032 VDD.t1244 3.20383
R24609 VDD.n11036 VDD.t3592 3.20383
R24610 VDD.n11021 VDD.t3694 3.20383
R24611 VDD.n11025 VDD.t2616 3.20383
R24612 VDD.n1778 VDD.t585 3.20383
R24613 VDD.n1774 VDD.t3947 3.20383
R24614 VDD.n1823 VDD.t4453 3.20383
R24615 VDD.n1819 VDD.t3317 3.20383
R24616 VDD.n1817 VDD.t1360 3.20383
R24617 VDD.n1808 VDD.t1556 3.20383
R24618 VDD.n5733 VDD.t3649 3.20383
R24619 VDD.n5729 VDD.t1228 3.20383
R24620 VDD.n5727 VDD.t733 3.20383
R24621 VDD.n5723 VDD.t1618 3.20383
R24622 VDD.n5776 VDD.t1319 3.20383
R24623 VDD.n5750 VDD.t1663 3.20383
R24624 VDD.n5748 VDD.t2658 3.20383
R24625 VDD.n5744 VDD.t3491 3.20383
R24626 VDD.n5765 VDD.t369 3.20383
R24627 VDD.n5767 VDD.t421 3.20383
R24628 VDD.n10982 VDD.t1504 3.20383
R24629 VDD.n10978 VDD.t1388 3.20383
R24630 VDD.n1829 VDD.t2693 3.20383
R24631 VDD.n1825 VDD.t2889 3.20383
R24632 VDD.n10966 VDD.t1139 3.20383
R24633 VDD.n10970 VDD.t1332 3.20383
R24634 VDD.n10972 VDD.t3629 3.20383
R24635 VDD.n10976 VDD.t2521 3.20383
R24636 VDD.n5788 VDD.t1364 3.20383
R24637 VDD.n5784 VDD.t2367 3.20383
R24638 VDD.n5782 VDD.t2144 3.20383
R24639 VDD.n5778 VDD.t3525 3.20383
R24640 VDD.n5809 VDD.t872 3.20383
R24641 VDD.n5805 VDD.t1729 3.20383
R24642 VDD.n5803 VDD.t3985 3.20383
R24643 VDD.n5799 VDD.t1178 3.20383
R24644 VDD.n1879 VDD.t1902 3.20383
R24645 VDD.n1875 VDD.t2120 3.20383
R24646 VDD.n1873 VDD.t706 3.20383
R24647 VDD.n1864 VDD.t3655 3.20383
R24648 VDD.n10927 VDD.t3201 3.20383
R24649 VDD.n10923 VDD.t3356 3.20383
R24650 VDD.n1894 VDD.t1446 3.20383
R24651 VDD.n1890 VDD.t4403 3.20383
R24652 VDD.n5843 VDD.t2777 3.20383
R24653 VDD.n5817 VDD.t3594 3.20383
R24654 VDD.n5815 VDD.t3459 3.20383
R24655 VDD.n5811 VDD.t648 3.20383
R24656 VDD.n5832 VDD.t4799 3.20383
R24657 VDD.n5834 VDD.t4798 3.20383
R24658 VDD.n5864 VDD.t2927 3.20383
R24659 VDD.n5860 VDD.t3751 3.20383
R24660 VDD.n5858 VDD.t4627 3.20383
R24661 VDD.n5854 VDD.t1844 3.20383
R24662 VDD.n10911 VDD.t3370 3.20383
R24663 VDD.n10915 VDD.t3572 3.20383
R24664 VDD.n10917 VDD.t576 3.20383
R24665 VDD.n10921 VDD.t3569 3.20383
R24666 VDD.n5527 VDD.t4563 3.20383
R24667 VDD.n5523 VDD.t3400 3.20383
R24668 VDD.n5521 VDD.t2975 3.20383
R24669 VDD.n5512 VDD.t612 3.20383
R24670 VDD.n5876 VDD.t4677 3.20383
R24671 VDD.n5872 VDD.t1889 3.20383
R24672 VDD.n5870 VDD.t936 3.20383
R24673 VDD.n5866 VDD.t3698 3.20383
R24674 VDD.n5637 VDD.t2819 3.20383
R24675 VDD.n5660 VDD.t1342 3.20383
R24676 VDD.n5662 VDD.t870 3.20383
R24677 VDD.n5666 VDD.t3215 3.20383
R24678 VDD.n5649 VDD.t4752 3.20383
R24679 VDD.n5651 VDD.t4751 3.20383
R24680 VDD.n10872 VDD.t2265 3.20383
R24681 VDD.n10868 VDD.t4165 3.20383
R24682 VDD.n5505 VDD.t2262 3.20383
R24683 VDD.n5509 VDD.t1382 3.20383
R24684 VDD.n10856 VDD.t2545 3.20383
R24685 VDD.n10860 VDD.t668 3.20383
R24686 VDD.n10862 VDD.t3015 3.20383
R24687 VDD.n10866 VDD.t2098 3.20383
R24688 VDD.n5616 VDD.t2985 3.20383
R24689 VDD.n5620 VDD.t3907 3.20383
R24690 VDD.n5622 VDD.t3392 3.20383
R24691 VDD.n5626 VDD.t1515 3.20383
R24692 VDD.n5595 VDD.t4725 3.20383
R24693 VDD.n5599 VDD.t3366 3.20383
R24694 VDD.n5601 VDD.t2924 3.20383
R24695 VDD.n5605 VDD.t3749 3.20383
R24696 VDD.n1971 VDD.t3680 3.20383
R24697 VDD.n1967 VDD.t1409 3.20383
R24698 VDD.n1965 VDD.t3677 3.20383
R24699 VDD.n1956 VDD.t3889 3.20383
R24700 VDD.n10814 VDD.t4437 3.20383
R24701 VDD.n10810 VDD.t3291 3.20383
R24702 VDD.n1986 VDD.t4433 3.20383
R24703 VDD.n1982 VDD.t4635 3.20383
R24704 VDD.t4211 VDD.n2104 3.20383
R24705 VDD.n5578 VDD.t1394 3.20383
R24706 VDD.n5580 VDD.t2381 3.20383
R24707 VDD.n5584 VDD.t3267 3.20383
R24708 VDD.n5567 VDD.t499 3.20383
R24709 VDD.n5569 VDD.t513 3.20383
R24710 VDD.n8109 VDD.t4107 3.20383
R24711 VDD.n8105 VDD.t865 3.20383
R24712 VDD.n8103 VDD.t675 3.20383
R24713 VDD.n8099 VDD.t2085 3.20383
R24714 VDD.n10798 VDD.t2742 3.20383
R24715 VDD.n10802 VDD.t2939 3.20383
R24716 VDD.n10804 VDD.t1004 3.20383
R24717 VDD.n10808 VDD.t3939 3.20383
R24718 VDD.n2053 VDD.t3425 3.20383
R24719 VDD.n2049 VDD.t3615 3.20383
R24720 VDD.n2047 VDD.t1714 3.20383
R24721 VDD.n2038 VDD.t4683 3.20383
R24722 VDD.n8121 VDD.t3551 3.20383
R24723 VDD.n8117 VDD.t4451 3.20383
R24724 VDD.n8115 VDD.t4299 3.20383
R24725 VDD.n8111 VDD.t1498 3.20383
R24726 VDD.n8164 VDD.t1207 3.20383
R24727 VDD.n8138 VDD.t2151 3.20383
R24728 VDD.n8136 VDD.t1982 3.20383
R24729 VDD.n8132 VDD.t3368 3.20383
R24730 VDD.n8153 VDD.t4767 3.20383
R24731 VDD.n8155 VDD.t4766 3.20383
R24732 VDD.n10767 VDD.t4617 3.20383
R24733 VDD.n10771 VDD.t673 3.20383
R24734 VDD.n2059 VDD.t3041 3.20383
R24735 VDD.n2055 VDD.t1733 3.20383
R24736 VDD.t2333 VDD.n2241 3.20383
R24737 VDD.n7095 VDD.t2333 3.20383
R24738 VDD.n7096 VDD.t3109 3.20383
R24739 VDD.n7105 VDD.t3971 3.20383
R24740 VDD.t3047 VDD.n7106 3.20383
R24741 VDD.n7113 VDD.t1922 3.20383
R24742 VDD.n7114 VDD.t2428 3.20383
R24743 VDD.n7123 VDD.t2250 3.20383
R24744 VDD.t4337 VDD.n2241 3.20383
R24745 VDD.n7095 VDD.t4337 3.20383
R24746 VDD.n7096 VDD.t973 3.20383
R24747 VDD.n7105 VDD.t1841 3.20383
R24748 VDD.n7106 VDD.t904 3.20383
R24749 VDD.n7113 VDD.t4005 3.20383
R24750 VDD.n7114 VDD.t4393 3.20383
R24751 VDD.n7123 VDD.t4285 3.20383
R24752 VDD.t1816 VDD.n2265 3.20383
R24753 VDD.n7079 VDD.t2841 3.20383
R24754 VDD.t1737 VDD.n7080 3.20383
R24755 VDD.t735 VDD.n7064 3.20383
R24756 VDD.n7061 VDD.t1135 3.20383
R24757 VDD.n7051 VDD.t1025 3.20383
R24758 VDD.n7050 VDD.t1064 3.20383
R24759 VDD.t1064 VDD.n7049 3.20383
R24760 VDD.t698 VDD.n2342 3.20383
R24761 VDD.n6656 VDD.t698 3.20383
R24762 VDD.n6657 VDD.t1438 3.20383
R24763 VDD.n6666 VDD.t1317 3.20383
R24764 VDD.t834 VDD.n6667 3.20383
R24765 VDD.n6674 VDD.t4493 3.20383
R24766 VDD.n6675 VDD.t4013 3.20383
R24767 VDD.n6684 VDD.t3416 3.20383
R24768 VDD.t1835 VDD.n2265 3.20383
R24769 VDD.n7079 VDD.t2855 3.20383
R24770 VDD.n7080 VDD.t1752 3.20383
R24771 VDD.n7064 VDD.t761 3.20383
R24772 VDD.n7061 VDD.t1148 3.20383
R24773 VDD.t1037 VDD.n7051 3.20383
R24774 VDD.n7050 VDD.t1074 3.20383
R24775 VDD.n7049 VDD.t1074 3.20383
R24776 VDD.t719 VDD.n2342 3.20383
R24777 VDD.n6656 VDD.t719 3.20383
R24778 VDD.n6657 VDD.t1470 3.20383
R24779 VDD.n6666 VDD.t1330 3.20383
R24780 VDD.n6667 VDD.t861 3.20383
R24781 VDD.n6674 VDD.t4507 3.20383
R24782 VDD.n6675 VDD.t4027 3.20383
R24783 VDD.n6684 VDD.t3431 3.20383
R24784 VDD.n2396 VDD.t3271 3.20383
R24785 VDD.n7033 VDD.t3151 3.20383
R24786 VDD.t2652 VDD.n7034 3.20383
R24787 VDD.n6718 VDD.t2106 3.20383
R24788 VDD.t1554 VDD.n6719 3.20383
R24789 VDD.n6875 VDD.t3590 3.20383
R24790 VDD.n6866 VDD.t4479 3.20383
R24791 VDD.n6865 VDD.t3515 3.20383
R24792 VDD.t2557 VDD.n6858 3.20383
R24793 VDD.n6857 VDD.t2977 3.20383
R24794 VDD.n2403 VDD.t2845 3.20383
R24795 VDD.t2764 VDD.n2322 3.20383
R24796 VDD.n5244 VDD.t2638 3.20383
R24797 VDD.t2042 VDD.n5245 3.20383
R24798 VDD.n5252 VDD.t1534 3.20383
R24799 VDD.n5253 VDD.t1048 3.20383
R24800 VDD.n5262 VDD.t4573 3.20383
R24801 VDD.t4727 VDD.n2322 3.20383
R24802 VDD.n5244 VDD.t4579 3.20383
R24803 VDD.n5245 VDD.t4103 3.20383
R24804 VDD.n5252 VDD.t3623 3.20383
R24805 VDD.n5253 VDD.t3163 3.20383
R24806 VDD.n5262 VDD.t2594 3.20383
R24807 VDD.n6360 VDD.t4419 3.20383
R24808 VDD.n6350 VDD.t4301 3.20383
R24809 VDD.n6349 VDD.t3789 3.20383
R24810 VDD.t2337 VDD.n6342 3.20383
R24811 VDD.n6341 VDD.t3231 3.20383
R24812 VDD.n6331 VDD.t4097 3.20383
R24813 VDD.n6330 VDD.t4373 3.20383
R24814 VDD.t4373 VDD.n6329 3.20383
R24815 VDD.n6360 VDD.t3339 3.20383
R24816 VDD.t3265 VDD.n6350 3.20383
R24817 VDD.n6349 VDD.t2788 3.20383
R24818 VDD.n6342 VDD.t1170 3.20383
R24819 VDD.n6341 VDD.t2089 3.20383
R24820 VDD.t3057 VDD.n6331 3.20383
R24821 VDD.n6330 VDD.t3311 3.20383
R24822 VDD.n6329 VDD.t3311 3.20383
R24823 VDD.n5445 VDD.t632 3.20383
R24824 VDD.n5454 VDD.t4669 3.20383
R24825 VDD.t4177 VDD.n5455 3.20383
R24826 VDD.n5462 VDD.t3690 3.20383
R24827 VDD.n5463 VDD.t4543 3.20383
R24828 VDD.n5472 VDD.t3995 3.20383
R24829 VDD.n5445 VDD.t3702 3.20383
R24830 VDD.n5454 VDD.t3584 3.20383
R24831 VDD.n5455 VDD.t3123 3.20383
R24832 VDD.n5462 VDD.t2680 3.20383
R24833 VDD.n5463 VDD.t3501 3.20383
R24834 VDD.n5472 VDD.t2973 3.20383
R24835 VDD.n6593 VDD.t2461 3.20383
R24836 VDD.n6584 VDD.t2285 3.20383
R24837 VDD.n6583 VDD.t1702 3.20383
R24838 VDD.n5926 VDD.t1246 3.20383
R24839 VDD.n5927 VDD.t2175 3.20383
R24840 VDD.n5936 VDD.t1530 3.20383
R24841 VDD.t3901 VDD.n5265 3.20383
R24842 VDD.n6242 VDD.t3771 3.20383
R24843 VDD.t3293 VDD.n6243 3.20383
R24844 VDD.n6250 VDD.t2867 3.20383
R24845 VDD.n6251 VDD.t3665 3.20383
R24846 VDD.n6260 VDD.t3143 3.20383
R24847 VDD.t737 VDD.n6261 3.20383
R24848 VDD.n6262 VDD.t737 3.20383
R24849 VDD.t1692 VDD.n6267 3.20383
R24850 VDD.n6268 VDD.t1692 3.20383
R24851 VDD.n6269 VDD.t3535 3.20383
R24852 VDD.n6278 VDD.t3412 3.20383
R24853 VDD.t2965 VDD.n6279 3.20383
R24854 VDD.n6286 VDD.t1350 3.20383
R24855 VDD.n6287 VDD.t2312 3.20383
R24856 VDD.n6296 VDD.t3235 3.20383
R24857 VDD.t3493 VDD.n6297 3.20383
R24858 VDD.n6298 VDD.t3493 3.20383
R24859 VDD.t3919 VDD.n5265 3.20383
R24860 VDD.n6242 VDD.t3787 3.20383
R24861 VDD.n6243 VDD.t3301 3.20383
R24862 VDD.n6250 VDD.t2879 3.20383
R24863 VDD.n6251 VDD.t3684 3.20383
R24864 VDD.n6260 VDD.t3157 3.20383
R24865 VDD.n6261 VDD.t763 3.20383
R24866 VDD.n6262 VDD.t763 3.20383
R24867 VDD.n6267 VDD.t1708 3.20383
R24868 VDD.n6268 VDD.t1708 3.20383
R24869 VDD.n6269 VDD.t3545 3.20383
R24870 VDD.n6278 VDD.t3433 3.20383
R24871 VDD.n6279 VDD.t2981 3.20383
R24872 VDD.n6286 VDD.t1366 3.20383
R24873 VDD.n6287 VDD.t2335 3.20383
R24874 VDD.n6296 VDD.t3249 3.20383
R24875 VDD.n6297 VDD.t3503 3.20383
R24876 VDD.n6298 VDD.t3503 3.20383
R24877 VDD.n5951 VDD.t2011 3.20383
R24878 VDD.n5960 VDD.t1865 3.20383
R24879 VDD.t1339 VDD.n5961 3.20383
R24880 VDD.n5968 VDD.t4025 3.20383
R24881 VDD.n5969 VDD.t765 3.20383
R24882 VDD.n5978 VDD.t1647 3.20383
R24883 VDD.n6380 VDD.t4721 3.20383
R24884 VDD.n6389 VDD.t4571 3.20383
R24885 VDD.t4095 VDD.n6390 3.20383
R24886 VDD.n5997 VDD.t2662 3.20383
R24887 VDD.n5998 VDD.t3483 3.20383
R24888 VDD.n6007 VDD.t4369 3.20383
R24889 VDD.n6009 VDD.t4673 3.20383
R24890 VDD.t4673 VDD.n6008 3.20383
R24891 VDD.n6380 VDD.t2719 3.20383
R24892 VDD.n6389 VDD.t2592 3.20383
R24893 VDD.n6390 VDD.t1980 3.20383
R24894 VDD.n5997 VDD.t4615 3.20383
R24895 VDD.n5998 VDD.t1346 3.20383
R24896 VDD.n6007 VDD.t2341 3.20383
R24897 VDD.n6009 VDD.t2668 3.20383
R24898 VDD.n6008 VDD.t2668 3.20383
R24899 VDD.t963 VDD.n5263 3.20383
R24900 VDD.n5343 VDD.t824 3.20383
R24901 VDD.t4443 VDD.n5344 3.20383
R24902 VDD.n5351 VDD.t3999 3.20383
R24903 VDD.n5352 VDD.t717 3.20383
R24904 VDD.n5361 VDD.t4279 3.20383
R24905 VDD.t3079 VDD.n5263 3.20383
R24906 VDD.n5343 VDD.t2963 3.20383
R24907 VDD.n5344 VDD.t2434 3.20383
R24908 VDD.n5351 VDD.t1874 3.20383
R24909 VDD.n5352 VDD.t2863 3.20383
R24910 VDD.n5361 VDD.t2204 3.20383
R24911 VDD.n6412 VDD.t1111 3.20383
R24912 VDD.n6403 VDD.t1006 3.20383
R24913 VDD.n6402 VDD.t4597 3.20383
R24914 VDD.n6161 VDD.t3171 3.20383
R24915 VDD.n6162 VDD.t4015 3.20383
R24916 VDD.n6171 VDD.t779 3.20383
R24917 VDD.t1454 VDD.n2410 3.20383
R24918 VDD.n6570 VDD.t1321 3.20383
R24919 VDD.t853 VDD.n6571 3.20383
R24920 VDD.n6028 VDD.t4501 3.20383
R24921 VDD.t1234 VDD.n6029 3.20383
R24922 VDD.t650 VDD.n6024 3.20383
R24923 VDD.n2216 VDD.t1217 3.20383
R24924 VDD.n2227 VDD.t4387 3.20383
R24925 VDD.n2219 VDD.t3380 3.20383
R24926 VDD.n2218 VDD.t3793 3.20383
R24927 VDD.t3647 VDD.n7980 3.20383
R24928 VDD.n7976 VDD.t3688 3.20383
R24929 VDD.t3688 VDD.n7975 3.20383
R24930 VDD.n7969 VDD.t3351 3.20383
R24931 VDD.t3351 VDD.n7968 3.20383
R24932 VDD.n7965 VDD.t4133 3.20383
R24933 VDD.n7851 VDD.t2786 3.20383
R24934 VDD.t2786 VDD.n7850 3.20383
R24935 VDD.n2215 VDD.t4481 3.20383
R24936 VDD.t4361 VDD.n2193 3.20383
R24937 VDD.n7986 VDD.t1109 3.20383
R24938 VDD.t3402 VDD.n7983 3.20383
R24939 VDD.n7979 VDD.t1432 3.20383
R24940 VDD.n7966 VDD.t1884 3.20383
R24941 VDD.t2758 VDD.n2202 3.20383
R24942 VDD.n2203 VDD.t2758 3.20383
R24943 VDD.n6605 VDD.t3991 3.20383
R24944 VDD.t3481 VDD.n6606 3.20383
R24945 VDD.n6613 VDD.t3073 3.20383
R24946 VDD.n6614 VDD.t2566 3.20383
R24947 VDD.n6623 VDD.t1867 3.20383
R24948 VDD.t2463 VDD.n2310 3.20383
R24949 VDD.n5415 VDD.t2287 3.20383
R24950 VDD.t1704 VDD.n5416 3.20383
R24951 VDD.n5423 VDD.t1248 3.20383
R24952 VDD.n5424 VDD.t769 3.20383
R24953 VDD.n5433 VDD.t4303 3.20383
R24954 VDD.t1261 VDD.n2310 3.20383
R24955 VDD.n5415 VDD.t1137 3.20383
R24956 VDD.n5416 VDD.t605 3.20383
R24957 VDD.n5423 VDD.t4319 3.20383
R24958 VDD.n5424 VDD.t3809 3.20383
R24959 VDD.n5433 VDD.t3263 3.20383
R24960 VDD.n7174 VDD.t1978 3.20383
R24961 VDD.t1978 VDD.n7173 3.20383
R24962 VDD.n7172 VDD.t2835 3.20383
R24963 VDD.n7162 VDD.t3653 3.20383
R24964 VDD.n7161 VDD.t2762 3.20383
R24965 VDD.t1622 VDD.n7154 3.20383
R24966 VDD.n7153 VDD.t2077 3.20383
R24967 VDD.n7143 VDD.t1917 3.20383
R24968 VDD.n7174 VDD.t916 3.20383
R24969 VDD.n7173 VDD.t916 3.20383
R24970 VDD.n7172 VDD.t1636 3.20383
R24971 VDD.t2656 VDD.n7162 3.20383
R24972 VDD.n7161 VDD.t1549 3.20383
R24973 VDD.n7154 VDD.t4689 3.20383
R24974 VDD.n7153 VDD.t989 3.20383
R24975 VDD.t851 VDD.n7143 3.20383
R24976 VDD.n7843 VDD.t4467 3.20383
R24977 VDD.n2173 VDD.t2804 3.20383
R24978 VDD.n2182 VDD.t2672 3.20383
R24979 VDD.t3495 VDD.n2183 3.20383
R24980 VDD.n8000 VDD.t1587 3.20383
R24981 VDD.n8001 VDD.t3835 3.20383
R24982 VDD.n8010 VDD.t4277 3.20383
R24983 VDD.t3519 VDD.n8459 3.20383
R24984 VDD.t3323 VDD.n9130 3.20383
R24985 VDD.t3001 VDD.n8459 3.20383
R24986 VDD.n9130 VDD.t2796 3.20383
R24987 VDD.n9139 VDD.t2549 3.20383
R24988 VDD.n9143 VDD.t4043 3.20383
R24989 VDD.n9145 VDD.t3899 3.20383
R24990 VDD.n9149 VDD.t3673 3.20383
R24991 VDD.n9166 VDD.t3103 3.20383
R24992 VDD.n9162 VDD.t4569 3.20383
R24993 VDD.t4461 VDD.n8472 3.20383
R24994 VDD.n8488 VDD.t4257 3.20383
R24995 VDD.n9109 VDD.t4790 3.20383
R24996 VDD.n9111 VDD.t4791 3.20383
R24997 VDD.n8763 VDD.t4061 3.20383
R24998 VDD.n8759 VDD.t3841 3.20383
R24999 VDD.n8757 VDD.t4517 3.20383
R25000 VDD.n8582 VDD.t3861 3.20383
R25001 VDD.n8559 VDD.t2255 3.20383
R25002 VDD.n8555 VDD.t2024 3.20383
R25003 VDD.n8553 VDD.t2815 3.20383
R25004 VDD.t2062 VDD.n184 3.20383
R25005 VDD.n8822 VDD.t9 3.20383
R25006 VDD.n8824 VDD.t4 3.20383
R25007 VDD.n8836 VDD.t2871 3.20383
R25008 VDD.n8810 VDD.t2112 3.20383
R25009 VDD.t1035 VDD.n8526 3.20383
R25010 VDD.n8547 VDD.t2134 3.20383
R25011 VDD.n8799 VDD.t4585 3.20383
R25012 VDD.n8803 VDD.t3935 3.20383
R25013 VDD.n8769 VDD.t2943 3.20383
R25014 VDD.n8765 VDD.t3959 3.20383
R25015 VDD.n8889 VDD.t2523 3.20383
R25016 VDD.n8885 VDD.t3447 3.20383
R25017 VDD.t2440 VDD.n8518 3.20383
R25018 VDD.n8775 VDD.t3471 3.20383
R25019 VDD.n8872 VDD.t581 3.20383
R25020 VDD.n8876 VDD.t1593 3.20383
R25021 VDD.n8842 VDD.t4693 3.20383
R25022 VDD.n8838 VDD.t1620 3.20383
R25023 VDD.n8945 VDD.t2470 3.20383
R25024 VDD.n8941 VDD.t1678 3.20383
R25025 VDD.t600 VDD.n8507 3.20383
R25026 VDD.n8848 VDD.t2214 3.20383
R25027 VDD.n8930 VDD.t4227 3.20383
R25028 VDD.n8934 VDD.t3527 3.20383
R25029 VDD.n8900 VDD.t2531 3.20383
R25030 VDD.n8513 VDD.t4019 3.20383
R25031 VDD.n9020 VDD.t4291 3.20383
R25032 VDD.n9016 VDD.t4083 3.20383
R25033 VDD.t2626 VDD.n8499 3.20383
R25034 VDD.n8906 VDD.t4111 3.20383
R25035 VDD.n8962 VDD.t4804 3.20383
R25036 VDD.n8964 VDD.t4800 3.20383
R25037 VDD.n8999 VDD.t2562 3.20383
R25038 VDD.n9007 VDD.t2292 3.20383
R25039 VDD.n8951 VDD.t711 3.20383
R25040 VDD.n8947 VDD.t2329 3.20383
R25041 VDD.n9042 VDD.t3025 3.20383
R25042 VDD.n9038 VDD.t4487 3.20383
R25043 VDD.t4367 VDD.n8490 3.20383
R25044 VDD.n8975 VDD.t4179 3.20383
R25045 VDD.t565 VDD.n8476 3.20383
R25046 VDD.n9031 VDD.t2194 3.20383
R25047 VDD.n9026 VDD.t2065 3.20383
R25048 VDD.n9022 VDD.t1799 3.20383
R25049 VDD.n9151 VDD.t684 3.20383
R25050 VDD.n9155 VDD.t2306 3.20383
R25051 VDD.n9073 VDD.t2132 3.20383
R25052 VDD.n8475 VDD.t1896 3.20383
R25053 VDD.n190 VDD.t4605 3.20383
R25054 VDD.n186 VDD.t2047 3.20383
R25055 VDD.n174 VDD.t4631 3.20383
R25056 VDD.n170 VDD.t4407 3.20383
R25057 VDD.n9123 VDD.t627 3.20383
R25058 VDD.n9097 VDD.t2232 3.20383
R25059 VDD.n9095 VDD.t2092 3.20383
R25060 VDD.t1839 VDD.n8470 3.20383
R25061 VDD.n1162 VDD.t4199 3.20383
R25062 VDD.t4199 VDD.n1161 3.20383
R25063 VDD.n1160 VDD.t1680 3.20383
R25064 VDD.n1748 VDD.t741 3.20383
R25065 VDD.t3051 VDD.n1749 3.20383
R25066 VDD.n1750 VDD.t3051 3.20383
R25067 VDD.t2913 VDD.n1711 3.20383
R25068 VDD.n1712 VDD.t2913 3.20383
R25069 VDD.t3137 VDD.n1713 3.20383
R25070 VDD.n722 VDD.t2723 3.20383
R25071 VDD.n721 VDD.t4287 3.20383
R25072 VDD.t4287 VDD.n720 3.20383
R25073 VDD.n719 VDD.t2537 3.20383
R25074 VDD.t2537 VDD.n700 3.20383
R25075 VDD.t1785 VDD.n1733 3.20383
R25076 VDD.n1734 VDD.t1785 3.20383
R25077 VDD.n1711 VDD.t2701 3.20383
R25078 VDD.n1712 VDD.t2701 3.20383
R25079 VDD.n1713 VDD.t2941 3.20383
R25080 VDD.t2509 VDD.n722 3.20383
R25081 VDD.n721 VDD.t4069 3.20383
R25082 VDD.n720 VDD.t4069 3.20383
R25083 VDD.n719 VDD.t2252 3.20383
R25084 VDD.t2252 VDD.n700 3.20383
R25085 VDD.n1733 VDD.t1575 3.20383
R25086 VDD.n1734 VDD.t1575 3.20383
R25087 VDD.t1371 VDD.n1735 3.20383
R25088 VDD.n1736 VDD.t1371 3.20383
R25089 VDD.t1506 VDD.n1737 3.20383
R25090 VDD.n948 VDD.t3817 3.20383
R25091 VDD.t2831 VDD.n950 3.20383
R25092 VDD.n951 VDD.t2831 3.20383
R25093 VDD.n916 VDD.t4463 3.20383
R25094 VDD.t4463 VDD.n915 3.20383
R25095 VDD.n914 VDD.t4583 3.20383
R25096 VDD.t2827 VDD.n907 3.20383
R25097 VDD.n906 VDD.t1649 3.20383
R25098 VDD.t1649 VDD.n905 3.20383
R25099 VDD.n1071 VDD.t1725 3.20383
R25100 VDD.t1725 VDD.n1070 3.20383
R25101 VDD.n1069 VDD.t1986 3.20383
R25102 VDD.t1528 VDD.n1062 3.20383
R25103 VDD.n1061 VDD.t3259 3.20383
R25104 VDD.t3259 VDD.n1060 3.20383
R25105 VDD.n1494 VDD.t4639 3.20383
R25106 VDD.t4639 VDD.n1493 3.20383
R25107 VDD.n1492 VDD.t739 3.20383
R25108 VDD.t1684 VDD.n1485 3.20383
R25109 VDD.n1484 VDD.t1930 3.20383
R25110 VDD.t1930 VDD.n1483 3.20383
R25111 VDD.n1482 VDD.t1772 3.20383
R25112 VDD.t1772 VDD.n1481 3.20383
R25113 VDD.n1461 VDD.t2660 3.20383
R25114 VDD.t2660 VDD.n1460 3.20383
R25115 VDD.n1459 VDD.t743 3.20383
R25116 VDD.t743 VDD.n1458 3.20383
R25117 VDD.n1457 VDD.t4739 3.20383
R25118 VDD.t1934 VDD.n1450 3.20383
R25119 VDD.t4529 VDD.n821 3.20383
R25120 VDD.n1445 VDD.t4529 3.20383
R25121 VDD.n1444 VDD.t4157 3.20383
R25122 VDD.t4157 VDD.n1443 3.20383
R25123 VDD.t3511 VDD.n824 3.20383
R25124 VDD.n1406 VDD.t3511 3.20383
R25125 VDD.t3147 VDD.n1407 3.20383
R25126 VDD.n1408 VDD.t3147 3.20383
R25127 VDD.t1511 VDD.n1409 3.20383
R25128 VDD.n1400 VDD.t1676 3.20383
R25129 VDD.n1399 VDD.t4313 3.20383
R25130 VDD.t4313 VDD.n1398 3.20383
R25131 VDD.n1397 VDD.t3891 3.20383
R25132 VDD.t3891 VDD.n729 3.20383
R25133 VDD.t3297 VDD.n1709 3.20383
R25134 VDD.n1710 VDD.t3297 3.20383
R25135 VDD.n1494 VDD.t4409 3.20383
R25136 VDD.n1493 VDD.t4409 3.20383
R25137 VDD.n1492 VDD.t4655 3.20383
R25138 VDD.n1485 VDD.t1472 3.20383
R25139 VDD.n1484 VDD.t1696 3.20383
R25140 VDD.n1483 VDD.t1696 3.20383
R25141 VDD.n1482 VDD.t1547 3.20383
R25142 VDD.n1481 VDD.t1547 3.20383
R25143 VDD.n1461 VDD.t2423 3.20383
R25144 VDD.n1460 VDD.t2423 3.20383
R25145 VDD.n1459 VDD.t4661 3.20383
R25146 VDD.n1458 VDD.t4661 3.20383
R25147 VDD.n1457 VDD.t4511 3.20383
R25148 VDD.n1450 VDD.t1700 3.20383
R25149 VDD.t4345 VDD.n821 3.20383
R25150 VDD.n1445 VDD.t4345 3.20383
R25151 VDD.n1444 VDD.t3933 3.20383
R25152 VDD.n1443 VDD.t3933 3.20383
R25153 VDD.t3313 VDD.n824 3.20383
R25154 VDD.n1406 VDD.t3313 3.20383
R25155 VDD.n1407 VDD.t2955 3.20383
R25156 VDD.n1408 VDD.t2955 3.20383
R25157 VDD.n1409 VDD.t1298 3.20383
R25158 VDD.t1450 VDD.n1400 3.20383
R25159 VDD.n1399 VDD.t4117 3.20383
R25160 VDD.n1398 VDD.t4117 3.20383
R25161 VDD.n1397 VDD.t3663 3.20383
R25162 VDD.t3663 VDD.n729 3.20383
R25163 VDD.n1709 VDD.t3107 3.20383
R25164 VDD.n1710 VDD.t3107 3.20383
R25165 VDD.n1218 VDD.t2480 3.20383
R25166 VDD.t2480 VDD.n1217 3.20383
R25167 VDD.n1216 VDD.t4671 3.20383
R25168 VDD.t3659 VDD.n1209 3.20383
R25169 VDD.n1208 VDD.t721 3.20383
R25170 VDD.t721 VDD.n1207 3.20383
R25171 VDD.t3420 VDD.n1270 3.20383
R25172 VDD.n1271 VDD.t3420 3.20383
R25173 VDD.t1846 VDD.n1272 3.20383
R25174 VDD.n1239 VDD.t4675 3.20383
R25175 VDD.n1238 VDD.t3195 3.20383
R25176 VDD.t3195 VDD.n1237 3.20383
R25177 VDD.t4151 VDD.n1593 3.20383
R25178 VDD.n1594 VDD.t4151 3.20383
R25179 VDD.t3708 VDD.n1595 3.20383
R25180 VDD.n1596 VDD.t3708 3.20383
R25181 VDD.t2189 VDD.n1597 3.20383
R25182 VDD.n1604 VDD.t786 3.20383
R25183 VDD.t3396 VDD.n1605 3.20383
R25184 VDD.n1606 VDD.t3396 3.20383
R25185 VDD.t1524 VDD.n1607 3.20383
R25186 VDD.n1608 VDD.t1524 3.20383
R25187 VDD.n1496 VDD.t2409 3.20383
R25188 VDD.t2409 VDD.n1495 3.20383
R25189 VDD.n1593 VDD.t3925 3.20383
R25190 VDD.n1594 VDD.t3925 3.20383
R25191 VDD.n1595 VDD.t3507 3.20383
R25192 VDD.n1596 VDD.t3507 3.20383
R25193 VDD.n1597 VDD.t1943 3.20383
R25194 VDD.n1604 VDD.t4697 3.20383
R25195 VDD.n1605 VDD.t3221 3.20383
R25196 VDD.n1606 VDD.t3221 3.20383
R25197 VDD.n1607 VDD.t1311 3.20383
R25198 VDD.n1608 VDD.t1311 3.20383
R25199 VDD.n1496 VDD.t2114 3.20383
R25200 VDD.n1495 VDD.t2114 3.20383
R25201 VDD.n1528 VDD.t1626 3.20383
R25202 VDD.t1872 VDD.n1518 3.20383
R25203 VDD.n1517 VDD.t696 3.20383
R25204 VDD.t2432 VDD.n771 3.20383
R25205 VDD.n1555 VDD.t4779 3.20383
R25206 VDD.n1555 VDD.t4776 3.20383
R25207 VDD.n1556 VDD.t4781 3.20383
R25208 VDD.n1556 VDD.t4778 3.20383
R25209 VDD.n1557 VDD.t4780 3.20383
R25210 VDD.n1557 VDD.t4777 3.20383
R25211 VDD.n1541 VDD.t998 3.20383
R25212 VDD.n1537 VDD.t1192 3.20383
R25213 VDD.n1559 VDD.t4207 3.20383
R25214 VDD.n1563 VDD.t1668 3.20383
R25215 VDD.n1175 VDD.t1480 3.20383
R25216 VDD.t1480 VDD.n1174 3.20383
R25217 VDD.n1173 VDD.t4141 3.20383
R25218 VDD.t1686 VDD.n1166 3.20383
R25219 VDD.n1165 VDD.t1219 3.20383
R25220 VDD.t1219 VDD.n1164 3.20383
R25221 VDD.n1188 VDD.t4731 3.20383
R25222 VDD.t4731 VDD.n1187 3.20383
R25223 VDD.n1186 VDD.t1762 3.20383
R25224 VDD.t4567 VDD.n1179 3.20383
R25225 VDD.n1178 VDD.t1630 3.20383
R25226 VDD.t1630 VDD.n1177 3.20383
R25227 VDD.t3574 VDD.n1337 3.20383
R25228 VDD.n1338 VDD.t3574 3.20383
R25229 VDD.t3799 VDD.n1339 3.20383
R25230 VDD.n1307 VDD.t593 3.20383
R25231 VDD.n1306 VDD.t884 3.20383
R25232 VDD.t884 VDD.n1305 3.20383
R25233 VDD.t3119 VDD.n1660 3.20383
R25234 VDD.n1659 VDD.t2711 3.20383
R25235 VDD.t2711 VDD.n1658 3.20383
R25236 VDD.n1657 VDD.t1092 3.20383
R25237 VDD.n1316 VDD.t3849 3.20383
R25238 VDD.t2379 VDD.n1317 3.20383
R25239 VDD.n1318 VDD.t2379 3.20383
R25240 VDD.t1996 VDD.n1384 3.20383
R25241 VDD.n1385 VDD.t1996 3.20383
R25242 VDD.t4593 VDD.n1386 3.20383
R25243 VDD.n1075 VDD.t583 3.20383
R25244 VDD.n1074 VDD.t3287 3.20383
R25245 VDD.t3287 VDD.n1073 3.20383
R25246 VDD.n1286 VDD.t3813 3.20383
R25247 VDD.t3813 VDD.n1285 3.20383
R25248 VDD.n1284 VDD.t3669 3.20383
R25249 VDD.n1362 VDD.t892 3.20383
R25250 VDD.t3499 VDD.n1363 3.20383
R25251 VDD.n1364 VDD.t3499 3.20383
R25252 VDD.n1644 VDD.t2937 3.20383
R25253 VDD.t2140 VDD.n1645 3.20383
R25254 VDD.n1646 VDD.t2140 3.20383
R25255 VDD.t3343 VDD.n1647 3.20383
R25256 VDD.n1248 VDD.t3435 3.20383
R25257 VDD.t4599 VDD.n1249 3.20383
R25258 VDD.n1250 VDD.t4599 3.20383
R25259 VDD.n1735 VDD.t1154 3.20383
R25260 VDD.n1736 VDD.t1154 3.20383
R25261 VDD.n1737 VDD.t1289 3.20383
R25262 VDD.n948 VDD.t3600 3.20383
R25263 VDD.n950 VDD.t2622 3.20383
R25264 VDD.n951 VDD.t2622 3.20383
R25265 VDD.n71 VDD.n70 3.2012
R25266 VDD.n160 VDD.n159 3.2012
R25267 VDD.n5770 VDD.n5769 3.2012
R25268 VDD.n5837 VDD.n5836 3.2012
R25269 VDD.n5654 VDD.n5653 3.2012
R25270 VDD.n5572 VDD.n5571 3.2012
R25271 VDD.n8158 VDD.n8157 3.2012
R25272 VDD.n9115 VDD.n9114 3.2012
R25273 VDD.n8828 VDD.n8827 3.2012
R25274 VDD.n8968 VDD.n8967 3.2012
R25275 VDD.n5766 VDD.n5765 3.1154
R25276 VDD.n5833 VDD.n5832 3.1154
R25277 VDD.n5650 VDD.n5649 3.1154
R25278 VDD.n5568 VDD.n5567 3.1154
R25279 VDD.n8154 VDD.n8153 3.1154
R25280 VDD.n66 VDD.n65 3.11413
R25281 VDD.n155 VDD.n154 3.11413
R25282 VDD.n9110 VDD.n9109 3.11413
R25283 VDD.n8823 VDD.n8822 3.11413
R25284 VDD.n8963 VDD.n8962 3.11413
R25285 VDD.n6152 VDD.n6021 3.00663
R25286 VDD.n6095 VDD.n6094 3.00663
R25287 VDD.n6847 VDD.n6846 3.00663
R25288 VDD.n6797 VDD.n6796 3.00663
R25289 VDD.n1425 VDD.n1424 2.89741
R25290 VDD.n1418 VDD.n858 2.89677
R25291 VDD.n1679 VDD.n1678 2.89677
R25292 VDD.n1692 VDD.n1691 2.89677
R25293 VDD.n1626 VDD.n1625 2.89677
R25294 VDD.n1673 VDD.n1672 2.89677
R25295 VDD.n1619 VDD.n784 2.89677
R25296 VDD.n1106 VDD.n1091 2.89677
R25297 VDD.n1685 VDD.n1684 2.89677
R25298 VDD.n1697 VDD.n735 2.89677
R25299 VDD.n1045 VDD.n1039 2.89677
R25300 VDD.n979 VDD.n706 2.89677
R25301 VDD.n1086 VDD.n844 2.89406
R25302 VDD.n1419 VDD.n1418 2.89406
R25303 VDD.n1678 VDD.n1677 2.89406
R25304 VDD.n1690 VDD.n1689 2.89406
R25305 VDD.n1620 VDD.n1619 2.89406
R25306 VDD.n1106 VDD.n1105 2.89406
R25307 VDD.n1684 VDD.n1683 2.89406
R25308 VDD.n1697 VDD.n1696 2.89406
R25309 VDD.n1045 VDD.n1044 2.89406
R25310 VDD.n853 VDD.n706 2.89406
R25311 VDD.n984 VDD.n983 2.89406
R25312 VDD.n1034 VDD.n1033 2.89406
R25313 VDD.n6136 VDD.n6134 2.7866
R25314 VDD.n6139 VDD.n6137 2.7866
R25315 VDD.n6143 VDD.n6141 2.7866
R25316 VDD.n6147 VDD.n6145 2.7866
R25317 VDD.n6132 VDD.n6130 2.7866
R25318 VDD.n6128 VDD.n6126 2.7866
R25319 VDD.n6124 VDD.n6122 2.7866
R25320 VDD.n6120 VDD.n6118 2.7866
R25321 VDD.n6044 VDD.n6042 2.7866
R25322 VDD.n6047 VDD.n6045 2.7866
R25323 VDD.n6051 VDD.n6049 2.7866
R25324 VDD.n6055 VDD.n6053 2.7866
R25325 VDD.n6078 VDD.n6076 2.7866
R25326 VDD.n6082 VDD.n6080 2.7866
R25327 VDD.n6086 VDD.n6084 2.7866
R25328 VDD.n6090 VDD.n6088 2.7866
R25329 VDD.n6810 VDD.n6808 2.7866
R25330 VDD.n6813 VDD.n6811 2.7866
R25331 VDD.n6817 VDD.n6815 2.7866
R25332 VDD.n6821 VDD.n6819 2.7866
R25333 VDD.n6826 VDD.n6824 2.7866
R25334 VDD.n6830 VDD.n6828 2.7866
R25335 VDD.n6834 VDD.n6832 2.7866
R25336 VDD.n6838 VDD.n6836 2.7866
R25337 VDD.n6777 VDD.n6775 2.7866
R25338 VDD.n6780 VDD.n6778 2.7866
R25339 VDD.n6784 VDD.n6782 2.7866
R25340 VDD.n6788 VDD.n6786 2.7866
R25341 VDD.n6773 VDD.n6771 2.7866
R25342 VDD.n6769 VDD.n6767 2.7866
R25343 VDD.n6765 VDD.n6763 2.7866
R25344 VDD.n6761 VDD.n6759 2.7866
R25345 VDD.n7004 VDD.n7002 2.73714
R25346 VDD.n6926 VDD.n6924 2.73714
R25347 VDD.n6541 VDD.n6539 2.73714
R25348 VDD.n6452 VDD.n6450 2.73714
R25349 VDD.n6140 VDD.n6136 2.73672
R25350 VDD.n6048 VDD.n6044 2.73672
R25351 VDD.n6814 VDD.n6810 2.73672
R25352 VDD.n6781 VDD.n6777 2.73672
R25353 VDD.n58 VDD.n57 2.65954
R25354 VDD.n64 VDD.n63 2.65954
R25355 VDD.n147 VDD.n146 2.65954
R25356 VDD.n153 VDD.n152 2.65954
R25357 VDD.n9102 VDD.n9101 2.65954
R25358 VDD.n9108 VDD.n9107 2.65954
R25359 VDD.n8815 VDD.n8814 2.65954
R25360 VDD.n8821 VDD.n8820 2.65954
R25361 VDD.n8955 VDD.n8954 2.65954
R25362 VDD.n8961 VDD.n8960 2.65954
R25363 VDD.n5764 VDD.n5762 2.65924
R25364 VDD.n5757 VDD.n5756 2.65924
R25365 VDD.n5831 VDD.n5829 2.65924
R25366 VDD.n5824 VDD.n5823 2.65924
R25367 VDD.n5648 VDD.n5646 2.65924
R25368 VDD.n5641 VDD.n5640 2.65924
R25369 VDD.n5566 VDD.n5564 2.65924
R25370 VDD.n5559 VDD.n5558 2.65924
R25371 VDD.n8152 VDD.n8150 2.65924
R25372 VDD.n8145 VDD.n8144 2.65924
R25373 VDD.n5767 VDD.n5766 2.61766
R25374 VDD.n5834 VDD.n5833 2.61766
R25375 VDD.n5651 VDD.n5650 2.61766
R25376 VDD.n5569 VDD.n5568 2.61766
R25377 VDD.n8155 VDD.n8154 2.61766
R25378 VDD.n67 VDD.n66 2.61737
R25379 VDD.n156 VDD.n155 2.61737
R25380 VDD.n9111 VDD.n9110 2.61737
R25381 VDD.n8824 VDD.n8823 2.61737
R25382 VDD.n8964 VDD.n8963 2.61737
R25383 VDD.n8064 VDD.n8063 2.60496
R25384 VDD.n7959 VDD.n7958 2.60386
R25385 VDD.n8082 VDD.n8081 2.6005
R25386 VDD.n8083 VDD.n2120 2.6005
R25387 VDD.n8074 VDD.n8073 2.6005
R25388 VDD.n8072 VDD.n8071 2.6005
R25389 VDD.n8054 VDD.n8052 2.59852
R25390 VDD.n7949 VDD.n7947 2.59742
R25391 VDD.n6956 VDD.n6954 2.59712
R25392 VDD.n6924 VDD.n6922 2.59712
R25393 VDD.n7008 VDD.n7006 2.59712
R25394 VDD.n7002 VDD.n7000 2.59712
R25395 VDD.n6500 VDD.n6498 2.59712
R25396 VDD.n6450 VDD.n6448 2.59712
R25397 VDD.n6546 VDD.n6544 2.59712
R25398 VDD.n6539 VDD.n6537 2.59712
R25399 VDD.t3016 VDD.n1529 2.55028
R25400 VDD.t2301 VDD.n1542 2.55022
R25401 VDD.n772 VDD.t4522 2.54061
R25402 VDD.t4522 VDD.n770 2.54061
R25403 VDD.t4588 VDD.n1635 2.54061
R25404 VDD.n1636 VDD.t4588 2.54061
R25405 VDD.t1079 VDD.n1632 2.54061
R25406 VDD.n1633 VDD.t1079 2.54061
R25407 VDD.t922 VDD.n1629 2.54061
R25408 VDD.n1630 VDD.t922 2.54061
R25409 VDD.n1510 VDD.t3874 2.54061
R25410 VDD.t3874 VDD.n782 2.54061
R25411 VDD.n1530 VDD.t3016 2.54061
R25412 VDD.n1532 VDD.t3060 2.54061
R25413 VDD.t3060 VDD.n1531 2.54061
R25414 VDD.n1546 VDD.t3603 2.54061
R25415 VDD.t3603 VDD.n1533 2.54061
R25416 VDD.t3444 VDD.n1544 2.54061
R25417 VDD.n1545 VDD.t3444 2.54061
R25418 VDD.n1543 VDD.t2301 2.54061
R25419 VDD.n2142 VDD.t1027 2.5255
R25420 VDD.n2140 VDD.t2413 2.5255
R25421 VDD.n2137 VDD.t3327 2.5255
R25422 VDD.n2137 VDD.t2300 2.5255
R25423 VDD.n2135 VDD.t775 2.5255
R25424 VDD.n2135 VDD.t3871 2.5255
R25425 VDD.n2132 VDD.t3803 2.5255
R25426 VDD.n2132 VDD.t2847 2.5255
R25427 VDD.n2129 VDD.t1992 2.5255
R25428 VDD.n2129 VDD.t966 2.5255
R25429 VDD.n8067 VDD.t573 2.5255
R25430 VDD.n2147 VDD.t1913 2.5255
R25431 VDD.n2160 VDD.t1831 2.5255
R25432 VDD.n2164 VDD.t3475 2.5255
R25433 VDD.n8015 VDD.t2430 2.5255
R25434 VDD.n2121 VDD.t4687 2.5255
R25435 VDD.n7913 VDD.n7912 2.46986
R25436 VDD.n7909 VDD.n7908 2.46873
R25437 VDD.n8018 VDD.n8017 2.46873
R25438 VDD.n8047 VDD.n8046 2.46198
R25439 VDD.n7891 VDD.n7890 2.46198
R25440 VDD.n7942 VDD.n7941 2.46086
R25441 VDD.n7005 VDD.n7004 2.46014
R25442 VDD.n6958 VDD.n6926 2.46014
R25443 VDD.n6548 VDD.n6541 2.46014
R25444 VDD.n6497 VDD.n6452 2.46014
R25445 VDD.t2843 VDD.n8072 2.4505
R25446 VDD.n8072 VDD.t1362 2.4505
R25447 VDD.n8073 VDD.t945 2.4505
R25448 VDD.n8073 VDD.t2843 2.4505
R25449 VDD.n8083 VDD.t2772 2.4505
R25450 VDD.t1279 VDD.n8083 2.4505
R25451 VDD.n8082 VDD.t863 2.4505
R25452 VDD.t2772 VDD.n8082 2.4505
R25453 VDD.n6956 VDD.n6955 2.39107
R25454 VDD.n6924 VDD.n6923 2.39107
R25455 VDD.n7008 VDD.n7007 2.39107
R25456 VDD.n7002 VDD.n7001 2.39107
R25457 VDD.n6500 VDD.n6499 2.39107
R25458 VDD.n6450 VDD.n6449 2.39107
R25459 VDD.n6546 VDD.n6545 2.39107
R25460 VDD.n6539 VDD.n6538 2.39107
R25461 VDD.n6751 VDD.n6750 2.37568
R25462 VDD.n6064 VDD.n6063 2.37568
R25463 VDD.n6107 VDD.n6106 2.37568
R25464 VDD.n6733 VDD.n6732 2.37568
R25465 VDD.n7892 VDD.n7886 2.37449
R25466 VDD.n7895 VDD.n7882 2.37449
R25467 VDD.n7898 VDD.n7878 2.37449
R25468 VDD.n7904 VDD.n7872 2.37449
R25469 VDD.n7907 VDD.n7868 2.37449
R25470 VDD.n1448 VDD.n1447 2.30715
R25471 VDD.n7024 VDD.n2375 2.30165
R25472 VDD.n6877 VDD.n6876 2.30165
R25473 VDD.n6414 VDD.n6413 2.30165
R25474 VDD.n6561 VDD.n5288 2.30165
R25475 VDD.n5906 VDD.n5905 2.26828
R25476 VDD.n12582 VDD.n12560 2.26741
R25477 VDD.n6172 VDD.n6016 2.26689
R25478 VDD.n3630 VDD.n2745 2.2505
R25479 VDD.n3632 VDD.n3631 2.2505
R25480 VDD.n3633 VDD.n2744 2.2505
R25481 VDD.n3635 VDD.n3634 2.2505
R25482 VDD.n3636 VDD.n2743 2.2505
R25483 VDD.n3638 VDD.n3637 2.2505
R25484 VDD.n3639 VDD.n2742 2.2505
R25485 VDD.n3641 VDD.n3640 2.2505
R25486 VDD.n3642 VDD.n2741 2.2505
R25487 VDD.n3644 VDD.n3643 2.2505
R25488 VDD.n3645 VDD.n2740 2.2505
R25489 VDD.n3647 VDD.n3646 2.2505
R25490 VDD.n3648 VDD.n2739 2.2505
R25491 VDD.n3650 VDD.n3649 2.2505
R25492 VDD.n3651 VDD.n2738 2.2505
R25493 VDD.n3653 VDD.n3652 2.2505
R25494 VDD.n3654 VDD.n2737 2.2505
R25495 VDD.n3656 VDD.n3655 2.2505
R25496 VDD.n3657 VDD.n2736 2.2505
R25497 VDD.n3659 VDD.n3658 2.2505
R25498 VDD.n3660 VDD.n2735 2.2505
R25499 VDD.n3662 VDD.n3661 2.2505
R25500 VDD.n3663 VDD.n2734 2.2505
R25501 VDD.n3665 VDD.n3664 2.2505
R25502 VDD.n3666 VDD.n2733 2.2505
R25503 VDD.n3668 VDD.n3667 2.2505
R25504 VDD.n3669 VDD.n2732 2.2505
R25505 VDD.n3671 VDD.n3670 2.2505
R25506 VDD.n3672 VDD.n2731 2.2505
R25507 VDD.n3674 VDD.n3673 2.2505
R25508 VDD.n3675 VDD.n2730 2.2505
R25509 VDD.n3677 VDD.n3676 2.2505
R25510 VDD.n3678 VDD.n2729 2.2505
R25511 VDD.n3680 VDD.n3679 2.2505
R25512 VDD.n3681 VDD.n2728 2.2505
R25513 VDD.n3683 VDD.n3682 2.2505
R25514 VDD.n3684 VDD.n2727 2.2505
R25515 VDD.n3686 VDD.n3685 2.2505
R25516 VDD.n3687 VDD.n2726 2.2505
R25517 VDD.n3689 VDD.n3688 2.2505
R25518 VDD.n3690 VDD.n2725 2.2505
R25519 VDD.n3692 VDD.n3691 2.2505
R25520 VDD.n3693 VDD.n2724 2.2505
R25521 VDD.n3695 VDD.n3694 2.2505
R25522 VDD.n3696 VDD.n2723 2.2505
R25523 VDD.n3698 VDD.n3697 2.2505
R25524 VDD.n3699 VDD.n2722 2.2505
R25525 VDD.n3701 VDD.n3700 2.2505
R25526 VDD.n3702 VDD.n2721 2.2505
R25527 VDD.n3704 VDD.n3703 2.2505
R25528 VDD.n3705 VDD.n2720 2.2505
R25529 VDD.n3707 VDD.n3706 2.2505
R25530 VDD.n3708 VDD.n2719 2.2505
R25531 VDD.n3710 VDD.n3709 2.2505
R25532 VDD.n3711 VDD.n2718 2.2505
R25533 VDD.n3713 VDD.n3712 2.2505
R25534 VDD.n3714 VDD.n2717 2.2505
R25535 VDD.n3716 VDD.n3715 2.2505
R25536 VDD.n3717 VDD.n2716 2.2505
R25537 VDD.n3719 VDD.n3718 2.2505
R25538 VDD.n3720 VDD.n2715 2.2505
R25539 VDD.n3722 VDD.n3721 2.2505
R25540 VDD.n3723 VDD.n2714 2.2505
R25541 VDD.n3725 VDD.n3724 2.2505
R25542 VDD.n3726 VDD.n2713 2.2505
R25543 VDD.n3728 VDD.n3727 2.2505
R25544 VDD.n3729 VDD.n2712 2.2505
R25545 VDD.n3731 VDD.n3730 2.2505
R25546 VDD.n3732 VDD.n2711 2.2505
R25547 VDD.n3734 VDD.n3733 2.2505
R25548 VDD.n3735 VDD.n2710 2.2505
R25549 VDD.n3737 VDD.n3736 2.2505
R25550 VDD.n3738 VDD.n2709 2.2505
R25551 VDD.n3740 VDD.n3739 2.2505
R25552 VDD.n3741 VDD.n2708 2.2505
R25553 VDD.n3743 VDD.n3742 2.2505
R25554 VDD.n3744 VDD.n2707 2.2505
R25555 VDD.n3746 VDD.n3745 2.2505
R25556 VDD.n3747 VDD.n2706 2.2505
R25557 VDD.n3749 VDD.n3748 2.2505
R25558 VDD.n3750 VDD.n2705 2.2505
R25559 VDD.n3752 VDD.n3751 2.2505
R25560 VDD.n3753 VDD.n2704 2.2505
R25561 VDD.n3755 VDD.n3754 2.2505
R25562 VDD.n3756 VDD.n2703 2.2505
R25563 VDD.n3758 VDD.n3757 2.2505
R25564 VDD.n3759 VDD.n2702 2.2505
R25565 VDD.n3761 VDD.n3760 2.2505
R25566 VDD.n3762 VDD.n2701 2.2505
R25567 VDD.n3764 VDD.n3763 2.2505
R25568 VDD.n3765 VDD.n2700 2.2505
R25569 VDD.n3767 VDD.n3766 2.2505
R25570 VDD.n3768 VDD.n2699 2.2505
R25571 VDD.n3770 VDD.n3769 2.2505
R25572 VDD.n3771 VDD.n2698 2.2505
R25573 VDD.n3773 VDD.n3772 2.2505
R25574 VDD.n3774 VDD.n2697 2.2505
R25575 VDD.n3776 VDD.n3775 2.2505
R25576 VDD.n3777 VDD.n2696 2.2505
R25577 VDD.n3779 VDD.n3778 2.2505
R25578 VDD.n3780 VDD.n2695 2.2505
R25579 VDD.n3782 VDD.n3781 2.2505
R25580 VDD.n3783 VDD.n2694 2.2505
R25581 VDD.n3785 VDD.n3784 2.2505
R25582 VDD.n3786 VDD.n2693 2.2505
R25583 VDD.n3788 VDD.n3787 2.2505
R25584 VDD.n3789 VDD.n2692 2.2505
R25585 VDD.n3791 VDD.n3790 2.2505
R25586 VDD.n3792 VDD.n2691 2.2505
R25587 VDD.n3794 VDD.n3793 2.2505
R25588 VDD.n3795 VDD.n2690 2.2505
R25589 VDD.n3797 VDD.n3796 2.2505
R25590 VDD.n3798 VDD.n2689 2.2505
R25591 VDD.n3800 VDD.n3799 2.2505
R25592 VDD.n3801 VDD.n2688 2.2505
R25593 VDD.n3803 VDD.n3802 2.2505
R25594 VDD.n3804 VDD.n2687 2.2505
R25595 VDD.n3806 VDD.n3805 2.2505
R25596 VDD.n3807 VDD.n2686 2.2505
R25597 VDD.n3809 VDD.n3808 2.2505
R25598 VDD.n3810 VDD.n2685 2.2505
R25599 VDD.n3812 VDD.n3811 2.2505
R25600 VDD.n3813 VDD.n2684 2.2505
R25601 VDD.n3815 VDD.n3814 2.2505
R25602 VDD.n3816 VDD.n2683 2.2505
R25603 VDD.n3818 VDD.n3817 2.2505
R25604 VDD.n3819 VDD.n2682 2.2505
R25605 VDD.n3821 VDD.n3820 2.2505
R25606 VDD.n3822 VDD.n2681 2.2505
R25607 VDD.n3824 VDD.n3823 2.2505
R25608 VDD.n3825 VDD.n2680 2.2505
R25609 VDD.n3827 VDD.n3826 2.2505
R25610 VDD.n3828 VDD.n2679 2.2505
R25611 VDD.n3830 VDD.n3829 2.2505
R25612 VDD.n3831 VDD.n2678 2.2505
R25613 VDD.n3833 VDD.n3832 2.2505
R25614 VDD.n3834 VDD.n2677 2.2505
R25615 VDD.n3836 VDD.n3835 2.2505
R25616 VDD.n3837 VDD.n2676 2.2505
R25617 VDD.n3839 VDD.n3838 2.2505
R25618 VDD.n3840 VDD.n2675 2.2505
R25619 VDD.n3842 VDD.n3841 2.2505
R25620 VDD.n3843 VDD.n2674 2.2505
R25621 VDD.n3845 VDD.n3844 2.2505
R25622 VDD.n3846 VDD.n2673 2.2505
R25623 VDD.n3848 VDD.n3847 2.2505
R25624 VDD.n3849 VDD.n2672 2.2505
R25625 VDD.n3851 VDD.n3850 2.2505
R25626 VDD.n3852 VDD.n2671 2.2505
R25627 VDD.n3854 VDD.n3853 2.2505
R25628 VDD.n3855 VDD.n2670 2.2505
R25629 VDD.n3857 VDD.n3856 2.2505
R25630 VDD.n3858 VDD.n2669 2.2505
R25631 VDD.n3860 VDD.n3859 2.2505
R25632 VDD.n3861 VDD.n2668 2.2505
R25633 VDD.n3863 VDD.n3862 2.2505
R25634 VDD.n3864 VDD.n2667 2.2505
R25635 VDD.n3866 VDD.n3865 2.2505
R25636 VDD.n3867 VDD.n2666 2.2505
R25637 VDD.n3869 VDD.n3868 2.2505
R25638 VDD.n3870 VDD.n2665 2.2505
R25639 VDD.n3872 VDD.n3871 2.2505
R25640 VDD.n3873 VDD.n2664 2.2505
R25641 VDD.n3875 VDD.n3874 2.2505
R25642 VDD.n3876 VDD.n2663 2.2505
R25643 VDD.n3878 VDD.n3877 2.2505
R25644 VDD.n3879 VDD.n2662 2.2505
R25645 VDD.n3881 VDD.n3880 2.2505
R25646 VDD.n3882 VDD.n2661 2.2505
R25647 VDD.n3884 VDD.n3883 2.2505
R25648 VDD.n3885 VDD.n2660 2.2505
R25649 VDD.n3887 VDD.n3886 2.2505
R25650 VDD.n3888 VDD.n2659 2.2505
R25651 VDD.n3890 VDD.n3889 2.2505
R25652 VDD.n3891 VDD.n2658 2.2505
R25653 VDD.n3893 VDD.n3892 2.2505
R25654 VDD.n3894 VDD.n2657 2.2505
R25655 VDD.n3896 VDD.n3895 2.2505
R25656 VDD.n3897 VDD.n2656 2.2505
R25657 VDD.n3899 VDD.n3898 2.2505
R25658 VDD.n3900 VDD.n2655 2.2505
R25659 VDD.n3902 VDD.n3901 2.2505
R25660 VDD.n3903 VDD.n2654 2.2505
R25661 VDD.n3905 VDD.n3904 2.2505
R25662 VDD.n3906 VDD.n2653 2.2505
R25663 VDD.n3908 VDD.n3907 2.2505
R25664 VDD.n3909 VDD.n2652 2.2505
R25665 VDD.n3911 VDD.n3910 2.2505
R25666 VDD.n3912 VDD.n2651 2.2505
R25667 VDD.n3914 VDD.n3913 2.2505
R25668 VDD.n3915 VDD.n2650 2.2505
R25669 VDD.n3917 VDD.n3916 2.2505
R25670 VDD.n3918 VDD.n2649 2.2505
R25671 VDD.n3920 VDD.n3919 2.2505
R25672 VDD.n3921 VDD.n2648 2.2505
R25673 VDD.n3923 VDD.n3922 2.2505
R25674 VDD.n3924 VDD.n2647 2.2505
R25675 VDD.n3926 VDD.n3925 2.2505
R25676 VDD.n3927 VDD.n2646 2.2505
R25677 VDD.n3929 VDD.n3928 2.2505
R25678 VDD.n3930 VDD.n2645 2.2505
R25679 VDD.n3932 VDD.n3931 2.2505
R25680 VDD.n3933 VDD.n2644 2.2505
R25681 VDD.n3935 VDD.n3934 2.2505
R25682 VDD.n3936 VDD.n2643 2.2505
R25683 VDD.n3938 VDD.n3937 2.2505
R25684 VDD.n3939 VDD.n2642 2.2505
R25685 VDD.n3941 VDD.n3940 2.2505
R25686 VDD.n3942 VDD.n2641 2.2505
R25687 VDD.n3944 VDD.n3943 2.2505
R25688 VDD.n3945 VDD.n2640 2.2505
R25689 VDD.n3947 VDD.n3946 2.2505
R25690 VDD.n3948 VDD.n2639 2.2505
R25691 VDD.n3950 VDD.n3949 2.2505
R25692 VDD.n3951 VDD.n2638 2.2505
R25693 VDD.n3953 VDD.n3952 2.2505
R25694 VDD.n3954 VDD.n2637 2.2505
R25695 VDD.n3956 VDD.n3955 2.2505
R25696 VDD.n3957 VDD.n2636 2.2505
R25697 VDD.n3959 VDD.n3958 2.2505
R25698 VDD.n3960 VDD.n2635 2.2505
R25699 VDD.n3962 VDD.n3961 2.2505
R25700 VDD.n3963 VDD.n2634 2.2505
R25701 VDD.n3965 VDD.n3964 2.2505
R25702 VDD.n3966 VDD.n2633 2.2505
R25703 VDD.n3968 VDD.n3967 2.2505
R25704 VDD.n3969 VDD.n2632 2.2505
R25705 VDD.n3971 VDD.n3970 2.2505
R25706 VDD.n3972 VDD.n2631 2.2505
R25707 VDD.n3974 VDD.n3973 2.2505
R25708 VDD.n3975 VDD.n2630 2.2505
R25709 VDD.n3977 VDD.n3976 2.2505
R25710 VDD.n3978 VDD.n2629 2.2505
R25711 VDD.n3980 VDD.n3979 2.2505
R25712 VDD.n3981 VDD.n2628 2.2505
R25713 VDD.n3983 VDD.n3982 2.2505
R25714 VDD.n3984 VDD.n2627 2.2505
R25715 VDD.n3986 VDD.n3985 2.2505
R25716 VDD.n3987 VDD.n2626 2.2505
R25717 VDD.n3989 VDD.n3988 2.2505
R25718 VDD.n3990 VDD.n2625 2.2505
R25719 VDD.n3992 VDD.n3991 2.2505
R25720 VDD.n3993 VDD.n2624 2.2505
R25721 VDD.n3995 VDD.n3994 2.2505
R25722 VDD.n3996 VDD.n2623 2.2505
R25723 VDD.n3998 VDD.n3997 2.2505
R25724 VDD.n3999 VDD.n2622 2.2505
R25725 VDD.n4001 VDD.n4000 2.2505
R25726 VDD.n4002 VDD.n2621 2.2505
R25727 VDD.n4004 VDD.n4003 2.2505
R25728 VDD.n4005 VDD.n2620 2.2505
R25729 VDD.n4007 VDD.n4006 2.2505
R25730 VDD.n4008 VDD.n2619 2.2505
R25731 VDD.n4010 VDD.n4009 2.2505
R25732 VDD.n4011 VDD.n2618 2.2505
R25733 VDD.n4013 VDD.n4012 2.2505
R25734 VDD.n4014 VDD.n2617 2.2505
R25735 VDD.n4016 VDD.n4015 2.2505
R25736 VDD.n4017 VDD.n2616 2.2505
R25737 VDD.n4019 VDD.n4018 2.2505
R25738 VDD.n4020 VDD.n2615 2.2505
R25739 VDD.n4022 VDD.n4021 2.2505
R25740 VDD.n4023 VDD.n2614 2.2505
R25741 VDD.n4025 VDD.n4024 2.2505
R25742 VDD.n4026 VDD.n2613 2.2505
R25743 VDD.n4028 VDD.n4027 2.2505
R25744 VDD.n4029 VDD.n2612 2.2505
R25745 VDD.n4031 VDD.n4030 2.2505
R25746 VDD.n4032 VDD.n2611 2.2505
R25747 VDD.n4034 VDD.n4033 2.2505
R25748 VDD.n4035 VDD.n2610 2.2505
R25749 VDD.n4037 VDD.n4036 2.2505
R25750 VDD.n4038 VDD.n2609 2.2505
R25751 VDD.n4040 VDD.n4039 2.2505
R25752 VDD.n4041 VDD.n2608 2.2505
R25753 VDD.n4043 VDD.n4042 2.2505
R25754 VDD.n4044 VDD.n2607 2.2505
R25755 VDD.n4046 VDD.n4045 2.2505
R25756 VDD.n4047 VDD.n2606 2.2505
R25757 VDD.n4049 VDD.n4048 2.2505
R25758 VDD.n4050 VDD.n2605 2.2505
R25759 VDD.n4052 VDD.n4051 2.2505
R25760 VDD.n4053 VDD.n2604 2.2505
R25761 VDD.n4055 VDD.n4054 2.2505
R25762 VDD.n4056 VDD.n2603 2.2505
R25763 VDD.n4058 VDD.n4057 2.2505
R25764 VDD.n4059 VDD.n2602 2.2505
R25765 VDD.n4061 VDD.n4060 2.2505
R25766 VDD.n4062 VDD.n2601 2.2505
R25767 VDD.n4064 VDD.n4063 2.2505
R25768 VDD.n4065 VDD.n2600 2.2505
R25769 VDD.n4067 VDD.n4066 2.2505
R25770 VDD.n4068 VDD.n2599 2.2505
R25771 VDD.n4070 VDD.n4069 2.2505
R25772 VDD.n4071 VDD.n2598 2.2505
R25773 VDD.n4073 VDD.n4072 2.2505
R25774 VDD.n4074 VDD.n2597 2.2505
R25775 VDD.n4076 VDD.n4075 2.2505
R25776 VDD.n4077 VDD.n2596 2.2505
R25777 VDD.n4079 VDD.n4078 2.2505
R25778 VDD.n4080 VDD.n2595 2.2505
R25779 VDD.n4082 VDD.n4081 2.2505
R25780 VDD.n4083 VDD.n2594 2.2505
R25781 VDD.n4085 VDD.n4084 2.2505
R25782 VDD.n4086 VDD.n2593 2.2505
R25783 VDD.n4088 VDD.n4087 2.2505
R25784 VDD.n4089 VDD.n2592 2.2505
R25785 VDD.n4091 VDD.n4090 2.2505
R25786 VDD.n4092 VDD.n2591 2.2505
R25787 VDD.n4094 VDD.n4093 2.2505
R25788 VDD.n4095 VDD.n2590 2.2505
R25789 VDD.n4097 VDD.n4096 2.2505
R25790 VDD.n4098 VDD.n2589 2.2505
R25791 VDD.n4100 VDD.n4099 2.2505
R25792 VDD.n4101 VDD.n2588 2.2505
R25793 VDD.n4103 VDD.n4102 2.2505
R25794 VDD.n4104 VDD.n2587 2.2505
R25795 VDD.n4106 VDD.n4105 2.2505
R25796 VDD.n4107 VDD.n2586 2.2505
R25797 VDD.n4109 VDD.n4108 2.2505
R25798 VDD.n4110 VDD.n2585 2.2505
R25799 VDD.n4112 VDD.n4111 2.2505
R25800 VDD.n4113 VDD.n2584 2.2505
R25801 VDD.n4115 VDD.n4114 2.2505
R25802 VDD.n4116 VDD.n2583 2.2505
R25803 VDD.n4118 VDD.n4117 2.2505
R25804 VDD.n4119 VDD.n2582 2.2505
R25805 VDD.n4121 VDD.n4120 2.2505
R25806 VDD.n4122 VDD.n2581 2.2505
R25807 VDD.n4124 VDD.n4123 2.2505
R25808 VDD.n4125 VDD.n2580 2.2505
R25809 VDD.n4127 VDD.n4126 2.2505
R25810 VDD.n4128 VDD.n2579 2.2505
R25811 VDD.n4130 VDD.n4129 2.2505
R25812 VDD.n4131 VDD.n2578 2.2505
R25813 VDD.n4133 VDD.n4132 2.2505
R25814 VDD.n4134 VDD.n2577 2.2505
R25815 VDD.n4136 VDD.n4135 2.2505
R25816 VDD.n4137 VDD.n2576 2.2505
R25817 VDD.n4139 VDD.n4138 2.2505
R25818 VDD.n4140 VDD.n2575 2.2505
R25819 VDD.n4142 VDD.n4141 2.2505
R25820 VDD.n4143 VDD.n2574 2.2505
R25821 VDD.n4145 VDD.n4144 2.2505
R25822 VDD.n4146 VDD.n2573 2.2505
R25823 VDD.n4148 VDD.n4147 2.2505
R25824 VDD.n4149 VDD.n2572 2.2505
R25825 VDD.n4151 VDD.n4150 2.2505
R25826 VDD.n4152 VDD.n2571 2.2505
R25827 VDD.n4154 VDD.n4153 2.2505
R25828 VDD.n4155 VDD.n2570 2.2505
R25829 VDD.n4157 VDD.n4156 2.2505
R25830 VDD.n4158 VDD.n2569 2.2505
R25831 VDD.n4160 VDD.n4159 2.2505
R25832 VDD.n4161 VDD.n2568 2.2505
R25833 VDD.n4163 VDD.n4162 2.2505
R25834 VDD.n4164 VDD.n2567 2.2505
R25835 VDD.n4166 VDD.n4165 2.2505
R25836 VDD.n4167 VDD.n2566 2.2505
R25837 VDD.n4169 VDD.n4168 2.2505
R25838 VDD.n4170 VDD.n2565 2.2505
R25839 VDD.n4172 VDD.n4171 2.2505
R25840 VDD.n4173 VDD.n2564 2.2505
R25841 VDD.n4175 VDD.n4174 2.2505
R25842 VDD.n4176 VDD.n2563 2.2505
R25843 VDD.n4178 VDD.n4177 2.2505
R25844 VDD.n4179 VDD.n2562 2.2505
R25845 VDD.n4181 VDD.n4180 2.2505
R25846 VDD.n4182 VDD.n2561 2.2505
R25847 VDD.n4184 VDD.n4183 2.2505
R25848 VDD.n4185 VDD.n2560 2.2505
R25849 VDD.n4187 VDD.n4186 2.2505
R25850 VDD.n4188 VDD.n2559 2.2505
R25851 VDD.n4190 VDD.n4189 2.2505
R25852 VDD.n4191 VDD.n2558 2.2505
R25853 VDD.n4193 VDD.n4192 2.2505
R25854 VDD.n4194 VDD.n2557 2.2505
R25855 VDD.n4196 VDD.n4195 2.2505
R25856 VDD.n4197 VDD.n2556 2.2505
R25857 VDD.n4199 VDD.n4198 2.2505
R25858 VDD.n4200 VDD.n2555 2.2505
R25859 VDD.n4202 VDD.n4201 2.2505
R25860 VDD.n4203 VDD.n2554 2.2505
R25861 VDD.n4205 VDD.n4204 2.2505
R25862 VDD.n4206 VDD.n2553 2.2505
R25863 VDD.n4208 VDD.n4207 2.2505
R25864 VDD.n4209 VDD.n2552 2.2505
R25865 VDD.n4211 VDD.n4210 2.2505
R25866 VDD.n4212 VDD.n2551 2.2505
R25867 VDD.n4214 VDD.n4213 2.2505
R25868 VDD.n4215 VDD.n2550 2.2505
R25869 VDD.n4217 VDD.n4216 2.2505
R25870 VDD.n4218 VDD.n2549 2.2505
R25871 VDD.n4220 VDD.n4219 2.2505
R25872 VDD.n4221 VDD.n2548 2.2505
R25873 VDD.n4223 VDD.n4222 2.2505
R25874 VDD.n4224 VDD.n2547 2.2505
R25875 VDD.n4226 VDD.n4225 2.2505
R25876 VDD.n4227 VDD.n2546 2.2505
R25877 VDD.n4229 VDD.n4228 2.2505
R25878 VDD.n4230 VDD.n2545 2.2505
R25879 VDD.n4232 VDD.n4231 2.2505
R25880 VDD.n4233 VDD.n2544 2.2505
R25881 VDD.n4235 VDD.n4234 2.2505
R25882 VDD.n4236 VDD.n2543 2.2505
R25883 VDD.n4238 VDD.n4237 2.2505
R25884 VDD.n4239 VDD.n2542 2.2505
R25885 VDD.n4241 VDD.n4240 2.2505
R25886 VDD.n4242 VDD.n2541 2.2505
R25887 VDD.n4244 VDD.n4243 2.2505
R25888 VDD.n4245 VDD.n2540 2.2505
R25889 VDD.n4247 VDD.n4246 2.2505
R25890 VDD.n4248 VDD.n2539 2.2505
R25891 VDD.n4250 VDD.n4249 2.2505
R25892 VDD.n4251 VDD.n2538 2.2505
R25893 VDD.n4253 VDD.n4252 2.2505
R25894 VDD.n4254 VDD.n2537 2.2505
R25895 VDD.n4256 VDD.n4255 2.2505
R25896 VDD.n4257 VDD.n2536 2.2505
R25897 VDD.n4259 VDD.n4258 2.2505
R25898 VDD.n4260 VDD.n2535 2.2505
R25899 VDD.n4262 VDD.n4261 2.2505
R25900 VDD.n4263 VDD.n2534 2.2505
R25901 VDD.n4265 VDD.n4264 2.2505
R25902 VDD.n4266 VDD.n2533 2.2505
R25903 VDD.n4268 VDD.n4267 2.2505
R25904 VDD.n4269 VDD.n2532 2.2505
R25905 VDD.n4271 VDD.n4270 2.2505
R25906 VDD.n4272 VDD.n2531 2.2505
R25907 VDD.n4274 VDD.n4273 2.2505
R25908 VDD.n4275 VDD.n2530 2.2505
R25909 VDD.n4277 VDD.n4276 2.2505
R25910 VDD.n4278 VDD.n2529 2.2505
R25911 VDD.n4280 VDD.n4279 2.2505
R25912 VDD.n4281 VDD.n2528 2.2505
R25913 VDD.n4283 VDD.n4282 2.2505
R25914 VDD.n4284 VDD.n2527 2.2505
R25915 VDD.n4286 VDD.n4285 2.2505
R25916 VDD.n4287 VDD.n2526 2.2505
R25917 VDD.n4289 VDD.n4288 2.2505
R25918 VDD.n4290 VDD.n2525 2.2505
R25919 VDD.n4292 VDD.n4291 2.2505
R25920 VDD.n4293 VDD.n2524 2.2505
R25921 VDD.n4295 VDD.n4294 2.2505
R25922 VDD.n4296 VDD.n2523 2.2505
R25923 VDD.n4298 VDD.n4297 2.2505
R25924 VDD.n4299 VDD.n2522 2.2505
R25925 VDD.n4301 VDD.n4300 2.2505
R25926 VDD.n4302 VDD.n2521 2.2505
R25927 VDD.n4304 VDD.n4303 2.2505
R25928 VDD.n4305 VDD.n2520 2.2505
R25929 VDD.n4307 VDD.n4306 2.2505
R25930 VDD.n4308 VDD.n2519 2.2505
R25931 VDD.n4310 VDD.n4309 2.2505
R25932 VDD.n4311 VDD.n2518 2.2505
R25933 VDD.n4313 VDD.n4312 2.2505
R25934 VDD.n4314 VDD.n2517 2.2505
R25935 VDD.n4316 VDD.n4315 2.2505
R25936 VDD.n4317 VDD.n2516 2.2505
R25937 VDD.n4319 VDD.n4318 2.2505
R25938 VDD.n4320 VDD.n2515 2.2505
R25939 VDD.n4322 VDD.n4321 2.2505
R25940 VDD.n4323 VDD.n2514 2.2505
R25941 VDD.n4325 VDD.n4324 2.2505
R25942 VDD.n4326 VDD.n2513 2.2505
R25943 VDD.n4328 VDD.n4327 2.2505
R25944 VDD.n4329 VDD.n2512 2.2505
R25945 VDD.n4331 VDD.n4330 2.2505
R25946 VDD.n4332 VDD.n2511 2.2505
R25947 VDD.n4334 VDD.n4333 2.2505
R25948 VDD.n4335 VDD.n2510 2.2505
R25949 VDD.n4337 VDD.n4336 2.2505
R25950 VDD.n4338 VDD.n2509 2.2505
R25951 VDD.n4340 VDD.n4339 2.2505
R25952 VDD.n4341 VDD.n2508 2.2505
R25953 VDD.n4343 VDD.n4342 2.2505
R25954 VDD.n4344 VDD.n2507 2.2505
R25955 VDD.n4346 VDD.n4345 2.2505
R25956 VDD.n4347 VDD.n2506 2.2505
R25957 VDD.n4349 VDD.n4348 2.2505
R25958 VDD.n4350 VDD.n2505 2.2505
R25959 VDD.n4352 VDD.n4351 2.2505
R25960 VDD.n4353 VDD.n2504 2.2505
R25961 VDD.n4355 VDD.n4354 2.2505
R25962 VDD.n4356 VDD.n2503 2.2505
R25963 VDD.n4358 VDD.n4357 2.2505
R25964 VDD.n4359 VDD.n2502 2.2505
R25965 VDD.n4361 VDD.n4360 2.2505
R25966 VDD.n4362 VDD.n2501 2.2505
R25967 VDD.n4364 VDD.n4363 2.2505
R25968 VDD.n4365 VDD.n2500 2.2505
R25969 VDD.n4367 VDD.n4366 2.2505
R25970 VDD.n4368 VDD.n2499 2.2505
R25971 VDD.n4370 VDD.n4369 2.2505
R25972 VDD.n4371 VDD.n2498 2.2505
R25973 VDD.n4373 VDD.n4372 2.2505
R25974 VDD.n4374 VDD.n2497 2.2505
R25975 VDD.n4376 VDD.n4375 2.2505
R25976 VDD.n4377 VDD.n2496 2.2505
R25977 VDD.n4379 VDD.n4378 2.2505
R25978 VDD.n4380 VDD.n2495 2.2505
R25979 VDD.n4382 VDD.n4381 2.2505
R25980 VDD.n4383 VDD.n2494 2.2505
R25981 VDD.n4385 VDD.n4384 2.2505
R25982 VDD.n4386 VDD.n2493 2.2505
R25983 VDD.n4388 VDD.n4387 2.2505
R25984 VDD.n4389 VDD.n2492 2.2505
R25985 VDD.n4391 VDD.n4390 2.2505
R25986 VDD.n4392 VDD.n2491 2.2505
R25987 VDD.n4394 VDD.n4393 2.2505
R25988 VDD.n4395 VDD.n2490 2.2505
R25989 VDD.n4397 VDD.n4396 2.2505
R25990 VDD.n4398 VDD.n2489 2.2505
R25991 VDD.n4400 VDD.n4399 2.2505
R25992 VDD.n4401 VDD.n2488 2.2505
R25993 VDD.n4403 VDD.n4402 2.2505
R25994 VDD.n4404 VDD.n2487 2.2505
R25995 VDD.n4406 VDD.n4405 2.2505
R25996 VDD.n4407 VDD.n2486 2.2505
R25997 VDD.n4409 VDD.n4408 2.2505
R25998 VDD.n4410 VDD.n2485 2.2505
R25999 VDD.n4412 VDD.n4411 2.2505
R26000 VDD.n4413 VDD.n2484 2.2505
R26001 VDD.n4415 VDD.n4414 2.2505
R26002 VDD.n4416 VDD.n2483 2.2505
R26003 VDD.n4418 VDD.n4417 2.2505
R26004 VDD.n4419 VDD.n2482 2.2505
R26005 VDD.n4421 VDD.n4420 2.2505
R26006 VDD.n4422 VDD.n2481 2.2505
R26007 VDD.n4424 VDD.n4423 2.2505
R26008 VDD.n4425 VDD.n2480 2.2505
R26009 VDD.n4427 VDD.n4426 2.2505
R26010 VDD.n4428 VDD.n2479 2.2505
R26011 VDD.n4430 VDD.n4429 2.2505
R26012 VDD.n4431 VDD.n2478 2.2505
R26013 VDD.n4433 VDD.n4432 2.2505
R26014 VDD.n4434 VDD.n2477 2.2505
R26015 VDD.n4436 VDD.n4435 2.2505
R26016 VDD.n4437 VDD.n2476 2.2505
R26017 VDD.n4439 VDD.n4438 2.2505
R26018 VDD.n4440 VDD.n2475 2.2505
R26019 VDD.n4442 VDD.n4441 2.2505
R26020 VDD.n4443 VDD.n2474 2.2505
R26021 VDD.n4445 VDD.n4444 2.2505
R26022 VDD.n4446 VDD.n2473 2.2505
R26023 VDD.n4448 VDD.n4447 2.2505
R26024 VDD.n4449 VDD.n2472 2.2505
R26025 VDD.n4451 VDD.n4450 2.2505
R26026 VDD.n4452 VDD.n2471 2.2505
R26027 VDD.n4454 VDD.n4453 2.2505
R26028 VDD.n4455 VDD.n2470 2.2505
R26029 VDD.n4457 VDD.n4456 2.2505
R26030 VDD.n4458 VDD.n2469 2.2505
R26031 VDD.n4460 VDD.n4459 2.2505
R26032 VDD.n4461 VDD.n2468 2.2505
R26033 VDD.n4463 VDD.n4462 2.2505
R26034 VDD.n4464 VDD.n2467 2.2505
R26035 VDD.n4466 VDD.n4465 2.2505
R26036 VDD.n4467 VDD.n2466 2.2505
R26037 VDD.n4469 VDD.n4468 2.2505
R26038 VDD.n4470 VDD.n2465 2.2505
R26039 VDD.n4472 VDD.n4471 2.2505
R26040 VDD.n4473 VDD.n2464 2.2505
R26041 VDD.n4475 VDD.n4474 2.2505
R26042 VDD.n4476 VDD.n2463 2.2505
R26043 VDD.n4478 VDD.n4477 2.2505
R26044 VDD.n4479 VDD.n2462 2.2505
R26045 VDD.n4481 VDD.n4480 2.2505
R26046 VDD.n4482 VDD.n2461 2.2505
R26047 VDD.n4484 VDD.n4483 2.2505
R26048 VDD.n4485 VDD.n2460 2.2505
R26049 VDD.n4487 VDD.n4486 2.2505
R26050 VDD.n4488 VDD.n2459 2.2505
R26051 VDD.n4490 VDD.n4489 2.2505
R26052 VDD.n4491 VDD.n2458 2.2505
R26053 VDD.n4493 VDD.n4492 2.2505
R26054 VDD.n4494 VDD.n2457 2.2505
R26055 VDD.n4496 VDD.n4495 2.2505
R26056 VDD.n4497 VDD.n2456 2.2505
R26057 VDD.n4499 VDD.n4498 2.2505
R26058 VDD.n4500 VDD.n2455 2.2505
R26059 VDD.n4502 VDD.n4501 2.2505
R26060 VDD.n4503 VDD.n2454 2.2505
R26061 VDD.n4505 VDD.n4504 2.2505
R26062 VDD.n4506 VDD.n2453 2.2505
R26063 VDD.n4508 VDD.n4507 2.2505
R26064 VDD.n4509 VDD.n2452 2.2505
R26065 VDD.n4511 VDD.n4510 2.2505
R26066 VDD.n4512 VDD.n2451 2.2505
R26067 VDD.n4514 VDD.n4513 2.2505
R26068 VDD.n4515 VDD.n2450 2.2505
R26069 VDD.n4517 VDD.n4516 2.2505
R26070 VDD.n4518 VDD.n2449 2.2505
R26071 VDD.n4520 VDD.n4519 2.2505
R26072 VDD.n4521 VDD.n2448 2.2505
R26073 VDD.n4523 VDD.n4522 2.2505
R26074 VDD.n4524 VDD.n2447 2.2505
R26075 VDD.n4526 VDD.n4525 2.2505
R26076 VDD.n4527 VDD.n2446 2.2505
R26077 VDD.n4529 VDD.n4528 2.2505
R26078 VDD.n4530 VDD.n2445 2.2505
R26079 VDD.n4532 VDD.n4531 2.2505
R26080 VDD.n4533 VDD.n2444 2.2505
R26081 VDD.n4535 VDD.n4534 2.2505
R26082 VDD.n4536 VDD.n2443 2.2505
R26083 VDD.n4538 VDD.n4537 2.2505
R26084 VDD.n4539 VDD.n2442 2.2505
R26085 VDD.n4541 VDD.n4540 2.2505
R26086 VDD.n4542 VDD.n2441 2.2505
R26087 VDD.n4544 VDD.n4543 2.2505
R26088 VDD.n4545 VDD.n2440 2.2505
R26089 VDD.n4547 VDD.n4546 2.2505
R26090 VDD.n4548 VDD.n2439 2.2505
R26091 VDD.n4550 VDD.n4549 2.2505
R26092 VDD.n4551 VDD.n2438 2.2505
R26093 VDD.n4553 VDD.n4552 2.2505
R26094 VDD.n4554 VDD.n2437 2.2505
R26095 VDD.n4556 VDD.n4555 2.2505
R26096 VDD.n4557 VDD.n2436 2.2505
R26097 VDD.n4559 VDD.n4558 2.2505
R26098 VDD.n4560 VDD.n2435 2.2505
R26099 VDD.n4562 VDD.n4561 2.2505
R26100 VDD.n4563 VDD.n2434 2.2505
R26101 VDD.n4565 VDD.n4564 2.2505
R26102 VDD.n4566 VDD.n2433 2.2505
R26103 VDD.n4568 VDD.n4567 2.2505
R26104 VDD.n4569 VDD.n2432 2.2505
R26105 VDD.n4571 VDD.n4570 2.2505
R26106 VDD.n4572 VDD.n2431 2.2505
R26107 VDD.n4574 VDD.n4573 2.2505
R26108 VDD.n4575 VDD.n2430 2.2505
R26109 VDD.n4577 VDD.n4576 2.2505
R26110 VDD.n4578 VDD.n2429 2.2505
R26111 VDD.n4580 VDD.n4579 2.2505
R26112 VDD.n4581 VDD.n2428 2.2505
R26113 VDD.n4583 VDD.n4582 2.2505
R26114 VDD.n4584 VDD.n2427 2.2505
R26115 VDD.n4586 VDD.n4585 2.2505
R26116 VDD.n4587 VDD.n2426 2.2505
R26117 VDD.n4589 VDD.n4588 2.2505
R26118 VDD.n5200 VDD.n5199 2.2505
R26119 VDD.n5198 VDD.n4598 2.2505
R26120 VDD.n5197 VDD.n5196 2.2505
R26121 VDD.n5195 VDD.n4600 2.2505
R26122 VDD.n5194 VDD.n5193 2.2505
R26123 VDD.n5192 VDD.n4601 2.2505
R26124 VDD.n5191 VDD.n5190 2.2505
R26125 VDD.n5189 VDD.n4602 2.2505
R26126 VDD.n5188 VDD.n5187 2.2505
R26127 VDD.n5186 VDD.n4603 2.2505
R26128 VDD.n5185 VDD.n5184 2.2505
R26129 VDD.n5183 VDD.n4604 2.2505
R26130 VDD.n5182 VDD.n5181 2.2505
R26131 VDD.n5180 VDD.n4605 2.2505
R26132 VDD.n5179 VDD.n5178 2.2505
R26133 VDD.n5177 VDD.n4606 2.2505
R26134 VDD.n5176 VDD.n5175 2.2505
R26135 VDD.n5174 VDD.n4607 2.2505
R26136 VDD.n5173 VDD.n5172 2.2505
R26137 VDD.n5171 VDD.n4608 2.2505
R26138 VDD.n5170 VDD.n5169 2.2505
R26139 VDD.n5168 VDD.n4609 2.2505
R26140 VDD.n5167 VDD.n5166 2.2505
R26141 VDD.n5165 VDD.n4610 2.2505
R26142 VDD.n5164 VDD.n5163 2.2505
R26143 VDD.n5162 VDD.n4611 2.2505
R26144 VDD.n5161 VDD.n5160 2.2505
R26145 VDD.n5159 VDD.n4612 2.2505
R26146 VDD.n5158 VDD.n5157 2.2505
R26147 VDD.n5156 VDD.n4613 2.2505
R26148 VDD.n5155 VDD.n5154 2.2505
R26149 VDD.n5153 VDD.n4614 2.2505
R26150 VDD.n5152 VDD.n5151 2.2505
R26151 VDD.n5150 VDD.n4615 2.2505
R26152 VDD.n5149 VDD.n5148 2.2505
R26153 VDD.n5147 VDD.n4616 2.2505
R26154 VDD.n5146 VDD.n5145 2.2505
R26155 VDD.n5144 VDD.n4617 2.2505
R26156 VDD.n5143 VDD.n5142 2.2505
R26157 VDD.n5141 VDD.n4618 2.2505
R26158 VDD.n5140 VDD.n5139 2.2505
R26159 VDD.n5138 VDD.n4619 2.2505
R26160 VDD.n5137 VDD.n5136 2.2505
R26161 VDD.n5135 VDD.n4620 2.2505
R26162 VDD.n5134 VDD.n5133 2.2505
R26163 VDD.n5132 VDD.n4621 2.2505
R26164 VDD.n5131 VDD.n5130 2.2505
R26165 VDD.n5129 VDD.n4622 2.2505
R26166 VDD.n5128 VDD.n5127 2.2505
R26167 VDD.n5126 VDD.n4623 2.2505
R26168 VDD.n5125 VDD.n5124 2.2505
R26169 VDD.n5123 VDD.n4624 2.2505
R26170 VDD.n5122 VDD.n5121 2.2505
R26171 VDD.n5120 VDD.n4625 2.2505
R26172 VDD.n5119 VDD.n5118 2.2505
R26173 VDD.n5117 VDD.n4626 2.2505
R26174 VDD.n5116 VDD.n5115 2.2505
R26175 VDD.n5114 VDD.n4627 2.2505
R26176 VDD.n5113 VDD.n5112 2.2505
R26177 VDD.n5111 VDD.n4628 2.2505
R26178 VDD.n5110 VDD.n5109 2.2505
R26179 VDD.n5108 VDD.n4629 2.2505
R26180 VDD.n5107 VDD.n5106 2.2505
R26181 VDD.n5105 VDD.n4630 2.2505
R26182 VDD.n5104 VDD.n5103 2.2505
R26183 VDD.n5102 VDD.n4631 2.2505
R26184 VDD.n5101 VDD.n5100 2.2505
R26185 VDD.n5099 VDD.n4632 2.2505
R26186 VDD.n5098 VDD.n5097 2.2505
R26187 VDD.n5096 VDD.n4633 2.2505
R26188 VDD.n5095 VDD.n5094 2.2505
R26189 VDD.n5093 VDD.n4634 2.2505
R26190 VDD.n5092 VDD.n5091 2.2505
R26191 VDD.n5090 VDD.n4635 2.2505
R26192 VDD.n5089 VDD.n5088 2.2505
R26193 VDD.n5087 VDD.n4636 2.2505
R26194 VDD.n5086 VDD.n5085 2.2505
R26195 VDD.n5084 VDD.n4637 2.2505
R26196 VDD.n5083 VDD.n5082 2.2505
R26197 VDD.n5081 VDD.n4638 2.2505
R26198 VDD.n5080 VDD.n5079 2.2505
R26199 VDD.n5078 VDD.n4639 2.2505
R26200 VDD.n5077 VDD.n5076 2.2505
R26201 VDD.n5075 VDD.n4640 2.2505
R26202 VDD.n5074 VDD.n5073 2.2505
R26203 VDD.n5072 VDD.n4641 2.2505
R26204 VDD.n5071 VDD.n5070 2.2505
R26205 VDD.n5069 VDD.n4642 2.2505
R26206 VDD.n5068 VDD.n5067 2.2505
R26207 VDD.n5066 VDD.n4643 2.2505
R26208 VDD.n5065 VDD.n5064 2.2505
R26209 VDD.n5063 VDD.n4644 2.2505
R26210 VDD.n5062 VDD.n5061 2.2505
R26211 VDD.n5060 VDD.n4645 2.2505
R26212 VDD.n5059 VDD.n5058 2.2505
R26213 VDD.n5057 VDD.n4646 2.2505
R26214 VDD.n5056 VDD.n5055 2.2505
R26215 VDD.n5054 VDD.n4647 2.2505
R26216 VDD.n5053 VDD.n5052 2.2505
R26217 VDD.n5051 VDD.n4648 2.2505
R26218 VDD.n5050 VDD.n5049 2.2505
R26219 VDD.n5048 VDD.n4649 2.2505
R26220 VDD.n5047 VDD.n5046 2.2505
R26221 VDD.n5045 VDD.n4650 2.2505
R26222 VDD.n5044 VDD.n5043 2.2505
R26223 VDD.n5042 VDD.n4651 2.2505
R26224 VDD.n5041 VDD.n5040 2.2505
R26225 VDD.n5039 VDD.n4652 2.2505
R26226 VDD.n5038 VDD.n5037 2.2505
R26227 VDD.n5036 VDD.n4653 2.2505
R26228 VDD.n5035 VDD.n5034 2.2505
R26229 VDD.n5033 VDD.n4654 2.2505
R26230 VDD.n5032 VDD.n5031 2.2505
R26231 VDD.n5030 VDD.n4655 2.2505
R26232 VDD.n5029 VDD.n5028 2.2505
R26233 VDD.n5027 VDD.n4656 2.2505
R26234 VDD.n5026 VDD.n5025 2.2505
R26235 VDD.n5024 VDD.n4657 2.2505
R26236 VDD.n5023 VDD.n5022 2.2505
R26237 VDD.n5021 VDD.n4658 2.2505
R26238 VDD.n5020 VDD.n5019 2.2505
R26239 VDD.n5018 VDD.n4659 2.2505
R26240 VDD.n5017 VDD.n5016 2.2505
R26241 VDD.n5015 VDD.n4660 2.2505
R26242 VDD.n5014 VDD.n5013 2.2505
R26243 VDD.n5012 VDD.n4661 2.2505
R26244 VDD.n5011 VDD.n5010 2.2505
R26245 VDD.n5009 VDD.n4662 2.2505
R26246 VDD.n5008 VDD.n5007 2.2505
R26247 VDD.n5006 VDD.n4663 2.2505
R26248 VDD.n5005 VDD.n5004 2.2505
R26249 VDD.n5003 VDD.n4664 2.2505
R26250 VDD.n5002 VDD.n5001 2.2505
R26251 VDD.n5000 VDD.n4665 2.2505
R26252 VDD.n4999 VDD.n4998 2.2505
R26253 VDD.n4997 VDD.n4666 2.2505
R26254 VDD.n4996 VDD.n4995 2.2505
R26255 VDD.n4994 VDD.n4667 2.2505
R26256 VDD.n4993 VDD.n4992 2.2505
R26257 VDD.n4991 VDD.n4668 2.2505
R26258 VDD.n4990 VDD.n4989 2.2505
R26259 VDD.n4988 VDD.n4669 2.2505
R26260 VDD.n4987 VDD.n4986 2.2505
R26261 VDD.n4985 VDD.n4670 2.2505
R26262 VDD.n4984 VDD.n4983 2.2505
R26263 VDD.n4982 VDD.n4671 2.2505
R26264 VDD.n4981 VDD.n4980 2.2505
R26265 VDD.n4979 VDD.n4672 2.2505
R26266 VDD.n4978 VDD.n4977 2.2505
R26267 VDD.n4976 VDD.n4673 2.2505
R26268 VDD.n4975 VDD.n4974 2.2505
R26269 VDD.n4973 VDD.n4674 2.2505
R26270 VDD.n4972 VDD.n4971 2.2505
R26271 VDD.n4970 VDD.n4675 2.2505
R26272 VDD.n4969 VDD.n4968 2.2505
R26273 VDD.n4967 VDD.n4676 2.2505
R26274 VDD.n4966 VDD.n4965 2.2505
R26275 VDD.n4964 VDD.n4677 2.2505
R26276 VDD.n4963 VDD.n4962 2.2505
R26277 VDD.n4961 VDD.n4678 2.2505
R26278 VDD.n4960 VDD.n4959 2.2505
R26279 VDD.n4958 VDD.n4679 2.2505
R26280 VDD.n4957 VDD.n4956 2.2505
R26281 VDD.n4955 VDD.n4680 2.2505
R26282 VDD.n4954 VDD.n4953 2.2505
R26283 VDD.n4952 VDD.n4681 2.2505
R26284 VDD.n4951 VDD.n4950 2.2505
R26285 VDD.n4949 VDD.n4682 2.2505
R26286 VDD.n4948 VDD.n4947 2.2505
R26287 VDD.n4946 VDD.n4683 2.2505
R26288 VDD.n4945 VDD.n4944 2.2505
R26289 VDD.n4943 VDD.n4684 2.2505
R26290 VDD.n4942 VDD.n4941 2.2505
R26291 VDD.n4940 VDD.n4685 2.2505
R26292 VDD.n4939 VDD.n4938 2.2505
R26293 VDD.n4937 VDD.n4686 2.2505
R26294 VDD.n4936 VDD.n4935 2.2505
R26295 VDD.n4934 VDD.n4687 2.2505
R26296 VDD.n4933 VDD.n4932 2.2505
R26297 VDD.n4931 VDD.n4688 2.2505
R26298 VDD.n4930 VDD.n4929 2.2505
R26299 VDD.n4928 VDD.n4689 2.2505
R26300 VDD.n4927 VDD.n4926 2.2505
R26301 VDD.n4925 VDD.n4690 2.2505
R26302 VDD.n4924 VDD.n4923 2.2505
R26303 VDD.n4922 VDD.n4691 2.2505
R26304 VDD.n4921 VDD.n4920 2.2505
R26305 VDD.n4919 VDD.n4692 2.2505
R26306 VDD.n4918 VDD.n4917 2.2505
R26307 VDD.n4916 VDD.n4693 2.2505
R26308 VDD.n4915 VDD.n4914 2.2505
R26309 VDD.n4913 VDD.n4694 2.2505
R26310 VDD.n4912 VDD.n4911 2.2505
R26311 VDD.n4910 VDD.n4695 2.2505
R26312 VDD.n4909 VDD.n4908 2.2505
R26313 VDD.n4907 VDD.n4696 2.2505
R26314 VDD.n4906 VDD.n4905 2.2505
R26315 VDD.n1768 VDD.n1767 2.2505
R26316 VDD.n11039 VDD.n11038 2.2505
R26317 VDD.n11043 VDD.n11042 2.2505
R26318 VDD.n11041 VDD.n673 2.2505
R26319 VDD.n11040 VDD.n676 2.2505
R26320 VDD.n11049 VDD.n668 2.2505
R26321 VDD.n11051 VDD.n11050 2.2505
R26322 VDD.n11052 VDD.n667 2.2505
R26323 VDD.n11054 VDD.n11053 2.2505
R26324 VDD.n11055 VDD.n666 2.2505
R26325 VDD.n11059 VDD.n11058 2.2505
R26326 VDD.n11060 VDD.n665 2.2505
R26327 VDD.n11062 VDD.n11061 2.2505
R26328 VDD.n11064 VDD.n664 2.2505
R26329 VDD.n11066 VDD.n11065 2.2505
R26330 VDD.n11067 VDD.n663 2.2505
R26331 VDD.n11069 VDD.n11068 2.2505
R26332 VDD.n11070 VDD.n662 2.2505
R26333 VDD.n11072 VDD.n11071 2.2505
R26334 VDD.n11074 VDD.n11073 2.2505
R26335 VDD.n11075 VDD.n660 2.2505
R26336 VDD.n11079 VDD.n11078 2.2505
R26337 VDD.n11080 VDD.n659 2.2505
R26338 VDD.n11082 VDD.n11081 2.2505
R26339 VDD.n11083 VDD.n658 2.2505
R26340 VDD.n11085 VDD.n11084 2.2505
R26341 VDD.n11087 VDD.n11086 2.2505
R26342 VDD.n11088 VDD.n656 2.2505
R26343 VDD.n11092 VDD.n11091 2.2505
R26344 VDD.n11093 VDD.n655 2.2505
R26345 VDD.n11095 VDD.n11094 2.2505
R26346 VDD.n11096 VDD.n654 2.2505
R26347 VDD.n11099 VDD.n11098 2.2505
R26348 VDD.n11100 VDD.n653 2.2505
R26349 VDD.n11102 VDD.n11101 2.2505
R26350 VDD.n11103 VDD.n652 2.2505
R26351 VDD.n11105 VDD.n11104 2.2505
R26352 VDD.n11107 VDD.n11106 2.2505
R26353 VDD.n11108 VDD.n650 2.2505
R26354 VDD.n11110 VDD.n11109 2.2505
R26355 VDD.n11112 VDD.n11111 2.2505
R26356 VDD.n11113 VDD.n647 2.2505
R26357 VDD.n11115 VDD.n11114 2.2505
R26358 VDD.n11116 VDD.n646 2.2505
R26359 VDD.n11118 VDD.n11117 2.2505
R26360 VDD.n11120 VDD.n645 2.2505
R26361 VDD.n11122 VDD.n11121 2.2505
R26362 VDD.n11124 VDD.n11123 2.2505
R26363 VDD.n11126 VDD.n11125 2.2505
R26364 VDD.n633 VDD.n632 2.2505
R26365 VDD.n11132 VDD.n11131 2.2505
R26366 VDD.n11133 VDD.n631 2.2505
R26367 VDD.n3629 VDD.n3628 2.2505
R26368 VDD.n3627 VDD.n2746 2.2505
R26369 VDD.n3626 VDD.n3625 2.2505
R26370 VDD.n3624 VDD.n2747 2.2505
R26371 VDD.n3623 VDD.n3622 2.2505
R26372 VDD.n3621 VDD.n2748 2.2505
R26373 VDD.n3620 VDD.n3619 2.2505
R26374 VDD.n3618 VDD.n2749 2.2505
R26375 VDD.n3617 VDD.n3616 2.2505
R26376 VDD.n3615 VDD.n2750 2.2505
R26377 VDD.n3614 VDD.n3613 2.2505
R26378 VDD.n3612 VDD.n2751 2.2505
R26379 VDD.n3611 VDD.n3610 2.2505
R26380 VDD.n3609 VDD.n2752 2.2505
R26381 VDD.n3608 VDD.n3607 2.2505
R26382 VDD.n3606 VDD.n2753 2.2505
R26383 VDD.n3605 VDD.n3604 2.2505
R26384 VDD.n3603 VDD.n2754 2.2505
R26385 VDD.n3602 VDD.n3601 2.2505
R26386 VDD.n3600 VDD.n2755 2.2505
R26387 VDD.n3599 VDD.n3598 2.2505
R26388 VDD.n3597 VDD.n2756 2.2505
R26389 VDD.n3596 VDD.n3595 2.2505
R26390 VDD.n3594 VDD.n2757 2.2505
R26391 VDD.n3593 VDD.n3592 2.2505
R26392 VDD.n3591 VDD.n2758 2.2505
R26393 VDD.n3590 VDD.n3589 2.2505
R26394 VDD.n3588 VDD.n2759 2.2505
R26395 VDD.n3587 VDD.n3586 2.2505
R26396 VDD.n3585 VDD.n2760 2.2505
R26397 VDD.n3584 VDD.n3583 2.2505
R26398 VDD.n3582 VDD.n2761 2.2505
R26399 VDD.n3581 VDD.n3580 2.2505
R26400 VDD.n3579 VDD.n2762 2.2505
R26401 VDD.n3578 VDD.n3577 2.2505
R26402 VDD.n3576 VDD.n2763 2.2505
R26403 VDD.n3575 VDD.n3574 2.2505
R26404 VDD.n3573 VDD.n2764 2.2505
R26405 VDD.n3572 VDD.n3571 2.2505
R26406 VDD.n3570 VDD.n2765 2.2505
R26407 VDD.n3569 VDD.n3568 2.2505
R26408 VDD.n3567 VDD.n2766 2.2505
R26409 VDD.n3566 VDD.n3565 2.2505
R26410 VDD.n3564 VDD.n2767 2.2505
R26411 VDD.n3563 VDD.n3562 2.2505
R26412 VDD.n3561 VDD.n2768 2.2505
R26413 VDD.n3560 VDD.n3559 2.2505
R26414 VDD.n3558 VDD.n2769 2.2505
R26415 VDD.n3557 VDD.n3556 2.2505
R26416 VDD.n3555 VDD.n2770 2.2505
R26417 VDD.n3554 VDD.n3553 2.2505
R26418 VDD.n3552 VDD.n2771 2.2505
R26419 VDD.n3551 VDD.n3550 2.2505
R26420 VDD.n3549 VDD.n2772 2.2505
R26421 VDD.n3548 VDD.n3547 2.2505
R26422 VDD.n3546 VDD.n2773 2.2505
R26423 VDD.n3545 VDD.n3544 2.2505
R26424 VDD.n3543 VDD.n2774 2.2505
R26425 VDD.n3542 VDD.n3541 2.2505
R26426 VDD.n3540 VDD.n2775 2.2505
R26427 VDD.n3539 VDD.n3538 2.2505
R26428 VDD.n3537 VDD.n2776 2.2505
R26429 VDD.n3536 VDD.n3535 2.2505
R26430 VDD.n3534 VDD.n2777 2.2505
R26431 VDD.n3533 VDD.n3532 2.2505
R26432 VDD.n3531 VDD.n2778 2.2505
R26433 VDD.n3530 VDD.n3529 2.2505
R26434 VDD.n3528 VDD.n2779 2.2505
R26435 VDD.n3527 VDD.n3526 2.2505
R26436 VDD.n3525 VDD.n2780 2.2505
R26437 VDD.n3524 VDD.n3523 2.2505
R26438 VDD.n3522 VDD.n2781 2.2505
R26439 VDD.n3521 VDD.n3520 2.2505
R26440 VDD.n3519 VDD.n2782 2.2505
R26441 VDD.n3518 VDD.n3517 2.2505
R26442 VDD.n3516 VDD.n2783 2.2505
R26443 VDD.n3515 VDD.n3514 2.2505
R26444 VDD.n3513 VDD.n2784 2.2505
R26445 VDD.n3512 VDD.n3511 2.2505
R26446 VDD.n3510 VDD.n2785 2.2505
R26447 VDD.n3509 VDD.n3508 2.2505
R26448 VDD.n3507 VDD.n2786 2.2505
R26449 VDD.n3506 VDD.n3505 2.2505
R26450 VDD.n3504 VDD.n2787 2.2505
R26451 VDD.n3503 VDD.n3502 2.2505
R26452 VDD.n3501 VDD.n2788 2.2505
R26453 VDD.n3500 VDD.n3499 2.2505
R26454 VDD.n3498 VDD.n2789 2.2505
R26455 VDD.n3497 VDD.n3496 2.2505
R26456 VDD.n3495 VDD.n2790 2.2505
R26457 VDD.n3494 VDD.n3493 2.2505
R26458 VDD.n3492 VDD.n2791 2.2505
R26459 VDD.n3491 VDD.n3490 2.2505
R26460 VDD.n3489 VDD.n2792 2.2505
R26461 VDD.n3488 VDD.n3487 2.2505
R26462 VDD.n3486 VDD.n2793 2.2505
R26463 VDD.n3485 VDD.n3484 2.2505
R26464 VDD.n3483 VDD.n2794 2.2505
R26465 VDD.n3482 VDD.n3481 2.2505
R26466 VDD.n3480 VDD.n2795 2.2505
R26467 VDD.n3479 VDD.n3478 2.2505
R26468 VDD.n3477 VDD.n2796 2.2505
R26469 VDD.n3476 VDD.n3475 2.2505
R26470 VDD.n3474 VDD.n2797 2.2505
R26471 VDD.n3473 VDD.n3472 2.2505
R26472 VDD.n3471 VDD.n2798 2.2505
R26473 VDD.n3470 VDD.n3469 2.2505
R26474 VDD.n3468 VDD.n2799 2.2505
R26475 VDD.n3467 VDD.n3466 2.2505
R26476 VDD.n3465 VDD.n2800 2.2505
R26477 VDD.n3464 VDD.n3463 2.2505
R26478 VDD.n3462 VDD.n2801 2.2505
R26479 VDD.n3461 VDD.n3460 2.2505
R26480 VDD.n3459 VDD.n2802 2.2505
R26481 VDD.n3458 VDD.n3457 2.2505
R26482 VDD.n3456 VDD.n2803 2.2505
R26483 VDD.n3455 VDD.n3454 2.2505
R26484 VDD.n3453 VDD.n2804 2.2505
R26485 VDD.n3452 VDD.n3451 2.2505
R26486 VDD.n3450 VDD.n2805 2.2505
R26487 VDD.n3449 VDD.n3448 2.2505
R26488 VDD.n3447 VDD.n2806 2.2505
R26489 VDD.n3446 VDD.n3445 2.2505
R26490 VDD.n3444 VDD.n2807 2.2505
R26491 VDD.n3443 VDD.n3442 2.2505
R26492 VDD.n3441 VDD.n2808 2.2505
R26493 VDD.n3440 VDD.n3439 2.2505
R26494 VDD.n3438 VDD.n2809 2.2505
R26495 VDD.n3437 VDD.n3436 2.2505
R26496 VDD.n3435 VDD.n2810 2.2505
R26497 VDD.n3434 VDD.n3433 2.2505
R26498 VDD.n3432 VDD.n2811 2.2505
R26499 VDD.n3431 VDD.n3430 2.2505
R26500 VDD.n3429 VDD.n2812 2.2505
R26501 VDD.n3428 VDD.n3427 2.2505
R26502 VDD.n3426 VDD.n2813 2.2505
R26503 VDD.n3425 VDD.n3424 2.2505
R26504 VDD.n3423 VDD.n2814 2.2505
R26505 VDD.n3422 VDD.n3421 2.2505
R26506 VDD.n3420 VDD.n2815 2.2505
R26507 VDD.n3419 VDD.n3418 2.2505
R26508 VDD.n3417 VDD.n2816 2.2505
R26509 VDD.n3416 VDD.n3415 2.2505
R26510 VDD.n3414 VDD.n2817 2.2505
R26511 VDD.n3413 VDD.n3412 2.2505
R26512 VDD.n3411 VDD.n2818 2.2505
R26513 VDD.n3410 VDD.n3409 2.2505
R26514 VDD.n3408 VDD.n2819 2.2505
R26515 VDD.n3407 VDD.n3406 2.2505
R26516 VDD.n3405 VDD.n2820 2.2505
R26517 VDD.n3404 VDD.n3403 2.2505
R26518 VDD.n3402 VDD.n2821 2.2505
R26519 VDD.n3401 VDD.n3400 2.2505
R26520 VDD.n3399 VDD.n2822 2.2505
R26521 VDD.n3398 VDD.n3397 2.2505
R26522 VDD.n3396 VDD.n2823 2.2505
R26523 VDD.n3395 VDD.n3394 2.2505
R26524 VDD.n3393 VDD.n2824 2.2505
R26525 VDD.n3392 VDD.n3391 2.2505
R26526 VDD.n3390 VDD.n2825 2.2505
R26527 VDD.n3389 VDD.n3388 2.2505
R26528 VDD.n3387 VDD.n2826 2.2505
R26529 VDD.n3386 VDD.n3385 2.2505
R26530 VDD.n3384 VDD.n2827 2.2505
R26531 VDD.n3383 VDD.n3382 2.2505
R26532 VDD.n3381 VDD.n2828 2.2505
R26533 VDD.n3380 VDD.n3379 2.2505
R26534 VDD.n3378 VDD.n2829 2.2505
R26535 VDD.n3377 VDD.n3376 2.2505
R26536 VDD.n3375 VDD.n2830 2.2505
R26537 VDD.n3374 VDD.n3373 2.2505
R26538 VDD.n3372 VDD.n2831 2.2505
R26539 VDD.n3371 VDD.n3370 2.2505
R26540 VDD.n3369 VDD.n2832 2.2505
R26541 VDD.n3368 VDD.n3367 2.2505
R26542 VDD.n3366 VDD.n2833 2.2505
R26543 VDD.n3365 VDD.n3364 2.2505
R26544 VDD.n3363 VDD.n2834 2.2505
R26545 VDD.n3362 VDD.n3361 2.2505
R26546 VDD.n3360 VDD.n2835 2.2505
R26547 VDD.n3359 VDD.n3358 2.2505
R26548 VDD.n3357 VDD.n2836 2.2505
R26549 VDD.n3356 VDD.n3355 2.2505
R26550 VDD.n3354 VDD.n2837 2.2505
R26551 VDD.n3353 VDD.n3352 2.2505
R26552 VDD.n3351 VDD.n2838 2.2505
R26553 VDD.n3350 VDD.n3349 2.2505
R26554 VDD.n3348 VDD.n2839 2.2505
R26555 VDD.n3347 VDD.n3346 2.2505
R26556 VDD.n3345 VDD.n2840 2.2505
R26557 VDD.n3344 VDD.n3343 2.2505
R26558 VDD.n3342 VDD.n2841 2.2505
R26559 VDD.n3341 VDD.n3340 2.2505
R26560 VDD.n3339 VDD.n2842 2.2505
R26561 VDD.n3338 VDD.n3337 2.2505
R26562 VDD.n3336 VDD.n2843 2.2505
R26563 VDD.n3335 VDD.n3334 2.2505
R26564 VDD.n3333 VDD.n2844 2.2505
R26565 VDD.n3332 VDD.n3331 2.2505
R26566 VDD.n3330 VDD.n2845 2.2505
R26567 VDD.n3329 VDD.n3328 2.2505
R26568 VDD.n3327 VDD.n2846 2.2505
R26569 VDD.n3326 VDD.n3325 2.2505
R26570 VDD.n3324 VDD.n2847 2.2505
R26571 VDD.n3323 VDD.n3322 2.2505
R26572 VDD.n3321 VDD.n2848 2.2505
R26573 VDD.n3320 VDD.n3319 2.2505
R26574 VDD.n3318 VDD.n2849 2.2505
R26575 VDD.n3317 VDD.n3316 2.2505
R26576 VDD.n3315 VDD.n2850 2.2505
R26577 VDD.n3314 VDD.n3313 2.2505
R26578 VDD.n3312 VDD.n2851 2.2505
R26579 VDD.n3311 VDD.n3310 2.2505
R26580 VDD.n3309 VDD.n2852 2.2505
R26581 VDD.n3308 VDD.n3307 2.2505
R26582 VDD.n3306 VDD.n2853 2.2505
R26583 VDD.n3305 VDD.n3304 2.2505
R26584 VDD.n3303 VDD.n2854 2.2505
R26585 VDD.n3302 VDD.n3301 2.2505
R26586 VDD.n3300 VDD.n2855 2.2505
R26587 VDD.n3299 VDD.n3298 2.2505
R26588 VDD.n3297 VDD.n2856 2.2505
R26589 VDD.n3296 VDD.n3295 2.2505
R26590 VDD.n3294 VDD.n2857 2.2505
R26591 VDD.n3293 VDD.n3292 2.2505
R26592 VDD.n3291 VDD.n2858 2.2505
R26593 VDD.n3290 VDD.n3289 2.2505
R26594 VDD.n3288 VDD.n2859 2.2505
R26595 VDD.n3287 VDD.n3286 2.2505
R26596 VDD.n3285 VDD.n2860 2.2505
R26597 VDD.n3284 VDD.n3283 2.2505
R26598 VDD.n3282 VDD.n2861 2.2505
R26599 VDD.n3281 VDD.n3280 2.2505
R26600 VDD.n3279 VDD.n2862 2.2505
R26601 VDD.n3278 VDD.n3277 2.2505
R26602 VDD.n3276 VDD.n2863 2.2505
R26603 VDD.n3275 VDD.n3274 2.2505
R26604 VDD.n3273 VDD.n2864 2.2505
R26605 VDD.n3272 VDD.n3271 2.2505
R26606 VDD.n3270 VDD.n2865 2.2505
R26607 VDD.n3269 VDD.n3268 2.2505
R26608 VDD.n3267 VDD.n2866 2.2505
R26609 VDD.n3266 VDD.n3265 2.2505
R26610 VDD.n3264 VDD.n2867 2.2505
R26611 VDD.n3263 VDD.n3262 2.2505
R26612 VDD.n3261 VDD.n2868 2.2505
R26613 VDD.n3260 VDD.n3259 2.2505
R26614 VDD.n3258 VDD.n2869 2.2505
R26615 VDD.n3257 VDD.n3256 2.2505
R26616 VDD.n3255 VDD.n2870 2.2505
R26617 VDD.n3254 VDD.n3253 2.2505
R26618 VDD.n3252 VDD.n2871 2.2505
R26619 VDD.n3251 VDD.n3250 2.2505
R26620 VDD.n3249 VDD.n2872 2.2505
R26621 VDD.n3248 VDD.n3247 2.2505
R26622 VDD.n3246 VDD.n2873 2.2505
R26623 VDD.n3245 VDD.n3244 2.2505
R26624 VDD.n3243 VDD.n2874 2.2505
R26625 VDD.n3242 VDD.n3241 2.2505
R26626 VDD.n3240 VDD.n2875 2.2505
R26627 VDD.n3239 VDD.n3238 2.2505
R26628 VDD.n3237 VDD.n2876 2.2505
R26629 VDD.n3236 VDD.n3235 2.2505
R26630 VDD.n3234 VDD.n2877 2.2505
R26631 VDD.n3233 VDD.n3232 2.2505
R26632 VDD.n3231 VDD.n2878 2.2505
R26633 VDD.n3230 VDD.n3229 2.2505
R26634 VDD.n3228 VDD.n2879 2.2505
R26635 VDD.n3227 VDD.n3226 2.2505
R26636 VDD.n3225 VDD.n2880 2.2505
R26637 VDD.n3224 VDD.n3223 2.2505
R26638 VDD.n3222 VDD.n2881 2.2505
R26639 VDD.n3221 VDD.n3220 2.2505
R26640 VDD.n3219 VDD.n2882 2.2505
R26641 VDD.n3218 VDD.n3217 2.2505
R26642 VDD.n3216 VDD.n2883 2.2505
R26643 VDD.n3215 VDD.n3214 2.2505
R26644 VDD.n3213 VDD.n2884 2.2505
R26645 VDD.n3212 VDD.n3211 2.2505
R26646 VDD.n3210 VDD.n2885 2.2505
R26647 VDD.n3209 VDD.n3208 2.2505
R26648 VDD.n3207 VDD.n2886 2.2505
R26649 VDD.n3206 VDD.n3205 2.2505
R26650 VDD.n3204 VDD.n2887 2.2505
R26651 VDD.n3203 VDD.n3202 2.2505
R26652 VDD.n3201 VDD.n2888 2.2505
R26653 VDD.n3200 VDD.n3199 2.2505
R26654 VDD.n3198 VDD.n2889 2.2505
R26655 VDD.n3197 VDD.n3196 2.2505
R26656 VDD.n3195 VDD.n2890 2.2505
R26657 VDD.n3194 VDD.n3193 2.2505
R26658 VDD.n3192 VDD.n2891 2.2505
R26659 VDD.n3191 VDD.n3190 2.2505
R26660 VDD.n3189 VDD.n2892 2.2505
R26661 VDD.n3188 VDD.n3187 2.2505
R26662 VDD.n3186 VDD.n2893 2.2505
R26663 VDD.n3185 VDD.n3184 2.2505
R26664 VDD.n3183 VDD.n2894 2.2505
R26665 VDD.n3182 VDD.n3181 2.2505
R26666 VDD.n3180 VDD.n2895 2.2505
R26667 VDD.n3179 VDD.n3178 2.2505
R26668 VDD.n3177 VDD.n2896 2.2505
R26669 VDD.n3176 VDD.n3175 2.2505
R26670 VDD.n3174 VDD.n2897 2.2505
R26671 VDD.n3173 VDD.n3172 2.2505
R26672 VDD.n3171 VDD.n2898 2.2505
R26673 VDD.n3170 VDD.n3169 2.2505
R26674 VDD.n3168 VDD.n2899 2.2505
R26675 VDD.n3167 VDD.n3166 2.2505
R26676 VDD.n3165 VDD.n2900 2.2505
R26677 VDD.n3164 VDD.n3163 2.2505
R26678 VDD.n3162 VDD.n2901 2.2505
R26679 VDD.n3161 VDD.n3160 2.2505
R26680 VDD.n3159 VDD.n2902 2.2505
R26681 VDD.n3158 VDD.n3157 2.2505
R26682 VDD.n3156 VDD.n2903 2.2505
R26683 VDD.n3155 VDD.n3154 2.2505
R26684 VDD.n3153 VDD.n2904 2.2505
R26685 VDD.n3152 VDD.n3151 2.2505
R26686 VDD.n3150 VDD.n2905 2.2505
R26687 VDD.n3149 VDD.n3148 2.2505
R26688 VDD.n3147 VDD.n2906 2.2505
R26689 VDD.n3146 VDD.n3145 2.2505
R26690 VDD.n3144 VDD.n2907 2.2505
R26691 VDD.n3143 VDD.n3142 2.2505
R26692 VDD.n3141 VDD.n2908 2.2505
R26693 VDD.n3140 VDD.n3139 2.2505
R26694 VDD.n3138 VDD.n2909 2.2505
R26695 VDD.n3137 VDD.n3136 2.2505
R26696 VDD.n3135 VDD.n2910 2.2505
R26697 VDD.n3134 VDD.n3133 2.2505
R26698 VDD.n3132 VDD.n2911 2.2505
R26699 VDD.n3131 VDD.n3130 2.2505
R26700 VDD.n3129 VDD.n2912 2.2505
R26701 VDD.n3128 VDD.n3127 2.2505
R26702 VDD.n3126 VDD.n2913 2.2505
R26703 VDD.n3125 VDD.n3124 2.2505
R26704 VDD.n3123 VDD.n2914 2.2505
R26705 VDD.n3122 VDD.n3121 2.2505
R26706 VDD.n3120 VDD.n2915 2.2505
R26707 VDD.n3119 VDD.n3118 2.2505
R26708 VDD.n3117 VDD.n2916 2.2505
R26709 VDD.n3116 VDD.n3115 2.2505
R26710 VDD.n3114 VDD.n2917 2.2505
R26711 VDD.n3113 VDD.n3112 2.2505
R26712 VDD.n3111 VDD.n2918 2.2505
R26713 VDD.n3110 VDD.n3109 2.2505
R26714 VDD.n3108 VDD.n2919 2.2505
R26715 VDD.n3107 VDD.n3106 2.2505
R26716 VDD.n3105 VDD.n2920 2.2505
R26717 VDD.n3104 VDD.n3103 2.2505
R26718 VDD.n3102 VDD.n2921 2.2505
R26719 VDD.n3101 VDD.n3100 2.2505
R26720 VDD.n3099 VDD.n2922 2.2505
R26721 VDD.n3098 VDD.n3097 2.2505
R26722 VDD.n3096 VDD.n2923 2.2505
R26723 VDD.n3095 VDD.n3094 2.2505
R26724 VDD.n3093 VDD.n2924 2.2505
R26725 VDD.n3092 VDD.n3091 2.2505
R26726 VDD.n3090 VDD.n2925 2.2505
R26727 VDD.n3089 VDD.n3088 2.2505
R26728 VDD.n3087 VDD.n2926 2.2505
R26729 VDD.n3086 VDD.n3085 2.2505
R26730 VDD.n3084 VDD.n2927 2.2505
R26731 VDD.n3083 VDD.n3082 2.2505
R26732 VDD.n3081 VDD.n2928 2.2505
R26733 VDD.n3080 VDD.n3079 2.2505
R26734 VDD.n3078 VDD.n2929 2.2505
R26735 VDD.n3077 VDD.n3076 2.2505
R26736 VDD.n3075 VDD.n2930 2.2505
R26737 VDD.n3074 VDD.n3073 2.2505
R26738 VDD.n3072 VDD.n2931 2.2505
R26739 VDD.n3071 VDD.n3070 2.2505
R26740 VDD.n3069 VDD.n2932 2.2505
R26741 VDD.n3068 VDD.n3067 2.2505
R26742 VDD.n3066 VDD.n2933 2.2505
R26743 VDD.n3065 VDD.n3064 2.2505
R26744 VDD.n3063 VDD.n2934 2.2505
R26745 VDD.n3062 VDD.n3061 2.2505
R26746 VDD.n3060 VDD.n2935 2.2505
R26747 VDD.n3059 VDD.n3058 2.2505
R26748 VDD.n3057 VDD.n2936 2.2505
R26749 VDD.n3056 VDD.n3055 2.2505
R26750 VDD.n3054 VDD.n2937 2.2505
R26751 VDD.n3053 VDD.n3052 2.2505
R26752 VDD.n3051 VDD.n2938 2.2505
R26753 VDD.n3050 VDD.n3049 2.2505
R26754 VDD.n3048 VDD.n2939 2.2505
R26755 VDD.n3047 VDD.n3046 2.2505
R26756 VDD.n3045 VDD.n2940 2.2505
R26757 VDD.n3044 VDD.n3043 2.2505
R26758 VDD.n3042 VDD.n2941 2.2505
R26759 VDD.n3041 VDD.n3040 2.2505
R26760 VDD.n3039 VDD.n2942 2.2505
R26761 VDD.n3038 VDD.n3037 2.2505
R26762 VDD.n3036 VDD.n2943 2.2505
R26763 VDD.n3035 VDD.n3034 2.2505
R26764 VDD.n3033 VDD.n2944 2.2505
R26765 VDD.n3032 VDD.n3031 2.2505
R26766 VDD.n3030 VDD.n2945 2.2505
R26767 VDD.n3029 VDD.n3028 2.2505
R26768 VDD.n3027 VDD.n2946 2.2505
R26769 VDD.n3026 VDD.n3025 2.2505
R26770 VDD.n3024 VDD.n2947 2.2505
R26771 VDD.n3023 VDD.n3022 2.2505
R26772 VDD.n3021 VDD.n2948 2.2505
R26773 VDD.n3020 VDD.n3019 2.2505
R26774 VDD.n3018 VDD.n2949 2.2505
R26775 VDD.n3017 VDD.n3016 2.2505
R26776 VDD.n3015 VDD.n2950 2.2505
R26777 VDD.n3014 VDD.n3013 2.2505
R26778 VDD.n3012 VDD.n2951 2.2505
R26779 VDD.n3011 VDD.n3010 2.2505
R26780 VDD.n3009 VDD.n2952 2.2505
R26781 VDD.n3008 VDD.n3007 2.2505
R26782 VDD.n3006 VDD.n2953 2.2505
R26783 VDD.n3005 VDD.n3004 2.2505
R26784 VDD.n3003 VDD.n2954 2.2505
R26785 VDD.n3002 VDD.n3001 2.2505
R26786 VDD.n3000 VDD.n2955 2.2505
R26787 VDD.n2999 VDD.n2998 2.2505
R26788 VDD.n2997 VDD.n2956 2.2505
R26789 VDD.n2996 VDD.n2995 2.2505
R26790 VDD.n2994 VDD.n2957 2.2505
R26791 VDD.n2993 VDD.n2992 2.2505
R26792 VDD.n2991 VDD.n2958 2.2505
R26793 VDD.n2990 VDD.n2989 2.2505
R26794 VDD.n2988 VDD.n2959 2.2505
R26795 VDD.n2987 VDD.n2986 2.2505
R26796 VDD.n2985 VDD.n2960 2.2505
R26797 VDD.n2984 VDD.n2983 2.2505
R26798 VDD.n2982 VDD.n2961 2.2505
R26799 VDD.n2981 VDD.n2980 2.2505
R26800 VDD.n2979 VDD.n2962 2.2505
R26801 VDD.n2978 VDD.n2977 2.2505
R26802 VDD.n2976 VDD.n2963 2.2505
R26803 VDD.n2975 VDD.n2974 2.2505
R26804 VDD.n2973 VDD.n2964 2.2505
R26805 VDD.n2972 VDD.n2971 2.2505
R26806 VDD.n2970 VDD.n2965 2.2505
R26807 VDD.n2969 VDD.n2968 2.2505
R26808 VDD.n11135 VDD.n11134 2.2505
R26809 VDD.n11136 VDD.n630 2.2505
R26810 VDD.n11138 VDD.n11137 2.2505
R26811 VDD.n11139 VDD.n629 2.2505
R26812 VDD.n11141 VDD.n11140 2.2505
R26813 VDD.n11142 VDD.n628 2.2505
R26814 VDD.n11144 VDD.n11143 2.2505
R26815 VDD.n11145 VDD.n627 2.2505
R26816 VDD.n11147 VDD.n11146 2.2505
R26817 VDD.n11148 VDD.n626 2.2505
R26818 VDD.n11150 VDD.n11149 2.2505
R26819 VDD.n11151 VDD.n625 2.2505
R26820 VDD.n11153 VDD.n11152 2.2505
R26821 VDD.n11154 VDD.n624 2.2505
R26822 VDD.n11156 VDD.n11155 2.2505
R26823 VDD.n11157 VDD.n623 2.2505
R26824 VDD.n11159 VDD.n11158 2.2505
R26825 VDD.n11160 VDD.n622 2.2505
R26826 VDD.n11162 VDD.n11161 2.2505
R26827 VDD.n11163 VDD.n621 2.2505
R26828 VDD.n11165 VDD.n11164 2.2505
R26829 VDD.n11166 VDD.n620 2.2505
R26830 VDD.n11168 VDD.n11167 2.2505
R26831 VDD.n11169 VDD.n619 2.2505
R26832 VDD.n11171 VDD.n11170 2.2505
R26833 VDD.n11172 VDD.n618 2.2505
R26834 VDD.n11174 VDD.n11173 2.2505
R26835 VDD.n11175 VDD.n617 2.2505
R26836 VDD.n11177 VDD.n11176 2.2505
R26837 VDD.n11178 VDD.n616 2.2505
R26838 VDD.n11180 VDD.n11179 2.2505
R26839 VDD.n11181 VDD.n615 2.2505
R26840 VDD.n11183 VDD.n11182 2.2505
R26841 VDD.n11184 VDD.n614 2.2505
R26842 VDD.n11186 VDD.n11185 2.2505
R26843 VDD.n11187 VDD.n613 2.2505
R26844 VDD.n11189 VDD.n11188 2.2505
R26845 VDD.n11190 VDD.n612 2.2505
R26846 VDD.n11192 VDD.n11191 2.2505
R26847 VDD.n11193 VDD.n611 2.2505
R26848 VDD.n11195 VDD.n11194 2.2505
R26849 VDD.n11196 VDD.n610 2.2505
R26850 VDD.n11198 VDD.n11197 2.2505
R26851 VDD.n11199 VDD.n609 2.2505
R26852 VDD.n11201 VDD.n11200 2.2505
R26853 VDD.n11202 VDD.n608 2.2505
R26854 VDD.n11204 VDD.n11203 2.2505
R26855 VDD.n11205 VDD.n607 2.2505
R26856 VDD.n11207 VDD.n11206 2.2505
R26857 VDD.n11208 VDD.n606 2.2505
R26858 VDD.n11210 VDD.n11209 2.2505
R26859 VDD.n11211 VDD.n605 2.2505
R26860 VDD.n11213 VDD.n11212 2.2505
R26861 VDD.n11214 VDD.n604 2.2505
R26862 VDD.n11216 VDD.n11215 2.2505
R26863 VDD.n11217 VDD.n603 2.2505
R26864 VDD.n11219 VDD.n11218 2.2505
R26865 VDD.n11220 VDD.n602 2.2505
R26866 VDD.n11222 VDD.n11221 2.2505
R26867 VDD.n11223 VDD.n601 2.2505
R26868 VDD.n11225 VDD.n11224 2.2505
R26869 VDD.n11226 VDD.n600 2.2505
R26870 VDD.n11228 VDD.n11227 2.2505
R26871 VDD.n11229 VDD.n599 2.2505
R26872 VDD.n11231 VDD.n11230 2.2505
R26873 VDD.n11232 VDD.n598 2.2505
R26874 VDD.n11234 VDD.n11233 2.2505
R26875 VDD.n11235 VDD.n597 2.2505
R26876 VDD.n11237 VDD.n11236 2.2505
R26877 VDD.n11238 VDD.n596 2.2505
R26878 VDD.n11240 VDD.n11239 2.2505
R26879 VDD.n11241 VDD.n595 2.2505
R26880 VDD.n11243 VDD.n11242 2.2505
R26881 VDD.n11244 VDD.n594 2.2505
R26882 VDD.n11246 VDD.n11245 2.2505
R26883 VDD.n11247 VDD.n593 2.2505
R26884 VDD.n11249 VDD.n11248 2.2505
R26885 VDD.n11250 VDD.n592 2.2505
R26886 VDD.n11252 VDD.n11251 2.2505
R26887 VDD.n11253 VDD.n591 2.2505
R26888 VDD.n11255 VDD.n11254 2.2505
R26889 VDD.n11256 VDD.n590 2.2505
R26890 VDD.n11258 VDD.n11257 2.2505
R26891 VDD.n11259 VDD.n589 2.2505
R26892 VDD.n11261 VDD.n11260 2.2505
R26893 VDD.n11262 VDD.n588 2.2505
R26894 VDD.n11264 VDD.n11263 2.2505
R26895 VDD.n11265 VDD.n587 2.2505
R26896 VDD.n11267 VDD.n11266 2.2505
R26897 VDD.n11268 VDD.n586 2.2505
R26898 VDD.n11270 VDD.n11269 2.2505
R26899 VDD.n11271 VDD.n585 2.2505
R26900 VDD.n11273 VDD.n11272 2.2505
R26901 VDD.n11274 VDD.n584 2.2505
R26902 VDD.n11276 VDD.n11275 2.2505
R26903 VDD.n11277 VDD.n583 2.2505
R26904 VDD.n11279 VDD.n11278 2.2505
R26905 VDD.n11280 VDD.n582 2.2505
R26906 VDD.n11282 VDD.n11281 2.2505
R26907 VDD.n11283 VDD.n581 2.2505
R26908 VDD.n11285 VDD.n11284 2.2505
R26909 VDD.n11286 VDD.n580 2.2505
R26910 VDD.n11288 VDD.n11287 2.2505
R26911 VDD.n11289 VDD.n579 2.2505
R26912 VDD.n11291 VDD.n11290 2.2505
R26913 VDD.n11292 VDD.n578 2.2505
R26914 VDD.n11294 VDD.n11293 2.2505
R26915 VDD.n11295 VDD.n577 2.2505
R26916 VDD.n11297 VDD.n11296 2.2505
R26917 VDD.n11298 VDD.n576 2.2505
R26918 VDD.n11300 VDD.n11299 2.2505
R26919 VDD.n11301 VDD.n575 2.2505
R26920 VDD.n11303 VDD.n11302 2.2505
R26921 VDD.n11304 VDD.n574 2.2505
R26922 VDD.n11306 VDD.n11305 2.2505
R26923 VDD.n11307 VDD.n573 2.2505
R26924 VDD.n11309 VDD.n11308 2.2505
R26925 VDD.n11310 VDD.n572 2.2505
R26926 VDD.n11312 VDD.n11311 2.2505
R26927 VDD.n11313 VDD.n571 2.2505
R26928 VDD.n11315 VDD.n11314 2.2505
R26929 VDD.n11316 VDD.n570 2.2505
R26930 VDD.n11318 VDD.n11317 2.2505
R26931 VDD.n11319 VDD.n569 2.2505
R26932 VDD.n11321 VDD.n11320 2.2505
R26933 VDD.n11322 VDD.n568 2.2505
R26934 VDD.n11324 VDD.n11323 2.2505
R26935 VDD.n11325 VDD.n567 2.2505
R26936 VDD.n11327 VDD.n11326 2.2505
R26937 VDD.n11328 VDD.n566 2.2505
R26938 VDD.n11330 VDD.n11329 2.2505
R26939 VDD.n11331 VDD.n565 2.2505
R26940 VDD.n11333 VDD.n11332 2.2505
R26941 VDD.n11334 VDD.n564 2.2505
R26942 VDD.n11336 VDD.n11335 2.2505
R26943 VDD.n11337 VDD.n563 2.2505
R26944 VDD.n11339 VDD.n11338 2.2505
R26945 VDD.n11340 VDD.n562 2.2505
R26946 VDD.n11342 VDD.n11341 2.2505
R26947 VDD.n11343 VDD.n561 2.2505
R26948 VDD.n11345 VDD.n11344 2.2505
R26949 VDD.n11346 VDD.n560 2.2505
R26950 VDD.n11348 VDD.n11347 2.2505
R26951 VDD.n11349 VDD.n559 2.2505
R26952 VDD.n11351 VDD.n11350 2.2505
R26953 VDD.n11352 VDD.n558 2.2505
R26954 VDD.n11354 VDD.n11353 2.2505
R26955 VDD.n11355 VDD.n557 2.2505
R26956 VDD.n11357 VDD.n11356 2.2505
R26957 VDD.n11358 VDD.n556 2.2505
R26958 VDD.n11360 VDD.n11359 2.2505
R26959 VDD.n11361 VDD.n555 2.2505
R26960 VDD.n11363 VDD.n11362 2.2505
R26961 VDD.n11364 VDD.n554 2.2505
R26962 VDD.n11366 VDD.n11365 2.2505
R26963 VDD.n11367 VDD.n553 2.2505
R26964 VDD.n11369 VDD.n11368 2.2505
R26965 VDD.n11370 VDD.n552 2.2505
R26966 VDD.n11372 VDD.n11371 2.2505
R26967 VDD.n11373 VDD.n551 2.2505
R26968 VDD.n11375 VDD.n11374 2.2505
R26969 VDD.n11376 VDD.n550 2.2505
R26970 VDD.n11378 VDD.n11377 2.2505
R26971 VDD.n11379 VDD.n549 2.2505
R26972 VDD.n11381 VDD.n11380 2.2505
R26973 VDD.n11382 VDD.n548 2.2505
R26974 VDD.n11384 VDD.n11383 2.2505
R26975 VDD.n11385 VDD.n547 2.2505
R26976 VDD.n11387 VDD.n11386 2.2505
R26977 VDD.n11388 VDD.n546 2.2505
R26978 VDD.n11390 VDD.n11389 2.2505
R26979 VDD.n11391 VDD.n545 2.2505
R26980 VDD.n11393 VDD.n11392 2.2505
R26981 VDD.n11394 VDD.n544 2.2505
R26982 VDD.n11396 VDD.n11395 2.2505
R26983 VDD.n11397 VDD.n543 2.2505
R26984 VDD.n11399 VDD.n11398 2.2505
R26985 VDD.n11400 VDD.n542 2.2505
R26986 VDD.n11402 VDD.n11401 2.2505
R26987 VDD.n11403 VDD.n541 2.2505
R26988 VDD.n11405 VDD.n11404 2.2505
R26989 VDD.n11406 VDD.n540 2.2505
R26990 VDD.n11408 VDD.n11407 2.2505
R26991 VDD.n11409 VDD.n539 2.2505
R26992 VDD.n11411 VDD.n11410 2.2505
R26993 VDD.n11412 VDD.n538 2.2505
R26994 VDD.n11414 VDD.n11413 2.2505
R26995 VDD.n11415 VDD.n537 2.2505
R26996 VDD.n11417 VDD.n11416 2.2505
R26997 VDD.n11418 VDD.n536 2.2505
R26998 VDD.n11420 VDD.n11419 2.2505
R26999 VDD.n11421 VDD.n535 2.2505
R27000 VDD.n11423 VDD.n11422 2.2505
R27001 VDD.n11424 VDD.n534 2.2505
R27002 VDD.n11426 VDD.n11425 2.2505
R27003 VDD.n11427 VDD.n533 2.2505
R27004 VDD.n11429 VDD.n11428 2.2505
R27005 VDD.n11430 VDD.n532 2.2505
R27006 VDD.n11432 VDD.n11431 2.2505
R27007 VDD.n11433 VDD.n531 2.2505
R27008 VDD.n11435 VDD.n11434 2.2505
R27009 VDD.n11436 VDD.n530 2.2505
R27010 VDD.n11438 VDD.n11437 2.2505
R27011 VDD.n11439 VDD.n529 2.2505
R27012 VDD.n11441 VDD.n11440 2.2505
R27013 VDD.n11442 VDD.n528 2.2505
R27014 VDD.n11444 VDD.n11443 2.2505
R27015 VDD.n11445 VDD.n527 2.2505
R27016 VDD.n11447 VDD.n11446 2.2505
R27017 VDD.n11448 VDD.n526 2.2505
R27018 VDD.n11450 VDD.n11449 2.2505
R27019 VDD.n11451 VDD.n525 2.2505
R27020 VDD.n11453 VDD.n11452 2.2505
R27021 VDD.n11454 VDD.n524 2.2505
R27022 VDD.n11456 VDD.n11455 2.2505
R27023 VDD.n11457 VDD.n523 2.2505
R27024 VDD.n11459 VDD.n11458 2.2505
R27025 VDD.n11460 VDD.n522 2.2505
R27026 VDD.n11462 VDD.n11461 2.2505
R27027 VDD.n11463 VDD.n521 2.2505
R27028 VDD.n11465 VDD.n11464 2.2505
R27029 VDD.n11466 VDD.n520 2.2505
R27030 VDD.n11468 VDD.n11467 2.2505
R27031 VDD.n11469 VDD.n519 2.2505
R27032 VDD.n11471 VDD.n11470 2.2505
R27033 VDD.n11472 VDD.n518 2.2505
R27034 VDD.n11474 VDD.n11473 2.2505
R27035 VDD.n11475 VDD.n517 2.2505
R27036 VDD.n11477 VDD.n11476 2.2505
R27037 VDD.n11478 VDD.n516 2.2505
R27038 VDD.n11480 VDD.n11479 2.2505
R27039 VDD.n11481 VDD.n515 2.2505
R27040 VDD.n11483 VDD.n11482 2.2505
R27041 VDD.n11484 VDD.n514 2.2505
R27042 VDD.n11486 VDD.n11485 2.2505
R27043 VDD.n11487 VDD.n513 2.2505
R27044 VDD.n11489 VDD.n11488 2.2505
R27045 VDD.n11490 VDD.n512 2.2505
R27046 VDD.n11492 VDD.n11491 2.2505
R27047 VDD.n11493 VDD.n511 2.2505
R27048 VDD.n11495 VDD.n11494 2.2505
R27049 VDD.n11496 VDD.n510 2.2505
R27050 VDD.n11498 VDD.n11497 2.2505
R27051 VDD.n11499 VDD.n509 2.2505
R27052 VDD.n11501 VDD.n11500 2.2505
R27053 VDD.n11502 VDD.n508 2.2505
R27054 VDD.n11504 VDD.n11503 2.2505
R27055 VDD.n11505 VDD.n507 2.2505
R27056 VDD.n11507 VDD.n11506 2.2505
R27057 VDD.n11508 VDD.n506 2.2505
R27058 VDD.n11510 VDD.n11509 2.2505
R27059 VDD.n11511 VDD.n505 2.2505
R27060 VDD.n11513 VDD.n11512 2.2505
R27061 VDD.n11514 VDD.n504 2.2505
R27062 VDD.n11516 VDD.n11515 2.2505
R27063 VDD.n11517 VDD.n503 2.2505
R27064 VDD.n11519 VDD.n11518 2.2505
R27065 VDD.n11520 VDD.n502 2.2505
R27066 VDD.n11522 VDD.n11521 2.2505
R27067 VDD.n11523 VDD.n501 2.2505
R27068 VDD.n11525 VDD.n11524 2.2505
R27069 VDD.n11526 VDD.n500 2.2505
R27070 VDD.n11528 VDD.n11527 2.2505
R27071 VDD.n11529 VDD.n499 2.2505
R27072 VDD.n11531 VDD.n11530 2.2505
R27073 VDD.n11532 VDD.n498 2.2505
R27074 VDD.n11534 VDD.n11533 2.2505
R27075 VDD.n11535 VDD.n497 2.2505
R27076 VDD.n11537 VDD.n11536 2.2505
R27077 VDD.n11538 VDD.n496 2.2505
R27078 VDD.n11540 VDD.n11539 2.2505
R27079 VDD.n11541 VDD.n495 2.2505
R27080 VDD.n11543 VDD.n11542 2.2505
R27081 VDD.n11544 VDD.n494 2.2505
R27082 VDD.n11546 VDD.n11545 2.2505
R27083 VDD.n11547 VDD.n493 2.2505
R27084 VDD.n11549 VDD.n11548 2.2505
R27085 VDD.n11550 VDD.n492 2.2505
R27086 VDD.n11552 VDD.n11551 2.2505
R27087 VDD.n11553 VDD.n491 2.2505
R27088 VDD.n11555 VDD.n11554 2.2505
R27089 VDD.n11556 VDD.n490 2.2505
R27090 VDD.n11558 VDD.n11557 2.2505
R27091 VDD.n11559 VDD.n489 2.2505
R27092 VDD.n11561 VDD.n11560 2.2505
R27093 VDD.n11562 VDD.n488 2.2505
R27094 VDD.n11564 VDD.n11563 2.2505
R27095 VDD.n11565 VDD.n487 2.2505
R27096 VDD.n11567 VDD.n11566 2.2505
R27097 VDD.n11568 VDD.n486 2.2505
R27098 VDD.n11570 VDD.n11569 2.2505
R27099 VDD.n11571 VDD.n485 2.2505
R27100 VDD.n11573 VDD.n11572 2.2505
R27101 VDD.n11574 VDD.n484 2.2505
R27102 VDD.n11576 VDD.n11575 2.2505
R27103 VDD.n11577 VDD.n483 2.2505
R27104 VDD.n11579 VDD.n11578 2.2505
R27105 VDD.n11580 VDD.n482 2.2505
R27106 VDD.n11582 VDD.n11581 2.2505
R27107 VDD.n11583 VDD.n481 2.2505
R27108 VDD.n11585 VDD.n11584 2.2505
R27109 VDD.n11586 VDD.n480 2.2505
R27110 VDD.n11588 VDD.n11587 2.2505
R27111 VDD.n11589 VDD.n479 2.2505
R27112 VDD.n11591 VDD.n11590 2.2505
R27113 VDD.n11592 VDD.n478 2.2505
R27114 VDD.n11594 VDD.n11593 2.2505
R27115 VDD.n11595 VDD.n477 2.2505
R27116 VDD.n11597 VDD.n11596 2.2505
R27117 VDD.n11598 VDD.n476 2.2505
R27118 VDD.n11600 VDD.n11599 2.2505
R27119 VDD.n11601 VDD.n475 2.2505
R27120 VDD.n11603 VDD.n11602 2.2505
R27121 VDD.n11604 VDD.n474 2.2505
R27122 VDD.n11606 VDD.n11605 2.2505
R27123 VDD.n11607 VDD.n473 2.2505
R27124 VDD.n11609 VDD.n11608 2.2505
R27125 VDD.n11610 VDD.n472 2.2505
R27126 VDD.n11612 VDD.n11611 2.2505
R27127 VDD.n11613 VDD.n471 2.2505
R27128 VDD.n11615 VDD.n11614 2.2505
R27129 VDD.n11616 VDD.n470 2.2505
R27130 VDD.n11618 VDD.n11617 2.2505
R27131 VDD.n11619 VDD.n469 2.2505
R27132 VDD.n11621 VDD.n11620 2.2505
R27133 VDD.n11622 VDD.n468 2.2505
R27134 VDD.n11624 VDD.n11623 2.2505
R27135 VDD.n11625 VDD.n467 2.2505
R27136 VDD.n11627 VDD.n11626 2.2505
R27137 VDD.n11628 VDD.n466 2.2505
R27138 VDD.n11630 VDD.n11629 2.2505
R27139 VDD.n11631 VDD.n465 2.2505
R27140 VDD.n11633 VDD.n11632 2.2505
R27141 VDD.n11634 VDD.n464 2.2505
R27142 VDD.n11636 VDD.n11635 2.2505
R27143 VDD.n11637 VDD.n463 2.2505
R27144 VDD.n11639 VDD.n11638 2.2505
R27145 VDD.n11640 VDD.n462 2.2505
R27146 VDD.n11642 VDD.n11641 2.2505
R27147 VDD.n11643 VDD.n461 2.2505
R27148 VDD.n11645 VDD.n11644 2.2505
R27149 VDD.n11646 VDD.n460 2.2505
R27150 VDD.n11648 VDD.n11647 2.2505
R27151 VDD.n11649 VDD.n459 2.2505
R27152 VDD.n11651 VDD.n11650 2.2505
R27153 VDD.n11652 VDD.n458 2.2505
R27154 VDD.n11654 VDD.n11653 2.2505
R27155 VDD.n11655 VDD.n457 2.2505
R27156 VDD.n11657 VDD.n11656 2.2505
R27157 VDD.n11658 VDD.n456 2.2505
R27158 VDD.n11660 VDD.n11659 2.2505
R27159 VDD.n11661 VDD.n455 2.2505
R27160 VDD.n11663 VDD.n11662 2.2505
R27161 VDD.n11664 VDD.n454 2.2505
R27162 VDD.n11666 VDD.n11665 2.2505
R27163 VDD.n11667 VDD.n453 2.2505
R27164 VDD.n11669 VDD.n11668 2.2505
R27165 VDD.n11670 VDD.n452 2.2505
R27166 VDD.n11672 VDD.n11671 2.2505
R27167 VDD.n11673 VDD.n451 2.2505
R27168 VDD.n11675 VDD.n11674 2.2505
R27169 VDD.n11676 VDD.n450 2.2505
R27170 VDD.n11678 VDD.n11677 2.2505
R27171 VDD.n11679 VDD.n449 2.2505
R27172 VDD.n11681 VDD.n11680 2.2505
R27173 VDD.n11682 VDD.n448 2.2505
R27174 VDD.n11684 VDD.n11683 2.2505
R27175 VDD.n11685 VDD.n447 2.2505
R27176 VDD.n11687 VDD.n11686 2.2505
R27177 VDD.n11688 VDD.n446 2.2505
R27178 VDD.n11690 VDD.n11689 2.2505
R27179 VDD.n11691 VDD.n445 2.2505
R27180 VDD.n11693 VDD.n11692 2.2505
R27181 VDD.n11694 VDD.n444 2.2505
R27182 VDD.n11696 VDD.n11695 2.2505
R27183 VDD.n11697 VDD.n443 2.2505
R27184 VDD.n11699 VDD.n11698 2.2505
R27185 VDD.n11700 VDD.n442 2.2505
R27186 VDD.n11702 VDD.n11701 2.2505
R27187 VDD.n11703 VDD.n441 2.2505
R27188 VDD.n11705 VDD.n11704 2.2505
R27189 VDD.n11706 VDD.n440 2.2505
R27190 VDD.n11708 VDD.n11707 2.2505
R27191 VDD.n11709 VDD.n439 2.2505
R27192 VDD.n11711 VDD.n11710 2.2505
R27193 VDD.n11712 VDD.n438 2.2505
R27194 VDD.n11714 VDD.n11713 2.2505
R27195 VDD.n11715 VDD.n437 2.2505
R27196 VDD.n11717 VDD.n11716 2.2505
R27197 VDD.n11718 VDD.n436 2.2505
R27198 VDD.n11720 VDD.n11719 2.2505
R27199 VDD.n11721 VDD.n435 2.2505
R27200 VDD.n11723 VDD.n11722 2.2505
R27201 VDD.n11724 VDD.n434 2.2505
R27202 VDD.n11726 VDD.n11725 2.2505
R27203 VDD.n11727 VDD.n433 2.2505
R27204 VDD.n11729 VDD.n11728 2.2505
R27205 VDD.n11730 VDD.n432 2.2505
R27206 VDD.n11732 VDD.n11731 2.2505
R27207 VDD.n11733 VDD.n431 2.2505
R27208 VDD.n11735 VDD.n11734 2.2505
R27209 VDD.n11736 VDD.n430 2.2505
R27210 VDD.n11738 VDD.n11737 2.2505
R27211 VDD.n11739 VDD.n429 2.2505
R27212 VDD.n11741 VDD.n11740 2.2505
R27213 VDD.n11742 VDD.n428 2.2505
R27214 VDD.n11744 VDD.n11743 2.2505
R27215 VDD.n11745 VDD.n427 2.2505
R27216 VDD.n11747 VDD.n11746 2.2505
R27217 VDD.n11748 VDD.n426 2.2505
R27218 VDD.n11750 VDD.n11749 2.2505
R27219 VDD.n11751 VDD.n425 2.2505
R27220 VDD.n11753 VDD.n11752 2.2505
R27221 VDD.n11754 VDD.n424 2.2505
R27222 VDD.n11756 VDD.n11755 2.2505
R27223 VDD.n11757 VDD.n423 2.2505
R27224 VDD.n11759 VDD.n11758 2.2505
R27225 VDD.n11760 VDD.n422 2.2505
R27226 VDD.n11762 VDD.n11761 2.2505
R27227 VDD.n11763 VDD.n421 2.2505
R27228 VDD.n11765 VDD.n11764 2.2505
R27229 VDD.n11766 VDD.n420 2.2505
R27230 VDD.n11768 VDD.n11767 2.2505
R27231 VDD.n11769 VDD.n419 2.2505
R27232 VDD.n11771 VDD.n11770 2.2505
R27233 VDD.n11772 VDD.n418 2.2505
R27234 VDD.n11774 VDD.n11773 2.2505
R27235 VDD.n11775 VDD.n417 2.2505
R27236 VDD.n11777 VDD.n11776 2.2505
R27237 VDD.n11778 VDD.n416 2.2505
R27238 VDD.n11780 VDD.n11779 2.2505
R27239 VDD.n11781 VDD.n415 2.2505
R27240 VDD.n11783 VDD.n11782 2.2505
R27241 VDD.n11784 VDD.n414 2.2505
R27242 VDD.n11786 VDD.n11785 2.2505
R27243 VDD.n11787 VDD.n413 2.2505
R27244 VDD.n11789 VDD.n11788 2.2505
R27245 VDD.n11790 VDD.n412 2.2505
R27246 VDD.n11792 VDD.n11791 2.2505
R27247 VDD.n11793 VDD.n411 2.2505
R27248 VDD.n11795 VDD.n11794 2.2505
R27249 VDD.n11796 VDD.n410 2.2505
R27250 VDD.n11798 VDD.n11797 2.2505
R27251 VDD.n11799 VDD.n409 2.2505
R27252 VDD.n11801 VDD.n11800 2.2505
R27253 VDD.n11802 VDD.n408 2.2505
R27254 VDD.n11804 VDD.n11803 2.2505
R27255 VDD.n11805 VDD.n407 2.2505
R27256 VDD.n11807 VDD.n11806 2.2505
R27257 VDD.n11808 VDD.n406 2.2505
R27258 VDD.n11810 VDD.n11809 2.2505
R27259 VDD.n11811 VDD.n405 2.2505
R27260 VDD.n2967 VDD.n2966 2.2505
R27261 VDD.n10762 VDD.n10761 2.2505
R27262 VDD.n10763 VDD.n2062 2.2505
R27263 VDD.n10765 VDD.n10764 2.2505
R27264 VDD.n8253 VDD.n2061 2.2505
R27265 VDD.n8252 VDD.n8251 2.2505
R27266 VDD.n8248 VDD.n2063 2.2505
R27267 VDD.n8247 VDD.n8246 2.2505
R27268 VDD.n8245 VDD.n8244 2.2505
R27269 VDD.n8243 VDD.n2065 2.2505
R27270 VDD.n8242 VDD.n8241 2.2505
R27271 VDD.n8240 VDD.n2066 2.2505
R27272 VDD.n8239 VDD.n8238 2.2505
R27273 VDD.n8235 VDD.n2067 2.2505
R27274 VDD.n8234 VDD.n8233 2.2505
R27275 VDD.n8232 VDD.n2068 2.2505
R27276 VDD.n8231 VDD.n8230 2.2505
R27277 VDD.n8228 VDD.n2069 2.2505
R27278 VDD.n8227 VDD.n8226 2.2505
R27279 VDD.n8225 VDD.n2070 2.2505
R27280 VDD.n8224 VDD.n8223 2.2505
R27281 VDD.n8221 VDD.n2071 2.2505
R27282 VDD.n8220 VDD.n8219 2.2505
R27283 VDD.n8218 VDD.n2072 2.2505
R27284 VDD.n8217 VDD.n8216 2.2505
R27285 VDD.n8213 VDD.n2073 2.2505
R27286 VDD.n8212 VDD.n8211 2.2505
R27287 VDD.n8210 VDD.n8209 2.2505
R27288 VDD.n8208 VDD.n2075 2.2505
R27289 VDD.n8207 VDD.n8206 2.2505
R27290 VDD.n8205 VDD.n2076 2.2505
R27291 VDD.n8204 VDD.n8203 2.2505
R27292 VDD.n8200 VDD.n2077 2.2505
R27293 VDD.n8199 VDD.n8198 2.2505
R27294 VDD.n8197 VDD.n8196 2.2505
R27295 VDD.n8195 VDD.n2079 2.2505
R27296 VDD.n8194 VDD.n8193 2.2505
R27297 VDD.n8192 VDD.n2080 2.2505
R27298 VDD.n8191 VDD.n8190 2.2505
R27299 VDD.n8189 VDD.n2081 2.2505
R27300 VDD.n8187 VDD.n8186 2.2505
R27301 VDD.n8185 VDD.n2082 2.2505
R27302 VDD.n8184 VDD.n8183 2.2505
R27303 VDD.n8180 VDD.n2083 2.2505
R27304 VDD.n8179 VDD.n8178 2.2505
R27305 VDD.n8177 VDD.n2084 2.2505
R27306 VDD.n8176 VDD.n8175 2.2505
R27307 VDD.n8174 VDD.n2085 2.2505
R27308 VDD.n8172 VDD.n8171 2.2505
R27309 VDD.n8170 VDD.n2086 2.2505
R27310 VDD.n8169 VDD.n8168 2.2505
R27311 VDD.n2088 VDD.n2087 2.2505
R27312 VDD.n7304 VDD.n7303 2.2505
R27313 VDD.n7306 VDD.n7305 2.2505
R27314 VDD.n7307 VDD.n7302 2.2505
R27315 VDD.n7309 VDD.n7308 2.2505
R27316 VDD.n7310 VDD.n7301 2.2505
R27317 VDD.n7312 VDD.n7311 2.2505
R27318 VDD.n7313 VDD.n7300 2.2505
R27319 VDD.n7315 VDD.n7314 2.2505
R27320 VDD.n7316 VDD.n7299 2.2505
R27321 VDD.n7318 VDD.n7317 2.2505
R27322 VDD.n7319 VDD.n7298 2.2505
R27323 VDD.n7321 VDD.n7320 2.2505
R27324 VDD.n7322 VDD.n7297 2.2505
R27325 VDD.n7324 VDD.n7323 2.2505
R27326 VDD.n7325 VDD.n7296 2.2505
R27327 VDD.n7327 VDD.n7326 2.2505
R27328 VDD.n7328 VDD.n7295 2.2505
R27329 VDD.n7330 VDD.n7329 2.2505
R27330 VDD.n7331 VDD.n7294 2.2505
R27331 VDD.n7333 VDD.n7332 2.2505
R27332 VDD.n7334 VDD.n7293 2.2505
R27333 VDD.n7336 VDD.n7335 2.2505
R27334 VDD.n7337 VDD.n7292 2.2505
R27335 VDD.n7339 VDD.n7338 2.2505
R27336 VDD.n7340 VDD.n7291 2.2505
R27337 VDD.n7342 VDD.n7341 2.2505
R27338 VDD.n7343 VDD.n7290 2.2505
R27339 VDD.n7345 VDD.n7344 2.2505
R27340 VDD.n7346 VDD.n7289 2.2505
R27341 VDD.n7348 VDD.n7347 2.2505
R27342 VDD.n7349 VDD.n7288 2.2505
R27343 VDD.n7351 VDD.n7350 2.2505
R27344 VDD.n7352 VDD.n7287 2.2505
R27345 VDD.n7354 VDD.n7353 2.2505
R27346 VDD.n7355 VDD.n7286 2.2505
R27347 VDD.n7357 VDD.n7356 2.2505
R27348 VDD.n7358 VDD.n7285 2.2505
R27349 VDD.n7360 VDD.n7359 2.2505
R27350 VDD.n7361 VDD.n7284 2.2505
R27351 VDD.n7363 VDD.n7362 2.2505
R27352 VDD.n7364 VDD.n7283 2.2505
R27353 VDD.n7366 VDD.n7365 2.2505
R27354 VDD.n7367 VDD.n7282 2.2505
R27355 VDD.n7369 VDD.n7368 2.2505
R27356 VDD.n7370 VDD.n7281 2.2505
R27357 VDD.n7372 VDD.n7371 2.2505
R27358 VDD.n7373 VDD.n7280 2.2505
R27359 VDD.n7375 VDD.n7374 2.2505
R27360 VDD.n7376 VDD.n7279 2.2505
R27361 VDD.n7378 VDD.n7377 2.2505
R27362 VDD.n7379 VDD.n7278 2.2505
R27363 VDD.n7381 VDD.n7380 2.2505
R27364 VDD.n7382 VDD.n7277 2.2505
R27365 VDD.n7384 VDD.n7383 2.2505
R27366 VDD.n7385 VDD.n7276 2.2505
R27367 VDD.n7387 VDD.n7386 2.2505
R27368 VDD.n7388 VDD.n7275 2.2505
R27369 VDD.n7390 VDD.n7389 2.2505
R27370 VDD.n7391 VDD.n7274 2.2505
R27371 VDD.n7393 VDD.n7392 2.2505
R27372 VDD.n7394 VDD.n7273 2.2505
R27373 VDD.n7396 VDD.n7395 2.2505
R27374 VDD.n7397 VDD.n7272 2.2505
R27375 VDD.n7399 VDD.n7398 2.2505
R27376 VDD.n7400 VDD.n7271 2.2505
R27377 VDD.n7402 VDD.n7401 2.2505
R27378 VDD.n7403 VDD.n7270 2.2505
R27379 VDD.n7405 VDD.n7404 2.2505
R27380 VDD.n7406 VDD.n7269 2.2505
R27381 VDD.n7408 VDD.n7407 2.2505
R27382 VDD.n7409 VDD.n7268 2.2505
R27383 VDD.n7411 VDD.n7410 2.2505
R27384 VDD.n7412 VDD.n7267 2.2505
R27385 VDD.n7414 VDD.n7413 2.2505
R27386 VDD.n7415 VDD.n7266 2.2505
R27387 VDD.n7417 VDD.n7416 2.2505
R27388 VDD.n7418 VDD.n7265 2.2505
R27389 VDD.n7420 VDD.n7419 2.2505
R27390 VDD.n7421 VDD.n7264 2.2505
R27391 VDD.n7423 VDD.n7422 2.2505
R27392 VDD.n7424 VDD.n7263 2.2505
R27393 VDD.n7426 VDD.n7425 2.2505
R27394 VDD.n7427 VDD.n7262 2.2505
R27395 VDD.n7429 VDD.n7428 2.2505
R27396 VDD.n7430 VDD.n7261 2.2505
R27397 VDD.n7432 VDD.n7431 2.2505
R27398 VDD.n7433 VDD.n7260 2.2505
R27399 VDD.n7435 VDD.n7434 2.2505
R27400 VDD.n7436 VDD.n7259 2.2505
R27401 VDD.n7438 VDD.n7437 2.2505
R27402 VDD.n7439 VDD.n7258 2.2505
R27403 VDD.n7441 VDD.n7440 2.2505
R27404 VDD.n7442 VDD.n7257 2.2505
R27405 VDD.n7444 VDD.n7443 2.2505
R27406 VDD.n7445 VDD.n7256 2.2505
R27407 VDD.n7447 VDD.n7446 2.2505
R27408 VDD.n7448 VDD.n7255 2.2505
R27409 VDD.n7450 VDD.n7449 2.2505
R27410 VDD.n7451 VDD.n7254 2.2505
R27411 VDD.n7453 VDD.n7452 2.2505
R27412 VDD.n7454 VDD.n7253 2.2505
R27413 VDD.n7456 VDD.n7455 2.2505
R27414 VDD.n7457 VDD.n7252 2.2505
R27415 VDD.n7459 VDD.n7458 2.2505
R27416 VDD.n7460 VDD.n7251 2.2505
R27417 VDD.n7462 VDD.n7461 2.2505
R27418 VDD.n7463 VDD.n7250 2.2505
R27419 VDD.n7465 VDD.n7464 2.2505
R27420 VDD.n7466 VDD.n7249 2.2505
R27421 VDD.n7468 VDD.n7467 2.2505
R27422 VDD.n7469 VDD.n7248 2.2505
R27423 VDD.n7471 VDD.n7470 2.2505
R27424 VDD.n7472 VDD.n7247 2.2505
R27425 VDD.n7474 VDD.n7473 2.2505
R27426 VDD.n7475 VDD.n7246 2.2505
R27427 VDD.n7477 VDD.n7476 2.2505
R27428 VDD.n7478 VDD.n7245 2.2505
R27429 VDD.n7480 VDD.n7479 2.2505
R27430 VDD.n7481 VDD.n7244 2.2505
R27431 VDD.n7483 VDD.n7482 2.2505
R27432 VDD.n7484 VDD.n7243 2.2505
R27433 VDD.n7486 VDD.n7485 2.2505
R27434 VDD.n7487 VDD.n7242 2.2505
R27435 VDD.n7489 VDD.n7488 2.2505
R27436 VDD.n7490 VDD.n7241 2.2505
R27437 VDD.n7492 VDD.n7491 2.2505
R27438 VDD.n7493 VDD.n7240 2.2505
R27439 VDD.n7495 VDD.n7494 2.2505
R27440 VDD.n7496 VDD.n7239 2.2505
R27441 VDD.n7498 VDD.n7497 2.2505
R27442 VDD.n7499 VDD.n7238 2.2505
R27443 VDD.n7501 VDD.n7500 2.2505
R27444 VDD.n7502 VDD.n7237 2.2505
R27445 VDD.n7504 VDD.n7503 2.2505
R27446 VDD.n7505 VDD.n7236 2.2505
R27447 VDD.n7507 VDD.n7506 2.2505
R27448 VDD.n7508 VDD.n7235 2.2505
R27449 VDD.n7510 VDD.n7509 2.2505
R27450 VDD.n7511 VDD.n7234 2.2505
R27451 VDD.n7513 VDD.n7512 2.2505
R27452 VDD.n7514 VDD.n7233 2.2505
R27453 VDD.n7516 VDD.n7515 2.2505
R27454 VDD.n7517 VDD.n7232 2.2505
R27455 VDD.n7519 VDD.n7518 2.2505
R27456 VDD.n7520 VDD.n7231 2.2505
R27457 VDD.n7522 VDD.n7521 2.2505
R27458 VDD.n7523 VDD.n7230 2.2505
R27459 VDD.n7525 VDD.n7524 2.2505
R27460 VDD.n7526 VDD.n7229 2.2505
R27461 VDD.n7528 VDD.n7527 2.2505
R27462 VDD.n7529 VDD.n7228 2.2505
R27463 VDD.n7531 VDD.n7530 2.2505
R27464 VDD.n7532 VDD.n7227 2.2505
R27465 VDD.n7534 VDD.n7533 2.2505
R27466 VDD.n7535 VDD.n7226 2.2505
R27467 VDD.n7537 VDD.n7536 2.2505
R27468 VDD.n7538 VDD.n7225 2.2505
R27469 VDD.n7540 VDD.n7539 2.2505
R27470 VDD.n7541 VDD.n7224 2.2505
R27471 VDD.n7543 VDD.n7542 2.2505
R27472 VDD.n7544 VDD.n7223 2.2505
R27473 VDD.n7546 VDD.n7545 2.2505
R27474 VDD.n7547 VDD.n7222 2.2505
R27475 VDD.n7549 VDD.n7548 2.2505
R27476 VDD.n7550 VDD.n7221 2.2505
R27477 VDD.n7552 VDD.n7551 2.2505
R27478 VDD.n7553 VDD.n7220 2.2505
R27479 VDD.n7555 VDD.n7554 2.2505
R27480 VDD.n7556 VDD.n7219 2.2505
R27481 VDD.n7558 VDD.n7557 2.2505
R27482 VDD.n7559 VDD.n7218 2.2505
R27483 VDD.n7561 VDD.n7560 2.2505
R27484 VDD.n7562 VDD.n7217 2.2505
R27485 VDD.n7564 VDD.n7563 2.2505
R27486 VDD.n7565 VDD.n7216 2.2505
R27487 VDD.n7567 VDD.n7566 2.2505
R27488 VDD.n7568 VDD.n7215 2.2505
R27489 VDD.n7570 VDD.n7569 2.2505
R27490 VDD.n7571 VDD.n7214 2.2505
R27491 VDD.n7573 VDD.n7572 2.2505
R27492 VDD.n7574 VDD.n7213 2.2505
R27493 VDD.n7576 VDD.n7575 2.2505
R27494 VDD.n7577 VDD.n7212 2.2505
R27495 VDD.n7579 VDD.n7578 2.2505
R27496 VDD.n7580 VDD.n7211 2.2505
R27497 VDD.n7582 VDD.n7581 2.2505
R27498 VDD.n7583 VDD.n7210 2.2505
R27499 VDD.n7585 VDD.n7584 2.2505
R27500 VDD.n7586 VDD.n7209 2.2505
R27501 VDD.n7588 VDD.n7587 2.2505
R27502 VDD.n7589 VDD.n7208 2.2505
R27503 VDD.n7591 VDD.n7590 2.2505
R27504 VDD.n7592 VDD.n7207 2.2505
R27505 VDD.n7594 VDD.n7593 2.2505
R27506 VDD.n7595 VDD.n7206 2.2505
R27507 VDD.n7597 VDD.n7596 2.2505
R27508 VDD.n7598 VDD.n7205 2.2505
R27509 VDD.n7600 VDD.n7599 2.2505
R27510 VDD.n7601 VDD.n7204 2.2505
R27511 VDD.n7603 VDD.n7602 2.2505
R27512 VDD.n7604 VDD.n7203 2.2505
R27513 VDD.n7606 VDD.n7605 2.2505
R27514 VDD.n7607 VDD.n7202 2.2505
R27515 VDD.n7609 VDD.n7608 2.2505
R27516 VDD.n7610 VDD.n7201 2.2505
R27517 VDD.n7612 VDD.n7611 2.2505
R27518 VDD.n7613 VDD.n7200 2.2505
R27519 VDD.n7615 VDD.n7614 2.2505
R27520 VDD.n7616 VDD.n7199 2.2505
R27521 VDD.n7618 VDD.n7617 2.2505
R27522 VDD.n7619 VDD.n7198 2.2505
R27523 VDD.n7621 VDD.n7620 2.2505
R27524 VDD.n7622 VDD.n7197 2.2505
R27525 VDD.n7624 VDD.n7623 2.2505
R27526 VDD.n7625 VDD.n7196 2.2505
R27527 VDD.n7627 VDD.n7626 2.2505
R27528 VDD.n7628 VDD.n7195 2.2505
R27529 VDD.n7630 VDD.n7629 2.2505
R27530 VDD.n7631 VDD.n7194 2.2505
R27531 VDD.n7633 VDD.n7632 2.2505
R27532 VDD.n7634 VDD.n7193 2.2505
R27533 VDD.n7636 VDD.n7635 2.2505
R27534 VDD.n7637 VDD.n7192 2.2505
R27535 VDD.n7639 VDD.n7638 2.2505
R27536 VDD.n7640 VDD.n7191 2.2505
R27537 VDD.n7642 VDD.n7641 2.2505
R27538 VDD.n7643 VDD.n7190 2.2505
R27539 VDD.n7645 VDD.n7644 2.2505
R27540 VDD.n7646 VDD.n7189 2.2505
R27541 VDD.n7648 VDD.n7647 2.2505
R27542 VDD.n7649 VDD.n7188 2.2505
R27543 VDD.n7651 VDD.n7650 2.2505
R27544 VDD.n7652 VDD.n7187 2.2505
R27545 VDD.n7654 VDD.n7653 2.2505
R27546 VDD.n7655 VDD.n7186 2.2505
R27547 VDD.n7657 VDD.n7656 2.2505
R27548 VDD.n7658 VDD.n7185 2.2505
R27549 VDD.n7660 VDD.n7659 2.2505
R27550 VDD.n7661 VDD.n7184 2.2505
R27551 VDD.n7663 VDD.n7662 2.2505
R27552 VDD.n7664 VDD.n7183 2.2505
R27553 VDD.n7666 VDD.n7665 2.2505
R27554 VDD.n7667 VDD.n7182 2.2505
R27555 VDD.n7669 VDD.n7668 2.2505
R27556 VDD.n7670 VDD.n7181 2.2505
R27557 VDD.n7672 VDD.n7671 2.2505
R27558 VDD.n7673 VDD.n7180 2.2505
R27559 VDD.n7675 VDD.n7674 2.2505
R27560 VDD.n7676 VDD.n7179 2.2505
R27561 VDD.n7678 VDD.n7677 2.2505
R27562 VDD.n7679 VDD.n7178 2.2505
R27563 VDD.n7681 VDD.n7680 2.2505
R27564 VDD.n7682 VDD.n2293 2.2505
R27565 VDD.n7685 VDD.n7684 2.2505
R27566 VDD.n7750 VDD.n7749 2.2505
R27567 VDD.n7751 VDD.n2268 2.2505
R27568 VDD.n7753 VDD.n7752 2.2505
R27569 VDD.n7754 VDD.n2267 2.2505
R27570 VDD.n7756 VDD.n7755 2.2505
R27571 VDD.n7757 VDD.n2266 2.2505
R27572 VDD.n7759 VDD.n7758 2.2505
R27573 VDD.n7761 VDD.n2264 2.2505
R27574 VDD.n7763 VDD.n7762 2.2505
R27575 VDD.n7764 VDD.n2263 2.2505
R27576 VDD.n7766 VDD.n7765 2.2505
R27577 VDD.n7767 VDD.n2262 2.2505
R27578 VDD.n7769 VDD.n7768 2.2505
R27579 VDD.n7770 VDD.n2261 2.2505
R27580 VDD.n7772 VDD.n7771 2.2505
R27581 VDD.n7773 VDD.n2259 2.2505
R27582 VDD.n7775 VDD.n7774 2.2505
R27583 VDD.n7776 VDD.n2258 2.2505
R27584 VDD.n7778 VDD.n7777 2.2505
R27585 VDD.n7779 VDD.n2257 2.2505
R27586 VDD.n7782 VDD.n7781 2.2505
R27587 VDD.n7783 VDD.n2256 2.2505
R27588 VDD.n7785 VDD.n7784 2.2505
R27589 VDD.n7786 VDD.n2255 2.2505
R27590 VDD.n7788 VDD.n7787 2.2505
R27591 VDD.n7789 VDD.n2254 2.2505
R27592 VDD.n7791 VDD.n7790 2.2505
R27593 VDD.n7792 VDD.n2253 2.2505
R27594 VDD.n7794 VDD.n7793 2.2505
R27595 VDD.n7796 VDD.n7795 2.2505
R27596 VDD.n7797 VDD.n2251 2.2505
R27597 VDD.n7799 VDD.n7798 2.2505
R27598 VDD.n7801 VDD.n7800 2.2505
R27599 VDD.n7802 VDD.n2249 2.2505
R27600 VDD.n7804 VDD.n7803 2.2505
R27601 VDD.n7805 VDD.n2248 2.2505
R27602 VDD.n7807 VDD.n7806 2.2505
R27603 VDD.n7808 VDD.n2247 2.2505
R27604 VDD.n7811 VDD.n7810 2.2505
R27605 VDD.n7812 VDD.n2246 2.2505
R27606 VDD.n7814 VDD.n7813 2.2505
R27607 VDD.n7815 VDD.n2245 2.2505
R27608 VDD.n7817 VDD.n7816 2.2505
R27609 VDD.n7818 VDD.n2243 2.2505
R27610 VDD.n7820 VDD.n7819 2.2505
R27611 VDD.n2244 VDD.n2242 2.2505
R27612 VDD.n4750 VDD.n4749 2.2505
R27613 VDD.n4751 VDD.n4748 2.2505
R27614 VDD.n4753 VDD.n4752 2.2505
R27615 VDD.n4754 VDD.n4747 2.2505
R27616 VDD.n4756 VDD.n4755 2.2505
R27617 VDD.n4757 VDD.n4746 2.2505
R27618 VDD.n4759 VDD.n4758 2.2505
R27619 VDD.n4760 VDD.n4745 2.2505
R27620 VDD.n4762 VDD.n4761 2.2505
R27621 VDD.n4763 VDD.n4744 2.2505
R27622 VDD.n4765 VDD.n4764 2.2505
R27623 VDD.n4766 VDD.n4743 2.2505
R27624 VDD.n4768 VDD.n4767 2.2505
R27625 VDD.n4769 VDD.n4742 2.2505
R27626 VDD.n4771 VDD.n4770 2.2505
R27627 VDD.n4772 VDD.n4741 2.2505
R27628 VDD.n4774 VDD.n4773 2.2505
R27629 VDD.n4775 VDD.n4740 2.2505
R27630 VDD.n4777 VDD.n4776 2.2505
R27631 VDD.n4778 VDD.n4739 2.2505
R27632 VDD.n4780 VDD.n4779 2.2505
R27633 VDD.n4781 VDD.n4738 2.2505
R27634 VDD.n4783 VDD.n4782 2.2505
R27635 VDD.n4784 VDD.n4737 2.2505
R27636 VDD.n4786 VDD.n4785 2.2505
R27637 VDD.n4787 VDD.n4736 2.2505
R27638 VDD.n4789 VDD.n4788 2.2505
R27639 VDD.n4790 VDD.n4735 2.2505
R27640 VDD.n4792 VDD.n4791 2.2505
R27641 VDD.n4793 VDD.n4734 2.2505
R27642 VDD.n4795 VDD.n4794 2.2505
R27643 VDD.n4796 VDD.n4733 2.2505
R27644 VDD.n4798 VDD.n4797 2.2505
R27645 VDD.n4799 VDD.n4732 2.2505
R27646 VDD.n4801 VDD.n4800 2.2505
R27647 VDD.n4802 VDD.n4731 2.2505
R27648 VDD.n4804 VDD.n4803 2.2505
R27649 VDD.n4805 VDD.n4730 2.2505
R27650 VDD.n4807 VDD.n4806 2.2505
R27651 VDD.n4808 VDD.n4729 2.2505
R27652 VDD.n4810 VDD.n4809 2.2505
R27653 VDD.n4811 VDD.n4728 2.2505
R27654 VDD.n4813 VDD.n4812 2.2505
R27655 VDD.n4814 VDD.n4727 2.2505
R27656 VDD.n4816 VDD.n4815 2.2505
R27657 VDD.n4817 VDD.n4726 2.2505
R27658 VDD.n4819 VDD.n4818 2.2505
R27659 VDD.n4820 VDD.n4725 2.2505
R27660 VDD.n4822 VDD.n4821 2.2505
R27661 VDD.n4823 VDD.n4724 2.2505
R27662 VDD.n4825 VDD.n4824 2.2505
R27663 VDD.n4826 VDD.n4723 2.2505
R27664 VDD.n4828 VDD.n4827 2.2505
R27665 VDD.n4829 VDD.n4722 2.2505
R27666 VDD.n4831 VDD.n4830 2.2505
R27667 VDD.n4832 VDD.n4721 2.2505
R27668 VDD.n4834 VDD.n4833 2.2505
R27669 VDD.n4835 VDD.n4720 2.2505
R27670 VDD.n4837 VDD.n4836 2.2505
R27671 VDD.n4838 VDD.n4719 2.2505
R27672 VDD.n4840 VDD.n4839 2.2505
R27673 VDD.n4841 VDD.n4718 2.2505
R27674 VDD.n4843 VDD.n4842 2.2505
R27675 VDD.n4844 VDD.n4717 2.2505
R27676 VDD.n4846 VDD.n4845 2.2505
R27677 VDD.n4847 VDD.n4716 2.2505
R27678 VDD.n4849 VDD.n4848 2.2505
R27679 VDD.n4850 VDD.n4715 2.2505
R27680 VDD.n4852 VDD.n4851 2.2505
R27681 VDD.n4853 VDD.n4714 2.2505
R27682 VDD.n4855 VDD.n4854 2.2505
R27683 VDD.n4856 VDD.n4713 2.2505
R27684 VDD.n4858 VDD.n4857 2.2505
R27685 VDD.n4859 VDD.n4712 2.2505
R27686 VDD.n4861 VDD.n4860 2.2505
R27687 VDD.n4862 VDD.n4711 2.2505
R27688 VDD.n4864 VDD.n4863 2.2505
R27689 VDD.n4865 VDD.n4710 2.2505
R27690 VDD.n4867 VDD.n4866 2.2505
R27691 VDD.n4868 VDD.n4709 2.2505
R27692 VDD.n4870 VDD.n4869 2.2505
R27693 VDD.n4871 VDD.n4708 2.2505
R27694 VDD.n4873 VDD.n4872 2.2505
R27695 VDD.n4874 VDD.n4707 2.2505
R27696 VDD.n4876 VDD.n4875 2.2505
R27697 VDD.n4877 VDD.n4706 2.2505
R27698 VDD.n4879 VDD.n4878 2.2505
R27699 VDD.n4880 VDD.n4705 2.2505
R27700 VDD.n4882 VDD.n4881 2.2505
R27701 VDD.n4883 VDD.n4704 2.2505
R27702 VDD.n4885 VDD.n4884 2.2505
R27703 VDD.n4886 VDD.n4703 2.2505
R27704 VDD.n4888 VDD.n4887 2.2505
R27705 VDD.n4889 VDD.n4702 2.2505
R27706 VDD.n4891 VDD.n4890 2.2505
R27707 VDD.n4892 VDD.n4701 2.2505
R27708 VDD.n4894 VDD.n4893 2.2505
R27709 VDD.n4895 VDD.n4700 2.2505
R27710 VDD.n4897 VDD.n4896 2.2505
R27711 VDD.n4898 VDD.n4699 2.2505
R27712 VDD.n4900 VDD.n4899 2.2505
R27713 VDD.n4901 VDD.n4698 2.2505
R27714 VDD.n4903 VDD.n4902 2.2505
R27715 VDD.n4904 VDD.n4697 2.2505
R27716 VDD.n7748 VDD.n2269 2.2505
R27717 VDD.n7747 VDD.n7746 2.2505
R27718 VDD.n7745 VDD.n7744 2.2505
R27719 VDD.n7743 VDD.n2271 2.2505
R27720 VDD.n7742 VDD.n7741 2.2505
R27721 VDD.n7740 VDD.n7739 2.2505
R27722 VDD.n7738 VDD.n2273 2.2505
R27723 VDD.n7737 VDD.n7736 2.2505
R27724 VDD.n7735 VDD.n2274 2.2505
R27725 VDD.n7734 VDD.n7733 2.2505
R27726 VDD.n7732 VDD.n2275 2.2505
R27727 VDD.n7731 VDD.n7730 2.2505
R27728 VDD.n7729 VDD.n2276 2.2505
R27729 VDD.n7728 VDD.n7727 2.2505
R27730 VDD.n7726 VDD.n2277 2.2505
R27731 VDD.n7724 VDD.n7723 2.2505
R27732 VDD.n7722 VDD.n2278 2.2505
R27733 VDD.n7721 VDD.n7720 2.2505
R27734 VDD.n7718 VDD.n2279 2.2505
R27735 VDD.n7717 VDD.n7716 2.2505
R27736 VDD.n7715 VDD.n2280 2.2505
R27737 VDD.n7714 VDD.n7713 2.2505
R27738 VDD.n7712 VDD.n2281 2.2505
R27739 VDD.n7711 VDD.n7710 2.2505
R27740 VDD.n7709 VDD.n7708 2.2505
R27741 VDD.n7707 VDD.n2284 2.2505
R27742 VDD.n7706 VDD.n7705 2.2505
R27743 VDD.n7704 VDD.n2285 2.2505
R27744 VDD.n7703 VDD.n7702 2.2505
R27745 VDD.n7701 VDD.n2286 2.2505
R27746 VDD.n7699 VDD.n7698 2.2505
R27747 VDD.n7697 VDD.n2287 2.2505
R27748 VDD.n7696 VDD.n7695 2.2505
R27749 VDD.n7694 VDD.n2288 2.2505
R27750 VDD.n7693 VDD.n7692 2.2505
R27751 VDD.n7691 VDD.n2289 2.2505
R27752 VDD.n7690 VDD.n7689 2.2505
R27753 VDD.n7688 VDD.n2290 2.2505
R27754 VDD.n7687 VDD.n7686 2.2505
R27755 VDD.n10760 VDD.n8254 2.2505
R27756 VDD.n10759 VDD.n10758 2.2505
R27757 VDD.n10150 VDD.n10149 2.2505
R27758 VDD.n10151 VDD.n8457 2.2505
R27759 VDD.n10153 VDD.n10152 2.2505
R27760 VDD.n10154 VDD.n8456 2.2505
R27761 VDD.n10156 VDD.n10155 2.2505
R27762 VDD.n10157 VDD.n8455 2.2505
R27763 VDD.n10159 VDD.n10158 2.2505
R27764 VDD.n10160 VDD.n8454 2.2505
R27765 VDD.n10162 VDD.n10161 2.2505
R27766 VDD.n10163 VDD.n8453 2.2505
R27767 VDD.n10165 VDD.n10164 2.2505
R27768 VDD.n10166 VDD.n8452 2.2505
R27769 VDD.n10168 VDD.n10167 2.2505
R27770 VDD.n10169 VDD.n8451 2.2505
R27771 VDD.n10171 VDD.n10170 2.2505
R27772 VDD.n10172 VDD.n8450 2.2505
R27773 VDD.n10174 VDD.n10173 2.2505
R27774 VDD.n10175 VDD.n8449 2.2505
R27775 VDD.n10177 VDD.n10176 2.2505
R27776 VDD.n10178 VDD.n8448 2.2505
R27777 VDD.n10180 VDD.n10179 2.2505
R27778 VDD.n10181 VDD.n8447 2.2505
R27779 VDD.n10183 VDD.n10182 2.2505
R27780 VDD.n10184 VDD.n8446 2.2505
R27781 VDD.n10186 VDD.n10185 2.2505
R27782 VDD.n10187 VDD.n8445 2.2505
R27783 VDD.n10189 VDD.n10188 2.2505
R27784 VDD.n10190 VDD.n8444 2.2505
R27785 VDD.n10192 VDD.n10191 2.2505
R27786 VDD.n10193 VDD.n8443 2.2505
R27787 VDD.n10195 VDD.n10194 2.2505
R27788 VDD.n10196 VDD.n8442 2.2505
R27789 VDD.n10198 VDD.n10197 2.2505
R27790 VDD.n10199 VDD.n8441 2.2505
R27791 VDD.n10201 VDD.n10200 2.2505
R27792 VDD.n10202 VDD.n8440 2.2505
R27793 VDD.n10204 VDD.n10203 2.2505
R27794 VDD.n10205 VDD.n8439 2.2505
R27795 VDD.n10207 VDD.n10206 2.2505
R27796 VDD.n10208 VDD.n8438 2.2505
R27797 VDD.n10210 VDD.n10209 2.2505
R27798 VDD.n10211 VDD.n8437 2.2505
R27799 VDD.n10213 VDD.n10212 2.2505
R27800 VDD.n10214 VDD.n8436 2.2505
R27801 VDD.n10216 VDD.n10215 2.2505
R27802 VDD.n10217 VDD.n8435 2.2505
R27803 VDD.n10219 VDD.n10218 2.2505
R27804 VDD.n10220 VDD.n8434 2.2505
R27805 VDD.n10222 VDD.n10221 2.2505
R27806 VDD.n10223 VDD.n8433 2.2505
R27807 VDD.n10225 VDD.n10224 2.2505
R27808 VDD.n10226 VDD.n8432 2.2505
R27809 VDD.n10228 VDD.n10227 2.2505
R27810 VDD.n10229 VDD.n8431 2.2505
R27811 VDD.n10231 VDD.n10230 2.2505
R27812 VDD.n10232 VDD.n8430 2.2505
R27813 VDD.n10234 VDD.n10233 2.2505
R27814 VDD.n10235 VDD.n8429 2.2505
R27815 VDD.n10237 VDD.n10236 2.2505
R27816 VDD.n10238 VDD.n8428 2.2505
R27817 VDD.n10240 VDD.n10239 2.2505
R27818 VDD.n10241 VDD.n8427 2.2505
R27819 VDD.n10243 VDD.n10242 2.2505
R27820 VDD.n10244 VDD.n8426 2.2505
R27821 VDD.n10246 VDD.n10245 2.2505
R27822 VDD.n10247 VDD.n8425 2.2505
R27823 VDD.n10249 VDD.n10248 2.2505
R27824 VDD.n10250 VDD.n8424 2.2505
R27825 VDD.n10252 VDD.n10251 2.2505
R27826 VDD.n10253 VDD.n8423 2.2505
R27827 VDD.n10255 VDD.n10254 2.2505
R27828 VDD.n10256 VDD.n8422 2.2505
R27829 VDD.n10258 VDD.n10257 2.2505
R27830 VDD.n10259 VDD.n8421 2.2505
R27831 VDD.n10261 VDD.n10260 2.2505
R27832 VDD.n10262 VDD.n8420 2.2505
R27833 VDD.n10264 VDD.n10263 2.2505
R27834 VDD.n10265 VDD.n8419 2.2505
R27835 VDD.n10267 VDD.n10266 2.2505
R27836 VDD.n10268 VDD.n8418 2.2505
R27837 VDD.n10270 VDD.n10269 2.2505
R27838 VDD.n10271 VDD.n8417 2.2505
R27839 VDD.n10273 VDD.n10272 2.2505
R27840 VDD.n10274 VDD.n8416 2.2505
R27841 VDD.n10276 VDD.n10275 2.2505
R27842 VDD.n10277 VDD.n8415 2.2505
R27843 VDD.n10279 VDD.n10278 2.2505
R27844 VDD.n10280 VDD.n8414 2.2505
R27845 VDD.n10282 VDD.n10281 2.2505
R27846 VDD.n10283 VDD.n8413 2.2505
R27847 VDD.n10285 VDD.n10284 2.2505
R27848 VDD.n10286 VDD.n8412 2.2505
R27849 VDD.n10288 VDD.n10287 2.2505
R27850 VDD.n10289 VDD.n8411 2.2505
R27851 VDD.n10291 VDD.n10290 2.2505
R27852 VDD.n10292 VDD.n8410 2.2505
R27853 VDD.n10294 VDD.n10293 2.2505
R27854 VDD.n10295 VDD.n8409 2.2505
R27855 VDD.n10297 VDD.n10296 2.2505
R27856 VDD.n10298 VDD.n8408 2.2505
R27857 VDD.n10300 VDD.n10299 2.2505
R27858 VDD.n10301 VDD.n8407 2.2505
R27859 VDD.n10303 VDD.n10302 2.2505
R27860 VDD.n10304 VDD.n8406 2.2505
R27861 VDD.n10306 VDD.n10305 2.2505
R27862 VDD.n10307 VDD.n8405 2.2505
R27863 VDD.n10309 VDD.n10308 2.2505
R27864 VDD.n10310 VDD.n8404 2.2505
R27865 VDD.n10312 VDD.n10311 2.2505
R27866 VDD.n10313 VDD.n8403 2.2505
R27867 VDD.n10315 VDD.n10314 2.2505
R27868 VDD.n10316 VDD.n8402 2.2505
R27869 VDD.n10318 VDD.n10317 2.2505
R27870 VDD.n10319 VDD.n8401 2.2505
R27871 VDD.n10321 VDD.n10320 2.2505
R27872 VDD.n10322 VDD.n8400 2.2505
R27873 VDD.n10324 VDD.n10323 2.2505
R27874 VDD.n10325 VDD.n8399 2.2505
R27875 VDD.n10327 VDD.n10326 2.2505
R27876 VDD.n10328 VDD.n8398 2.2505
R27877 VDD.n10330 VDD.n10329 2.2505
R27878 VDD.n10331 VDD.n8397 2.2505
R27879 VDD.n10333 VDD.n10332 2.2505
R27880 VDD.n10334 VDD.n8396 2.2505
R27881 VDD.n10336 VDD.n10335 2.2505
R27882 VDD.n10337 VDD.n8395 2.2505
R27883 VDD.n10339 VDD.n10338 2.2505
R27884 VDD.n10340 VDD.n8394 2.2505
R27885 VDD.n10342 VDD.n10341 2.2505
R27886 VDD.n10343 VDD.n8393 2.2505
R27887 VDD.n10345 VDD.n10344 2.2505
R27888 VDD.n10346 VDD.n8392 2.2505
R27889 VDD.n10348 VDD.n10347 2.2505
R27890 VDD.n10349 VDD.n8391 2.2505
R27891 VDD.n10351 VDD.n10350 2.2505
R27892 VDD.n10352 VDD.n8390 2.2505
R27893 VDD.n10354 VDD.n10353 2.2505
R27894 VDD.n10355 VDD.n8389 2.2505
R27895 VDD.n10357 VDD.n10356 2.2505
R27896 VDD.n10358 VDD.n8388 2.2505
R27897 VDD.n10360 VDD.n10359 2.2505
R27898 VDD.n10361 VDD.n8387 2.2505
R27899 VDD.n10363 VDD.n10362 2.2505
R27900 VDD.n10364 VDD.n8386 2.2505
R27901 VDD.n10366 VDD.n10365 2.2505
R27902 VDD.n10367 VDD.n8385 2.2505
R27903 VDD.n10369 VDD.n10368 2.2505
R27904 VDD.n10370 VDD.n8384 2.2505
R27905 VDD.n10372 VDD.n10371 2.2505
R27906 VDD.n10373 VDD.n8383 2.2505
R27907 VDD.n10375 VDD.n10374 2.2505
R27908 VDD.n10376 VDD.n8382 2.2505
R27909 VDD.n10378 VDD.n10377 2.2505
R27910 VDD.n10379 VDD.n8381 2.2505
R27911 VDD.n10381 VDD.n10380 2.2505
R27912 VDD.n10382 VDD.n8380 2.2505
R27913 VDD.n10384 VDD.n10383 2.2505
R27914 VDD.n10385 VDD.n8379 2.2505
R27915 VDD.n10387 VDD.n10386 2.2505
R27916 VDD.n10388 VDD.n8378 2.2505
R27917 VDD.n10390 VDD.n10389 2.2505
R27918 VDD.n10391 VDD.n8377 2.2505
R27919 VDD.n10393 VDD.n10392 2.2505
R27920 VDD.n10394 VDD.n8376 2.2505
R27921 VDD.n10396 VDD.n10395 2.2505
R27922 VDD.n10397 VDD.n8375 2.2505
R27923 VDD.n10399 VDD.n10398 2.2505
R27924 VDD.n10400 VDD.n8374 2.2505
R27925 VDD.n10402 VDD.n10401 2.2505
R27926 VDD.n10403 VDD.n8373 2.2505
R27927 VDD.n10405 VDD.n10404 2.2505
R27928 VDD.n10406 VDD.n8372 2.2505
R27929 VDD.n10408 VDD.n10407 2.2505
R27930 VDD.n10409 VDD.n8371 2.2505
R27931 VDD.n10411 VDD.n10410 2.2505
R27932 VDD.n10412 VDD.n8370 2.2505
R27933 VDD.n10414 VDD.n10413 2.2505
R27934 VDD.n10415 VDD.n8369 2.2505
R27935 VDD.n10417 VDD.n10416 2.2505
R27936 VDD.n10418 VDD.n8368 2.2505
R27937 VDD.n10420 VDD.n10419 2.2505
R27938 VDD.n10421 VDD.n8367 2.2505
R27939 VDD.n10423 VDD.n10422 2.2505
R27940 VDD.n10424 VDD.n8366 2.2505
R27941 VDD.n10426 VDD.n10425 2.2505
R27942 VDD.n10427 VDD.n8365 2.2505
R27943 VDD.n10429 VDD.n10428 2.2505
R27944 VDD.n10430 VDD.n8364 2.2505
R27945 VDD.n10432 VDD.n10431 2.2505
R27946 VDD.n10433 VDD.n8363 2.2505
R27947 VDD.n10435 VDD.n10434 2.2505
R27948 VDD.n10436 VDD.n8362 2.2505
R27949 VDD.n10438 VDD.n10437 2.2505
R27950 VDD.n10439 VDD.n8361 2.2505
R27951 VDD.n10441 VDD.n10440 2.2505
R27952 VDD.n10442 VDD.n8360 2.2505
R27953 VDD.n10444 VDD.n10443 2.2505
R27954 VDD.n10445 VDD.n8359 2.2505
R27955 VDD.n10447 VDD.n10446 2.2505
R27956 VDD.n10448 VDD.n8358 2.2505
R27957 VDD.n10450 VDD.n10449 2.2505
R27958 VDD.n10451 VDD.n8357 2.2505
R27959 VDD.n10453 VDD.n10452 2.2505
R27960 VDD.n10454 VDD.n8356 2.2505
R27961 VDD.n10456 VDD.n10455 2.2505
R27962 VDD.n10457 VDD.n8355 2.2505
R27963 VDD.n10459 VDD.n10458 2.2505
R27964 VDD.n10460 VDD.n8354 2.2505
R27965 VDD.n10462 VDD.n10461 2.2505
R27966 VDD.n10463 VDD.n8353 2.2505
R27967 VDD.n10465 VDD.n10464 2.2505
R27968 VDD.n10466 VDD.n8352 2.2505
R27969 VDD.n10468 VDD.n10467 2.2505
R27970 VDD.n10469 VDD.n8351 2.2505
R27971 VDD.n10471 VDD.n10470 2.2505
R27972 VDD.n10472 VDD.n8350 2.2505
R27973 VDD.n10474 VDD.n10473 2.2505
R27974 VDD.n10475 VDD.n8349 2.2505
R27975 VDD.n10477 VDD.n10476 2.2505
R27976 VDD.n10478 VDD.n8348 2.2505
R27977 VDD.n10480 VDD.n10479 2.2505
R27978 VDD.n10481 VDD.n8347 2.2505
R27979 VDD.n10483 VDD.n10482 2.2505
R27980 VDD.n10484 VDD.n8346 2.2505
R27981 VDD.n10486 VDD.n10485 2.2505
R27982 VDD.n10487 VDD.n8345 2.2505
R27983 VDD.n10489 VDD.n10488 2.2505
R27984 VDD.n10490 VDD.n8344 2.2505
R27985 VDD.n10492 VDD.n10491 2.2505
R27986 VDD.n10493 VDD.n8343 2.2505
R27987 VDD.n10495 VDD.n10494 2.2505
R27988 VDD.n10496 VDD.n8342 2.2505
R27989 VDD.n10498 VDD.n10497 2.2505
R27990 VDD.n10499 VDD.n8341 2.2505
R27991 VDD.n10501 VDD.n10500 2.2505
R27992 VDD.n10502 VDD.n8340 2.2505
R27993 VDD.n10504 VDD.n10503 2.2505
R27994 VDD.n10505 VDD.n8339 2.2505
R27995 VDD.n10507 VDD.n10506 2.2505
R27996 VDD.n10508 VDD.n8338 2.2505
R27997 VDD.n10510 VDD.n10509 2.2505
R27998 VDD.n10511 VDD.n8337 2.2505
R27999 VDD.n10513 VDD.n10512 2.2505
R28000 VDD.n10514 VDD.n8336 2.2505
R28001 VDD.n10516 VDD.n10515 2.2505
R28002 VDD.n10517 VDD.n8335 2.2505
R28003 VDD.n10519 VDD.n10518 2.2505
R28004 VDD.n10520 VDD.n8334 2.2505
R28005 VDD.n10522 VDD.n10521 2.2505
R28006 VDD.n10523 VDD.n8333 2.2505
R28007 VDD.n10525 VDD.n10524 2.2505
R28008 VDD.n10526 VDD.n8332 2.2505
R28009 VDD.n10528 VDD.n10527 2.2505
R28010 VDD.n10529 VDD.n8331 2.2505
R28011 VDD.n10531 VDD.n10530 2.2505
R28012 VDD.n10532 VDD.n8330 2.2505
R28013 VDD.n10534 VDD.n10533 2.2505
R28014 VDD.n10535 VDD.n8329 2.2505
R28015 VDD.n10537 VDD.n10536 2.2505
R28016 VDD.n10538 VDD.n8328 2.2505
R28017 VDD.n10540 VDD.n10539 2.2505
R28018 VDD.n10541 VDD.n8327 2.2505
R28019 VDD.n10543 VDD.n10542 2.2505
R28020 VDD.n10544 VDD.n8326 2.2505
R28021 VDD.n10546 VDD.n10545 2.2505
R28022 VDD.n10547 VDD.n8325 2.2505
R28023 VDD.n10549 VDD.n10548 2.2505
R28024 VDD.n10550 VDD.n8324 2.2505
R28025 VDD.n10552 VDD.n10551 2.2505
R28026 VDD.n10553 VDD.n8323 2.2505
R28027 VDD.n10555 VDD.n10554 2.2505
R28028 VDD.n10556 VDD.n8322 2.2505
R28029 VDD.n10558 VDD.n10557 2.2505
R28030 VDD.n10559 VDD.n8321 2.2505
R28031 VDD.n10561 VDD.n10560 2.2505
R28032 VDD.n10562 VDD.n8320 2.2505
R28033 VDD.n10564 VDD.n10563 2.2505
R28034 VDD.n10565 VDD.n8319 2.2505
R28035 VDD.n10567 VDD.n10566 2.2505
R28036 VDD.n10568 VDD.n8318 2.2505
R28037 VDD.n10570 VDD.n10569 2.2505
R28038 VDD.n10571 VDD.n8317 2.2505
R28039 VDD.n10573 VDD.n10572 2.2505
R28040 VDD.n10574 VDD.n8316 2.2505
R28041 VDD.n10576 VDD.n10575 2.2505
R28042 VDD.n10577 VDD.n8315 2.2505
R28043 VDD.n10579 VDD.n10578 2.2505
R28044 VDD.n10580 VDD.n8314 2.2505
R28045 VDD.n10582 VDD.n10581 2.2505
R28046 VDD.n10583 VDD.n8313 2.2505
R28047 VDD.n10585 VDD.n10584 2.2505
R28048 VDD.n10586 VDD.n8312 2.2505
R28049 VDD.n10588 VDD.n10587 2.2505
R28050 VDD.n10589 VDD.n8311 2.2505
R28051 VDD.n10591 VDD.n10590 2.2505
R28052 VDD.n10592 VDD.n8310 2.2505
R28053 VDD.n10594 VDD.n10593 2.2505
R28054 VDD.n10595 VDD.n8309 2.2505
R28055 VDD.n10597 VDD.n10596 2.2505
R28056 VDD.n10598 VDD.n8308 2.2505
R28057 VDD.n10600 VDD.n10599 2.2505
R28058 VDD.n10601 VDD.n8307 2.2505
R28059 VDD.n10603 VDD.n10602 2.2505
R28060 VDD.n10604 VDD.n8306 2.2505
R28061 VDD.n10606 VDD.n10605 2.2505
R28062 VDD.n10607 VDD.n8305 2.2505
R28063 VDD.n10609 VDD.n10608 2.2505
R28064 VDD.n10610 VDD.n8304 2.2505
R28065 VDD.n10612 VDD.n10611 2.2505
R28066 VDD.n10613 VDD.n8303 2.2505
R28067 VDD.n10615 VDD.n10614 2.2505
R28068 VDD.n10616 VDD.n8302 2.2505
R28069 VDD.n10618 VDD.n10617 2.2505
R28070 VDD.n10619 VDD.n8301 2.2505
R28071 VDD.n10621 VDD.n10620 2.2505
R28072 VDD.n10622 VDD.n8300 2.2505
R28073 VDD.n10624 VDD.n10623 2.2505
R28074 VDD.n10625 VDD.n8299 2.2505
R28075 VDD.n10627 VDD.n10626 2.2505
R28076 VDD.n10628 VDD.n8298 2.2505
R28077 VDD.n10630 VDD.n10629 2.2505
R28078 VDD.n10631 VDD.n8297 2.2505
R28079 VDD.n10633 VDD.n10632 2.2505
R28080 VDD.n10634 VDD.n8296 2.2505
R28081 VDD.n10636 VDD.n10635 2.2505
R28082 VDD.n10637 VDD.n8295 2.2505
R28083 VDD.n10639 VDD.n10638 2.2505
R28084 VDD.n10640 VDD.n8294 2.2505
R28085 VDD.n10642 VDD.n10641 2.2505
R28086 VDD.n10643 VDD.n8293 2.2505
R28087 VDD.n10645 VDD.n10644 2.2505
R28088 VDD.n10646 VDD.n8292 2.2505
R28089 VDD.n10648 VDD.n10647 2.2505
R28090 VDD.n10649 VDD.n8291 2.2505
R28091 VDD.n10651 VDD.n10650 2.2505
R28092 VDD.n10652 VDD.n8290 2.2505
R28093 VDD.n10654 VDD.n10653 2.2505
R28094 VDD.n10655 VDD.n8289 2.2505
R28095 VDD.n10657 VDD.n10656 2.2505
R28096 VDD.n10658 VDD.n8288 2.2505
R28097 VDD.n10660 VDD.n10659 2.2505
R28098 VDD.n10661 VDD.n8287 2.2505
R28099 VDD.n10663 VDD.n10662 2.2505
R28100 VDD.n10664 VDD.n8286 2.2505
R28101 VDD.n10666 VDD.n10665 2.2505
R28102 VDD.n10667 VDD.n8285 2.2505
R28103 VDD.n10669 VDD.n10668 2.2505
R28104 VDD.n10670 VDD.n8284 2.2505
R28105 VDD.n10672 VDD.n10671 2.2505
R28106 VDD.n10673 VDD.n8283 2.2505
R28107 VDD.n10675 VDD.n10674 2.2505
R28108 VDD.n10676 VDD.n8282 2.2505
R28109 VDD.n10678 VDD.n10677 2.2505
R28110 VDD.n10679 VDD.n8281 2.2505
R28111 VDD.n10681 VDD.n10680 2.2505
R28112 VDD.n10682 VDD.n8280 2.2505
R28113 VDD.n10684 VDD.n10683 2.2505
R28114 VDD.n10685 VDD.n8279 2.2505
R28115 VDD.n10687 VDD.n10686 2.2505
R28116 VDD.n10688 VDD.n8278 2.2505
R28117 VDD.n10690 VDD.n10689 2.2505
R28118 VDD.n10691 VDD.n8277 2.2505
R28119 VDD.n10693 VDD.n10692 2.2505
R28120 VDD.n10694 VDD.n8276 2.2505
R28121 VDD.n10696 VDD.n10695 2.2505
R28122 VDD.n10697 VDD.n8275 2.2505
R28123 VDD.n10699 VDD.n10698 2.2505
R28124 VDD.n10700 VDD.n8274 2.2505
R28125 VDD.n10702 VDD.n10701 2.2505
R28126 VDD.n10703 VDD.n8273 2.2505
R28127 VDD.n10705 VDD.n10704 2.2505
R28128 VDD.n10706 VDD.n8272 2.2505
R28129 VDD.n10708 VDD.n10707 2.2505
R28130 VDD.n10709 VDD.n8271 2.2505
R28131 VDD.n10711 VDD.n10710 2.2505
R28132 VDD.n10712 VDD.n8270 2.2505
R28133 VDD.n10714 VDD.n10713 2.2505
R28134 VDD.n10715 VDD.n8269 2.2505
R28135 VDD.n10717 VDD.n10716 2.2505
R28136 VDD.n10718 VDD.n8268 2.2505
R28137 VDD.n10720 VDD.n10719 2.2505
R28138 VDD.n10721 VDD.n8267 2.2505
R28139 VDD.n10723 VDD.n10722 2.2505
R28140 VDD.n10724 VDD.n8266 2.2505
R28141 VDD.n10726 VDD.n10725 2.2505
R28142 VDD.n10727 VDD.n8265 2.2505
R28143 VDD.n10729 VDD.n10728 2.2505
R28144 VDD.n10730 VDD.n8264 2.2505
R28145 VDD.n10732 VDD.n10731 2.2505
R28146 VDD.n10733 VDD.n8263 2.2505
R28147 VDD.n10735 VDD.n10734 2.2505
R28148 VDD.n10736 VDD.n8262 2.2505
R28149 VDD.n10738 VDD.n10737 2.2505
R28150 VDD.n10739 VDD.n8261 2.2505
R28151 VDD.n10741 VDD.n10740 2.2505
R28152 VDD.n10742 VDD.n8260 2.2505
R28153 VDD.n10744 VDD.n10743 2.2505
R28154 VDD.n10745 VDD.n8259 2.2505
R28155 VDD.n10747 VDD.n10746 2.2505
R28156 VDD.n10748 VDD.n8258 2.2505
R28157 VDD.n10750 VDD.n10749 2.2505
R28158 VDD.n10751 VDD.n8257 2.2505
R28159 VDD.n10753 VDD.n10752 2.2505
R28160 VDD.n10754 VDD.n8256 2.2505
R28161 VDD.n10756 VDD.n10755 2.2505
R28162 VDD.n10757 VDD.n8255 2.2505
R28163 VDD.n10103 VDD.n9214 2.2505
R28164 VDD.n10105 VDD.n10104 2.2505
R28165 VDD.n10106 VDD.n9213 2.2505
R28166 VDD.n10108 VDD.n10107 2.2505
R28167 VDD.n10109 VDD.n9212 2.2505
R28168 VDD.n10111 VDD.n10110 2.2505
R28169 VDD.n10112 VDD.n9211 2.2505
R28170 VDD.n10114 VDD.n10113 2.2505
R28171 VDD.n10115 VDD.n9210 2.2505
R28172 VDD.n10117 VDD.n10116 2.2505
R28173 VDD.n10118 VDD.n9209 2.2505
R28174 VDD.n10120 VDD.n10119 2.2505
R28175 VDD.n10121 VDD.n9208 2.2505
R28176 VDD.n10123 VDD.n10122 2.2505
R28177 VDD.n10124 VDD.n9207 2.2505
R28178 VDD.n10126 VDD.n10125 2.2505
R28179 VDD.n10127 VDD.n9206 2.2505
R28180 VDD.n10129 VDD.n10128 2.2505
R28181 VDD.n10130 VDD.n9205 2.2505
R28182 VDD.n10132 VDD.n10131 2.2505
R28183 VDD.n10133 VDD.n9204 2.2505
R28184 VDD.n10135 VDD.n10134 2.2505
R28185 VDD.n10136 VDD.n9203 2.2505
R28186 VDD.n10138 VDD.n10137 2.2505
R28187 VDD.n10139 VDD.n9202 2.2505
R28188 VDD.n10141 VDD.n10140 2.2505
R28189 VDD.n10142 VDD.n9201 2.2505
R28190 VDD.n10144 VDD.n10143 2.2505
R28191 VDD.n10145 VDD.n9186 2.2505
R28192 VDD.n10147 VDD.n10146 2.2505
R28193 VDD.n10102 VDD.n10101 2.2505
R28194 VDD.n10100 VDD.n9215 2.2505
R28195 VDD.n10099 VDD.n10098 2.2505
R28196 VDD.n10097 VDD.n9216 2.2505
R28197 VDD.n10096 VDD.n10095 2.2505
R28198 VDD.n10094 VDD.n9217 2.2505
R28199 VDD.n10093 VDD.n10092 2.2505
R28200 VDD.n10091 VDD.n9218 2.2505
R28201 VDD.n10090 VDD.n10089 2.2505
R28202 VDD.n10088 VDD.n9219 2.2505
R28203 VDD.n10087 VDD.n10086 2.2505
R28204 VDD.n10085 VDD.n9220 2.2505
R28205 VDD.n10084 VDD.n10083 2.2505
R28206 VDD.n10082 VDD.n9221 2.2505
R28207 VDD.n10081 VDD.n10080 2.2505
R28208 VDD.n10079 VDD.n9222 2.2505
R28209 VDD.n10078 VDD.n10077 2.2505
R28210 VDD.n10076 VDD.n9223 2.2505
R28211 VDD.n10075 VDD.n10074 2.2505
R28212 VDD.n10073 VDD.n9224 2.2505
R28213 VDD.n10072 VDD.n10071 2.2505
R28214 VDD.n10070 VDD.n9225 2.2505
R28215 VDD.n10069 VDD.n10068 2.2505
R28216 VDD.n10067 VDD.n9226 2.2505
R28217 VDD.n10066 VDD.n10065 2.2505
R28218 VDD.n10064 VDD.n9227 2.2505
R28219 VDD.n10063 VDD.n10062 2.2505
R28220 VDD.n10061 VDD.n9228 2.2505
R28221 VDD.n10060 VDD.n10059 2.2505
R28222 VDD.n10058 VDD.n9229 2.2505
R28223 VDD.n10057 VDD.n10056 2.2505
R28224 VDD.n10055 VDD.n9230 2.2505
R28225 VDD.n10054 VDD.n10053 2.2505
R28226 VDD.n10052 VDD.n9231 2.2505
R28227 VDD.n10051 VDD.n10050 2.2505
R28228 VDD.n10049 VDD.n9232 2.2505
R28229 VDD.n10048 VDD.n10047 2.2505
R28230 VDD.n10046 VDD.n9233 2.2505
R28231 VDD.n10045 VDD.n10044 2.2505
R28232 VDD.n10043 VDD.n9234 2.2505
R28233 VDD.n10042 VDD.n10041 2.2505
R28234 VDD.n10040 VDD.n9235 2.2505
R28235 VDD.n10039 VDD.n10038 2.2505
R28236 VDD.n10037 VDD.n9236 2.2505
R28237 VDD.n10036 VDD.n10035 2.2505
R28238 VDD.n10034 VDD.n9237 2.2505
R28239 VDD.n10033 VDD.n10032 2.2505
R28240 VDD.n10031 VDD.n9238 2.2505
R28241 VDD.n10030 VDD.n10029 2.2505
R28242 VDD.n10028 VDD.n9239 2.2505
R28243 VDD.n10027 VDD.n10026 2.2505
R28244 VDD.n10025 VDD.n9240 2.2505
R28245 VDD.n10024 VDD.n10023 2.2505
R28246 VDD.n10022 VDD.n9241 2.2505
R28247 VDD.n10021 VDD.n10020 2.2505
R28248 VDD.n10019 VDD.n9242 2.2505
R28249 VDD.n10018 VDD.n10017 2.2505
R28250 VDD.n10016 VDD.n9243 2.2505
R28251 VDD.n10015 VDD.n10014 2.2505
R28252 VDD.n10013 VDD.n9244 2.2505
R28253 VDD.n10012 VDD.n10011 2.2505
R28254 VDD.n10010 VDD.n9245 2.2505
R28255 VDD.n10009 VDD.n10008 2.2505
R28256 VDD.n10007 VDD.n9246 2.2505
R28257 VDD.n10006 VDD.n10005 2.2505
R28258 VDD.n10004 VDD.n9247 2.2505
R28259 VDD.n10003 VDD.n10002 2.2505
R28260 VDD.n10001 VDD.n9248 2.2505
R28261 VDD.n10000 VDD.n9999 2.2505
R28262 VDD.n9998 VDD.n9249 2.2505
R28263 VDD.n9997 VDD.n9996 2.2505
R28264 VDD.n9995 VDD.n9250 2.2505
R28265 VDD.n9994 VDD.n9993 2.2505
R28266 VDD.n9992 VDD.n9251 2.2505
R28267 VDD.n9991 VDD.n9990 2.2505
R28268 VDD.n9989 VDD.n9252 2.2505
R28269 VDD.n9988 VDD.n9987 2.2505
R28270 VDD.n9986 VDD.n9253 2.2505
R28271 VDD.n9985 VDD.n9984 2.2505
R28272 VDD.n9983 VDD.n9254 2.2505
R28273 VDD.n9982 VDD.n9981 2.2505
R28274 VDD.n9980 VDD.n9255 2.2505
R28275 VDD.n9979 VDD.n9978 2.2505
R28276 VDD.n9977 VDD.n9256 2.2505
R28277 VDD.n9976 VDD.n9975 2.2505
R28278 VDD.n9974 VDD.n9257 2.2505
R28279 VDD.n9973 VDD.n9972 2.2505
R28280 VDD.n9971 VDD.n9258 2.2505
R28281 VDD.n9970 VDD.n9969 2.2505
R28282 VDD.n9968 VDD.n9259 2.2505
R28283 VDD.n9967 VDD.n9966 2.2505
R28284 VDD.n9965 VDD.n9260 2.2505
R28285 VDD.n9964 VDD.n9963 2.2505
R28286 VDD.n9962 VDD.n9261 2.2505
R28287 VDD.n9961 VDD.n9960 2.2505
R28288 VDD.n9959 VDD.n9262 2.2505
R28289 VDD.n9958 VDD.n9957 2.2505
R28290 VDD.n9956 VDD.n9263 2.2505
R28291 VDD.n9955 VDD.n9954 2.2505
R28292 VDD.n9953 VDD.n9264 2.2505
R28293 VDD.n9952 VDD.n9951 2.2505
R28294 VDD.n9950 VDD.n9265 2.2505
R28295 VDD.n9949 VDD.n9948 2.2505
R28296 VDD.n9947 VDD.n9266 2.2505
R28297 VDD.n9946 VDD.n9945 2.2505
R28298 VDD.n9944 VDD.n9267 2.2505
R28299 VDD.n9943 VDD.n9942 2.2505
R28300 VDD.n9941 VDD.n9268 2.2505
R28301 VDD.n9940 VDD.n9939 2.2505
R28302 VDD.n9938 VDD.n9269 2.2505
R28303 VDD.n9937 VDD.n9936 2.2505
R28304 VDD.n9935 VDD.n9270 2.2505
R28305 VDD.n9934 VDD.n9933 2.2505
R28306 VDD.n9932 VDD.n9271 2.2505
R28307 VDD.n9931 VDD.n9930 2.2505
R28308 VDD.n9929 VDD.n9272 2.2505
R28309 VDD.n9928 VDD.n9927 2.2505
R28310 VDD.n9926 VDD.n9273 2.2505
R28311 VDD.n9925 VDD.n9924 2.2505
R28312 VDD.n9923 VDD.n9274 2.2505
R28313 VDD.n9922 VDD.n9921 2.2505
R28314 VDD.n9920 VDD.n9275 2.2505
R28315 VDD.n9919 VDD.n9918 2.2505
R28316 VDD.n9917 VDD.n9276 2.2505
R28317 VDD.n9916 VDD.n9915 2.2505
R28318 VDD.n9914 VDD.n9277 2.2505
R28319 VDD.n9913 VDD.n9912 2.2505
R28320 VDD.n9911 VDD.n9278 2.2505
R28321 VDD.n9910 VDD.n9909 2.2505
R28322 VDD.n9908 VDD.n9279 2.2505
R28323 VDD.n9907 VDD.n9906 2.2505
R28324 VDD.n9905 VDD.n9280 2.2505
R28325 VDD.n9904 VDD.n9903 2.2505
R28326 VDD.n9902 VDD.n9281 2.2505
R28327 VDD.n9901 VDD.n9900 2.2505
R28328 VDD.n9899 VDD.n9282 2.2505
R28329 VDD.n9898 VDD.n9897 2.2505
R28330 VDD.n9896 VDD.n9283 2.2505
R28331 VDD.n9895 VDD.n9894 2.2505
R28332 VDD.n9893 VDD.n9284 2.2505
R28333 VDD.n9892 VDD.n9891 2.2505
R28334 VDD.n9890 VDD.n9285 2.2505
R28335 VDD.n9889 VDD.n9888 2.2505
R28336 VDD.n9887 VDD.n9286 2.2505
R28337 VDD.n9886 VDD.n9885 2.2505
R28338 VDD.n9884 VDD.n9287 2.2505
R28339 VDD.n9883 VDD.n9882 2.2505
R28340 VDD.n9881 VDD.n9288 2.2505
R28341 VDD.n9880 VDD.n9879 2.2505
R28342 VDD.n9878 VDD.n9289 2.2505
R28343 VDD.n9877 VDD.n9876 2.2505
R28344 VDD.n9875 VDD.n9290 2.2505
R28345 VDD.n9874 VDD.n9873 2.2505
R28346 VDD.n9872 VDD.n9291 2.2505
R28347 VDD.n9871 VDD.n9870 2.2505
R28348 VDD.n9869 VDD.n9292 2.2505
R28349 VDD.n9868 VDD.n9867 2.2505
R28350 VDD.n9866 VDD.n9293 2.2505
R28351 VDD.n9865 VDD.n9864 2.2505
R28352 VDD.n9863 VDD.n9294 2.2505
R28353 VDD.n9862 VDD.n9861 2.2505
R28354 VDD.n9860 VDD.n9295 2.2505
R28355 VDD.n9859 VDD.n9858 2.2505
R28356 VDD.n9857 VDD.n9296 2.2505
R28357 VDD.n9856 VDD.n9855 2.2505
R28358 VDD.n9854 VDD.n9297 2.2505
R28359 VDD.n9853 VDD.n9852 2.2505
R28360 VDD.n9851 VDD.n9298 2.2505
R28361 VDD.n9850 VDD.n9849 2.2505
R28362 VDD.n9848 VDD.n9299 2.2505
R28363 VDD.n9847 VDD.n9846 2.2505
R28364 VDD.n9845 VDD.n9300 2.2505
R28365 VDD.n9844 VDD.n9843 2.2505
R28366 VDD.n9842 VDD.n9301 2.2505
R28367 VDD.n9841 VDD.n9840 2.2505
R28368 VDD.n9839 VDD.n9302 2.2505
R28369 VDD.n9838 VDD.n9837 2.2505
R28370 VDD.n9836 VDD.n9303 2.2505
R28371 VDD.n9835 VDD.n9834 2.2505
R28372 VDD.n9833 VDD.n9304 2.2505
R28373 VDD.n9832 VDD.n9831 2.2505
R28374 VDD.n9830 VDD.n9305 2.2505
R28375 VDD.n9829 VDD.n9828 2.2505
R28376 VDD.n9827 VDD.n9306 2.2505
R28377 VDD.n9826 VDD.n9825 2.2505
R28378 VDD.n9824 VDD.n9307 2.2505
R28379 VDD.n9823 VDD.n9822 2.2505
R28380 VDD.n9821 VDD.n9308 2.2505
R28381 VDD.n9820 VDD.n9819 2.2505
R28382 VDD.n9818 VDD.n9309 2.2505
R28383 VDD.n9817 VDD.n9816 2.2505
R28384 VDD.n9815 VDD.n9310 2.2505
R28385 VDD.n9814 VDD.n9813 2.2505
R28386 VDD.n9812 VDD.n9311 2.2505
R28387 VDD.n9811 VDD.n9810 2.2505
R28388 VDD.n9809 VDD.n9312 2.2505
R28389 VDD.n9808 VDD.n9807 2.2505
R28390 VDD.n9806 VDD.n9313 2.2505
R28391 VDD.n9805 VDD.n9804 2.2505
R28392 VDD.n9803 VDD.n9314 2.2505
R28393 VDD.n9802 VDD.n9801 2.2505
R28394 VDD.n9800 VDD.n9315 2.2505
R28395 VDD.n9799 VDD.n9798 2.2505
R28396 VDD.n9797 VDD.n9316 2.2505
R28397 VDD.n9796 VDD.n9795 2.2505
R28398 VDD.n9794 VDD.n9317 2.2505
R28399 VDD.n9793 VDD.n9792 2.2505
R28400 VDD.n9791 VDD.n9318 2.2505
R28401 VDD.n9790 VDD.n9789 2.2505
R28402 VDD.n9788 VDD.n9319 2.2505
R28403 VDD.n9787 VDD.n9786 2.2505
R28404 VDD.n9785 VDD.n9320 2.2505
R28405 VDD.n9784 VDD.n9783 2.2505
R28406 VDD.n9782 VDD.n9321 2.2505
R28407 VDD.n9781 VDD.n9780 2.2505
R28408 VDD.n9779 VDD.n9322 2.2505
R28409 VDD.n9778 VDD.n9777 2.2505
R28410 VDD.n9776 VDD.n9323 2.2505
R28411 VDD.n9775 VDD.n9774 2.2505
R28412 VDD.n9773 VDD.n9324 2.2505
R28413 VDD.n9772 VDD.n9771 2.2505
R28414 VDD.n9770 VDD.n9325 2.2505
R28415 VDD.n9769 VDD.n9768 2.2505
R28416 VDD.n9767 VDD.n9326 2.2505
R28417 VDD.n9766 VDD.n9765 2.2505
R28418 VDD.n9764 VDD.n9327 2.2505
R28419 VDD.n9763 VDD.n9762 2.2505
R28420 VDD.n9761 VDD.n9328 2.2505
R28421 VDD.n9760 VDD.n9759 2.2505
R28422 VDD.n9758 VDD.n9329 2.2505
R28423 VDD.n9757 VDD.n9756 2.2505
R28424 VDD.n9755 VDD.n9330 2.2505
R28425 VDD.n9754 VDD.n9753 2.2505
R28426 VDD.n9752 VDD.n9331 2.2505
R28427 VDD.n9751 VDD.n9750 2.2505
R28428 VDD.n9749 VDD.n9332 2.2505
R28429 VDD.n9748 VDD.n9747 2.2505
R28430 VDD.n9746 VDD.n9333 2.2505
R28431 VDD.n9745 VDD.n9744 2.2505
R28432 VDD.n9743 VDD.n9334 2.2505
R28433 VDD.n9742 VDD.n9741 2.2505
R28434 VDD.n9740 VDD.n9335 2.2505
R28435 VDD.n9739 VDD.n9738 2.2505
R28436 VDD.n9737 VDD.n9336 2.2505
R28437 VDD.n9736 VDD.n9735 2.2505
R28438 VDD.n9734 VDD.n9337 2.2505
R28439 VDD.n9733 VDD.n9732 2.2505
R28440 VDD.n9731 VDD.n9338 2.2505
R28441 VDD.n9730 VDD.n9729 2.2505
R28442 VDD.n9728 VDD.n9339 2.2505
R28443 VDD.n9727 VDD.n9726 2.2505
R28444 VDD.n9725 VDD.n9340 2.2505
R28445 VDD.n9724 VDD.n9723 2.2505
R28446 VDD.n9722 VDD.n9341 2.2505
R28447 VDD.n9721 VDD.n9720 2.2505
R28448 VDD.n9719 VDD.n9342 2.2505
R28449 VDD.n9718 VDD.n9717 2.2505
R28450 VDD.n9716 VDD.n9343 2.2505
R28451 VDD.n9715 VDD.n9714 2.2505
R28452 VDD.n9713 VDD.n9344 2.2505
R28453 VDD.n9712 VDD.n9711 2.2505
R28454 VDD.n9710 VDD.n9345 2.2505
R28455 VDD.n9709 VDD.n9708 2.2505
R28456 VDD.n9707 VDD.n9346 2.2505
R28457 VDD.n9706 VDD.n9705 2.2505
R28458 VDD.n9704 VDD.n9347 2.2505
R28459 VDD.n9703 VDD.n9702 2.2505
R28460 VDD.n9701 VDD.n9348 2.2505
R28461 VDD.n9700 VDD.n9699 2.2505
R28462 VDD.n9698 VDD.n9349 2.2505
R28463 VDD.n9697 VDD.n9696 2.2505
R28464 VDD.n9695 VDD.n9350 2.2505
R28465 VDD.n9694 VDD.n9693 2.2505
R28466 VDD.n9692 VDD.n9351 2.2505
R28467 VDD.n9691 VDD.n9690 2.2505
R28468 VDD.n9689 VDD.n9352 2.2505
R28469 VDD.n9688 VDD.n9687 2.2505
R28470 VDD.n9686 VDD.n9353 2.2505
R28471 VDD.n9685 VDD.n9684 2.2505
R28472 VDD.n9683 VDD.n9354 2.2505
R28473 VDD.n9682 VDD.n9681 2.2505
R28474 VDD.n9680 VDD.n9355 2.2505
R28475 VDD.n9679 VDD.n9678 2.2505
R28476 VDD.n9677 VDD.n9356 2.2505
R28477 VDD.n9676 VDD.n9675 2.2505
R28478 VDD.n9674 VDD.n9357 2.2505
R28479 VDD.n9673 VDD.n9672 2.2505
R28480 VDD.n9671 VDD.n9358 2.2505
R28481 VDD.n9670 VDD.n9669 2.2505
R28482 VDD.n9668 VDD.n9359 2.2505
R28483 VDD.n9667 VDD.n9666 2.2505
R28484 VDD.n9665 VDD.n9360 2.2505
R28485 VDD.n9664 VDD.n9663 2.2505
R28486 VDD.n9662 VDD.n9361 2.2505
R28487 VDD.n9661 VDD.n9660 2.2505
R28488 VDD.n9659 VDD.n9362 2.2505
R28489 VDD.n9658 VDD.n9657 2.2505
R28490 VDD.n9656 VDD.n9363 2.2505
R28491 VDD.n9655 VDD.n9654 2.2505
R28492 VDD.n9653 VDD.n9364 2.2505
R28493 VDD.n9652 VDD.n9651 2.2505
R28494 VDD.n9650 VDD.n9365 2.2505
R28495 VDD.n9649 VDD.n9648 2.2505
R28496 VDD.n9647 VDD.n9366 2.2505
R28497 VDD.n9646 VDD.n9645 2.2505
R28498 VDD.n9644 VDD.n9367 2.2505
R28499 VDD.n9643 VDD.n9642 2.2505
R28500 VDD.n9641 VDD.n9368 2.2505
R28501 VDD.n9640 VDD.n9639 2.2505
R28502 VDD.n9638 VDD.n9369 2.2505
R28503 VDD.n9637 VDD.n9636 2.2505
R28504 VDD.n9635 VDD.n9370 2.2505
R28505 VDD.n9634 VDD.n9633 2.2505
R28506 VDD.n9632 VDD.n9371 2.2505
R28507 VDD.n9631 VDD.n9630 2.2505
R28508 VDD.n9629 VDD.n9372 2.2505
R28509 VDD.n9628 VDD.n9627 2.2505
R28510 VDD.n9626 VDD.n9373 2.2505
R28511 VDD.n9625 VDD.n9624 2.2505
R28512 VDD.n9623 VDD.n9374 2.2505
R28513 VDD.n9622 VDD.n9621 2.2505
R28514 VDD.n9620 VDD.n9375 2.2505
R28515 VDD.n9619 VDD.n9618 2.2505
R28516 VDD.n9617 VDD.n9376 2.2505
R28517 VDD.n9616 VDD.n9615 2.2505
R28518 VDD.n9614 VDD.n9377 2.2505
R28519 VDD.n9613 VDD.n9612 2.2505
R28520 VDD.n9611 VDD.n9378 2.2505
R28521 VDD.n9610 VDD.n9609 2.2505
R28522 VDD.n9608 VDD.n9379 2.2505
R28523 VDD.n9607 VDD.n9606 2.2505
R28524 VDD.n9605 VDD.n9380 2.2505
R28525 VDD.n9604 VDD.n9603 2.2505
R28526 VDD.n9602 VDD.n9381 2.2505
R28527 VDD.n9601 VDD.n9600 2.2505
R28528 VDD.n9599 VDD.n9382 2.2505
R28529 VDD.n9598 VDD.n9597 2.2505
R28530 VDD.n9596 VDD.n9383 2.2505
R28531 VDD.n9595 VDD.n9594 2.2505
R28532 VDD.n9593 VDD.n9384 2.2505
R28533 VDD.n9592 VDD.n9591 2.2505
R28534 VDD.n9590 VDD.n9385 2.2505
R28535 VDD.n9589 VDD.n9588 2.2505
R28536 VDD.n9587 VDD.n9386 2.2505
R28537 VDD.n9586 VDD.n9585 2.2505
R28538 VDD.n9584 VDD.n9387 2.2505
R28539 VDD.n9583 VDD.n9582 2.2505
R28540 VDD.n9581 VDD.n9388 2.2505
R28541 VDD.n9580 VDD.n9579 2.2505
R28542 VDD.n9578 VDD.n9389 2.2505
R28543 VDD.n9577 VDD.n9576 2.2505
R28544 VDD.n9575 VDD.n9390 2.2505
R28545 VDD.n9574 VDD.n9573 2.2505
R28546 VDD.n9572 VDD.n9391 2.2505
R28547 VDD.n9571 VDD.n9570 2.2505
R28548 VDD.n9569 VDD.n9392 2.2505
R28549 VDD.n9568 VDD.n9567 2.2505
R28550 VDD.n9566 VDD.n9393 2.2505
R28551 VDD.n9565 VDD.n9564 2.2505
R28552 VDD.n9563 VDD.n9394 2.2505
R28553 VDD.n9562 VDD.n9561 2.2505
R28554 VDD.n9560 VDD.n9395 2.2505
R28555 VDD.n9559 VDD.n9558 2.2505
R28556 VDD.n9557 VDD.n9396 2.2505
R28557 VDD.n9556 VDD.n9555 2.2505
R28558 VDD.n9554 VDD.n9397 2.2505
R28559 VDD.n9553 VDD.n9552 2.2505
R28560 VDD.n9551 VDD.n9398 2.2505
R28561 VDD.n9550 VDD.n9549 2.2505
R28562 VDD.n9548 VDD.n9399 2.2505
R28563 VDD.n9547 VDD.n9546 2.2505
R28564 VDD.n9545 VDD.n9400 2.2505
R28565 VDD.n9544 VDD.n9543 2.2505
R28566 VDD.n9542 VDD.n9401 2.2505
R28567 VDD.n9541 VDD.n9540 2.2505
R28568 VDD.n9539 VDD.n9402 2.2505
R28569 VDD.n9538 VDD.n9537 2.2505
R28570 VDD.n9536 VDD.n9403 2.2505
R28571 VDD.n9535 VDD.n9534 2.2505
R28572 VDD.n9533 VDD.n9404 2.2505
R28573 VDD.n9532 VDD.n9531 2.2505
R28574 VDD.n9530 VDD.n9405 2.2505
R28575 VDD.n9529 VDD.n9528 2.2505
R28576 VDD.n9527 VDD.n9406 2.2505
R28577 VDD.n9526 VDD.n9525 2.2505
R28578 VDD.n9524 VDD.n9407 2.2505
R28579 VDD.n9523 VDD.n9522 2.2505
R28580 VDD.n9521 VDD.n9408 2.2505
R28581 VDD.n9520 VDD.n9519 2.2505
R28582 VDD.n9518 VDD.n9409 2.2505
R28583 VDD.n9517 VDD.n9516 2.2505
R28584 VDD.n9515 VDD.n9410 2.2505
R28585 VDD.n9514 VDD.n9513 2.2505
R28586 VDD.n9512 VDD.n9411 2.2505
R28587 VDD.n9511 VDD.n9510 2.2505
R28588 VDD.n9509 VDD.n9412 2.2505
R28589 VDD.n9508 VDD.n9507 2.2505
R28590 VDD.n9506 VDD.n9413 2.2505
R28591 VDD.n9505 VDD.n9504 2.2505
R28592 VDD.n9503 VDD.n9414 2.2505
R28593 VDD.n9502 VDD.n9501 2.2505
R28594 VDD.n9500 VDD.n9415 2.2505
R28595 VDD.n9499 VDD.n9498 2.2505
R28596 VDD.n9497 VDD.n9416 2.2505
R28597 VDD.n9496 VDD.n9495 2.2505
R28598 VDD.n9494 VDD.n9417 2.2505
R28599 VDD.n9493 VDD.n9492 2.2505
R28600 VDD.n9491 VDD.n9418 2.2505
R28601 VDD.n9490 VDD.n9489 2.2505
R28602 VDD.n9488 VDD.n9419 2.2505
R28603 VDD.n9487 VDD.n9486 2.2505
R28604 VDD.n9485 VDD.n9420 2.2505
R28605 VDD.n9484 VDD.n9483 2.2505
R28606 VDD.n9482 VDD.n9421 2.2505
R28607 VDD.n9481 VDD.n9480 2.2505
R28608 VDD.n9479 VDD.n9422 2.2505
R28609 VDD.n9478 VDD.n9477 2.2505
R28610 VDD.n9476 VDD.n9423 2.2505
R28611 VDD.n9475 VDD.n9474 2.2505
R28612 VDD.n9473 VDD.n9424 2.2505
R28613 VDD.n9472 VDD.n9471 2.2505
R28614 VDD.n9470 VDD.n9425 2.2505
R28615 VDD.n9469 VDD.n9468 2.2505
R28616 VDD.n9467 VDD.n9426 2.2505
R28617 VDD.n9466 VDD.n9465 2.2505
R28618 VDD.n9464 VDD.n9427 2.2505
R28619 VDD.n9463 VDD.n9462 2.2505
R28620 VDD.n9461 VDD.n9428 2.2505
R28621 VDD.n9460 VDD.n9459 2.2505
R28622 VDD.n9458 VDD.n9429 2.2505
R28623 VDD.n9457 VDD.n9456 2.2505
R28624 VDD.n9455 VDD.n9430 2.2505
R28625 VDD.n9454 VDD.n9453 2.2505
R28626 VDD.n9452 VDD.n9431 2.2505
R28627 VDD.n9451 VDD.n9450 2.2505
R28628 VDD.n9449 VDD.n9432 2.2505
R28629 VDD.n9448 VDD.n9447 2.2505
R28630 VDD.n9446 VDD.n9433 2.2505
R28631 VDD.n9445 VDD.n9444 2.2505
R28632 VDD.n9443 VDD.n9434 2.2505
R28633 VDD.n9442 VDD.n9441 2.2505
R28634 VDD.n9440 VDD.n9435 2.2505
R28635 VDD.n9439 VDD.n9438 2.2505
R28636 VDD.n9437 VDD.n9436 2.2505
R28637 VDD.n12441 VDD.n12440 2.2505
R28638 VDD.n12439 VDD.n196 2.2505
R28639 VDD.n12438 VDD.n12437 2.2505
R28640 VDD.n12436 VDD.n197 2.2505
R28641 VDD.n12435 VDD.n12434 2.2505
R28642 VDD.n12433 VDD.n198 2.2505
R28643 VDD.n12432 VDD.n12431 2.2505
R28644 VDD.n12430 VDD.n199 2.2505
R28645 VDD.n12429 VDD.n12428 2.2505
R28646 VDD.n12427 VDD.n200 2.2505
R28647 VDD.n12426 VDD.n12425 2.2505
R28648 VDD.n12424 VDD.n201 2.2505
R28649 VDD.n12423 VDD.n12422 2.2505
R28650 VDD.n12421 VDD.n202 2.2505
R28651 VDD.n12420 VDD.n12419 2.2505
R28652 VDD.n12418 VDD.n203 2.2505
R28653 VDD.n12417 VDD.n12416 2.2505
R28654 VDD.n12415 VDD.n204 2.2505
R28655 VDD.n12414 VDD.n12413 2.2505
R28656 VDD.n12412 VDD.n205 2.2505
R28657 VDD.n12411 VDD.n12410 2.2505
R28658 VDD.n12409 VDD.n206 2.2505
R28659 VDD.n12408 VDD.n12407 2.2505
R28660 VDD.n12406 VDD.n207 2.2505
R28661 VDD.n12405 VDD.n12404 2.2505
R28662 VDD.n12403 VDD.n208 2.2505
R28663 VDD.n12402 VDD.n12401 2.2505
R28664 VDD.n12400 VDD.n209 2.2505
R28665 VDD.n12399 VDD.n12398 2.2505
R28666 VDD.n12397 VDD.n210 2.2505
R28667 VDD.n12396 VDD.n12395 2.2505
R28668 VDD.n12394 VDD.n211 2.2505
R28669 VDD.n12393 VDD.n12392 2.2505
R28670 VDD.n12391 VDD.n212 2.2505
R28671 VDD.n12390 VDD.n12389 2.2505
R28672 VDD.n12388 VDD.n213 2.2505
R28673 VDD.n12387 VDD.n12386 2.2505
R28674 VDD.n12385 VDD.n214 2.2505
R28675 VDD.n12384 VDD.n12383 2.2505
R28676 VDD.n12382 VDD.n215 2.2505
R28677 VDD.n12381 VDD.n12380 2.2505
R28678 VDD.n12379 VDD.n216 2.2505
R28679 VDD.n12378 VDD.n12377 2.2505
R28680 VDD.n12376 VDD.n217 2.2505
R28681 VDD.n12375 VDD.n12374 2.2505
R28682 VDD.n12373 VDD.n218 2.2505
R28683 VDD.n12372 VDD.n12371 2.2505
R28684 VDD.n12370 VDD.n219 2.2505
R28685 VDD.n12369 VDD.n12368 2.2505
R28686 VDD.n12367 VDD.n220 2.2505
R28687 VDD.n12366 VDD.n12365 2.2505
R28688 VDD.n12364 VDD.n221 2.2505
R28689 VDD.n12363 VDD.n12362 2.2505
R28690 VDD.n12361 VDD.n222 2.2505
R28691 VDD.n12360 VDD.n12359 2.2505
R28692 VDD.n12358 VDD.n223 2.2505
R28693 VDD.n12357 VDD.n12356 2.2505
R28694 VDD.n12355 VDD.n224 2.2505
R28695 VDD.n12354 VDD.n12353 2.2505
R28696 VDD.n12352 VDD.n225 2.2505
R28697 VDD.n12351 VDD.n12350 2.2505
R28698 VDD.n12349 VDD.n226 2.2505
R28699 VDD.n12348 VDD.n12347 2.2505
R28700 VDD.n12346 VDD.n227 2.2505
R28701 VDD.n12345 VDD.n12344 2.2505
R28702 VDD.n12343 VDD.n228 2.2505
R28703 VDD.n12342 VDD.n12341 2.2505
R28704 VDD.n12340 VDD.n229 2.2505
R28705 VDD.n12339 VDD.n12338 2.2505
R28706 VDD.n12337 VDD.n230 2.2505
R28707 VDD.n12336 VDD.n12335 2.2505
R28708 VDD.n12334 VDD.n231 2.2505
R28709 VDD.n12333 VDD.n12332 2.2505
R28710 VDD.n12331 VDD.n232 2.2505
R28711 VDD.n12330 VDD.n12329 2.2505
R28712 VDD.n12328 VDD.n233 2.2505
R28713 VDD.n12327 VDD.n12326 2.2505
R28714 VDD.n12325 VDD.n234 2.2505
R28715 VDD.n12324 VDD.n12323 2.2505
R28716 VDD.n12322 VDD.n235 2.2505
R28717 VDD.n12321 VDD.n12320 2.2505
R28718 VDD.n12319 VDD.n236 2.2505
R28719 VDD.n12318 VDD.n12317 2.2505
R28720 VDD.n12316 VDD.n237 2.2505
R28721 VDD.n12315 VDD.n12314 2.2505
R28722 VDD.n12313 VDD.n238 2.2505
R28723 VDD.n12312 VDD.n12311 2.2505
R28724 VDD.n12310 VDD.n239 2.2505
R28725 VDD.n12309 VDD.n12308 2.2505
R28726 VDD.n12307 VDD.n240 2.2505
R28727 VDD.n12306 VDD.n12305 2.2505
R28728 VDD.n12304 VDD.n241 2.2505
R28729 VDD.n12303 VDD.n12302 2.2505
R28730 VDD.n12301 VDD.n242 2.2505
R28731 VDD.n12300 VDD.n12299 2.2505
R28732 VDD.n12298 VDD.n243 2.2505
R28733 VDD.n12297 VDD.n12296 2.2505
R28734 VDD.n12295 VDD.n244 2.2505
R28735 VDD.n12294 VDD.n12293 2.2505
R28736 VDD.n12292 VDD.n245 2.2505
R28737 VDD.n12291 VDD.n12290 2.2505
R28738 VDD.n12289 VDD.n246 2.2505
R28739 VDD.n12288 VDD.n12287 2.2505
R28740 VDD.n12286 VDD.n247 2.2505
R28741 VDD.n12285 VDD.n12284 2.2505
R28742 VDD.n12283 VDD.n248 2.2505
R28743 VDD.n12282 VDD.n12281 2.2505
R28744 VDD.n12280 VDD.n249 2.2505
R28745 VDD.n12279 VDD.n12278 2.2505
R28746 VDD.n12277 VDD.n250 2.2505
R28747 VDD.n12276 VDD.n12275 2.2505
R28748 VDD.n12274 VDD.n251 2.2505
R28749 VDD.n12273 VDD.n12272 2.2505
R28750 VDD.n12271 VDD.n252 2.2505
R28751 VDD.n12270 VDD.n12269 2.2505
R28752 VDD.n12268 VDD.n253 2.2505
R28753 VDD.n12267 VDD.n12266 2.2505
R28754 VDD.n12265 VDD.n254 2.2505
R28755 VDD.n12264 VDD.n12263 2.2505
R28756 VDD.n12262 VDD.n255 2.2505
R28757 VDD.n12261 VDD.n12260 2.2505
R28758 VDD.n12259 VDD.n256 2.2505
R28759 VDD.n12258 VDD.n12257 2.2505
R28760 VDD.n12256 VDD.n257 2.2505
R28761 VDD.n12255 VDD.n12254 2.2505
R28762 VDD.n12253 VDD.n258 2.2505
R28763 VDD.n12252 VDD.n12251 2.2505
R28764 VDD.n12250 VDD.n259 2.2505
R28765 VDD.n12249 VDD.n12248 2.2505
R28766 VDD.n12247 VDD.n260 2.2505
R28767 VDD.n12246 VDD.n12245 2.2505
R28768 VDD.n12244 VDD.n261 2.2505
R28769 VDD.n12243 VDD.n12242 2.2505
R28770 VDD.n12241 VDD.n262 2.2505
R28771 VDD.n12240 VDD.n12239 2.2505
R28772 VDD.n12238 VDD.n263 2.2505
R28773 VDD.n12237 VDD.n12236 2.2505
R28774 VDD.n12235 VDD.n264 2.2505
R28775 VDD.n12234 VDD.n12233 2.2505
R28776 VDD.n12232 VDD.n265 2.2505
R28777 VDD.n12231 VDD.n12230 2.2505
R28778 VDD.n12229 VDD.n266 2.2505
R28779 VDD.n12228 VDD.n12227 2.2505
R28780 VDD.n12226 VDD.n267 2.2505
R28781 VDD.n12225 VDD.n12224 2.2505
R28782 VDD.n12223 VDD.n268 2.2505
R28783 VDD.n12222 VDD.n12221 2.2505
R28784 VDD.n12220 VDD.n269 2.2505
R28785 VDD.n12219 VDD.n12218 2.2505
R28786 VDD.n12217 VDD.n270 2.2505
R28787 VDD.n12216 VDD.n12215 2.2505
R28788 VDD.n12214 VDD.n271 2.2505
R28789 VDD.n12213 VDD.n12212 2.2505
R28790 VDD.n12211 VDD.n272 2.2505
R28791 VDD.n12210 VDD.n12209 2.2505
R28792 VDD.n12208 VDD.n273 2.2505
R28793 VDD.n12207 VDD.n12206 2.2505
R28794 VDD.n12205 VDD.n274 2.2505
R28795 VDD.n12204 VDD.n12203 2.2505
R28796 VDD.n12202 VDD.n275 2.2505
R28797 VDD.n12201 VDD.n12200 2.2505
R28798 VDD.n12199 VDD.n276 2.2505
R28799 VDD.n12198 VDD.n12197 2.2505
R28800 VDD.n12196 VDD.n277 2.2505
R28801 VDD.n12195 VDD.n12194 2.2505
R28802 VDD.n12193 VDD.n278 2.2505
R28803 VDD.n12192 VDD.n12191 2.2505
R28804 VDD.n12190 VDD.n279 2.2505
R28805 VDD.n12189 VDD.n12188 2.2505
R28806 VDD.n12187 VDD.n280 2.2505
R28807 VDD.n12186 VDD.n12185 2.2505
R28808 VDD.n12184 VDD.n281 2.2505
R28809 VDD.n12183 VDD.n12182 2.2505
R28810 VDD.n12181 VDD.n282 2.2505
R28811 VDD.n12180 VDD.n12179 2.2505
R28812 VDD.n12178 VDD.n283 2.2505
R28813 VDD.n12177 VDD.n12176 2.2505
R28814 VDD.n12175 VDD.n284 2.2505
R28815 VDD.n12174 VDD.n12173 2.2505
R28816 VDD.n12172 VDD.n285 2.2505
R28817 VDD.n12171 VDD.n12170 2.2505
R28818 VDD.n12169 VDD.n286 2.2505
R28819 VDD.n12168 VDD.n12167 2.2505
R28820 VDD.n12166 VDD.n287 2.2505
R28821 VDD.n12165 VDD.n12164 2.2505
R28822 VDD.n12163 VDD.n288 2.2505
R28823 VDD.n12162 VDD.n12161 2.2505
R28824 VDD.n12160 VDD.n289 2.2505
R28825 VDD.n12159 VDD.n12158 2.2505
R28826 VDD.n12157 VDD.n290 2.2505
R28827 VDD.n12156 VDD.n12155 2.2505
R28828 VDD.n12154 VDD.n291 2.2505
R28829 VDD.n12153 VDD.n12152 2.2505
R28830 VDD.n12151 VDD.n292 2.2505
R28831 VDD.n12150 VDD.n12149 2.2505
R28832 VDD.n12148 VDD.n293 2.2505
R28833 VDD.n12147 VDD.n12146 2.2505
R28834 VDD.n12145 VDD.n294 2.2505
R28835 VDD.n12144 VDD.n12143 2.2505
R28836 VDD.n12142 VDD.n295 2.2505
R28837 VDD.n12141 VDD.n12140 2.2505
R28838 VDD.n12139 VDD.n296 2.2505
R28839 VDD.n12138 VDD.n12137 2.2505
R28840 VDD.n12136 VDD.n297 2.2505
R28841 VDD.n12135 VDD.n12134 2.2505
R28842 VDD.n12133 VDD.n298 2.2505
R28843 VDD.n12132 VDD.n12131 2.2505
R28844 VDD.n12130 VDD.n299 2.2505
R28845 VDD.n12129 VDD.n12128 2.2505
R28846 VDD.n12127 VDD.n300 2.2505
R28847 VDD.n12126 VDD.n12125 2.2505
R28848 VDD.n12124 VDD.n301 2.2505
R28849 VDD.n12123 VDD.n12122 2.2505
R28850 VDD.n12121 VDD.n302 2.2505
R28851 VDD.n12120 VDD.n12119 2.2505
R28852 VDD.n12118 VDD.n303 2.2505
R28853 VDD.n12117 VDD.n12116 2.2505
R28854 VDD.n12115 VDD.n304 2.2505
R28855 VDD.n12114 VDD.n12113 2.2505
R28856 VDD.n12112 VDD.n305 2.2505
R28857 VDD.n12111 VDD.n12110 2.2505
R28858 VDD.n12109 VDD.n306 2.2505
R28859 VDD.n12108 VDD.n12107 2.2505
R28860 VDD.n12106 VDD.n307 2.2505
R28861 VDD.n12105 VDD.n12104 2.2505
R28862 VDD.n12103 VDD.n308 2.2505
R28863 VDD.n12102 VDD.n12101 2.2505
R28864 VDD.n12100 VDD.n309 2.2505
R28865 VDD.n12099 VDD.n12098 2.2505
R28866 VDD.n12097 VDD.n310 2.2505
R28867 VDD.n12096 VDD.n12095 2.2505
R28868 VDD.n12094 VDD.n311 2.2505
R28869 VDD.n12093 VDD.n12092 2.2505
R28870 VDD.n12091 VDD.n312 2.2505
R28871 VDD.n12090 VDD.n12089 2.2505
R28872 VDD.n12088 VDD.n313 2.2505
R28873 VDD.n12087 VDD.n12086 2.2505
R28874 VDD.n12085 VDD.n314 2.2505
R28875 VDD.n12084 VDD.n12083 2.2505
R28876 VDD.n12082 VDD.n315 2.2505
R28877 VDD.n12081 VDD.n12080 2.2505
R28878 VDD.n12079 VDD.n316 2.2505
R28879 VDD.n12078 VDD.n12077 2.2505
R28880 VDD.n12076 VDD.n317 2.2505
R28881 VDD.n12075 VDD.n12074 2.2505
R28882 VDD.n12073 VDD.n318 2.2505
R28883 VDD.n12072 VDD.n12071 2.2505
R28884 VDD.n12070 VDD.n319 2.2505
R28885 VDD.n12069 VDD.n12068 2.2505
R28886 VDD.n12067 VDD.n320 2.2505
R28887 VDD.n12066 VDD.n12065 2.2505
R28888 VDD.n12064 VDD.n321 2.2505
R28889 VDD.n12063 VDD.n12062 2.2505
R28890 VDD.n12061 VDD.n322 2.2505
R28891 VDD.n12060 VDD.n12059 2.2505
R28892 VDD.n12058 VDD.n323 2.2505
R28893 VDD.n12057 VDD.n12056 2.2505
R28894 VDD.n12055 VDD.n324 2.2505
R28895 VDD.n12054 VDD.n12053 2.2505
R28896 VDD.n12052 VDD.n325 2.2505
R28897 VDD.n12051 VDD.n12050 2.2505
R28898 VDD.n12049 VDD.n326 2.2505
R28899 VDD.n12048 VDD.n12047 2.2505
R28900 VDD.n12046 VDD.n327 2.2505
R28901 VDD.n12045 VDD.n12044 2.2505
R28902 VDD.n12043 VDD.n328 2.2505
R28903 VDD.n12042 VDD.n12041 2.2505
R28904 VDD.n12040 VDD.n329 2.2505
R28905 VDD.n12039 VDD.n12038 2.2505
R28906 VDD.n12037 VDD.n330 2.2505
R28907 VDD.n12036 VDD.n12035 2.2505
R28908 VDD.n12034 VDD.n331 2.2505
R28909 VDD.n12033 VDD.n12032 2.2505
R28910 VDD.n12031 VDD.n332 2.2505
R28911 VDD.n12030 VDD.n12029 2.2505
R28912 VDD.n12028 VDD.n333 2.2505
R28913 VDD.n12027 VDD.n12026 2.2505
R28914 VDD.n12025 VDD.n334 2.2505
R28915 VDD.n12024 VDD.n12023 2.2505
R28916 VDD.n12022 VDD.n335 2.2505
R28917 VDD.n12021 VDD.n12020 2.2505
R28918 VDD.n12019 VDD.n336 2.2505
R28919 VDD.n12018 VDD.n12017 2.2505
R28920 VDD.n12016 VDD.n337 2.2505
R28921 VDD.n12015 VDD.n12014 2.2505
R28922 VDD.n12013 VDD.n338 2.2505
R28923 VDD.n12012 VDD.n12011 2.2505
R28924 VDD.n12010 VDD.n339 2.2505
R28925 VDD.n12009 VDD.n12008 2.2505
R28926 VDD.n12007 VDD.n340 2.2505
R28927 VDD.n12006 VDD.n12005 2.2505
R28928 VDD.n12004 VDD.n341 2.2505
R28929 VDD.n12003 VDD.n12002 2.2505
R28930 VDD.n12001 VDD.n342 2.2505
R28931 VDD.n12000 VDD.n11999 2.2505
R28932 VDD.n11998 VDD.n343 2.2505
R28933 VDD.n11997 VDD.n11996 2.2505
R28934 VDD.n11995 VDD.n344 2.2505
R28935 VDD.n11994 VDD.n11993 2.2505
R28936 VDD.n11992 VDD.n345 2.2505
R28937 VDD.n11991 VDD.n11990 2.2505
R28938 VDD.n11989 VDD.n346 2.2505
R28939 VDD.n11988 VDD.n11987 2.2505
R28940 VDD.n11986 VDD.n347 2.2505
R28941 VDD.n11985 VDD.n11984 2.2505
R28942 VDD.n11983 VDD.n348 2.2505
R28943 VDD.n11982 VDD.n11981 2.2505
R28944 VDD.n11980 VDD.n349 2.2505
R28945 VDD.n11979 VDD.n11978 2.2505
R28946 VDD.n11977 VDD.n350 2.2505
R28947 VDD.n11976 VDD.n11975 2.2505
R28948 VDD.n11974 VDD.n351 2.2505
R28949 VDD.n11973 VDD.n11972 2.2505
R28950 VDD.n11971 VDD.n352 2.2505
R28951 VDD.n11970 VDD.n11969 2.2505
R28952 VDD.n11968 VDD.n353 2.2505
R28953 VDD.n11967 VDD.n11966 2.2505
R28954 VDD.n11965 VDD.n354 2.2505
R28955 VDD.n11964 VDD.n11963 2.2505
R28956 VDD.n11962 VDD.n355 2.2505
R28957 VDD.n11961 VDD.n11960 2.2505
R28958 VDD.n11959 VDD.n356 2.2505
R28959 VDD.n11958 VDD.n11957 2.2505
R28960 VDD.n11956 VDD.n357 2.2505
R28961 VDD.n11955 VDD.n11954 2.2505
R28962 VDD.n11953 VDD.n358 2.2505
R28963 VDD.n11952 VDD.n11951 2.2505
R28964 VDD.n11950 VDD.n359 2.2505
R28965 VDD.n11949 VDD.n11948 2.2505
R28966 VDD.n11947 VDD.n360 2.2505
R28967 VDD.n11946 VDD.n11945 2.2505
R28968 VDD.n11944 VDD.n361 2.2505
R28969 VDD.n11943 VDD.n11942 2.2505
R28970 VDD.n11941 VDD.n362 2.2505
R28971 VDD.n11940 VDD.n11939 2.2505
R28972 VDD.n11938 VDD.n363 2.2505
R28973 VDD.n11937 VDD.n11936 2.2505
R28974 VDD.n11935 VDD.n364 2.2505
R28975 VDD.n11934 VDD.n11933 2.2505
R28976 VDD.n11932 VDD.n365 2.2505
R28977 VDD.n11931 VDD.n11930 2.2505
R28978 VDD.n11929 VDD.n366 2.2505
R28979 VDD.n11928 VDD.n11927 2.2505
R28980 VDD.n11926 VDD.n367 2.2505
R28981 VDD.n11925 VDD.n11924 2.2505
R28982 VDD.n11923 VDD.n368 2.2505
R28983 VDD.n11922 VDD.n11921 2.2505
R28984 VDD.n11920 VDD.n369 2.2505
R28985 VDD.n11919 VDD.n11918 2.2505
R28986 VDD.n11917 VDD.n370 2.2505
R28987 VDD.n11916 VDD.n11915 2.2505
R28988 VDD.n11914 VDD.n371 2.2505
R28989 VDD.n11913 VDD.n11912 2.2505
R28990 VDD.n11911 VDD.n372 2.2505
R28991 VDD.n11910 VDD.n11909 2.2505
R28992 VDD.n11908 VDD.n373 2.2505
R28993 VDD.n11907 VDD.n11906 2.2505
R28994 VDD.n11905 VDD.n374 2.2505
R28995 VDD.n11904 VDD.n11903 2.2505
R28996 VDD.n11902 VDD.n375 2.2505
R28997 VDD.n11901 VDD.n11900 2.2505
R28998 VDD.n11899 VDD.n376 2.2505
R28999 VDD.n11898 VDD.n11897 2.2505
R29000 VDD.n11896 VDD.n377 2.2505
R29001 VDD.n11895 VDD.n11894 2.2505
R29002 VDD.n11893 VDD.n378 2.2505
R29003 VDD.n11892 VDD.n11891 2.2505
R29004 VDD.n11890 VDD.n379 2.2505
R29005 VDD.n11889 VDD.n11888 2.2505
R29006 VDD.n11887 VDD.n380 2.2505
R29007 VDD.n11886 VDD.n11885 2.2505
R29008 VDD.n11884 VDD.n381 2.2505
R29009 VDD.n11883 VDD.n11882 2.2505
R29010 VDD.n11881 VDD.n382 2.2505
R29011 VDD.n11880 VDD.n11879 2.2505
R29012 VDD.n11878 VDD.n383 2.2505
R29013 VDD.n11877 VDD.n11876 2.2505
R29014 VDD.n11875 VDD.n384 2.2505
R29015 VDD.n11874 VDD.n11873 2.2505
R29016 VDD.n11871 VDD.n385 2.2505
R29017 VDD.n11870 VDD.n11869 2.2505
R29018 VDD.n11868 VDD.n386 2.2505
R29019 VDD.n11867 VDD.n11866 2.2505
R29020 VDD.n11865 VDD.n387 2.2505
R29021 VDD.n11864 VDD.n11863 2.2505
R29022 VDD.n11862 VDD.n388 2.2505
R29023 VDD.n11861 VDD.n11860 2.2505
R29024 VDD.n11859 VDD.n389 2.2505
R29025 VDD.n11858 VDD.n11857 2.2505
R29026 VDD.n11856 VDD.n390 2.2505
R29027 VDD.n11855 VDD.n11854 2.2505
R29028 VDD.n11853 VDD.n391 2.2505
R29029 VDD.n11852 VDD.n11851 2.2505
R29030 VDD.n11850 VDD.n392 2.2505
R29031 VDD.n11849 VDD.n11848 2.2505
R29032 VDD.n11847 VDD.n393 2.2505
R29033 VDD.n11846 VDD.n11845 2.2505
R29034 VDD.n11844 VDD.n394 2.2505
R29035 VDD.n11843 VDD.n11842 2.2505
R29036 VDD.n11841 VDD.n395 2.2505
R29037 VDD.n11840 VDD.n11839 2.2505
R29038 VDD.n11838 VDD.n396 2.2505
R29039 VDD.n11837 VDD.n11836 2.2505
R29040 VDD.n11835 VDD.n397 2.2505
R29041 VDD.n11834 VDD.n11833 2.2505
R29042 VDD.n11832 VDD.n398 2.2505
R29043 VDD.n11831 VDD.n11830 2.2505
R29044 VDD.n11829 VDD.n399 2.2505
R29045 VDD.n11828 VDD.n11827 2.2505
R29046 VDD.n11826 VDD.n400 2.2505
R29047 VDD.n11825 VDD.n11824 2.2505
R29048 VDD.n11823 VDD.n401 2.2505
R29049 VDD.n11822 VDD.n11821 2.2505
R29050 VDD.n11820 VDD.n402 2.2505
R29051 VDD.n11819 VDD.n11818 2.2505
R29052 VDD.n11817 VDD.n403 2.2505
R29053 VDD.n11816 VDD.n11815 2.2505
R29054 VDD.n11814 VDD.n404 2.2505
R29055 VDD.n11813 VDD.n11812 2.2505
R29056 VDD.n1449 VDD.n1448 2.2505
R29057 VDD.n1754 VDD.n681 2.25019
R29058 VDD.n998 VDD.n957 2.25019
R29059 VDD.n12638 VDD.n2 2.25019
R29060 VDD.n4595 VDD.n2411 2.25018
R29061 VDD.n2118 VDD.n2108 2.25015
R29062 VDD.n5537 VDD.n5490 2.25014
R29063 VDD.n5910 VDD.n5541 2.25014
R29064 VDD.n5889 VDD.n5888 2.25014
R29065 VDD.n6319 VDD.n5913 2.24874
R29066 VDD.n6321 VDD.n6320 2.24218
R29067 VDD.n6323 VDD.n5982 2.24218
R29068 VDD.n6320 VDD.n5915 2.24218
R29069 VDD.n6173 VDD.n6172 2.24218
R29070 VDD.n6177 VDD.n6176 2.24218
R29071 VDD.n6173 VDD.n6017 2.24218
R29072 VDD.n10817 VDD.n10816 2.24218
R29073 VDD.n10818 VDD.n10817 2.24218
R29074 VDD.n8093 VDD.n8092 2.24218
R29075 VDD.n8095 VDD.n2107 2.24218
R29076 VDD.n2117 VDD.n2105 2.24218
R29077 VDD.n2004 VDD.n2003 2.24218
R29078 VDD.n5907 VDD.n5906 2.24218
R29079 VDD.n5534 VDD.n5530 2.24218
R29080 VDD.n5532 VDD.n5529 2.24218
R29081 VDD.n5887 VDD.n1919 2.24218
R29082 VDD.n5882 VDD.n1918 2.24218
R29083 VDD.n5909 VDD.n5901 2.24218
R29084 VDD.n5903 VDD.n5901 2.24218
R29085 VDD.n5884 VDD.n1918 2.24218
R29086 VDD.n5536 VDD.n5503 2.24218
R29087 VDD.n11048 VDD.n671 2.24218
R29088 VDD.n11048 VDD.n670 2.24218
R29089 VDD.n11044 VDD.n672 2.24218
R29090 VDD.n11128 VDD.n11127 2.24218
R29091 VDD.n640 VDD.n639 2.24218
R29092 VDD.n11127 VDD.n643 2.24218
R29093 VDD.n12583 VDD.n12578 2.24218
R29094 VDD.n12585 VDD.n12560 2.24218
R29095 VDD.n12581 VDD.n12562 2.24218
R29096 VDD.n12626 VDD.n10 2.24218
R29097 VDD.n12627 VDD.n12626 2.24218
R29098 VDD.n12622 VDD.n9 2.24218
R29099 VDD.n1753 VDD.n680 2.24218
R29100 VDD.n1758 VDD.n1756 2.24218
R29101 VDD.n1002 VDD.n999 2.24218
R29102 VDD.n1004 VDD.n955 2.24218
R29103 VDD.n4 VDD.n1 2.24218
R29104 VDD.n12637 VDD.n1 2.24218
R29105 VDD.n2424 VDD.n2409 2.24111
R29106 VDD.n5220 VDD.n2423 2.24111
R29107 VDD.n5220 VDD.n2422 2.24111
R29108 VDD.n5220 VDD.n2421 2.24111
R29109 VDD.n5220 VDD.n2420 2.24111
R29110 VDD.n5220 VDD.n2419 2.24111
R29111 VDD.n5220 VDD.n2418 2.24111
R29112 VDD.n5220 VDD.n2417 2.24111
R29113 VDD.n5220 VDD.n2416 2.24111
R29114 VDD.n5220 VDD.n2415 2.24111
R29115 VDD.n5220 VDD.n2414 2.24111
R29116 VDD.n5220 VDD.n2413 2.24111
R29117 VDD.n5220 VDD.n2412 2.24111
R29118 VDD.n4596 VDD.n2408 2.24111
R29119 VDD.n5218 VDD.n5217 2.24111
R29120 VDD.n5218 VDD.n5216 2.24111
R29121 VDD.n5218 VDD.n5215 2.24111
R29122 VDD.n5218 VDD.n5214 2.24111
R29123 VDD.n5218 VDD.n5213 2.24111
R29124 VDD.n5218 VDD.n5212 2.24111
R29125 VDD.n5218 VDD.n5211 2.24111
R29126 VDD.n5218 VDD.n5210 2.24111
R29127 VDD.n5218 VDD.n5209 2.24111
R29128 VDD.n5218 VDD.n5208 2.24111
R29129 VDD.n5218 VDD.n5207 2.24111
R29130 VDD.n5218 VDD.n5206 2.24111
R29131 VDD.n5218 VDD.n5205 2.24111
R29132 VDD.n5203 VDD.n5202 2.24111
R29133 VDD.n5202 VDD.n4597 2.24111
R29134 VDD.n9199 VDD.n9185 2.24111
R29135 VDD.n9198 VDD.n9184 2.24111
R29136 VDD.n9187 VDD.n9185 2.24111
R29137 VDD.n9188 VDD.n9184 2.24111
R29138 VDD.n9189 VDD.n9185 2.24111
R29139 VDD.n9190 VDD.n9184 2.24111
R29140 VDD.n9191 VDD.n9185 2.24111
R29141 VDD.n9192 VDD.n9184 2.24111
R29142 VDD.n9193 VDD.n9185 2.24111
R29143 VDD.n9194 VDD.n9184 2.24111
R29144 VDD.n9195 VDD.n9185 2.24111
R29145 VDD.n9196 VDD.n9184 2.24111
R29146 VDD.n9197 VDD.n9185 2.24111
R29147 VDD.n12448 VDD.n193 2.24111
R29148 VDD.n12448 VDD.n192 2.24111
R29149 VDD.n12448 VDD.n191 2.24111
R29150 VDD.n12445 VDD.n12444 2.24111
R29151 VDD.n12445 VDD.n12443 2.24111
R29152 VDD.n12445 VDD.n12442 2.24111
R29153 VDD.n12446 VDD.n12445 2.24111
R29154 VDD.n6116 VDD.n6115 2.24038
R29155 VDD.n6073 VDD.n6072 2.24038
R29156 VDD.n6800 VDD.n6739 2.24038
R29157 VDD.n6746 VDD.n6745 2.24038
R29158 VDD.n7885 VDD.n7884 2.21344
R29159 VDD.n7881 VDD.n7880 2.21344
R29160 VDD.n7877 VDD.n7876 2.21344
R29161 VDD.n7871 VDD.n7870 2.21344
R29162 VDD.n7867 VDD.n7866 2.21344
R29163 VDD.n6136 VDD.n6135 2.2016
R29164 VDD.n6139 VDD.n6138 2.2016
R29165 VDD.n6143 VDD.n6142 2.2016
R29166 VDD.n6147 VDD.n6146 2.2016
R29167 VDD.n6132 VDD.n6131 2.2016
R29168 VDD.n6128 VDD.n6127 2.2016
R29169 VDD.n6124 VDD.n6123 2.2016
R29170 VDD.n6120 VDD.n6119 2.2016
R29171 VDD.n6044 VDD.n6043 2.2016
R29172 VDD.n6047 VDD.n6046 2.2016
R29173 VDD.n6051 VDD.n6050 2.2016
R29174 VDD.n6055 VDD.n6054 2.2016
R29175 VDD.n6078 VDD.n6077 2.2016
R29176 VDD.n6082 VDD.n6081 2.2016
R29177 VDD.n6086 VDD.n6085 2.2016
R29178 VDD.n6090 VDD.n6089 2.2016
R29179 VDD.n6810 VDD.n6809 2.2016
R29180 VDD.n6813 VDD.n6812 2.2016
R29181 VDD.n6817 VDD.n6816 2.2016
R29182 VDD.n6821 VDD.n6820 2.2016
R29183 VDD.n6826 VDD.n6825 2.2016
R29184 VDD.n6830 VDD.n6829 2.2016
R29185 VDD.n6834 VDD.n6833 2.2016
R29186 VDD.n6838 VDD.n6837 2.2016
R29187 VDD.n6777 VDD.n6776 2.2016
R29188 VDD.n6780 VDD.n6779 2.2016
R29189 VDD.n6784 VDD.n6783 2.2016
R29190 VDD.n6788 VDD.n6787 2.2016
R29191 VDD.n6773 VDD.n6772 2.2016
R29192 VDD.n6769 VDD.n6768 2.2016
R29193 VDD.n6765 VDD.n6764 2.2016
R29194 VDD.n6761 VDD.n6760 2.2016
R29195 VDD.n6951 VDD.n6950 2.18645
R29196 VDD.n6504 VDD.n6447 2.18645
R29197 VDD.n6996 VDD.n6995 2.18502
R29198 VDD.n6991 VDD.n6990 2.18502
R29199 VDD.n6986 VDD.n6985 2.18502
R29200 VDD.n6981 VDD.n6980 2.18502
R29201 VDD.n6899 VDD.n6898 2.18502
R29202 VDD.n6894 VDD.n6893 2.18502
R29203 VDD.n6889 VDD.n6888 2.18502
R29204 VDD.n6948 VDD.n6947 2.18502
R29205 VDD.n6943 VDD.n6942 2.18502
R29206 VDD.n6938 VDD.n6937 2.18502
R29207 VDD.n6933 VDD.n6932 2.18502
R29208 VDD.n6918 VDD.n6917 2.18502
R29209 VDD.n6913 VDD.n6912 2.18502
R29210 VDD.n6908 VDD.n6907 2.18502
R29211 VDD.n6446 VDD.n6445 2.18502
R29212 VDD.n6443 VDD.n6442 2.18502
R29213 VDD.n6440 VDD.n6439 2.18502
R29214 VDD.n6437 VDD.n6436 2.18502
R29215 VDD.n6432 VDD.n6431 2.18502
R29216 VDD.n6427 VDD.n6426 2.18502
R29217 VDD.n6422 VDD.n6421 2.18502
R29218 VDD.n6483 VDD.n6482 2.18502
R29219 VDD.n6480 VDD.n6479 2.18502
R29220 VDD.n6477 VDD.n6476 2.18502
R29221 VDD.n6474 VDD.n6473 2.18502
R29222 VDD.n6469 VDD.n6468 2.18502
R29223 VDD.n6464 VDD.n6463 2.18502
R29224 VDD.n6459 VDD.n6458 2.18502
R29225 VDD.n8044 VDD.n8043 2.1566
R29226 VDD.n8039 VDD.n8038 2.1566
R29227 VDD.n8034 VDD.n8033 2.1566
R29228 VDD.n8025 VDD.n8024 2.1566
R29229 VDD.n8020 VDD.n8019 2.1566
R29230 VDD.n7939 VDD.n7938 2.14594
R29231 VDD.n7934 VDD.n7933 2.14594
R29232 VDD.n7929 VDD.n7928 2.14594
R29233 VDD.n7920 VDD.n7919 2.14594
R29234 VDD.n7915 VDD.n7914 2.14594
R29235 VDD.n6959 VDD.n6921 2.0852
R29236 VDD.n6496 VDD.n6495 2.0852
R29237 VDD.n6074 VDD.n6073 2.0852
R29238 VDD.n6791 VDD.n6746 2.0852
R29239 VDD.n1761 VDD.n6 1.9774
R29240 VDD.n12634 VDD.n6 1.9617
R29241 VDD.n12634 VDD.n12633 1.84997
R29242 VDD.n1762 VDD.n1761 1.83884
R29243 VDD.n8089 VDD.n8087 1.78866
R29244 VDD.n7015 VDD.n7013 1.73609
R29245 VDD.n6968 VDD.n6878 1.73609
R29246 VDD.n6560 VDD.n6559 1.73609
R29247 VDD.n6521 VDD.n6520 1.73609
R29248 VDD.n2058 VDD.n2057 1.73383
R29249 VDD.n10770 VDD.n10769 1.73383
R29250 VDD.n5260 VDD.n5223 1.73383
R29251 VDD.n5258 VDD.n5224 1.73383
R29252 VDD.n5255 VDD.n5226 1.73383
R29253 VDD.n5250 VDD.n5228 1.73383
R29254 VDD.n5247 VDD.n5229 1.73383
R29255 VDD.n5242 VDD.n5232 1.73383
R29256 VDD.n5240 VDD.n5233 1.73383
R29257 VDD.n5237 VDD.n5235 1.73383
R29258 VDD.n5261 VDD.n5260 1.73383
R29259 VDD.n5258 VDD.n5257 1.73383
R29260 VDD.n5256 VDD.n5255 1.73383
R29261 VDD.n5251 VDD.n5250 1.73383
R29262 VDD.n5247 VDD.n5246 1.73383
R29263 VDD.n5243 VDD.n5242 1.73383
R29264 VDD.n5240 VDD.n5239 1.73383
R29265 VDD.n5238 VDD.n5237 1.73383
R29266 VDD.n5470 VDD.n5380 1.73383
R29267 VDD.n5468 VDD.n5381 1.73383
R29268 VDD.n5465 VDD.n5383 1.73383
R29269 VDD.n5460 VDD.n5385 1.73383
R29270 VDD.n5457 VDD.n5386 1.73383
R29271 VDD.n5452 VDD.n5389 1.73383
R29272 VDD.n5450 VDD.n5390 1.73383
R29273 VDD.n5447 VDD.n5392 1.73383
R29274 VDD.n5471 VDD.n5470 1.73383
R29275 VDD.n5468 VDD.n5467 1.73383
R29276 VDD.n5466 VDD.n5465 1.73383
R29277 VDD.n5461 VDD.n5460 1.73383
R29278 VDD.n5457 VDD.n5456 1.73383
R29279 VDD.n5453 VDD.n5452 1.73383
R29280 VDD.n5450 VDD.n5449 1.73383
R29281 VDD.n5448 VDD.n5447 1.73383
R29282 VDD.n5935 VDD.n5934 1.73383
R29283 VDD.n5932 VDD.n5931 1.73383
R29284 VDD.n5930 VDD.n5929 1.73383
R29285 VDD.n5925 VDD.n5274 1.73383
R29286 VDD.n6582 VDD.n6581 1.73383
R29287 VDD.n6587 VDD.n6586 1.73383
R29288 VDD.n6589 VDD.n6588 1.73383
R29289 VDD.n6592 VDD.n6591 1.73383
R29290 VDD.n5977 VDD.n5976 1.73383
R29291 VDD.n5974 VDD.n5973 1.73383
R29292 VDD.n5972 VDD.n5971 1.73383
R29293 VDD.n5967 VDD.n5966 1.73383
R29294 VDD.n5963 VDD.n5962 1.73383
R29295 VDD.n5959 VDD.n5958 1.73383
R29296 VDD.n5956 VDD.n5955 1.73383
R29297 VDD.n5954 VDD.n5953 1.73383
R29298 VDD.n5359 VDD.n5322 1.73383
R29299 VDD.n5357 VDD.n5323 1.73383
R29300 VDD.n5354 VDD.n5325 1.73383
R29301 VDD.n5349 VDD.n5327 1.73383
R29302 VDD.n5346 VDD.n5328 1.73383
R29303 VDD.n5341 VDD.n5331 1.73383
R29304 VDD.n5339 VDD.n5332 1.73383
R29305 VDD.n5336 VDD.n5334 1.73383
R29306 VDD.n5360 VDD.n5359 1.73383
R29307 VDD.n5357 VDD.n5356 1.73383
R29308 VDD.n5355 VDD.n5354 1.73383
R29309 VDD.n5350 VDD.n5349 1.73383
R29310 VDD.n5346 VDD.n5345 1.73383
R29311 VDD.n5342 VDD.n5341 1.73383
R29312 VDD.n5339 VDD.n5338 1.73383
R29313 VDD.n5337 VDD.n5336 1.73383
R29314 VDD.n6036 VDD.n6035 1.73383
R29315 VDD.n6034 VDD.n6033 1.73383
R29316 VDD.n6031 VDD.n6030 1.73383
R29317 VDD.n6027 VDD.n5283 1.73383
R29318 VDD.n6573 VDD.n6572 1.73383
R29319 VDD.n6569 VDD.n6568 1.73383
R29320 VDD.n6566 VDD.n6565 1.73383
R29321 VDD.n6564 VDD.n6563 1.73383
R29322 VDD.n6170 VDD.n6169 1.73383
R29323 VDD.n6167 VDD.n6166 1.73383
R29324 VDD.n6165 VDD.n6164 1.73383
R29325 VDD.n6160 VDD.n5302 1.73383
R29326 VDD.n6401 VDD.n6400 1.73383
R29327 VDD.n6406 VDD.n6405 1.73383
R29328 VDD.n6408 VDD.n6407 1.73383
R29329 VDD.n6411 VDD.n6410 1.73383
R29330 VDD.n6005 VDD.n5990 1.73383
R29331 VDD.n6003 VDD.n5991 1.73383
R29332 VDD.n6000 VDD.n5993 1.73383
R29333 VDD.n5994 VDD.n5313 1.73383
R29334 VDD.n6392 VDD.n5314 1.73383
R29335 VDD.n6387 VDD.n5317 1.73383
R29336 VDD.n6385 VDD.n5318 1.73383
R29337 VDD.n6382 VDD.n5320 1.73383
R29338 VDD.n6006 VDD.n6005 1.73383
R29339 VDD.n6003 VDD.n6002 1.73383
R29340 VDD.n6001 VDD.n6000 1.73383
R29341 VDD.n5996 VDD.n5313 1.73383
R29342 VDD.n6392 VDD.n6391 1.73383
R29343 VDD.n6388 VDD.n6387 1.73383
R29344 VDD.n6385 VDD.n6384 1.73383
R29345 VDD.n6383 VDD.n6382 1.73383
R29346 VDD.n6294 VDD.n6202 1.73383
R29347 VDD.n6292 VDD.n6203 1.73383
R29348 VDD.n6289 VDD.n6205 1.73383
R29349 VDD.n6284 VDD.n6207 1.73383
R29350 VDD.n6281 VDD.n6208 1.73383
R29351 VDD.n6276 VDD.n6211 1.73383
R29352 VDD.n6274 VDD.n6212 1.73383
R29353 VDD.n6271 VDD.n6214 1.73383
R29354 VDD.n6258 VDD.n6221 1.73383
R29355 VDD.n6256 VDD.n6222 1.73383
R29356 VDD.n6253 VDD.n6224 1.73383
R29357 VDD.n6248 VDD.n6226 1.73383
R29358 VDD.n6245 VDD.n6227 1.73383
R29359 VDD.n6240 VDD.n6230 1.73383
R29360 VDD.n6238 VDD.n6231 1.73383
R29361 VDD.n6235 VDD.n6233 1.73383
R29362 VDD.n6295 VDD.n6294 1.73383
R29363 VDD.n6292 VDD.n6291 1.73383
R29364 VDD.n6290 VDD.n6289 1.73383
R29365 VDD.n6285 VDD.n6284 1.73383
R29366 VDD.n6281 VDD.n6280 1.73383
R29367 VDD.n6277 VDD.n6276 1.73383
R29368 VDD.n6274 VDD.n6273 1.73383
R29369 VDD.n6272 VDD.n6271 1.73383
R29370 VDD.n6259 VDD.n6258 1.73383
R29371 VDD.n6256 VDD.n6255 1.73383
R29372 VDD.n6254 VDD.n6253 1.73383
R29373 VDD.n6249 VDD.n6248 1.73383
R29374 VDD.n6245 VDD.n6244 1.73383
R29375 VDD.n6241 VDD.n6240 1.73383
R29376 VDD.n6238 VDD.n6237 1.73383
R29377 VDD.n6236 VDD.n6235 1.73383
R29378 VDD.n6333 VDD.n6332 1.73383
R29379 VDD.n6337 VDD.n6336 1.73383
R29380 VDD.n6339 VDD.n6338 1.73383
R29381 VDD.n6345 VDD.n6344 1.73383
R29382 VDD.n6347 VDD.n6346 1.73383
R29383 VDD.n6352 VDD.n6351 1.73383
R29384 VDD.n6356 VDD.n6355 1.73383
R29385 VDD.n6358 VDD.n6357 1.73383
R29386 VDD.n6334 VDD.n6333 1.73383
R29387 VDD.n6336 VDD.n6335 1.73383
R29388 VDD.n6340 VDD.n6339 1.73383
R29389 VDD.n6344 VDD.n6343 1.73383
R29390 VDD.n6348 VDD.n6347 1.73383
R29391 VDD.n6353 VDD.n6352 1.73383
R29392 VDD.n6355 VDD.n6354 1.73383
R29393 VDD.n6359 VDD.n6358 1.73383
R29394 VDD.n6622 VDD.n6621 1.73383
R29395 VDD.n6619 VDD.n6618 1.73383
R29396 VDD.n6617 VDD.n6616 1.73383
R29397 VDD.n6612 VDD.n6611 1.73383
R29398 VDD.n6608 VDD.n6607 1.73383
R29399 VDD.n6604 VDD.n6603 1.73383
R29400 VDD.n6601 VDD.n6600 1.73383
R29401 VDD.n7846 VDD.n7845 1.73383
R29402 VDD.n7145 VDD.n7144 1.73383
R29403 VDD.n7149 VDD.n7148 1.73383
R29404 VDD.n7151 VDD.n7150 1.73383
R29405 VDD.n7157 VDD.n7156 1.73383
R29406 VDD.n7159 VDD.n7158 1.73383
R29407 VDD.n7164 VDD.n7163 1.73383
R29408 VDD.n7168 VDD.n7167 1.73383
R29409 VDD.n7170 VDD.n7169 1.73383
R29410 VDD.n7146 VDD.n7145 1.73383
R29411 VDD.n7148 VDD.n7147 1.73383
R29412 VDD.n7152 VDD.n7151 1.73383
R29413 VDD.n7156 VDD.n7155 1.73383
R29414 VDD.n7160 VDD.n7159 1.73383
R29415 VDD.n7165 VDD.n7164 1.73383
R29416 VDD.n7167 VDD.n7166 1.73383
R29417 VDD.n7171 VDD.n7170 1.73383
R29418 VDD.n5431 VDD.n5394 1.73383
R29419 VDD.n5429 VDD.n5395 1.73383
R29420 VDD.n5426 VDD.n5397 1.73383
R29421 VDD.n5421 VDD.n5399 1.73383
R29422 VDD.n5418 VDD.n5400 1.73383
R29423 VDD.n5413 VDD.n5403 1.73383
R29424 VDD.n5411 VDD.n5404 1.73383
R29425 VDD.n5408 VDD.n5406 1.73383
R29426 VDD.n5432 VDD.n5431 1.73383
R29427 VDD.n5429 VDD.n5428 1.73383
R29428 VDD.n5427 VDD.n5426 1.73383
R29429 VDD.n5422 VDD.n5421 1.73383
R29430 VDD.n5418 VDD.n5417 1.73383
R29431 VDD.n5414 VDD.n5413 1.73383
R29432 VDD.n5411 VDD.n5410 1.73383
R29433 VDD.n5409 VDD.n5408 1.73383
R29434 VDD.n8009 VDD.n8008 1.73383
R29435 VDD.n8006 VDD.n8005 1.73383
R29436 VDD.n8004 VDD.n8003 1.73383
R29437 VDD.n7999 VDD.n7998 1.73383
R29438 VDD.n2185 VDD.n2184 1.73383
R29439 VDD.n2181 VDD.n2180 1.73383
R29440 VDD.n2178 VDD.n2177 1.73383
R29441 VDD.n2176 VDD.n2175 1.73383
R29442 VDD.n7971 VDD.n7970 1.73383
R29443 VDD.n7973 VDD.n7972 1.73383
R29444 VDD.n7978 VDD.n7977 1.73383
R29445 VDD.n7984 VDD.n2189 1.73383
R29446 VDD.n7985 VDD.n2192 1.73383
R29447 VDD.n2223 VDD.n2222 1.73383
R29448 VDD.n2231 VDD.n2230 1.73383
R29449 VDD.n2229 VDD.n2228 1.73383
R29450 VDD.n7964 VDD.n7963 1.73383
R29451 VDD.n7982 VDD.n7981 1.73383
R29452 VDD.n7992 VDD.n7991 1.73383
R29453 VDD.n7990 VDD.n7989 1.73383
R29454 VDD.n2225 VDD.n2224 1.73383
R29455 VDD.n2226 VDD.n2212 1.73383
R29456 VDD.n7849 VDD.n7848 1.73383
R29457 VDD.n7847 VDD.n2206 1.73383
R29458 VDD.n6851 VDD.n6850 1.73383
R29459 VDD.n6853 VDD.n6852 1.73383
R29460 VDD.n6856 VDD.n6855 1.73383
R29461 VDD.n6860 VDD.n6859 1.73383
R29462 VDD.n6864 VDD.n6863 1.73383
R29463 VDD.n6869 VDD.n6868 1.73383
R29464 VDD.n6871 VDD.n6870 1.73383
R29465 VDD.n6874 VDD.n6873 1.73383
R29466 VDD.n6726 VDD.n6725 1.73383
R29467 VDD.n6724 VDD.n6723 1.73383
R29468 VDD.n6721 VDD.n6720 1.73383
R29469 VDD.n6717 VDD.n2370 1.73383
R29470 VDD.n7036 VDD.n7035 1.73383
R29471 VDD.n7032 VDD.n7031 1.73383
R29472 VDD.n7029 VDD.n7028 1.73383
R29473 VDD.n7027 VDD.n7026 1.73383
R29474 VDD.n6682 VDD.n6643 1.73383
R29475 VDD.n6680 VDD.n6644 1.73383
R29476 VDD.n6677 VDD.n6646 1.73383
R29477 VDD.n6672 VDD.n6671 1.73383
R29478 VDD.n6670 VDD.n6669 1.73383
R29479 VDD.n6664 VDD.n6651 1.73383
R29480 VDD.n6662 VDD.n6652 1.73383
R29481 VDD.n6659 VDD.n6654 1.73383
R29482 VDD.n7053 VDD.n7052 1.73383
R29483 VDD.n7057 VDD.n7056 1.73383
R29484 VDD.n7059 VDD.n7058 1.73383
R29485 VDD.n7062 VDD.n2333 1.73383
R29486 VDD.n7082 VDD.n2334 1.73383
R29487 VDD.n7077 VDD.n7067 1.73383
R29488 VDD.n7075 VDD.n7068 1.73383
R29489 VDD.n7072 VDD.n7070 1.73383
R29490 VDD.n6683 VDD.n6682 1.73383
R29491 VDD.n6680 VDD.n6679 1.73383
R29492 VDD.n6678 VDD.n6677 1.73383
R29493 VDD.n6673 VDD.n6672 1.73383
R29494 VDD.n6669 VDD.n6668 1.73383
R29495 VDD.n6665 VDD.n6664 1.73383
R29496 VDD.n6662 VDD.n6661 1.73383
R29497 VDD.n6660 VDD.n6659 1.73383
R29498 VDD.n7054 VDD.n7053 1.73383
R29499 VDD.n7056 VDD.n7055 1.73383
R29500 VDD.n7060 VDD.n7059 1.73383
R29501 VDD.n7065 VDD.n2333 1.73383
R29502 VDD.n7082 VDD.n7081 1.73383
R29503 VDD.n7078 VDD.n7077 1.73383
R29504 VDD.n7075 VDD.n7074 1.73383
R29505 VDD.n7073 VDD.n7072 1.73383
R29506 VDD.n7121 VDD.n2325 1.73383
R29507 VDD.n7119 VDD.n2326 1.73383
R29508 VDD.n7116 VDD.n2328 1.73383
R29509 VDD.n7111 VDD.n2330 1.73383
R29510 VDD.n7108 VDD.n7088 1.73383
R29511 VDD.n7103 VDD.n7091 1.73383
R29512 VDD.n7101 VDD.n7092 1.73383
R29513 VDD.n7098 VDD.n7094 1.73383
R29514 VDD.n7122 VDD.n7121 1.73383
R29515 VDD.n7119 VDD.n7118 1.73383
R29516 VDD.n7117 VDD.n7116 1.73383
R29517 VDD.n7112 VDD.n7111 1.73383
R29518 VDD.n7108 VDD.n7107 1.73383
R29519 VDD.n7104 VDD.n7103 1.73383
R29520 VDD.n7101 VDD.n7100 1.73383
R29521 VDD.n7099 VDD.n7098 1.73383
R29522 VDD.n8135 VDD.n8134 1.73383
R29523 VDD.n8163 VDD.n8162 1.73383
R29524 VDD.n8114 VDD.n8113 1.73383
R29525 VDD.n8120 VDD.n8119 1.73383
R29526 VDD.n2046 VDD.n2045 1.73383
R29527 VDD.n2052 VDD.n2051 1.73383
R29528 VDD.n10807 VDD.n10806 1.73383
R29529 VDD.n10801 VDD.n10800 1.73383
R29530 VDD.n8102 VDD.n8101 1.73383
R29531 VDD.n8108 VDD.n8107 1.73383
R29532 VDD.n5583 VDD.n5582 1.73383
R29533 VDD.n5577 VDD.n5576 1.73383
R29534 VDD.n1985 VDD.n1984 1.73383
R29535 VDD.n10813 VDD.n10812 1.73383
R29536 VDD.n1964 VDD.n1963 1.73383
R29537 VDD.n1970 VDD.n1969 1.73383
R29538 VDD.n5604 VDD.n5603 1.73383
R29539 VDD.n5598 VDD.n5597 1.73383
R29540 VDD.n5625 VDD.n5624 1.73383
R29541 VDD.n5619 VDD.n5618 1.73383
R29542 VDD.n10865 VDD.n10864 1.73383
R29543 VDD.n10859 VDD.n10858 1.73383
R29544 VDD.n5508 VDD.n5507 1.73383
R29545 VDD.n10871 VDD.n10870 1.73383
R29546 VDD.n5665 VDD.n5664 1.73383
R29547 VDD.n5659 VDD.n5658 1.73383
R29548 VDD.n5869 VDD.n5868 1.73383
R29549 VDD.n5875 VDD.n5874 1.73383
R29550 VDD.n5520 VDD.n5519 1.73383
R29551 VDD.n5526 VDD.n5525 1.73383
R29552 VDD.n10920 VDD.n10919 1.73383
R29553 VDD.n10914 VDD.n10913 1.73383
R29554 VDD.n5857 VDD.n5856 1.73383
R29555 VDD.n5863 VDD.n5862 1.73383
R29556 VDD.n5814 VDD.n5813 1.73383
R29557 VDD.n5842 VDD.n5841 1.73383
R29558 VDD.n1893 VDD.n1892 1.73383
R29559 VDD.n10926 VDD.n10925 1.73383
R29560 VDD.n1872 VDD.n1871 1.73383
R29561 VDD.n1878 VDD.n1877 1.73383
R29562 VDD.n5802 VDD.n5801 1.73383
R29563 VDD.n5808 VDD.n5807 1.73383
R29564 VDD.n5781 VDD.n5780 1.73383
R29565 VDD.n5787 VDD.n5786 1.73383
R29566 VDD.n10975 VDD.n10974 1.73383
R29567 VDD.n10969 VDD.n10968 1.73383
R29568 VDD.n1828 VDD.n1827 1.73383
R29569 VDD.n10981 VDD.n10980 1.73383
R29570 VDD.n5747 VDD.n5746 1.73383
R29571 VDD.n5775 VDD.n5774 1.73383
R29572 VDD.n5726 VDD.n5725 1.73383
R29573 VDD.n5732 VDD.n5731 1.73383
R29574 VDD.n1816 VDD.n1815 1.73383
R29575 VDD.n1822 VDD.n1821 1.73383
R29576 VDD.n1777 VDD.n1776 1.73383
R29577 VDD.n11024 VDD.n11023 1.73383
R29578 VDD.n11035 VDD.n11034 1.73383
R29579 VDD.n5720 VDD.n5719 1.73383
R29580 VDD.n9072 VDD.n9071 1.73383
R29581 VDD.n9154 VDD.n9153 1.73383
R29582 VDD.n9025 VDD.n9024 1.73383
R29583 VDD.n9030 VDD.n9029 1.73383
R29584 VDD.n8974 VDD.n8973 1.73383
R29585 VDD.n9041 VDD.n9040 1.73383
R29586 VDD.n8950 VDD.n8949 1.73383
R29587 VDD.n9006 VDD.n9005 1.73383
R29588 VDD.n8905 VDD.n8904 1.73383
R29589 VDD.n9019 VDD.n9018 1.73383
R29590 VDD.n8899 VDD.n8898 1.73383
R29591 VDD.n8933 VDD.n8932 1.73383
R29592 VDD.n8847 VDD.n8846 1.73383
R29593 VDD.n8944 VDD.n8943 1.73383
R29594 VDD.n8841 VDD.n8840 1.73383
R29595 VDD.n8875 VDD.n8874 1.73383
R29596 VDD.n8774 VDD.n8773 1.73383
R29597 VDD.n8888 VDD.n8887 1.73383
R29598 VDD.n8768 VDD.n8767 1.73383
R29599 VDD.n8802 VDD.n8801 1.73383
R29600 VDD.n8546 VDD.n8545 1.73383
R29601 VDD.n8835 VDD.n8834 1.73383
R29602 VDD.n8552 VDD.n8551 1.73383
R29603 VDD.n8558 VDD.n8557 1.73383
R29604 VDD.n8756 VDD.n8755 1.73383
R29605 VDD.n8762 VDD.n8761 1.73383
R29606 VDD.n173 VDD.n172 1.73383
R29607 VDD.n189 VDD.n188 1.73383
R29608 VDD.n9094 VDD.n9093 1.73383
R29609 VDD.n9122 VDD.n9121 1.73383
R29610 VDD.n8487 VDD.n8486 1.73383
R29611 VDD.n9165 VDD.n9164 1.73383
R29612 VDD.n9148 VDD.n9147 1.73383
R29613 VDD.n9142 VDD.n9141 1.73383
R29614 VDD.n9132 VDD.n9129 1.73383
R29615 VDD.n9132 VDD.n9131 1.73383
R29616 VDD.n8739 VDD.n8738 1.73383
R29617 VDD.n8745 VDD.n8744 1.73383
R29618 VDD.n8718 VDD.n8717 1.73383
R29619 VDD.n8724 VDD.n8723 1.73383
R29620 VDD.n139 VDD.n138 1.73383
R29621 VDD.n167 VDD.n166 1.73383
R29622 VDD.n12497 VDD.n12496 1.73383
R29623 VDD.n12491 VDD.n12490 1.73383
R29624 VDD.n8706 VDD.n8705 1.73383
R29625 VDD.n8712 VDD.n8711 1.73383
R29626 VDD.n8680 VDD.n8679 1.73383
R29627 VDD.n8686 VDD.n8685 1.73383
R29628 VDD.n93 VDD.n92 1.73383
R29629 VDD.n12503 VDD.n12502 1.73383
R29630 VDD.n50 VDD.n49 1.73383
R29631 VDD.n78 VDD.n77 1.73383
R29632 VDD.n8668 VDD.n8667 1.73383
R29633 VDD.n8674 VDD.n8673 1.73383
R29634 VDD.n8647 VDD.n8646 1.73383
R29635 VDD.n8653 VDD.n8652 1.73383
R29636 VDD.n12553 VDD.n12552 1.73383
R29637 VDD.n12547 VDD.n12546 1.73383
R29638 VDD.n12590 VDD.n12589 1.73383
R29639 VDD.n12597 VDD.n12596 1.73383
R29640 VDD.n12619 VDD.n12618 1.73383
R29641 VDD.n8636 VDD.n8635 1.73383
R29642 VDD.n1562 VDD.n1561 1.73383
R29643 VDD.n1540 VDD.n1539 1.73383
R29644 VDD.n1516 VDD.n1515 1.73383
R29645 VDD.n1527 VDD.n1526 1.73383
R29646 VDD.n1181 VDD.n1180 1.73383
R29647 VDD.n1185 VDD.n1184 1.73383
R29648 VDD.n1168 VDD.n1167 1.73383
R29649 VDD.n1172 VDD.n1171 1.73383
R29650 VDD.n1315 VDD.n1314 1.73383
R29651 VDD.n1656 VDD.n1655 1.73383
R29652 VDD.n1310 VDD.n1309 1.73383
R29653 VDD.n1341 VDD.n1340 1.73383
R29654 VDD.n1361 VDD.n1360 1.73383
R29655 VDD.n1283 VDD.n1082 1.73383
R29656 VDD.n1078 VDD.n1077 1.73383
R29657 VDD.n1388 VDD.n1387 1.73383
R29658 VDD.n1247 VDD.n1246 1.73383
R29659 VDD.n1649 VDD.n1648 1.73383
R29660 VDD.n1602 VDD.n1500 1.73383
R29661 VDD.n1599 VDD.n1501 1.73383
R29662 VDD.n1603 VDD.n1602 1.73383
R29663 VDD.n1599 VDD.n1598 1.73383
R29664 VDD.n1242 VDD.n1241 1.73383
R29665 VDD.n1274 VDD.n1273 1.73383
R29666 VDD.n1211 VDD.n1210 1.73383
R29667 VDD.n1215 VDD.n1214 1.73383
R29668 VDD.n1402 VDD.n1401 1.73383
R29669 VDD.n1411 VDD.n1392 1.73383
R29670 VDD.n1453 VDD.n1452 1.73383
R29671 VDD.n1455 VDD.n1454 1.73383
R29672 VDD.n1488 VDD.n1487 1.73383
R29673 VDD.n1490 VDD.n1489 1.73383
R29674 VDD.n1403 VDD.n1402 1.73383
R29675 VDD.n1411 VDD.n1410 1.73383
R29676 VDD.n1452 VDD.n1451 1.73383
R29677 VDD.n1456 VDD.n1455 1.73383
R29678 VDD.n1487 VDD.n1486 1.73383
R29679 VDD.n1491 VDD.n1490 1.73383
R29680 VDD.n1064 VDD.n1063 1.73383
R29681 VDD.n1068 VDD.n1067 1.73383
R29682 VDD.n909 VDD.n908 1.73383
R29683 VDD.n913 VDD.n912 1.73383
R29684 VDD.n946 VDD.n945 1.73383
R29685 VDD.n1739 VDD.n694 1.73383
R29686 VDD.n947 VDD.n946 1.73383
R29687 VDD.n1739 VDD.n1738 1.73383
R29688 VDD.n724 VDD.n723 1.73383
R29689 VDD.n1715 VDD.n714 1.73383
R29690 VDD.n725 VDD.n724 1.73383
R29691 VDD.n1715 VDD.n1714 1.73383
R29692 VDD.n1747 VDD.n1746 1.73383
R29693 VDD.n1159 VDD.n685 1.73383
R29694 VDD.n1442 VDD.t2748 1.7314
R29695 VDD.n1610 VDD.t2802 1.7314
R29696 VDD.n1610 VDD.t1070 1.7314
R29697 VDD.n1480 VDD.t1532 1.7314
R29698 VDD.n1480 VDD.t4071 1.7314
R29699 VDD.n6157 VDD.n6156 1.69136
R29700 VDD.n6151 VDD.n6037 1.69136
R29701 VDD.n6849 VDD.n6848 1.69136
R29702 VDD.n6841 VDD.n6727 1.69136
R29703 VDD.n6121 VDD.n6019 1.65018
R29704 VDD.n6092 VDD.n6091 1.65018
R29705 VDD.n6840 VDD.n6839 1.65018
R29706 VDD.n6762 VDD.n6758 1.65018
R29707 VDD.n679 VDD.t1172 1.60217
R29708 VDD.n968 VDD.t3582 1.60217
R29709 VDD.n967 VDD.t2547 1.60217
R29710 VDD.n966 VDD.t2670 1.60217
R29711 VDD.n965 VDD.t1434 1.60217
R29712 VDD.n964 VDD.t1562 1.60217
R29713 VDD.n963 VDD.t4611 1.60217
R29714 VDD.n962 VDD.t809 1.60217
R29715 VDD.n961 VDD.t3847 1.60217
R29716 VDD.n960 VDD.t3979 1.60217
R29717 VDD.n959 VDD.t2933 1.60217
R29718 VDD.n958 VDD.t941 1.60217
R29719 VDD.n942 VDD.t687 1.60217
R29720 VDD.n941 VDD.t3331 1.60217
R29721 VDD.n940 VDD.t2228 1.60217
R29722 VDD.n939 VDD.t2624 1.60217
R29723 VDD.n938 VDD.t2501 1.60217
R29724 VDD.n937 VDD.t2630 1.60217
R29725 VDD.n1017 VDD.t1400 1.60217
R29726 VDD.n1018 VDD.t1513 1.60217
R29727 VDD.n1019 VDD.t4545 1.60217
R29728 VDD.n1020 VDD.t2568 1.60217
R29729 VDD.n1021 VDD.t1344 1.60217
R29730 VDD.n12639 VDD.t4001 1.60217
R29731 VDD.n7809 VDD.t3955 1.60217
R29732 VDD.n2252 VDD.t3588 1.60217
R29733 VDD.n2260 VDD.t1082 1.60217
R29734 VDD.n2270 VDD.t1094 1.60217
R29735 VDD.n7725 VDD.t2829 1.60217
R29736 VDD.n2283 VDD.t2455 1.60217
R29737 VDD.n2291 VDD.t2713 1.60217
R29738 VDD.n7826 VDD.t2055 1.60217
R29739 VDD.n7823 VDD.t1665 1.60217
R29740 VDD.n2401 VDD.t2875 1.60217
R29741 VDD.n2399 VDD.t4427 1.60217
R29742 VDD.n2320 VDD.t4093 1.60217
R29743 VDD.n7130 VDD.t995 1.60217
R29744 VDD.n7127 VDD.t4743 1.60217
R29745 VDD.n7125 VDD.t2296 1.60217
R29746 VDD.n2401 VDD.t2529 1.60217
R29747 VDD.n2399 VDD.t4115 1.60217
R29748 VDD.n2320 VDD.t3734 1.60217
R29749 VDD.n7130 VDD.t588 1.60217
R29750 VDD.n7127 VDD.t4397 1.60217
R29751 VDD.n7125 VDD.t1891 1.60217
R29752 VDD.n2323 VDD.t4311 1.60217
R29753 VDD.n2344 VDD.t2019 1.60217
R29754 VDD.n2347 VDD.t1642 1.60217
R29755 VDD.n7044 VDD.t3931 1.60217
R29756 VDD.n7047 VDD.t3563 1.60217
R29757 VDD.n2323 VDD.t3981 1.60217
R29758 VDD.n2344 VDD.t1658 1.60217
R29759 VDD.n2347 VDD.t1287 1.60217
R29760 VDD.n7044 VDD.t3578 1.60217
R29761 VDD.n7047 VDD.t3269 1.60217
R29762 VDD.n6712 VDD.t2873 1.60217
R29763 VDD.n6710 VDD.t4425 1.60217
R29764 VDD.n6707 VDD.t4091 1.60217
R29765 VDD.n6705 VDD.t993 1.60217
R29766 VDD.n6702 VDD.t4741 1.60217
R29767 VDD.n6700 VDD.t2294 1.60217
R29768 VDD.n6712 VDD.t708 1.60217
R29769 VDD.n6710 VDD.t2448 1.60217
R29770 VDD.n6707 VDD.t2001 1.60217
R29771 VDD.n6705 VDD.t3111 1.60217
R29772 VDD.n6702 VDD.t2782 1.60217
R29773 VDD.n6700 VDD.t4331 1.60217
R29774 VDD.n6698 VDD.t4309 1.60217
R29775 VDD.n6696 VDD.t2017 1.60217
R29776 VDD.n6693 VDD.t1640 1.60217
R29777 VDD.n6691 VDD.t3929 1.60217
R29778 VDD.n6688 VDD.t3561 1.60217
R29779 VDD.n6686 VDD.t1062 1.60217
R29780 VDD.n6698 VDD.t2260 1.60217
R29781 VDD.n6696 VDD.t4113 1.60217
R29782 VDD.n6693 VDD.t3732 1.60217
R29783 VDD.n6691 VDD.t1818 1.60217
R29784 VDD.n6688 VDD.t1452 1.60217
R29785 VDD.n6686 VDD.t3189 1.60217
R29786 VDD.n6641 VDD.t1076 1.60217
R29787 VDD.n6639 VDD.t2808 1.60217
R29788 VDD.n6636 VDD.t2438 1.60217
R29789 VDD.n5267 VDD.t2691 1.60217
R29790 VDD.n5436 VDD.t2277 1.60217
R29791 VDD.n5438 VDD.t1955 1.60217
R29792 VDD.n6641 VDD.t3207 1.60217
R29793 VDD.n6639 VDD.t618 1.60217
R29794 VDD.n6636 VDD.t4411 1.60217
R29795 VDD.n5267 VDD.t4679 1.60217
R29796 VDD.n5436 VDD.t4317 1.60217
R29797 VDD.n5438 VDD.t4051 1.60217
R29798 VDD.n5443 VDD.t890 1.60217
R29799 VDD.n5441 VDD.t2606 1.60217
R29800 VDD.n5269 VDD.t2169 1.60217
R29801 VDD.n6630 VDD.t2220 1.60217
R29802 VDD.n6627 VDD.t1808 1.60217
R29803 VDD.n6625 VDD.t3686 1.60217
R29804 VDD.n5443 VDD.t3023 1.60217
R29805 VDD.n5441 VDD.t4559 1.60217
R29806 VDD.n5269 VDD.t4243 1.60217
R29807 VDD.n6630 VDD.t4275 1.60217
R29808 VDD.n6627 VDD.t3921 1.60217
R29809 VDD.n6625 VDD.t1595 1.60217
R29810 VDD.n6265 VDD.t2482 1.60217
R29811 VDD.n5377 VDD.t2051 1.60217
R29812 VDD.n6367 VDD.t2345 1.60217
R29813 VDD.n6364 VDD.t1911 1.60217
R29814 VDD.n6362 VDD.t1624 1.60217
R29815 VDD.n6265 VDD.t3390 1.60217
R29816 VDD.n5377 VDD.t3091 1.60217
R29817 VDD.n6367 VDD.t3305 1.60217
R29818 VDD.n6364 VDD.t3003 1.60217
R29819 VDD.n6362 VDD.t2709 1.60217
R29820 VDD.n5473 VDD.t4691 1.60217
R29821 VDD.n5938 VDD.t2216 1.60217
R29822 VDD.n5941 VDD.t1804 1.60217
R29823 VDD.n5944 VDD.t1857 1.60217
R29824 VDD.n5947 VDD.t1487 1.60217
R29825 VDD.n5949 VDD.t3382 1.60217
R29826 VDD.n5473 VDD.t1502 1.60217
R29827 VDD.n5938 VDD.t3239 1.60217
R29828 VDD.n5941 VDD.t2899 1.60217
R29829 VDD.n5944 VDD.t2953 1.60217
R29830 VDD.n5947 VDD.t2586 1.60217
R29831 VDD.n5949 VDD.t4353 1.60217
R29832 VDD.n6301 VDD.t1010 1.60217
R29833 VDD.n6304 VDD.t591 1.60217
R29834 VDD.n6308 VDD.t899 1.60217
R29835 VDD.n6305 VDD.t4653 1.60217
R29836 VDD.n5984 VDD.t790 1.60217
R29837 VDD.n5987 VDD.t4537 1.60217
R29838 VDD.n6314 VDD.t4595 1.60217
R29839 VDD.n6317 VDD.t4263 1.60217
R29840 VDD.n5979 VDD.t1951 1.60217
R29841 VDD.n6175 VDD.t1068 1.60217
R29842 VDD.n6181 VDD.t2798 1.60217
R29843 VDD.n6184 VDD.t2421 1.60217
R29844 VDD.n6186 VDD.t3406 1.60217
R29845 VDD.n6189 VDD.t3093 1.60217
R29846 VDD.n6191 VDD.t4421 1.60217
R29847 VDD.n6194 VDD.t4087 1.60217
R29848 VDD.n6196 VDD.t2210 1.60217
R29849 VDD.n6199 VDD.t1794 1.60217
R29850 VDD.n5362 VDD.t2559 1.60217
R29851 VDD.n5364 VDD.t4139 1.60217
R29852 VDD.n5367 VDD.t3765 1.60217
R29853 VDD.n5369 VDD.t621 1.60217
R29854 VDD.n5372 VDD.t4423 1.60217
R29855 VDD.n5374 VDD.t1924 1.60217
R29856 VDD.n5362 VDD.t3473 1.60217
R29857 VDD.n5364 VDD.t977 1.60217
R29858 VDD.n5367 VDD.t4735 1.60217
R29859 VDD.n5369 VDD.t1611 1.60217
R29860 VDD.n5372 VDD.t1252 1.60217
R29861 VDD.n5374 VDD.t3011 1.60217
R29862 VDD.n6378 VDD.t4007 1.60217
R29863 VDD.n6376 VDD.t1674 1.60217
R29864 VDD.n6373 VDD.t1309 1.60217
R29865 VDD.n5375 VDD.t3598 1.60217
R29866 VDD.n6218 VDD.t3289 1.60217
R29867 VDD.n6378 VDD.t843 1.60217
R29868 VDD.n6376 VDD.t2774 1.60217
R29869 VDD.n6373 VDD.t2398 1.60217
R29870 VDD.n5375 VDD.t4547 1.60217
R29871 VDD.n6218 VDD.t4239 1.60217
R29872 VDD.n2146 VDD.t1100 1.60217
R29873 VDD.n2157 VDD.t3753 1.60217
R29874 VDD.n2163 VDD.t2173 1.60217
R29875 VDD.n8012 VDD.t914 1.60217
R29876 VDD.n2204 VDD.t1384 1.60217
R29877 VDD.n7863 VDD.t3967 1.60217
R29878 VDD.n7910 VDD.t2308 1.60217
R29879 VDD.n2341 VDD.t2806 1.60217
R29880 VDD.n2360 VDD.t2436 1.60217
R29881 VDD.n2365 VDD.t2689 1.60217
R29882 VDD.n2362 VDD.t2275 1.60217
R29883 VDD.n2311 VDD.t1953 1.60217
R29884 VDD.n2341 VDD.t2453 1.60217
R29885 VDD.n2360 VDD.t2007 1.60217
R29886 VDD.n2365 VDD.t2310 1.60217
R29887 VDD.n2362 VDD.t1882 1.60217
R29888 VDD.n2311 VDD.t1597 1.60217
R29889 VDD.n7141 VDD.t887 1.60217
R29890 VDD.n7139 VDD.t2604 1.60217
R29891 VDD.n7136 VDD.t2167 1.60217
R29892 VDD.n2316 VDD.t2218 1.60217
R29893 VDD.n2313 VDD.t1806 1.60217
R29894 VDD.n7141 VDD.t4665 1.60217
R29895 VDD.n7139 VDD.t2181 1.60217
R29896 VDD.n7136 VDD.t1776 1.60217
R29897 VDD.n2316 VDD.t1829 1.60217
R29898 VDD.n2313 VDD.t1466 1.60217
R29899 VDD.n2296 VDD.t2628 1.60217
R29900 VDD.n2209 VDD.t2196 1.60217
R29901 VDD.n7837 VDD.t2246 1.60217
R29902 VDD.n7840 VDD.t1837 1.60217
R29903 VDD.n7842 VDD.t3712 1.60217
R29904 VDD.n7176 VDD.t2316 1.60217
R29905 VDD.n7946 VDD.t1398 1.60217
R29906 VDD.n7943 VDD.t3987 1.60217
R29907 VDD.n7887 VDD.t2339 1.60217
R29908 VDD.n7888 VDD.t1120 1.60217
R29909 VDD.n8051 VDD.t3781 1.60217
R29910 VDD.n8048 VDD.t2200 1.60217
R29911 VDD.n2172 VDD.t929 1.60217
R29912 VDD.n2390 VDD.t2897 1.60217
R29913 VDD.n2388 VDD.t4459 1.60217
R29914 VDD.n2239 VDD.t4121 1.60217
R29915 VDD.n7831 VDD.t1012 1.60217
R29916 VDD.n7828 VDD.t598 1.60217
R29917 VDD.n1156 VDD.t3608 1.60217
R29918 VDD.n1140 VDD.t4265 1.60217
R29919 VDD.n1141 VDD.t3197 1.60217
R29920 VDD.n1142 VDD.t3303 1.60217
R29921 VDD.n1143 VDD.t2162 1.60217
R29922 VDD.n1144 VDD.t2324 1.60217
R29923 VDD.n705 VDD.t1143 1.60217
R29924 VDD.n704 VDD.t1460 1.60217
R29925 VDD.n703 VDD.t4503 1.60217
R29926 VDD.n702 VDD.t4637 1.60217
R29927 VDD.n701 VDD.t3537 1.60217
R29928 VDD.n1156 VDD.t754 1.60217
R29929 VDD.n1140 VDD.t3915 1.60217
R29930 VDD.n1141 VDD.t2877 1.60217
R29931 VDD.n1142 VDD.t3007 1.60217
R29932 VDD.n1143 VDD.t1774 1.60217
R29933 VDD.n1144 VDD.t1915 1.60217
R29934 VDD.n705 VDD.t819 1.60217
R29935 VDD.n704 VDD.t1133 1.60217
R29936 VDD.n703 VDD.t4193 1.60217
R29937 VDD.n702 VDD.t4295 1.60217
R29938 VDD.n701 VDD.t3245 1.60217
R29939 VDD.n927 VDD.t693 1.60217
R29940 VDD.n926 VDD.t3740 1.60217
R29941 VDD.n925 VDD.t4073 1.60217
R29942 VDD.n924 VDD.t3963 1.60217
R29943 VDD.n923 VDD.t4081 1.60217
R29944 VDD.n922 VDD.t3035 1.60217
R29945 VDD.n921 VDD.t3145 1.60217
R29946 VDD.n920 VDD.t1964 1.60217
R29947 VDD.n919 VDD.t4037 1.60217
R29948 VDD.n918 VDD.t2995 1.60217
R29949 VDD.n917 VDD.t1348 1.60217
R29950 VDD.n927 VDD.t4233 1.60217
R29951 VDD.n926 VDD.t3161 1.60217
R29952 VDD.n925 VDD.t3453 1.60217
R29953 VDD.n924 VDD.t3329 1.60217
R29954 VDD.n923 VDD.t3457 1.60217
R29955 VDD.n922 VDD.t2400 1.60217
R29956 VDD.n921 VDD.t2527 1.60217
R29957 VDD.n920 VDD.t1300 1.60217
R29958 VDD.n919 VDD.t3398 1.60217
R29959 VDD.n918 VDD.t2318 1.60217
R29960 VDD.n917 VDD.t746 1.60217
R29961 VDD.n730 VDD.t2149 1.60217
R29962 VDD.n731 VDD.t1029 1.60217
R29963 VDD.n732 VDD.t1323 1.60217
R29964 VDD.n733 VDD.t1215 1.60217
R29965 VDD.n734 VDD.t1328 1.60217
R29966 VDD.n884 VDD.t4381 1.60217
R29967 VDD.n883 VDD.t4499 1.60217
R29968 VDD.n882 VDD.t3422 1.60217
R29969 VDD.n881 VDD.t1283 1.60217
R29970 VDD.n880 VDD.t4347 1.60217
R29971 VDD.n879 VDD.t2891 1.60217
R29972 VDD.n730 VDD.t1476 1.60217
R29973 VDD.n731 VDD.t4515 1.60217
R29974 VDD.n732 VDD.t713 1.60217
R29975 VDD.n733 VDD.t4737 1.60217
R29976 VDD.n734 VDD.t715 1.60217
R29977 VDD.n884 VDD.t3767 1.60217
R29978 VDD.n883 VDD.t3887 1.60217
R29979 VDD.n882 VDD.t2853 1.60217
R29980 VDD.n881 VDD.t661 1.60217
R29981 VDD.n880 VDD.t3706 1.60217
R29982 VDD.n879 VDD.t2198 1.60217
R29983 VDD.n1462 VDD.t4215 1.60217
R29984 VDD.n1463 VDD.t3149 1.60217
R29985 VDD.n1464 VDD.t3429 1.60217
R29986 VDD.n1465 VDD.t3325 1.60217
R29987 VDD.n1466 VDD.t3437 1.60217
R29988 VDD.n1292 VDD.t2371 1.60217
R29989 VDD.n1291 VDD.t2511 1.60217
R29990 VDD.n1290 VDD.t1281 1.60217
R29991 VDD.n1289 VDD.t3364 1.60217
R29992 VDD.n1288 VDD.t2279 1.60217
R29993 VDD.n1287 VDD.t704 1.60217
R29994 VDD.n1462 VDD.t822 1.60217
R29995 VDD.n1463 VDD.t3857 1.60217
R29996 VDD.n1464 VDD.t4201 1.60217
R29997 VDD.n1465 VDD.t4067 1.60217
R29998 VDD.n1466 VDD.t4209 1.60217
R29999 VDD.n1292 VDD.t3139 1.60217
R30000 VDD.n1291 VDD.t3253 1.60217
R30001 VDD.n1290 VDD.t2094 1.60217
R30002 VDD.n1289 VDD.t4155 1.60217
R30003 VDD.n1288 VDD.t3089 1.60217
R30004 VDD.n1287 VDD.t1458 1.60217
R30005 VDD.n1235 VDD.t1787 1.60217
R30006 VDD.n1220 VDD.t3671 1.60217
R30007 VDD.n1221 VDD.t2650 1.60217
R30008 VDD.n1222 VDD.t2784 1.60217
R30009 VDD.n1223 VDD.t1536 1.60217
R30010 VDD.n1224 VDD.t1670 1.60217
R30011 VDD.n1092 VDD.t4719 1.60217
R30012 VDD.n1093 VDD.t926 1.60217
R30013 VDD.n1094 VDD.t3957 1.60217
R30014 VDD.n1235 VDD.t4205 1.60217
R30015 VDD.n1220 VDD.t2361 1.60217
R30016 VDD.n1221 VDD.t1152 1.60217
R30017 VDD.n1222 VDD.t1271 1.60217
R30018 VDD.n1223 VDD.t4335 1.60217
R30019 VDD.n1224 VDD.t4447 1.60217
R30020 VDD.n1092 VDD.t3345 1.60217
R30021 VDD.n1093 VDD.t3657 1.60217
R30022 VDD.n1094 VDD.t2640 1.60217
R30023 VDD.n1268 VDD.t2907 1.60217
R30024 VDD.n1252 VDD.t666 1.60217
R30025 VDD.n1253 VDD.t3716 1.60217
R30026 VDD.n1254 VDD.t3839 1.60217
R30027 VDD.n1255 VDD.t2812 1.60217
R30028 VDD.n1256 VDD.t2919 1.60217
R30029 VDD.n785 VDD.t1698 1.60217
R30030 VDD.n786 VDD.t2073 1.60217
R30031 VDD.n787 VDD.t961 1.60217
R30032 VDD.n1268 VDD.t1043 1.60217
R30033 VDD.n1252 VDD.t3467 1.60217
R30034 VDD.n1253 VDD.t2407 1.60217
R30035 VDD.n1254 VDD.t2533 1.60217
R30036 VDD.n1255 VDD.t1305 1.60217
R30037 VDD.n1256 VDD.t1430 1.60217
R30038 VDD.n785 VDD.t4477 1.60217
R30039 VDD.n786 VDD.t658 1.60217
R30040 VDD.n787 VDD.t3700 1.60217
R30041 VDD.n1577 VDD.t2465 1.60217
R30042 VDD.n1578 VDD.t1240 1.60217
R30043 VDD.n1579 VDD.t1570 1.60217
R30044 VDD.n1580 VDD.t1448 1.60217
R30045 VDD.n1581 VDD.t1581 1.60217
R30046 VDD.n748 VDD.t4621 1.60217
R30047 VDD.n749 VDD.t4745 1.60217
R30048 VDD.n750 VDD.t3633 1.60217
R30049 VDD.n1505 VDD.t2756 1.60217
R30050 VDD.n1509 VDD.t579 1.60217
R30051 VDD.n1508 VDD.t3643 1.60217
R30052 VDD.n1639 VDD.t4523 1.60217
R30053 VDD.n775 VDD.t4589 1.60217
R30054 VDD.n1519 VDD.t1080 1.60217
R30055 VDD.n780 VDD.t924 1.60217
R30056 VDD.n1566 VDD.t3875 1.60217
R30057 VDD.n769 VDD.t3410 1.60217
R30058 VDD.n773 VDD.t2326 1.60217
R30059 VDD.n776 VDD.t2484 1.60217
R30060 VDD.n778 VDD.t1259 1.60217
R30061 VDD.n781 VDD.t1390 1.60217
R30062 VDD.n1565 VDD.t4429 1.60217
R30063 VDD.n1523 VDD.t3017 1.60217
R30064 VDD.n1522 VDD.t3061 1.60217
R30065 VDD.n1547 VDD.t3604 1.60217
R30066 VDD.n1534 VDD.t3445 1.60217
R30067 VDD.n1535 VDD.t2303 1.60217
R30068 VDD.n1134 VDD.t954 1.60217
R30069 VDD.n1119 VDD.t3627 1.60217
R30070 VDD.n1120 VDD.t2608 1.60217
R30071 VDD.n1121 VDD.t2727 1.60217
R30072 VDD.n1122 VDD.t1500 1.60217
R30073 VDD.n1123 VDD.t1632 1.60217
R30074 VDD.n860 VDD.t4681 1.60217
R30075 VDD.n861 VDD.t882 1.60217
R30076 VDD.n862 VDD.t3905 1.60217
R30077 VDD.n863 VDD.t4039 1.60217
R30078 VDD.n864 VDD.t2999 1.60217
R30079 VDD.n1134 VDD.t2248 1.60217
R30080 VDD.n1119 VDD.t3319 1.60217
R30081 VDD.n1120 VDD.t2191 1.60217
R30082 VDD.n1121 VDD.t2369 1.60217
R30083 VDD.n1122 VDD.t1163 1.60217
R30084 VDD.n1123 VDD.t1277 1.60217
R30085 VDD.n860 VDD.t4339 1.60217
R30086 VDD.n861 VDD.t4659 1.60217
R30087 VDD.n862 VDD.t3555 1.60217
R30088 VDD.n863 VDD.t3667 1.60217
R30089 VDD.n864 VDD.t2648 1.60217
R30090 VDD.n1205 VDD.t4181 1.60217
R30091 VDD.n1190 VDD.t3724 1.60217
R30092 VDD.n1191 VDD.t2699 1.60217
R30093 VDD.n1192 VDD.t2821 1.60217
R30094 VDD.n1193 VDD.t1601 1.60217
R30095 VDD.n1194 VDD.t1719 1.60217
R30096 VDD.n843 VDD.t595 1.60217
R30097 VDD.n842 VDD.t985 1.60217
R30098 VDD.n841 VDD.t4011 1.60217
R30099 VDD.n840 VDD.t4137 1.60217
R30100 VDD.n1205 VDD.t1273 1.60217
R30101 VDD.n1190 VDD.t3388 1.60217
R30102 VDD.n1191 VDD.t2314 1.60217
R30103 VDD.n1192 VDD.t2478 1.60217
R30104 VDD.n1193 VDD.t1257 1.60217
R30105 VDD.n1194 VDD.t1379 1.60217
R30106 VDD.n843 VDD.t4415 1.60217
R30107 VDD.n842 VDD.t562 1.60217
R30108 VDD.n841 VDD.t3635 1.60217
R30109 VDD.n840 VDD.t3775 1.60217
R30110 VDD.n788 VDD.t3969 1.60217
R30111 VDD.n789 VDD.t2917 1.60217
R30112 VDD.n790 VDD.t3227 1.60217
R30113 VDD.n791 VDD.t3117 1.60217
R30114 VDD.n792 VDD.t3233 1.60217
R30115 VDD.n1324 VDD.t2075 1.60217
R30116 VDD.n1323 VDD.t2202 1.60217
R30117 VDD.n1322 VDD.t1072 1.60217
R30118 VDD.n1321 VDD.t3181 1.60217
R30119 VDD.n1320 VDD.t2003 1.60217
R30120 VDD.n1319 VDD.t4609 1.60217
R30121 VDD.n788 VDD.t4717 1.60217
R30122 VDD.n789 VDD.t3619 1.60217
R30123 VDD.n790 VDD.t3953 1.60217
R30124 VDD.n791 VDD.t3823 1.60217
R30125 VDD.n792 VDD.t3961 1.60217
R30126 VDD.n1324 VDD.t2911 1.60217
R30127 VDD.n1323 VDD.t3033 1.60217
R30128 VDD.n1322 VDD.t1814 1.60217
R30129 VDD.n1321 VDD.t3895 1.60217
R30130 VDD.n1320 VDD.t2859 1.60217
R30131 VDD.n1319 VDD.t1224 1.60217
R30132 VDD.n753 VDD.t4553 1.60217
R30133 VDD.n825 VDD.t2476 1.60217
R30134 VDD.n826 VDD.t1250 1.60217
R30135 VDD.n827 VDD.t1585 1.60217
R30136 VDD.n828 VDD.t1456 1.60217
R30137 VDD.n829 VDD.t1589 1.60217
R30138 VDD.n1370 VDD.t4633 1.60217
R30139 VDD.n1369 VDD.t568 1.60217
R30140 VDD.n1368 VDD.t3637 1.60217
R30141 VDD.n1367 VDD.t1526 1.60217
R30142 VDD.n1366 VDD.t4565 1.60217
R30143 VDD.n1365 VDD.t3121 1.60217
R30144 VDD.n825 VDD.t1723 1.60217
R30145 VDD.n826 VDD.t610 1.60217
R30146 VDD.n827 VDD.t991 1.60217
R30147 VDD.n828 VDD.t874 1.60217
R30148 VDD.n829 VDD.t1000 1.60217
R30149 VDD.n1370 VDD.t4023 1.60217
R30150 VDD.n1369 VDD.t4147 1.60217
R30151 VDD.n1368 VDD.t3087 1.60217
R30152 VDD.n1367 VDD.t943 1.60217
R30153 VDD.n1366 VDD.t3973 1.60217
R30154 VDD.n1365 VDD.t2515 1.60217
R30155 VDD.n6999 VDD.n6998 1.60175
R30156 VDD.n6523 VDD.n6522 1.60175
R30157 VDD.n72 VDD.n71 1.59478
R30158 VDD.n161 VDD.n160 1.59478
R30159 VDD.n5771 VDD.n5770 1.59478
R30160 VDD.n5838 VDD.n5837 1.59478
R30161 VDD.n5655 VDD.n5654 1.59478
R30162 VDD.n5573 VDD.n5572 1.59478
R30163 VDD.n8159 VDD.n8158 1.59478
R30164 VDD.n9116 VDD.n9115 1.59478
R30165 VDD.n8829 VDD.n8828 1.59478
R30166 VDD.n8969 VDD.n8968 1.59478
R30167 VDD.n751 VDD.t1522 1.58642
R30168 VDD.n1506 VDD.t3785 1.58642
R30169 VDD.n7956 VDD.n7954 1.57603
R30170 VDD.n8061 VDD.n8059 1.57603
R30171 VDD.n2356 VDD.n2317 1.56483
R30172 VDD.n1441 VDD.t3075 1.55829
R30173 VDD.n804 VDD.t4125 1.55829
R30174 VDD.n803 VDD.t3837 1.55829
R30175 VDD.n1479 VDD.t3031 1.55829
R30176 VDD.n814 VDD.t2766 1.55829
R30177 VDD.n6014 VDD.n6013 1.52779
R30178 VDD.n7005 VDD.n2376 1.5005
R30179 VDD.n6976 VDD.n6975 1.5005
R30180 VDD.n6978 VDD.n6977 1.5005
R30181 VDD.n7023 VDD.n7022 1.5005
R30182 VDD.n6959 VDD.n6958 1.5005
R30183 VDD.n6549 VDD.n6548 1.5005
R30184 VDD.n6512 VDD.n6415 1.5005
R30185 VDD.n6536 VDD.n6535 1.5005
R30186 VDD.n6551 VDD.n6550 1.5005
R30187 VDD.n6497 VDD.n6496 1.5005
R30188 VDD.n6095 VDD.n6038 1.5005
R30189 VDD.n6117 VDD.n6116 1.5005
R30190 VDD.n6152 VDD.n6151 1.5005
R30191 VDD.n6075 VDD.n6074 1.5005
R30192 VDD.n6150 VDD.n6149 1.5005
R30193 VDD.n6798 VDD.n6797 1.5005
R30194 VDD.n6800 VDD.n6799 1.5005
R30195 VDD.n6848 VDD.n6847 1.5005
R30196 VDD.n6791 VDD.n6790 1.5005
R30197 VDD.n6823 VDD.n2405 1.5005
R30198 VDD.n8642 VDD.n8640 1.49396
R30199 VDD.n8701 VDD.n8699 1.49396
R30200 VDD.n1811 VDD.n1809 1.49396
R30201 VDD.n1867 VDD.n1865 1.49396
R30202 VDD.n5515 VDD.n5513 1.49396
R30203 VDD.n1959 VDD.n1957 1.49396
R30204 VDD.n2041 VDD.n2039 1.49396
R30205 VDD.n8751 VDD.n8749 1.49396
R30206 VDD.n8894 VDD.n8892 1.49396
R30207 VDD.n9067 VDD.n9065 1.49396
R30208 VDD.n8636 VDD.t2642 1.4705
R30209 VDD.t1810 VDD.n8636 1.4705
R30210 VDD.t2666 VDD.n12619 1.4705
R30211 VDD.n12619 VDD.t1468 1.4705
R30212 VDD.n12597 VDD.t756 1.4705
R30213 VDD.t4189 VDD.n12597 1.4705
R30214 VDD.n12590 VDD.t781 1.4705
R30215 VDD.t3829 VDD.n12590 1.4705
R30216 VDD.t849 VDD.n12547 1.4705
R30217 VDD.n12547 VDD.t4267 1.4705
R30218 VDD.t1294 VDD.n12553 1.4705
R30219 VDD.n12553 VDD.t3917 1.4705
R30220 VDD.n8653 VDD.t2736 1.4705
R30221 VDD.t1907 VDD.n8653 1.4705
R30222 VDD.n8647 VDD.t3191 1.4705
R30223 VDD.t1543 VDD.n8647 1.4705
R30224 VDD.n8674 VDD.t731 1.4705
R30225 VDD.t3682 VDD.n8674 1.4705
R30226 VDD.n8668 VDD.t767 1.4705
R30227 VDD.t3347 VDD.n8668 1.4705
R30228 VDD.n78 VDD.t3129 1.4705
R30229 VDD.t1855 VDD.n78 1.4705
R30230 VDD.n50 VDD.t3153 1.4705
R30231 VDD.t1495 VDD.n50 1.4705
R30232 VDD.n12503 VDD.t2426 1.4705
R30233 VDD.t799 VDD.n12503 1.4705
R30234 VDD.n93 VDD.t1999 1.4705
R30235 VDD.t2244 VDD.n93 1.4705
R30236 VDD.n8686 VDD.t4183 1.4705
R30237 VDD.t2685 VDD.n8686 1.4705
R30238 VDD.n8680 VDD.t3819 1.4705
R30239 VDD.t4049 VDD.n8680 1.4705
R30240 VDD.n8712 VDD.t4261 1.4705
R30241 VDD.t2790 VDD.n8712 1.4705
R30242 VDD.n8706 VDD.t1406 1.4705
R30243 VDD.t1634 VDD.n8706 1.4705
R30244 VDD.t2525 VDD.n12491 1.4705
R30245 VDD.n12491 VDD.t906 1.4705
R30246 VDD.t3773 VDD.n12497 1.4705
R30247 VDD.n12497 VDD.t3997 1.4705
R30248 VDD.n167 VDD.t4229 1.4705
R30249 VDD.t2732 VDD.n167 1.4705
R30250 VDD.n139 VDD.t3859 1.4705
R30251 VDD.t4079 VDD.n139 1.4705
R30252 VDD.n8724 VDD.t1853 1.4705
R30253 VDD.t4455 VDD.n8724 1.4705
R30254 VDD.n8718 VDD.t1490 1.4705
R30255 VDD.t1711 VDD.n8718 1.4705
R30256 VDD.n8745 VDD.t3851 1.4705
R30257 VDD.t2348 VDD.n8745 1.4705
R30258 VDD.n8739 VDD.t2101 1.4705
R30259 VDD.t2386 VDD.n8739 1.4705
R30260 VDD.n5720 VDD.t1756 1.4705
R30261 VDD.t4223 VDD.n5720 1.4705
R30262 VDD.t3592 VDD.n11035 1.4705
R30263 VDD.n11035 VDD.t1244 1.4705
R30264 VDD.t2616 VDD.n11024 1.4705
R30265 VDD.n11024 VDD.t3694 1.4705
R30266 VDD.n1777 VDD.t3947 1.4705
R30267 VDD.t585 VDD.n1777 1.4705
R30268 VDD.n1822 VDD.t3317 1.4705
R30269 VDD.t4453 VDD.n1822 1.4705
R30270 VDD.n1816 VDD.t1556 1.4705
R30271 VDD.t1360 VDD.n1816 1.4705
R30272 VDD.n5732 VDD.t1228 1.4705
R30273 VDD.t3649 VDD.n5732 1.4705
R30274 VDD.n5726 VDD.t1618 1.4705
R30275 VDD.t733 VDD.n5726 1.4705
R30276 VDD.n5775 VDD.t1663 1.4705
R30277 VDD.t1319 VDD.n5775 1.4705
R30278 VDD.n5747 VDD.t3491 1.4705
R30279 VDD.t2658 VDD.n5747 1.4705
R30280 VDD.n10981 VDD.t1388 1.4705
R30281 VDD.t1504 VDD.n10981 1.4705
R30282 VDD.n1828 VDD.t2889 1.4705
R30283 VDD.t2693 VDD.n1828 1.4705
R30284 VDD.t1332 VDD.n10969 1.4705
R30285 VDD.n10969 VDD.t1139 1.4705
R30286 VDD.t2521 VDD.n10975 1.4705
R30287 VDD.n10975 VDD.t3629 1.4705
R30288 VDD.n5787 VDD.t2367 1.4705
R30289 VDD.t1364 VDD.n5787 1.4705
R30290 VDD.n5781 VDD.t3525 1.4705
R30291 VDD.t2144 VDD.n5781 1.4705
R30292 VDD.n5808 VDD.t1729 1.4705
R30293 VDD.t872 VDD.n5808 1.4705
R30294 VDD.n5802 VDD.t1178 1.4705
R30295 VDD.t3985 VDD.n5802 1.4705
R30296 VDD.n1878 VDD.t2120 1.4705
R30297 VDD.t1902 VDD.n1878 1.4705
R30298 VDD.n1872 VDD.t3655 1.4705
R30299 VDD.t706 VDD.n1872 1.4705
R30300 VDD.n10926 VDD.t3356 1.4705
R30301 VDD.t3201 VDD.n10926 1.4705
R30302 VDD.n1893 VDD.t4403 1.4705
R30303 VDD.t1446 VDD.n1893 1.4705
R30304 VDD.n5842 VDD.t3594 1.4705
R30305 VDD.t2777 VDD.n5842 1.4705
R30306 VDD.n5814 VDD.t648 1.4705
R30307 VDD.t3459 VDD.n5814 1.4705
R30308 VDD.n5863 VDD.t3751 1.4705
R30309 VDD.t2927 VDD.n5863 1.4705
R30310 VDD.n5857 VDD.t1844 1.4705
R30311 VDD.t4627 VDD.n5857 1.4705
R30312 VDD.t3572 VDD.n10914 1.4705
R30313 VDD.n10914 VDD.t3370 1.4705
R30314 VDD.t3569 VDD.n10920 1.4705
R30315 VDD.n10920 VDD.t576 1.4705
R30316 VDD.n5526 VDD.t3400 1.4705
R30317 VDD.t4563 VDD.n5526 1.4705
R30318 VDD.n5520 VDD.t612 1.4705
R30319 VDD.t2975 VDD.n5520 1.4705
R30320 VDD.n5875 VDD.t1889 1.4705
R30321 VDD.t4677 VDD.n5875 1.4705
R30322 VDD.n5869 VDD.t3698 1.4705
R30323 VDD.t936 VDD.n5869 1.4705
R30324 VDD.t1342 VDD.n5659 1.4705
R30325 VDD.n5659 VDD.t2819 1.4705
R30326 VDD.t3215 VDD.n5665 1.4705
R30327 VDD.n5665 VDD.t870 1.4705
R30328 VDD.n10871 VDD.t4165 1.4705
R30329 VDD.t2265 VDD.n10871 1.4705
R30330 VDD.t1382 VDD.n5508 1.4705
R30331 VDD.n5508 VDD.t2262 1.4705
R30332 VDD.t668 VDD.n10859 1.4705
R30333 VDD.n10859 VDD.t2545 1.4705
R30334 VDD.t2098 VDD.n10865 1.4705
R30335 VDD.n10865 VDD.t3015 1.4705
R30336 VDD.t3907 VDD.n5619 1.4705
R30337 VDD.n5619 VDD.t2985 1.4705
R30338 VDD.t1515 VDD.n5625 1.4705
R30339 VDD.n5625 VDD.t3392 1.4705
R30340 VDD.t3366 VDD.n5598 1.4705
R30341 VDD.n5598 VDD.t4725 1.4705
R30342 VDD.t3749 VDD.n5604 1.4705
R30343 VDD.n5604 VDD.t2924 1.4705
R30344 VDD.n1970 VDD.t1409 1.4705
R30345 VDD.t3680 VDD.n1970 1.4705
R30346 VDD.n1964 VDD.t3889 1.4705
R30347 VDD.t3677 VDD.n1964 1.4705
R30348 VDD.n10813 VDD.t3291 1.4705
R30349 VDD.t4437 VDD.n10813 1.4705
R30350 VDD.n1985 VDD.t4635 1.4705
R30351 VDD.t4433 VDD.n1985 1.4705
R30352 VDD.t1394 VDD.n5577 1.4705
R30353 VDD.n5577 VDD.t4211 1.4705
R30354 VDD.t3267 VDD.n5583 1.4705
R30355 VDD.n5583 VDD.t2381 1.4705
R30356 VDD.n8108 VDD.t865 1.4705
R30357 VDD.t4107 VDD.n8108 1.4705
R30358 VDD.n8102 VDD.t2085 1.4705
R30359 VDD.t675 VDD.n8102 1.4705
R30360 VDD.t2939 VDD.n10801 1.4705
R30361 VDD.n10801 VDD.t2742 1.4705
R30362 VDD.t3939 VDD.n10807 1.4705
R30363 VDD.n10807 VDD.t1004 1.4705
R30364 VDD.n2052 VDD.t3615 1.4705
R30365 VDD.t3425 VDD.n2052 1.4705
R30366 VDD.n2046 VDD.t4683 1.4705
R30367 VDD.t1714 VDD.n2046 1.4705
R30368 VDD.n8120 VDD.t4451 1.4705
R30369 VDD.t3551 VDD.n8120 1.4705
R30370 VDD.n8114 VDD.t1498 1.4705
R30371 VDD.t4299 VDD.n8114 1.4705
R30372 VDD.n8163 VDD.t2151 1.4705
R30373 VDD.t1207 VDD.n8163 1.4705
R30374 VDD.n8135 VDD.t3368 1.4705
R30375 VDD.t1982 VDD.n8135 1.4705
R30376 VDD.t673 VDD.n10770 1.4705
R30377 VDD.n10770 VDD.t4617 1.4705
R30378 VDD.n2058 VDD.t1733 1.4705
R30379 VDD.t3041 VDD.n2058 1.4705
R30380 VDD.t3965 VDD.n7099 1.4705
R30381 VDD.n7099 VDD.t3109 1.4705
R30382 VDD.n7100 VDD.t1150 1.4705
R30383 VDD.n7100 VDD.t3965 1.4705
R30384 VDD.t3971 VDD.n7104 1.4705
R30385 VDD.n7104 VDD.t1150 1.4705
R30386 VDD.n7107 VDD.t4701 1.4705
R30387 VDD.n7107 VDD.t3047 1.4705
R30388 VDD.t1922 VDD.n7112 1.4705
R30389 VDD.n7112 VDD.t4701 1.4705
R30390 VDD.t3726 VDD.n7117 1.4705
R30391 VDD.n7117 VDD.t2428 1.4705
R30392 VDD.n7118 VDD.t975 1.4705
R30393 VDD.n7118 VDD.t3726 1.4705
R30394 VDD.t2250 VDD.n7122 1.4705
R30395 VDD.n7122 VDD.t975 1.4705
R30396 VDD.n7094 VDD.t1833 1.4705
R30397 VDD.t973 VDD.n7094 1.4705
R30398 VDD.n7092 VDD.t3283 1.4705
R30399 VDD.t1833 VDD.n7092 1.4705
R30400 VDD.n7091 VDD.t1841 1.4705
R30401 VDD.t3283 VDD.n7091 1.4705
R30402 VDD.n7088 VDD.t2703 1.4705
R30403 VDD.t904 VDD.n7088 1.4705
R30404 VDD.n2330 VDD.t4005 1.4705
R30405 VDD.t2703 VDD.n2330 1.4705
R30406 VDD.n2328 VDD.t1616 1.4705
R30407 VDD.t4393 VDD.n2328 1.4705
R30408 VDD.n2326 VDD.t3083 1.4705
R30409 VDD.t1616 VDD.n2326 1.4705
R30410 VDD.n2325 VDD.t4285 1.4705
R30411 VDD.t3083 VDD.n2325 1.4705
R30412 VDD.t2833 VDD.n7073 1.4705
R30413 VDD.n7073 VDD.t1816 1.4705
R30414 VDD.n7074 VDD.t4143 1.4705
R30415 VDD.n7074 VDD.t2833 1.4705
R30416 VDD.t2841 VDD.n7078 1.4705
R30417 VDD.n7078 VDD.t4143 1.4705
R30418 VDD.n7081 VDD.t3521 1.4705
R30419 VDD.n7081 VDD.t1737 1.4705
R30420 VDD.n7065 VDD.t735 1.4705
R30421 VDD.t3521 VDD.n7065 1.4705
R30422 VDD.n7060 VDD.t2618 1.4705
R30423 VDD.t1135 VDD.n7060 1.4705
R30424 VDD.n7055 VDD.t3909 1.4705
R30425 VDD.n7055 VDD.t2618 1.4705
R30426 VDD.n7054 VDD.t1025 1.4705
R30427 VDD.t3909 VDD.n7054 1.4705
R30428 VDD.t2931 VDD.n6660 1.4705
R30429 VDD.n6660 VDD.t1438 1.4705
R30430 VDD.n6661 VDD.t3757 1.4705
R30431 VDD.n6661 VDD.t2931 1.4705
R30432 VDD.t1317 VDD.n6665 1.4705
R30433 VDD.n6665 VDD.t3757 1.4705
R30434 VDD.n6668 VDD.t3193 1.4705
R30435 VDD.n6668 VDD.t834 1.4705
R30436 VDD.t4493 VDD.n6673 1.4705
R30437 VDD.n6673 VDD.t3193 1.4705
R30438 VDD.t1113 VDD.n6678 1.4705
R30439 VDD.n6678 VDD.t4013 1.4705
R30440 VDD.n6679 VDD.t2578 1.4705
R30441 VDD.n6679 VDD.t1113 1.4705
R30442 VDD.t3416 VDD.n6683 1.4705
R30443 VDD.n6683 VDD.t2578 1.4705
R30444 VDD.n7070 VDD.t2849 1.4705
R30445 VDD.n7070 VDD.t1835 1.4705
R30446 VDD.n7068 VDD.t4159 1.4705
R30447 VDD.t2849 VDD.n7068 1.4705
R30448 VDD.n7067 VDD.t2855 1.4705
R30449 VDD.t4159 VDD.n7067 1.4705
R30450 VDD.t3533 VDD.n2334 1.4705
R30451 VDD.t1752 VDD.n2334 1.4705
R30452 VDD.t761 VDD.n7062 1.4705
R30453 VDD.n7062 VDD.t3533 1.4705
R30454 VDD.n7058 VDD.t2634 1.4705
R30455 VDD.n7058 VDD.t1148 1.4705
R30456 VDD.n7057 VDD.t3927 1.4705
R30457 VDD.t2634 VDD.n7057 1.4705
R30458 VDD.n7052 VDD.t1037 1.4705
R30459 VDD.n7052 VDD.t3927 1.4705
R30460 VDD.n6654 VDD.t2959 1.4705
R30461 VDD.t1470 VDD.n6654 1.4705
R30462 VDD.n6652 VDD.t3777 1.4705
R30463 VDD.t2959 VDD.n6652 1.4705
R30464 VDD.n6651 VDD.t1330 1.4705
R30465 VDD.t3777 VDD.n6651 1.4705
R30466 VDD.t3213 VDD.n6670 1.4705
R30467 VDD.n6670 VDD.t861 1.4705
R30468 VDD.n6671 VDD.t4507 1.4705
R30469 VDD.n6671 VDD.t3213 1.4705
R30470 VDD.n6646 VDD.t1124 1.4705
R30471 VDD.t4027 VDD.n6646 1.4705
R30472 VDD.n6644 VDD.t2596 1.4705
R30473 VDD.t1124 VDD.n6644 1.4705
R30474 VDD.n6643 VDD.t3431 1.4705
R30475 VDD.t2596 VDD.n6643 1.4705
R30476 VDD.t4555 VDD.n7027 1.4705
R30477 VDD.n7027 VDD.t3271 1.4705
R30478 VDD.n7028 VDD.t1315 1.4705
R30479 VDD.n7028 VDD.t4555 1.4705
R30480 VDD.t3151 VDD.n7032 1.4705
R30481 VDD.n7032 VDD.t1315 1.4705
R30482 VDD.n7035 VDD.t726 1.4705
R30483 VDD.n7035 VDD.t2652 1.4705
R30484 VDD.t2106 VDD.n6717 1.4705
R30485 VDD.n6717 VDD.t726 1.4705
R30486 VDD.n6720 VDD.t2947 1.4705
R30487 VDD.n6720 VDD.t1554 1.4705
R30488 VDD.t4245 VDD.n6724 1.4705
R30489 VDD.n6724 VDD.t2947 1.4705
R30490 VDD.n6725 VDD.t1008 1.4705
R30491 VDD.n6725 VDD.t4245 1.4705
R30492 VDD.n6742 VDD.t226 1.4705
R30493 VDD.n6742 VDD.t92 1.4705
R30494 VDD.n6750 VDD.t246 1.4705
R30495 VDD.n6750 VDD.t149 1.4705
R30496 VDD.n6874 VDD.t4475 1.4705
R30497 VDD.t3590 VDD.n6874 1.4705
R30498 VDD.n6870 VDD.t1690 1.4705
R30499 VDD.n6870 VDD.t4475 1.4705
R30500 VDD.n6869 VDD.t4479 1.4705
R30501 VDD.t1690 VDD.n6869 1.4705
R30502 VDD.n6864 VDD.t1096 1.4705
R30503 VDD.t3515 VDD.n6864 1.4705
R30504 VDD.n6859 VDD.t2557 1.4705
R30505 VDD.n6859 VDD.t1096 1.4705
R30506 VDD.n6856 VDD.t4269 1.4705
R30507 VDD.t2977 VDD.n6856 1.4705
R30508 VDD.n6852 VDD.t1464 1.4705
R30509 VDD.n6852 VDD.t4269 1.4705
R30510 VDD.n6851 VDD.t2845 1.4705
R30511 VDD.t1464 VDD.n6851 1.4705
R30512 VDD.n6954 VDD.t256 1.4705
R30513 VDD.n6954 VDD.t98 1.4705
R30514 VDD.n6955 VDD.t133 1.4705
R30515 VDD.n6955 VDD.t208 1.4705
R30516 VDD.n6922 VDD.t273 1.4705
R30517 VDD.n6922 VDD.t122 1.4705
R30518 VDD.n6923 VDD.t155 1.4705
R30519 VDD.n6923 VDD.t227 1.4705
R30520 VDD.n7014 VDD.t223 1.4705
R30521 VDD.n7014 VDD.t267 1.4705
R30522 VDD.n7016 VDD.t221 1.4705
R30523 VDD.n7016 VDD.t146 1.4705
R30524 VDD.n7018 VDD.t229 1.4705
R30525 VDD.n7018 VDD.t66 1.4705
R30526 VDD.n7020 VDD.t83 1.4705
R30527 VDD.n7020 VDD.t157 1.4705
R30528 VDD.n2382 VDD.t214 1.4705
R30529 VDD.n2382 VDD.t285 1.4705
R30530 VDD.n2380 VDD.t51 1.4705
R30531 VDD.n2380 VDD.t165 1.4705
R30532 VDD.n2378 VDD.t72 1.4705
R30533 VDD.n2378 VDD.t154 1.4705
R30534 VDD.n2377 VDD.t185 1.4705
R30535 VDD.n2377 VDD.t233 1.4705
R30536 VDD.n6995 VDD.t204 1.4705
R30537 VDD.n6995 VDD.t253 1.4705
R30538 VDD.n6990 VDD.t202 1.4705
R30539 VDD.n6990 VDD.t128 1.4705
R30540 VDD.n6985 VDD.t215 1.4705
R30541 VDD.n6985 VDD.t286 1.4705
R30542 VDD.n6980 VDD.t53 1.4705
R30543 VDD.n6980 VDD.t139 1.4705
R30544 VDD.n6898 VDD.t196 1.4705
R30545 VDD.n6898 VDD.t271 1.4705
R30546 VDD.n6893 VDD.t276 1.4705
R30547 VDD.n6893 VDD.t151 1.4705
R30548 VDD.n6888 VDD.t287 1.4705
R30549 VDD.n6888 VDD.t135 1.4705
R30550 VDD.n6886 VDD.t167 1.4705
R30551 VDD.n6886 VDD.t219 1.4705
R30552 VDD.n6967 VDD.t126 1.4705
R30553 VDD.n6967 VDD.t173 1.4705
R30554 VDD.n6969 VDD.t124 1.4705
R30555 VDD.n6969 VDD.t275 1.4705
R30556 VDD.n6971 VDD.t138 1.4705
R30557 VDD.n6971 VDD.t211 1.4705
R30558 VDD.n6973 VDD.t222 1.4705
R30559 VDD.n6973 VDD.t284 1.4705
R30560 VDD.n6965 VDD.t119 1.4705
R30561 VDD.n6965 VDD.t194 1.4705
R30562 VDD.n6963 VDD.t203 1.4705
R30563 VDD.n6963 VDD.t57 1.4705
R30564 VDD.n6961 VDD.t216 1.4705
R30565 VDD.n6961 VDD.t279 1.4705
R30566 VDD.n6960 VDD.t86 1.4705
R30567 VDD.n6960 VDD.t141 1.4705
R30568 VDD.n6947 VDD.t266 1.4705
R30569 VDD.n6947 VDD.t88 1.4705
R30570 VDD.n6942 VDD.t265 1.4705
R30571 VDD.n6942 VDD.t190 1.4705
R30572 VDD.n6937 VDD.t277 1.4705
R30573 VDD.n6937 VDD.t130 1.4705
R30574 VDD.n6932 VDD.t136 1.4705
R30575 VDD.n6932 VDD.t207 1.4705
R30576 VDD.n6917 VDD.t264 1.4705
R30577 VDD.n6917 VDD.t111 1.4705
R30578 VDD.n6912 VDD.t116 1.4705
R30579 VDD.n6912 VDD.t213 1.4705
R30580 VDD.n6907 VDD.t132 1.4705
R30581 VDD.n6907 VDD.t201 1.4705
R30582 VDD.n6905 VDD.t232 1.4705
R30583 VDD.n6905 VDD.t278 1.4705
R30584 VDD.n7006 VDD.t120 1.4705
R30585 VDD.n7006 VDD.t198 1.4705
R30586 VDD.n7007 VDD.t288 1.4705
R30587 VDD.n7007 VDD.t144 1.4705
R30588 VDD.n7000 VDD.t145 1.4705
R30589 VDD.n7000 VDD.t220 1.4705
R30590 VDD.n7001 VDD.t82 1.4705
R30591 VDD.n7001 VDD.t162 1.4705
R30592 VDD.t4059 VDD.n5238 1.4705
R30593 VDD.n5238 VDD.t2764 1.4705
R30594 VDD.n5239 VDD.t811 1.4705
R30595 VDD.n5239 VDD.t4059 1.4705
R30596 VDD.t2638 VDD.n5243 1.4705
R30597 VDD.n5243 VDD.t811 1.4705
R30598 VDD.n5246 VDD.t4341 1.4705
R30599 VDD.n5246 VDD.t2042 1.4705
R30600 VDD.t1534 VDD.n5251 1.4705
R30601 VDD.n5251 VDD.t4341 1.4705
R30602 VDD.t2392 VDD.n5256 1.4705
R30603 VDD.n5256 VDD.t1048 1.4705
R30604 VDD.n5257 VDD.t3692 1.4705
R30605 VDD.n5257 VDD.t2392 1.4705
R30606 VDD.t4573 VDD.n5261 1.4705
R30607 VDD.n5261 VDD.t3692 1.4705
R30608 VDD.n5235 VDD.t1949 1.4705
R30609 VDD.n5235 VDD.t4727 1.4705
R30610 VDD.n5233 VDD.t2957 1.4705
R30611 VDD.t1949 VDD.n5233 1.4705
R30612 VDD.n5232 VDD.t4579 1.4705
R30613 VDD.t2957 VDD.n5232 1.4705
R30614 VDD.n5229 VDD.t2281 1.4705
R30615 VDD.t4103 VDD.n5229 1.4705
R30616 VDD.n5228 VDD.t3623 1.4705
R30617 VDD.t2281 VDD.n5228 1.4705
R30618 VDD.n5226 VDD.t4365 1.4705
R30619 VDD.t3163 VDD.n5226 1.4705
R30620 VDD.n5224 VDD.t1577 1.4705
R30621 VDD.t4365 VDD.n5224 1.4705
R30622 VDD.n5223 VDD.t2594 1.4705
R30623 VDD.t1577 VDD.n5223 1.4705
R30624 VDD.n6359 VDD.t570 1.4705
R30625 VDD.t4419 VDD.n6359 1.4705
R30626 VDD.n6354 VDD.t1988 1.4705
R30627 VDD.n6354 VDD.t570 1.4705
R30628 VDD.n6353 VDD.t4301 1.4705
R30629 VDD.t1988 VDD.n6353 1.4705
R30630 VDD.n6348 VDD.t1936 1.4705
R30631 VDD.t3789 VDD.n6348 1.4705
R30632 VDD.n6343 VDD.t2337 1.4705
R30633 VDD.n6343 VDD.t1936 1.4705
R30634 VDD.n6340 VDD.t4089 1.4705
R30635 VDD.t3231 VDD.n6340 1.4705
R30636 VDD.n6335 VDD.t1275 1.4705
R30637 VDD.n6335 VDD.t4089 1.4705
R30638 VDD.n6334 VDD.t4097 1.4705
R30639 VDD.t1275 VDD.n6334 1.4705
R30640 VDD.n6357 VDD.t3661 1.4705
R30641 VDD.n6357 VDD.t3339 1.4705
R30642 VDD.n6356 VDD.t918 1.4705
R30643 VDD.t3661 VDD.n6356 1.4705
R30644 VDD.n6351 VDD.t3265 1.4705
R30645 VDD.n6351 VDD.t918 1.4705
R30646 VDD.n6346 VDD.t876 1.4705
R30647 VDD.n6346 VDD.t2788 1.4705
R30648 VDD.n6345 VDD.t1170 1.4705
R30649 VDD.t876 VDD.n6345 1.4705
R30650 VDD.n6338 VDD.t3053 1.4705
R30651 VDD.n6338 VDD.t2089 1.4705
R30652 VDD.n6337 VDD.t4351 1.4705
R30653 VDD.t3053 VDD.n6337 1.4705
R30654 VDD.n6332 VDD.t3057 1.4705
R30655 VDD.n6332 VDD.t4351 1.4705
R30656 VDD.t2040 VDD.n5448 1.4705
R30657 VDD.n5448 VDD.t632 1.4705
R30658 VDD.n5449 VDD.t3019 1.4705
R30659 VDD.n5449 VDD.t2040 1.4705
R30660 VDD.t4669 VDD.n5453 1.4705
R30661 VDD.n5453 VDD.t3019 1.4705
R30662 VDD.n5456 VDD.t2390 1.4705
R30663 VDD.n5456 VDD.t4177 1.4705
R30664 VDD.t3690 VDD.n5461 1.4705
R30665 VDD.n5461 VDD.t2390 1.4705
R30666 VDD.t4439 VDD.n5466 1.4705
R30667 VDD.n5466 VDD.t4543 1.4705
R30668 VDD.n5467 VDD.t1653 1.4705
R30669 VDD.n5467 VDD.t4439 1.4705
R30670 VDD.t3995 VDD.n5471 1.4705
R30671 VDD.n5471 VDD.t1653 1.4705
R30672 VDD.n5392 VDD.t952 1.4705
R30673 VDD.t3702 VDD.n5392 1.4705
R30674 VDD.n5390 VDD.t1812 1.4705
R30675 VDD.t952 VDD.n5390 1.4705
R30676 VDD.n5389 VDD.t3584 1.4705
R30677 VDD.t1812 VDD.n5389 1.4705
R30678 VDD.n5386 VDD.t1196 1.4705
R30679 VDD.t3123 VDD.n5386 1.4705
R30680 VDD.n5385 VDD.t2680 1.4705
R30681 VDD.t1196 VDD.n5385 1.4705
R30682 VDD.n5383 VDD.t3360 1.4705
R30683 VDD.t3501 VDD.n5383 1.4705
R30684 VDD.n5381 VDD.t4715 1.4705
R30685 VDD.t3360 VDD.n5381 1.4705
R30686 VDD.n5380 VDD.t2973 1.4705
R30687 VDD.t4715 VDD.n5380 1.4705
R30688 VDD.n6592 VDD.t3759 1.4705
R30689 VDD.t2461 VDD.n6592 1.4705
R30690 VDD.n6588 VDD.t4649 1.4705
R30691 VDD.n6588 VDD.t3759 1.4705
R30692 VDD.n6587 VDD.t2285 1.4705
R30693 VDD.t4649 VDD.n6587 1.4705
R30694 VDD.n6582 VDD.t4053 1.4705
R30695 VDD.t1702 VDD.n6582 1.4705
R30696 VDD.t1246 VDD.n5925 1.4705
R30697 VDD.n5925 VDD.t4053 1.4705
R30698 VDD.t2030 VDD.n5930 1.4705
R30699 VDD.n5930 VDD.t2175 1.4705
R30700 VDD.n5931 VDD.t3414 1.4705
R30701 VDD.n5931 VDD.t2030 1.4705
R30702 VDD.t1530 VDD.n5935 1.4705
R30703 VDD.n5935 VDD.t3414 1.4705
R30704 VDD.t1118 VDD.n6236 1.4705
R30705 VDD.n6236 VDD.t3901 1.4705
R30706 VDD.n6237 VDD.t2038 1.4705
R30707 VDD.n6237 VDD.t1118 1.4705
R30708 VDD.t3771 VDD.n6241 1.4705
R30709 VDD.n6241 VDD.t2038 1.4705
R30710 VDD.n6244 VDD.t1392 1.4705
R30711 VDD.n6244 VDD.t3293 1.4705
R30712 VDD.t2867 VDD.n6249 1.4705
R30713 VDD.n6249 VDD.t1392 1.4705
R30714 VDD.t3541 VDD.n6254 1.4705
R30715 VDD.n6254 VDD.t3665 1.4705
R30716 VDD.n6255 VDD.t777 1.4705
R30717 VDD.n6255 VDD.t3541 1.4705
R30718 VDD.t3143 VDD.n6259 1.4705
R30719 VDD.n6259 VDD.t777 1.4705
R30720 VDD.t3863 VDD.n6272 1.4705
R30721 VDD.n6272 VDD.t3535 1.4705
R30722 VDD.n6273 VDD.t1087 1.4705
R30723 VDD.n6273 VDD.t3863 1.4705
R30724 VDD.t3412 VDD.n6277 1.4705
R30725 VDD.n6277 VDD.t1087 1.4705
R30726 VDD.n6280 VDD.t1041 1.4705
R30727 VDD.n6280 VDD.t2965 1.4705
R30728 VDD.t1350 VDD.n6285 1.4705
R30729 VDD.n6285 VDD.t1041 1.4705
R30730 VDD.t3229 VDD.n6290 1.4705
R30731 VDD.n6290 VDD.t2312 1.4705
R30732 VDD.n6291 VDD.t4521 1.4705
R30733 VDD.n6291 VDD.t3229 1.4705
R30734 VDD.t3235 VDD.n6295 1.4705
R30735 VDD.n6295 VDD.t4521 1.4705
R30736 VDD.n6233 VDD.t1128 1.4705
R30737 VDD.n6233 VDD.t3919 1.4705
R30738 VDD.n6231 VDD.t2059 1.4705
R30739 VDD.t1128 VDD.n6231 1.4705
R30740 VDD.n6230 VDD.t3787 1.4705
R30741 VDD.t2059 VDD.n6230 1.4705
R30742 VDD.n6227 VDD.t1404 1.4705
R30743 VDD.t3301 VDD.n6227 1.4705
R30744 VDD.n6226 VDD.t2879 1.4705
R30745 VDD.t1404 VDD.n6226 1.4705
R30746 VDD.n6224 VDD.t3553 1.4705
R30747 VDD.t3684 VDD.n6224 1.4705
R30748 VDD.n6222 VDD.t788 1.4705
R30749 VDD.t3553 VDD.n6222 1.4705
R30750 VDD.n6221 VDD.t3157 1.4705
R30751 VDD.t788 VDD.n6221 1.4705
R30752 VDD.n6214 VDD.t3877 1.4705
R30753 VDD.t3545 VDD.n6214 1.4705
R30754 VDD.n6212 VDD.t1105 1.4705
R30755 VDD.t3877 VDD.n6212 1.4705
R30756 VDD.n6211 VDD.t3433 1.4705
R30757 VDD.t1105 VDD.n6211 1.4705
R30758 VDD.n6208 VDD.t1066 1.4705
R30759 VDD.t2981 VDD.n6208 1.4705
R30760 VDD.n6207 VDD.t1366 1.4705
R30761 VDD.t1066 VDD.n6207 1.4705
R30762 VDD.n6205 VDD.t3243 1.4705
R30763 VDD.t2335 VDD.n6205 1.4705
R30764 VDD.n6203 VDD.t4527 1.4705
R30765 VDD.t3243 VDD.n6203 1.4705
R30766 VDD.n6202 VDD.t3249 1.4705
R30767 VDD.t4527 VDD.n6202 1.4705
R30768 VDD.t2419 VDD.n5954 1.4705
R30769 VDD.n5954 VDD.t2011 1.4705
R30770 VDD.n5955 VDD.t3722 1.4705
R30771 VDD.n5955 VDD.t2419 1.4705
R30772 VDD.t1865 VDD.n5959 1.4705
R30773 VDD.n5959 VDD.t3722 1.4705
R30774 VDD.n5962 VDD.t3675 1.4705
R30775 VDD.n5962 VDD.t1339 1.4705
R30776 VDD.t4025 VDD.n5967 1.4705
R30777 VDD.n5967 VDD.t3675 1.4705
R30778 VDD.t1638 VDD.n5972 1.4705
R30779 VDD.n5972 VDD.t765 1.4705
R30780 VDD.n5973 VDD.t3099 1.4705
R30781 VDD.n5973 VDD.t1638 1.4705
R30782 VDD.t1647 VDD.n5977 1.4705
R30783 VDD.n5977 VDD.t3099 1.4705
R30784 VDD.t931 VDD.n6383 1.4705
R30785 VDD.n6383 VDD.t4721 1.4705
R30786 VDD.n6384 VDD.t2343 1.4705
R30787 VDD.n6384 VDD.t931 1.4705
R30788 VDD.t4571 VDD.n6388 1.4705
R30789 VDD.n6388 VDD.t2343 1.4705
R30790 VDD.n6391 VDD.t2273 1.4705
R30791 VDD.n6391 VDD.t4095 1.4705
R30792 VDD.t2662 VDD.n5996 1.4705
R30793 VDD.n5996 VDD.t2273 1.4705
R30794 VDD.t4363 VDD.n6001 1.4705
R30795 VDD.n6001 VDD.t3483 1.4705
R30796 VDD.n6002 VDD.t1568 1.4705
R30797 VDD.n6002 VDD.t4363 1.4705
R30798 VDD.t4369 VDD.n6006 1.4705
R30799 VDD.n6006 VDD.t1568 1.4705
R30800 VDD.n5320 VDD.t3045 1.4705
R30801 VDD.t2719 VDD.n5320 1.4705
R30802 VDD.n5318 VDD.t4343 1.4705
R30803 VDD.t3045 VDD.n5318 1.4705
R30804 VDD.n5317 VDD.t2592 1.4705
R30805 VDD.t4343 VDD.n5317 1.4705
R30806 VDD.t4297 VDD.n5314 1.4705
R30807 VDD.t1980 VDD.n5314 1.4705
R30808 VDD.t4615 VDD.n5994 1.4705
R30809 VDD.n5994 VDD.t4297 1.4705
R30810 VDD.n5993 VDD.t2331 1.4705
R30811 VDD.t1346 VDD.n5993 1.4705
R30812 VDD.n5991 VDD.t3641 1.4705
R30813 VDD.t2331 VDD.n5991 1.4705
R30814 VDD.n5990 VDD.t2341 1.4705
R30815 VDD.t3641 VDD.n5990 1.4705
R30816 VDD.t2396 VDD.n5337 1.4705
R30817 VDD.n5337 VDD.t963 1.4705
R30818 VDD.n5338 VDD.t3279 1.4705
R30819 VDD.n5338 VDD.t2396 1.4705
R30820 VDD.t824 VDD.n5342 1.4705
R30821 VDD.n5342 VDD.t3279 1.4705
R30822 VDD.n5345 VDD.t2697 1.4705
R30823 VDD.n5345 VDD.t4443 1.4705
R30824 VDD.t3999 VDD.n5350 1.4705
R30825 VDD.n5350 VDD.t2697 1.4705
R30826 VDD.t4733 VDD.n5355 1.4705
R30827 VDD.n5355 VDD.t717 1.4705
R30828 VDD.n5356 VDD.t1962 1.4705
R30829 VDD.n5356 VDD.t4733 1.4705
R30830 VDD.t4279 VDD.n5360 1.4705
R30831 VDD.n5360 VDD.t1962 1.4705
R30832 VDD.n5334 VDD.t4371 1.4705
R30833 VDD.n5334 VDD.t3079 1.4705
R30834 VDD.n5332 VDD.t1126 1.4705
R30835 VDD.t4371 VDD.n5332 1.4705
R30836 VDD.n5331 VDD.t2963 1.4705
R30837 VDD.t1126 VDD.n5331 1.4705
R30838 VDD.n5328 VDD.t4663 1.4705
R30839 VDD.t2434 VDD.n5328 1.4705
R30840 VDD.n5327 VDD.t1874 1.4705
R30841 VDD.t4663 VDD.n5327 1.4705
R30842 VDD.n5325 VDD.t2738 1.4705
R30843 VDD.t2863 VDD.n5325 1.4705
R30844 VDD.n5323 VDD.t4041 1.4705
R30845 VDD.t2738 VDD.n5323 1.4705
R30846 VDD.n5322 VDD.t2204 1.4705
R30847 VDD.t4041 VDD.n5322 1.4705
R30848 VDD.n6411 VDD.t1420 1.4705
R30849 VDD.t1111 VDD.n6411 1.4705
R30850 VDD.n6407 VDD.t2901 1.4705
R30851 VDD.n6407 VDD.t1420 1.4705
R30852 VDD.n6406 VDD.t1006 1.4705
R30853 VDD.t2901 VDD.n6406 1.4705
R30854 VDD.n6401 VDD.t2861 1.4705
R30855 VDD.t4597 VDD.n6401 1.4705
R30856 VDD.t3171 VDD.n6160 1.4705
R30857 VDD.n6160 VDD.t2861 1.4705
R30858 VDD.t771 VDD.n6165 1.4705
R30859 VDD.n6165 VDD.t4015 1.4705
R30860 VDD.n6166 VDD.t2136 1.4705
R30861 VDD.n6166 VDD.t771 1.4705
R30862 VDD.t779 VDD.n6170 1.4705
R30863 VDD.n6170 VDD.t2136 1.4705
R30864 VDD.t2949 VDD.n6564 1.4705
R30865 VDD.n6564 VDD.t1454 1.4705
R30866 VDD.n6565 VDD.t3769 1.4705
R30867 VDD.n6565 VDD.t2949 1.4705
R30868 VDD.t1321 VDD.n6569 1.4705
R30869 VDD.n6569 VDD.t3769 1.4705
R30870 VDD.n6572 VDD.t3211 1.4705
R30871 VDD.n6572 VDD.t853 1.4705
R30872 VDD.t4501 VDD.n6027 1.4705
R30873 VDD.n6027 VDD.t3211 1.4705
R30874 VDD.n6030 VDD.t1122 1.4705
R30875 VDD.n6030 VDD.t1234 1.4705
R30876 VDD.t2584 VDD.n6034 1.4705
R30877 VDD.n6034 VDD.t1122 1.4705
R30878 VDD.n6035 VDD.t650 1.4705
R30879 VDD.n6035 VDD.t2584 1.4705
R30880 VDD.n6498 VDD.t4923 1.4705
R30881 VDD.n6498 VDD.t4858 1.4705
R30882 VDD.n6499 VDD.t4834 1.4705
R30883 VDD.n6499 VDD.t4964 1.4705
R30884 VDD.n6448 VDD.t4856 1.4705
R30885 VDD.n6448 VDD.t4840 1.4705
R30886 VDD.n6449 VDD.t4963 1.4705
R30887 VDD.n6449 VDD.t4947 1.4705
R30888 VDD.n6558 VDD.t4978 1.4705
R30889 VDD.n6558 VDD.t4915 1.4705
R30890 VDD.n6556 VDD.t4909 1.4705
R30891 VDD.n6556 VDD.t4827 1.4705
R30892 VDD.n6554 VDD.t4900 1.4705
R30893 VDD.n6554 VDD.t4905 1.4705
R30894 VDD.n6552 VDD.t4875 1.4705
R30895 VDD.n6552 VDD.t4961 1.4705
R30896 VDD.n5295 VDD.t4914 1.4705
R30897 VDD.n5295 VDD.t4898 1.4705
R30898 VDD.n5293 VDD.t4892 1.4705
R30899 VDD.n5293 VDD.t4974 1.4705
R30900 VDD.n5291 VDD.t4881 1.4705
R30901 VDD.n5291 VDD.t4833 1.4705
R30902 VDD.n5290 VDD.t4882 1.4705
R30903 VDD.n5290 VDD.t4941 1.4705
R30904 VDD.n6445 VDD.t4812 1.4705
R30905 VDD.n6445 VDD.t4927 1.4705
R30906 VDD.n6442 VDD.t4922 1.4705
R30907 VDD.n6442 VDD.t4837 1.4705
R30908 VDD.n6439 VDD.t4913 1.4705
R30909 VDD.n6439 VDD.t4918 1.4705
R30910 VDD.n6436 VDD.t4891 1.4705
R30911 VDD.n6436 VDD.t4973 1.4705
R30912 VDD.n6431 VDD.t4924 1.4705
R30913 VDD.n6431 VDD.t4910 1.4705
R30914 VDD.n6426 VDD.t4906 1.4705
R30915 VDD.n6426 VDD.t4809 1.4705
R30916 VDD.n6421 VDD.t4895 1.4705
R30917 VDD.n6421 VDD.t4848 1.4705
R30918 VDD.n6419 VDD.t4896 1.4705
R30919 VDD.n6419 VDD.t4954 1.4705
R30920 VDD.n6519 VDD.t4864 1.4705
R30921 VDD.n6519 VDD.t4814 1.4705
R30922 VDD.n6517 VDD.t4981 1.4705
R30923 VDD.n6517 VDD.t4907 1.4705
R30924 VDD.n6515 VDD.t4977 1.4705
R30925 VDD.n6515 VDD.t4980 1.4705
R30926 VDD.n6513 VDD.t4952 1.4705
R30927 VDD.n6513 VDD.t4844 1.4705
R30928 VDD.n6510 VDD.t4811 1.4705
R30929 VDD.n6510 VDD.t4975 1.4705
R30930 VDD.n6508 VDD.t4966 1.4705
R30931 VDD.n6508 VDD.t4862 1.4705
R30932 VDD.n6506 VDD.t4957 1.4705
R30933 VDD.n6506 VDD.t4917 1.4705
R30934 VDD.n6505 VDD.t4958 1.4705
R30935 VDD.n6505 VDD.t4830 1.4705
R30936 VDD.n6482 VDD.t4933 1.4705
R30937 VDD.n6482 VDD.t4872 1.4705
R30938 VDD.n6479 VDD.t4867 1.4705
R30939 VDD.n6479 VDD.t4979 1.4705
R30940 VDD.n6476 VDD.t4852 1.4705
R30941 VDD.n6476 VDD.t4860 1.4705
R30942 VDD.n6473 VDD.t4832 1.4705
R30943 VDD.n6473 VDD.t4920 1.4705
R30944 VDD.n6468 VDD.t4870 1.4705
R30945 VDD.n6468 VDD.t4849 1.4705
R30946 VDD.n6463 VDD.t4845 1.4705
R30947 VDD.n6463 VDD.t4931 1.4705
R30948 VDD.n6458 VDD.t4835 1.4705
R30949 VDD.n6458 VDD.t4808 1.4705
R30950 VDD.n6456 VDD.t4836 1.4705
R30951 VDD.n6456 VDD.t4904 1.4705
R30952 VDD.n6544 VDD.t4841 1.4705
R30953 VDD.n6544 VDD.t4970 1.4705
R30954 VDD.n6545 VDD.t4894 1.4705
R30955 VDD.n6545 VDD.t4829 1.4705
R30956 VDD.n6537 VDD.t4968 1.4705
R30957 VDD.n6537 VDD.t4953 1.4705
R30958 VDD.n6538 VDD.t4828 1.4705
R30959 VDD.n6538 VDD.t4818 1.4705
R30960 VDD.n6069 VDD.t4948 1.4705
R30961 VDD.n6069 VDD.t4839 1.4705
R30962 VDD.n6063 VDD.t4930 1.4705
R30963 VDD.n6063 VDD.t4826 1.4705
R30964 VDD.n6134 VDD.t4960 1.4705
R30965 VDD.n6134 VDD.t4899 1.4705
R30966 VDD.n6135 VDD.t4823 1.4705
R30967 VDD.n6135 VDD.t4943 1.4705
R30968 VDD.n6137 VDD.t4893 1.4705
R30969 VDD.n6137 VDD.t4816 1.4705
R30970 VDD.n6138 VDD.t4936 1.4705
R30971 VDD.n6138 VDD.t4853 1.4705
R30972 VDD.n6141 VDD.t4883 1.4705
R30973 VDD.n6141 VDD.t4887 1.4705
R30974 VDD.n6142 VDD.t4928 1.4705
R30975 VDD.n6142 VDD.t4932 1.4705
R30976 VDD.n6145 VDD.t4854 1.4705
R30977 VDD.n6145 VDD.t4942 1.4705
R30978 VDD.n6146 VDD.t4908 1.4705
R30979 VDD.n6146 VDD.t4813 1.4705
R30980 VDD.n6130 VDD.t4897 1.4705
R30981 VDD.n6130 VDD.t4880 1.4705
R30982 VDD.n6131 VDD.t4939 1.4705
R30983 VDD.n6131 VDD.t4926 1.4705
R30984 VDD.n6126 VDD.t4874 1.4705
R30985 VDD.n6126 VDD.t4955 1.4705
R30986 VDD.n6127 VDD.t4921 1.4705
R30987 VDD.n6127 VDD.t4822 1.4705
R30988 VDD.n6122 VDD.t4861 1.4705
R30989 VDD.n6122 VDD.t4824 1.4705
R30990 VDD.n6123 VDD.t4911 1.4705
R30991 VDD.n6123 VDD.t4869 1.4705
R30992 VDD.n6118 VDD.t4863 1.4705
R30993 VDD.n6118 VDD.t4925 1.4705
R30994 VDD.n6119 VDD.t4912 1.4705
R30995 VDD.n6119 VDD.t4971 1.4705
R30996 VDD.n6042 VDD.t4843 1.4705
R30997 VDD.n6042 VDD.t4976 1.4705
R30998 VDD.n6043 VDD.t4950 1.4705
R30999 VDD.n6043 VDD.t4889 1.4705
R31000 VDD.n6045 VDD.t4967 1.4705
R31001 VDD.n6045 VDD.t4890 1.4705
R31002 VDD.n6046 VDD.t4885 1.4705
R31003 VDD.n6046 VDD.t4815 1.4705
R31004 VDD.n6049 VDD.t4959 1.4705
R31005 VDD.n6049 VDD.t4965 1.4705
R31006 VDD.n6050 VDD.t4873 1.4705
R31007 VDD.n6050 VDD.t4879 1.4705
R31008 VDD.n6053 VDD.t4935 1.4705
R31009 VDD.n6053 VDD.t4831 1.4705
R31010 VDD.n6054 VDD.t4847 1.4705
R31011 VDD.n6054 VDD.t4934 1.4705
R31012 VDD.n6076 VDD.t4972 1.4705
R31013 VDD.n6076 VDD.t4956 1.4705
R31014 VDD.n6077 VDD.t4888 1.4705
R31015 VDD.n6077 VDD.t4871 1.4705
R31016 VDD.n6080 VDD.t4951 1.4705
R31017 VDD.n6080 VDD.t4842 1.4705
R31018 VDD.n6081 VDD.t4865 1.4705
R31019 VDD.n6081 VDD.t4949 1.4705
R31020 VDD.n6084 VDD.t4938 1.4705
R31021 VDD.n6084 VDD.t4903 1.4705
R31022 VDD.n6085 VDD.t4850 1.4705
R31023 VDD.n6085 VDD.t4820 1.4705
R31024 VDD.n6088 VDD.t4940 1.4705
R31025 VDD.n6088 VDD.t4821 1.4705
R31026 VDD.n6089 VDD.t4851 1.4705
R31027 VDD.n6089 VDD.t4919 1.4705
R31028 VDD.n6020 VDD.t4859 1.4705
R31029 VDD.n6020 VDD.t4810 1.4705
R31030 VDD.n6154 VDD.t4983 1.4705
R31031 VDD.n6154 VDD.t4969 1.4705
R31032 VDD.n6112 VDD.t4819 1.4705
R31033 VDD.n6112 VDD.t4902 1.4705
R31034 VDD.n6106 VDD.t4982 1.4705
R31035 VDD.n6106 VDD.t4884 1.4705
R31036 VDD.n6093 VDD.t4937 1.4705
R31037 VDD.n6093 VDD.t4878 1.4705
R31038 VDD.n6097 VDD.t4876 1.4705
R31039 VDD.n6097 VDD.t4857 1.4705
R31040 VDD.t2695 VDD.n7847 1.4705
R31041 VDD.n7847 VDD.t1205 1.4705
R31042 VDD.n7848 VDD.t1217 1.4705
R31043 VDD.n7848 VDD.t2695 1.4705
R31044 VDD.n2226 VDD.t1994 1.4705
R31045 VDD.t4387 VDD.n2226 1.4705
R31046 VDD.n2225 VDD.t3380 1.4705
R31047 VDD.t1994 VDD.n2225 1.4705
R31048 VDD.t1021 VDD.n7990 1.4705
R31049 VDD.n7990 VDD.t3793 1.4705
R31050 VDD.n7991 VDD.t2474 1.4705
R31051 VDD.n7991 VDD.t1021 1.4705
R31052 VDD.n7981 VDD.t3647 1.4705
R31053 VDD.n7981 VDD.t2474 1.4705
R31054 VDD.n7964 VDD.t1307 1.4705
R31055 VDD.t4133 VDD.n7964 1.4705
R31056 VDD.t1694 VDD.n2229 1.4705
R31057 VDD.n2229 VDD.t4481 1.4705
R31058 VDD.n2230 VDD.t3063 1.4705
R31059 VDD.n2230 VDD.t1694 1.4705
R31060 VDD.n2222 VDD.t4361 1.4705
R31061 VDD.n2222 VDD.t3063 1.4705
R31062 VDD.n7985 VDD.t2009 1.4705
R31063 VDD.t1109 VDD.n7985 1.4705
R31064 VDD.n7984 VDD.t3402 1.4705
R31065 VDD.t2009 VDD.n7984 1.4705
R31066 VDD.n7978 VDD.t2442 1.4705
R31067 VDD.t1432 VDD.n7978 1.4705
R31068 VDD.n7972 VDD.t1014 1.4705
R31069 VDD.n7972 VDD.t2442 1.4705
R31070 VDD.n7971 VDD.t1884 1.4705
R31071 VDD.t1014 VDD.n7971 1.4705
R31072 VDD.n6600 VDD.t2269 1.4705
R31073 VDD.n6600 VDD.t1307 1.4705
R31074 VDD.t3991 VDD.n6604 1.4705
R31075 VDD.n6604 VDD.t2269 1.4705
R31076 VDD.n6607 VDD.t1605 1.4705
R31077 VDD.n6607 VDD.t3481 1.4705
R31078 VDD.t3073 VDD.n6612 1.4705
R31079 VDD.n6612 VDD.t1605 1.4705
R31080 VDD.t3755 VDD.n6617 1.4705
R31081 VDD.n6617 VDD.t2566 1.4705
R31082 VDD.n6618 VDD.t1002 1.4705
R31083 VDD.n6618 VDD.t3755 1.4705
R31084 VDD.t1867 VDD.n6622 1.4705
R31085 VDD.n6622 VDD.t1002 1.4705
R31086 VDD.t3763 VDD.n5409 1.4705
R31087 VDD.n5409 VDD.t2463 1.4705
R31088 VDD.n5410 VDD.t4651 1.4705
R31089 VDD.n5410 VDD.t3763 1.4705
R31090 VDD.t2287 VDD.n5414 1.4705
R31091 VDD.n5414 VDD.t4651 1.4705
R31092 VDD.n5417 VDD.t4055 1.4705
R31093 VDD.n5417 VDD.t1704 1.4705
R31094 VDD.t1248 VDD.n5422 1.4705
R31095 VDD.n5422 VDD.t4055 1.4705
R31096 VDD.t2032 VDD.n5427 1.4705
R31097 VDD.n5427 VDD.t769 1.4705
R31098 VDD.n5428 VDD.t3418 1.4705
R31099 VDD.n5428 VDD.t2032 1.4705
R31100 VDD.t4303 VDD.n5432 1.4705
R31101 VDD.n5432 VDD.t3418 1.4705
R31102 VDD.n5406 VDD.t2752 1.4705
R31103 VDD.n5406 VDD.t1261 1.4705
R31104 VDD.n5404 VDD.t3576 1.4705
R31105 VDD.t2752 VDD.n5404 1.4705
R31106 VDD.n5403 VDD.t1137 1.4705
R31107 VDD.t3576 VDD.n5403 1.4705
R31108 VDD.n5400 VDD.t3027 1.4705
R31109 VDD.t605 VDD.n5400 1.4705
R31110 VDD.n5399 VDD.t4319 1.4705
R31111 VDD.t3027 VDD.n5399 1.4705
R31112 VDD.n5397 VDD.t950 1.4705
R31113 VDD.t3809 VDD.n5397 1.4705
R31114 VDD.n5395 VDD.t2373 1.4705
R31115 VDD.t950 VDD.n5395 1.4705
R31116 VDD.n5394 VDD.t3263 1.4705
R31117 VDD.t2373 VDD.n5394 1.4705
R31118 VDD.n7171 VDD.t3645 1.4705
R31119 VDD.t2835 VDD.n7171 1.4705
R31120 VDD.n7166 VDD.t911 1.4705
R31121 VDD.n7166 VDD.t3645 1.4705
R31122 VDD.n7165 VDD.t3653 1.4705
R31123 VDD.t911 VDD.n7165 1.4705
R31124 VDD.n7160 VDD.t4399 1.4705
R31125 VDD.t2762 VDD.n7160 1.4705
R31126 VDD.n7155 VDD.t1622 1.4705
R31127 VDD.n7155 VDD.t4399 1.4705
R31128 VDD.n7152 VDD.t3455 1.4705
R31129 VDD.t2077 VDD.n7152 1.4705
R31130 VDD.n7147 VDD.t645 1.4705
R31131 VDD.n7147 VDD.t3455 1.4705
R31132 VDD.n7146 VDD.t1917 1.4705
R31133 VDD.t645 VDD.n7146 1.4705
R31134 VDD.n7169 VDD.t2644 1.4705
R31135 VDD.n7169 VDD.t1636 1.4705
R31136 VDD.n7168 VDD.t3951 1.4705
R31137 VDD.t2644 VDD.n7168 1.4705
R31138 VDD.n7163 VDD.t2656 1.4705
R31139 VDD.n7163 VDD.t3951 1.4705
R31140 VDD.n7158 VDD.t3333 1.4705
R31141 VDD.n7158 VDD.t1549 1.4705
R31142 VDD.n7157 VDD.t4689 1.4705
R31143 VDD.t3333 VDD.n7157 1.4705
R31144 VDD.n7150 VDD.t2415 1.4705
R31145 VDD.n7150 VDD.t989 1.4705
R31146 VDD.n7149 VDD.t3714 1.4705
R31147 VDD.t2415 VDD.n7149 1.4705
R31148 VDD.n7144 VDD.t851 1.4705
R31149 VDD.n7144 VDD.t3714 1.4705
R31150 VDD.t1205 VDD.n7846 1.4705
R31151 VDD.n7846 VDD.t4467 1.4705
R31152 VDD.n7948 VDD.t46 1.4705
R31153 VDD.n7948 VDD.t38 1.4705
R31154 VDD.n7950 VDD.t36 1.4705
R31155 VDD.n7950 VDD.t29 1.4705
R31156 VDD.n7953 VDD.t210 1.4705
R31157 VDD.n7953 VDD.t281 1.4705
R31158 VDD.n7955 VDD.t22 1.4705
R31159 VDD.n7955 VDD.t44 1.4705
R31160 VDD.n7957 VDD.t16 1.4705
R31161 VDD.n7957 VDD.t42 1.4705
R31162 VDD.n7938 VDD.t163 1.4705
R31163 VDD.n7938 VDD.t238 1.4705
R31164 VDD.n7933 VDD.t243 1.4705
R31165 VDD.n7933 VDD.t91 1.4705
R31166 VDD.n7928 VDD.t152 1.4705
R31167 VDD.n7928 VDD.t197 1.4705
R31168 VDD.n7919 VDD.t131 1.4705
R31169 VDD.n7919 VDD.t178 1.4705
R31170 VDD.n7914 VDD.t156 1.4705
R31171 VDD.n7914 VDD.t205 1.4705
R31172 VDD.n7884 VDD.t259 1.4705
R31173 VDD.n7884 VDD.t101 1.4705
R31174 VDD.n7886 VDD.t90 1.4705
R31175 VDD.n7886 VDD.t168 1.4705
R31176 VDD.n7880 VDD.t112 1.4705
R31177 VDD.n7880 VDD.t188 1.4705
R31178 VDD.n7882 VDD.t175 1.4705
R31179 VDD.n7882 VDD.t251 1.4705
R31180 VDD.n7876 VDD.t27 1.4705
R31181 VDD.n7876 VDD.t18 1.4705
R31182 VDD.n7878 VDD.t45 1.4705
R31183 VDD.n7878 VDD.t39 1.4705
R31184 VDD.n7870 VDD.t224 1.4705
R31185 VDD.n7870 VDD.t269 1.4705
R31186 VDD.n7872 VDD.t280 1.4705
R31187 VDD.n7872 VDD.t105 1.4705
R31188 VDD.n7866 VDD.t245 1.4705
R31189 VDD.n7866 VDD.t49 1.4705
R31190 VDD.n7868 VDD.t75 1.4705
R31191 VDD.n7868 VDD.t134 1.4705
R31192 VDD.n8053 VDD.t174 1.4705
R31193 VDD.n8053 VDD.t249 1.4705
R31194 VDD.n8055 VDD.t260 1.4705
R31195 VDD.n8055 VDD.t102 1.4705
R31196 VDD.n8058 VDD.t78 1.4705
R31197 VDD.n8058 VDD.t159 1.4705
R31198 VDD.n8060 VDD.t143 1.4705
R31199 VDD.n8060 VDD.t189 1.4705
R31200 VDD.n8062 VDD.t166 1.4705
R31201 VDD.n8062 VDD.t217 1.4705
R31202 VDD.n8043 VDD.t24 1.4705
R31203 VDD.n8043 VDD.t43 1.4705
R31204 VDD.n8038 VDD.t40 1.4705
R31205 VDD.n8038 VDD.t33 1.4705
R31206 VDD.n8033 VDD.t244 1.4705
R31207 VDD.n8033 VDD.t48 1.4705
R31208 VDD.n8024 VDD.t32 1.4705
R31209 VDD.n8024 VDD.t20 1.4705
R31210 VDD.n8019 VDD.t25 1.4705
R31211 VDD.n8019 VDD.t47 1.4705
R31212 VDD.t4109 VDD.n2176 1.4705
R31213 VDD.n2176 VDD.t2804 1.4705
R31214 VDD.n2177 VDD.t1189 1.4705
R31215 VDD.n2177 VDD.t4109 1.4705
R31216 VDD.t2672 VDD.n2181 1.4705
R31217 VDD.n2181 VDD.t1189 1.4705
R31218 VDD.n2184 VDD.t4375 1.4705
R31219 VDD.n2184 VDD.t3495 1.4705
R31220 VDD.t1587 VDD.n7999 1.4705
R31221 VDD.n7999 VDD.t4375 1.4705
R31222 VDD.t4729 VDD.n8004 1.4705
R31223 VDD.n8004 VDD.t3835 1.4705
R31224 VDD.n8005 VDD.t3378 1.4705
R31225 VDD.n8005 VDD.t4729 1.4705
R31226 VDD.t4277 VDD.n8009 1.4705
R31227 VDD.n8009 VDD.t3378 1.4705
R31228 VDD.n6808 VDD.t241 1.4705
R31229 VDD.n6808 VDD.t283 1.4705
R31230 VDD.n6809 VDD.t184 1.4705
R31231 VDD.n6809 VDD.t230 1.4705
R31232 VDD.n6811 VDD.t239 1.4705
R31233 VDD.n6811 VDD.t164 1.4705
R31234 VDD.n6812 VDD.t183 1.4705
R31235 VDD.n6812 VDD.t106 1.4705
R31236 VDD.n6815 VDD.t252 1.4705
R31237 VDD.n6815 VDD.t95 1.4705
R31238 VDD.n6816 VDD.t193 1.4705
R31239 VDD.n6816 VDD.t268 1.4705
R31240 VDD.n6819 VDD.t104 1.4705
R31241 VDD.n6819 VDD.t176 1.4705
R31242 VDD.n6820 VDD.t274 1.4705
R31243 VDD.n6820 VDD.t117 1.4705
R31244 VDD.n6824 VDD.t234 1.4705
R31245 VDD.n6824 VDD.t74 1.4705
R31246 VDD.n6825 VDD.t177 1.4705
R31247 VDD.n6825 VDD.t254 1.4705
R31248 VDD.n6828 VDD.t84 1.4705
R31249 VDD.n6828 VDD.t186 1.4705
R31250 VDD.n6829 VDD.t261 1.4705
R31251 VDD.n6829 VDD.t129 1.4705
R31252 VDD.n6832 VDD.t96 1.4705
R31253 VDD.n6832 VDD.t170 1.4705
R31254 VDD.n6833 VDD.t270 1.4705
R31255 VDD.n6833 VDD.t113 1.4705
R31256 VDD.n6836 VDD.t206 1.4705
R31257 VDD.n6836 VDD.t255 1.4705
R31258 VDD.n6837 VDD.t150 1.4705
R31259 VDD.n6837 VDD.t195 1.4705
R31260 VDD.n6775 VDD.t148 1.4705
R31261 VDD.n6775 VDD.t192 1.4705
R31262 VDD.n6776 VDD.t248 1.4705
R31263 VDD.n6776 VDD.t59 1.4705
R31264 VDD.n6778 VDD.t147 1.4705
R31265 VDD.n6778 VDD.t55 1.4705
R31266 VDD.n6779 VDD.t247 1.4705
R31267 VDD.n6779 VDD.t172 1.4705
R31268 VDD.n6782 VDD.t158 1.4705
R31269 VDD.n6782 VDD.t231 1.4705
R31270 VDD.n6783 VDD.t262 1.4705
R31271 VDD.n6783 VDD.t107 1.4705
R31272 VDD.n6786 VDD.t240 1.4705
R31273 VDD.n6786 VDD.t70 1.4705
R31274 VDD.n6787 VDD.t114 1.4705
R31275 VDD.n6787 VDD.t187 1.4705
R31276 VDD.n6771 VDD.t142 1.4705
R31277 VDD.n6771 VDD.t218 1.4705
R31278 VDD.n6772 VDD.t242 1.4705
R31279 VDD.n6772 VDD.t89 1.4705
R31280 VDD.n6767 VDD.t225 1.4705
R31281 VDD.n6767 VDD.t87 1.4705
R31282 VDD.n6768 VDD.t94 1.4705
R31283 VDD.n6768 VDD.t191 1.4705
R31284 VDD.n6763 VDD.t235 1.4705
R31285 VDD.n6763 VDD.t64 1.4705
R31286 VDD.n6764 VDD.t110 1.4705
R31287 VDD.n6764 VDD.t181 1.4705
R31288 VDD.n6759 VDD.t108 1.4705
R31289 VDD.n6759 VDD.t160 1.4705
R31290 VDD.n6760 VDD.t212 1.4705
R31291 VDD.n6760 VDD.t263 1.4705
R31292 VDD.n6845 VDD.t97 1.4705
R31293 VDD.n6845 VDD.t179 1.4705
R31294 VDD.n6842 VDD.t121 1.4705
R31295 VDD.n6842 VDD.t199 1.4705
R31296 VDD.n6736 VDD.t161 1.4705
R31297 VDD.n6736 VDD.t258 1.4705
R31298 VDD.n6732 VDD.t182 1.4705
R31299 VDD.n6732 VDD.t68 1.4705
R31300 VDD.n6795 VDD.t236 1.4705
R31301 VDD.n6795 VDD.t77 1.4705
R31302 VDD.n6792 VDD.t257 1.4705
R31303 VDD.n6792 VDD.t100 1.4705
R31304 VDD.n9131 VDD.t3323 1.4705
R31305 VDD.n9131 VDD.t3519 1.4705
R31306 VDD.t2796 VDD.n9129 1.4705
R31307 VDD.n9129 VDD.t3001 1.4705
R31308 VDD.t4043 VDD.n9142 1.4705
R31309 VDD.n9142 VDD.t2549 1.4705
R31310 VDD.t3673 VDD.n9148 1.4705
R31311 VDD.n9148 VDD.t3899 1.4705
R31312 VDD.n9165 VDD.t4569 1.4705
R31313 VDD.t3103 VDD.n9165 1.4705
R31314 VDD.t4257 VDD.n8487 1.4705
R31315 VDD.n8487 VDD.t4461 1.4705
R31316 VDD.n8762 VDD.t3841 1.4705
R31317 VDD.t4061 VDD.n8762 1.4705
R31318 VDD.n8756 VDD.t3861 1.4705
R31319 VDD.t4517 VDD.n8756 1.4705
R31320 VDD.n8558 VDD.t2024 1.4705
R31321 VDD.t2255 VDD.n8558 1.4705
R31322 VDD.n8552 VDD.t2062 1.4705
R31323 VDD.t2815 VDD.n8552 1.4705
R31324 VDD.n8835 VDD.t2112 1.4705
R31325 VDD.t2871 VDD.n8835 1.4705
R31326 VDD.t2134 VDD.n8546 1.4705
R31327 VDD.n8546 VDD.t1035 1.4705
R31328 VDD.t3935 VDD.n8802 1.4705
R31329 VDD.n8802 VDD.t4585 1.4705
R31330 VDD.n8768 VDD.t3959 1.4705
R31331 VDD.t2943 VDD.n8768 1.4705
R31332 VDD.n8888 VDD.t3447 1.4705
R31333 VDD.t2523 VDD.n8888 1.4705
R31334 VDD.t3471 VDD.n8774 1.4705
R31335 VDD.n8774 VDD.t2440 1.4705
R31336 VDD.t1593 VDD.n8875 1.4705
R31337 VDD.n8875 VDD.t581 1.4705
R31338 VDD.n8841 VDD.t1620 1.4705
R31339 VDD.t4693 VDD.n8841 1.4705
R31340 VDD.n8944 VDD.t1678 1.4705
R31341 VDD.t2470 VDD.n8944 1.4705
R31342 VDD.t2214 VDD.n8847 1.4705
R31343 VDD.n8847 VDD.t600 1.4705
R31344 VDD.t3527 VDD.n8933 1.4705
R31345 VDD.n8933 VDD.t4227 1.4705
R31346 VDD.n8899 VDD.t4019 1.4705
R31347 VDD.t2531 VDD.n8899 1.4705
R31348 VDD.n9019 VDD.t4083 1.4705
R31349 VDD.t4291 VDD.n9019 1.4705
R31350 VDD.t4111 VDD.n8905 1.4705
R31351 VDD.n8905 VDD.t2626 1.4705
R31352 VDD.t2292 VDD.n9006 1.4705
R31353 VDD.n9006 VDD.t2562 1.4705
R31354 VDD.n8950 VDD.t2329 1.4705
R31355 VDD.t711 VDD.n8950 1.4705
R31356 VDD.n9041 VDD.t4487 1.4705
R31357 VDD.t3025 VDD.n9041 1.4705
R31358 VDD.t4179 VDD.n8974 1.4705
R31359 VDD.n8974 VDD.t4367 1.4705
R31360 VDD.t2194 VDD.n9030 1.4705
R31361 VDD.n9030 VDD.t565 1.4705
R31362 VDD.n9025 VDD.t1799 1.4705
R31363 VDD.t2065 VDD.n9025 1.4705
R31364 VDD.t2306 VDD.n9154 1.4705
R31365 VDD.n9154 VDD.t684 1.4705
R31366 VDD.n9072 VDD.t1896 1.4705
R31367 VDD.t2132 VDD.n9072 1.4705
R31368 VDD.n189 VDD.t2047 1.4705
R31369 VDD.t4605 VDD.n189 1.4705
R31370 VDD.n173 VDD.t4407 1.4705
R31371 VDD.t4631 VDD.n173 1.4705
R31372 VDD.n9122 VDD.t2232 1.4705
R31373 VDD.t627 VDD.n9122 1.4705
R31374 VDD.n9094 VDD.t1839 1.4705
R31375 VDD.t2092 VDD.n9094 1.4705
R31376 VDD.n1159 VDD.t4641 1.4705
R31377 VDD.t1680 VDD.n1159 1.4705
R31378 VDD.t741 VDD.n1747 1.4705
R31379 VDD.n1747 VDD.t4641 1.4705
R31380 VDD.n981 VDD.t463 1.4705
R31381 VDD.n981 VDD.t451 1.4705
R31382 VDD.n978 VDD.t437 1.4705
R31383 VDD.n978 VDD.t423 1.4705
R31384 VDD.n1714 VDD.t2945 1.4705
R31385 VDD.n1714 VDD.t3137 1.4705
R31386 VDD.n725 VDD.t2723 1.4705
R31387 VDD.t2945 VDD.n725 1.4705
R31388 VDD.t2721 VDD.n714 1.4705
R31389 VDD.t2941 VDD.n714 1.4705
R31390 VDD.n723 VDD.t2509 1.4705
R31391 VDD.n723 VDD.t2721 1.4705
R31392 VDD.n1738 VDD.t1291 1.4705
R31393 VDD.n1738 VDD.t1506 1.4705
R31394 VDD.t3817 VDD.n947 1.4705
R31395 VDD.n947 VDD.t1291 1.4705
R31396 VDD.n1035 VDD.t427 1.4705
R31397 VDD.n1035 VDD.t445 1.4705
R31398 VDD.n1037 VDD.t432 1.4705
R31399 VDD.n1037 VDD.t435 1.4705
R31400 VDD.n913 VDD.t4379 1.4705
R31401 VDD.t4583 VDD.n913 1.4705
R31402 VDD.n908 VDD.t2827 1.4705
R31403 VDD.n908 VDD.t4379 1.4705
R31404 VDD.n1068 VDD.t1747 1.4705
R31405 VDD.t1986 VDD.n1068 1.4705
R31406 VDD.n1063 VDD.t1528 1.4705
R31407 VDD.n1063 VDD.t1747 1.4705
R31408 VDD.n1042 VDD.t461 1.4705
R31409 VDD.n1042 VDD.t464 1.4705
R31410 VDD.n1040 VDD.t454 1.4705
R31411 VDD.n1040 VDD.t455 1.4705
R31412 VDD.n1491 VDD.t1909 1.4705
R31413 VDD.t739 VDD.n1491 1.4705
R31414 VDD.n1486 VDD.t1684 1.4705
R31415 VDD.n1486 VDD.t1909 1.4705
R31416 VDD.n1456 VDD.t4513 1.4705
R31417 VDD.t4739 VDD.n1456 1.4705
R31418 VDD.n1451 VDD.t1934 1.4705
R31419 VDD.n1451 VDD.t4513 1.4705
R31420 VDD.n1410 VDD.t3159 1.4705
R31421 VDD.n1410 VDD.t1511 1.4705
R31422 VDD.n1403 VDD.t1676 1.4705
R31423 VDD.t3159 VDD.n1403 1.4705
R31424 VDD.n1489 VDD.t1682 1.4705
R31425 VDD.n1489 VDD.t4655 1.4705
R31426 VDD.n1488 VDD.t1472 1.4705
R31427 VDD.t1682 VDD.n1488 1.4705
R31428 VDD.n1454 VDD.t4315 1.4705
R31429 VDD.n1454 VDD.t4511 1.4705
R31430 VDD.n1453 VDD.t1700 1.4705
R31431 VDD.t4315 VDD.n1453 1.4705
R31432 VDD.t2969 VDD.n1392 1.4705
R31433 VDD.t1298 VDD.n1392 1.4705
R31434 VDD.n1401 VDD.t1450 1.4705
R31435 VDD.n1401 VDD.t2969 1.4705
R31436 VDD.n1215 VDD.t3485 1.4705
R31437 VDD.t4671 VDD.n1215 1.4705
R31438 VDD.n1210 VDD.t3659 1.4705
R31439 VDD.n1210 VDD.t3485 1.4705
R31440 VDD.n1273 VDD.t1706 1.4705
R31441 VDD.n1273 VDD.t1846 1.4705
R31442 VDD.n1242 VDD.t4675 1.4705
R31443 VDD.t1706 VDD.n1242 1.4705
R31444 VDD.n1101 VDD.t362 1.4705
R31445 VDD.n1101 VDD.t372 1.4705
R31446 VDD.n1103 VDD.t370 1.4705
R31447 VDD.n1103 VDD.t335 1.4705
R31448 VDD.n1598 VDD.t3728 1.4705
R31449 VDD.n1598 VDD.t2189 1.4705
R31450 VDD.t786 VDD.n1603 1.4705
R31451 VDD.n1603 VDD.t3728 1.4705
R31452 VDD.n1501 VDD.t3523 1.4705
R31453 VDD.t1943 VDD.n1501 1.4705
R31454 VDD.n1500 VDD.t4697 1.4705
R31455 VDD.t3523 VDD.n1500 1.4705
R31456 VDD.n1623 VDD.t354 1.4705
R31457 VDD.n1623 VDD.t349 1.4705
R31458 VDD.n1621 VDD.t337 1.4705
R31459 VDD.n1621 VDD.t338 1.4705
R31460 VDD.n1527 VDD.t1872 1.4705
R31461 VDD.t1626 VDD.n1527 1.4705
R31462 VDD.n1516 VDD.t2432 1.4705
R31463 VDD.t696 VDD.n1516 1.4705
R31464 VDD.n1540 VDD.t1192 1.4705
R31465 VDD.t998 VDD.n1540 1.4705
R31466 VDD.t1668 VDD.n1562 1.4705
R31467 VDD.n1562 VDD.t4207 1.4705
R31468 VDD.n1172 VDD.t3005 1.4705
R31469 VDD.t4141 VDD.n1172 1.4705
R31470 VDD.n1167 VDD.t1686 1.4705
R31471 VDD.n1167 VDD.t3005 1.4705
R31472 VDD.n1185 VDD.t1990 1.4705
R31473 VDD.t1762 VDD.n1185 1.4705
R31474 VDD.n1180 VDD.t4567 1.4705
R31475 VDD.n1180 VDD.t1990 1.4705
R31476 VDD.n1089 VDD.t340 1.4705
R31477 VDD.n1089 VDD.t358 1.4705
R31478 VDD.n1087 VDD.t347 1.4705
R31479 VDD.n1087 VDD.t357 1.4705
R31480 VDD.n1420 VDD.t460 1.4705
R31481 VDD.n1420 VDD.t458 1.4705
R31482 VDD.n1422 VDD.t444 1.4705
R31483 VDD.n1422 VDD.t434 1.4705
R31484 VDD.n854 VDD.t425 1.4705
R31485 VDD.n854 VDD.t457 1.4705
R31486 VDD.n856 VDD.t442 1.4705
R31487 VDD.n856 VDD.t429 1.4705
R31488 VDD.n746 VDD.t342 1.4705
R31489 VDD.n746 VDD.t356 1.4705
R31490 VDD.n1675 VDD.t345 1.4705
R31491 VDD.n1675 VDD.t361 1.4705
R31492 VDD.n743 VDD.t336 1.4705
R31493 VDD.n743 VDD.t341 1.4705
R31494 VDD.n1681 VDD.t344 1.4705
R31495 VDD.n1681 VDD.t377 1.4705
R31496 VDD.n1340 VDD.t867 1.4705
R31497 VDD.n1340 VDD.t3799 1.4705
R31498 VDD.n1310 VDD.t593 1.4705
R31499 VDD.t867 VDD.n1310 1.4705
R31500 VDD.n1656 VDD.t2746 1.4705
R31501 VDD.t1092 VDD.n1656 1.4705
R31502 VDD.t3849 VDD.n1315 1.4705
R31503 VDD.n1315 VDD.t2746 1.4705
R31504 VDD.n740 VDD.t353 1.4705
R31505 VDD.n740 VDD.t346 1.4705
R31506 VDD.n1687 VDD.t355 1.4705
R31507 VDD.n1687 VDD.t4984 1.4705
R31508 VDD.n1694 VDD.t452 1.4705
R31509 VDD.n1694 VDD.t466 1.4705
R31510 VDD.n737 VDD.t456 1.4705
R31511 VDD.n737 VDD.t436 1.4705
R31512 VDD.n1387 VDD.t2028 1.4705
R31513 VDD.n1387 VDD.t4593 1.4705
R31514 VDD.n1078 VDD.t583 1.4705
R31515 VDD.t2028 VDD.n1078 1.4705
R31516 VDD.n1283 VDD.t3479 1.4705
R31517 VDD.t3669 VDD.n1283 1.4705
R31518 VDD.t892 VDD.n1361 1.4705
R31519 VDD.n1361 VDD.t3479 1.4705
R31520 VDD.n1648 VDD.t3543 1.4705
R31521 VDD.n1648 VDD.t3343 1.4705
R31522 VDD.t3435 VDD.n1247 1.4705
R31523 VDD.n1247 VDD.t3543 1.4705
R31524 VDD.t1107 VDD.n694 1.4705
R31525 VDD.t1289 VDD.n694 1.4705
R31526 VDD.n945 VDD.t3600 1.4705
R31527 VDD.n945 VDD.t1107 1.4705
R31528 VDD.n6953 VDD.n6952 1.46537
R31529 VDD.n6957 VDD.n6956 1.46537
R31530 VDD.n6926 VDD.n6925 1.46537
R31531 VDD.n7011 VDD.n7010 1.46537
R31532 VDD.n7009 VDD.n7008 1.46537
R31533 VDD.n7004 VDD.n7003 1.46537
R31534 VDD.n6503 VDD.n6502 1.46537
R31535 VDD.n6501 VDD.n6500 1.46537
R31536 VDD.n6452 VDD.n6451 1.46537
R31537 VDD.n6543 VDD.n6542 1.46537
R31538 VDD.n6547 VDD.n6546 1.46537
R31539 VDD.n6541 VDD.n6540 1.46537
R31540 VDD.n6140 VDD.n6139 1.46537
R31541 VDD.n6144 VDD.n6143 1.46537
R31542 VDD.n6148 VDD.n6147 1.46537
R31543 VDD.n6133 VDD.n6132 1.46537
R31544 VDD.n6129 VDD.n6128 1.46537
R31545 VDD.n6125 VDD.n6124 1.46537
R31546 VDD.n6121 VDD.n6120 1.46537
R31547 VDD.n6048 VDD.n6047 1.46537
R31548 VDD.n6052 VDD.n6051 1.46537
R31549 VDD.n6056 VDD.n6055 1.46537
R31550 VDD.n6079 VDD.n6078 1.46537
R31551 VDD.n6083 VDD.n6082 1.46537
R31552 VDD.n6087 VDD.n6086 1.46537
R31553 VDD.n6091 VDD.n6090 1.46537
R31554 VDD.n6814 VDD.n6813 1.46537
R31555 VDD.n6818 VDD.n6817 1.46537
R31556 VDD.n6822 VDD.n6821 1.46537
R31557 VDD.n6827 VDD.n6826 1.46537
R31558 VDD.n6831 VDD.n6830 1.46537
R31559 VDD.n6835 VDD.n6834 1.46537
R31560 VDD.n6839 VDD.n6838 1.46537
R31561 VDD.n6781 VDD.n6780 1.46537
R31562 VDD.n6785 VDD.n6784 1.46537
R31563 VDD.n6789 VDD.n6788 1.46537
R31564 VDD.n6774 VDD.n6773 1.46537
R31565 VDD.n6770 VDD.n6769 1.46537
R31566 VDD.n6766 VDD.n6765 1.46537
R31567 VDD.n6762 VDD.n6761 1.46537
R31568 VDD.n6327 VDD.n5488 1.3379
R31569 VDD.n6013 VDD.n5488 1.3306
R31570 VDD.n7932 VDD.n7931 1.30325
R31571 VDD.n7897 VDD.n7896 1.30325
R31572 VDD.n8037 VDD.n8036 1.30325
R31573 VDD.n7951 VDD.n7949 1.27338
R31574 VDD.n7958 VDD.n7956 1.27338
R31575 VDD.n7954 VDD.n7952 1.27228
R31576 VDD.n8063 VDD.n8061 1.27228
R31577 VDD.n8059 VDD.n8057 1.27228
R31578 VDD.n8056 VDD.n8054 1.27228
R31579 VDD.n2383 VDD.n2381 1.27228
R31580 VDD.n7021 VDD.n7019 1.27228
R31581 VDD.n7017 VDD.n7015 1.27228
R31582 VDD.n6966 VDD.n6964 1.27228
R31583 VDD.n6974 VDD.n6972 1.27228
R31584 VDD.n6970 VDD.n6968 1.27228
R31585 VDD.n7011 VDD.n7009 1.27228
R31586 VDD.n6957 VDD.n6953 1.27228
R31587 VDD.n5296 VDD.n5294 1.27228
R31588 VDD.n6555 VDD.n6553 1.27228
R31589 VDD.n6559 VDD.n6557 1.27228
R31590 VDD.n6511 VDD.n6509 1.27228
R31591 VDD.n6516 VDD.n6514 1.27228
R31592 VDD.n6520 VDD.n6518 1.27228
R31593 VDD.n6547 VDD.n6543 1.27228
R31594 VDD.n6503 VDD.n6501 1.27228
R31595 VDD.n6125 VDD.n6121 1.27228
R31596 VDD.n6133 VDD.n6129 1.27228
R31597 VDD.n6148 VDD.n6144 1.27228
R31598 VDD.n6091 VDD.n6087 1.27228
R31599 VDD.n6083 VDD.n6079 1.27228
R31600 VDD.n6056 VDD.n6052 1.27228
R31601 VDD.n6155 VDD.n6153 1.27228
R31602 VDD.n6098 VDD.n6096 1.27228
R31603 VDD.n6839 VDD.n6835 1.27228
R31604 VDD.n6831 VDD.n6827 1.27228
R31605 VDD.n6822 VDD.n6818 1.27228
R31606 VDD.n6766 VDD.n6762 1.27228
R31607 VDD.n6774 VDD.n6770 1.27228
R31608 VDD.n6789 VDD.n6785 1.27228
R31609 VDD.n6844 VDD.n6843 1.27228
R31610 VDD.n6794 VDD.n6793 1.27228
R31611 VDD.n1511 VDD.t1666 1.27155
R31612 VDD.n1560 VDD.t4206 1.27155
R31613 VDD.n1538 VDD.t1190 1.27155
R31614 VDD.n1536 VDD.t996 1.27155
R31615 VDD.n1514 VDD.t2431 1.27155
R31616 VDD.n1513 VDD.t694 1.27155
R31617 VDD.n1525 VDD.t1871 1.27155
R31618 VDD.n1524 VDD.t1625 1.27155
R31619 VDD.n8089 VDD.n8088 1.26911
R31620 VDD.n1763 VDD.n1762 1.23698
R31621 VDD.n6327 VDD.n6326 1.14768
R31622 VDD.n6396 VDD.t412 1.1382
R31623 VDD.n6577 VDD.t408 1.1382
R31624 VDD.n7040 VDD.t99 1.1382
R31625 VDD.n7086 VDD.t76 1.1382
R31626 VDD.n7025 VDD.n7024 1.13692
R31627 VDD.n6414 VDD.n5297 1.13692
R31628 VDD.n6562 VDD.n6561 1.13692
R31629 VDD.n6877 VDD.n2384 1.13692
R31630 VDD.n12624 VDD.t837 1.00929
R31631 VDD.n12564 VDD.t1165 1.00929
R31632 VDD.n12568 VDD.t1768 1.00929
R31633 VDD.n12571 VDD.t1176 1.00929
R31634 VDD.n12575 VDD.t1538 1.00929
R31635 VDD.n12557 VDD.t3219 1.00929
R31636 VDD.n8624 VDD.t3125 1.00929
R31637 VDD.n8625 VDD.t3439 1.00929
R31638 VDD.n18 VDD.t4045 1.00929
R31639 VDD.n21 VDD.t3449 1.00929
R31640 VDD.n22 VDD.t3807 1.00929
R31641 VDD.n23 VDD.t1222 1.00929
R31642 VDD.n8631 VDD.t2997 1.00929
R31643 VDD.n8628 VDD.t3299 1.00929
R31644 VDD.n19 VDD.t3873 1.00929
R31645 VDD.n12607 VDD.t3309 1.00929
R31646 VDD.n12603 VDD.t3639 1.00929
R31647 VDD.n12600 VDD.t1090 1.00929
R31648 VDD.n8655 VDD.t3209 1.00929
R31649 VDD.n8656 VDD.t3509 1.00929
R31650 VDD.n27 VDD.t4135 1.00929
R31651 VDD.n12531 VDD.t3529 1.00929
R31652 VDD.n12536 VDD.t3893 1.00929
R31653 VDD.n12540 VDD.t1303 1.00929
R31654 VDD.n8662 VDD.t3065 1.00929
R31655 VDD.n8659 VDD.t3358 1.00929
R31656 VDD.n28 VDD.t3975 1.00929
R31657 VDD.n12532 VDD.t3374 1.00929
R31658 VDD.n12537 VDD.t3742 1.00929
R31659 VDD.n12541 VDD.t1159 1.00929
R31660 VDD.n8610 VDD.t3843 1.00929
R31661 VDD.n8611 VDD.t4213 1.00929
R31662 VDD.n37 VDD.t640 1.00929
R31663 VDD.n40 VDD.t4231 1.00929
R31664 VDD.n82 VDD.t4551 1.00929
R31665 VDD.n86 VDD.t2034 1.00929
R31666 VDD.n8617 VDD.t3469 1.00929
R31667 VDD.n8614 VDD.t3801 1.00929
R31668 VDD.n38 VDD.t4401 1.00929
R31669 VDD.n41 VDD.t3821 1.00929
R31670 VDD.n83 VDD.t4221 1.00929
R31671 VDD.n87 VDD.t1614 1.00929
R31672 VDD.n8688 VDD.t1428 1.00929
R31673 VDD.n8689 VDD.t1778 1.00929
R31674 VDD.n98 VDD.t2513 1.00929
R31675 VDD.n101 VDD.t1792 1.00929
R31676 VDD.n102 VDD.t2224 1.00929
R31677 VDD.n103 VDD.t3795 1.00929
R31678 VDD.n8695 VDD.t4167 1.00929
R31679 VDD.n8692 VDD.t4483 1.00929
R31680 VDD.n99 VDD.t987 1.00929
R31681 VDD.n12513 VDD.t4491 1.00929
R31682 VDD.n12509 VDD.t752 1.00929
R31683 VDD.n12506 VDD.t2411 1.00929
R31684 VDD.n8596 VDD.t1509 1.00929
R31685 VDD.n8597 VDD.t1876 1.00929
R31686 VDD.n107 VDD.t2600 1.00929
R31687 VDD.n12475 VDD.t1893 1.00929
R31688 VDD.n12480 VDD.t2350 1.00929
R31689 VDD.n12484 VDD.t3879 1.00929
R31690 VDD.n8603 VDD.t4247 1.00929
R31691 VDD.n8600 VDD.t4549 1.00929
R31692 VDD.n108 VDD.t1050 1.00929
R31693 VDD.n12476 VDD.t4575 1.00929
R31694 VDD.n12481 VDD.t832 1.00929
R31695 VDD.n12485 VDD.t2499 1.00929
R31696 VDD.n8726 VDD.t1056 1.00929
R31697 VDD.n8727 VDD.t1386 1.00929
R31698 VDD.n117 VDD.t2015 1.00929
R31699 VDD.n120 VDD.t1396 1.00929
R31700 VDD.n128 VDD.t1766 1.00929
R31701 VDD.n132 VDD.t3394 1.00929
R31702 VDD.n8733 VDD.t1824 1.00929
R31703 VDD.n8730 VDD.t2222 1.00929
R31704 VDD.n118 VDD.t2893 1.00929
R31705 VDD.n121 VDD.t2239 1.00929
R31706 VDD.n129 VDD.t2674 1.00929
R31707 VDD.n133 VDD.t4197 1.00929
R31708 VDD.n8583 VDD.t1131 1.00929
R31709 VDD.n8584 VDD.t1462 1.00929
R31710 VDD.n178 VDD.t2110 1.00929
R31711 VDD.n181 VDD.t1478 1.00929
R31712 VDD.n182 VDD.t1861 1.00929
R31713 VDD.n183 VDD.t3487 1.00929
R31714 VDD.n8590 VDD.t3827 1.00929
R31715 VDD.n8587 VDD.t4195 1.00929
R31716 VDD.n179 VDD.t615 1.00929
R31717 VDD.n12457 VDD.t4217 1.00929
R31718 VDD.n12453 VDD.t4535 1.00929
R31719 VDD.n12450 VDD.t2005 1.00929
R31720 VDD.n1765 VDD.t1672 1.00929
R31721 VDD.n11056 VDD.t1313 1.00929
R31722 VDD.n11076 VDD.t3883 1.00929
R31723 VDD.n11089 VDD.t1296 1.00929
R31724 VDD.n648 VDD.t969 1.00929
R31725 VDD.n641 VDD.t3943 1.00929
R31726 VDD.n5708 VDD.t2129 1.00929
R31727 VDD.n5709 VDD.t1741 1.00929
R31728 VDD.n1781 VDD.t4307 1.00929
R31729 VDD.n11008 VDD.t1731 1.00929
R31730 VDD.n11013 VDD.t1358 1.00929
R31731 VDD.n11017 VDD.t2071 1.00929
R31732 VDD.n5715 VDD.t4707 1.00929
R31733 VDD.n5712 VDD.t4359 1.00929
R31734 VDD.n1782 VDD.t2837 1.00929
R31735 VDD.n11009 VDD.t4349 1.00929
R31736 VDD.n11014 VDD.t3983 1.00929
R31737 VDD.n11018 VDD.t1423 1.00929
R31738 VDD.n5734 VDD.t1560 1.00929
R31739 VDD.n5735 VDD.t1203 1.00929
R31740 VDD.n1788 VDD.t3779 1.00929
R31741 VDD.n1791 VDD.t1194 1.00929
R31742 VDD.n1799 VDD.t856 1.00929
R31743 VDD.n1803 VDD.t2887 1.00929
R31744 VDD.n5741 VDD.t4191 1.00929
R31745 VDD.n5738 VDD.t3825 1.00929
R31746 VDD.n1789 VDD.t2237 1.00929
R31747 VDD.n1792 VDD.t3811 1.00929
R31748 VDD.n1800 VDD.t3451 1.00929
R31749 VDD.n1804 VDD.t2235 1.00929
R31750 VDD.n5695 VDD.t1141 1.00929
R31751 VDD.n5696 VDD.t807 1.00929
R31752 VDD.n1834 VDD.t3353 1.00929
R31753 VDD.n1837 VDD.t793 1.00929
R31754 VDD.n1838 VDD.t4531 1.00929
R31755 VDD.n1839 VDD.t3845 1.00929
R31756 VDD.n5702 VDD.t948 1.00929
R31757 VDD.n5699 VDD.t4713 1.00929
R31758 VDD.n1835 VDD.t3169 1.00929
R31759 VDD.n10991 VDD.t4699 1.00929
R31760 VDD.n10987 VDD.t4327 1.00929
R31761 VDD.n10984 VDD.t3141 1.00929
R31762 VDD.n5789 VDD.t3069 1.00929
R31763 VDD.n5790 VDD.t2729 1.00929
R31764 VDD.n1843 VDD.t1033 1.00929
R31765 VDD.n10953 VDD.t2707 1.00929
R31766 VDD.n10958 VDD.t2283 1.00929
R31767 VDD.n10962 VDD.t939 1.00929
R31768 VDD.n5796 VDD.t4643 1.00929
R31769 VDD.n5793 VDD.t4293 1.00929
R31770 VDD.n1844 VDD.t2780 1.00929
R31771 VDD.n10954 VDD.t4281 1.00929
R31772 VDD.n10959 VDD.t3911 1.00929
R31773 VDD.n10963 VDD.t4127 1.00929
R31774 VDD.n5682 VDD.t2543 1.00929
R31775 VDD.n5683 VDD.t2108 1.00929
R31776 VDD.n1853 VDD.t4629 1.00929
R31777 VDD.n1856 VDD.t2096 1.00929
R31778 VDD.n1882 VDD.t1688 1.00929
R31779 VDD.n1886 VDD.t1661 1.00929
R31780 VDD.n5689 VDD.t4131 1.00929
R31781 VDD.n5686 VDD.t3761 1.00929
R31782 VDD.n1854 VDD.t2157 1.00929
R31783 VDD.n1857 VDD.t3744 1.00929
R31784 VDD.n1883 VDD.t3376 1.00929
R31785 VDD.n1887 VDD.t701 1.00929
R31786 VDD.n5844 VDD.t859 1.00929
R31787 VDD.n5845 VDD.t4623 1.00929
R31788 VDD.n1899 VDD.t3095 1.00929
R31789 VDD.n1902 VDD.t4603 1.00929
R31790 VDD.n1903 VDD.t4255 1.00929
R31791 VDD.n1904 VDD.t2444 1.00929
R31792 VDD.n5851 VDD.t1770 1.00929
R31793 VDD.n5848 VDD.t1414 1.00929
R31794 VDD.n1900 VDD.t3993 1.00929
R31795 VDD.n10936 VDD.t1402 1.00929
R31796 VDD.n10932 VDD.t1053 1.00929
R31797 VDD.n10929 VDD.t1926 1.00929
R31798 VDD.n5669 VDD.t4445 1.00929
R31799 VDD.n5670 VDD.t4119 1.00929
R31800 VDD.n1908 VDD.t2573 1.00929
R31801 VDD.n10898 VDD.t4099 1.00929
R31802 VDD.n10903 VDD.t3704 1.00929
R31803 VDD.n10907 VDD.t3183 1.00929
R31804 VDD.n5676 VDD.t1947 1.00929
R31805 VDD.n5673 VDD.t1583 1.00929
R31806 VDD.n1909 VDD.t4161 1.00929
R31807 VDD.n10899 VDD.t1558 1.00929
R31808 VDD.n10904 VDD.t1187 1.00929
R31809 VDD.n10908 VDD.t2177 1.00929
R31810 VDD.n5877 VDD.t3923 1.00929
R31811 VDD.n5878 VDD.t3565 1.00929
R31812 VDD.n5879 VDD.t1939 1.00929
R31813 VDD.n5491 VDD.t3547 1.00929
R31814 VDD.n5496 VDD.t3225 1.00929
R31815 VDD.n5500 VDD.t3885 1.00929
R31816 VDD.n5898 VDD.t3797 1.00929
R31817 VDD.n5895 VDD.t3463 1.00929
R31818 VDD.n5891 VDD.t1802 1.00929
R31819 VDD.n5492 VDD.t3443 1.00929
R31820 VDD.n5497 VDD.t3113 1.00929
R31821 VDD.n5501 VDD.t3404 1.00929
R31822 VDD.n5627 VDD.t2851 1.00929
R31823 VDD.n5628 VDD.t2495 1.00929
R31824 VDD.n1926 VDD.t802 1.00929
R31825 VDD.n1929 VDD.t2486 1.00929
R31826 VDD.n1930 VDD.t2026 1.00929
R31827 VDD.n1931 VDD.t3217 1.00929
R31828 VDD.n5634 VDD.t3295 1.00929
R31829 VDD.n5631 VDD.t2989 1.00929
R31830 VDD.n1927 VDD.t1266 1.00929
R31831 VDD.n10881 VDD.t2967 1.00929
R31832 VDD.n10877 VDD.t2598 1.00929
R31833 VDD.n10874 VDD.t4169 1.00929
R31834 VDD.n5606 VDD.t829 1.00929
R31835 VDD.n5607 VDD.t4601 1.00929
R31836 VDD.n1935 VDD.t3081 1.00929
R31837 VDD.n10843 VDD.t4577 1.00929
R31838 VDD.n10848 VDD.t4241 1.00929
R31839 VDD.n10852 VDD.t817 1.00929
R31840 VDD.n5613 VDD.t4449 1.00929
R31841 VDD.n5610 VDD.t4123 1.00929
R31842 VDD.n1936 VDD.t2576 1.00929
R31843 VDD.n10844 VDD.t4101 1.00929
R31844 VDD.n10849 VDD.t3710 1.00929
R31845 VDD.n10853 VDD.t3321 1.00929
R31846 VDD.n5585 VDD.t2750 1.00929
R31847 VDD.n5586 VDD.t2377 1.00929
R31848 VDD.n1945 VDD.t678 1.00929
R31849 VDD.n1948 VDD.t2357 1.00929
R31850 VDD.n1974 VDD.t1898 1.00929
R31851 VDD.n1978 VDD.t2053 1.00929
R31852 VDD.n5592 VDD.t2153 1.00929
R31853 VDD.n5589 VDD.t1758 1.00929
R31854 VDD.n1946 VDD.t4323 1.00929
R31855 VDD.n1949 VDD.t1743 1.00929
R31856 VDD.n1975 VDD.t1374 1.00929
R31857 VDD.n1979 VDD.t4495 1.00929
R31858 VDD.n2106 VDD.t3865 1.00929
R31859 VDD.n2111 VDD.t3517 1.00929
R31860 VDD.n1991 VDD.t1878 1.00929
R31861 VDD.n1994 VDD.t3505 1.00929
R31862 VDD.n1995 VDD.t3175 1.00929
R31863 VDD.n1998 VDD.t1168 1.00929
R31864 VDD.n8096 VDD.t653 1.00929
R31865 VDD.n2114 VDD.t4457 1.00929
R31866 VDD.n1992 VDD.t2935 1.00929
R31867 VDD.n10826 VDD.t4431 1.00929
R31868 VDD.n10822 VDD.t4075 1.00929
R31869 VDD.n1999 VDD.t773 1.00929
R31870 VDD.n2093 VDD.t3335 1.00929
R31871 VDD.n2094 VDD.t3043 1.00929
R31872 VDD.n2008 VDD.t1326 1.00929
R31873 VDD.n10785 VDD.t3029 1.00929
R31874 VDD.n10790 VDD.t2664 1.00929
R31875 VDD.n10794 VDD.t1928 1.00929
R31876 VDD.n2100 VDD.t3257 1.00929
R31877 VDD.n2097 VDD.t2929 1.00929
R31878 VDD.n2009 VDD.t1210 1.00929
R31879 VDD.n10786 VDD.t2909 1.00929
R31880 VDD.n10791 VDD.t2541 1.00929
R31881 VDD.n10795 VDD.t1416 1.00929
R31882 VDD.n8122 VDD.t1016 1.00929
R31883 VDD.n8123 VDD.t637 1.00929
R31884 VDD.n2018 VDD.t3251 1.00929
R31885 VDD.n2021 VDD.t603 1.00929
R31886 VDD.n2029 VDD.t4395 1.00929
R31887 VDD.n2033 VDD.t3223 1.00929
R31888 VDD.n8129 VDD.t2754 1.00929
R31889 VDD.n8126 VDD.t2383 1.00929
R31890 VDD.n2019 VDD.t681 1.00929
R31891 VDD.n2022 VDD.t2363 1.00929
R31892 VDD.n2030 VDD.t1900 1.00929
R31893 VDD.n2034 VDD.t2230 1.00929
R31894 VDD.n8166 VDD.t2125 1.00929
R31895 VDD.n8181 VDD.t1735 1.00929
R31896 VDD.n8201 VDD.t4305 1.00929
R31897 VDD.n8214 VDD.t1721 1.00929
R31898 VDD.n8236 VDD.t1353 1.00929
R31899 VDD.n8249 VDD.t3037 1.00929
R31900 VDD.n9088 VDD.t3135 1.00929
R31901 VDD.n9089 VDD.t4647 1.00929
R31902 VDD.n9086 VDD.t2403 1.00929
R31903 VDD.n9087 VDD.t2768 1.00929
R31904 VDD.n9075 VDD.t3696 1.00929
R31905 VDD.n9076 VDD.t4063 1.00929
R31906 VDD.n8463 VDD.t4657 1.00929
R31907 VDD.n8467 VDD.t4077 1.00929
R31908 VDD.n8468 VDD.t4435 1.00929
R31909 VDD.n8469 VDD.t1870 1.00929
R31910 VDD.n9082 VDD.t2258 1.00929
R31911 VDD.n9079 VDD.t2676 1.00929
R31912 VDD.n8464 VDD.t3261 1.00929
R31913 VDD.n9175 VDD.t2687 1.00929
R31914 VDD.n9171 VDD.t3055 1.00929
R31915 VDD.n9168 VDD.t4541 1.00929
R31916 VDD.n8532 VDD.t1199 1.00929
R31917 VDD.n8533 VDD.t1540 1.00929
R31918 VDD.n8534 VDD.t2212 1.00929
R31919 VDD.n8540 VDD.t1564 1.00929
R31920 VDD.n8541 VDD.t1966 1.00929
R31921 VDD.n8542 VDD.t3559 1.00929
R31922 VDD.n8578 VDD.t1412 1.00929
R31923 VDD.n8575 VDD.t1764 1.00929
R31924 VDD.n8571 VDD.t2493 1.00929
R31925 VDD.n8568 VDD.t1780 1.00929
R31926 VDD.n8564 VDD.t2206 1.00929
R31927 VDD.n8561 VDD.t3783 1.00929
R31928 VDD.n8776 VDD.t3165 1.00929
R31929 VDD.n8777 VDD.t3477 1.00929
R31930 VDD.n8778 VDD.t4085 1.00929
R31931 VDD.n8779 VDD.t3497 1.00929
R31932 VDD.n8780 VDD.t3855 1.00929
R31933 VDD.n8522 VDD.t1269 1.00929
R31934 VDD.n8796 VDD.t1493 1.00929
R31935 VDD.n8793 VDD.t1859 1.00929
R31936 VDD.n8789 VDD.t2580 1.00929
R31937 VDD.n8786 VDD.t1880 1.00929
R31938 VDD.n8782 VDD.t2320 1.00929
R31939 VDD.n8523 VDD.t3867 1.00929
R31940 VDD.n8514 VDD.t3651 1.00929
R31941 VDD.n8850 VDD.t4033 1.00929
R31942 VDD.n8855 VDD.t4613 1.00929
R31943 VDD.n8859 VDD.t4047 1.00929
R31944 VDD.n8864 VDD.t4389 1.00929
R31945 VDD.n8868 VDD.t1821 1.00929
R31946 VDD.n8515 VDD.t2104 1.00929
R31947 VDD.n8851 VDD.t2535 1.00929
R31948 VDD.n8856 VDD.t3131 1.00929
R31949 VDD.n8860 VDD.t2553 1.00929
R31950 VDD.n8865 VDD.t2921 1.00929
R31951 VDD.n8869 VDD.t4417 1.00929
R31952 VDD.n8907 VDD.t1255 1.00929
R31953 VDD.n8908 VDD.t1609 1.00929
R31954 VDD.n8909 VDD.t2271 1.00929
R31955 VDD.n8910 VDD.t1628 1.00929
R31956 VDD.n8911 VDD.t2021 1.00929
R31957 VDD.n8503 VDD.t3612 1.00929
R31958 VDD.n8927 VDD.t3869 1.00929
R31959 VDD.n8924 VDD.t4237 1.00929
R31960 VDD.n8920 VDD.t671 1.00929
R31961 VDD.n8917 VDD.t4249 1.00929
R31962 VDD.n8913 VDD.t4591 1.00929
R31963 VDD.n8504 VDD.t2067 1.00929
R31964 VDD.n8495 VDD.t1827 1.00929
R31965 VDD.n8977 VDD.t2226 1.00929
R31966 VDD.n8982 VDD.t2895 1.00929
R31967 VDD.n8986 VDD.t2241 1.00929
R31968 VDD.n8991 VDD.t2678 1.00929
R31969 VDD.n8995 VDD.t4203 1.00929
R31970 VDD.n8496 VDD.t2734 1.00929
R31971 VDD.n8978 VDD.t3071 1.00929
R31972 VDD.n8983 VDD.t3617 1.00929
R31973 VDD.n8987 VDD.t3085 1.00929
R31974 VDD.n8992 VDD.t3408 1.00929
R31975 VDD.n8996 VDD.t840 1.00929
R31976 VDD.n8477 VDD.t1920 1.00929
R31977 VDD.n8478 VDD.t2355 1.00929
R31978 VDD.n8479 VDD.t2991 1.00929
R31979 VDD.n8481 VDD.t2375 1.00929
R31980 VDD.n8482 VDD.t2770 1.00929
R31981 VDD.n8483 VDD.t4271 1.00929
R31982 VDD.n9061 VDD.t2165 1.00929
R31983 VDD.n9058 VDD.t2590 1.00929
R31984 VDD.n9054 VDD.t3179 1.00929
R31985 VDD.n9051 VDD.t2612 1.00929
R31986 VDD.n9047 VDD.t2987 1.00929
R31987 VDD.n9044 VDD.t4473 1.00929
R31988 VDD.n12624 VDD.t1485 1.00871
R31989 VDD.n12564 VDD.t1850 1.00871
R31990 VDD.n12568 VDD.t2564 1.00871
R31991 VDD.n12571 VDD.t1863 1.00871
R31992 VDD.n12575 VDD.t2298 1.00871
R31993 VDD.n12557 VDD.t3853 1.00871
R31994 VDD.n8624 VDD.t1573 1.00871
R31995 VDD.n8625 VDD.t1941 1.00871
R31996 VDD.n18 VDD.t2654 1.00871
R31997 VDD.n21 VDD.t1968 1.00871
R31998 VDD.n22 VDD.t2417 1.00871
R31999 VDD.n23 VDD.t3945 1.00871
R32000 VDD.n8631 VDD.t1783 1.00871
R32001 VDD.n8628 VDD.t2185 1.00871
R32002 VDD.n19 VDD.t2865 1.00871
R32003 VDD.n12607 VDD.t2208 1.00871
R32004 VDD.n12603 VDD.t2646 1.00871
R32005 VDD.n12600 VDD.t4173 1.00871
R32006 VDD.n8655 VDD.t3372 1.00871
R32007 VDD.n8656 VDD.t3720 1.00871
R32008 VDD.n27 VDD.t4329 1.00871
R32009 VDD.n12531 VDD.t3736 1.00871
R32010 VDD.n12536 VDD.t4129 1.00871
R32011 VDD.n12540 VDD.t1518 1.00871
R32012 VDD.n8662 VDD.t1887 1.00871
R32013 VDD.n8659 VDD.t2289 1.00871
R32014 VDD.n28 VDD.t2961 1.00871
R32015 VDD.n12532 VDD.t2322 1.00871
R32016 VDD.n12537 VDD.t2740 1.00871
R32017 VDD.n12541 VDD.t4253 1.00871
R32018 VDD.n8610 VDD.t4065 1.00871
R32019 VDD.n8611 VDD.t4391 1.00871
R32020 VDD.n37 VDD.t894 1.00871
R32021 VDD.n40 VDD.t4405 1.00871
R32022 VDD.n82 VDD.t630 1.00871
R32023 VDD.n86 VDD.t2267 1.00871
R32024 VDD.n8617 VDD.t690 1.00871
R32025 VDD.n8614 VDD.t1060 1.00871
R32026 VDD.n38 VDD.t1651 1.00871
R32027 VDD.n41 VDD.t1078 1.00871
R32028 VDD.n83 VDD.t1418 1.00871
R32029 VDD.n87 VDD.t3105 1.00871
R32030 VDD.n8688 VDD.t1656 1.00871
R32031 VDD.n8689 VDD.t2036 1.00871
R32032 VDD.n98 VDD.t2725 1.00871
R32033 VDD.n101 VDD.t2057 1.00871
R32034 VDD.n102 VDD.t2503 1.00871
R32035 VDD.n103 VDD.t4017 1.00871
R32036 VDD.n8695 VDD.t4355 1.00871
R32037 VDD.n8692 VDD.t4705 1.00871
R32038 VDD.n99 VDD.t1156 1.00871
R32039 VDD.n12513 VDD.t4723 1.00871
R32040 VDD.n12509 VDD.t980 1.00871
R32041 VDD.n12506 VDD.t2636 1.00871
R32042 VDD.n8596 VDD.t4149 1.00871
R32043 VDD.n8597 VDD.t4471 1.00871
R32044 VDD.n107 VDD.t971 1.00871
R32045 VDD.n12475 VDD.t4485 1.00871
R32046 VDD.n12480 VDD.t729 1.00871
R32047 VDD.n12484 VDD.t2388 1.00871
R32048 VDD.n8603 VDD.t4441 1.00871
R32049 VDD.n8600 VDD.t624 1.00871
R32050 VDD.n108 VDD.t1236 1.00871
R32051 VDD.n12476 VDD.t655 1.00871
R32052 VDD.n12481 VDD.t1039 1.00871
R32053 VDD.n12485 VDD.t2715 1.00871
R32054 VDD.n8726 VDD.t3631 1.00871
R32055 VDD.n8727 VDD.t4009 1.00871
R32056 VDD.n117 VDD.t4587 1.00871
R32057 VDD.n120 VDD.t4031 1.00871
R32058 VDD.n128 VDD.t4377 1.00871
R32059 VDD.n132 VDD.t1790 1.00871
R32060 VDD.n8733 VDD.t2080 1.00871
R32061 VDD.n8730 VDD.t2497 1.00871
R32062 VDD.n118 VDD.t3097 1.00871
R32063 VDD.n121 VDD.t2517 1.00871
R32064 VDD.n129 VDD.t2881 1.00871
R32065 VDD.n133 VDD.t4383 1.00871
R32066 VDD.n8583 VDD.t4219 1.00871
R32067 VDD.n8584 VDD.t4525 1.00871
R32068 VDD.n178 VDD.t1023 1.00871
R32069 VDD.n181 VDD.t4533 1.00871
R32070 VDD.n182 VDD.t796 1.00871
R32071 VDD.n183 VDD.t2457 1.00871
R32072 VDD.n8590 VDD.t2717 1.00871
R32073 VDD.n8587 VDD.t3059 1.00871
R32074 VDD.n179 VDD.t3602 1.00871
R32075 VDD.n12457 VDD.t3077 1.00871
R32076 VDD.n12453 VDD.t3386 1.00871
R32077 VDD.n12450 VDD.t827 1.00871
R32078 VDD.n1765 VDD.t3127 1.00871
R32079 VDD.n11056 VDD.t2800 1.00871
R32080 VDD.n11076 VDD.t1103 1.00871
R32081 VDD.n11089 VDD.t2792 1.00871
R32082 VDD.n648 VDD.t2394 1.00871
R32083 VDD.n641 VDD.t2044 1.00871
R32084 VDD.n5708 VDD.t2614 1.00871
R32085 VDD.n5709 VDD.t2187 1.00871
R32086 VDD.n1781 VDD.t4703 1.00871
R32087 VDD.n11008 VDD.t2171 1.00871
R32088 VDD.n11013 VDD.t1750 1.00871
R32089 VDD.n11017 VDD.t2869 1.00871
R32090 VDD.n5715 VDD.t2491 1.00871
R32091 VDD.n5712 VDD.t2069 1.00871
R32092 VDD.n1782 VDD.t4561 1.00871
R32093 VDD.n11009 VDD.t2049 1.00871
R32094 VDD.n11014 VDD.t1645 1.00871
R32095 VDD.n11018 VDD.t2365 1.00871
R32096 VDD.n5734 VDD.t4357 1.00871
R32097 VDD.n5735 VDD.t4021 1.00871
R32098 VDD.n1788 VDD.t2489 1.00871
R32099 VDD.n1791 VDD.t4003 1.00871
R32100 VDD.n1799 VDD.t3621 1.00871
R32101 VDD.n1803 VDD.t4035 1.00871
R32102 VDD.n5741 VDD.t1848 1.00871
R32103 VDD.n5738 VDD.t1482 1.00871
R32104 VDD.n1789 VDD.t4057 1.00871
R32105 VDD.n1792 VDD.t1474 1.00871
R32106 VDD.n1800 VDD.t1116 1.00871
R32107 VDD.n1804 VDD.t3115 1.00871
R32108 VDD.n5695 VDD.t3949 1.00871
R32109 VDD.n5696 VDD.t3586 1.00871
R32110 VDD.n1834 VDD.t1970 1.00871
R32111 VDD.n1837 VDD.t3567 1.00871
R32112 VDD.n1838 VDD.t3247 1.00871
R32113 VDD.n1839 VDD.t921 1.00871
R32114 VDD.n5702 VDD.t749 1.00871
R32115 VDD.n5699 VDD.t4509 1.00871
R32116 VDD.n1835 VDD.t3013 1.00871
R32117 VDD.n10991 VDD.t4497 1.00871
R32118 VDD.n10987 VDD.t4163 1.00871
R32119 VDD.n10984 VDD.t4607 1.00871
R32120 VDD.n5789 VDD.t1599 1.00871
R32121 VDD.n5790 VDD.t1238 1.00871
R32122 VDD.n1843 VDD.t3805 1.00871
R32123 VDD.n10953 VDD.t1230 1.00871
R32124 VDD.n10958 VDD.t897 1.00871
R32125 VDD.n10962 VDD.t2127 1.00871
R32126 VDD.n5796 VDD.t3307 1.00871
R32127 VDD.n5793 VDD.t3009 1.00871
R32128 VDD.n1844 VDD.t1285 1.00871
R32129 VDD.n10954 VDD.t2993 1.00871
R32130 VDD.n10959 VDD.t2620 1.00871
R32131 VDD.n10963 VDD.t1146 1.00871
R32132 VDD.n5682 VDD.t1520 1.00871
R32133 VDD.n5683 VDD.t1174 1.00871
R32134 VDD.n1853 VDD.t3738 1.00871
R32135 VDD.n1856 VDD.t1161 1.00871
R32136 VDD.n1882 VDD.t805 1.00871
R32137 VDD.n1886 VDD.t1440 1.00871
R32138 VDD.n5689 VDD.t2817 1.00871
R32139 VDD.n5686 VDD.t2459 1.00871
R32140 VDD.n1854 VDD.t784 1.00871
R32141 VDD.n1857 VDD.t2446 1.00871
R32142 VDD.n1883 VDD.t1984 1.00871
R32143 VDD.n1887 VDD.t1904 1.00871
R32144 VDD.n5844 VDD.t4105 1.00871
R32145 VDD.n5845 VDD.t3730 1.00871
R32146 VDD.n1899 VDD.t2123 1.00871
R32147 VDD.n1902 VDD.t3718 1.00871
R32148 VDD.n1903 VDD.t3341 1.00871
R32149 VDD.n1904 VDD.t2179 1.00871
R32150 VDD.n5851 VDD.t4539 1.00871
R32151 VDD.n5848 VDD.t4235 1.00871
R32152 VDD.n1900 VDD.t2683 1.00871
R32153 VDD.n10936 VDD.t4225 1.00871
R32154 VDD.n10932 VDD.t3831 1.00871
R32155 VDD.n10929 VDD.t3203 1.00871
R32156 VDD.n5669 VDD.t2142 1.00871
R32157 VDD.n5670 VDD.t1754 1.00871
R32158 VDD.n1908 VDD.t4321 1.00871
R32159 VDD.n10898 VDD.t1739 1.00871
R32160 VDD.n10903 VDD.t1369 1.00871
R32161 VDD.n10907 VDD.t3977 1.00871
R32162 VDD.n5676 VDD.t1603 1.00871
R32163 VDD.n5673 VDD.t1242 1.00871
R32164 VDD.n1909 VDD.t3815 1.00871
R32165 VDD.n10899 VDD.t1232 1.00871
R32166 VDD.n10904 VDD.t909 1.00871
R32167 VDD.n10908 VDD.t2359 1.00871
R32168 VDD.n5877 VDD.t1579 1.00871
R32169 VDD.n5878 VDD.t1226 1.00871
R32170 VDD.n5879 VDD.t3791 1.00871
R32171 VDD.n5491 VDD.t1201 1.00871
R32172 VDD.n5496 VDD.t879 1.00871
R32173 VDD.n5500 VDD.t4711 1.00871
R32174 VDD.n5898 VDD.t3941 1.00871
R32175 VDD.n5895 VDD.t3580 1.00871
R32176 VDD.n5891 VDD.t1960 1.00871
R32177 VDD.n5492 VDD.t3557 1.00871
R32178 VDD.n5497 VDD.t3241 1.00871
R32179 VDD.n5501 VDD.t2116 1.00871
R32180 VDD.n5627 VDD.t1031 1.00871
R32181 VDD.n5628 VDD.t663 1.00871
R32182 VDD.n1926 VDD.t3275 1.00871
R32183 VDD.n1929 VDD.t643 1.00871
R32184 VDD.n1930 VDD.t4413 1.00871
R32185 VDD.n1931 VDD.t4333 1.00871
R32186 VDD.n5634 VDD.t1976 1.00871
R32187 VDD.n5631 VDD.t1607 1.00871
R32188 VDD.n1927 VDD.t4187 1.00871
R32189 VDD.n10881 VDD.t1591 1.00871
R32190 VDD.n10877 VDD.t1213 1.00871
R32191 VDD.n10874 VDD.t3913 1.00871
R32192 VDD.n5606 VDD.t4625 1.00871
R32193 VDD.n5607 VDD.t4289 1.00871
R32194 VDD.n1935 VDD.t2760 1.00871
R32195 VDD.n10843 VDD.t4273 1.00871
R32196 VDD.n10848 VDD.t3897 1.00871
R32197 VDD.n10852 VDD.t959 1.00871
R32198 VDD.n5613 VDD.t2155 1.00871
R32199 VDD.n5610 VDD.t1760 1.00871
R32200 VDD.n1936 VDD.t4325 1.00871
R32201 VDD.n10844 VDD.t1745 1.00871
R32202 VDD.n10849 VDD.t1377 1.00871
R32203 VDD.n10853 VDD.t4145 1.00871
R32204 VDD.n5585 VDD.t2405 1.00871
R32205 VDD.n5586 VDD.t1972 1.00871
R32206 VDD.n1945 VDD.t4489 1.00871
R32207 VDD.n1948 VDD.t1945 1.00871
R32208 VDD.n1974 VDD.t1552 1.00871
R32209 VDD.n1978 VDD.t2183 1.00871
R32210 VDD.n5592 VDD.t3989 1.00871
R32211 VDD.n5589 VDD.t3625 1.00871
R32212 VDD.n1946 VDD.t2013 1.00871
R32213 VDD.n1949 VDD.t3610 1.00871
R32214 VDD.n1975 VDD.t3285 1.00871
R32215 VDD.n1979 VDD.t1184 1.00871
R32216 VDD.n2106 VDD.t2570 1.00871
R32217 VDD.n2111 VDD.t2138 1.00871
R32218 VDD.n1991 VDD.t4667 1.00871
R32219 VDD.n1994 VDD.t2118 1.00871
R32220 VDD.n1995 VDD.t1717 1.00871
R32221 VDD.n1998 VDD.t2472 1.00871
R32222 VDD.n8096 VDD.t3465 1.00871
R32223 VDD.n2114 VDD.t3155 1.00871
R32224 VDD.n1992 VDD.t1443 1.00871
R32225 VDD.n10826 VDD.t3133 1.00871
R32226 VDD.n10822 VDD.t2794 1.00871
R32227 VDD.n1999 VDD.t1957 1.00871
R32228 VDD.n2093 VDD.t1932 1.00871
R32229 VDD.n2094 VDD.t1566 1.00871
R32230 VDD.n2008 VDD.t4153 1.00871
R32231 VDD.n10785 VDD.t1545 1.00871
R32232 VDD.n10790 VDD.t1181 1.00871
R32233 VDD.n10794 VDD.t3205 1.00871
R32234 VDD.n2100 VDD.t1796 1.00871
R32235 VDD.n2097 VDD.t1436 1.00871
R32236 VDD.n2009 VDD.t4029 1.00871
R32237 VDD.n10786 VDD.t1425 1.00871
R32238 VDD.n10791 VDD.t1085 1.00871
R32239 VDD.n10795 VDD.t2744 1.00871
R32240 VDD.n8122 VDD.t4259 1.00871
R32241 VDD.n8123 VDD.t3903 1.00871
R32242 VDD.n2018 VDD.t2353 1.00871
R32243 VDD.n2021 VDD.t3881 1.00871
R32244 VDD.n2029 VDD.t3513 1.00871
R32245 VDD.n2033 VDD.t3039 1.00871
R32246 VDD.n8129 VDD.t1263 1.00871
R32247 VDD.n8126 VDD.t956 1.00871
R32248 VDD.n2019 VDD.t3489 1.00871
R32249 VDD.n2022 VDD.t934 1.00871
R32250 VDD.n2030 VDD.t4685 1.00871
R32251 VDD.n2034 VDD.t3427 1.00871
R32252 VDD.n8166 VDD.t759 1.00871
R32253 VDD.n8181 VDD.t4519 1.00871
R32254 VDD.n8201 VDD.t3021 1.00871
R32255 VDD.n8214 VDD.t4505 1.00871
R32256 VDD.n8236 VDD.t4175 1.00871
R32257 VDD.n8249 VDD.t4185 1.00871
R32258 VDD.n9088 VDD.t3315 1.00871
R32259 VDD.n9089 VDD.t724 1.00871
R32260 VDD.n9086 VDD.t2632 1.00871
R32261 VDD.n9087 VDD.t2979 1.00871
R32262 VDD.n9075 VDD.t2147 1.00871
R32263 VDD.n9076 VDD.t2582 1.00871
R32264 VDD.n8463 VDD.t3167 1.00871
R32265 VDD.n8467 VDD.t2602 1.00871
R32266 VDD.n8468 VDD.t2971 1.00871
R32267 VDD.n8469 VDD.t4465 1.00871
R32268 VDD.n9082 VDD.t2539 1.00871
R32269 VDD.n9079 VDD.t2883 1.00871
R32270 VDD.n8464 VDD.t3441 1.00871
R32271 VDD.n9175 VDD.t2905 1.00871
R32272 VDD.n9171 VDD.t3255 1.00871
R32273 VDD.n9168 VDD.t608 1.00871
R32274 VDD.n8532 VDD.t4283 1.00871
R32275 VDD.n8533 VDD.t4619 1.00871
R32276 VDD.n8534 VDD.t1098 1.00871
R32277 VDD.n8540 VDD.t4645 1.00871
R32278 VDD.n8541 VDD.t902 1.00871
R32279 VDD.n8542 VDD.t2551 1.00871
R32280 VDD.n8578 VDD.t2705 1.00871
R32281 VDD.n8575 VDD.t3049 1.00871
R32282 VDD.n8571 VDD.t3596 1.00871
R32283 VDD.n8568 VDD.t3067 1.00871
R32284 VDD.n8564 VDD.t3384 1.00871
R32285 VDD.n8561 VDD.t814 1.00871
R32286 VDD.n8776 VDD.t2468 1.00871
R32287 VDD.n8777 VDD.t2823 1.00871
R32288 VDD.n8778 VDD.t3362 1.00871
R32289 VDD.n8779 VDD.t2839 1.00871
R32290 VDD.n8780 VDD.t3187 1.00871
R32291 VDD.n8522 VDD.t4709 1.00871
R32292 VDD.n8796 VDD.t3237 1.00871
R32293 VDD.n8793 VDD.t3539 1.00871
R32294 VDD.n8789 VDD.t4171 1.00871
R32295 VDD.n8786 VDD.t3549 1.00871
R32296 VDD.n8782 VDD.t3937 1.00871
R32297 VDD.n8523 VDD.t1337 1.00871
R32298 VDD.n8514 VDD.t2555 1.00871
R32299 VDD.n8850 VDD.t2903 1.00871
R32300 VDD.n8855 VDD.t3461 1.00871
R32301 VDD.n8859 VDD.t2915 1.00871
R32302 VDD.n8864 VDD.t3277 1.00871
R32303 VDD.n8868 VDD.t635 1.00871
R32304 VDD.n8515 VDD.t1019 1.00871
R32305 VDD.n8851 VDD.t1334 1.00871
R32306 VDD.n8856 VDD.t1974 1.00871
R32307 VDD.n8860 VDD.t1355 1.00871
R32308 VDD.n8865 VDD.t1727 1.00871
R32309 VDD.n8869 VDD.t3349 1.00871
R32310 VDD.n8907 VDD.t4251 1.00871
R32311 VDD.n8908 VDD.t4557 1.00871
R32312 VDD.n8909 VDD.t1058 1.00871
R32313 VDD.n8910 VDD.t4581 1.00871
R32314 VDD.n8911 VDD.t846 1.00871
R32315 VDD.n8503 VDD.t2507 1.00871
R32316 VDD.n8927 VDD.t2857 1.00871
R32317 VDD.n8924 VDD.t3185 1.00871
R32318 VDD.n8920 VDD.t3746 1.00871
R32319 VDD.n8917 VDD.t3199 1.00871
R32320 VDD.n8913 VDD.t3531 1.00871
R32321 VDD.n8504 VDD.t983 1.00871
R32322 VDD.n8495 VDD.t2083 1.00871
R32323 VDD.n8977 VDD.t2505 1.00871
R32324 VDD.n8982 VDD.t3101 1.00871
R32325 VDD.n8986 VDD.t2519 1.00871
R32326 VDD.n8991 VDD.t2885 1.00871
R32327 VDD.n8995 VDD.t4385 1.00871
R32328 VDD.n8496 VDD.t2951 1.00871
R32329 VDD.n8978 VDD.t3273 1.00871
R32330 VDD.n8983 VDD.t3833 1.00871
R32331 VDD.n8987 VDD.t3281 1.00871
R32332 VDD.n8992 VDD.t3606 1.00871
R32333 VDD.n8996 VDD.t1046 1.00871
R32334 VDD.n8477 VDD.t2160 1.00871
R32335 VDD.n8478 VDD.t2588 1.00871
R32336 VDD.n8479 VDD.t3177 1.00871
R32337 VDD.n8481 VDD.t2610 1.00871
R32338 VDD.n8482 VDD.t2983 1.00871
R32339 VDD.n8483 VDD.t4469 1.00871
R32340 VDD.n9061 VDD.t2451 1.00871
R32341 VDD.n9058 VDD.t2810 1.00871
R32342 VDD.n9054 VDD.t3337 1.00871
R32343 VDD.n9051 VDD.t2825 1.00871
R32344 VDD.n9047 VDD.t3173 1.00871
R32345 VDD.n9044 VDD.t4695 1.00871
R32346 VDD.n6897 VDD.n6896 0.9995
R32347 VDD.n6984 VDD.n6983 0.9995
R32348 VDD.n6994 VDD.n6993 0.9995
R32349 VDD.n6916 VDD.n6915 0.9995
R32350 VDD.n6936 VDD.n6935 0.9995
R32351 VDD.n6946 VDD.n6945 0.9995
R32352 VDD.n6430 VDD.n6429 0.9995
R32353 VDD.n6532 VDD.n6531 0.9995
R32354 VDD.n6526 VDD.n6525 0.9995
R32355 VDD.n6467 VDD.n6466 0.9995
R32356 VDD.n6492 VDD.n6491 0.9995
R32357 VDD.n6486 VDD.n6485 0.9995
R32358 VDD.n7918 VDD.n7917 0.9995
R32359 VDD.n7927 VDD.n7926 0.9995
R32360 VDD.n7937 VDD.n7936 0.9995
R32361 VDD.n7906 VDD.n7905 0.9995
R32362 VDD.n7900 VDD.n7899 0.9995
R32363 VDD.n7894 VDD.n7893 0.9995
R32364 VDD.n8023 VDD.n8022 0.9995
R32365 VDD.n8032 VDD.n8031 0.9995
R32366 VDD.n8042 VDD.n8041 0.9995
R32367 VDD.n6105 VDD.n6104 0.991625
R32368 VDD.n6062 VDD.n6061 0.991625
R32369 VDD.n6804 VDD.n6803 0.991625
R32370 VDD.n6755 VDD.n6754 0.991625
R32371 VDD.n7024 VDD.n7023 0.983405
R32372 VDD.n7013 VDD.n6877 0.983405
R32373 VDD.n6550 VDD.n6414 0.983405
R32374 VDD.n6561 VDD.n6560 0.983405
R32375 VDD.n7952 VDD.n7951 0.937025
R32376 VDD.n8057 VDD.n8056 0.937025
R32377 VDD.n12633 VDD.n7 0.897031
R32378 VDD.n11872 VDD.n7 0.884663
R32379 VDD.n5539 VDD.n5538 0.851788
R32380 VDD.n6977 VDD.n6976 0.822966
R32381 VDD.n6999 VDD.n6878 0.822966
R32382 VDD.n6536 VDD.n6415 0.822966
R32383 VDD.n6522 VDD.n6521 0.822966
R32384 VDD.n65 VDD.n64 0.805721
R32385 VDD.n154 VDD.n153 0.805721
R32386 VDD.n9109 VDD.n9108 0.805721
R32387 VDD.n8822 VDD.n8821 0.805721
R32388 VDD.n8962 VDD.n8961 0.805721
R32389 VDD.n5765 VDD.n5764 0.805146
R32390 VDD.n5832 VDD.n5831 0.805146
R32391 VDD.n5649 VDD.n5648 0.805146
R32392 VDD.n5567 VDD.n5566 0.805146
R32393 VDD.n8153 VDD.n8152 0.805146
R32394 VDD.n69 VDD.n67 0.803395
R32395 VDD.n158 VDD.n156 0.803395
R32396 VDD.n9113 VDD.n9111 0.803395
R32397 VDD.n8826 VDD.n8824 0.803395
R32398 VDD.n8966 VDD.n8964 0.803395
R32399 VDD.n5768 VDD.n5767 0.80221
R32400 VDD.n5835 VDD.n5834 0.80221
R32401 VDD.n5652 VDD.n5651 0.80221
R32402 VDD.n5570 VDD.n5569 0.80221
R32403 VDD.n8156 VDD.n8155 0.80221
R32404 VDD.n8087 VDD.n8086 0.789456
R32405 VDD.n6156 VDD.n6019 0.737223
R32406 VDD.n6099 VDD.n6092 0.737223
R32407 VDD.n6151 VDD.n6150 0.737223
R32408 VDD.n6074 VDD.n6038 0.737223
R32409 VDD.n6848 VDD.n2405 0.737223
R32410 VDD.n6798 VDD.n6791 0.737223
R32411 VDD.n6841 VDD.n6840 0.737223
R32412 VDD.n6758 VDD.n6728 0.737223
R32413 VDD.n6100 VDD.n6099 0.725061
R32414 VDD.n6117 VDD.n6038 0.725061
R32415 VDD.n6799 VDD.n6798 0.725061
R32416 VDD.n6807 VDD.n6728 0.725061
R32417 VDD.n6328 VDD.n6327 0.699146
R32418 VDD.n6013 VDD.n5988 0.697565
R32419 VDD.n6299 VDD.n5488 0.694506
R32420 VDD.n7923 VDD.n7922 0.66425
R32421 VDD.n7903 VDD.n7902 0.66425
R32422 VDD.n8028 VDD.n8027 0.66425
R32423 VDD.n7023 VDD.n2376 0.639318
R32424 VDD.n6976 VDD.n6959 0.639318
R32425 VDD.n7013 VDD.n7012 0.639318
R32426 VDD.n6951 VDD.n6878 0.639318
R32427 VDD.n6550 VDD.n6549 0.639318
R32428 VDD.n6496 VDD.n6415 0.639318
R32429 VDD.n6560 VDD.n5289 0.639318
R32430 VDD.n6521 VDD.n6504 0.639318
R32431 VDD.n980 VDD.n979 0.636255
R32432 VDD.n1039 VDD.n1038 0.636255
R32433 VDD.n1041 VDD.n735 0.636255
R32434 VDD.n1102 VDD.n784 0.636255
R32435 VDD.n1625 VDD.n1624 0.636255
R32436 VDD.n1091 VDD.n1090 0.636255
R32437 VDD.n1424 VDD.n1423 0.636255
R32438 VDD.n858 VDD.n857 0.636255
R32439 VDD.n1674 VDD.n1673 0.636255
R32440 VDD.n1680 VDD.n1679 0.636255
R32441 VDD.n1686 VDD.n1685 0.636255
R32442 VDD.n1693 VDD.n1692 0.636255
R32443 VDD.n983 VDD.n982 0.63334
R32444 VDD.n1036 VDD.n1034 0.63334
R32445 VDD.n1044 VDD.n1043 0.63334
R32446 VDD.n1105 VDD.n1104 0.63334
R32447 VDD.n1622 VDD.n1620 0.63334
R32448 VDD.n1088 VDD.n1086 0.63334
R32449 VDD.n1421 VDD.n1419 0.63334
R32450 VDD.n855 VDD.n853 0.63334
R32451 VDD.n1677 VDD.n1676 0.63334
R32452 VDD.n1683 VDD.n1682 0.63334
R32453 VDD.n1689 VDD.n1688 0.63334
R32454 VDD.n1696 VDD.n1695 0.63334
R32455 VDD.n982 VDD.n980 0.631515
R32456 VDD.n1038 VDD.n1036 0.631515
R32457 VDD.n1043 VDD.n1041 0.631515
R32458 VDD.n1104 VDD.n1102 0.631515
R32459 VDD.n1624 VDD.n1622 0.631515
R32460 VDD.n1090 VDD.n1088 0.631515
R32461 VDD.n1423 VDD.n1421 0.631515
R32462 VDD.n857 VDD.n855 0.631515
R32463 VDD.n1676 VDD.n1674 0.631515
R32464 VDD.n1682 VDD.n1680 0.631515
R32465 VDD.n1688 VDD.n1686 0.631515
R32466 VDD.n1695 VDD.n1693 0.631515
R32467 VDD.n1742 VDD.t431 0.60727
R32468 VDD.t441 VDD.n1718 0.60727
R32469 VDD.t443 VDD.n1414 0.60727
R32470 VDD.n1356 VDD.t319 0.60727
R32471 VDD.n1349 VDD.t320 0.60727
R32472 VDD.n1652 VDD.t314 0.60727
R32473 VDD.n6977 VDD.n2376 0.585196
R32474 VDD.n7012 VDD.n6999 0.585196
R32475 VDD.n6549 VDD.n6536 0.585196
R32476 VDD.n6522 VDD.n5289 0.585196
R32477 VDD.n6100 VDD.n6019 0.585196
R32478 VDD.n6150 VDD.n6117 0.585196
R32479 VDD.n6799 VDD.n2405 0.585196
R32480 VDD.n6840 VDD.n6807 0.585196
R32481 VDD.n8087 VDD.n2119 0.51351
R32482 VDD.n5912 VDD.n5539 0.48482
R32483 VDD.n8250 VDD.n8249 0.468749
R32484 VDD.n8237 VDD.n8236 0.468749
R32485 VDD.n8215 VDD.n8214 0.468749
R32486 VDD.n8202 VDD.n8201 0.468749
R32487 VDD.n8182 VDD.n8181 0.468749
R32488 VDD.n8167 VDD.n8166 0.468749
R32489 VDD.n2035 VDD.n2034 0.468749
R32490 VDD.n2031 VDD.n2030 0.468749
R32491 VDD.n2023 VDD.n2022 0.468749
R32492 VDD.n2020 VDD.n2019 0.468749
R32493 VDD.n8127 VDD.n8126 0.468749
R32494 VDD.n8130 VDD.n8129 0.468749
R32495 VDD.n2035 VDD.n2033 0.468749
R32496 VDD.n2031 VDD.n2029 0.468749
R32497 VDD.n2023 VDD.n2021 0.468749
R32498 VDD.n2020 VDD.n2018 0.468749
R32499 VDD.n8127 VDD.n8123 0.468749
R32500 VDD.n8130 VDD.n8122 0.468749
R32501 VDD.n10796 VDD.n10795 0.468749
R32502 VDD.n10792 VDD.n10791 0.468749
R32503 VDD.n10787 VDD.n10786 0.468749
R32504 VDD.n2010 VDD.n2009 0.468749
R32505 VDD.n2098 VDD.n2097 0.468749
R32506 VDD.n2101 VDD.n2100 0.468749
R32507 VDD.n10796 VDD.n10794 0.468749
R32508 VDD.n10792 VDD.n10790 0.468749
R32509 VDD.n10787 VDD.n10785 0.468749
R32510 VDD.n2010 VDD.n2008 0.468749
R32511 VDD.n2098 VDD.n2094 0.468749
R32512 VDD.n2101 VDD.n2093 0.468749
R32513 VDD.n2000 VDD.n1999 0.468749
R32514 VDD.n10823 VDD.n10822 0.468749
R32515 VDD.n10827 VDD.n10826 0.468749
R32516 VDD.n1993 VDD.n1992 0.468749
R32517 VDD.n2115 VDD.n2114 0.468749
R32518 VDD.n8097 VDD.n8096 0.468749
R32519 VDD.n2000 VDD.n1998 0.468749
R32520 VDD.n10823 VDD.n1995 0.468749
R32521 VDD.n10827 VDD.n1994 0.468749
R32522 VDD.n1993 VDD.n1991 0.468749
R32523 VDD.n2115 VDD.n2111 0.468749
R32524 VDD.n8097 VDD.n2106 0.468749
R32525 VDD.n1980 VDD.n1979 0.468749
R32526 VDD.n1976 VDD.n1975 0.468749
R32527 VDD.n1950 VDD.n1949 0.468749
R32528 VDD.n1947 VDD.n1946 0.468749
R32529 VDD.n5590 VDD.n5589 0.468749
R32530 VDD.n5593 VDD.n5592 0.468749
R32531 VDD.n1980 VDD.n1978 0.468749
R32532 VDD.n1976 VDD.n1974 0.468749
R32533 VDD.n1950 VDD.n1948 0.468749
R32534 VDD.n1947 VDD.n1945 0.468749
R32535 VDD.n5590 VDD.n5586 0.468749
R32536 VDD.n5593 VDD.n5585 0.468749
R32537 VDD.n10854 VDD.n10853 0.468749
R32538 VDD.n10850 VDD.n10849 0.468749
R32539 VDD.n10845 VDD.n10844 0.468749
R32540 VDD.n1937 VDD.n1936 0.468749
R32541 VDD.n5611 VDD.n5610 0.468749
R32542 VDD.n5614 VDD.n5613 0.468749
R32543 VDD.n10854 VDD.n10852 0.468749
R32544 VDD.n10850 VDD.n10848 0.468749
R32545 VDD.n10845 VDD.n10843 0.468749
R32546 VDD.n1937 VDD.n1935 0.468749
R32547 VDD.n5611 VDD.n5607 0.468749
R32548 VDD.n5614 VDD.n5606 0.468749
R32549 VDD.n10875 VDD.n10874 0.468749
R32550 VDD.n10878 VDD.n10877 0.468749
R32551 VDD.n10882 VDD.n10881 0.468749
R32552 VDD.n1928 VDD.n1927 0.468749
R32553 VDD.n5632 VDD.n5631 0.468749
R32554 VDD.n5635 VDD.n5634 0.468749
R32555 VDD.n10875 VDD.n1931 0.468749
R32556 VDD.n10878 VDD.n1930 0.468749
R32557 VDD.n10882 VDD.n1929 0.468749
R32558 VDD.n1928 VDD.n1926 0.468749
R32559 VDD.n5632 VDD.n5628 0.468749
R32560 VDD.n5635 VDD.n5627 0.468749
R32561 VDD.n5502 VDD.n5501 0.468749
R32562 VDD.n5498 VDD.n5497 0.468749
R32563 VDD.n5493 VDD.n5492 0.468749
R32564 VDD.n5892 VDD.n5891 0.468749
R32565 VDD.n5896 VDD.n5895 0.468749
R32566 VDD.n5899 VDD.n5898 0.468749
R32567 VDD.n5502 VDD.n5500 0.468749
R32568 VDD.n5498 VDD.n5496 0.468749
R32569 VDD.n5493 VDD.n5491 0.468749
R32570 VDD.n5892 VDD.n5879 0.468749
R32571 VDD.n5896 VDD.n5878 0.468749
R32572 VDD.n5899 VDD.n5877 0.468749
R32573 VDD.n10909 VDD.n10908 0.468749
R32574 VDD.n10905 VDD.n10904 0.468749
R32575 VDD.n10900 VDD.n10899 0.468749
R32576 VDD.n1910 VDD.n1909 0.468749
R32577 VDD.n5674 VDD.n5673 0.468749
R32578 VDD.n5677 VDD.n5676 0.468749
R32579 VDD.n10909 VDD.n10907 0.468749
R32580 VDD.n10905 VDD.n10903 0.468749
R32581 VDD.n10900 VDD.n10898 0.468749
R32582 VDD.n1910 VDD.n1908 0.468749
R32583 VDD.n5674 VDD.n5670 0.468749
R32584 VDD.n5677 VDD.n5669 0.468749
R32585 VDD.n10930 VDD.n10929 0.468749
R32586 VDD.n10933 VDD.n10932 0.468749
R32587 VDD.n10937 VDD.n10936 0.468749
R32588 VDD.n1901 VDD.n1900 0.468749
R32589 VDD.n5849 VDD.n5848 0.468749
R32590 VDD.n5852 VDD.n5851 0.468749
R32591 VDD.n10930 VDD.n1904 0.468749
R32592 VDD.n10933 VDD.n1903 0.468749
R32593 VDD.n10937 VDD.n1902 0.468749
R32594 VDD.n1901 VDD.n1899 0.468749
R32595 VDD.n5849 VDD.n5845 0.468749
R32596 VDD.n5852 VDD.n5844 0.468749
R32597 VDD.n1888 VDD.n1887 0.468749
R32598 VDD.n1884 VDD.n1883 0.468749
R32599 VDD.n1858 VDD.n1857 0.468749
R32600 VDD.n1855 VDD.n1854 0.468749
R32601 VDD.n5687 VDD.n5686 0.468749
R32602 VDD.n5690 VDD.n5689 0.468749
R32603 VDD.n1888 VDD.n1886 0.468749
R32604 VDD.n1884 VDD.n1882 0.468749
R32605 VDD.n1858 VDD.n1856 0.468749
R32606 VDD.n1855 VDD.n1853 0.468749
R32607 VDD.n5687 VDD.n5683 0.468749
R32608 VDD.n5690 VDD.n5682 0.468749
R32609 VDD.n10964 VDD.n10963 0.468749
R32610 VDD.n10960 VDD.n10959 0.468749
R32611 VDD.n10955 VDD.n10954 0.468749
R32612 VDD.n1845 VDD.n1844 0.468749
R32613 VDD.n5794 VDD.n5793 0.468749
R32614 VDD.n5797 VDD.n5796 0.468749
R32615 VDD.n10964 VDD.n10962 0.468749
R32616 VDD.n10960 VDD.n10958 0.468749
R32617 VDD.n10955 VDD.n10953 0.468749
R32618 VDD.n1845 VDD.n1843 0.468749
R32619 VDD.n5794 VDD.n5790 0.468749
R32620 VDD.n5797 VDD.n5789 0.468749
R32621 VDD.n10985 VDD.n10984 0.468749
R32622 VDD.n10988 VDD.n10987 0.468749
R32623 VDD.n10992 VDD.n10991 0.468749
R32624 VDD.n1836 VDD.n1835 0.468749
R32625 VDD.n5700 VDD.n5699 0.468749
R32626 VDD.n5703 VDD.n5702 0.468749
R32627 VDD.n10985 VDD.n1839 0.468749
R32628 VDD.n10988 VDD.n1838 0.468749
R32629 VDD.n10992 VDD.n1837 0.468749
R32630 VDD.n1836 VDD.n1834 0.468749
R32631 VDD.n5700 VDD.n5696 0.468749
R32632 VDD.n5703 VDD.n5695 0.468749
R32633 VDD.n1805 VDD.n1804 0.468749
R32634 VDD.n1801 VDD.n1800 0.468749
R32635 VDD.n1793 VDD.n1792 0.468749
R32636 VDD.n1790 VDD.n1789 0.468749
R32637 VDD.n5739 VDD.n5738 0.468749
R32638 VDD.n5742 VDD.n5741 0.468749
R32639 VDD.n1805 VDD.n1803 0.468749
R32640 VDD.n1801 VDD.n1799 0.468749
R32641 VDD.n1793 VDD.n1791 0.468749
R32642 VDD.n1790 VDD.n1788 0.468749
R32643 VDD.n5739 VDD.n5735 0.468749
R32644 VDD.n5742 VDD.n5734 0.468749
R32645 VDD.n11019 VDD.n11018 0.468749
R32646 VDD.n11015 VDD.n11014 0.468749
R32647 VDD.n11010 VDD.n11009 0.468749
R32648 VDD.n1783 VDD.n1782 0.468749
R32649 VDD.n5713 VDD.n5712 0.468749
R32650 VDD.n5716 VDD.n5715 0.468749
R32651 VDD.n11019 VDD.n11017 0.468749
R32652 VDD.n11015 VDD.n11013 0.468749
R32653 VDD.n11010 VDD.n11008 0.468749
R32654 VDD.n1783 VDD.n1781 0.468749
R32655 VDD.n5713 VDD.n5709 0.468749
R32656 VDD.n5716 VDD.n5708 0.468749
R32657 VDD.n642 VDD.n641 0.468749
R32658 VDD.n649 VDD.n648 0.468749
R32659 VDD.n11090 VDD.n11089 0.468749
R32660 VDD.n11077 VDD.n11076 0.468749
R32661 VDD.n11057 VDD.n11056 0.468749
R32662 VDD.n1766 VDD.n1765 0.468749
R32663 VDD.n9045 VDD.n9044 0.468749
R32664 VDD.n9048 VDD.n9047 0.468749
R32665 VDD.n9052 VDD.n9051 0.468749
R32666 VDD.n9055 VDD.n9054 0.468749
R32667 VDD.n9059 VDD.n9058 0.468749
R32668 VDD.n9062 VDD.n9061 0.468749
R32669 VDD.n9045 VDD.n8483 0.468749
R32670 VDD.n9048 VDD.n8482 0.468749
R32671 VDD.n9052 VDD.n8481 0.468749
R32672 VDD.n9055 VDD.n8479 0.468749
R32673 VDD.n9059 VDD.n8478 0.468749
R32674 VDD.n9062 VDD.n8477 0.468749
R32675 VDD.n8997 VDD.n8996 0.468749
R32676 VDD.n8993 VDD.n8992 0.468749
R32677 VDD.n8988 VDD.n8987 0.468749
R32678 VDD.n8984 VDD.n8983 0.468749
R32679 VDD.n8979 VDD.n8978 0.468749
R32680 VDD.n8497 VDD.n8496 0.468749
R32681 VDD.n8997 VDD.n8995 0.468749
R32682 VDD.n8993 VDD.n8991 0.468749
R32683 VDD.n8988 VDD.n8986 0.468749
R32684 VDD.n8984 VDD.n8982 0.468749
R32685 VDD.n8979 VDD.n8977 0.468749
R32686 VDD.n8497 VDD.n8495 0.468749
R32687 VDD.n8505 VDD.n8504 0.468749
R32688 VDD.n8914 VDD.n8913 0.468749
R32689 VDD.n8918 VDD.n8917 0.468749
R32690 VDD.n8921 VDD.n8920 0.468749
R32691 VDD.n8925 VDD.n8924 0.468749
R32692 VDD.n8928 VDD.n8927 0.468749
R32693 VDD.n8505 VDD.n8503 0.468749
R32694 VDD.n8914 VDD.n8911 0.468749
R32695 VDD.n8918 VDD.n8910 0.468749
R32696 VDD.n8921 VDD.n8909 0.468749
R32697 VDD.n8925 VDD.n8908 0.468749
R32698 VDD.n8928 VDD.n8907 0.468749
R32699 VDD.n8870 VDD.n8869 0.468749
R32700 VDD.n8866 VDD.n8865 0.468749
R32701 VDD.n8861 VDD.n8860 0.468749
R32702 VDD.n8857 VDD.n8856 0.468749
R32703 VDD.n8852 VDD.n8851 0.468749
R32704 VDD.n8516 VDD.n8515 0.468749
R32705 VDD.n8870 VDD.n8868 0.468749
R32706 VDD.n8866 VDD.n8864 0.468749
R32707 VDD.n8861 VDD.n8859 0.468749
R32708 VDD.n8857 VDD.n8855 0.468749
R32709 VDD.n8852 VDD.n8850 0.468749
R32710 VDD.n8516 VDD.n8514 0.468749
R32711 VDD.n8524 VDD.n8523 0.468749
R32712 VDD.n8783 VDD.n8782 0.468749
R32713 VDD.n8787 VDD.n8786 0.468749
R32714 VDD.n8790 VDD.n8789 0.468749
R32715 VDD.n8794 VDD.n8793 0.468749
R32716 VDD.n8797 VDD.n8796 0.468749
R32717 VDD.n8524 VDD.n8522 0.468749
R32718 VDD.n8783 VDD.n8780 0.468749
R32719 VDD.n8787 VDD.n8779 0.468749
R32720 VDD.n8790 VDD.n8778 0.468749
R32721 VDD.n8794 VDD.n8777 0.468749
R32722 VDD.n8797 VDD.n8776 0.468749
R32723 VDD.n8562 VDD.n8561 0.468749
R32724 VDD.n8565 VDD.n8564 0.468749
R32725 VDD.n8569 VDD.n8568 0.468749
R32726 VDD.n8572 VDD.n8571 0.468749
R32727 VDD.n8576 VDD.n8575 0.468749
R32728 VDD.n8579 VDD.n8578 0.468749
R32729 VDD.n8562 VDD.n8542 0.468749
R32730 VDD.n8565 VDD.n8541 0.468749
R32731 VDD.n8569 VDD.n8540 0.468749
R32732 VDD.n8572 VDD.n8534 0.468749
R32733 VDD.n8576 VDD.n8533 0.468749
R32734 VDD.n8579 VDD.n8532 0.468749
R32735 VDD.n9169 VDD.n9168 0.468749
R32736 VDD.n9172 VDD.n9171 0.468749
R32737 VDD.n9176 VDD.n9175 0.468749
R32738 VDD.n8465 VDD.n8464 0.468749
R32739 VDD.n9080 VDD.n9079 0.468749
R32740 VDD.n9083 VDD.n9082 0.468749
R32741 VDD.n9169 VDD.n8469 0.468749
R32742 VDD.n9172 VDD.n8468 0.468749
R32743 VDD.n9176 VDD.n8467 0.468749
R32744 VDD.n8465 VDD.n8463 0.468749
R32745 VDD.n9080 VDD.n9076 0.468749
R32746 VDD.n9083 VDD.n9075 0.468749
R32747 VDD.n9136 VDD.n9087 0.468749
R32748 VDD.n9138 VDD.n9086 0.468749
R32749 VDD.n9124 VDD.n9089 0.468749
R32750 VDD.n9126 VDD.n9088 0.468749
R32751 VDD.n12451 VDD.n12450 0.468749
R32752 VDD.n12454 VDD.n12453 0.468749
R32753 VDD.n12458 VDD.n12457 0.468749
R32754 VDD.n180 VDD.n179 0.468749
R32755 VDD.n8588 VDD.n8587 0.468749
R32756 VDD.n8591 VDD.n8590 0.468749
R32757 VDD.n12451 VDD.n183 0.468749
R32758 VDD.n12454 VDD.n182 0.468749
R32759 VDD.n12458 VDD.n181 0.468749
R32760 VDD.n180 VDD.n178 0.468749
R32761 VDD.n8588 VDD.n8584 0.468749
R32762 VDD.n8591 VDD.n8583 0.468749
R32763 VDD.n134 VDD.n133 0.468749
R32764 VDD.n130 VDD.n129 0.468749
R32765 VDD.n122 VDD.n121 0.468749
R32766 VDD.n119 VDD.n118 0.468749
R32767 VDD.n8731 VDD.n8730 0.468749
R32768 VDD.n8734 VDD.n8733 0.468749
R32769 VDD.n134 VDD.n132 0.468749
R32770 VDD.n130 VDD.n128 0.468749
R32771 VDD.n122 VDD.n120 0.468749
R32772 VDD.n119 VDD.n117 0.468749
R32773 VDD.n8731 VDD.n8727 0.468749
R32774 VDD.n8734 VDD.n8726 0.468749
R32775 VDD.n12486 VDD.n12485 0.468749
R32776 VDD.n12482 VDD.n12481 0.468749
R32777 VDD.n12477 VDD.n12476 0.468749
R32778 VDD.n109 VDD.n108 0.468749
R32779 VDD.n8601 VDD.n8600 0.468749
R32780 VDD.n8604 VDD.n8603 0.468749
R32781 VDD.n12486 VDD.n12484 0.468749
R32782 VDD.n12482 VDD.n12480 0.468749
R32783 VDD.n12477 VDD.n12475 0.468749
R32784 VDD.n109 VDD.n107 0.468749
R32785 VDD.n8601 VDD.n8597 0.468749
R32786 VDD.n8604 VDD.n8596 0.468749
R32787 VDD.n12507 VDD.n12506 0.468749
R32788 VDD.n12510 VDD.n12509 0.468749
R32789 VDD.n12514 VDD.n12513 0.468749
R32790 VDD.n100 VDD.n99 0.468749
R32791 VDD.n8693 VDD.n8692 0.468749
R32792 VDD.n8696 VDD.n8695 0.468749
R32793 VDD.n12507 VDD.n103 0.468749
R32794 VDD.n12510 VDD.n102 0.468749
R32795 VDD.n12514 VDD.n101 0.468749
R32796 VDD.n100 VDD.n98 0.468749
R32797 VDD.n8693 VDD.n8689 0.468749
R32798 VDD.n8696 VDD.n8688 0.468749
R32799 VDD.n88 VDD.n87 0.468749
R32800 VDD.n84 VDD.n83 0.468749
R32801 VDD.n42 VDD.n41 0.468749
R32802 VDD.n39 VDD.n38 0.468749
R32803 VDD.n8615 VDD.n8614 0.468749
R32804 VDD.n8618 VDD.n8617 0.468749
R32805 VDD.n88 VDD.n86 0.468749
R32806 VDD.n84 VDD.n82 0.468749
R32807 VDD.n42 VDD.n40 0.468749
R32808 VDD.n39 VDD.n37 0.468749
R32809 VDD.n8615 VDD.n8611 0.468749
R32810 VDD.n8618 VDD.n8610 0.468749
R32811 VDD.n12542 VDD.n12541 0.468749
R32812 VDD.n12538 VDD.n12537 0.468749
R32813 VDD.n12533 VDD.n12532 0.468749
R32814 VDD.n29 VDD.n28 0.468749
R32815 VDD.n8660 VDD.n8659 0.468749
R32816 VDD.n8663 VDD.n8662 0.468749
R32817 VDD.n12542 VDD.n12540 0.468749
R32818 VDD.n12538 VDD.n12536 0.468749
R32819 VDD.n12533 VDD.n12531 0.468749
R32820 VDD.n29 VDD.n27 0.468749
R32821 VDD.n8660 VDD.n8656 0.468749
R32822 VDD.n8663 VDD.n8655 0.468749
R32823 VDD.n12601 VDD.n12600 0.468749
R32824 VDD.n12604 VDD.n12603 0.468749
R32825 VDD.n12608 VDD.n12607 0.468749
R32826 VDD.n20 VDD.n19 0.468749
R32827 VDD.n8629 VDD.n8628 0.468749
R32828 VDD.n8632 VDD.n8631 0.468749
R32829 VDD.n12601 VDD.n23 0.468749
R32830 VDD.n12604 VDD.n22 0.468749
R32831 VDD.n12608 VDD.n21 0.468749
R32832 VDD.n20 VDD.n18 0.468749
R32833 VDD.n8629 VDD.n8625 0.468749
R32834 VDD.n8632 VDD.n8624 0.468749
R32835 VDD.n12558 VDD.n12557 0.468749
R32836 VDD.n12576 VDD.n12575 0.468749
R32837 VDD.n12572 VDD.n12571 0.468749
R32838 VDD.n12569 VDD.n12568 0.468749
R32839 VDD.n12565 VDD.n12564 0.468749
R32840 VDD.n12625 VDD.n12624 0.468749
R32841 VDD.n71 VDD.n62 0.3755
R32842 VDD.n160 VDD.n151 0.3755
R32843 VDD.n5770 VDD.n5761 0.3755
R32844 VDD.n5837 VDD.n5828 0.3755
R32845 VDD.n5654 VDD.n5645 0.3755
R32846 VDD.n5572 VDD.n5563 0.3755
R32847 VDD.n8158 VDD.n8149 0.3755
R32848 VDD.n5912 VDD.n5911 0.3755
R32849 VDD.n5886 VDD.n5539 0.3755
R32850 VDD.n6326 VDD.n6325 0.3755
R32851 VDD.n8090 VDD.n8089 0.3755
R32852 VDD.n9115 VDD.n9106 0.3755
R32853 VDD.n8828 VDD.n8819 0.3755
R32854 VDD.n8968 VDD.n8959 0.3755
R32855 VDD.n1000 VDD.n6 0.3755
R32856 VDD.n12635 VDD.n12634 0.3755
R32857 VDD.n12633 VDD.n12632 0.3755
R32858 VDD.n12579 VDD.n7 0.3755
R32859 VDD.n1762 VDD.n638 0.3755
R32860 VDD.n1761 VDD.n1760 0.3755
R32861 VDD.n6713 VDD.n2409 0.355763
R32862 VDD.n6713 VDD.n2410 0.281286
R32863 VDD.n1556 VDD.n1555 0.249951
R32864 VDD.n1557 VDD.n1556 0.249951
R32865 VDD.n7022 VDD.n2383 0.236091
R32866 VDD.n6975 VDD.n6966 0.236091
R32867 VDD.n6551 VDD.n5296 0.236091
R32868 VDD.n6512 VDD.n6511 0.236091
R32869 VDD.n1555 VDD.n1554 0.192465
R32870 VDD.n1558 VDD.n1557 0.192465
R32871 VDD.n6713 VDD.n2408 0.177356
R32872 VDD.n1442 VDD.n1441 0.174614
R32873 VDD.n1610 VDD.n804 0.174614
R32874 VDD.n1610 VDD.n803 0.174614
R32875 VDD.n1480 VDD.n814 0.174614
R32876 VDD.n1480 VDD.n1479 0.174614
R32877 VDD.n2136 VDD.n2123 0.166289
R32878 VDD.n2162 VDD.n2124 0.166289
R32879 VDD.n2354 VDD.n2124 0.166289
R32880 VDD.n61 VDD.n58 0.157683
R32881 VDD.n70 VDD.n63 0.157683
R32882 VDD.n150 VDD.n147 0.157683
R32883 VDD.n159 VDD.n152 0.157683
R32884 VDD.n5769 VDD.n5762 0.157683
R32885 VDD.n5760 VDD.n5757 0.157683
R32886 VDD.n5836 VDD.n5829 0.157683
R32887 VDD.n5827 VDD.n5824 0.157683
R32888 VDD.n5653 VDD.n5646 0.157683
R32889 VDD.n5644 VDD.n5641 0.157683
R32890 VDD.n5571 VDD.n5564 0.157683
R32891 VDD.n5562 VDD.n5559 0.157683
R32892 VDD.n8157 VDD.n8150 0.157683
R32893 VDD.n8148 VDD.n8145 0.157683
R32894 VDD.n9105 VDD.n9102 0.157683
R32895 VDD.n9114 VDD.n9107 0.157683
R32896 VDD.n8818 VDD.n8815 0.157683
R32897 VDD.n8827 VDD.n8820 0.157683
R32898 VDD.n8958 VDD.n8955 0.157683
R32899 VDD.n8967 VDD.n8960 0.157683
R32900 VDD.n6149 VDD.n6148 0.150184
R32901 VDD.n6075 VDD.n6056 0.150184
R32902 VDD.n6823 VDD.n6822 0.150184
R32903 VDD.n6790 VDD.n6789 0.150184
R32904 VDD.n12449 VDD.n12448 0.143306
R32905 VDD.n6887 VDD.n6885 0.14
R32906 VDD.n6891 VDD.n6885 0.14
R32907 VDD.n6892 VDD.n6884 0.14
R32908 VDD.n6896 VDD.n6884 0.14
R32909 VDD.n6897 VDD.n6883 0.14
R32910 VDD.n6901 VDD.n6883 0.14
R32911 VDD.n6979 VDD.n6882 0.14
R32912 VDD.n6983 VDD.n6882 0.14
R32913 VDD.n6984 VDD.n6881 0.14
R32914 VDD.n6988 VDD.n6881 0.14
R32915 VDD.n6989 VDD.n6880 0.14
R32916 VDD.n6993 VDD.n6880 0.14
R32917 VDD.n6994 VDD.n6879 0.14
R32918 VDD.n6998 VDD.n6879 0.14
R32919 VDD.n6906 VDD.n6904 0.14
R32920 VDD.n6910 VDD.n6904 0.14
R32921 VDD.n6911 VDD.n6903 0.14
R32922 VDD.n6915 VDD.n6903 0.14
R32923 VDD.n6916 VDD.n6902 0.14
R32924 VDD.n6920 VDD.n6902 0.14
R32925 VDD.n6931 VDD.n6930 0.14
R32926 VDD.n6935 VDD.n6930 0.14
R32927 VDD.n6936 VDD.n6929 0.14
R32928 VDD.n6940 VDD.n6929 0.14
R32929 VDD.n6941 VDD.n6928 0.14
R32930 VDD.n6945 VDD.n6928 0.14
R32931 VDD.n6946 VDD.n6927 0.14
R32932 VDD.n6950 VDD.n6927 0.14
R32933 VDD.n6420 VDD.n6418 0.14
R32934 VDD.n6424 VDD.n6418 0.14
R32935 VDD.n6425 VDD.n6417 0.14
R32936 VDD.n6429 VDD.n6417 0.14
R32937 VDD.n6430 VDD.n6416 0.14
R32938 VDD.n6434 VDD.n6416 0.14
R32939 VDD.n6534 VDD.n6435 0.14
R32940 VDD.n6532 VDD.n6435 0.14
R32941 VDD.n6531 VDD.n6438 0.14
R32942 VDD.n6529 VDD.n6438 0.14
R32943 VDD.n6528 VDD.n6441 0.14
R32944 VDD.n6526 VDD.n6441 0.14
R32945 VDD.n6525 VDD.n6444 0.14
R32946 VDD.n6523 VDD.n6444 0.14
R32947 VDD.n6457 VDD.n6455 0.14
R32948 VDD.n6461 VDD.n6455 0.14
R32949 VDD.n6462 VDD.n6454 0.14
R32950 VDD.n6466 VDD.n6454 0.14
R32951 VDD.n6467 VDD.n6453 0.14
R32952 VDD.n6471 VDD.n6453 0.14
R32953 VDD.n6494 VDD.n6472 0.14
R32954 VDD.n6492 VDD.n6472 0.14
R32955 VDD.n6491 VDD.n6475 0.14
R32956 VDD.n6489 VDD.n6475 0.14
R32957 VDD.n6488 VDD.n6478 0.14
R32958 VDD.n6486 VDD.n6478 0.14
R32959 VDD.n6485 VDD.n6481 0.14
R32960 VDD.n6481 VDD.n6447 0.14
R32961 VDD.n6101 VDD.n6040 0.14
R32962 VDD.n6104 VDD.n6040 0.14
R32963 VDD.n6105 VDD.n6039 0.14
R32964 VDD.n6109 VDD.n6039 0.14
R32965 VDD.n6115 VDD.n6110 0.14
R32966 VDD.n6113 VDD.n6110 0.14
R32967 VDD.n6058 VDD.n6041 0.14
R32968 VDD.n6061 VDD.n6058 0.14
R32969 VDD.n6062 VDD.n6057 0.14
R32970 VDD.n6066 VDD.n6057 0.14
R32971 VDD.n6072 VDD.n6067 0.14
R32972 VDD.n6070 VDD.n6067 0.14
R32973 VDD.n7913 VDD.n7860 0.14
R32974 VDD.n7917 VDD.n7860 0.14
R32975 VDD.n7918 VDD.n7859 0.14
R32976 VDD.n7922 VDD.n7859 0.14
R32977 VDD.n7923 VDD.n7858 0.14
R32978 VDD.n7926 VDD.n7858 0.14
R32979 VDD.n7927 VDD.n7857 0.14
R32980 VDD.n7931 VDD.n7857 0.14
R32981 VDD.n7932 VDD.n7856 0.14
R32982 VDD.n7936 VDD.n7856 0.14
R32983 VDD.n7937 VDD.n7855 0.14
R32984 VDD.n7941 VDD.n7855 0.14
R32985 VDD.n7908 VDD.n7865 0.14
R32986 VDD.n7906 VDD.n7865 0.14
R32987 VDD.n7905 VDD.n7869 0.14
R32988 VDD.n7903 VDD.n7869 0.14
R32989 VDD.n7902 VDD.n7873 0.14
R32990 VDD.n7900 VDD.n7873 0.14
R32991 VDD.n7899 VDD.n7875 0.14
R32992 VDD.n7897 VDD.n7875 0.14
R32993 VDD.n7896 VDD.n7879 0.14
R32994 VDD.n7894 VDD.n7879 0.14
R32995 VDD.n7893 VDD.n7883 0.14
R32996 VDD.n7891 VDD.n7883 0.14
R32997 VDD.n8018 VDD.n2155 0.14
R32998 VDD.n8022 VDD.n2155 0.14
R32999 VDD.n8023 VDD.n2154 0.14
R33000 VDD.n8027 VDD.n2154 0.14
R33001 VDD.n8028 VDD.n2153 0.14
R33002 VDD.n8031 VDD.n2153 0.14
R33003 VDD.n8032 VDD.n2152 0.14
R33004 VDD.n8036 VDD.n2152 0.14
R33005 VDD.n8037 VDD.n2151 0.14
R33006 VDD.n8041 VDD.n2151 0.14
R33007 VDD.n8042 VDD.n2150 0.14
R33008 VDD.n8046 VDD.n2150 0.14
R33009 VDD.n6806 VDD.n6729 0.14
R33010 VDD.n6804 VDD.n6729 0.14
R33011 VDD.n6803 VDD.n6731 0.14
R33012 VDD.n6801 VDD.n6731 0.14
R33013 VDD.n6739 VDD.n6734 0.14
R33014 VDD.n6737 VDD.n6734 0.14
R33015 VDD.n6757 VDD.n6747 0.14
R33016 VDD.n6755 VDD.n6747 0.14
R33017 VDD.n6754 VDD.n6749 0.14
R33018 VDD.n6752 VDD.n6749 0.14
R33019 VDD.n6745 VDD.n6740 0.14
R33020 VDD.n6743 VDD.n6740 0.14
R33021 VDD.n6714 VDD.n6713 0.136679
R33022 VDD.n8076 VDD.n8075 0.13175
R33023 VDD.n8077 VDD.n8076 0.13175
R33024 VDD.n8079 VDD.n8078 0.13175
R33025 VDD.n8078 VDD.n8077 0.13175
R33026 VDD.n1549 VDD.n1548 0.119368
R33027 VDD.n1521 VDD.n1520 0.119368
R33028 VDD.n4906 VDD.n4697 0.110375
R33029 VDD.n4905 VDD.n4904 0.110375
R33030 VDD.n3630 VDD.n3629 0.11
R33031 VDD.n3628 VDD.n2745 0.11
R33032 VDD.n10103 VDD.n10102 0.11
R33033 VDD.n10101 VDD.n9214 0.11
R33034 VDD.n11813 VDD.n405 0.109625
R33035 VDD.n11812 VDD.n11811 0.109625
R33036 VDD.n1390 VDD.n1389 0.109121
R33037 VDD.n1414 VDD.n1390 0.109121
R33038 VDD.n1358 VDD.n1357 0.109121
R33039 VDD.n1357 VDD.n1356 0.109121
R33040 VDD.n1343 VDD.n1342 0.109121
R33041 VDD.n1349 VDD.n1343 0.109121
R33042 VDD.n1654 VDD.n1653 0.109121
R33043 VDD.n1653 VDD.n1652 0.109121
R33044 VDD.n1170 VDD.n707 0.109121
R33045 VDD.n1718 VDD.n707 0.109121
R33046 VDD.n1183 VDD.n845 0.109121
R33047 VDD.n1414 VDD.n845 0.109121
R33048 VDD.n1651 VDD.n1650 0.109121
R33049 VDD.n1652 VDD.n1651 0.109121
R33050 VDD.n1600 VDD.n761 0.109121
R33051 VDD.n1652 VDD.n761 0.109121
R33052 VDD.n1600 VDD.n760 0.109121
R33053 VDD.n1652 VDD.n760 0.109121
R33054 VDD.n1276 VDD.n1275 0.109121
R33055 VDD.n1349 VDD.n1276 0.109121
R33056 VDD.n1213 VDD.n849 0.109121
R33057 VDD.n1356 VDD.n849 0.109121
R33058 VDD.n1413 VDD.n1412 0.109121
R33059 VDD.n1414 VDD.n1413 0.109121
R33060 VDD.n1355 VDD.n818 0.109121
R33061 VDD.n1356 VDD.n1355 0.109121
R33062 VDD.n1348 VDD.n808 0.109121
R33063 VDD.n1349 VDD.n1348 0.109121
R33064 VDD.n1412 VDD.n846 0.109121
R33065 VDD.n1414 VDD.n846 0.109121
R33066 VDD.n850 VDD.n818 0.109121
R33067 VDD.n1356 VDD.n850 0.109121
R33068 VDD.n1350 VDD.n808 0.109121
R33069 VDD.n1350 VDD.n1349 0.109121
R33070 VDD.n1066 VDD.n711 0.109121
R33071 VDD.n1718 VDD.n711 0.109121
R33072 VDD.n911 VDD.n689 0.109121
R33073 VDD.n1742 VDD.n689 0.109121
R33074 VDD.n1741 VDD.n1740 0.109121
R33075 VDD.n1742 VDD.n1741 0.109121
R33076 VDD.n1740 VDD.n688 0.109121
R33077 VDD.n1742 VDD.n688 0.109121
R33078 VDD.n1717 VDD.n1716 0.109121
R33079 VDD.n1718 VDD.n1717 0.109121
R33080 VDD.n1716 VDD.n708 0.109121
R33081 VDD.n1718 VDD.n708 0.109121
R33082 VDD.n1744 VDD.n1743 0.109121
R33083 VDD.n1743 VDD.n1742 0.109121
R33084 VDD.n2074 VDD.n2025 0.10728
R33085 VDD.n8137 VDD.n2024 0.10728
R33086 VDD.n10773 VDD.n2024 0.10728
R33087 VDD.n8116 VDD.n2012 0.10728
R33088 VDD.n10781 VDD.n2012 0.10728
R33089 VDD.n10778 VDD.n10777 0.10728
R33090 VDD.n10779 VDD.n10778 0.10728
R33091 VDD.n10777 VDD.n10776 0.10728
R33092 VDD.n10776 VDD.n2017 0.10728
R33093 VDD.n10784 VDD.n2011 0.10728
R33094 VDD.n2016 VDD.n2011 0.10728
R33095 VDD.n10784 VDD.n10783 0.10728
R33096 VDD.n10783 VDD.n10782 0.10728
R33097 VDD.n8104 VDD.n1989 0.10728
R33098 VDD.n2014 VDD.n1989 0.10728
R33099 VDD.n5579 VDD.n1951 0.10728
R33100 VDD.n1988 VDD.n1951 0.10728
R33101 VDD.n10828 VDD.n1952 0.10728
R33102 VDD.n10831 VDD.n1952 0.10728
R33103 VDD.n10829 VDD.n10828 0.10728
R33104 VDD.n10830 VDD.n10829 0.10728
R33105 VDD.n10836 VDD.n10835 0.10728
R33106 VDD.n10837 VDD.n10836 0.10728
R33107 VDD.n10835 VDD.n10834 0.10728
R33108 VDD.n10834 VDD.n1944 0.10728
R33109 VDD.n5600 VDD.n1939 0.10728
R33110 VDD.n10839 VDD.n1939 0.10728
R33111 VDD.n5621 VDD.n1924 0.10728
R33112 VDD.n1941 VDD.n1924 0.10728
R33113 VDD.n10842 VDD.n1938 0.10728
R33114 VDD.n1943 VDD.n1938 0.10728
R33115 VDD.n10842 VDD.n10841 0.10728
R33116 VDD.n10841 VDD.n10840 0.10728
R33117 VDD.n10883 VDD.n1921 0.10728
R33118 VDD.n10886 VDD.n1921 0.10728
R33119 VDD.n10884 VDD.n10883 0.10728
R33120 VDD.n10885 VDD.n10884 0.10728
R33121 VDD.n5661 VDD.n1920 0.10728
R33122 VDD.n1923 VDD.n1920 0.10728
R33123 VDD.n5871 VDD.n1912 0.10728
R33124 VDD.n10894 VDD.n1912 0.10728
R33125 VDD.n10891 VDD.n10890 0.10728
R33126 VDD.n10892 VDD.n10891 0.10728
R33127 VDD.n10890 VDD.n10889 0.10728
R33128 VDD.n10889 VDD.n1917 0.10728
R33129 VDD.n10897 VDD.n1911 0.10728
R33130 VDD.n1916 VDD.n1911 0.10728
R33131 VDD.n10897 VDD.n10896 0.10728
R33132 VDD.n10896 VDD.n10895 0.10728
R33133 VDD.n5859 VDD.n1897 0.10728
R33134 VDD.n1914 VDD.n1897 0.10728
R33135 VDD.n5816 VDD.n1859 0.10728
R33136 VDD.n1896 VDD.n1859 0.10728
R33137 VDD.n10938 VDD.n1860 0.10728
R33138 VDD.n10941 VDD.n1860 0.10728
R33139 VDD.n10939 VDD.n10938 0.10728
R33140 VDD.n10940 VDD.n10939 0.10728
R33141 VDD.n10946 VDD.n10945 0.10728
R33142 VDD.n10947 VDD.n10946 0.10728
R33143 VDD.n10945 VDD.n10944 0.10728
R33144 VDD.n10944 VDD.n1852 0.10728
R33145 VDD.n5804 VDD.n1847 0.10728
R33146 VDD.n10949 VDD.n1847 0.10728
R33147 VDD.n5783 VDD.n1832 0.10728
R33148 VDD.n1849 VDD.n1832 0.10728
R33149 VDD.n10952 VDD.n1846 0.10728
R33150 VDD.n1851 VDD.n1846 0.10728
R33151 VDD.n10952 VDD.n10951 0.10728
R33152 VDD.n10951 VDD.n10950 0.10728
R33153 VDD.n10993 VDD.n1795 0.10728
R33154 VDD.n10996 VDD.n1795 0.10728
R33155 VDD.n10994 VDD.n10993 0.10728
R33156 VDD.n10995 VDD.n10994 0.10728
R33157 VDD.n5749 VDD.n1794 0.10728
R33158 VDD.n1831 VDD.n1794 0.10728
R33159 VDD.n5728 VDD.n1784 0.10728
R33160 VDD.n11004 VDD.n1784 0.10728
R33161 VDD.n11001 VDD.n11000 0.10728
R33162 VDD.n11002 VDD.n11001 0.10728
R33163 VDD.n11000 VDD.n10999 0.10728
R33164 VDD.n10999 VDD.n1787 0.10728
R33165 VDD.n11007 VDD.n1772 0.10728
R33166 VDD.n1786 VDD.n1772 0.10728
R33167 VDD.n11007 VDD.n11006 0.10728
R33168 VDD.n11006 VDD.n11005 0.10728
R33169 VDD.n11031 VDD.n11030 0.10728
R33170 VDD.n11030 VDD.n11029 0.10728
R33171 VDD.n1771 VDD.n657 0.10728
R33172 VDD.n12465 VDD.n175 0.10728
R33173 VDD.n12465 VDD.n12464 0.10728
R33174 VDD.n8570 VDD.n8539 0.10728
R33175 VDD.n8539 VDD.n8538 0.10728
R33176 VDD.n8554 VDD.n177 0.10728
R33177 VDD.n8535 VDD.n177 0.10728
R33178 VDD.n8570 VDD.n8527 0.10728
R33179 VDD.n8537 VDD.n8527 0.10728
R33180 VDD.n8788 VDD.n8528 0.10728
R33181 VDD.n8530 VDD.n8528 0.10728
R33182 VDD.n8809 VDD.n8808 0.10728
R33183 VDD.n8808 VDD.n8807 0.10728
R33184 VDD.n8788 VDD.n8519 0.10728
R33185 VDD.n8529 VDD.n8519 0.10728
R33186 VDD.n8858 VDD.n8520 0.10728
R33187 VDD.n8881 VDD.n8520 0.10728
R33188 VDD.n8878 VDD.n8877 0.10728
R33189 VDD.n8879 VDD.n8878 0.10728
R33190 VDD.n8858 VDD.n8508 0.10728
R33191 VDD.n8880 VDD.n8508 0.10728
R33192 VDD.n8919 VDD.n8509 0.10728
R33193 VDD.n8511 VDD.n8509 0.10728
R33194 VDD.n8940 VDD.n8939 0.10728
R33195 VDD.n8939 VDD.n8938 0.10728
R33196 VDD.n8919 VDD.n8500 0.10728
R33197 VDD.n8510 VDD.n8500 0.10728
R33198 VDD.n8985 VDD.n8501 0.10728
R33199 VDD.n9012 VDD.n8501 0.10728
R33200 VDD.n9009 VDD.n9008 0.10728
R33201 VDD.n9010 VDD.n9009 0.10728
R33202 VDD.n8985 VDD.n8491 0.10728
R33203 VDD.n9011 VDD.n8491 0.10728
R33204 VDD.n9053 VDD.n8480 0.10728
R33205 VDD.n8493 VDD.n8480 0.10728
R33206 VDD.n9037 VDD.n9036 0.10728
R33207 VDD.n9036 VDD.n9035 0.10728
R33208 VDD.n9053 VDD.n8473 0.10728
R33209 VDD.n8492 VDD.n8473 0.10728
R33210 VDD.n9096 VDD.n8461 0.10728
R33211 VDD.n9180 VDD.n8461 0.10728
R33212 VDD.n9161 VDD.n9160 0.10728
R33213 VDD.n9160 VDD.n9159 0.10728
R33214 VDD.n9177 VDD.n8466 0.10728
R33215 VDD.n8466 VDD.n8462 0.10728
R33216 VDD.n9178 VDD.n9177 0.10728
R33217 VDD.n9179 VDD.n9178 0.10728
R33218 VDD.n9183 VDD.n9182 0.10728
R33219 VDD.n12459 VDD.n124 0.10728
R33220 VDD.n12462 VDD.n124 0.10728
R33221 VDD.n12460 VDD.n12459 0.10728
R33222 VDD.n12461 VDD.n12460 0.10728
R33223 VDD.n12468 VDD.n12467 0.10728
R33224 VDD.n12469 VDD.n12468 0.10728
R33225 VDD.n12467 VDD.n12466 0.10728
R33226 VDD.n12466 VDD.n116 0.10728
R33227 VDD.n141 VDD.n112 0.10728
R33228 VDD.n12471 VDD.n112 0.10728
R33229 VDD.n12493 VDD.n97 0.10728
R33230 VDD.n113 VDD.n97 0.10728
R33231 VDD.n12474 VDD.n110 0.10728
R33232 VDD.n115 VDD.n110 0.10728
R33233 VDD.n12474 VDD.n12473 0.10728
R33234 VDD.n12473 VDD.n12472 0.10728
R33235 VDD.n12515 VDD.n44 0.10728
R33236 VDD.n12518 VDD.n44 0.10728
R33237 VDD.n12516 VDD.n12515 0.10728
R33238 VDD.n12517 VDD.n12516 0.10728
R33239 VDD.n12521 VDD.n95 0.10728
R33240 VDD.n12521 VDD.n12520 0.10728
R33241 VDD.n52 VDD.n32 0.10728
R33242 VDD.n12527 VDD.n32 0.10728
R33243 VDD.n12524 VDD.n12523 0.10728
R33244 VDD.n12525 VDD.n12524 0.10728
R33245 VDD.n12523 VDD.n12522 0.10728
R33246 VDD.n12522 VDD.n36 0.10728
R33247 VDD.n12530 VDD.n30 0.10728
R33248 VDD.n35 VDD.n30 0.10728
R33249 VDD.n12530 VDD.n12529 0.10728
R33250 VDD.n12529 VDD.n12528 0.10728
R33251 VDD.n12549 VDD.n17 0.10728
R33252 VDD.n33 VDD.n17 0.10728
R33253 VDD.n12593 VDD.n12592 0.10728
R33254 VDD.n12592 VDD.n15 0.10728
R33255 VDD.n12609 VDD.n14 0.10728
R33256 VDD.n12612 VDD.n14 0.10728
R33257 VDD.n12610 VDD.n12609 0.10728
R33258 VDD.n12611 VDD.n12610 0.10728
R33259 VDD.n12570 VDD.n13 0.10728
R33260 VDD.n7841 VDD.n7840 0.105779
R33261 VDD.n2389 VDD.n2388 0.105779
R33262 VDD.n10775 VDD.n10772 0.1055
R33263 VDD.n10775 VDD.n10774 0.1055
R33264 VDD.n2048 VDD.n2013 0.1055
R33265 VDD.n10780 VDD.n2013 0.1055
R33266 VDD.n10803 VDD.n1990 0.1055
R33267 VDD.n2015 VDD.n1990 0.1055
R33268 VDD.n10833 VDD.n1987 0.1055
R33269 VDD.n10833 VDD.n10832 0.1055
R33270 VDD.n1966 VDD.n1940 0.1055
R33271 VDD.n10838 VDD.n1940 0.1055
R33272 VDD.n10861 VDD.n1925 0.1055
R33273 VDD.n1942 VDD.n1925 0.1055
R33274 VDD.n10888 VDD.n1922 0.1055
R33275 VDD.n10888 VDD.n10887 0.1055
R33276 VDD.n5522 VDD.n1913 0.1055
R33277 VDD.n10893 VDD.n1913 0.1055
R33278 VDD.n10916 VDD.n1898 0.1055
R33279 VDD.n1915 VDD.n1898 0.1055
R33280 VDD.n10943 VDD.n1895 0.1055
R33281 VDD.n10943 VDD.n10942 0.1055
R33282 VDD.n1874 VDD.n1848 0.1055
R33283 VDD.n10948 VDD.n1848 0.1055
R33284 VDD.n10971 VDD.n1833 0.1055
R33285 VDD.n1850 VDD.n1833 0.1055
R33286 VDD.n10998 VDD.n1830 0.1055
R33287 VDD.n10998 VDD.n10997 0.1055
R33288 VDD.n1818 VDD.n1785 0.1055
R33289 VDD.n11003 VDD.n1785 0.1055
R33290 VDD.n11027 VDD.n11026 0.1055
R33291 VDD.n11028 VDD.n11027 0.1055
R33292 VDD.n8758 VDD.n176 0.1055
R33293 VDD.n8536 VDD.n176 0.1055
R33294 VDD.n8805 VDD.n8804 0.1055
R33295 VDD.n8806 VDD.n8805 0.1055
R33296 VDD.n8884 VDD.n8883 0.1055
R33297 VDD.n8883 VDD.n8882 0.1055
R33298 VDD.n8936 VDD.n8935 0.1055
R33299 VDD.n8937 VDD.n8936 0.1055
R33300 VDD.n9015 VDD.n9014 0.1055
R33301 VDD.n9014 VDD.n9013 0.1055
R33302 VDD.n9033 VDD.n9032 0.1055
R33303 VDD.n9034 VDD.n9033 0.1055
R33304 VDD.n9157 VDD.n9156 0.1055
R33305 VDD.n9158 VDD.n9157 0.1055
R33306 VDD.n9144 VDD.n8460 0.1055
R33307 VDD.n9181 VDD.n8460 0.1055
R33308 VDD.n8741 VDD.n123 0.1055
R33309 VDD.n12463 VDD.n123 0.1055
R33310 VDD.n8720 VDD.n111 0.1055
R33311 VDD.n12470 VDD.n111 0.1055
R33312 VDD.n8708 VDD.n96 0.1055
R33313 VDD.n114 VDD.n96 0.1055
R33314 VDD.n8682 VDD.n43 0.1055
R33315 VDD.n12519 VDD.n43 0.1055
R33316 VDD.n8670 VDD.n31 0.1055
R33317 VDD.n12526 VDD.n31 0.1055
R33318 VDD.n8649 VDD.n16 0.1055
R33319 VDD.n34 VDD.n16 0.1055
R33320 VDD.n12615 VDD.n12614 0.1055
R33321 VDD.n12614 VDD.n12613 0.1055
R33322 VDD.n7176 VDD.n7175 0.101802
R33323 VDD.n7175 VDD.n2296 0.101802
R33324 VDD.n7828 VDD.n7827 0.101802
R33325 VDD.n7827 VDD.n7826 0.101802
R33326 VDD.n6978 VDD.n6901 0.10175
R33327 VDD.n6921 VDD.n6920 0.10175
R33328 VDD.n6535 VDD.n6434 0.10175
R33329 VDD.n6495 VDD.n6471 0.10175
R33330 VDD.n6313 VDD.n6312 0.0931471
R33331 VDD.n6312 VDD.n6311 0.0931471
R33332 VDD.n5943 VDD.n5942 0.0931471
R33333 VDD.n5942 VDD.n5376 0.0931471
R33334 VDD.n5943 VDD.n5275 0.0931471
R33335 VDD.n6370 VDD.n5275 0.0931471
R33336 VDD.n7135 VDD.n2312 0.0931471
R33337 VDD.n2317 VDD.n2312 0.0931471
R33338 VDD.n7135 VDD.n7134 0.0931471
R33339 VDD.n7134 VDD.n7133 0.0931471
R33340 VDD.n7836 VDD.n7835 0.0931471
R33341 VDD.n7835 VDD.n7834 0.0931471
R33342 VDD.n6310 VDD.n6309 0.0931471
R33343 VDD.n6311 VDD.n6310 0.0931471
R33344 VDD.n6368 VDD.n5378 0.0931471
R33345 VDD.n5378 VDD.n5376 0.0931471
R33346 VDD.n6369 VDD.n6368 0.0931471
R33347 VDD.n6370 VDD.n6369 0.0931471
R33348 VDD.n2367 VDD.n2366 0.0931471
R33349 VDD.n2367 VDD.n2317 0.0931471
R33350 VDD.n2366 VDD.n2319 0.0931471
R33351 VDD.n7133 VDD.n2319 0.0931471
R33352 VDD.n6195 VDD.n5311 0.0931471
R33353 VDD.n6311 VDD.n5311 0.0931471
R33354 VDD.n6372 VDD.n5312 0.0931471
R33355 VDD.n5376 VDD.n5312 0.0931471
R33356 VDD.n6372 VDD.n6371 0.0931471
R33357 VDD.n6371 VDD.n6370 0.0931471
R33358 VDD.n6185 VDD.n5303 0.0931471
R33359 VDD.n6311 VDD.n5303 0.0931471
R33360 VDD.n5368 VDD.n5304 0.0931471
R33361 VDD.n5376 VDD.n5304 0.0931471
R33362 VDD.n5368 VDD.n5282 0.0931471
R33363 VDD.n6370 VDD.n5282 0.0931471
R33364 VDD.n7833 VDD.n7832 0.0931471
R33365 VDD.n7834 VDD.n7833 0.0931471
R33366 VDD.n6631 VDD.n5270 0.0931471
R33367 VDD.n5270 VDD.n5268 0.0931471
R33368 VDD.n6632 VDD.n6631 0.0931471
R33369 VDD.n6633 VDD.n6632 0.0931471
R33370 VDD.n6635 VDD.n5266 0.0931471
R33371 VDD.n5268 VDD.n5266 0.0931471
R33372 VDD.n6635 VDD.n6634 0.0931471
R33373 VDD.n6634 VDD.n6633 0.0931471
R33374 VDD.n6692 VDD.n5264 0.0931471
R33375 VDD.n5268 VDD.n5264 0.0931471
R33376 VDD.n6692 VDD.n2349 0.0931471
R33377 VDD.n6633 VDD.n2349 0.0931471
R33378 VDD.n6706 VDD.n5221 0.0931471
R33379 VDD.n5268 VDD.n5221 0.0931471
R33380 VDD.n6706 VDD.n2369 0.0931471
R33381 VDD.n6633 VDD.n2369 0.0931471
R33382 VDD.n7043 VDD.n7042 0.0931471
R33383 VDD.n7042 VDD.n2317 0.0931471
R33384 VDD.n7043 VDD.n2318 0.0931471
R33385 VDD.n7133 VDD.n2318 0.0931471
R33386 VDD.n7131 VDD.n2321 0.0931471
R33387 VDD.n2321 VDD.n2317 0.0931471
R33388 VDD.n7132 VDD.n7131 0.0931471
R33389 VDD.n7133 VDD.n7132 0.0931471
R33390 VDD.n7700 VDD.n2236 0.0931471
R33391 VDD.n7834 VDD.n2236 0.0931471
R33392 VDD.n7821 VDD.n2235 0.0931471
R33393 VDD.n7834 VDD.n2235 0.0931471
R33394 VDD.n6318 VDD.n6317 0.0831095
R33395 VDD.n6181 VDD.n6180 0.0831095
R33396 VDD.n6301 VDD.n6300 0.0799891
R33397 VDD.n6305 VDD.n5487 0.0799891
R33398 VDD.n5984 VDD.n5487 0.0799891
R33399 VDD.n6191 VDD.n6190 0.0799891
R33400 VDD.n6300 VDD.n6199 0.0799891
R33401 VDD.n6190 VDD.n6189 0.0799891
R33402 VDD.n7864 VDD.n2187 0.0737558
R33403 VDD.n2355 VDD.n2187 0.0737558
R33404 VDD.n7889 VDD.n2188 0.0737558
R33405 VDD.n7837 VDD.n7836 0.0723953
R33406 VDD.n7832 VDD.n7831 0.0723953
R33407 VDD.n2130 VDD.n2128 0.0720299
R33408 VDD.n8047 VDD.n2149 0.0692176
R33409 VDD.n7994 VDD.n7993 0.0682419
R33410 VDD.n7995 VDD.n7994 0.0682419
R33411 VDD.n7997 VDD.n7996 0.0682419
R33412 VDD.n7996 VDD.n7995 0.0682419
R33413 VDD.n5481 VDD.n5309 0.0682419
R33414 VDD.n6396 VDD.n5309 0.0682419
R33415 VDD.n5459 VDD.n5279 0.0682419
R33416 VDD.n6577 VDD.n5279 0.0682419
R33417 VDD.n5420 VDD.n2357 0.0682419
R33418 VDD.n7040 VDD.n2357 0.0682419
R33419 VDD.n2305 VDD.n2210 0.0682419
R33420 VDD.n7086 VDD.n2210 0.0682419
R33421 VDD.n6283 VDD.n5310 0.0682419
R33422 VDD.n6396 VDD.n5310 0.0682419
R33423 VDD.n6247 VDD.n5280 0.0682419
R33424 VDD.n6577 VDD.n5280 0.0682419
R33425 VDD.n6395 VDD.n6394 0.0682419
R33426 VDD.n6396 VDD.n6395 0.0682419
R33427 VDD.n5348 VDD.n5281 0.0682419
R33428 VDD.n6577 VDD.n5281 0.0682419
R33429 VDD.n5249 VDD.n2348 0.0682419
R33430 VDD.n7040 VDD.n2348 0.0682419
R33431 VDD.n6398 VDD.n6397 0.0682419
R33432 VDD.n6397 VDD.n6396 0.0682419
R33433 VDD.n6576 VDD.n6575 0.0682419
R33434 VDD.n6577 VDD.n6576 0.0682419
R33435 VDD.n6861 VDD.n2237 0.0682419
R33436 VDD.n7086 VDD.n2237 0.0682419
R33437 VDD.n7039 VDD.n7038 0.0682419
R33438 VDD.n7040 VDD.n7039 0.0682419
R33439 VDD.n2368 VDD.n2350 0.0682419
R33440 VDD.n7040 VDD.n2368 0.0682419
R33441 VDD.n7085 VDD.n7084 0.0682419
R33442 VDD.n7086 VDD.n7085 0.0682419
R33443 VDD.n7110 VDD.n7087 0.0682419
R33444 VDD.n7087 VDD.n7086 0.0682419
R33445 VDD.n1563 VDD.n1511 0.0677787
R33446 VDD.n1561 VDD.n1511 0.0677787
R33447 VDD.n1561 VDD.n1560 0.0677787
R33448 VDD.n1560 VDD.n1559 0.0677787
R33449 VDD.n1538 VDD.n1537 0.0677787
R33450 VDD.n1539 VDD.n1538 0.0677787
R33451 VDD.n1539 VDD.n1536 0.0677787
R33452 VDD.n1541 VDD.n1536 0.0677787
R33453 VDD.n1514 VDD.n771 0.0677787
R33454 VDD.n1515 VDD.n1514 0.0677787
R33455 VDD.n1515 VDD.n1513 0.0677787
R33456 VDD.n1517 VDD.n1513 0.0677787
R33457 VDD.n1525 VDD.n1518 0.0677787
R33458 VDD.n1526 VDD.n1525 0.0677787
R33459 VDD.n1526 VDD.n1524 0.0677787
R33460 VDD.n1528 VDD.n1524 0.0677787
R33461 VDD.n5965 VDD.n5308 0.0668158
R33462 VDD.n6396 VDD.n5308 0.0668158
R33463 VDD.n6579 VDD.n6578 0.0668158
R33464 VDD.n6578 VDD.n6577 0.0668158
R33465 VDD.n6610 VDD.n2353 0.0668158
R33466 VDD.n7040 VDD.n2353 0.0668158
R33467 VDD.n2234 VDD.n2233 0.0668158
R33468 VDD.n7086 VDD.n2234 0.0668158
R33469 VDD.n5481 VDD.n5307 0.0668158
R33470 VDD.n6396 VDD.n5307 0.0668158
R33471 VDD.n5459 VDD.n5278 0.0668158
R33472 VDD.n6577 VDD.n5278 0.0668158
R33473 VDD.n5420 VDD.n2352 0.0668158
R33474 VDD.n7040 VDD.n2352 0.0668158
R33475 VDD.n2332 VDD.n2305 0.0668158
R33476 VDD.n7086 VDD.n2332 0.0668158
R33477 VDD.n6283 VDD.n5306 0.0668158
R33478 VDD.n6396 VDD.n5306 0.0668158
R33479 VDD.n6247 VDD.n5277 0.0668158
R33480 VDD.n6577 VDD.n5277 0.0668158
R33481 VDD.n6394 VDD.n5305 0.0668158
R33482 VDD.n6396 VDD.n5305 0.0668158
R33483 VDD.n5348 VDD.n5276 0.0668158
R33484 VDD.n6577 VDD.n5276 0.0668158
R33485 VDD.n5249 VDD.n2351 0.0668158
R33486 VDD.n7040 VDD.n2351 0.0668158
R33487 VDD.n7041 VDD.n2350 0.0668158
R33488 VDD.n7041 VDD.n7040 0.0668158
R33489 VDD.n7084 VDD.n2331 0.0668158
R33490 VDD.n7086 VDD.n2331 0.0668158
R33491 VDD.n7110 VDD.n2238 0.0668158
R33492 VDD.n7086 VDD.n2238 0.0668158
R33493 VDD.n7836 VDD.n2209 0.0629767
R33494 VDD.n7832 VDD.n2239 0.0629767
R33495 VDD.n1553 VDD.n1552 0.0628762
R33496 VDD.n1552 VDD.n1551 0.0628762
R33497 VDD.n752 VDD.n751 0.0627244
R33498 VDD.n1507 VDD.n1506 0.0627244
R33499 VDD.n7947 VDD.n7853 0.0619118
R33500 VDD.n1550 VDD.n1512 0.061665
R33501 VDD.n1551 VDD.n1550 0.061665
R33502 VDD.n7960 VDD.n7959 0.0616241
R33503 VDD.n7823 VDD.n7822 0.0585814
R33504 VDD.n6309 VDD.n6308 0.0569142
R33505 VDD.n6314 VDD.n6313 0.0569142
R33506 VDD.n6196 VDD.n6195 0.0569142
R33507 VDD.n6186 VDD.n6185 0.0569142
R33508 VDD.n847 VDD.n739 0.0543462
R33509 VDD.n1429 VDD.n847 0.0543462
R33510 VDD.n848 VDD.n738 0.0543462
R33511 VDD.n1428 VDD.n848 0.0543462
R33512 VDD.n1347 VDD.n744 0.0543462
R33513 VDD.n1347 VDD.n1346 0.0543462
R33514 VDD.n758 VDD.n744 0.0543462
R33515 VDD.n1345 VDD.n758 0.0543462
R33516 VDD.n1417 VDD.n859 0.0543462
R33517 VDD.n874 VDD.n859 0.0543462
R33518 VDD.n1417 VDD.n1416 0.0543462
R33519 VDD.n1416 VDD.n1415 0.0543462
R33520 VDD.n1431 VDD.n1430 0.0543462
R33521 VDD.n1430 VDD.n1429 0.0543462
R33522 VDD.n1427 VDD.n1426 0.0543462
R33523 VDD.n1428 VDD.n1427 0.0543462
R33524 VDD.n1627 VDD.n764 0.0543462
R33525 VDD.n764 VDD.n763 0.0543462
R33526 VDD.n759 VDD.n747 0.0543462
R33527 VDD.n763 VDD.n759 0.0543462
R33528 VDD.n1277 VDD.n783 0.0543462
R33529 VDD.n1346 VDD.n1277 0.0543462
R33530 VDD.n783 VDD.n762 0.0543462
R33531 VDD.n1345 VDD.n762 0.0543462
R33532 VDD.n1353 VDD.n1352 0.0543462
R33533 VDD.n1354 VDD.n1353 0.0543462
R33534 VDD.n1352 VDD.n1351 0.0543462
R33535 VDD.n1351 VDD.n1084 0.0543462
R33536 VDD.n1083 VDD.n741 0.0543462
R33537 VDD.n1354 VDD.n1083 0.0543462
R33538 VDD.n1344 VDD.n741 0.0543462
R33539 VDD.n1344 VDD.n1084 0.0543462
R33540 VDD.n736 VDD.n712 0.0543462
R33541 VDD.n874 VDD.n712 0.0543462
R33542 VDD.n875 VDD.n736 0.0543462
R33543 VDD.n1415 VDD.n875 0.0543462
R33544 VDD.n1046 VDD.n710 0.0543462
R33545 VDD.n1719 VDD.n710 0.0543462
R33546 VDD.n1046 VDD.n692 0.0543462
R33547 VDD.n709 VDD.n692 0.0543462
R33548 VDD.n1721 VDD.n687 0.0543462
R33549 VDD.n709 VDD.n687 0.0543462
R33550 VDD.n1721 VDD.n1720 0.0543462
R33551 VDD.n1720 VDD.n1719 0.0543462
R33552 VDD.n1032 VDD.n691 0.0543462
R33553 VDD.n691 VDD.n690 0.0543462
R33554 VDD.n985 VDD.n686 0.0543462
R33555 VDD.n690 VDD.n686 0.0543462
R33556 VDD.n5364 VDD.n5363 0.0525345
R33557 VDD.n5373 VDD.n5372 0.0525345
R33558 VDD.n6377 VDD.n6376 0.0525345
R33559 VDD.n6364 VDD.n6363 0.0525345
R33560 VDD.n5938 VDD.n5937 0.0525345
R33561 VDD.n5948 VDD.n5947 0.0525345
R33562 VDD.n2362 VDD.n2361 0.0525345
R33563 VDD.n7140 VDD.n7139 0.0525345
R33564 VDD.n2400 VDD.n2399 0.0525345
R33565 VDD.n7127 VDD.n7126 0.0525345
R33566 VDD.n2344 VDD.n2343 0.0525345
R33567 VDD.n2128 VDD.n2122 0.0513315
R33568 VDD.n7889 VDD.n7888 0.0507941
R33569 VDD.n6266 VDD.n6218 0.050569
R33570 VDD.n6266 VDD.n6265 0.050569
R33571 VDD.n7048 VDD.n2341 0.050569
R33572 VDD.n2313 VDD.n2199 0.050569
R33573 VDD.n7048 VDD.n7047 0.050569
R33574 VDD.n6309 VDD.n6304 0.0495237
R33575 VDD.n6313 VDD.n5987 0.0495237
R33576 VDD.n6195 VDD.n6194 0.0495237
R33577 VDD.n6185 VDD.n6184 0.0495237
R33578 VDD.n8084 VDD.n2121 0.0465048
R33579 VDD.n2141 VDD.n2140 0.0445515
R33580 VDD.n8069 VDD.n8068 0.0440678
R33581 VDD.n8081 VDD.n8080 0.0436757
R33582 VDD.n8085 VDD.n8084 0.0436757
R33583 VDD.n2143 VDD.n2127 0.0433141
R33584 VDD.n2144 VDD.n2127 0.0433141
R33585 VDD.n2145 VDD.n2125 0.0433141
R33586 VDD.n8074 VDD.n2126 0.0433141
R33587 VDD.n8071 VDD.n2126 0.0433141
R33588 VDD.n8071 VDD.n8070 0.0433141
R33589 VDD.n8070 VDD.n8069 0.0433141
R33590 VDD.n2143 VDD.n2142 0.0430669
R33591 VDD.n7890 VDD.n7887 0.0430647
R33592 VDD.n7910 VDD.n7909 0.0428653
R33593 VDD.n7945 VDD.n7944 0.0417941
R33594 VDD.n8050 VDD.n8049 0.0417941
R33595 VDD.n1662 VDD.n1661 0.0416398
R33596 VDD.n1643 VDD.n1642 0.0416398
R33597 VDD.n1592 VDD.n1576 0.0416398
R33598 VDD.n1592 VDD.n1591 0.0416398
R33599 VDD.n7862 VDD.n7861 0.0416007
R33600 VDD.n7947 VDD.n7946 0.0415824
R33601 VDD.n7959 VDD.n2204 0.0413899
R33602 VDD.n2295 VDD.n2294 0.041314
R33603 VDD.n7839 VDD.n7838 0.041314
R33604 VDD.n2387 VDD.n2386 0.041314
R33605 VDD.n7830 VDD.n7829 0.041314
R33606 VDD.n7825 VDD.n7824 0.041314
R33607 VDD.n5216 VDD.n2423 0.0410752
R33608 VDD.n5215 VDD.n2422 0.0410752
R33609 VDD.n5214 VDD.n2421 0.0410752
R33610 VDD.n5213 VDD.n2420 0.0410752
R33611 VDD.n5212 VDD.n2419 0.0410752
R33612 VDD.n5211 VDD.n2418 0.0410752
R33613 VDD.n5210 VDD.n2417 0.0410752
R33614 VDD.n5209 VDD.n2416 0.0410752
R33615 VDD.n5208 VDD.n2415 0.0410752
R33616 VDD.n5207 VDD.n2414 0.0410752
R33617 VDD.n5206 VDD.n2413 0.0410752
R33618 VDD.n5205 VDD.n2412 0.0410752
R33619 VDD.n4597 VDD.n4596 0.0410752
R33620 VDD.n5217 VDD.n2423 0.0410752
R33621 VDD.n5216 VDD.n2422 0.0410752
R33622 VDD.n5215 VDD.n2421 0.0410752
R33623 VDD.n5214 VDD.n2420 0.0410752
R33624 VDD.n5213 VDD.n2419 0.0410752
R33625 VDD.n5212 VDD.n2418 0.0410752
R33626 VDD.n5211 VDD.n2417 0.0410752
R33627 VDD.n5210 VDD.n2416 0.0410752
R33628 VDD.n5209 VDD.n2415 0.0410752
R33629 VDD.n5208 VDD.n2414 0.0410752
R33630 VDD.n5207 VDD.n2413 0.0410752
R33631 VDD.n5206 VDD.n2412 0.0410752
R33632 VDD.n5203 VDD.n4596 0.0410752
R33633 VDD.n12446 VDD.n191 0.0410752
R33634 VDD.n12442 VDD.n192 0.0410752
R33635 VDD.n12443 VDD.n193 0.0410752
R33636 VDD.n9188 VDD.n9187 0.0410752
R33637 VDD.n9190 VDD.n9189 0.0410752
R33638 VDD.n9192 VDD.n9191 0.0410752
R33639 VDD.n9194 VDD.n9193 0.0410752
R33640 VDD.n9196 VDD.n9195 0.0410752
R33641 VDD.n9198 VDD.n9197 0.0410752
R33642 VDD.n9199 VDD.n9198 0.0410752
R33643 VDD.n9189 VDD.n9188 0.0410752
R33644 VDD.n9191 VDD.n9190 0.0410752
R33645 VDD.n9193 VDD.n9192 0.0410752
R33646 VDD.n9195 VDD.n9194 0.0410752
R33647 VDD.n9197 VDD.n9196 0.0410752
R33648 VDD.n12444 VDD.n193 0.0410752
R33649 VDD.n12443 VDD.n192 0.0410752
R33650 VDD.n12442 VDD.n191 0.0410752
R33651 VDD.n2145 VDD.n2144 0.040902
R33652 VDD.n1480 VDD.n1477 0.0404831
R33653 VDD.n1611 VDD.n1610 0.0404831
R33654 VDD.n1610 VDD.n1609 0.0404831
R33655 VDD.n1480 VDD.n1478 0.0404831
R33656 VDD.n5200 VDD.n4598 0.04025
R33657 VDD.n5196 VDD.n4598 0.04025
R33658 VDD.n5196 VDD.n5195 0.04025
R33659 VDD.n5195 VDD.n5194 0.04025
R33660 VDD.n5194 VDD.n4601 0.04025
R33661 VDD.n5190 VDD.n4601 0.04025
R33662 VDD.n5190 VDD.n5189 0.04025
R33663 VDD.n5189 VDD.n5188 0.04025
R33664 VDD.n5188 VDD.n4603 0.04025
R33665 VDD.n5184 VDD.n4603 0.04025
R33666 VDD.n5184 VDD.n5183 0.04025
R33667 VDD.n5183 VDD.n5182 0.04025
R33668 VDD.n5182 VDD.n4605 0.04025
R33669 VDD.n5178 VDD.n4605 0.04025
R33670 VDD.n5178 VDD.n5177 0.04025
R33671 VDD.n5177 VDD.n5176 0.04025
R33672 VDD.n5176 VDD.n4607 0.04025
R33673 VDD.n5172 VDD.n4607 0.04025
R33674 VDD.n5172 VDD.n5171 0.04025
R33675 VDD.n5171 VDD.n5170 0.04025
R33676 VDD.n5170 VDD.n4609 0.04025
R33677 VDD.n5166 VDD.n4609 0.04025
R33678 VDD.n5166 VDD.n5165 0.04025
R33679 VDD.n5165 VDD.n5164 0.04025
R33680 VDD.n5164 VDD.n4611 0.04025
R33681 VDD.n5160 VDD.n4611 0.04025
R33682 VDD.n5160 VDD.n5159 0.04025
R33683 VDD.n5159 VDD.n5158 0.04025
R33684 VDD.n5158 VDD.n4613 0.04025
R33685 VDD.n5154 VDD.n4613 0.04025
R33686 VDD.n5154 VDD.n5153 0.04025
R33687 VDD.n5153 VDD.n5152 0.04025
R33688 VDD.n5152 VDD.n4615 0.04025
R33689 VDD.n5148 VDD.n4615 0.04025
R33690 VDD.n5148 VDD.n5147 0.04025
R33691 VDD.n5147 VDD.n5146 0.04025
R33692 VDD.n5146 VDD.n4617 0.04025
R33693 VDD.n5142 VDD.n4617 0.04025
R33694 VDD.n5142 VDD.n5141 0.04025
R33695 VDD.n5141 VDD.n5140 0.04025
R33696 VDD.n5140 VDD.n4619 0.04025
R33697 VDD.n5136 VDD.n4619 0.04025
R33698 VDD.n5136 VDD.n5135 0.04025
R33699 VDD.n5135 VDD.n5134 0.04025
R33700 VDD.n5134 VDD.n4621 0.04025
R33701 VDD.n5130 VDD.n4621 0.04025
R33702 VDD.n5130 VDD.n5129 0.04025
R33703 VDD.n5129 VDD.n5128 0.04025
R33704 VDD.n5128 VDD.n4623 0.04025
R33705 VDD.n5124 VDD.n4623 0.04025
R33706 VDD.n5124 VDD.n5123 0.04025
R33707 VDD.n5123 VDD.n5122 0.04025
R33708 VDD.n5122 VDD.n4625 0.04025
R33709 VDD.n5118 VDD.n4625 0.04025
R33710 VDD.n5118 VDD.n5117 0.04025
R33711 VDD.n5117 VDD.n5116 0.04025
R33712 VDD.n5116 VDD.n4627 0.04025
R33713 VDD.n5112 VDD.n4627 0.04025
R33714 VDD.n5112 VDD.n5111 0.04025
R33715 VDD.n5111 VDD.n5110 0.04025
R33716 VDD.n5110 VDD.n4629 0.04025
R33717 VDD.n5106 VDD.n4629 0.04025
R33718 VDD.n5106 VDD.n5105 0.04025
R33719 VDD.n5105 VDD.n5104 0.04025
R33720 VDD.n5104 VDD.n4631 0.04025
R33721 VDD.n5100 VDD.n4631 0.04025
R33722 VDD.n5100 VDD.n5099 0.04025
R33723 VDD.n5099 VDD.n5098 0.04025
R33724 VDD.n5098 VDD.n4633 0.04025
R33725 VDD.n5094 VDD.n4633 0.04025
R33726 VDD.n5094 VDD.n5093 0.04025
R33727 VDD.n5093 VDD.n5092 0.04025
R33728 VDD.n5092 VDD.n4635 0.04025
R33729 VDD.n5088 VDD.n4635 0.04025
R33730 VDD.n5088 VDD.n5087 0.04025
R33731 VDD.n5087 VDD.n5086 0.04025
R33732 VDD.n5086 VDD.n4637 0.04025
R33733 VDD.n5082 VDD.n4637 0.04025
R33734 VDD.n5082 VDD.n5081 0.04025
R33735 VDD.n5081 VDD.n5080 0.04025
R33736 VDD.n5080 VDD.n4639 0.04025
R33737 VDD.n5076 VDD.n4639 0.04025
R33738 VDD.n5076 VDD.n5075 0.04025
R33739 VDD.n5075 VDD.n5074 0.04025
R33740 VDD.n5074 VDD.n4641 0.04025
R33741 VDD.n5070 VDD.n4641 0.04025
R33742 VDD.n5070 VDD.n5069 0.04025
R33743 VDD.n5069 VDD.n5068 0.04025
R33744 VDD.n5068 VDD.n4643 0.04025
R33745 VDD.n5064 VDD.n4643 0.04025
R33746 VDD.n5064 VDD.n5063 0.04025
R33747 VDD.n5063 VDD.n5062 0.04025
R33748 VDD.n5062 VDD.n4645 0.04025
R33749 VDD.n5058 VDD.n4645 0.04025
R33750 VDD.n5058 VDD.n5057 0.04025
R33751 VDD.n5057 VDD.n5056 0.04025
R33752 VDD.n5056 VDD.n4647 0.04025
R33753 VDD.n5052 VDD.n4647 0.04025
R33754 VDD.n5052 VDD.n5051 0.04025
R33755 VDD.n5051 VDD.n5050 0.04025
R33756 VDD.n5050 VDD.n4649 0.04025
R33757 VDD.n5046 VDD.n4649 0.04025
R33758 VDD.n5046 VDD.n5045 0.04025
R33759 VDD.n5045 VDD.n5044 0.04025
R33760 VDD.n5044 VDD.n4651 0.04025
R33761 VDD.n5040 VDD.n4651 0.04025
R33762 VDD.n5040 VDD.n5039 0.04025
R33763 VDD.n5039 VDD.n5038 0.04025
R33764 VDD.n5038 VDD.n4653 0.04025
R33765 VDD.n5034 VDD.n4653 0.04025
R33766 VDD.n5034 VDD.n5033 0.04025
R33767 VDD.n5033 VDD.n5032 0.04025
R33768 VDD.n5032 VDD.n4655 0.04025
R33769 VDD.n5028 VDD.n4655 0.04025
R33770 VDD.n5028 VDD.n5027 0.04025
R33771 VDD.n5027 VDD.n5026 0.04025
R33772 VDD.n5026 VDD.n4657 0.04025
R33773 VDD.n5022 VDD.n4657 0.04025
R33774 VDD.n5022 VDD.n5021 0.04025
R33775 VDD.n5021 VDD.n5020 0.04025
R33776 VDD.n5020 VDD.n4659 0.04025
R33777 VDD.n5016 VDD.n4659 0.04025
R33778 VDD.n5016 VDD.n5015 0.04025
R33779 VDD.n5015 VDD.n5014 0.04025
R33780 VDD.n5014 VDD.n4661 0.04025
R33781 VDD.n5010 VDD.n4661 0.04025
R33782 VDD.n5010 VDD.n5009 0.04025
R33783 VDD.n5009 VDD.n5008 0.04025
R33784 VDD.n5008 VDD.n4663 0.04025
R33785 VDD.n5004 VDD.n4663 0.04025
R33786 VDD.n5004 VDD.n5003 0.04025
R33787 VDD.n5003 VDD.n5002 0.04025
R33788 VDD.n5002 VDD.n4665 0.04025
R33789 VDD.n4998 VDD.n4665 0.04025
R33790 VDD.n4998 VDD.n4997 0.04025
R33791 VDD.n4997 VDD.n4996 0.04025
R33792 VDD.n4996 VDD.n4667 0.04025
R33793 VDD.n4992 VDD.n4667 0.04025
R33794 VDD.n4992 VDD.n4991 0.04025
R33795 VDD.n4991 VDD.n4990 0.04025
R33796 VDD.n4990 VDD.n4669 0.04025
R33797 VDD.n4986 VDD.n4669 0.04025
R33798 VDD.n4986 VDD.n4985 0.04025
R33799 VDD.n4985 VDD.n4984 0.04025
R33800 VDD.n4984 VDD.n4671 0.04025
R33801 VDD.n4980 VDD.n4671 0.04025
R33802 VDD.n4980 VDD.n4979 0.04025
R33803 VDD.n4979 VDD.n4978 0.04025
R33804 VDD.n4978 VDD.n4673 0.04025
R33805 VDD.n4974 VDD.n4673 0.04025
R33806 VDD.n4974 VDD.n4973 0.04025
R33807 VDD.n4973 VDD.n4972 0.04025
R33808 VDD.n4972 VDD.n4675 0.04025
R33809 VDD.n4968 VDD.n4675 0.04025
R33810 VDD.n4968 VDD.n4967 0.04025
R33811 VDD.n4967 VDD.n4966 0.04025
R33812 VDD.n4966 VDD.n4677 0.04025
R33813 VDD.n4962 VDD.n4677 0.04025
R33814 VDD.n4962 VDD.n4961 0.04025
R33815 VDD.n4961 VDD.n4960 0.04025
R33816 VDD.n4960 VDD.n4679 0.04025
R33817 VDD.n4956 VDD.n4679 0.04025
R33818 VDD.n4956 VDD.n4955 0.04025
R33819 VDD.n4955 VDD.n4954 0.04025
R33820 VDD.n4954 VDD.n4681 0.04025
R33821 VDD.n4950 VDD.n4681 0.04025
R33822 VDD.n4950 VDD.n4949 0.04025
R33823 VDD.n4949 VDD.n4948 0.04025
R33824 VDD.n4948 VDD.n4683 0.04025
R33825 VDD.n4944 VDD.n4683 0.04025
R33826 VDD.n4944 VDD.n4943 0.04025
R33827 VDD.n4943 VDD.n4942 0.04025
R33828 VDD.n4942 VDD.n4685 0.04025
R33829 VDD.n4938 VDD.n4685 0.04025
R33830 VDD.n4938 VDD.n4937 0.04025
R33831 VDD.n4937 VDD.n4936 0.04025
R33832 VDD.n4936 VDD.n4687 0.04025
R33833 VDD.n4932 VDD.n4687 0.04025
R33834 VDD.n4932 VDD.n4931 0.04025
R33835 VDD.n4931 VDD.n4930 0.04025
R33836 VDD.n4930 VDD.n4689 0.04025
R33837 VDD.n4926 VDD.n4689 0.04025
R33838 VDD.n4926 VDD.n4925 0.04025
R33839 VDD.n4925 VDD.n4924 0.04025
R33840 VDD.n4924 VDD.n4691 0.04025
R33841 VDD.n4920 VDD.n4691 0.04025
R33842 VDD.n4920 VDD.n4919 0.04025
R33843 VDD.n4919 VDD.n4918 0.04025
R33844 VDD.n4918 VDD.n4693 0.04025
R33845 VDD.n4914 VDD.n4693 0.04025
R33846 VDD.n4914 VDD.n4913 0.04025
R33847 VDD.n4913 VDD.n4912 0.04025
R33848 VDD.n4912 VDD.n4695 0.04025
R33849 VDD.n4908 VDD.n4695 0.04025
R33850 VDD.n4908 VDD.n4907 0.04025
R33851 VDD.n4907 VDD.n4906 0.04025
R33852 VDD.n4902 VDD.n4697 0.04025
R33853 VDD.n4902 VDD.n4901 0.04025
R33854 VDD.n4901 VDD.n4900 0.04025
R33855 VDD.n4900 VDD.n4699 0.04025
R33856 VDD.n4896 VDD.n4699 0.04025
R33857 VDD.n4896 VDD.n4895 0.04025
R33858 VDD.n4895 VDD.n4894 0.04025
R33859 VDD.n4894 VDD.n4701 0.04025
R33860 VDD.n4890 VDD.n4701 0.04025
R33861 VDD.n4890 VDD.n4889 0.04025
R33862 VDD.n4889 VDD.n4888 0.04025
R33863 VDD.n4888 VDD.n4703 0.04025
R33864 VDD.n4884 VDD.n4703 0.04025
R33865 VDD.n4884 VDD.n4883 0.04025
R33866 VDD.n4883 VDD.n4882 0.04025
R33867 VDD.n4882 VDD.n4705 0.04025
R33868 VDD.n4878 VDD.n4705 0.04025
R33869 VDD.n4878 VDD.n4877 0.04025
R33870 VDD.n4877 VDD.n4876 0.04025
R33871 VDD.n4876 VDD.n4707 0.04025
R33872 VDD.n4872 VDD.n4707 0.04025
R33873 VDD.n4872 VDD.n4871 0.04025
R33874 VDD.n4871 VDD.n4870 0.04025
R33875 VDD.n4870 VDD.n4709 0.04025
R33876 VDD.n4866 VDD.n4709 0.04025
R33877 VDD.n4866 VDD.n4865 0.04025
R33878 VDD.n4865 VDD.n4864 0.04025
R33879 VDD.n4864 VDD.n4711 0.04025
R33880 VDD.n4860 VDD.n4711 0.04025
R33881 VDD.n4860 VDD.n4859 0.04025
R33882 VDD.n4859 VDD.n4858 0.04025
R33883 VDD.n4858 VDD.n4713 0.04025
R33884 VDD.n4854 VDD.n4713 0.04025
R33885 VDD.n4854 VDD.n4853 0.04025
R33886 VDD.n4853 VDD.n4852 0.04025
R33887 VDD.n4852 VDD.n4715 0.04025
R33888 VDD.n4848 VDD.n4715 0.04025
R33889 VDD.n4848 VDD.n4847 0.04025
R33890 VDD.n4847 VDD.n4846 0.04025
R33891 VDD.n4846 VDD.n4717 0.04025
R33892 VDD.n4842 VDD.n4717 0.04025
R33893 VDD.n4842 VDD.n4841 0.04025
R33894 VDD.n4841 VDD.n4840 0.04025
R33895 VDD.n4840 VDD.n4719 0.04025
R33896 VDD.n4836 VDD.n4719 0.04025
R33897 VDD.n4836 VDD.n4835 0.04025
R33898 VDD.n4835 VDD.n4834 0.04025
R33899 VDD.n4834 VDD.n4721 0.04025
R33900 VDD.n4830 VDD.n4721 0.04025
R33901 VDD.n4830 VDD.n4829 0.04025
R33902 VDD.n4829 VDD.n4828 0.04025
R33903 VDD.n4828 VDD.n4723 0.04025
R33904 VDD.n4824 VDD.n4723 0.04025
R33905 VDD.n4824 VDD.n4823 0.04025
R33906 VDD.n4823 VDD.n4822 0.04025
R33907 VDD.n4822 VDD.n4725 0.04025
R33908 VDD.n4818 VDD.n4725 0.04025
R33909 VDD.n4818 VDD.n4817 0.04025
R33910 VDD.n4817 VDD.n4816 0.04025
R33911 VDD.n4816 VDD.n4727 0.04025
R33912 VDD.n4812 VDD.n4727 0.04025
R33913 VDD.n4812 VDD.n4811 0.04025
R33914 VDD.n4811 VDD.n4810 0.04025
R33915 VDD.n4810 VDD.n4729 0.04025
R33916 VDD.n4806 VDD.n4729 0.04025
R33917 VDD.n4806 VDD.n4805 0.04025
R33918 VDD.n4805 VDD.n4804 0.04025
R33919 VDD.n4804 VDD.n4731 0.04025
R33920 VDD.n4800 VDD.n4731 0.04025
R33921 VDD.n4800 VDD.n4799 0.04025
R33922 VDD.n4799 VDD.n4798 0.04025
R33923 VDD.n4798 VDD.n4733 0.04025
R33924 VDD.n4794 VDD.n4733 0.04025
R33925 VDD.n4794 VDD.n4793 0.04025
R33926 VDD.n4793 VDD.n4792 0.04025
R33927 VDD.n4792 VDD.n4735 0.04025
R33928 VDD.n4788 VDD.n4735 0.04025
R33929 VDD.n4788 VDD.n4787 0.04025
R33930 VDD.n4787 VDD.n4786 0.04025
R33931 VDD.n4786 VDD.n4737 0.04025
R33932 VDD.n4782 VDD.n4737 0.04025
R33933 VDD.n4782 VDD.n4781 0.04025
R33934 VDD.n4781 VDD.n4780 0.04025
R33935 VDD.n4780 VDD.n4739 0.04025
R33936 VDD.n4776 VDD.n4739 0.04025
R33937 VDD.n4776 VDD.n4775 0.04025
R33938 VDD.n4775 VDD.n4774 0.04025
R33939 VDD.n4774 VDD.n4741 0.04025
R33940 VDD.n4770 VDD.n4741 0.04025
R33941 VDD.n4770 VDD.n4769 0.04025
R33942 VDD.n4769 VDD.n4768 0.04025
R33943 VDD.n4768 VDD.n4743 0.04025
R33944 VDD.n4764 VDD.n4743 0.04025
R33945 VDD.n4764 VDD.n4763 0.04025
R33946 VDD.n4763 VDD.n4762 0.04025
R33947 VDD.n4762 VDD.n4745 0.04025
R33948 VDD.n4758 VDD.n4745 0.04025
R33949 VDD.n4758 VDD.n4757 0.04025
R33950 VDD.n4757 VDD.n4756 0.04025
R33951 VDD.n4756 VDD.n4747 0.04025
R33952 VDD.n4752 VDD.n4747 0.04025
R33953 VDD.n4752 VDD.n4751 0.04025
R33954 VDD.n4751 VDD.n4750 0.04025
R33955 VDD.n4750 VDD.n2242 0.04025
R33956 VDD.n7682 VDD.n7681 0.04025
R33957 VDD.n7681 VDD.n7178 0.04025
R33958 VDD.n7677 VDD.n7178 0.04025
R33959 VDD.n7677 VDD.n7676 0.04025
R33960 VDD.n7676 VDD.n7675 0.04025
R33961 VDD.n7675 VDD.n7180 0.04025
R33962 VDD.n7671 VDD.n7180 0.04025
R33963 VDD.n7671 VDD.n7670 0.04025
R33964 VDD.n7670 VDD.n7669 0.04025
R33965 VDD.n7669 VDD.n7182 0.04025
R33966 VDD.n7665 VDD.n7182 0.04025
R33967 VDD.n7665 VDD.n7664 0.04025
R33968 VDD.n7664 VDD.n7663 0.04025
R33969 VDD.n7663 VDD.n7184 0.04025
R33970 VDD.n7659 VDD.n7184 0.04025
R33971 VDD.n7659 VDD.n7658 0.04025
R33972 VDD.n7658 VDD.n7657 0.04025
R33973 VDD.n7657 VDD.n7186 0.04025
R33974 VDD.n7653 VDD.n7186 0.04025
R33975 VDD.n7653 VDD.n7652 0.04025
R33976 VDD.n7652 VDD.n7651 0.04025
R33977 VDD.n7651 VDD.n7188 0.04025
R33978 VDD.n7647 VDD.n7188 0.04025
R33979 VDD.n7647 VDD.n7646 0.04025
R33980 VDD.n7646 VDD.n7645 0.04025
R33981 VDD.n7645 VDD.n7190 0.04025
R33982 VDD.n7641 VDD.n7190 0.04025
R33983 VDD.n7641 VDD.n7640 0.04025
R33984 VDD.n7640 VDD.n7639 0.04025
R33985 VDD.n7639 VDD.n7192 0.04025
R33986 VDD.n7635 VDD.n7192 0.04025
R33987 VDD.n7635 VDD.n7634 0.04025
R33988 VDD.n7634 VDD.n7633 0.04025
R33989 VDD.n7633 VDD.n7194 0.04025
R33990 VDD.n7629 VDD.n7194 0.04025
R33991 VDD.n7629 VDD.n7628 0.04025
R33992 VDD.n7628 VDD.n7627 0.04025
R33993 VDD.n7627 VDD.n7196 0.04025
R33994 VDD.n7623 VDD.n7196 0.04025
R33995 VDD.n7623 VDD.n7622 0.04025
R33996 VDD.n7622 VDD.n7621 0.04025
R33997 VDD.n7621 VDD.n7198 0.04025
R33998 VDD.n7617 VDD.n7198 0.04025
R33999 VDD.n7617 VDD.n7616 0.04025
R34000 VDD.n7616 VDD.n7615 0.04025
R34001 VDD.n7615 VDD.n7200 0.04025
R34002 VDD.n7611 VDD.n7200 0.04025
R34003 VDD.n7611 VDD.n7610 0.04025
R34004 VDD.n7610 VDD.n7609 0.04025
R34005 VDD.n7609 VDD.n7202 0.04025
R34006 VDD.n7605 VDD.n7202 0.04025
R34007 VDD.n7605 VDD.n7604 0.04025
R34008 VDD.n7604 VDD.n7603 0.04025
R34009 VDD.n7603 VDD.n7204 0.04025
R34010 VDD.n7599 VDD.n7204 0.04025
R34011 VDD.n7599 VDD.n7598 0.04025
R34012 VDD.n7598 VDD.n7597 0.04025
R34013 VDD.n7597 VDD.n7206 0.04025
R34014 VDD.n7593 VDD.n7206 0.04025
R34015 VDD.n7593 VDD.n7592 0.04025
R34016 VDD.n7592 VDD.n7591 0.04025
R34017 VDD.n7591 VDD.n7208 0.04025
R34018 VDD.n7587 VDD.n7208 0.04025
R34019 VDD.n7587 VDD.n7586 0.04025
R34020 VDD.n7586 VDD.n7585 0.04025
R34021 VDD.n7585 VDD.n7210 0.04025
R34022 VDD.n7581 VDD.n7210 0.04025
R34023 VDD.n7581 VDD.n7580 0.04025
R34024 VDD.n7580 VDD.n7579 0.04025
R34025 VDD.n7579 VDD.n7212 0.04025
R34026 VDD.n7575 VDD.n7212 0.04025
R34027 VDD.n7575 VDD.n7574 0.04025
R34028 VDD.n7574 VDD.n7573 0.04025
R34029 VDD.n7573 VDD.n7214 0.04025
R34030 VDD.n7569 VDD.n7214 0.04025
R34031 VDD.n7569 VDD.n7568 0.04025
R34032 VDD.n7568 VDD.n7567 0.04025
R34033 VDD.n7567 VDD.n7216 0.04025
R34034 VDD.n7563 VDD.n7216 0.04025
R34035 VDD.n7563 VDD.n7562 0.04025
R34036 VDD.n7562 VDD.n7561 0.04025
R34037 VDD.n7561 VDD.n7218 0.04025
R34038 VDD.n7557 VDD.n7218 0.04025
R34039 VDD.n7557 VDD.n7556 0.04025
R34040 VDD.n7556 VDD.n7555 0.04025
R34041 VDD.n7555 VDD.n7220 0.04025
R34042 VDD.n7551 VDD.n7220 0.04025
R34043 VDD.n7551 VDD.n7550 0.04025
R34044 VDD.n7550 VDD.n7549 0.04025
R34045 VDD.n7549 VDD.n7222 0.04025
R34046 VDD.n7545 VDD.n7222 0.04025
R34047 VDD.n7545 VDD.n7544 0.04025
R34048 VDD.n7544 VDD.n7543 0.04025
R34049 VDD.n7543 VDD.n7224 0.04025
R34050 VDD.n7539 VDD.n7224 0.04025
R34051 VDD.n7539 VDD.n7538 0.04025
R34052 VDD.n7538 VDD.n7537 0.04025
R34053 VDD.n7537 VDD.n7226 0.04025
R34054 VDD.n7533 VDD.n7226 0.04025
R34055 VDD.n7533 VDD.n7532 0.04025
R34056 VDD.n7532 VDD.n7531 0.04025
R34057 VDD.n7531 VDD.n7228 0.04025
R34058 VDD.n7527 VDD.n7228 0.04025
R34059 VDD.n7527 VDD.n7526 0.04025
R34060 VDD.n7526 VDD.n7525 0.04025
R34061 VDD.n7525 VDD.n7230 0.04025
R34062 VDD.n7521 VDD.n7230 0.04025
R34063 VDD.n7521 VDD.n7520 0.04025
R34064 VDD.n7520 VDD.n7519 0.04025
R34065 VDD.n7519 VDD.n7232 0.04025
R34066 VDD.n7515 VDD.n7232 0.04025
R34067 VDD.n7515 VDD.n7514 0.04025
R34068 VDD.n7514 VDD.n7513 0.04025
R34069 VDD.n7513 VDD.n7234 0.04025
R34070 VDD.n7509 VDD.n7234 0.04025
R34071 VDD.n7509 VDD.n7508 0.04025
R34072 VDD.n7508 VDD.n7507 0.04025
R34073 VDD.n7507 VDD.n7236 0.04025
R34074 VDD.n7503 VDD.n7236 0.04025
R34075 VDD.n7503 VDD.n7502 0.04025
R34076 VDD.n7502 VDD.n7501 0.04025
R34077 VDD.n7501 VDD.n7238 0.04025
R34078 VDD.n7497 VDD.n7238 0.04025
R34079 VDD.n7497 VDD.n7496 0.04025
R34080 VDD.n7496 VDD.n7495 0.04025
R34081 VDD.n7495 VDD.n7240 0.04025
R34082 VDD.n7491 VDD.n7240 0.04025
R34083 VDD.n7491 VDD.n7490 0.04025
R34084 VDD.n7490 VDD.n7489 0.04025
R34085 VDD.n7489 VDD.n7242 0.04025
R34086 VDD.n7485 VDD.n7242 0.04025
R34087 VDD.n7485 VDD.n7484 0.04025
R34088 VDD.n7484 VDD.n7483 0.04025
R34089 VDD.n7483 VDD.n7244 0.04025
R34090 VDD.n7479 VDD.n7244 0.04025
R34091 VDD.n7479 VDD.n7478 0.04025
R34092 VDD.n7478 VDD.n7477 0.04025
R34093 VDD.n7477 VDD.n7246 0.04025
R34094 VDD.n7473 VDD.n7246 0.04025
R34095 VDD.n7473 VDD.n7472 0.04025
R34096 VDD.n7472 VDD.n7471 0.04025
R34097 VDD.n7471 VDD.n7248 0.04025
R34098 VDD.n7467 VDD.n7248 0.04025
R34099 VDD.n7467 VDD.n7466 0.04025
R34100 VDD.n7466 VDD.n7465 0.04025
R34101 VDD.n7465 VDD.n7250 0.04025
R34102 VDD.n7461 VDD.n7250 0.04025
R34103 VDD.n7461 VDD.n7460 0.04025
R34104 VDD.n7460 VDD.n7459 0.04025
R34105 VDD.n7459 VDD.n7252 0.04025
R34106 VDD.n7455 VDD.n7252 0.04025
R34107 VDD.n7455 VDD.n7454 0.04025
R34108 VDD.n7454 VDD.n7453 0.04025
R34109 VDD.n7453 VDD.n7254 0.04025
R34110 VDD.n7449 VDD.n7254 0.04025
R34111 VDD.n7449 VDD.n7448 0.04025
R34112 VDD.n7448 VDD.n7447 0.04025
R34113 VDD.n7447 VDD.n7256 0.04025
R34114 VDD.n7443 VDD.n7256 0.04025
R34115 VDD.n7443 VDD.n7442 0.04025
R34116 VDD.n7442 VDD.n7441 0.04025
R34117 VDD.n7441 VDD.n7258 0.04025
R34118 VDD.n7437 VDD.n7258 0.04025
R34119 VDD.n7437 VDD.n7436 0.04025
R34120 VDD.n7436 VDD.n7435 0.04025
R34121 VDD.n7435 VDD.n7260 0.04025
R34122 VDD.n7431 VDD.n7260 0.04025
R34123 VDD.n7431 VDD.n7430 0.04025
R34124 VDD.n7430 VDD.n7429 0.04025
R34125 VDD.n7429 VDD.n7262 0.04025
R34126 VDD.n7425 VDD.n7262 0.04025
R34127 VDD.n7425 VDD.n7424 0.04025
R34128 VDD.n7424 VDD.n7423 0.04025
R34129 VDD.n7423 VDD.n7264 0.04025
R34130 VDD.n7419 VDD.n7264 0.04025
R34131 VDD.n7419 VDD.n7418 0.04025
R34132 VDD.n7418 VDD.n7417 0.04025
R34133 VDD.n7417 VDD.n7266 0.04025
R34134 VDD.n7413 VDD.n7266 0.04025
R34135 VDD.n7413 VDD.n7412 0.04025
R34136 VDD.n7412 VDD.n7411 0.04025
R34137 VDD.n7411 VDD.n7268 0.04025
R34138 VDD.n7407 VDD.n7268 0.04025
R34139 VDD.n7407 VDD.n7406 0.04025
R34140 VDD.n7406 VDD.n7405 0.04025
R34141 VDD.n7405 VDD.n7270 0.04025
R34142 VDD.n7401 VDD.n7270 0.04025
R34143 VDD.n7401 VDD.n7400 0.04025
R34144 VDD.n7400 VDD.n7399 0.04025
R34145 VDD.n7399 VDD.n7272 0.04025
R34146 VDD.n7395 VDD.n7272 0.04025
R34147 VDD.n7395 VDD.n7394 0.04025
R34148 VDD.n7394 VDD.n7393 0.04025
R34149 VDD.n7393 VDD.n7274 0.04025
R34150 VDD.n7389 VDD.n7274 0.04025
R34151 VDD.n7389 VDD.n7388 0.04025
R34152 VDD.n7388 VDD.n7387 0.04025
R34153 VDD.n7387 VDD.n7276 0.04025
R34154 VDD.n7383 VDD.n7276 0.04025
R34155 VDD.n7383 VDD.n7382 0.04025
R34156 VDD.n7382 VDD.n7381 0.04025
R34157 VDD.n7381 VDD.n7278 0.04025
R34158 VDD.n7377 VDD.n7278 0.04025
R34159 VDD.n7377 VDD.n7376 0.04025
R34160 VDD.n7376 VDD.n7375 0.04025
R34161 VDD.n7375 VDD.n7280 0.04025
R34162 VDD.n7371 VDD.n7280 0.04025
R34163 VDD.n7371 VDD.n7370 0.04025
R34164 VDD.n7370 VDD.n7369 0.04025
R34165 VDD.n7369 VDD.n7282 0.04025
R34166 VDD.n7365 VDD.n7282 0.04025
R34167 VDD.n7365 VDD.n7364 0.04025
R34168 VDD.n7364 VDD.n7363 0.04025
R34169 VDD.n7363 VDD.n7284 0.04025
R34170 VDD.n7359 VDD.n7284 0.04025
R34171 VDD.n7359 VDD.n7358 0.04025
R34172 VDD.n7358 VDD.n7357 0.04025
R34173 VDD.n7357 VDD.n7286 0.04025
R34174 VDD.n7353 VDD.n7286 0.04025
R34175 VDD.n7353 VDD.n7352 0.04025
R34176 VDD.n7352 VDD.n7351 0.04025
R34177 VDD.n7351 VDD.n7288 0.04025
R34178 VDD.n7347 VDD.n7288 0.04025
R34179 VDD.n7347 VDD.n7346 0.04025
R34180 VDD.n7346 VDD.n7345 0.04025
R34181 VDD.n7345 VDD.n7290 0.04025
R34182 VDD.n7341 VDD.n7290 0.04025
R34183 VDD.n7341 VDD.n7340 0.04025
R34184 VDD.n7340 VDD.n7339 0.04025
R34185 VDD.n7339 VDD.n7292 0.04025
R34186 VDD.n7335 VDD.n7292 0.04025
R34187 VDD.n7335 VDD.n7334 0.04025
R34188 VDD.n7334 VDD.n7333 0.04025
R34189 VDD.n7333 VDD.n7294 0.04025
R34190 VDD.n7329 VDD.n7294 0.04025
R34191 VDD.n7329 VDD.n7328 0.04025
R34192 VDD.n7328 VDD.n7327 0.04025
R34193 VDD.n7327 VDD.n7296 0.04025
R34194 VDD.n7323 VDD.n7296 0.04025
R34195 VDD.n7323 VDD.n7322 0.04025
R34196 VDD.n7322 VDD.n7321 0.04025
R34197 VDD.n7321 VDD.n7298 0.04025
R34198 VDD.n7317 VDD.n7298 0.04025
R34199 VDD.n7317 VDD.n7316 0.04025
R34200 VDD.n7316 VDD.n7315 0.04025
R34201 VDD.n7315 VDD.n7300 0.04025
R34202 VDD.n7311 VDD.n7300 0.04025
R34203 VDD.n7311 VDD.n7310 0.04025
R34204 VDD.n7310 VDD.n7309 0.04025
R34205 VDD.n10759 VDD.n8255 0.04025
R34206 VDD.n10755 VDD.n8255 0.04025
R34207 VDD.n10755 VDD.n10754 0.04025
R34208 VDD.n10754 VDD.n10753 0.04025
R34209 VDD.n10753 VDD.n8257 0.04025
R34210 VDD.n10749 VDD.n8257 0.04025
R34211 VDD.n10749 VDD.n10748 0.04025
R34212 VDD.n10748 VDD.n10747 0.04025
R34213 VDD.n10747 VDD.n8259 0.04025
R34214 VDD.n10743 VDD.n8259 0.04025
R34215 VDD.n10743 VDD.n10742 0.04025
R34216 VDD.n10742 VDD.n10741 0.04025
R34217 VDD.n10741 VDD.n8261 0.04025
R34218 VDD.n10737 VDD.n8261 0.04025
R34219 VDD.n10737 VDD.n10736 0.04025
R34220 VDD.n10736 VDD.n10735 0.04025
R34221 VDD.n10735 VDD.n8263 0.04025
R34222 VDD.n10731 VDD.n8263 0.04025
R34223 VDD.n10731 VDD.n10730 0.04025
R34224 VDD.n10730 VDD.n10729 0.04025
R34225 VDD.n10729 VDD.n8265 0.04025
R34226 VDD.n10725 VDD.n8265 0.04025
R34227 VDD.n10725 VDD.n10724 0.04025
R34228 VDD.n10724 VDD.n10723 0.04025
R34229 VDD.n10723 VDD.n8267 0.04025
R34230 VDD.n10719 VDD.n8267 0.04025
R34231 VDD.n10719 VDD.n10718 0.04025
R34232 VDD.n10718 VDD.n10717 0.04025
R34233 VDD.n10717 VDD.n8269 0.04025
R34234 VDD.n10713 VDD.n8269 0.04025
R34235 VDD.n10713 VDD.n10712 0.04025
R34236 VDD.n10712 VDD.n10711 0.04025
R34237 VDD.n10711 VDD.n8271 0.04025
R34238 VDD.n10707 VDD.n8271 0.04025
R34239 VDD.n10707 VDD.n10706 0.04025
R34240 VDD.n10706 VDD.n10705 0.04025
R34241 VDD.n10705 VDD.n8273 0.04025
R34242 VDD.n10701 VDD.n8273 0.04025
R34243 VDD.n10701 VDD.n10700 0.04025
R34244 VDD.n10700 VDD.n10699 0.04025
R34245 VDD.n10699 VDD.n8275 0.04025
R34246 VDD.n10695 VDD.n8275 0.04025
R34247 VDD.n10695 VDD.n10694 0.04025
R34248 VDD.n10694 VDD.n10693 0.04025
R34249 VDD.n10693 VDD.n8277 0.04025
R34250 VDD.n10689 VDD.n8277 0.04025
R34251 VDD.n10689 VDD.n10688 0.04025
R34252 VDD.n10688 VDD.n10687 0.04025
R34253 VDD.n10687 VDD.n8279 0.04025
R34254 VDD.n10683 VDD.n8279 0.04025
R34255 VDD.n10683 VDD.n10682 0.04025
R34256 VDD.n10682 VDD.n10681 0.04025
R34257 VDD.n10681 VDD.n8281 0.04025
R34258 VDD.n10677 VDD.n8281 0.04025
R34259 VDD.n10677 VDD.n10676 0.04025
R34260 VDD.n10676 VDD.n10675 0.04025
R34261 VDD.n10675 VDD.n8283 0.04025
R34262 VDD.n10671 VDD.n8283 0.04025
R34263 VDD.n10671 VDD.n10670 0.04025
R34264 VDD.n10670 VDD.n10669 0.04025
R34265 VDD.n10669 VDD.n8285 0.04025
R34266 VDD.n10665 VDD.n8285 0.04025
R34267 VDD.n10665 VDD.n10664 0.04025
R34268 VDD.n10664 VDD.n10663 0.04025
R34269 VDD.n10663 VDD.n8287 0.04025
R34270 VDD.n10659 VDD.n8287 0.04025
R34271 VDD.n10659 VDD.n10658 0.04025
R34272 VDD.n10658 VDD.n10657 0.04025
R34273 VDD.n10657 VDD.n8289 0.04025
R34274 VDD.n10653 VDD.n8289 0.04025
R34275 VDD.n10653 VDD.n10652 0.04025
R34276 VDD.n10652 VDD.n10651 0.04025
R34277 VDD.n10651 VDD.n8291 0.04025
R34278 VDD.n10647 VDD.n8291 0.04025
R34279 VDD.n10647 VDD.n10646 0.04025
R34280 VDD.n10646 VDD.n10645 0.04025
R34281 VDD.n10645 VDD.n8293 0.04025
R34282 VDD.n10641 VDD.n8293 0.04025
R34283 VDD.n10641 VDD.n10640 0.04025
R34284 VDD.n10640 VDD.n10639 0.04025
R34285 VDD.n10639 VDD.n8295 0.04025
R34286 VDD.n10635 VDD.n8295 0.04025
R34287 VDD.n10635 VDD.n10634 0.04025
R34288 VDD.n10634 VDD.n10633 0.04025
R34289 VDD.n10633 VDD.n8297 0.04025
R34290 VDD.n10629 VDD.n8297 0.04025
R34291 VDD.n10629 VDD.n10628 0.04025
R34292 VDD.n10628 VDD.n10627 0.04025
R34293 VDD.n10627 VDD.n8299 0.04025
R34294 VDD.n10623 VDD.n8299 0.04025
R34295 VDD.n10623 VDD.n10622 0.04025
R34296 VDD.n10622 VDD.n10621 0.04025
R34297 VDD.n10621 VDD.n8301 0.04025
R34298 VDD.n10617 VDD.n8301 0.04025
R34299 VDD.n10617 VDD.n10616 0.04025
R34300 VDD.n10616 VDD.n10615 0.04025
R34301 VDD.n10615 VDD.n8303 0.04025
R34302 VDD.n10611 VDD.n8303 0.04025
R34303 VDD.n10611 VDD.n10610 0.04025
R34304 VDD.n10610 VDD.n10609 0.04025
R34305 VDD.n10609 VDD.n8305 0.04025
R34306 VDD.n10605 VDD.n8305 0.04025
R34307 VDD.n10605 VDD.n10604 0.04025
R34308 VDD.n10604 VDD.n10603 0.04025
R34309 VDD.n10603 VDD.n8307 0.04025
R34310 VDD.n10599 VDD.n8307 0.04025
R34311 VDD.n10599 VDD.n10598 0.04025
R34312 VDD.n10598 VDD.n10597 0.04025
R34313 VDD.n10597 VDD.n8309 0.04025
R34314 VDD.n10593 VDD.n8309 0.04025
R34315 VDD.n10593 VDD.n10592 0.04025
R34316 VDD.n10592 VDD.n10591 0.04025
R34317 VDD.n10591 VDD.n8311 0.04025
R34318 VDD.n10587 VDD.n8311 0.04025
R34319 VDD.n10587 VDD.n10586 0.04025
R34320 VDD.n10586 VDD.n10585 0.04025
R34321 VDD.n10585 VDD.n8313 0.04025
R34322 VDD.n10581 VDD.n8313 0.04025
R34323 VDD.n10581 VDD.n10580 0.04025
R34324 VDD.n10580 VDD.n10579 0.04025
R34325 VDD.n10579 VDD.n8315 0.04025
R34326 VDD.n10575 VDD.n8315 0.04025
R34327 VDD.n10575 VDD.n10574 0.04025
R34328 VDD.n10574 VDD.n10573 0.04025
R34329 VDD.n10573 VDD.n8317 0.04025
R34330 VDD.n10569 VDD.n8317 0.04025
R34331 VDD.n10569 VDD.n10568 0.04025
R34332 VDD.n10568 VDD.n10567 0.04025
R34333 VDD.n10567 VDD.n8319 0.04025
R34334 VDD.n10563 VDD.n8319 0.04025
R34335 VDD.n10563 VDD.n10562 0.04025
R34336 VDD.n10562 VDD.n10561 0.04025
R34337 VDD.n10561 VDD.n8321 0.04025
R34338 VDD.n10557 VDD.n8321 0.04025
R34339 VDD.n10557 VDD.n10556 0.04025
R34340 VDD.n10556 VDD.n10555 0.04025
R34341 VDD.n10555 VDD.n8323 0.04025
R34342 VDD.n10551 VDD.n8323 0.04025
R34343 VDD.n10551 VDD.n10550 0.04025
R34344 VDD.n10550 VDD.n10549 0.04025
R34345 VDD.n10549 VDD.n8325 0.04025
R34346 VDD.n10545 VDD.n8325 0.04025
R34347 VDD.n10545 VDD.n10544 0.04025
R34348 VDD.n10544 VDD.n10543 0.04025
R34349 VDD.n10543 VDD.n8327 0.04025
R34350 VDD.n10539 VDD.n8327 0.04025
R34351 VDD.n10539 VDD.n10538 0.04025
R34352 VDD.n10538 VDD.n10537 0.04025
R34353 VDD.n10537 VDD.n8329 0.04025
R34354 VDD.n10533 VDD.n8329 0.04025
R34355 VDD.n10533 VDD.n10532 0.04025
R34356 VDD.n10532 VDD.n10531 0.04025
R34357 VDD.n10531 VDD.n8331 0.04025
R34358 VDD.n10527 VDD.n8331 0.04025
R34359 VDD.n10527 VDD.n10526 0.04025
R34360 VDD.n10526 VDD.n10525 0.04025
R34361 VDD.n10525 VDD.n8333 0.04025
R34362 VDD.n10521 VDD.n8333 0.04025
R34363 VDD.n10521 VDD.n10520 0.04025
R34364 VDD.n10520 VDD.n10519 0.04025
R34365 VDD.n10519 VDD.n8335 0.04025
R34366 VDD.n10515 VDD.n8335 0.04025
R34367 VDD.n10515 VDD.n10514 0.04025
R34368 VDD.n10514 VDD.n10513 0.04025
R34369 VDD.n10513 VDD.n8337 0.04025
R34370 VDD.n10509 VDD.n8337 0.04025
R34371 VDD.n10509 VDD.n10508 0.04025
R34372 VDD.n10508 VDD.n10507 0.04025
R34373 VDD.n10507 VDD.n8339 0.04025
R34374 VDD.n10503 VDD.n8339 0.04025
R34375 VDD.n10503 VDD.n10502 0.04025
R34376 VDD.n10502 VDD.n10501 0.04025
R34377 VDD.n10501 VDD.n8341 0.04025
R34378 VDD.n10497 VDD.n8341 0.04025
R34379 VDD.n10497 VDD.n10496 0.04025
R34380 VDD.n10496 VDD.n10495 0.04025
R34381 VDD.n10495 VDD.n8343 0.04025
R34382 VDD.n10491 VDD.n8343 0.04025
R34383 VDD.n10491 VDD.n10490 0.04025
R34384 VDD.n10490 VDD.n10489 0.04025
R34385 VDD.n10489 VDD.n8345 0.04025
R34386 VDD.n10485 VDD.n8345 0.04025
R34387 VDD.n10485 VDD.n10484 0.04025
R34388 VDD.n10484 VDD.n10483 0.04025
R34389 VDD.n10483 VDD.n8347 0.04025
R34390 VDD.n10479 VDD.n8347 0.04025
R34391 VDD.n10479 VDD.n10478 0.04025
R34392 VDD.n10478 VDD.n10477 0.04025
R34393 VDD.n10477 VDD.n8349 0.04025
R34394 VDD.n10473 VDD.n8349 0.04025
R34395 VDD.n10473 VDD.n10472 0.04025
R34396 VDD.n10472 VDD.n10471 0.04025
R34397 VDD.n10471 VDD.n8351 0.04025
R34398 VDD.n10467 VDD.n8351 0.04025
R34399 VDD.n10467 VDD.n10466 0.04025
R34400 VDD.n10466 VDD.n10465 0.04025
R34401 VDD.n10465 VDD.n8353 0.04025
R34402 VDD.n10461 VDD.n8353 0.04025
R34403 VDD.n10461 VDD.n10460 0.04025
R34404 VDD.n10460 VDD.n10459 0.04025
R34405 VDD.n10459 VDD.n8355 0.04025
R34406 VDD.n10455 VDD.n8355 0.04025
R34407 VDD.n10455 VDD.n10454 0.04025
R34408 VDD.n10454 VDD.n10453 0.04025
R34409 VDD.n10453 VDD.n8357 0.04025
R34410 VDD.n10449 VDD.n8357 0.04025
R34411 VDD.n10449 VDD.n10448 0.04025
R34412 VDD.n10448 VDD.n10447 0.04025
R34413 VDD.n10447 VDD.n8359 0.04025
R34414 VDD.n10443 VDD.n8359 0.04025
R34415 VDD.n10443 VDD.n10442 0.04025
R34416 VDD.n10442 VDD.n10441 0.04025
R34417 VDD.n10441 VDD.n8361 0.04025
R34418 VDD.n10437 VDD.n8361 0.04025
R34419 VDD.n10437 VDD.n10436 0.04025
R34420 VDD.n10436 VDD.n10435 0.04025
R34421 VDD.n10435 VDD.n8363 0.04025
R34422 VDD.n10431 VDD.n8363 0.04025
R34423 VDD.n10431 VDD.n10430 0.04025
R34424 VDD.n10430 VDD.n10429 0.04025
R34425 VDD.n10429 VDD.n8365 0.04025
R34426 VDD.n10425 VDD.n8365 0.04025
R34427 VDD.n10425 VDD.n10424 0.04025
R34428 VDD.n10424 VDD.n10423 0.04025
R34429 VDD.n10423 VDD.n8367 0.04025
R34430 VDD.n10419 VDD.n8367 0.04025
R34431 VDD.n10419 VDD.n10418 0.04025
R34432 VDD.n10418 VDD.n10417 0.04025
R34433 VDD.n10417 VDD.n8369 0.04025
R34434 VDD.n10413 VDD.n8369 0.04025
R34435 VDD.n10413 VDD.n10412 0.04025
R34436 VDD.n10412 VDD.n10411 0.04025
R34437 VDD.n10411 VDD.n8371 0.04025
R34438 VDD.n10407 VDD.n8371 0.04025
R34439 VDD.n10407 VDD.n10406 0.04025
R34440 VDD.n10406 VDD.n10405 0.04025
R34441 VDD.n10405 VDD.n8373 0.04025
R34442 VDD.n10401 VDD.n8373 0.04025
R34443 VDD.n10401 VDD.n10400 0.04025
R34444 VDD.n10400 VDD.n10399 0.04025
R34445 VDD.n10399 VDD.n8375 0.04025
R34446 VDD.n10395 VDD.n8375 0.04025
R34447 VDD.n10395 VDD.n10394 0.04025
R34448 VDD.n10394 VDD.n10393 0.04025
R34449 VDD.n10393 VDD.n8377 0.04025
R34450 VDD.n10389 VDD.n8377 0.04025
R34451 VDD.n10389 VDD.n10388 0.04025
R34452 VDD.n10388 VDD.n10387 0.04025
R34453 VDD.n10387 VDD.n8379 0.04025
R34454 VDD.n10383 VDD.n8379 0.04025
R34455 VDD.n10383 VDD.n10382 0.04025
R34456 VDD.n10382 VDD.n10381 0.04025
R34457 VDD.n10381 VDD.n8381 0.04025
R34458 VDD.n10377 VDD.n8381 0.04025
R34459 VDD.n10377 VDD.n10376 0.04025
R34460 VDD.n10376 VDD.n10375 0.04025
R34461 VDD.n10375 VDD.n8383 0.04025
R34462 VDD.n10371 VDD.n8383 0.04025
R34463 VDD.n10371 VDD.n10370 0.04025
R34464 VDD.n10370 VDD.n10369 0.04025
R34465 VDD.n10369 VDD.n8385 0.04025
R34466 VDD.n10365 VDD.n8385 0.04025
R34467 VDD.n10365 VDD.n10364 0.04025
R34468 VDD.n10364 VDD.n10363 0.04025
R34469 VDD.n10363 VDD.n8387 0.04025
R34470 VDD.n10359 VDD.n8387 0.04025
R34471 VDD.n10359 VDD.n10358 0.04025
R34472 VDD.n10358 VDD.n10357 0.04025
R34473 VDD.n10357 VDD.n8389 0.04025
R34474 VDD.n10353 VDD.n8389 0.04025
R34475 VDD.n10353 VDD.n10352 0.04025
R34476 VDD.n10352 VDD.n10351 0.04025
R34477 VDD.n10351 VDD.n8391 0.04025
R34478 VDD.n10347 VDD.n8391 0.04025
R34479 VDD.n10347 VDD.n10346 0.04025
R34480 VDD.n10346 VDD.n10345 0.04025
R34481 VDD.n10345 VDD.n8393 0.04025
R34482 VDD.n10341 VDD.n8393 0.04025
R34483 VDD.n10341 VDD.n10340 0.04025
R34484 VDD.n10340 VDD.n10339 0.04025
R34485 VDD.n10339 VDD.n8395 0.04025
R34486 VDD.n10335 VDD.n8395 0.04025
R34487 VDD.n10335 VDD.n10334 0.04025
R34488 VDD.n10334 VDD.n10333 0.04025
R34489 VDD.n10333 VDD.n8397 0.04025
R34490 VDD.n10329 VDD.n8397 0.04025
R34491 VDD.n10329 VDD.n10328 0.04025
R34492 VDD.n10328 VDD.n10327 0.04025
R34493 VDD.n10327 VDD.n8399 0.04025
R34494 VDD.n10323 VDD.n8399 0.04025
R34495 VDD.n10323 VDD.n10322 0.04025
R34496 VDD.n10322 VDD.n10321 0.04025
R34497 VDD.n10321 VDD.n8401 0.04025
R34498 VDD.n10317 VDD.n8401 0.04025
R34499 VDD.n10317 VDD.n10316 0.04025
R34500 VDD.n10316 VDD.n10315 0.04025
R34501 VDD.n10315 VDD.n8403 0.04025
R34502 VDD.n10311 VDD.n8403 0.04025
R34503 VDD.n10311 VDD.n10310 0.04025
R34504 VDD.n10310 VDD.n10309 0.04025
R34505 VDD.n10309 VDD.n8405 0.04025
R34506 VDD.n10305 VDD.n8405 0.04025
R34507 VDD.n10305 VDD.n10304 0.04025
R34508 VDD.n10304 VDD.n10303 0.04025
R34509 VDD.n10303 VDD.n8407 0.04025
R34510 VDD.n10299 VDD.n8407 0.04025
R34511 VDD.n10299 VDD.n10298 0.04025
R34512 VDD.n10298 VDD.n10297 0.04025
R34513 VDD.n10297 VDD.n8409 0.04025
R34514 VDD.n10293 VDD.n8409 0.04025
R34515 VDD.n10293 VDD.n10292 0.04025
R34516 VDD.n10292 VDD.n10291 0.04025
R34517 VDD.n10291 VDD.n8411 0.04025
R34518 VDD.n10287 VDD.n8411 0.04025
R34519 VDD.n10287 VDD.n10286 0.04025
R34520 VDD.n10286 VDD.n10285 0.04025
R34521 VDD.n10285 VDD.n8413 0.04025
R34522 VDD.n10281 VDD.n8413 0.04025
R34523 VDD.n10281 VDD.n10280 0.04025
R34524 VDD.n10280 VDD.n10279 0.04025
R34525 VDD.n10279 VDD.n8415 0.04025
R34526 VDD.n10275 VDD.n8415 0.04025
R34527 VDD.n10275 VDD.n10274 0.04025
R34528 VDD.n10274 VDD.n10273 0.04025
R34529 VDD.n10273 VDD.n8417 0.04025
R34530 VDD.n10269 VDD.n8417 0.04025
R34531 VDD.n10269 VDD.n10268 0.04025
R34532 VDD.n10268 VDD.n10267 0.04025
R34533 VDD.n10267 VDD.n8419 0.04025
R34534 VDD.n10263 VDD.n8419 0.04025
R34535 VDD.n10263 VDD.n10262 0.04025
R34536 VDD.n10262 VDD.n10261 0.04025
R34537 VDD.n10261 VDD.n8421 0.04025
R34538 VDD.n10257 VDD.n8421 0.04025
R34539 VDD.n10257 VDD.n10256 0.04025
R34540 VDD.n10256 VDD.n10255 0.04025
R34541 VDD.n10255 VDD.n8423 0.04025
R34542 VDD.n10251 VDD.n8423 0.04025
R34543 VDD.n10251 VDD.n10250 0.04025
R34544 VDD.n10250 VDD.n10249 0.04025
R34545 VDD.n10249 VDD.n8425 0.04025
R34546 VDD.n10245 VDD.n8425 0.04025
R34547 VDD.n10245 VDD.n10244 0.04025
R34548 VDD.n10244 VDD.n10243 0.04025
R34549 VDD.n10243 VDD.n8427 0.04025
R34550 VDD.n10239 VDD.n8427 0.04025
R34551 VDD.n10239 VDD.n10238 0.04025
R34552 VDD.n10238 VDD.n10237 0.04025
R34553 VDD.n10237 VDD.n8429 0.04025
R34554 VDD.n10233 VDD.n8429 0.04025
R34555 VDD.n10233 VDD.n10232 0.04025
R34556 VDD.n10232 VDD.n10231 0.04025
R34557 VDD.n10231 VDD.n8431 0.04025
R34558 VDD.n10227 VDD.n8431 0.04025
R34559 VDD.n10227 VDD.n10226 0.04025
R34560 VDD.n10226 VDD.n10225 0.04025
R34561 VDD.n10225 VDD.n8433 0.04025
R34562 VDD.n10221 VDD.n8433 0.04025
R34563 VDD.n10221 VDD.n10220 0.04025
R34564 VDD.n10220 VDD.n10219 0.04025
R34565 VDD.n10219 VDD.n8435 0.04025
R34566 VDD.n10215 VDD.n8435 0.04025
R34567 VDD.n10215 VDD.n10214 0.04025
R34568 VDD.n10214 VDD.n10213 0.04025
R34569 VDD.n10213 VDD.n8437 0.04025
R34570 VDD.n10209 VDD.n8437 0.04025
R34571 VDD.n10209 VDD.n10208 0.04025
R34572 VDD.n10208 VDD.n10207 0.04025
R34573 VDD.n10207 VDD.n8439 0.04025
R34574 VDD.n10203 VDD.n8439 0.04025
R34575 VDD.n10203 VDD.n10202 0.04025
R34576 VDD.n10202 VDD.n10201 0.04025
R34577 VDD.n10201 VDD.n8441 0.04025
R34578 VDD.n10197 VDD.n8441 0.04025
R34579 VDD.n10197 VDD.n10196 0.04025
R34580 VDD.n10196 VDD.n10195 0.04025
R34581 VDD.n10195 VDD.n8443 0.04025
R34582 VDD.n10191 VDD.n8443 0.04025
R34583 VDD.n10191 VDD.n10190 0.04025
R34584 VDD.n10190 VDD.n10189 0.04025
R34585 VDD.n10189 VDD.n8445 0.04025
R34586 VDD.n10185 VDD.n8445 0.04025
R34587 VDD.n10185 VDD.n10184 0.04025
R34588 VDD.n10184 VDD.n10183 0.04025
R34589 VDD.n10183 VDD.n8447 0.04025
R34590 VDD.n10179 VDD.n8447 0.04025
R34591 VDD.n10179 VDD.n10178 0.04025
R34592 VDD.n10178 VDD.n10177 0.04025
R34593 VDD.n10177 VDD.n8449 0.04025
R34594 VDD.n10173 VDD.n8449 0.04025
R34595 VDD.n10173 VDD.n10172 0.04025
R34596 VDD.n10172 VDD.n10171 0.04025
R34597 VDD.n10171 VDD.n8451 0.04025
R34598 VDD.n10167 VDD.n8451 0.04025
R34599 VDD.n10167 VDD.n10166 0.04025
R34600 VDD.n10166 VDD.n10165 0.04025
R34601 VDD.n10165 VDD.n8453 0.04025
R34602 VDD.n10161 VDD.n8453 0.04025
R34603 VDD.n10161 VDD.n10160 0.04025
R34604 VDD.n10160 VDD.n10159 0.04025
R34605 VDD.n10159 VDD.n8455 0.04025
R34606 VDD.n10155 VDD.n8455 0.04025
R34607 VDD.n10155 VDD.n10154 0.04025
R34608 VDD.n10154 VDD.n10153 0.04025
R34609 VDD.n10153 VDD.n8457 0.04025
R34610 VDD.n10149 VDD.n8457 0.04025
R34611 VDD.n11137 VDD.n11136 0.04025
R34612 VDD.n11137 VDD.n629 0.04025
R34613 VDD.n11141 VDD.n629 0.04025
R34614 VDD.n11142 VDD.n11141 0.04025
R34615 VDD.n11143 VDD.n11142 0.04025
R34616 VDD.n11143 VDD.n627 0.04025
R34617 VDD.n11147 VDD.n627 0.04025
R34618 VDD.n11148 VDD.n11147 0.04025
R34619 VDD.n11149 VDD.n11148 0.04025
R34620 VDD.n11149 VDD.n625 0.04025
R34621 VDD.n11153 VDD.n625 0.04025
R34622 VDD.n11154 VDD.n11153 0.04025
R34623 VDD.n11155 VDD.n11154 0.04025
R34624 VDD.n11155 VDD.n623 0.04025
R34625 VDD.n11159 VDD.n623 0.04025
R34626 VDD.n11160 VDD.n11159 0.04025
R34627 VDD.n11161 VDD.n11160 0.04025
R34628 VDD.n11161 VDD.n621 0.04025
R34629 VDD.n11165 VDD.n621 0.04025
R34630 VDD.n11166 VDD.n11165 0.04025
R34631 VDD.n11167 VDD.n11166 0.04025
R34632 VDD.n11167 VDD.n619 0.04025
R34633 VDD.n11171 VDD.n619 0.04025
R34634 VDD.n11172 VDD.n11171 0.04025
R34635 VDD.n11173 VDD.n11172 0.04025
R34636 VDD.n11173 VDD.n617 0.04025
R34637 VDD.n11177 VDD.n617 0.04025
R34638 VDD.n11178 VDD.n11177 0.04025
R34639 VDD.n11179 VDD.n11178 0.04025
R34640 VDD.n11179 VDD.n615 0.04025
R34641 VDD.n11183 VDD.n615 0.04025
R34642 VDD.n11184 VDD.n11183 0.04025
R34643 VDD.n11185 VDD.n11184 0.04025
R34644 VDD.n11185 VDD.n613 0.04025
R34645 VDD.n11189 VDD.n613 0.04025
R34646 VDD.n11190 VDD.n11189 0.04025
R34647 VDD.n11191 VDD.n11190 0.04025
R34648 VDD.n11191 VDD.n611 0.04025
R34649 VDD.n11195 VDD.n611 0.04025
R34650 VDD.n11196 VDD.n11195 0.04025
R34651 VDD.n11197 VDD.n11196 0.04025
R34652 VDD.n11197 VDD.n609 0.04025
R34653 VDD.n11201 VDD.n609 0.04025
R34654 VDD.n11202 VDD.n11201 0.04025
R34655 VDD.n11203 VDD.n11202 0.04025
R34656 VDD.n11203 VDD.n607 0.04025
R34657 VDD.n11207 VDD.n607 0.04025
R34658 VDD.n11208 VDD.n11207 0.04025
R34659 VDD.n11209 VDD.n11208 0.04025
R34660 VDD.n11209 VDD.n605 0.04025
R34661 VDD.n11213 VDD.n605 0.04025
R34662 VDD.n11214 VDD.n11213 0.04025
R34663 VDD.n11215 VDD.n11214 0.04025
R34664 VDD.n11215 VDD.n603 0.04025
R34665 VDD.n11219 VDD.n603 0.04025
R34666 VDD.n11220 VDD.n11219 0.04025
R34667 VDD.n11221 VDD.n11220 0.04025
R34668 VDD.n11221 VDD.n601 0.04025
R34669 VDD.n11225 VDD.n601 0.04025
R34670 VDD.n11226 VDD.n11225 0.04025
R34671 VDD.n11227 VDD.n11226 0.04025
R34672 VDD.n11227 VDD.n599 0.04025
R34673 VDD.n11231 VDD.n599 0.04025
R34674 VDD.n11232 VDD.n11231 0.04025
R34675 VDD.n11233 VDD.n11232 0.04025
R34676 VDD.n11233 VDD.n597 0.04025
R34677 VDD.n11237 VDD.n597 0.04025
R34678 VDD.n11238 VDD.n11237 0.04025
R34679 VDD.n11239 VDD.n11238 0.04025
R34680 VDD.n11239 VDD.n595 0.04025
R34681 VDD.n11243 VDD.n595 0.04025
R34682 VDD.n11244 VDD.n11243 0.04025
R34683 VDD.n11245 VDD.n11244 0.04025
R34684 VDD.n11245 VDD.n593 0.04025
R34685 VDD.n11249 VDD.n593 0.04025
R34686 VDD.n11250 VDD.n11249 0.04025
R34687 VDD.n11251 VDD.n11250 0.04025
R34688 VDD.n11251 VDD.n591 0.04025
R34689 VDD.n11255 VDD.n591 0.04025
R34690 VDD.n11256 VDD.n11255 0.04025
R34691 VDD.n11257 VDD.n11256 0.04025
R34692 VDD.n11257 VDD.n589 0.04025
R34693 VDD.n11261 VDD.n589 0.04025
R34694 VDD.n11262 VDD.n11261 0.04025
R34695 VDD.n11263 VDD.n11262 0.04025
R34696 VDD.n11263 VDD.n587 0.04025
R34697 VDD.n11267 VDD.n587 0.04025
R34698 VDD.n11268 VDD.n11267 0.04025
R34699 VDD.n11269 VDD.n11268 0.04025
R34700 VDD.n11269 VDD.n585 0.04025
R34701 VDD.n11273 VDD.n585 0.04025
R34702 VDD.n11274 VDD.n11273 0.04025
R34703 VDD.n11275 VDD.n11274 0.04025
R34704 VDD.n11275 VDD.n583 0.04025
R34705 VDD.n11279 VDD.n583 0.04025
R34706 VDD.n11280 VDD.n11279 0.04025
R34707 VDD.n11281 VDD.n11280 0.04025
R34708 VDD.n11281 VDD.n581 0.04025
R34709 VDD.n11285 VDD.n581 0.04025
R34710 VDD.n11286 VDD.n11285 0.04025
R34711 VDD.n11287 VDD.n11286 0.04025
R34712 VDD.n11287 VDD.n579 0.04025
R34713 VDD.n11291 VDD.n579 0.04025
R34714 VDD.n11292 VDD.n11291 0.04025
R34715 VDD.n11293 VDD.n11292 0.04025
R34716 VDD.n11293 VDD.n577 0.04025
R34717 VDD.n11297 VDD.n577 0.04025
R34718 VDD.n11298 VDD.n11297 0.04025
R34719 VDD.n11299 VDD.n11298 0.04025
R34720 VDD.n11299 VDD.n575 0.04025
R34721 VDD.n11303 VDD.n575 0.04025
R34722 VDD.n11304 VDD.n11303 0.04025
R34723 VDD.n11305 VDD.n11304 0.04025
R34724 VDD.n11305 VDD.n573 0.04025
R34725 VDD.n11309 VDD.n573 0.04025
R34726 VDD.n11310 VDD.n11309 0.04025
R34727 VDD.n11311 VDD.n11310 0.04025
R34728 VDD.n11311 VDD.n571 0.04025
R34729 VDD.n11315 VDD.n571 0.04025
R34730 VDD.n11316 VDD.n11315 0.04025
R34731 VDD.n11317 VDD.n11316 0.04025
R34732 VDD.n11317 VDD.n569 0.04025
R34733 VDD.n11321 VDD.n569 0.04025
R34734 VDD.n11322 VDD.n11321 0.04025
R34735 VDD.n11323 VDD.n11322 0.04025
R34736 VDD.n11323 VDD.n567 0.04025
R34737 VDD.n11327 VDD.n567 0.04025
R34738 VDD.n11328 VDD.n11327 0.04025
R34739 VDD.n11329 VDD.n11328 0.04025
R34740 VDD.n11329 VDD.n565 0.04025
R34741 VDD.n11333 VDD.n565 0.04025
R34742 VDD.n11334 VDD.n11333 0.04025
R34743 VDD.n11335 VDD.n11334 0.04025
R34744 VDD.n11335 VDD.n563 0.04025
R34745 VDD.n11339 VDD.n563 0.04025
R34746 VDD.n11340 VDD.n11339 0.04025
R34747 VDD.n11341 VDD.n11340 0.04025
R34748 VDD.n11341 VDD.n561 0.04025
R34749 VDD.n11345 VDD.n561 0.04025
R34750 VDD.n11346 VDD.n11345 0.04025
R34751 VDD.n11347 VDD.n11346 0.04025
R34752 VDD.n11347 VDD.n559 0.04025
R34753 VDD.n11351 VDD.n559 0.04025
R34754 VDD.n11352 VDD.n11351 0.04025
R34755 VDD.n11353 VDD.n11352 0.04025
R34756 VDD.n11353 VDD.n557 0.04025
R34757 VDD.n11357 VDD.n557 0.04025
R34758 VDD.n11358 VDD.n11357 0.04025
R34759 VDD.n11359 VDD.n11358 0.04025
R34760 VDD.n11359 VDD.n555 0.04025
R34761 VDD.n11363 VDD.n555 0.04025
R34762 VDD.n11364 VDD.n11363 0.04025
R34763 VDD.n11365 VDD.n11364 0.04025
R34764 VDD.n11365 VDD.n553 0.04025
R34765 VDD.n11369 VDD.n553 0.04025
R34766 VDD.n11370 VDD.n11369 0.04025
R34767 VDD.n11371 VDD.n11370 0.04025
R34768 VDD.n11371 VDD.n551 0.04025
R34769 VDD.n11375 VDD.n551 0.04025
R34770 VDD.n11376 VDD.n11375 0.04025
R34771 VDD.n11377 VDD.n11376 0.04025
R34772 VDD.n11377 VDD.n549 0.04025
R34773 VDD.n11381 VDD.n549 0.04025
R34774 VDD.n11382 VDD.n11381 0.04025
R34775 VDD.n11383 VDD.n11382 0.04025
R34776 VDD.n11383 VDD.n547 0.04025
R34777 VDD.n11387 VDD.n547 0.04025
R34778 VDD.n11388 VDD.n11387 0.04025
R34779 VDD.n11389 VDD.n11388 0.04025
R34780 VDD.n11389 VDD.n545 0.04025
R34781 VDD.n11393 VDD.n545 0.04025
R34782 VDD.n11394 VDD.n11393 0.04025
R34783 VDD.n11395 VDD.n11394 0.04025
R34784 VDD.n11395 VDD.n543 0.04025
R34785 VDD.n11399 VDD.n543 0.04025
R34786 VDD.n11400 VDD.n11399 0.04025
R34787 VDD.n11401 VDD.n11400 0.04025
R34788 VDD.n11401 VDD.n541 0.04025
R34789 VDD.n11405 VDD.n541 0.04025
R34790 VDD.n11406 VDD.n11405 0.04025
R34791 VDD.n11407 VDD.n11406 0.04025
R34792 VDD.n11407 VDD.n539 0.04025
R34793 VDD.n11411 VDD.n539 0.04025
R34794 VDD.n11412 VDD.n11411 0.04025
R34795 VDD.n11413 VDD.n11412 0.04025
R34796 VDD.n11413 VDD.n537 0.04025
R34797 VDD.n11417 VDD.n537 0.04025
R34798 VDD.n11418 VDD.n11417 0.04025
R34799 VDD.n11419 VDD.n11418 0.04025
R34800 VDD.n11419 VDD.n535 0.04025
R34801 VDD.n11423 VDD.n535 0.04025
R34802 VDD.n11424 VDD.n11423 0.04025
R34803 VDD.n11425 VDD.n11424 0.04025
R34804 VDD.n11425 VDD.n533 0.04025
R34805 VDD.n11429 VDD.n533 0.04025
R34806 VDD.n11430 VDD.n11429 0.04025
R34807 VDD.n11431 VDD.n11430 0.04025
R34808 VDD.n11431 VDD.n531 0.04025
R34809 VDD.n11435 VDD.n531 0.04025
R34810 VDD.n11436 VDD.n11435 0.04025
R34811 VDD.n11437 VDD.n11436 0.04025
R34812 VDD.n11437 VDD.n529 0.04025
R34813 VDD.n11441 VDD.n529 0.04025
R34814 VDD.n11442 VDD.n11441 0.04025
R34815 VDD.n11443 VDD.n11442 0.04025
R34816 VDD.n11443 VDD.n527 0.04025
R34817 VDD.n11447 VDD.n527 0.04025
R34818 VDD.n11448 VDD.n11447 0.04025
R34819 VDD.n11449 VDD.n11448 0.04025
R34820 VDD.n11449 VDD.n525 0.04025
R34821 VDD.n11453 VDD.n525 0.04025
R34822 VDD.n11454 VDD.n11453 0.04025
R34823 VDD.n11455 VDD.n11454 0.04025
R34824 VDD.n11455 VDD.n523 0.04025
R34825 VDD.n11459 VDD.n523 0.04025
R34826 VDD.n11460 VDD.n11459 0.04025
R34827 VDD.n11461 VDD.n11460 0.04025
R34828 VDD.n11461 VDD.n521 0.04025
R34829 VDD.n11465 VDD.n521 0.04025
R34830 VDD.n11466 VDD.n11465 0.04025
R34831 VDD.n11467 VDD.n11466 0.04025
R34832 VDD.n11467 VDD.n519 0.04025
R34833 VDD.n11471 VDD.n519 0.04025
R34834 VDD.n11472 VDD.n11471 0.04025
R34835 VDD.n11473 VDD.n11472 0.04025
R34836 VDD.n11473 VDD.n517 0.04025
R34837 VDD.n11477 VDD.n517 0.04025
R34838 VDD.n11478 VDD.n11477 0.04025
R34839 VDD.n11479 VDD.n11478 0.04025
R34840 VDD.n11479 VDD.n515 0.04025
R34841 VDD.n11483 VDD.n515 0.04025
R34842 VDD.n11484 VDD.n11483 0.04025
R34843 VDD.n11485 VDD.n11484 0.04025
R34844 VDD.n11485 VDD.n513 0.04025
R34845 VDD.n11489 VDD.n513 0.04025
R34846 VDD.n11490 VDD.n11489 0.04025
R34847 VDD.n11491 VDD.n11490 0.04025
R34848 VDD.n11491 VDD.n511 0.04025
R34849 VDD.n11495 VDD.n511 0.04025
R34850 VDD.n11496 VDD.n11495 0.04025
R34851 VDD.n11497 VDD.n11496 0.04025
R34852 VDD.n11497 VDD.n509 0.04025
R34853 VDD.n11501 VDD.n509 0.04025
R34854 VDD.n11502 VDD.n11501 0.04025
R34855 VDD.n11503 VDD.n11502 0.04025
R34856 VDD.n11503 VDD.n507 0.04025
R34857 VDD.n11507 VDD.n507 0.04025
R34858 VDD.n11508 VDD.n11507 0.04025
R34859 VDD.n11509 VDD.n11508 0.04025
R34860 VDD.n11509 VDD.n505 0.04025
R34861 VDD.n11513 VDD.n505 0.04025
R34862 VDD.n11514 VDD.n11513 0.04025
R34863 VDD.n11515 VDD.n11514 0.04025
R34864 VDD.n11515 VDD.n503 0.04025
R34865 VDD.n11519 VDD.n503 0.04025
R34866 VDD.n11520 VDD.n11519 0.04025
R34867 VDD.n11521 VDD.n11520 0.04025
R34868 VDD.n11521 VDD.n501 0.04025
R34869 VDD.n11525 VDD.n501 0.04025
R34870 VDD.n11526 VDD.n11525 0.04025
R34871 VDD.n11527 VDD.n11526 0.04025
R34872 VDD.n11527 VDD.n499 0.04025
R34873 VDD.n11531 VDD.n499 0.04025
R34874 VDD.n11532 VDD.n11531 0.04025
R34875 VDD.n11533 VDD.n11532 0.04025
R34876 VDD.n11533 VDD.n497 0.04025
R34877 VDD.n11537 VDD.n497 0.04025
R34878 VDD.n11538 VDD.n11537 0.04025
R34879 VDD.n11539 VDD.n11538 0.04025
R34880 VDD.n11539 VDD.n495 0.04025
R34881 VDD.n11543 VDD.n495 0.04025
R34882 VDD.n11544 VDD.n11543 0.04025
R34883 VDD.n11545 VDD.n11544 0.04025
R34884 VDD.n11545 VDD.n493 0.04025
R34885 VDD.n11549 VDD.n493 0.04025
R34886 VDD.n11550 VDD.n11549 0.04025
R34887 VDD.n11551 VDD.n11550 0.04025
R34888 VDD.n11551 VDD.n491 0.04025
R34889 VDD.n11555 VDD.n491 0.04025
R34890 VDD.n11556 VDD.n11555 0.04025
R34891 VDD.n11557 VDD.n11556 0.04025
R34892 VDD.n11557 VDD.n489 0.04025
R34893 VDD.n11561 VDD.n489 0.04025
R34894 VDD.n11562 VDD.n11561 0.04025
R34895 VDD.n11563 VDD.n11562 0.04025
R34896 VDD.n11563 VDD.n487 0.04025
R34897 VDD.n11567 VDD.n487 0.04025
R34898 VDD.n11568 VDD.n11567 0.04025
R34899 VDD.n11569 VDD.n11568 0.04025
R34900 VDD.n11569 VDD.n485 0.04025
R34901 VDD.n11573 VDD.n485 0.04025
R34902 VDD.n11574 VDD.n11573 0.04025
R34903 VDD.n11575 VDD.n11574 0.04025
R34904 VDD.n11575 VDD.n483 0.04025
R34905 VDD.n11579 VDD.n483 0.04025
R34906 VDD.n11580 VDD.n11579 0.04025
R34907 VDD.n11581 VDD.n11580 0.04025
R34908 VDD.n11581 VDD.n481 0.04025
R34909 VDD.n11585 VDD.n481 0.04025
R34910 VDD.n11586 VDD.n11585 0.04025
R34911 VDD.n11587 VDD.n11586 0.04025
R34912 VDD.n11587 VDD.n479 0.04025
R34913 VDD.n11591 VDD.n479 0.04025
R34914 VDD.n11592 VDD.n11591 0.04025
R34915 VDD.n11593 VDD.n11592 0.04025
R34916 VDD.n11593 VDD.n477 0.04025
R34917 VDD.n11597 VDD.n477 0.04025
R34918 VDD.n11598 VDD.n11597 0.04025
R34919 VDD.n11599 VDD.n11598 0.04025
R34920 VDD.n11599 VDD.n475 0.04025
R34921 VDD.n11603 VDD.n475 0.04025
R34922 VDD.n11604 VDD.n11603 0.04025
R34923 VDD.n11605 VDD.n11604 0.04025
R34924 VDD.n11605 VDD.n473 0.04025
R34925 VDD.n11609 VDD.n473 0.04025
R34926 VDD.n11610 VDD.n11609 0.04025
R34927 VDD.n11611 VDD.n11610 0.04025
R34928 VDD.n11611 VDD.n471 0.04025
R34929 VDD.n11615 VDD.n471 0.04025
R34930 VDD.n11616 VDD.n11615 0.04025
R34931 VDD.n11617 VDD.n11616 0.04025
R34932 VDD.n11617 VDD.n469 0.04025
R34933 VDD.n11621 VDD.n469 0.04025
R34934 VDD.n11622 VDD.n11621 0.04025
R34935 VDD.n11623 VDD.n11622 0.04025
R34936 VDD.n11623 VDD.n467 0.04025
R34937 VDD.n11627 VDD.n467 0.04025
R34938 VDD.n11628 VDD.n11627 0.04025
R34939 VDD.n11629 VDD.n11628 0.04025
R34940 VDD.n11629 VDD.n465 0.04025
R34941 VDD.n11633 VDD.n465 0.04025
R34942 VDD.n11634 VDD.n11633 0.04025
R34943 VDD.n11635 VDD.n11634 0.04025
R34944 VDD.n11635 VDD.n463 0.04025
R34945 VDD.n11639 VDD.n463 0.04025
R34946 VDD.n11640 VDD.n11639 0.04025
R34947 VDD.n11641 VDD.n11640 0.04025
R34948 VDD.n11641 VDD.n461 0.04025
R34949 VDD.n11645 VDD.n461 0.04025
R34950 VDD.n11646 VDD.n11645 0.04025
R34951 VDD.n11647 VDD.n11646 0.04025
R34952 VDD.n11647 VDD.n459 0.04025
R34953 VDD.n11651 VDD.n459 0.04025
R34954 VDD.n11652 VDD.n11651 0.04025
R34955 VDD.n11653 VDD.n11652 0.04025
R34956 VDD.n11653 VDD.n457 0.04025
R34957 VDD.n11657 VDD.n457 0.04025
R34958 VDD.n11658 VDD.n11657 0.04025
R34959 VDD.n11659 VDD.n11658 0.04025
R34960 VDD.n11659 VDD.n455 0.04025
R34961 VDD.n11663 VDD.n455 0.04025
R34962 VDD.n11664 VDD.n11663 0.04025
R34963 VDD.n11665 VDD.n11664 0.04025
R34964 VDD.n11665 VDD.n453 0.04025
R34965 VDD.n11669 VDD.n453 0.04025
R34966 VDD.n11670 VDD.n11669 0.04025
R34967 VDD.n11671 VDD.n11670 0.04025
R34968 VDD.n11671 VDD.n451 0.04025
R34969 VDD.n11675 VDD.n451 0.04025
R34970 VDD.n11676 VDD.n11675 0.04025
R34971 VDD.n11677 VDD.n11676 0.04025
R34972 VDD.n11677 VDD.n449 0.04025
R34973 VDD.n11681 VDD.n449 0.04025
R34974 VDD.n11682 VDD.n11681 0.04025
R34975 VDD.n11683 VDD.n11682 0.04025
R34976 VDD.n11683 VDD.n447 0.04025
R34977 VDD.n11687 VDD.n447 0.04025
R34978 VDD.n11688 VDD.n11687 0.04025
R34979 VDD.n11689 VDD.n11688 0.04025
R34980 VDD.n11689 VDD.n445 0.04025
R34981 VDD.n11693 VDD.n445 0.04025
R34982 VDD.n11694 VDD.n11693 0.04025
R34983 VDD.n11695 VDD.n11694 0.04025
R34984 VDD.n11695 VDD.n443 0.04025
R34985 VDD.n11699 VDD.n443 0.04025
R34986 VDD.n11700 VDD.n11699 0.04025
R34987 VDD.n11701 VDD.n11700 0.04025
R34988 VDD.n11701 VDD.n441 0.04025
R34989 VDD.n11705 VDD.n441 0.04025
R34990 VDD.n11706 VDD.n11705 0.04025
R34991 VDD.n11707 VDD.n11706 0.04025
R34992 VDD.n11707 VDD.n439 0.04025
R34993 VDD.n11711 VDD.n439 0.04025
R34994 VDD.n11712 VDD.n11711 0.04025
R34995 VDD.n11713 VDD.n11712 0.04025
R34996 VDD.n11713 VDD.n437 0.04025
R34997 VDD.n11717 VDD.n437 0.04025
R34998 VDD.n11718 VDD.n11717 0.04025
R34999 VDD.n11719 VDD.n11718 0.04025
R35000 VDD.n11719 VDD.n435 0.04025
R35001 VDD.n11723 VDD.n435 0.04025
R35002 VDD.n11724 VDD.n11723 0.04025
R35003 VDD.n11725 VDD.n11724 0.04025
R35004 VDD.n11725 VDD.n433 0.04025
R35005 VDD.n11729 VDD.n433 0.04025
R35006 VDD.n11730 VDD.n11729 0.04025
R35007 VDD.n11731 VDD.n11730 0.04025
R35008 VDD.n11731 VDD.n431 0.04025
R35009 VDD.n11735 VDD.n431 0.04025
R35010 VDD.n11736 VDD.n11735 0.04025
R35011 VDD.n11737 VDD.n11736 0.04025
R35012 VDD.n11737 VDD.n429 0.04025
R35013 VDD.n11741 VDD.n429 0.04025
R35014 VDD.n11742 VDD.n11741 0.04025
R35015 VDD.n11743 VDD.n11742 0.04025
R35016 VDD.n11743 VDD.n427 0.04025
R35017 VDD.n11747 VDD.n427 0.04025
R35018 VDD.n11748 VDD.n11747 0.04025
R35019 VDD.n11749 VDD.n11748 0.04025
R35020 VDD.n11749 VDD.n425 0.04025
R35021 VDD.n11753 VDD.n425 0.04025
R35022 VDD.n11754 VDD.n11753 0.04025
R35023 VDD.n11755 VDD.n11754 0.04025
R35024 VDD.n11755 VDD.n423 0.04025
R35025 VDD.n11759 VDD.n423 0.04025
R35026 VDD.n11760 VDD.n11759 0.04025
R35027 VDD.n11761 VDD.n11760 0.04025
R35028 VDD.n11761 VDD.n421 0.04025
R35029 VDD.n11765 VDD.n421 0.04025
R35030 VDD.n11766 VDD.n11765 0.04025
R35031 VDD.n11767 VDD.n11766 0.04025
R35032 VDD.n11767 VDD.n419 0.04025
R35033 VDD.n11771 VDD.n419 0.04025
R35034 VDD.n11772 VDD.n11771 0.04025
R35035 VDD.n11773 VDD.n11772 0.04025
R35036 VDD.n11773 VDD.n417 0.04025
R35037 VDD.n11777 VDD.n417 0.04025
R35038 VDD.n11778 VDD.n11777 0.04025
R35039 VDD.n11779 VDD.n11778 0.04025
R35040 VDD.n11779 VDD.n415 0.04025
R35041 VDD.n11783 VDD.n415 0.04025
R35042 VDD.n11784 VDD.n11783 0.04025
R35043 VDD.n11785 VDD.n11784 0.04025
R35044 VDD.n11785 VDD.n413 0.04025
R35045 VDD.n11789 VDD.n413 0.04025
R35046 VDD.n11790 VDD.n11789 0.04025
R35047 VDD.n11791 VDD.n11790 0.04025
R35048 VDD.n11791 VDD.n411 0.04025
R35049 VDD.n11795 VDD.n411 0.04025
R35050 VDD.n11796 VDD.n11795 0.04025
R35051 VDD.n11797 VDD.n11796 0.04025
R35052 VDD.n11797 VDD.n409 0.04025
R35053 VDD.n11801 VDD.n409 0.04025
R35054 VDD.n11802 VDD.n11801 0.04025
R35055 VDD.n11803 VDD.n11802 0.04025
R35056 VDD.n11803 VDD.n407 0.04025
R35057 VDD.n11807 VDD.n407 0.04025
R35058 VDD.n11808 VDD.n11807 0.04025
R35059 VDD.n11809 VDD.n11808 0.04025
R35060 VDD.n11809 VDD.n405 0.04025
R35061 VDD.n3629 VDD.n2746 0.04025
R35062 VDD.n3625 VDD.n2746 0.04025
R35063 VDD.n3625 VDD.n3624 0.04025
R35064 VDD.n3624 VDD.n3623 0.04025
R35065 VDD.n3623 VDD.n2748 0.04025
R35066 VDD.n3619 VDD.n2748 0.04025
R35067 VDD.n3619 VDD.n3618 0.04025
R35068 VDD.n3618 VDD.n3617 0.04025
R35069 VDD.n3617 VDD.n2750 0.04025
R35070 VDD.n3613 VDD.n2750 0.04025
R35071 VDD.n3613 VDD.n3612 0.04025
R35072 VDD.n3612 VDD.n3611 0.04025
R35073 VDD.n3611 VDD.n2752 0.04025
R35074 VDD.n3607 VDD.n2752 0.04025
R35075 VDD.n3607 VDD.n3606 0.04025
R35076 VDD.n3606 VDD.n3605 0.04025
R35077 VDD.n3605 VDD.n2754 0.04025
R35078 VDD.n3601 VDD.n2754 0.04025
R35079 VDD.n3601 VDD.n3600 0.04025
R35080 VDD.n3600 VDD.n3599 0.04025
R35081 VDD.n3599 VDD.n2756 0.04025
R35082 VDD.n3595 VDD.n2756 0.04025
R35083 VDD.n3595 VDD.n3594 0.04025
R35084 VDD.n3594 VDD.n3593 0.04025
R35085 VDD.n3593 VDD.n2758 0.04025
R35086 VDD.n3589 VDD.n2758 0.04025
R35087 VDD.n3589 VDD.n3588 0.04025
R35088 VDD.n3588 VDD.n3587 0.04025
R35089 VDD.n3587 VDD.n2760 0.04025
R35090 VDD.n3583 VDD.n2760 0.04025
R35091 VDD.n3583 VDD.n3582 0.04025
R35092 VDD.n3582 VDD.n3581 0.04025
R35093 VDD.n3581 VDD.n2762 0.04025
R35094 VDD.n3577 VDD.n2762 0.04025
R35095 VDD.n3577 VDD.n3576 0.04025
R35096 VDD.n3576 VDD.n3575 0.04025
R35097 VDD.n3575 VDD.n2764 0.04025
R35098 VDD.n3571 VDD.n2764 0.04025
R35099 VDD.n3571 VDD.n3570 0.04025
R35100 VDD.n3570 VDD.n3569 0.04025
R35101 VDD.n3569 VDD.n2766 0.04025
R35102 VDD.n3565 VDD.n2766 0.04025
R35103 VDD.n3565 VDD.n3564 0.04025
R35104 VDD.n3564 VDD.n3563 0.04025
R35105 VDD.n3563 VDD.n2768 0.04025
R35106 VDD.n3559 VDD.n2768 0.04025
R35107 VDD.n3559 VDD.n3558 0.04025
R35108 VDD.n3558 VDD.n3557 0.04025
R35109 VDD.n3557 VDD.n2770 0.04025
R35110 VDD.n3553 VDD.n2770 0.04025
R35111 VDD.n3553 VDD.n3552 0.04025
R35112 VDD.n3552 VDD.n3551 0.04025
R35113 VDD.n3551 VDD.n2772 0.04025
R35114 VDD.n3547 VDD.n2772 0.04025
R35115 VDD.n3547 VDD.n3546 0.04025
R35116 VDD.n3546 VDD.n3545 0.04025
R35117 VDD.n3545 VDD.n2774 0.04025
R35118 VDD.n3541 VDD.n2774 0.04025
R35119 VDD.n3541 VDD.n3540 0.04025
R35120 VDD.n3540 VDD.n3539 0.04025
R35121 VDD.n3539 VDD.n2776 0.04025
R35122 VDD.n3535 VDD.n2776 0.04025
R35123 VDD.n3535 VDD.n3534 0.04025
R35124 VDD.n3534 VDD.n3533 0.04025
R35125 VDD.n3533 VDD.n2778 0.04025
R35126 VDD.n3529 VDD.n2778 0.04025
R35127 VDD.n3529 VDD.n3528 0.04025
R35128 VDD.n3528 VDD.n3527 0.04025
R35129 VDD.n3527 VDD.n2780 0.04025
R35130 VDD.n3523 VDD.n2780 0.04025
R35131 VDD.n3523 VDD.n3522 0.04025
R35132 VDD.n3522 VDD.n3521 0.04025
R35133 VDD.n3521 VDD.n2782 0.04025
R35134 VDD.n3517 VDD.n2782 0.04025
R35135 VDD.n3517 VDD.n3516 0.04025
R35136 VDD.n3516 VDD.n3515 0.04025
R35137 VDD.n3515 VDD.n2784 0.04025
R35138 VDD.n3511 VDD.n2784 0.04025
R35139 VDD.n3511 VDD.n3510 0.04025
R35140 VDD.n3510 VDD.n3509 0.04025
R35141 VDD.n3509 VDD.n2786 0.04025
R35142 VDD.n3505 VDD.n2786 0.04025
R35143 VDD.n3505 VDD.n3504 0.04025
R35144 VDD.n3504 VDD.n3503 0.04025
R35145 VDD.n3503 VDD.n2788 0.04025
R35146 VDD.n3499 VDD.n2788 0.04025
R35147 VDD.n3499 VDD.n3498 0.04025
R35148 VDD.n3498 VDD.n3497 0.04025
R35149 VDD.n3497 VDD.n2790 0.04025
R35150 VDD.n3493 VDD.n2790 0.04025
R35151 VDD.n3493 VDD.n3492 0.04025
R35152 VDD.n3492 VDD.n3491 0.04025
R35153 VDD.n3491 VDD.n2792 0.04025
R35154 VDD.n3487 VDD.n2792 0.04025
R35155 VDD.n3487 VDD.n3486 0.04025
R35156 VDD.n3486 VDD.n3485 0.04025
R35157 VDD.n3485 VDD.n2794 0.04025
R35158 VDD.n3481 VDD.n2794 0.04025
R35159 VDD.n3481 VDD.n3480 0.04025
R35160 VDD.n3480 VDD.n3479 0.04025
R35161 VDD.n3479 VDD.n2796 0.04025
R35162 VDD.n3475 VDD.n2796 0.04025
R35163 VDD.n3475 VDD.n3474 0.04025
R35164 VDD.n3474 VDD.n3473 0.04025
R35165 VDD.n3473 VDD.n2798 0.04025
R35166 VDD.n3469 VDD.n2798 0.04025
R35167 VDD.n3469 VDD.n3468 0.04025
R35168 VDD.n3468 VDD.n3467 0.04025
R35169 VDD.n3467 VDD.n2800 0.04025
R35170 VDD.n3463 VDD.n2800 0.04025
R35171 VDD.n3463 VDD.n3462 0.04025
R35172 VDD.n3462 VDD.n3461 0.04025
R35173 VDD.n3461 VDD.n2802 0.04025
R35174 VDD.n3457 VDD.n2802 0.04025
R35175 VDD.n3457 VDD.n3456 0.04025
R35176 VDD.n3456 VDD.n3455 0.04025
R35177 VDD.n3455 VDD.n2804 0.04025
R35178 VDD.n3451 VDD.n2804 0.04025
R35179 VDD.n3451 VDD.n3450 0.04025
R35180 VDD.n3450 VDD.n3449 0.04025
R35181 VDD.n3449 VDD.n2806 0.04025
R35182 VDD.n3445 VDD.n2806 0.04025
R35183 VDD.n3445 VDD.n3444 0.04025
R35184 VDD.n3444 VDD.n3443 0.04025
R35185 VDD.n3443 VDD.n2808 0.04025
R35186 VDD.n3439 VDD.n2808 0.04025
R35187 VDD.n3439 VDD.n3438 0.04025
R35188 VDD.n3438 VDD.n3437 0.04025
R35189 VDD.n3437 VDD.n2810 0.04025
R35190 VDD.n3433 VDD.n2810 0.04025
R35191 VDD.n3433 VDD.n3432 0.04025
R35192 VDD.n3432 VDD.n3431 0.04025
R35193 VDD.n3431 VDD.n2812 0.04025
R35194 VDD.n3427 VDD.n2812 0.04025
R35195 VDD.n3427 VDD.n3426 0.04025
R35196 VDD.n3426 VDD.n3425 0.04025
R35197 VDD.n3425 VDD.n2814 0.04025
R35198 VDD.n3421 VDD.n2814 0.04025
R35199 VDD.n3421 VDD.n3420 0.04025
R35200 VDD.n3420 VDD.n3419 0.04025
R35201 VDD.n3419 VDD.n2816 0.04025
R35202 VDD.n3415 VDD.n2816 0.04025
R35203 VDD.n3415 VDD.n3414 0.04025
R35204 VDD.n3414 VDD.n3413 0.04025
R35205 VDD.n3413 VDD.n2818 0.04025
R35206 VDD.n3409 VDD.n2818 0.04025
R35207 VDD.n3409 VDD.n3408 0.04025
R35208 VDD.n3408 VDD.n3407 0.04025
R35209 VDD.n3407 VDD.n2820 0.04025
R35210 VDD.n3403 VDD.n2820 0.04025
R35211 VDD.n3403 VDD.n3402 0.04025
R35212 VDD.n3402 VDD.n3401 0.04025
R35213 VDD.n3401 VDD.n2822 0.04025
R35214 VDD.n3397 VDD.n2822 0.04025
R35215 VDD.n3397 VDD.n3396 0.04025
R35216 VDD.n3396 VDD.n3395 0.04025
R35217 VDD.n3395 VDD.n2824 0.04025
R35218 VDD.n3391 VDD.n2824 0.04025
R35219 VDD.n3391 VDD.n3390 0.04025
R35220 VDD.n3390 VDD.n3389 0.04025
R35221 VDD.n3389 VDD.n2826 0.04025
R35222 VDD.n3385 VDD.n2826 0.04025
R35223 VDD.n3385 VDD.n3384 0.04025
R35224 VDD.n3384 VDD.n3383 0.04025
R35225 VDD.n3383 VDD.n2828 0.04025
R35226 VDD.n3379 VDD.n2828 0.04025
R35227 VDD.n3379 VDD.n3378 0.04025
R35228 VDD.n3378 VDD.n3377 0.04025
R35229 VDD.n3377 VDD.n2830 0.04025
R35230 VDD.n3373 VDD.n2830 0.04025
R35231 VDD.n3373 VDD.n3372 0.04025
R35232 VDD.n3372 VDD.n3371 0.04025
R35233 VDD.n3371 VDD.n2832 0.04025
R35234 VDD.n3367 VDD.n2832 0.04025
R35235 VDD.n3367 VDD.n3366 0.04025
R35236 VDD.n3366 VDD.n3365 0.04025
R35237 VDD.n3365 VDD.n2834 0.04025
R35238 VDD.n3361 VDD.n2834 0.04025
R35239 VDD.n3361 VDD.n3360 0.04025
R35240 VDD.n3360 VDD.n3359 0.04025
R35241 VDD.n3359 VDD.n2836 0.04025
R35242 VDD.n3355 VDD.n2836 0.04025
R35243 VDD.n3355 VDD.n3354 0.04025
R35244 VDD.n3354 VDD.n3353 0.04025
R35245 VDD.n3353 VDD.n2838 0.04025
R35246 VDD.n3349 VDD.n2838 0.04025
R35247 VDD.n3349 VDD.n3348 0.04025
R35248 VDD.n3348 VDD.n3347 0.04025
R35249 VDD.n3347 VDD.n2840 0.04025
R35250 VDD.n3343 VDD.n2840 0.04025
R35251 VDD.n3343 VDD.n3342 0.04025
R35252 VDD.n3342 VDD.n3341 0.04025
R35253 VDD.n3341 VDD.n2842 0.04025
R35254 VDD.n3337 VDD.n2842 0.04025
R35255 VDD.n3337 VDD.n3336 0.04025
R35256 VDD.n3336 VDD.n3335 0.04025
R35257 VDD.n3335 VDD.n2844 0.04025
R35258 VDD.n3331 VDD.n2844 0.04025
R35259 VDD.n3331 VDD.n3330 0.04025
R35260 VDD.n3330 VDD.n3329 0.04025
R35261 VDD.n3329 VDD.n2846 0.04025
R35262 VDD.n3325 VDD.n2846 0.04025
R35263 VDD.n3325 VDD.n3324 0.04025
R35264 VDD.n3324 VDD.n3323 0.04025
R35265 VDD.n3323 VDD.n2848 0.04025
R35266 VDD.n3319 VDD.n2848 0.04025
R35267 VDD.n3319 VDD.n3318 0.04025
R35268 VDD.n3318 VDD.n3317 0.04025
R35269 VDD.n3317 VDD.n2850 0.04025
R35270 VDD.n3313 VDD.n2850 0.04025
R35271 VDD.n3313 VDD.n3312 0.04025
R35272 VDD.n3312 VDD.n3311 0.04025
R35273 VDD.n3311 VDD.n2852 0.04025
R35274 VDD.n3307 VDD.n2852 0.04025
R35275 VDD.n3307 VDD.n3306 0.04025
R35276 VDD.n3306 VDD.n3305 0.04025
R35277 VDD.n3305 VDD.n2854 0.04025
R35278 VDD.n3301 VDD.n2854 0.04025
R35279 VDD.n3301 VDD.n3300 0.04025
R35280 VDD.n3300 VDD.n3299 0.04025
R35281 VDD.n3299 VDD.n2856 0.04025
R35282 VDD.n3295 VDD.n2856 0.04025
R35283 VDD.n3295 VDD.n3294 0.04025
R35284 VDD.n3294 VDD.n3293 0.04025
R35285 VDD.n3293 VDD.n2858 0.04025
R35286 VDD.n3289 VDD.n2858 0.04025
R35287 VDD.n3289 VDD.n3288 0.04025
R35288 VDD.n3288 VDD.n3287 0.04025
R35289 VDD.n3287 VDD.n2860 0.04025
R35290 VDD.n3283 VDD.n2860 0.04025
R35291 VDD.n3283 VDD.n3282 0.04025
R35292 VDD.n3282 VDD.n3281 0.04025
R35293 VDD.n3281 VDD.n2862 0.04025
R35294 VDD.n3277 VDD.n2862 0.04025
R35295 VDD.n3277 VDD.n3276 0.04025
R35296 VDD.n3276 VDD.n3275 0.04025
R35297 VDD.n3275 VDD.n2864 0.04025
R35298 VDD.n3271 VDD.n2864 0.04025
R35299 VDD.n3271 VDD.n3270 0.04025
R35300 VDD.n3270 VDD.n3269 0.04025
R35301 VDD.n3269 VDD.n2866 0.04025
R35302 VDD.n3265 VDD.n2866 0.04025
R35303 VDD.n3265 VDD.n3264 0.04025
R35304 VDD.n3264 VDD.n3263 0.04025
R35305 VDD.n3263 VDD.n2868 0.04025
R35306 VDD.n3259 VDD.n2868 0.04025
R35307 VDD.n3259 VDD.n3258 0.04025
R35308 VDD.n3258 VDD.n3257 0.04025
R35309 VDD.n3257 VDD.n2870 0.04025
R35310 VDD.n3253 VDD.n2870 0.04025
R35311 VDD.n3253 VDD.n3252 0.04025
R35312 VDD.n3252 VDD.n3251 0.04025
R35313 VDD.n3251 VDD.n2872 0.04025
R35314 VDD.n3247 VDD.n2872 0.04025
R35315 VDD.n3247 VDD.n3246 0.04025
R35316 VDD.n3246 VDD.n3245 0.04025
R35317 VDD.n3245 VDD.n2874 0.04025
R35318 VDD.n3241 VDD.n2874 0.04025
R35319 VDD.n3241 VDD.n3240 0.04025
R35320 VDD.n3240 VDD.n3239 0.04025
R35321 VDD.n3239 VDD.n2876 0.04025
R35322 VDD.n3235 VDD.n2876 0.04025
R35323 VDD.n3235 VDD.n3234 0.04025
R35324 VDD.n3234 VDD.n3233 0.04025
R35325 VDD.n3233 VDD.n2878 0.04025
R35326 VDD.n3229 VDD.n2878 0.04025
R35327 VDD.n3229 VDD.n3228 0.04025
R35328 VDD.n3228 VDD.n3227 0.04025
R35329 VDD.n3227 VDD.n2880 0.04025
R35330 VDD.n3223 VDD.n2880 0.04025
R35331 VDD.n3223 VDD.n3222 0.04025
R35332 VDD.n3222 VDD.n3221 0.04025
R35333 VDD.n3221 VDD.n2882 0.04025
R35334 VDD.n3217 VDD.n2882 0.04025
R35335 VDD.n3217 VDD.n3216 0.04025
R35336 VDD.n3216 VDD.n3215 0.04025
R35337 VDD.n3215 VDD.n2884 0.04025
R35338 VDD.n3211 VDD.n2884 0.04025
R35339 VDD.n3211 VDD.n3210 0.04025
R35340 VDD.n3210 VDD.n3209 0.04025
R35341 VDD.n3209 VDD.n2886 0.04025
R35342 VDD.n3205 VDD.n2886 0.04025
R35343 VDD.n3205 VDD.n3204 0.04025
R35344 VDD.n3204 VDD.n3203 0.04025
R35345 VDD.n3203 VDD.n2888 0.04025
R35346 VDD.n3199 VDD.n2888 0.04025
R35347 VDD.n3199 VDD.n3198 0.04025
R35348 VDD.n3198 VDD.n3197 0.04025
R35349 VDD.n3197 VDD.n2890 0.04025
R35350 VDD.n3193 VDD.n2890 0.04025
R35351 VDD.n3193 VDD.n3192 0.04025
R35352 VDD.n3192 VDD.n3191 0.04025
R35353 VDD.n3191 VDD.n2892 0.04025
R35354 VDD.n3187 VDD.n2892 0.04025
R35355 VDD.n3187 VDD.n3186 0.04025
R35356 VDD.n3186 VDD.n3185 0.04025
R35357 VDD.n3185 VDD.n2894 0.04025
R35358 VDD.n3181 VDD.n2894 0.04025
R35359 VDD.n3181 VDD.n3180 0.04025
R35360 VDD.n3180 VDD.n3179 0.04025
R35361 VDD.n3179 VDD.n2896 0.04025
R35362 VDD.n3175 VDD.n2896 0.04025
R35363 VDD.n3175 VDD.n3174 0.04025
R35364 VDD.n3174 VDD.n3173 0.04025
R35365 VDD.n3173 VDD.n2898 0.04025
R35366 VDD.n3169 VDD.n2898 0.04025
R35367 VDD.n3169 VDD.n3168 0.04025
R35368 VDD.n3168 VDD.n3167 0.04025
R35369 VDD.n3167 VDD.n2900 0.04025
R35370 VDD.n3163 VDD.n2900 0.04025
R35371 VDD.n3163 VDD.n3162 0.04025
R35372 VDD.n3162 VDD.n3161 0.04025
R35373 VDD.n3161 VDD.n2902 0.04025
R35374 VDD.n3157 VDD.n2902 0.04025
R35375 VDD.n3157 VDD.n3156 0.04025
R35376 VDD.n3156 VDD.n3155 0.04025
R35377 VDD.n3155 VDD.n2904 0.04025
R35378 VDD.n3151 VDD.n2904 0.04025
R35379 VDD.n3151 VDD.n3150 0.04025
R35380 VDD.n3150 VDD.n3149 0.04025
R35381 VDD.n3149 VDD.n2906 0.04025
R35382 VDD.n3145 VDD.n2906 0.04025
R35383 VDD.n3145 VDD.n3144 0.04025
R35384 VDD.n3144 VDD.n3143 0.04025
R35385 VDD.n3143 VDD.n2908 0.04025
R35386 VDD.n3139 VDD.n2908 0.04025
R35387 VDD.n3139 VDD.n3138 0.04025
R35388 VDD.n3138 VDD.n3137 0.04025
R35389 VDD.n3137 VDD.n2910 0.04025
R35390 VDD.n3133 VDD.n2910 0.04025
R35391 VDD.n3133 VDD.n3132 0.04025
R35392 VDD.n3132 VDD.n3131 0.04025
R35393 VDD.n3131 VDD.n2912 0.04025
R35394 VDD.n3127 VDD.n2912 0.04025
R35395 VDD.n3127 VDD.n3126 0.04025
R35396 VDD.n3126 VDD.n3125 0.04025
R35397 VDD.n3125 VDD.n2914 0.04025
R35398 VDD.n3121 VDD.n2914 0.04025
R35399 VDD.n3121 VDD.n3120 0.04025
R35400 VDD.n3120 VDD.n3119 0.04025
R35401 VDD.n3119 VDD.n2916 0.04025
R35402 VDD.n3115 VDD.n2916 0.04025
R35403 VDD.n3115 VDD.n3114 0.04025
R35404 VDD.n3114 VDD.n3113 0.04025
R35405 VDD.n3113 VDD.n2918 0.04025
R35406 VDD.n3109 VDD.n2918 0.04025
R35407 VDD.n3109 VDD.n3108 0.04025
R35408 VDD.n3108 VDD.n3107 0.04025
R35409 VDD.n3107 VDD.n2920 0.04025
R35410 VDD.n3103 VDD.n2920 0.04025
R35411 VDD.n3103 VDD.n3102 0.04025
R35412 VDD.n3102 VDD.n3101 0.04025
R35413 VDD.n3101 VDD.n2922 0.04025
R35414 VDD.n3097 VDD.n2922 0.04025
R35415 VDD.n3097 VDD.n3096 0.04025
R35416 VDD.n3096 VDD.n3095 0.04025
R35417 VDD.n3095 VDD.n2924 0.04025
R35418 VDD.n3091 VDD.n2924 0.04025
R35419 VDD.n3091 VDD.n3090 0.04025
R35420 VDD.n3090 VDD.n3089 0.04025
R35421 VDD.n3089 VDD.n2926 0.04025
R35422 VDD.n3085 VDD.n2926 0.04025
R35423 VDD.n3085 VDD.n3084 0.04025
R35424 VDD.n3084 VDD.n3083 0.04025
R35425 VDD.n3083 VDD.n2928 0.04025
R35426 VDD.n3079 VDD.n2928 0.04025
R35427 VDD.n3079 VDD.n3078 0.04025
R35428 VDD.n3078 VDD.n3077 0.04025
R35429 VDD.n3077 VDD.n2930 0.04025
R35430 VDD.n3073 VDD.n2930 0.04025
R35431 VDD.n3073 VDD.n3072 0.04025
R35432 VDD.n3072 VDD.n3071 0.04025
R35433 VDD.n3071 VDD.n2932 0.04025
R35434 VDD.n3067 VDD.n2932 0.04025
R35435 VDD.n3067 VDD.n3066 0.04025
R35436 VDD.n3066 VDD.n3065 0.04025
R35437 VDD.n3065 VDD.n2934 0.04025
R35438 VDD.n3061 VDD.n2934 0.04025
R35439 VDD.n3061 VDD.n3060 0.04025
R35440 VDD.n3060 VDD.n3059 0.04025
R35441 VDD.n3059 VDD.n2936 0.04025
R35442 VDD.n3055 VDD.n2936 0.04025
R35443 VDD.n3055 VDD.n3054 0.04025
R35444 VDD.n3054 VDD.n3053 0.04025
R35445 VDD.n3053 VDD.n2938 0.04025
R35446 VDD.n3049 VDD.n2938 0.04025
R35447 VDD.n3049 VDD.n3048 0.04025
R35448 VDD.n3048 VDD.n3047 0.04025
R35449 VDD.n3047 VDD.n2940 0.04025
R35450 VDD.n3043 VDD.n2940 0.04025
R35451 VDD.n3043 VDD.n3042 0.04025
R35452 VDD.n3042 VDD.n3041 0.04025
R35453 VDD.n3041 VDD.n2942 0.04025
R35454 VDD.n3037 VDD.n2942 0.04025
R35455 VDD.n3037 VDD.n3036 0.04025
R35456 VDD.n3036 VDD.n3035 0.04025
R35457 VDD.n3035 VDD.n2944 0.04025
R35458 VDD.n3031 VDD.n2944 0.04025
R35459 VDD.n3031 VDD.n3030 0.04025
R35460 VDD.n3030 VDD.n3029 0.04025
R35461 VDD.n3029 VDD.n2946 0.04025
R35462 VDD.n3025 VDD.n2946 0.04025
R35463 VDD.n3025 VDD.n3024 0.04025
R35464 VDD.n3024 VDD.n3023 0.04025
R35465 VDD.n3023 VDD.n2948 0.04025
R35466 VDD.n3019 VDD.n2948 0.04025
R35467 VDD.n3019 VDD.n3018 0.04025
R35468 VDD.n3018 VDD.n3017 0.04025
R35469 VDD.n3017 VDD.n2950 0.04025
R35470 VDD.n3013 VDD.n2950 0.04025
R35471 VDD.n3013 VDD.n3012 0.04025
R35472 VDD.n3012 VDD.n3011 0.04025
R35473 VDD.n3011 VDD.n2952 0.04025
R35474 VDD.n3007 VDD.n2952 0.04025
R35475 VDD.n3007 VDD.n3006 0.04025
R35476 VDD.n3006 VDD.n3005 0.04025
R35477 VDD.n3005 VDD.n2954 0.04025
R35478 VDD.n3001 VDD.n2954 0.04025
R35479 VDD.n3001 VDD.n3000 0.04025
R35480 VDD.n3000 VDD.n2999 0.04025
R35481 VDD.n2999 VDD.n2956 0.04025
R35482 VDD.n2995 VDD.n2956 0.04025
R35483 VDD.n2995 VDD.n2994 0.04025
R35484 VDD.n2994 VDD.n2993 0.04025
R35485 VDD.n2993 VDD.n2958 0.04025
R35486 VDD.n2989 VDD.n2958 0.04025
R35487 VDD.n2989 VDD.n2988 0.04025
R35488 VDD.n2988 VDD.n2987 0.04025
R35489 VDD.n2987 VDD.n2960 0.04025
R35490 VDD.n2983 VDD.n2960 0.04025
R35491 VDD.n2983 VDD.n2982 0.04025
R35492 VDD.n2982 VDD.n2981 0.04025
R35493 VDD.n2981 VDD.n2962 0.04025
R35494 VDD.n2977 VDD.n2962 0.04025
R35495 VDD.n2977 VDD.n2976 0.04025
R35496 VDD.n2976 VDD.n2975 0.04025
R35497 VDD.n2975 VDD.n2964 0.04025
R35498 VDD.n2971 VDD.n2964 0.04025
R35499 VDD.n2971 VDD.n2970 0.04025
R35500 VDD.n3631 VDD.n3630 0.04025
R35501 VDD.n3631 VDD.n2744 0.04025
R35502 VDD.n3635 VDD.n2744 0.04025
R35503 VDD.n3636 VDD.n3635 0.04025
R35504 VDD.n3637 VDD.n3636 0.04025
R35505 VDD.n3637 VDD.n2742 0.04025
R35506 VDD.n3641 VDD.n2742 0.04025
R35507 VDD.n3642 VDD.n3641 0.04025
R35508 VDD.n3643 VDD.n3642 0.04025
R35509 VDD.n3643 VDD.n2740 0.04025
R35510 VDD.n3647 VDD.n2740 0.04025
R35511 VDD.n3648 VDD.n3647 0.04025
R35512 VDD.n3649 VDD.n3648 0.04025
R35513 VDD.n3649 VDD.n2738 0.04025
R35514 VDD.n3653 VDD.n2738 0.04025
R35515 VDD.n3654 VDD.n3653 0.04025
R35516 VDD.n3655 VDD.n3654 0.04025
R35517 VDD.n3655 VDD.n2736 0.04025
R35518 VDD.n3659 VDD.n2736 0.04025
R35519 VDD.n3660 VDD.n3659 0.04025
R35520 VDD.n3661 VDD.n3660 0.04025
R35521 VDD.n3661 VDD.n2734 0.04025
R35522 VDD.n3665 VDD.n2734 0.04025
R35523 VDD.n3666 VDD.n3665 0.04025
R35524 VDD.n3667 VDD.n3666 0.04025
R35525 VDD.n3667 VDD.n2732 0.04025
R35526 VDD.n3671 VDD.n2732 0.04025
R35527 VDD.n3672 VDD.n3671 0.04025
R35528 VDD.n3673 VDD.n3672 0.04025
R35529 VDD.n3673 VDD.n2730 0.04025
R35530 VDD.n3677 VDD.n2730 0.04025
R35531 VDD.n3678 VDD.n3677 0.04025
R35532 VDD.n3679 VDD.n3678 0.04025
R35533 VDD.n3679 VDD.n2728 0.04025
R35534 VDD.n3683 VDD.n2728 0.04025
R35535 VDD.n3684 VDD.n3683 0.04025
R35536 VDD.n3685 VDD.n3684 0.04025
R35537 VDD.n3685 VDD.n2726 0.04025
R35538 VDD.n3689 VDD.n2726 0.04025
R35539 VDD.n3690 VDD.n3689 0.04025
R35540 VDD.n3691 VDD.n3690 0.04025
R35541 VDD.n3691 VDD.n2724 0.04025
R35542 VDD.n3695 VDD.n2724 0.04025
R35543 VDD.n3696 VDD.n3695 0.04025
R35544 VDD.n3697 VDD.n3696 0.04025
R35545 VDD.n3697 VDD.n2722 0.04025
R35546 VDD.n3701 VDD.n2722 0.04025
R35547 VDD.n3702 VDD.n3701 0.04025
R35548 VDD.n3703 VDD.n3702 0.04025
R35549 VDD.n3703 VDD.n2720 0.04025
R35550 VDD.n3707 VDD.n2720 0.04025
R35551 VDD.n3708 VDD.n3707 0.04025
R35552 VDD.n3709 VDD.n3708 0.04025
R35553 VDD.n3709 VDD.n2718 0.04025
R35554 VDD.n3713 VDD.n2718 0.04025
R35555 VDD.n3714 VDD.n3713 0.04025
R35556 VDD.n3715 VDD.n3714 0.04025
R35557 VDD.n3715 VDD.n2716 0.04025
R35558 VDD.n3719 VDD.n2716 0.04025
R35559 VDD.n3720 VDD.n3719 0.04025
R35560 VDD.n3721 VDD.n3720 0.04025
R35561 VDD.n3721 VDD.n2714 0.04025
R35562 VDD.n3725 VDD.n2714 0.04025
R35563 VDD.n3726 VDD.n3725 0.04025
R35564 VDD.n3727 VDD.n3726 0.04025
R35565 VDD.n3727 VDD.n2712 0.04025
R35566 VDD.n3731 VDD.n2712 0.04025
R35567 VDD.n3732 VDD.n3731 0.04025
R35568 VDD.n3733 VDD.n3732 0.04025
R35569 VDD.n3733 VDD.n2710 0.04025
R35570 VDD.n3737 VDD.n2710 0.04025
R35571 VDD.n3738 VDD.n3737 0.04025
R35572 VDD.n3739 VDD.n3738 0.04025
R35573 VDD.n3739 VDD.n2708 0.04025
R35574 VDD.n3743 VDD.n2708 0.04025
R35575 VDD.n3744 VDD.n3743 0.04025
R35576 VDD.n3745 VDD.n3744 0.04025
R35577 VDD.n3745 VDD.n2706 0.04025
R35578 VDD.n3749 VDD.n2706 0.04025
R35579 VDD.n3750 VDD.n3749 0.04025
R35580 VDD.n3751 VDD.n3750 0.04025
R35581 VDD.n3751 VDD.n2704 0.04025
R35582 VDD.n3755 VDD.n2704 0.04025
R35583 VDD.n3756 VDD.n3755 0.04025
R35584 VDD.n3757 VDD.n3756 0.04025
R35585 VDD.n3757 VDD.n2702 0.04025
R35586 VDD.n3761 VDD.n2702 0.04025
R35587 VDD.n3762 VDD.n3761 0.04025
R35588 VDD.n3763 VDD.n3762 0.04025
R35589 VDD.n3763 VDD.n2700 0.04025
R35590 VDD.n3767 VDD.n2700 0.04025
R35591 VDD.n3768 VDD.n3767 0.04025
R35592 VDD.n3769 VDD.n3768 0.04025
R35593 VDD.n3769 VDD.n2698 0.04025
R35594 VDD.n3773 VDD.n2698 0.04025
R35595 VDD.n3774 VDD.n3773 0.04025
R35596 VDD.n3775 VDD.n3774 0.04025
R35597 VDD.n3775 VDD.n2696 0.04025
R35598 VDD.n3779 VDD.n2696 0.04025
R35599 VDD.n3780 VDD.n3779 0.04025
R35600 VDD.n3781 VDD.n3780 0.04025
R35601 VDD.n3781 VDD.n2694 0.04025
R35602 VDD.n3785 VDD.n2694 0.04025
R35603 VDD.n3786 VDD.n3785 0.04025
R35604 VDD.n3787 VDD.n3786 0.04025
R35605 VDD.n3787 VDD.n2692 0.04025
R35606 VDD.n3791 VDD.n2692 0.04025
R35607 VDD.n3792 VDD.n3791 0.04025
R35608 VDD.n3793 VDD.n3792 0.04025
R35609 VDD.n3793 VDD.n2690 0.04025
R35610 VDD.n3797 VDD.n2690 0.04025
R35611 VDD.n3798 VDD.n3797 0.04025
R35612 VDD.n3799 VDD.n3798 0.04025
R35613 VDD.n3799 VDD.n2688 0.04025
R35614 VDD.n3803 VDD.n2688 0.04025
R35615 VDD.n3804 VDD.n3803 0.04025
R35616 VDD.n3805 VDD.n3804 0.04025
R35617 VDD.n3805 VDD.n2686 0.04025
R35618 VDD.n3809 VDD.n2686 0.04025
R35619 VDD.n3810 VDD.n3809 0.04025
R35620 VDD.n3811 VDD.n3810 0.04025
R35621 VDD.n3811 VDD.n2684 0.04025
R35622 VDD.n3815 VDD.n2684 0.04025
R35623 VDD.n3816 VDD.n3815 0.04025
R35624 VDD.n3817 VDD.n3816 0.04025
R35625 VDD.n3817 VDD.n2682 0.04025
R35626 VDD.n3821 VDD.n2682 0.04025
R35627 VDD.n3822 VDD.n3821 0.04025
R35628 VDD.n3823 VDD.n3822 0.04025
R35629 VDD.n3823 VDD.n2680 0.04025
R35630 VDD.n3827 VDD.n2680 0.04025
R35631 VDD.n3828 VDD.n3827 0.04025
R35632 VDD.n3829 VDD.n3828 0.04025
R35633 VDD.n3829 VDD.n2678 0.04025
R35634 VDD.n3833 VDD.n2678 0.04025
R35635 VDD.n3834 VDD.n3833 0.04025
R35636 VDD.n3835 VDD.n3834 0.04025
R35637 VDD.n3835 VDD.n2676 0.04025
R35638 VDD.n3839 VDD.n2676 0.04025
R35639 VDD.n3840 VDD.n3839 0.04025
R35640 VDD.n3841 VDD.n3840 0.04025
R35641 VDD.n3841 VDD.n2674 0.04025
R35642 VDD.n3845 VDD.n2674 0.04025
R35643 VDD.n3846 VDD.n3845 0.04025
R35644 VDD.n3847 VDD.n3846 0.04025
R35645 VDD.n3847 VDD.n2672 0.04025
R35646 VDD.n3851 VDD.n2672 0.04025
R35647 VDD.n3852 VDD.n3851 0.04025
R35648 VDD.n3853 VDD.n3852 0.04025
R35649 VDD.n3853 VDD.n2670 0.04025
R35650 VDD.n3857 VDD.n2670 0.04025
R35651 VDD.n3858 VDD.n3857 0.04025
R35652 VDD.n3859 VDD.n3858 0.04025
R35653 VDD.n3859 VDD.n2668 0.04025
R35654 VDD.n3863 VDD.n2668 0.04025
R35655 VDD.n3864 VDD.n3863 0.04025
R35656 VDD.n3865 VDD.n3864 0.04025
R35657 VDD.n3865 VDD.n2666 0.04025
R35658 VDD.n3869 VDD.n2666 0.04025
R35659 VDD.n3870 VDD.n3869 0.04025
R35660 VDD.n3871 VDD.n3870 0.04025
R35661 VDD.n3871 VDD.n2664 0.04025
R35662 VDD.n3875 VDD.n2664 0.04025
R35663 VDD.n3876 VDD.n3875 0.04025
R35664 VDD.n3877 VDD.n3876 0.04025
R35665 VDD.n3877 VDD.n2662 0.04025
R35666 VDD.n3881 VDD.n2662 0.04025
R35667 VDD.n3882 VDD.n3881 0.04025
R35668 VDD.n3883 VDD.n3882 0.04025
R35669 VDD.n3883 VDD.n2660 0.04025
R35670 VDD.n3887 VDD.n2660 0.04025
R35671 VDD.n3888 VDD.n3887 0.04025
R35672 VDD.n3889 VDD.n3888 0.04025
R35673 VDD.n3889 VDD.n2658 0.04025
R35674 VDD.n3893 VDD.n2658 0.04025
R35675 VDD.n3894 VDD.n3893 0.04025
R35676 VDD.n3895 VDD.n3894 0.04025
R35677 VDD.n3895 VDD.n2656 0.04025
R35678 VDD.n3899 VDD.n2656 0.04025
R35679 VDD.n3900 VDD.n3899 0.04025
R35680 VDD.n3901 VDD.n3900 0.04025
R35681 VDD.n3901 VDD.n2654 0.04025
R35682 VDD.n3905 VDD.n2654 0.04025
R35683 VDD.n3906 VDD.n3905 0.04025
R35684 VDD.n3907 VDD.n3906 0.04025
R35685 VDD.n3907 VDD.n2652 0.04025
R35686 VDD.n3911 VDD.n2652 0.04025
R35687 VDD.n3912 VDD.n3911 0.04025
R35688 VDD.n3913 VDD.n3912 0.04025
R35689 VDD.n3913 VDD.n2650 0.04025
R35690 VDD.n3917 VDD.n2650 0.04025
R35691 VDD.n3918 VDD.n3917 0.04025
R35692 VDD.n3919 VDD.n3918 0.04025
R35693 VDD.n3919 VDD.n2648 0.04025
R35694 VDD.n3923 VDD.n2648 0.04025
R35695 VDD.n3924 VDD.n3923 0.04025
R35696 VDD.n3925 VDD.n3924 0.04025
R35697 VDD.n3925 VDD.n2646 0.04025
R35698 VDD.n3929 VDD.n2646 0.04025
R35699 VDD.n3930 VDD.n3929 0.04025
R35700 VDD.n3931 VDD.n3930 0.04025
R35701 VDD.n3931 VDD.n2644 0.04025
R35702 VDD.n3935 VDD.n2644 0.04025
R35703 VDD.n3936 VDD.n3935 0.04025
R35704 VDD.n3937 VDD.n3936 0.04025
R35705 VDD.n3937 VDD.n2642 0.04025
R35706 VDD.n3941 VDD.n2642 0.04025
R35707 VDD.n3942 VDD.n3941 0.04025
R35708 VDD.n3943 VDD.n3942 0.04025
R35709 VDD.n3943 VDD.n2640 0.04025
R35710 VDD.n3947 VDD.n2640 0.04025
R35711 VDD.n3948 VDD.n3947 0.04025
R35712 VDD.n3949 VDD.n3948 0.04025
R35713 VDD.n3949 VDD.n2638 0.04025
R35714 VDD.n3953 VDD.n2638 0.04025
R35715 VDD.n3954 VDD.n3953 0.04025
R35716 VDD.n3955 VDD.n3954 0.04025
R35717 VDD.n3955 VDD.n2636 0.04025
R35718 VDD.n3959 VDD.n2636 0.04025
R35719 VDD.n3960 VDD.n3959 0.04025
R35720 VDD.n3961 VDD.n3960 0.04025
R35721 VDD.n3961 VDD.n2634 0.04025
R35722 VDD.n3965 VDD.n2634 0.04025
R35723 VDD.n3966 VDD.n3965 0.04025
R35724 VDD.n3967 VDD.n3966 0.04025
R35725 VDD.n3967 VDD.n2632 0.04025
R35726 VDD.n3971 VDD.n2632 0.04025
R35727 VDD.n3972 VDD.n3971 0.04025
R35728 VDD.n3973 VDD.n3972 0.04025
R35729 VDD.n3973 VDD.n2630 0.04025
R35730 VDD.n3977 VDD.n2630 0.04025
R35731 VDD.n3978 VDD.n3977 0.04025
R35732 VDD.n3979 VDD.n3978 0.04025
R35733 VDD.n3979 VDD.n2628 0.04025
R35734 VDD.n3983 VDD.n2628 0.04025
R35735 VDD.n3984 VDD.n3983 0.04025
R35736 VDD.n3985 VDD.n3984 0.04025
R35737 VDD.n3985 VDD.n2626 0.04025
R35738 VDD.n3989 VDD.n2626 0.04025
R35739 VDD.n3990 VDD.n3989 0.04025
R35740 VDD.n3991 VDD.n3990 0.04025
R35741 VDD.n3991 VDD.n2624 0.04025
R35742 VDD.n3995 VDD.n2624 0.04025
R35743 VDD.n3996 VDD.n3995 0.04025
R35744 VDD.n3997 VDD.n3996 0.04025
R35745 VDD.n3997 VDD.n2622 0.04025
R35746 VDD.n4001 VDD.n2622 0.04025
R35747 VDD.n4002 VDD.n4001 0.04025
R35748 VDD.n4003 VDD.n4002 0.04025
R35749 VDD.n4003 VDD.n2620 0.04025
R35750 VDD.n4007 VDD.n2620 0.04025
R35751 VDD.n4008 VDD.n4007 0.04025
R35752 VDD.n4009 VDD.n4008 0.04025
R35753 VDD.n4009 VDD.n2618 0.04025
R35754 VDD.n4013 VDD.n2618 0.04025
R35755 VDD.n4014 VDD.n4013 0.04025
R35756 VDD.n4015 VDD.n4014 0.04025
R35757 VDD.n4015 VDD.n2616 0.04025
R35758 VDD.n4019 VDD.n2616 0.04025
R35759 VDD.n4020 VDD.n4019 0.04025
R35760 VDD.n4021 VDD.n4020 0.04025
R35761 VDD.n4021 VDD.n2614 0.04025
R35762 VDD.n4025 VDD.n2614 0.04025
R35763 VDD.n4026 VDD.n4025 0.04025
R35764 VDD.n4027 VDD.n4026 0.04025
R35765 VDD.n4027 VDD.n2612 0.04025
R35766 VDD.n4031 VDD.n2612 0.04025
R35767 VDD.n4032 VDD.n4031 0.04025
R35768 VDD.n4033 VDD.n4032 0.04025
R35769 VDD.n4033 VDD.n2610 0.04025
R35770 VDD.n4037 VDD.n2610 0.04025
R35771 VDD.n4038 VDD.n4037 0.04025
R35772 VDD.n4039 VDD.n4038 0.04025
R35773 VDD.n4039 VDD.n2608 0.04025
R35774 VDD.n4043 VDD.n2608 0.04025
R35775 VDD.n4044 VDD.n4043 0.04025
R35776 VDD.n4045 VDD.n4044 0.04025
R35777 VDD.n4045 VDD.n2606 0.04025
R35778 VDD.n4049 VDD.n2606 0.04025
R35779 VDD.n4050 VDD.n4049 0.04025
R35780 VDD.n4051 VDD.n4050 0.04025
R35781 VDD.n4051 VDD.n2604 0.04025
R35782 VDD.n4055 VDD.n2604 0.04025
R35783 VDD.n4056 VDD.n4055 0.04025
R35784 VDD.n4057 VDD.n4056 0.04025
R35785 VDD.n4057 VDD.n2602 0.04025
R35786 VDD.n4061 VDD.n2602 0.04025
R35787 VDD.n4062 VDD.n4061 0.04025
R35788 VDD.n4063 VDD.n4062 0.04025
R35789 VDD.n4063 VDD.n2600 0.04025
R35790 VDD.n4067 VDD.n2600 0.04025
R35791 VDD.n4068 VDD.n4067 0.04025
R35792 VDD.n4069 VDD.n4068 0.04025
R35793 VDD.n4069 VDD.n2598 0.04025
R35794 VDD.n4073 VDD.n2598 0.04025
R35795 VDD.n4074 VDD.n4073 0.04025
R35796 VDD.n4075 VDD.n4074 0.04025
R35797 VDD.n4075 VDD.n2596 0.04025
R35798 VDD.n4079 VDD.n2596 0.04025
R35799 VDD.n4080 VDD.n4079 0.04025
R35800 VDD.n4081 VDD.n4080 0.04025
R35801 VDD.n4081 VDD.n2594 0.04025
R35802 VDD.n4085 VDD.n2594 0.04025
R35803 VDD.n4086 VDD.n4085 0.04025
R35804 VDD.n4087 VDD.n4086 0.04025
R35805 VDD.n4087 VDD.n2592 0.04025
R35806 VDD.n4091 VDD.n2592 0.04025
R35807 VDD.n4092 VDD.n4091 0.04025
R35808 VDD.n4093 VDD.n4092 0.04025
R35809 VDD.n4093 VDD.n2590 0.04025
R35810 VDD.n4097 VDD.n2590 0.04025
R35811 VDD.n4098 VDD.n4097 0.04025
R35812 VDD.n4099 VDD.n4098 0.04025
R35813 VDD.n4099 VDD.n2588 0.04025
R35814 VDD.n4103 VDD.n2588 0.04025
R35815 VDD.n4104 VDD.n4103 0.04025
R35816 VDD.n4105 VDD.n4104 0.04025
R35817 VDD.n4105 VDD.n2586 0.04025
R35818 VDD.n4109 VDD.n2586 0.04025
R35819 VDD.n4110 VDD.n4109 0.04025
R35820 VDD.n4111 VDD.n4110 0.04025
R35821 VDD.n4111 VDD.n2584 0.04025
R35822 VDD.n4115 VDD.n2584 0.04025
R35823 VDD.n4116 VDD.n4115 0.04025
R35824 VDD.n4117 VDD.n4116 0.04025
R35825 VDD.n4117 VDD.n2582 0.04025
R35826 VDD.n4121 VDD.n2582 0.04025
R35827 VDD.n4122 VDD.n4121 0.04025
R35828 VDD.n4123 VDD.n4122 0.04025
R35829 VDD.n4123 VDD.n2580 0.04025
R35830 VDD.n4127 VDD.n2580 0.04025
R35831 VDD.n4128 VDD.n4127 0.04025
R35832 VDD.n4129 VDD.n4128 0.04025
R35833 VDD.n4129 VDD.n2578 0.04025
R35834 VDD.n4133 VDD.n2578 0.04025
R35835 VDD.n4134 VDD.n4133 0.04025
R35836 VDD.n4135 VDD.n4134 0.04025
R35837 VDD.n4135 VDD.n2576 0.04025
R35838 VDD.n4139 VDD.n2576 0.04025
R35839 VDD.n4140 VDD.n4139 0.04025
R35840 VDD.n4141 VDD.n4140 0.04025
R35841 VDD.n4141 VDD.n2574 0.04025
R35842 VDD.n4145 VDD.n2574 0.04025
R35843 VDD.n4146 VDD.n4145 0.04025
R35844 VDD.n4147 VDD.n4146 0.04025
R35845 VDD.n4147 VDD.n2572 0.04025
R35846 VDD.n4151 VDD.n2572 0.04025
R35847 VDD.n4152 VDD.n4151 0.04025
R35848 VDD.n4153 VDD.n4152 0.04025
R35849 VDD.n4153 VDD.n2570 0.04025
R35850 VDD.n4157 VDD.n2570 0.04025
R35851 VDD.n4158 VDD.n4157 0.04025
R35852 VDD.n4159 VDD.n4158 0.04025
R35853 VDD.n4159 VDD.n2568 0.04025
R35854 VDD.n4163 VDD.n2568 0.04025
R35855 VDD.n4164 VDD.n4163 0.04025
R35856 VDD.n4165 VDD.n4164 0.04025
R35857 VDD.n4165 VDD.n2566 0.04025
R35858 VDD.n4169 VDD.n2566 0.04025
R35859 VDD.n4170 VDD.n4169 0.04025
R35860 VDD.n4171 VDD.n4170 0.04025
R35861 VDD.n4171 VDD.n2564 0.04025
R35862 VDD.n4175 VDD.n2564 0.04025
R35863 VDD.n4176 VDD.n4175 0.04025
R35864 VDD.n4177 VDD.n4176 0.04025
R35865 VDD.n4177 VDD.n2562 0.04025
R35866 VDD.n4181 VDD.n2562 0.04025
R35867 VDD.n4182 VDD.n4181 0.04025
R35868 VDD.n4183 VDD.n4182 0.04025
R35869 VDD.n4183 VDD.n2560 0.04025
R35870 VDD.n4187 VDD.n2560 0.04025
R35871 VDD.n4188 VDD.n4187 0.04025
R35872 VDD.n4189 VDD.n4188 0.04025
R35873 VDD.n4189 VDD.n2558 0.04025
R35874 VDD.n4193 VDD.n2558 0.04025
R35875 VDD.n4194 VDD.n4193 0.04025
R35876 VDD.n4195 VDD.n4194 0.04025
R35877 VDD.n4195 VDD.n2556 0.04025
R35878 VDD.n4199 VDD.n2556 0.04025
R35879 VDD.n4200 VDD.n4199 0.04025
R35880 VDD.n4201 VDD.n4200 0.04025
R35881 VDD.n4201 VDD.n2554 0.04025
R35882 VDD.n4205 VDD.n2554 0.04025
R35883 VDD.n4206 VDD.n4205 0.04025
R35884 VDD.n4207 VDD.n4206 0.04025
R35885 VDD.n4207 VDD.n2552 0.04025
R35886 VDD.n4211 VDD.n2552 0.04025
R35887 VDD.n4212 VDD.n4211 0.04025
R35888 VDD.n4213 VDD.n4212 0.04025
R35889 VDD.n4213 VDD.n2550 0.04025
R35890 VDD.n4217 VDD.n2550 0.04025
R35891 VDD.n4218 VDD.n4217 0.04025
R35892 VDD.n4219 VDD.n4218 0.04025
R35893 VDD.n4219 VDD.n2548 0.04025
R35894 VDD.n4223 VDD.n2548 0.04025
R35895 VDD.n4224 VDD.n4223 0.04025
R35896 VDD.n4225 VDD.n4224 0.04025
R35897 VDD.n4225 VDD.n2546 0.04025
R35898 VDD.n4229 VDD.n2546 0.04025
R35899 VDD.n4230 VDD.n4229 0.04025
R35900 VDD.n4231 VDD.n4230 0.04025
R35901 VDD.n4231 VDD.n2544 0.04025
R35902 VDD.n4235 VDD.n2544 0.04025
R35903 VDD.n4236 VDD.n4235 0.04025
R35904 VDD.n4237 VDD.n4236 0.04025
R35905 VDD.n4237 VDD.n2542 0.04025
R35906 VDD.n4241 VDD.n2542 0.04025
R35907 VDD.n4242 VDD.n4241 0.04025
R35908 VDD.n4243 VDD.n4242 0.04025
R35909 VDD.n4243 VDD.n2540 0.04025
R35910 VDD.n4247 VDD.n2540 0.04025
R35911 VDD.n4248 VDD.n4247 0.04025
R35912 VDD.n4249 VDD.n4248 0.04025
R35913 VDD.n4249 VDD.n2538 0.04025
R35914 VDD.n4253 VDD.n2538 0.04025
R35915 VDD.n4254 VDD.n4253 0.04025
R35916 VDD.n4255 VDD.n4254 0.04025
R35917 VDD.n4255 VDD.n2536 0.04025
R35918 VDD.n4259 VDD.n2536 0.04025
R35919 VDD.n4260 VDD.n4259 0.04025
R35920 VDD.n4261 VDD.n4260 0.04025
R35921 VDD.n4261 VDD.n2534 0.04025
R35922 VDD.n4265 VDD.n2534 0.04025
R35923 VDD.n4266 VDD.n4265 0.04025
R35924 VDD.n4267 VDD.n4266 0.04025
R35925 VDD.n4267 VDD.n2532 0.04025
R35926 VDD.n4271 VDD.n2532 0.04025
R35927 VDD.n4272 VDD.n4271 0.04025
R35928 VDD.n4273 VDD.n4272 0.04025
R35929 VDD.n4273 VDD.n2530 0.04025
R35930 VDD.n4277 VDD.n2530 0.04025
R35931 VDD.n4278 VDD.n4277 0.04025
R35932 VDD.n4279 VDD.n4278 0.04025
R35933 VDD.n4279 VDD.n2528 0.04025
R35934 VDD.n4283 VDD.n2528 0.04025
R35935 VDD.n4284 VDD.n4283 0.04025
R35936 VDD.n4285 VDD.n4284 0.04025
R35937 VDD.n4285 VDD.n2526 0.04025
R35938 VDD.n4289 VDD.n2526 0.04025
R35939 VDD.n4290 VDD.n4289 0.04025
R35940 VDD.n4291 VDD.n4290 0.04025
R35941 VDD.n4291 VDD.n2524 0.04025
R35942 VDD.n4295 VDD.n2524 0.04025
R35943 VDD.n4296 VDD.n4295 0.04025
R35944 VDD.n4297 VDD.n4296 0.04025
R35945 VDD.n4297 VDD.n2522 0.04025
R35946 VDD.n4301 VDD.n2522 0.04025
R35947 VDD.n4302 VDD.n4301 0.04025
R35948 VDD.n4303 VDD.n4302 0.04025
R35949 VDD.n4303 VDD.n2520 0.04025
R35950 VDD.n4307 VDD.n2520 0.04025
R35951 VDD.n4308 VDD.n4307 0.04025
R35952 VDD.n4309 VDD.n4308 0.04025
R35953 VDD.n4309 VDD.n2518 0.04025
R35954 VDD.n4313 VDD.n2518 0.04025
R35955 VDD.n4314 VDD.n4313 0.04025
R35956 VDD.n4315 VDD.n4314 0.04025
R35957 VDD.n4315 VDD.n2516 0.04025
R35958 VDD.n4319 VDD.n2516 0.04025
R35959 VDD.n4320 VDD.n4319 0.04025
R35960 VDD.n4321 VDD.n4320 0.04025
R35961 VDD.n4321 VDD.n2514 0.04025
R35962 VDD.n4325 VDD.n2514 0.04025
R35963 VDD.n4326 VDD.n4325 0.04025
R35964 VDD.n4327 VDD.n4326 0.04025
R35965 VDD.n4327 VDD.n2512 0.04025
R35966 VDD.n4331 VDD.n2512 0.04025
R35967 VDD.n4332 VDD.n4331 0.04025
R35968 VDD.n4333 VDD.n4332 0.04025
R35969 VDD.n4333 VDD.n2510 0.04025
R35970 VDD.n4337 VDD.n2510 0.04025
R35971 VDD.n4338 VDD.n4337 0.04025
R35972 VDD.n4339 VDD.n4338 0.04025
R35973 VDD.n4339 VDD.n2508 0.04025
R35974 VDD.n4343 VDD.n2508 0.04025
R35975 VDD.n4344 VDD.n4343 0.04025
R35976 VDD.n4345 VDD.n4344 0.04025
R35977 VDD.n4345 VDD.n2506 0.04025
R35978 VDD.n4349 VDD.n2506 0.04025
R35979 VDD.n4350 VDD.n4349 0.04025
R35980 VDD.n4351 VDD.n4350 0.04025
R35981 VDD.n4351 VDD.n2504 0.04025
R35982 VDD.n4355 VDD.n2504 0.04025
R35983 VDD.n4356 VDD.n4355 0.04025
R35984 VDD.n4357 VDD.n4356 0.04025
R35985 VDD.n4357 VDD.n2502 0.04025
R35986 VDD.n4361 VDD.n2502 0.04025
R35987 VDD.n4362 VDD.n4361 0.04025
R35988 VDD.n4363 VDD.n4362 0.04025
R35989 VDD.n4363 VDD.n2500 0.04025
R35990 VDD.n4367 VDD.n2500 0.04025
R35991 VDD.n4368 VDD.n4367 0.04025
R35992 VDD.n4369 VDD.n4368 0.04025
R35993 VDD.n4369 VDD.n2498 0.04025
R35994 VDD.n4373 VDD.n2498 0.04025
R35995 VDD.n4374 VDD.n4373 0.04025
R35996 VDD.n4375 VDD.n4374 0.04025
R35997 VDD.n4375 VDD.n2496 0.04025
R35998 VDD.n4379 VDD.n2496 0.04025
R35999 VDD.n4380 VDD.n4379 0.04025
R36000 VDD.n4381 VDD.n4380 0.04025
R36001 VDD.n4381 VDD.n2494 0.04025
R36002 VDD.n4385 VDD.n2494 0.04025
R36003 VDD.n4386 VDD.n4385 0.04025
R36004 VDD.n4387 VDD.n4386 0.04025
R36005 VDD.n4387 VDD.n2492 0.04025
R36006 VDD.n4391 VDD.n2492 0.04025
R36007 VDD.n4392 VDD.n4391 0.04025
R36008 VDD.n4393 VDD.n4392 0.04025
R36009 VDD.n4393 VDD.n2490 0.04025
R36010 VDD.n4397 VDD.n2490 0.04025
R36011 VDD.n4398 VDD.n4397 0.04025
R36012 VDD.n4399 VDD.n4398 0.04025
R36013 VDD.n4399 VDD.n2488 0.04025
R36014 VDD.n4403 VDD.n2488 0.04025
R36015 VDD.n4404 VDD.n4403 0.04025
R36016 VDD.n4405 VDD.n4404 0.04025
R36017 VDD.n4405 VDD.n2486 0.04025
R36018 VDD.n4409 VDD.n2486 0.04025
R36019 VDD.n4410 VDD.n4409 0.04025
R36020 VDD.n4411 VDD.n4410 0.04025
R36021 VDD.n4411 VDD.n2484 0.04025
R36022 VDD.n4415 VDD.n2484 0.04025
R36023 VDD.n4416 VDD.n4415 0.04025
R36024 VDD.n4417 VDD.n4416 0.04025
R36025 VDD.n4417 VDD.n2482 0.04025
R36026 VDD.n4421 VDD.n2482 0.04025
R36027 VDD.n4422 VDD.n4421 0.04025
R36028 VDD.n4423 VDD.n4422 0.04025
R36029 VDD.n4423 VDD.n2480 0.04025
R36030 VDD.n4427 VDD.n2480 0.04025
R36031 VDD.n4428 VDD.n4427 0.04025
R36032 VDD.n4429 VDD.n4428 0.04025
R36033 VDD.n4429 VDD.n2478 0.04025
R36034 VDD.n4433 VDD.n2478 0.04025
R36035 VDD.n4434 VDD.n4433 0.04025
R36036 VDD.n4435 VDD.n4434 0.04025
R36037 VDD.n4435 VDD.n2476 0.04025
R36038 VDD.n4439 VDD.n2476 0.04025
R36039 VDD.n4440 VDD.n4439 0.04025
R36040 VDD.n4441 VDD.n4440 0.04025
R36041 VDD.n4441 VDD.n2474 0.04025
R36042 VDD.n4445 VDD.n2474 0.04025
R36043 VDD.n4446 VDD.n4445 0.04025
R36044 VDD.n4447 VDD.n4446 0.04025
R36045 VDD.n4447 VDD.n2472 0.04025
R36046 VDD.n4451 VDD.n2472 0.04025
R36047 VDD.n4452 VDD.n4451 0.04025
R36048 VDD.n4453 VDD.n4452 0.04025
R36049 VDD.n4453 VDD.n2470 0.04025
R36050 VDD.n4457 VDD.n2470 0.04025
R36051 VDD.n4458 VDD.n4457 0.04025
R36052 VDD.n4459 VDD.n4458 0.04025
R36053 VDD.n4459 VDD.n2468 0.04025
R36054 VDD.n4463 VDD.n2468 0.04025
R36055 VDD.n4464 VDD.n4463 0.04025
R36056 VDD.n4465 VDD.n4464 0.04025
R36057 VDD.n4465 VDD.n2466 0.04025
R36058 VDD.n4469 VDD.n2466 0.04025
R36059 VDD.n4470 VDD.n4469 0.04025
R36060 VDD.n4471 VDD.n4470 0.04025
R36061 VDD.n4471 VDD.n2464 0.04025
R36062 VDD.n4475 VDD.n2464 0.04025
R36063 VDD.n4476 VDD.n4475 0.04025
R36064 VDD.n4477 VDD.n4476 0.04025
R36065 VDD.n4477 VDD.n2462 0.04025
R36066 VDD.n4481 VDD.n2462 0.04025
R36067 VDD.n4482 VDD.n4481 0.04025
R36068 VDD.n4483 VDD.n4482 0.04025
R36069 VDD.n4483 VDD.n2460 0.04025
R36070 VDD.n4487 VDD.n2460 0.04025
R36071 VDD.n4488 VDD.n4487 0.04025
R36072 VDD.n4489 VDD.n4488 0.04025
R36073 VDD.n4489 VDD.n2458 0.04025
R36074 VDD.n4493 VDD.n2458 0.04025
R36075 VDD.n4494 VDD.n4493 0.04025
R36076 VDD.n4495 VDD.n4494 0.04025
R36077 VDD.n4495 VDD.n2456 0.04025
R36078 VDD.n4499 VDD.n2456 0.04025
R36079 VDD.n4500 VDD.n4499 0.04025
R36080 VDD.n4501 VDD.n4500 0.04025
R36081 VDD.n4501 VDD.n2454 0.04025
R36082 VDD.n4505 VDD.n2454 0.04025
R36083 VDD.n4506 VDD.n4505 0.04025
R36084 VDD.n4507 VDD.n4506 0.04025
R36085 VDD.n4507 VDD.n2452 0.04025
R36086 VDD.n4511 VDD.n2452 0.04025
R36087 VDD.n4512 VDD.n4511 0.04025
R36088 VDD.n4513 VDD.n4512 0.04025
R36089 VDD.n4513 VDD.n2450 0.04025
R36090 VDD.n4517 VDD.n2450 0.04025
R36091 VDD.n4518 VDD.n4517 0.04025
R36092 VDD.n4519 VDD.n4518 0.04025
R36093 VDD.n4519 VDD.n2448 0.04025
R36094 VDD.n4523 VDD.n2448 0.04025
R36095 VDD.n4524 VDD.n4523 0.04025
R36096 VDD.n4525 VDD.n4524 0.04025
R36097 VDD.n4525 VDD.n2446 0.04025
R36098 VDD.n4529 VDD.n2446 0.04025
R36099 VDD.n4530 VDD.n4529 0.04025
R36100 VDD.n4531 VDD.n4530 0.04025
R36101 VDD.n4531 VDD.n2444 0.04025
R36102 VDD.n4535 VDD.n2444 0.04025
R36103 VDD.n4536 VDD.n4535 0.04025
R36104 VDD.n4537 VDD.n4536 0.04025
R36105 VDD.n4537 VDD.n2442 0.04025
R36106 VDD.n4541 VDD.n2442 0.04025
R36107 VDD.n4542 VDD.n4541 0.04025
R36108 VDD.n4543 VDD.n4542 0.04025
R36109 VDD.n4543 VDD.n2440 0.04025
R36110 VDD.n4547 VDD.n2440 0.04025
R36111 VDD.n4548 VDD.n4547 0.04025
R36112 VDD.n4549 VDD.n4548 0.04025
R36113 VDD.n4549 VDD.n2438 0.04025
R36114 VDD.n4553 VDD.n2438 0.04025
R36115 VDD.n4554 VDD.n4553 0.04025
R36116 VDD.n4555 VDD.n4554 0.04025
R36117 VDD.n4555 VDD.n2436 0.04025
R36118 VDD.n4559 VDD.n2436 0.04025
R36119 VDD.n4560 VDD.n4559 0.04025
R36120 VDD.n4561 VDD.n4560 0.04025
R36121 VDD.n4561 VDD.n2434 0.04025
R36122 VDD.n4565 VDD.n2434 0.04025
R36123 VDD.n4566 VDD.n4565 0.04025
R36124 VDD.n4567 VDD.n4566 0.04025
R36125 VDD.n4567 VDD.n2432 0.04025
R36126 VDD.n4571 VDD.n2432 0.04025
R36127 VDD.n4572 VDD.n4571 0.04025
R36128 VDD.n4573 VDD.n4572 0.04025
R36129 VDD.n4573 VDD.n2430 0.04025
R36130 VDD.n4577 VDD.n2430 0.04025
R36131 VDD.n4578 VDD.n4577 0.04025
R36132 VDD.n4579 VDD.n4578 0.04025
R36133 VDD.n4579 VDD.n2428 0.04025
R36134 VDD.n4583 VDD.n2428 0.04025
R36135 VDD.n4584 VDD.n4583 0.04025
R36136 VDD.n4585 VDD.n4584 0.04025
R36137 VDD.n4585 VDD.n2426 0.04025
R36138 VDD.n4589 VDD.n2426 0.04025
R36139 VDD.n3632 VDD.n2745 0.04025
R36140 VDD.n3633 VDD.n3632 0.04025
R36141 VDD.n3634 VDD.n3633 0.04025
R36142 VDD.n3634 VDD.n2743 0.04025
R36143 VDD.n3638 VDD.n2743 0.04025
R36144 VDD.n3639 VDD.n3638 0.04025
R36145 VDD.n3640 VDD.n3639 0.04025
R36146 VDD.n3640 VDD.n2741 0.04025
R36147 VDD.n3644 VDD.n2741 0.04025
R36148 VDD.n3645 VDD.n3644 0.04025
R36149 VDD.n3646 VDD.n3645 0.04025
R36150 VDD.n3646 VDD.n2739 0.04025
R36151 VDD.n3650 VDD.n2739 0.04025
R36152 VDD.n3651 VDD.n3650 0.04025
R36153 VDD.n3652 VDD.n3651 0.04025
R36154 VDD.n3652 VDD.n2737 0.04025
R36155 VDD.n3656 VDD.n2737 0.04025
R36156 VDD.n3657 VDD.n3656 0.04025
R36157 VDD.n3658 VDD.n3657 0.04025
R36158 VDD.n3658 VDD.n2735 0.04025
R36159 VDD.n3662 VDD.n2735 0.04025
R36160 VDD.n3663 VDD.n3662 0.04025
R36161 VDD.n3664 VDD.n3663 0.04025
R36162 VDD.n3664 VDD.n2733 0.04025
R36163 VDD.n3668 VDD.n2733 0.04025
R36164 VDD.n3669 VDD.n3668 0.04025
R36165 VDD.n3670 VDD.n3669 0.04025
R36166 VDD.n3670 VDD.n2731 0.04025
R36167 VDD.n3674 VDD.n2731 0.04025
R36168 VDD.n3675 VDD.n3674 0.04025
R36169 VDD.n3676 VDD.n3675 0.04025
R36170 VDD.n3676 VDD.n2729 0.04025
R36171 VDD.n3680 VDD.n2729 0.04025
R36172 VDD.n3681 VDD.n3680 0.04025
R36173 VDD.n3682 VDD.n3681 0.04025
R36174 VDD.n3682 VDD.n2727 0.04025
R36175 VDD.n3686 VDD.n2727 0.04025
R36176 VDD.n3687 VDD.n3686 0.04025
R36177 VDD.n3688 VDD.n3687 0.04025
R36178 VDD.n3688 VDD.n2725 0.04025
R36179 VDD.n3692 VDD.n2725 0.04025
R36180 VDD.n3693 VDD.n3692 0.04025
R36181 VDD.n3694 VDD.n3693 0.04025
R36182 VDD.n3694 VDD.n2723 0.04025
R36183 VDD.n3698 VDD.n2723 0.04025
R36184 VDD.n3699 VDD.n3698 0.04025
R36185 VDD.n3700 VDD.n3699 0.04025
R36186 VDD.n3700 VDD.n2721 0.04025
R36187 VDD.n3704 VDD.n2721 0.04025
R36188 VDD.n3705 VDD.n3704 0.04025
R36189 VDD.n3706 VDD.n3705 0.04025
R36190 VDD.n3706 VDD.n2719 0.04025
R36191 VDD.n3710 VDD.n2719 0.04025
R36192 VDD.n3711 VDD.n3710 0.04025
R36193 VDD.n3712 VDD.n3711 0.04025
R36194 VDD.n3712 VDD.n2717 0.04025
R36195 VDD.n3716 VDD.n2717 0.04025
R36196 VDD.n3717 VDD.n3716 0.04025
R36197 VDD.n3718 VDD.n3717 0.04025
R36198 VDD.n3718 VDD.n2715 0.04025
R36199 VDD.n3722 VDD.n2715 0.04025
R36200 VDD.n3723 VDD.n3722 0.04025
R36201 VDD.n3724 VDD.n3723 0.04025
R36202 VDD.n3724 VDD.n2713 0.04025
R36203 VDD.n3728 VDD.n2713 0.04025
R36204 VDD.n3729 VDD.n3728 0.04025
R36205 VDD.n3730 VDD.n3729 0.04025
R36206 VDD.n3730 VDD.n2711 0.04025
R36207 VDD.n3734 VDD.n2711 0.04025
R36208 VDD.n3735 VDD.n3734 0.04025
R36209 VDD.n3736 VDD.n3735 0.04025
R36210 VDD.n3736 VDD.n2709 0.04025
R36211 VDD.n3740 VDD.n2709 0.04025
R36212 VDD.n3741 VDD.n3740 0.04025
R36213 VDD.n3742 VDD.n3741 0.04025
R36214 VDD.n3742 VDD.n2707 0.04025
R36215 VDD.n3746 VDD.n2707 0.04025
R36216 VDD.n3747 VDD.n3746 0.04025
R36217 VDD.n3748 VDD.n3747 0.04025
R36218 VDD.n3748 VDD.n2705 0.04025
R36219 VDD.n3752 VDD.n2705 0.04025
R36220 VDD.n3753 VDD.n3752 0.04025
R36221 VDD.n3754 VDD.n3753 0.04025
R36222 VDD.n3754 VDD.n2703 0.04025
R36223 VDD.n3758 VDD.n2703 0.04025
R36224 VDD.n3759 VDD.n3758 0.04025
R36225 VDD.n3760 VDD.n3759 0.04025
R36226 VDD.n3760 VDD.n2701 0.04025
R36227 VDD.n3764 VDD.n2701 0.04025
R36228 VDD.n3765 VDD.n3764 0.04025
R36229 VDD.n3766 VDD.n3765 0.04025
R36230 VDD.n3766 VDD.n2699 0.04025
R36231 VDD.n3770 VDD.n2699 0.04025
R36232 VDD.n3771 VDD.n3770 0.04025
R36233 VDD.n3772 VDD.n3771 0.04025
R36234 VDD.n3772 VDD.n2697 0.04025
R36235 VDD.n3776 VDD.n2697 0.04025
R36236 VDD.n3777 VDD.n3776 0.04025
R36237 VDD.n3778 VDD.n3777 0.04025
R36238 VDD.n3778 VDD.n2695 0.04025
R36239 VDD.n3782 VDD.n2695 0.04025
R36240 VDD.n3783 VDD.n3782 0.04025
R36241 VDD.n3784 VDD.n3783 0.04025
R36242 VDD.n3784 VDD.n2693 0.04025
R36243 VDD.n3788 VDD.n2693 0.04025
R36244 VDD.n3789 VDD.n3788 0.04025
R36245 VDD.n3790 VDD.n3789 0.04025
R36246 VDD.n3790 VDD.n2691 0.04025
R36247 VDD.n3794 VDD.n2691 0.04025
R36248 VDD.n3795 VDD.n3794 0.04025
R36249 VDD.n3796 VDD.n3795 0.04025
R36250 VDD.n3796 VDD.n2689 0.04025
R36251 VDD.n3800 VDD.n2689 0.04025
R36252 VDD.n3801 VDD.n3800 0.04025
R36253 VDD.n3802 VDD.n3801 0.04025
R36254 VDD.n3802 VDD.n2687 0.04025
R36255 VDD.n3806 VDD.n2687 0.04025
R36256 VDD.n3807 VDD.n3806 0.04025
R36257 VDD.n3808 VDD.n3807 0.04025
R36258 VDD.n3808 VDD.n2685 0.04025
R36259 VDD.n3812 VDD.n2685 0.04025
R36260 VDD.n3813 VDD.n3812 0.04025
R36261 VDD.n3814 VDD.n3813 0.04025
R36262 VDD.n3814 VDD.n2683 0.04025
R36263 VDD.n3818 VDD.n2683 0.04025
R36264 VDD.n3819 VDD.n3818 0.04025
R36265 VDD.n3820 VDD.n3819 0.04025
R36266 VDD.n3820 VDD.n2681 0.04025
R36267 VDD.n3824 VDD.n2681 0.04025
R36268 VDD.n3825 VDD.n3824 0.04025
R36269 VDD.n3826 VDD.n3825 0.04025
R36270 VDD.n3826 VDD.n2679 0.04025
R36271 VDD.n3830 VDD.n2679 0.04025
R36272 VDD.n3831 VDD.n3830 0.04025
R36273 VDD.n3832 VDD.n3831 0.04025
R36274 VDD.n3832 VDD.n2677 0.04025
R36275 VDD.n3836 VDD.n2677 0.04025
R36276 VDD.n3837 VDD.n3836 0.04025
R36277 VDD.n3838 VDD.n3837 0.04025
R36278 VDD.n3838 VDD.n2675 0.04025
R36279 VDD.n3842 VDD.n2675 0.04025
R36280 VDD.n3843 VDD.n3842 0.04025
R36281 VDD.n3844 VDD.n3843 0.04025
R36282 VDD.n3844 VDD.n2673 0.04025
R36283 VDD.n3848 VDD.n2673 0.04025
R36284 VDD.n3849 VDD.n3848 0.04025
R36285 VDD.n3850 VDD.n3849 0.04025
R36286 VDD.n3850 VDD.n2671 0.04025
R36287 VDD.n3854 VDD.n2671 0.04025
R36288 VDD.n3855 VDD.n3854 0.04025
R36289 VDD.n3856 VDD.n3855 0.04025
R36290 VDD.n3856 VDD.n2669 0.04025
R36291 VDD.n3860 VDD.n2669 0.04025
R36292 VDD.n3861 VDD.n3860 0.04025
R36293 VDD.n3862 VDD.n3861 0.04025
R36294 VDD.n3862 VDD.n2667 0.04025
R36295 VDD.n3866 VDD.n2667 0.04025
R36296 VDD.n3867 VDD.n3866 0.04025
R36297 VDD.n3868 VDD.n3867 0.04025
R36298 VDD.n3868 VDD.n2665 0.04025
R36299 VDD.n3872 VDD.n2665 0.04025
R36300 VDD.n3873 VDD.n3872 0.04025
R36301 VDD.n3874 VDD.n3873 0.04025
R36302 VDD.n3874 VDD.n2663 0.04025
R36303 VDD.n3878 VDD.n2663 0.04025
R36304 VDD.n3879 VDD.n3878 0.04025
R36305 VDD.n3880 VDD.n3879 0.04025
R36306 VDD.n3880 VDD.n2661 0.04025
R36307 VDD.n3884 VDD.n2661 0.04025
R36308 VDD.n3885 VDD.n3884 0.04025
R36309 VDD.n3886 VDD.n3885 0.04025
R36310 VDD.n3886 VDD.n2659 0.04025
R36311 VDD.n3890 VDD.n2659 0.04025
R36312 VDD.n3891 VDD.n3890 0.04025
R36313 VDD.n3892 VDD.n3891 0.04025
R36314 VDD.n3892 VDD.n2657 0.04025
R36315 VDD.n3896 VDD.n2657 0.04025
R36316 VDD.n3897 VDD.n3896 0.04025
R36317 VDD.n3898 VDD.n3897 0.04025
R36318 VDD.n3898 VDD.n2655 0.04025
R36319 VDD.n3902 VDD.n2655 0.04025
R36320 VDD.n3903 VDD.n3902 0.04025
R36321 VDD.n3904 VDD.n3903 0.04025
R36322 VDD.n3904 VDD.n2653 0.04025
R36323 VDD.n3908 VDD.n2653 0.04025
R36324 VDD.n3909 VDD.n3908 0.04025
R36325 VDD.n3910 VDD.n3909 0.04025
R36326 VDD.n3910 VDD.n2651 0.04025
R36327 VDD.n3914 VDD.n2651 0.04025
R36328 VDD.n3915 VDD.n3914 0.04025
R36329 VDD.n3916 VDD.n3915 0.04025
R36330 VDD.n3916 VDD.n2649 0.04025
R36331 VDD.n3920 VDD.n2649 0.04025
R36332 VDD.n3921 VDD.n3920 0.04025
R36333 VDD.n3922 VDD.n3921 0.04025
R36334 VDD.n3922 VDD.n2647 0.04025
R36335 VDD.n3926 VDD.n2647 0.04025
R36336 VDD.n3927 VDD.n3926 0.04025
R36337 VDD.n3928 VDD.n3927 0.04025
R36338 VDD.n3928 VDD.n2645 0.04025
R36339 VDD.n3932 VDD.n2645 0.04025
R36340 VDD.n3933 VDD.n3932 0.04025
R36341 VDD.n3934 VDD.n3933 0.04025
R36342 VDD.n3934 VDD.n2643 0.04025
R36343 VDD.n3938 VDD.n2643 0.04025
R36344 VDD.n3939 VDD.n3938 0.04025
R36345 VDD.n3940 VDD.n3939 0.04025
R36346 VDD.n3940 VDD.n2641 0.04025
R36347 VDD.n3944 VDD.n2641 0.04025
R36348 VDD.n3945 VDD.n3944 0.04025
R36349 VDD.n3946 VDD.n3945 0.04025
R36350 VDD.n3946 VDD.n2639 0.04025
R36351 VDD.n3950 VDD.n2639 0.04025
R36352 VDD.n3951 VDD.n3950 0.04025
R36353 VDD.n3952 VDD.n3951 0.04025
R36354 VDD.n3952 VDD.n2637 0.04025
R36355 VDD.n3956 VDD.n2637 0.04025
R36356 VDD.n3957 VDD.n3956 0.04025
R36357 VDD.n3958 VDD.n3957 0.04025
R36358 VDD.n3958 VDD.n2635 0.04025
R36359 VDD.n3962 VDD.n2635 0.04025
R36360 VDD.n3963 VDD.n3962 0.04025
R36361 VDD.n3964 VDD.n3963 0.04025
R36362 VDD.n3964 VDD.n2633 0.04025
R36363 VDD.n3968 VDD.n2633 0.04025
R36364 VDD.n3969 VDD.n3968 0.04025
R36365 VDD.n3970 VDD.n3969 0.04025
R36366 VDD.n3970 VDD.n2631 0.04025
R36367 VDD.n3974 VDD.n2631 0.04025
R36368 VDD.n3975 VDD.n3974 0.04025
R36369 VDD.n3976 VDD.n3975 0.04025
R36370 VDD.n3976 VDD.n2629 0.04025
R36371 VDD.n3980 VDD.n2629 0.04025
R36372 VDD.n3981 VDD.n3980 0.04025
R36373 VDD.n3982 VDD.n3981 0.04025
R36374 VDD.n3982 VDD.n2627 0.04025
R36375 VDD.n3986 VDD.n2627 0.04025
R36376 VDD.n3987 VDD.n3986 0.04025
R36377 VDD.n3988 VDD.n3987 0.04025
R36378 VDD.n3988 VDD.n2625 0.04025
R36379 VDD.n3992 VDD.n2625 0.04025
R36380 VDD.n3993 VDD.n3992 0.04025
R36381 VDD.n3994 VDD.n3993 0.04025
R36382 VDD.n3994 VDD.n2623 0.04025
R36383 VDD.n3998 VDD.n2623 0.04025
R36384 VDD.n3999 VDD.n3998 0.04025
R36385 VDD.n4000 VDD.n3999 0.04025
R36386 VDD.n4000 VDD.n2621 0.04025
R36387 VDD.n4004 VDD.n2621 0.04025
R36388 VDD.n4005 VDD.n4004 0.04025
R36389 VDD.n4006 VDD.n4005 0.04025
R36390 VDD.n4006 VDD.n2619 0.04025
R36391 VDD.n4010 VDD.n2619 0.04025
R36392 VDD.n4011 VDD.n4010 0.04025
R36393 VDD.n4012 VDD.n4011 0.04025
R36394 VDD.n4012 VDD.n2617 0.04025
R36395 VDD.n4016 VDD.n2617 0.04025
R36396 VDD.n4017 VDD.n4016 0.04025
R36397 VDD.n4018 VDD.n4017 0.04025
R36398 VDD.n4018 VDD.n2615 0.04025
R36399 VDD.n4022 VDD.n2615 0.04025
R36400 VDD.n4023 VDD.n4022 0.04025
R36401 VDD.n4024 VDD.n4023 0.04025
R36402 VDD.n4024 VDD.n2613 0.04025
R36403 VDD.n4028 VDD.n2613 0.04025
R36404 VDD.n4029 VDD.n4028 0.04025
R36405 VDD.n4030 VDD.n4029 0.04025
R36406 VDD.n4030 VDD.n2611 0.04025
R36407 VDD.n4034 VDD.n2611 0.04025
R36408 VDD.n4035 VDD.n4034 0.04025
R36409 VDD.n4036 VDD.n4035 0.04025
R36410 VDD.n4036 VDD.n2609 0.04025
R36411 VDD.n4040 VDD.n2609 0.04025
R36412 VDD.n4041 VDD.n4040 0.04025
R36413 VDD.n4042 VDD.n4041 0.04025
R36414 VDD.n4042 VDD.n2607 0.04025
R36415 VDD.n4046 VDD.n2607 0.04025
R36416 VDD.n4047 VDD.n4046 0.04025
R36417 VDD.n4048 VDD.n4047 0.04025
R36418 VDD.n4048 VDD.n2605 0.04025
R36419 VDD.n4052 VDD.n2605 0.04025
R36420 VDD.n4053 VDD.n4052 0.04025
R36421 VDD.n4054 VDD.n4053 0.04025
R36422 VDD.n4054 VDD.n2603 0.04025
R36423 VDD.n4058 VDD.n2603 0.04025
R36424 VDD.n4059 VDD.n4058 0.04025
R36425 VDD.n4060 VDD.n4059 0.04025
R36426 VDD.n4060 VDD.n2601 0.04025
R36427 VDD.n4064 VDD.n2601 0.04025
R36428 VDD.n4065 VDD.n4064 0.04025
R36429 VDD.n4066 VDD.n4065 0.04025
R36430 VDD.n4066 VDD.n2599 0.04025
R36431 VDD.n4070 VDD.n2599 0.04025
R36432 VDD.n4071 VDD.n4070 0.04025
R36433 VDD.n4072 VDD.n4071 0.04025
R36434 VDD.n4072 VDD.n2597 0.04025
R36435 VDD.n4076 VDD.n2597 0.04025
R36436 VDD.n4077 VDD.n4076 0.04025
R36437 VDD.n4078 VDD.n4077 0.04025
R36438 VDD.n4078 VDD.n2595 0.04025
R36439 VDD.n4082 VDD.n2595 0.04025
R36440 VDD.n4083 VDD.n4082 0.04025
R36441 VDD.n4084 VDD.n4083 0.04025
R36442 VDD.n4084 VDD.n2593 0.04025
R36443 VDD.n4088 VDD.n2593 0.04025
R36444 VDD.n4089 VDD.n4088 0.04025
R36445 VDD.n4090 VDD.n4089 0.04025
R36446 VDD.n4090 VDD.n2591 0.04025
R36447 VDD.n4094 VDD.n2591 0.04025
R36448 VDD.n4095 VDD.n4094 0.04025
R36449 VDD.n4096 VDD.n4095 0.04025
R36450 VDD.n4096 VDD.n2589 0.04025
R36451 VDD.n4100 VDD.n2589 0.04025
R36452 VDD.n4101 VDD.n4100 0.04025
R36453 VDD.n4102 VDD.n4101 0.04025
R36454 VDD.n4102 VDD.n2587 0.04025
R36455 VDD.n4106 VDD.n2587 0.04025
R36456 VDD.n4107 VDD.n4106 0.04025
R36457 VDD.n4108 VDD.n4107 0.04025
R36458 VDD.n4108 VDD.n2585 0.04025
R36459 VDD.n4112 VDD.n2585 0.04025
R36460 VDD.n4113 VDD.n4112 0.04025
R36461 VDD.n4114 VDD.n4113 0.04025
R36462 VDD.n4114 VDD.n2583 0.04025
R36463 VDD.n4118 VDD.n2583 0.04025
R36464 VDD.n4119 VDD.n4118 0.04025
R36465 VDD.n4120 VDD.n4119 0.04025
R36466 VDD.n4120 VDD.n2581 0.04025
R36467 VDD.n4124 VDD.n2581 0.04025
R36468 VDD.n4125 VDD.n4124 0.04025
R36469 VDD.n4126 VDD.n4125 0.04025
R36470 VDD.n4126 VDD.n2579 0.04025
R36471 VDD.n4130 VDD.n2579 0.04025
R36472 VDD.n4131 VDD.n4130 0.04025
R36473 VDD.n4132 VDD.n4131 0.04025
R36474 VDD.n4132 VDD.n2577 0.04025
R36475 VDD.n4136 VDD.n2577 0.04025
R36476 VDD.n4137 VDD.n4136 0.04025
R36477 VDD.n4138 VDD.n4137 0.04025
R36478 VDD.n4138 VDD.n2575 0.04025
R36479 VDD.n4142 VDD.n2575 0.04025
R36480 VDD.n4143 VDD.n4142 0.04025
R36481 VDD.n4144 VDD.n4143 0.04025
R36482 VDD.n4144 VDD.n2573 0.04025
R36483 VDD.n4148 VDD.n2573 0.04025
R36484 VDD.n4149 VDD.n4148 0.04025
R36485 VDD.n4150 VDD.n4149 0.04025
R36486 VDD.n4150 VDD.n2571 0.04025
R36487 VDD.n4154 VDD.n2571 0.04025
R36488 VDD.n4155 VDD.n4154 0.04025
R36489 VDD.n4156 VDD.n4155 0.04025
R36490 VDD.n4156 VDD.n2569 0.04025
R36491 VDD.n4160 VDD.n2569 0.04025
R36492 VDD.n4161 VDD.n4160 0.04025
R36493 VDD.n4162 VDD.n4161 0.04025
R36494 VDD.n4162 VDD.n2567 0.04025
R36495 VDD.n4166 VDD.n2567 0.04025
R36496 VDD.n4167 VDD.n4166 0.04025
R36497 VDD.n4168 VDD.n4167 0.04025
R36498 VDD.n4168 VDD.n2565 0.04025
R36499 VDD.n4172 VDD.n2565 0.04025
R36500 VDD.n4173 VDD.n4172 0.04025
R36501 VDD.n4174 VDD.n4173 0.04025
R36502 VDD.n4174 VDD.n2563 0.04025
R36503 VDD.n4178 VDD.n2563 0.04025
R36504 VDD.n4179 VDD.n4178 0.04025
R36505 VDD.n4180 VDD.n4179 0.04025
R36506 VDD.n4180 VDD.n2561 0.04025
R36507 VDD.n4184 VDD.n2561 0.04025
R36508 VDD.n4185 VDD.n4184 0.04025
R36509 VDD.n4186 VDD.n4185 0.04025
R36510 VDD.n4186 VDD.n2559 0.04025
R36511 VDD.n4190 VDD.n2559 0.04025
R36512 VDD.n4191 VDD.n4190 0.04025
R36513 VDD.n4192 VDD.n4191 0.04025
R36514 VDD.n4192 VDD.n2557 0.04025
R36515 VDD.n4196 VDD.n2557 0.04025
R36516 VDD.n4197 VDD.n4196 0.04025
R36517 VDD.n4198 VDD.n4197 0.04025
R36518 VDD.n4198 VDD.n2555 0.04025
R36519 VDD.n4202 VDD.n2555 0.04025
R36520 VDD.n4203 VDD.n4202 0.04025
R36521 VDD.n4204 VDD.n4203 0.04025
R36522 VDD.n4204 VDD.n2553 0.04025
R36523 VDD.n4208 VDD.n2553 0.04025
R36524 VDD.n4209 VDD.n4208 0.04025
R36525 VDD.n4210 VDD.n4209 0.04025
R36526 VDD.n4210 VDD.n2551 0.04025
R36527 VDD.n4214 VDD.n2551 0.04025
R36528 VDD.n4215 VDD.n4214 0.04025
R36529 VDD.n4216 VDD.n4215 0.04025
R36530 VDD.n4216 VDD.n2549 0.04025
R36531 VDD.n4220 VDD.n2549 0.04025
R36532 VDD.n4221 VDD.n4220 0.04025
R36533 VDD.n4222 VDD.n4221 0.04025
R36534 VDD.n4222 VDD.n2547 0.04025
R36535 VDD.n4226 VDD.n2547 0.04025
R36536 VDD.n4227 VDD.n4226 0.04025
R36537 VDD.n4228 VDD.n4227 0.04025
R36538 VDD.n4228 VDD.n2545 0.04025
R36539 VDD.n4232 VDD.n2545 0.04025
R36540 VDD.n4233 VDD.n4232 0.04025
R36541 VDD.n4234 VDD.n4233 0.04025
R36542 VDD.n4234 VDD.n2543 0.04025
R36543 VDD.n4238 VDD.n2543 0.04025
R36544 VDD.n4239 VDD.n4238 0.04025
R36545 VDD.n4240 VDD.n4239 0.04025
R36546 VDD.n4240 VDD.n2541 0.04025
R36547 VDD.n4244 VDD.n2541 0.04025
R36548 VDD.n4245 VDD.n4244 0.04025
R36549 VDD.n4246 VDD.n4245 0.04025
R36550 VDD.n4246 VDD.n2539 0.04025
R36551 VDD.n4250 VDD.n2539 0.04025
R36552 VDD.n4251 VDD.n4250 0.04025
R36553 VDD.n4252 VDD.n4251 0.04025
R36554 VDD.n4252 VDD.n2537 0.04025
R36555 VDD.n4256 VDD.n2537 0.04025
R36556 VDD.n4257 VDD.n4256 0.04025
R36557 VDD.n4258 VDD.n4257 0.04025
R36558 VDD.n4258 VDD.n2535 0.04025
R36559 VDD.n4262 VDD.n2535 0.04025
R36560 VDD.n4263 VDD.n4262 0.04025
R36561 VDD.n4264 VDD.n4263 0.04025
R36562 VDD.n4264 VDD.n2533 0.04025
R36563 VDD.n4268 VDD.n2533 0.04025
R36564 VDD.n4269 VDD.n4268 0.04025
R36565 VDD.n4270 VDD.n4269 0.04025
R36566 VDD.n4270 VDD.n2531 0.04025
R36567 VDD.n4274 VDD.n2531 0.04025
R36568 VDD.n4275 VDD.n4274 0.04025
R36569 VDD.n4276 VDD.n4275 0.04025
R36570 VDD.n4276 VDD.n2529 0.04025
R36571 VDD.n4280 VDD.n2529 0.04025
R36572 VDD.n4281 VDD.n4280 0.04025
R36573 VDD.n4282 VDD.n4281 0.04025
R36574 VDD.n4282 VDD.n2527 0.04025
R36575 VDD.n4286 VDD.n2527 0.04025
R36576 VDD.n4287 VDD.n4286 0.04025
R36577 VDD.n4288 VDD.n4287 0.04025
R36578 VDD.n4288 VDD.n2525 0.04025
R36579 VDD.n4292 VDD.n2525 0.04025
R36580 VDD.n4293 VDD.n4292 0.04025
R36581 VDD.n4294 VDD.n4293 0.04025
R36582 VDD.n4294 VDD.n2523 0.04025
R36583 VDD.n4298 VDD.n2523 0.04025
R36584 VDD.n4299 VDD.n4298 0.04025
R36585 VDD.n4300 VDD.n4299 0.04025
R36586 VDD.n4300 VDD.n2521 0.04025
R36587 VDD.n4304 VDD.n2521 0.04025
R36588 VDD.n4305 VDD.n4304 0.04025
R36589 VDD.n4306 VDD.n4305 0.04025
R36590 VDD.n4306 VDD.n2519 0.04025
R36591 VDD.n4310 VDD.n2519 0.04025
R36592 VDD.n4311 VDD.n4310 0.04025
R36593 VDD.n4312 VDD.n4311 0.04025
R36594 VDD.n4312 VDD.n2517 0.04025
R36595 VDD.n4316 VDD.n2517 0.04025
R36596 VDD.n4317 VDD.n4316 0.04025
R36597 VDD.n4318 VDD.n4317 0.04025
R36598 VDD.n4318 VDD.n2515 0.04025
R36599 VDD.n4322 VDD.n2515 0.04025
R36600 VDD.n4323 VDD.n4322 0.04025
R36601 VDD.n4324 VDD.n4323 0.04025
R36602 VDD.n4324 VDD.n2513 0.04025
R36603 VDD.n4328 VDD.n2513 0.04025
R36604 VDD.n4329 VDD.n4328 0.04025
R36605 VDD.n4330 VDD.n4329 0.04025
R36606 VDD.n4330 VDD.n2511 0.04025
R36607 VDD.n4334 VDD.n2511 0.04025
R36608 VDD.n4335 VDD.n4334 0.04025
R36609 VDD.n4336 VDD.n4335 0.04025
R36610 VDD.n4336 VDD.n2509 0.04025
R36611 VDD.n4340 VDD.n2509 0.04025
R36612 VDD.n4341 VDD.n4340 0.04025
R36613 VDD.n4342 VDD.n4341 0.04025
R36614 VDD.n4342 VDD.n2507 0.04025
R36615 VDD.n4346 VDD.n2507 0.04025
R36616 VDD.n4347 VDD.n4346 0.04025
R36617 VDD.n4348 VDD.n4347 0.04025
R36618 VDD.n4348 VDD.n2505 0.04025
R36619 VDD.n4352 VDD.n2505 0.04025
R36620 VDD.n4353 VDD.n4352 0.04025
R36621 VDD.n4354 VDD.n4353 0.04025
R36622 VDD.n4354 VDD.n2503 0.04025
R36623 VDD.n4358 VDD.n2503 0.04025
R36624 VDD.n4359 VDD.n4358 0.04025
R36625 VDD.n4360 VDD.n4359 0.04025
R36626 VDD.n4360 VDD.n2501 0.04025
R36627 VDD.n4364 VDD.n2501 0.04025
R36628 VDD.n4365 VDD.n4364 0.04025
R36629 VDD.n4366 VDD.n4365 0.04025
R36630 VDD.n4366 VDD.n2499 0.04025
R36631 VDD.n4370 VDD.n2499 0.04025
R36632 VDD.n4371 VDD.n4370 0.04025
R36633 VDD.n4372 VDD.n4371 0.04025
R36634 VDD.n4372 VDD.n2497 0.04025
R36635 VDD.n4376 VDD.n2497 0.04025
R36636 VDD.n4377 VDD.n4376 0.04025
R36637 VDD.n4378 VDD.n4377 0.04025
R36638 VDD.n4378 VDD.n2495 0.04025
R36639 VDD.n4382 VDD.n2495 0.04025
R36640 VDD.n4383 VDD.n4382 0.04025
R36641 VDD.n4384 VDD.n4383 0.04025
R36642 VDD.n4384 VDD.n2493 0.04025
R36643 VDD.n4388 VDD.n2493 0.04025
R36644 VDD.n4389 VDD.n4388 0.04025
R36645 VDD.n4390 VDD.n4389 0.04025
R36646 VDD.n4390 VDD.n2491 0.04025
R36647 VDD.n4394 VDD.n2491 0.04025
R36648 VDD.n4395 VDD.n4394 0.04025
R36649 VDD.n4396 VDD.n4395 0.04025
R36650 VDD.n4396 VDD.n2489 0.04025
R36651 VDD.n4400 VDD.n2489 0.04025
R36652 VDD.n4401 VDD.n4400 0.04025
R36653 VDD.n4402 VDD.n4401 0.04025
R36654 VDD.n4402 VDD.n2487 0.04025
R36655 VDD.n4406 VDD.n2487 0.04025
R36656 VDD.n4407 VDD.n4406 0.04025
R36657 VDD.n4408 VDD.n4407 0.04025
R36658 VDD.n4408 VDD.n2485 0.04025
R36659 VDD.n4412 VDD.n2485 0.04025
R36660 VDD.n4413 VDD.n4412 0.04025
R36661 VDD.n4414 VDD.n4413 0.04025
R36662 VDD.n4414 VDD.n2483 0.04025
R36663 VDD.n4418 VDD.n2483 0.04025
R36664 VDD.n4419 VDD.n4418 0.04025
R36665 VDD.n4420 VDD.n4419 0.04025
R36666 VDD.n4420 VDD.n2481 0.04025
R36667 VDD.n4424 VDD.n2481 0.04025
R36668 VDD.n4425 VDD.n4424 0.04025
R36669 VDD.n4426 VDD.n4425 0.04025
R36670 VDD.n4426 VDD.n2479 0.04025
R36671 VDD.n4430 VDD.n2479 0.04025
R36672 VDD.n4431 VDD.n4430 0.04025
R36673 VDD.n4432 VDD.n4431 0.04025
R36674 VDD.n4432 VDD.n2477 0.04025
R36675 VDD.n4436 VDD.n2477 0.04025
R36676 VDD.n4437 VDD.n4436 0.04025
R36677 VDD.n4438 VDD.n4437 0.04025
R36678 VDD.n4438 VDD.n2475 0.04025
R36679 VDD.n4442 VDD.n2475 0.04025
R36680 VDD.n4443 VDD.n4442 0.04025
R36681 VDD.n4444 VDD.n4443 0.04025
R36682 VDD.n4444 VDD.n2473 0.04025
R36683 VDD.n4448 VDD.n2473 0.04025
R36684 VDD.n4449 VDD.n4448 0.04025
R36685 VDD.n4450 VDD.n4449 0.04025
R36686 VDD.n4450 VDD.n2471 0.04025
R36687 VDD.n4454 VDD.n2471 0.04025
R36688 VDD.n4455 VDD.n4454 0.04025
R36689 VDD.n4456 VDD.n4455 0.04025
R36690 VDD.n4456 VDD.n2469 0.04025
R36691 VDD.n4460 VDD.n2469 0.04025
R36692 VDD.n4461 VDD.n4460 0.04025
R36693 VDD.n4462 VDD.n4461 0.04025
R36694 VDD.n4462 VDD.n2467 0.04025
R36695 VDD.n4466 VDD.n2467 0.04025
R36696 VDD.n4467 VDD.n4466 0.04025
R36697 VDD.n4468 VDD.n4467 0.04025
R36698 VDD.n4468 VDD.n2465 0.04025
R36699 VDD.n4472 VDD.n2465 0.04025
R36700 VDD.n4473 VDD.n4472 0.04025
R36701 VDD.n4474 VDD.n4473 0.04025
R36702 VDD.n4474 VDD.n2463 0.04025
R36703 VDD.n4478 VDD.n2463 0.04025
R36704 VDD.n4479 VDD.n4478 0.04025
R36705 VDD.n4480 VDD.n4479 0.04025
R36706 VDD.n4480 VDD.n2461 0.04025
R36707 VDD.n4484 VDD.n2461 0.04025
R36708 VDD.n4485 VDD.n4484 0.04025
R36709 VDD.n4486 VDD.n4485 0.04025
R36710 VDD.n4486 VDD.n2459 0.04025
R36711 VDD.n4490 VDD.n2459 0.04025
R36712 VDD.n4491 VDD.n4490 0.04025
R36713 VDD.n4492 VDD.n4491 0.04025
R36714 VDD.n4492 VDD.n2457 0.04025
R36715 VDD.n4496 VDD.n2457 0.04025
R36716 VDD.n4497 VDD.n4496 0.04025
R36717 VDD.n4498 VDD.n4497 0.04025
R36718 VDD.n4498 VDD.n2455 0.04025
R36719 VDD.n4502 VDD.n2455 0.04025
R36720 VDD.n4503 VDD.n4502 0.04025
R36721 VDD.n4504 VDD.n4503 0.04025
R36722 VDD.n4504 VDD.n2453 0.04025
R36723 VDD.n4508 VDD.n2453 0.04025
R36724 VDD.n4509 VDD.n4508 0.04025
R36725 VDD.n4510 VDD.n4509 0.04025
R36726 VDD.n4510 VDD.n2451 0.04025
R36727 VDD.n4514 VDD.n2451 0.04025
R36728 VDD.n4515 VDD.n4514 0.04025
R36729 VDD.n4516 VDD.n4515 0.04025
R36730 VDD.n4516 VDD.n2449 0.04025
R36731 VDD.n4520 VDD.n2449 0.04025
R36732 VDD.n4521 VDD.n4520 0.04025
R36733 VDD.n4522 VDD.n4521 0.04025
R36734 VDD.n4522 VDD.n2447 0.04025
R36735 VDD.n4526 VDD.n2447 0.04025
R36736 VDD.n4527 VDD.n4526 0.04025
R36737 VDD.n4528 VDD.n4527 0.04025
R36738 VDD.n4528 VDD.n2445 0.04025
R36739 VDD.n4532 VDD.n2445 0.04025
R36740 VDD.n4533 VDD.n4532 0.04025
R36741 VDD.n4534 VDD.n4533 0.04025
R36742 VDD.n4534 VDD.n2443 0.04025
R36743 VDD.n4538 VDD.n2443 0.04025
R36744 VDD.n4539 VDD.n4538 0.04025
R36745 VDD.n4540 VDD.n4539 0.04025
R36746 VDD.n4540 VDD.n2441 0.04025
R36747 VDD.n4544 VDD.n2441 0.04025
R36748 VDD.n4545 VDD.n4544 0.04025
R36749 VDD.n4546 VDD.n4545 0.04025
R36750 VDD.n4546 VDD.n2439 0.04025
R36751 VDD.n4550 VDD.n2439 0.04025
R36752 VDD.n4551 VDD.n4550 0.04025
R36753 VDD.n4552 VDD.n4551 0.04025
R36754 VDD.n4552 VDD.n2437 0.04025
R36755 VDD.n4556 VDD.n2437 0.04025
R36756 VDD.n4557 VDD.n4556 0.04025
R36757 VDD.n4558 VDD.n4557 0.04025
R36758 VDD.n4558 VDD.n2435 0.04025
R36759 VDD.n4562 VDD.n2435 0.04025
R36760 VDD.n4563 VDD.n4562 0.04025
R36761 VDD.n4564 VDD.n4563 0.04025
R36762 VDD.n4564 VDD.n2433 0.04025
R36763 VDD.n4568 VDD.n2433 0.04025
R36764 VDD.n4569 VDD.n4568 0.04025
R36765 VDD.n4570 VDD.n4569 0.04025
R36766 VDD.n4570 VDD.n2431 0.04025
R36767 VDD.n4574 VDD.n2431 0.04025
R36768 VDD.n4575 VDD.n4574 0.04025
R36769 VDD.n4576 VDD.n4575 0.04025
R36770 VDD.n4576 VDD.n2429 0.04025
R36771 VDD.n4580 VDD.n2429 0.04025
R36772 VDD.n4581 VDD.n4580 0.04025
R36773 VDD.n4582 VDD.n4581 0.04025
R36774 VDD.n4582 VDD.n2427 0.04025
R36775 VDD.n4586 VDD.n2427 0.04025
R36776 VDD.n4587 VDD.n4586 0.04025
R36777 VDD.n4588 VDD.n4587 0.04025
R36778 VDD.n4588 VDD.n2425 0.04025
R36779 VDD.n4593 VDD.n4592 0.04025
R36780 VDD.n4595 VDD.n4594 0.04025
R36781 VDD.n5219 VDD.n4595 0.04025
R36782 VDD.n5219 VDD.n5204 0.04025
R36783 VDD.n5199 VDD.n4599 0.04025
R36784 VDD.n5199 VDD.n5198 0.04025
R36785 VDD.n5198 VDD.n5197 0.04025
R36786 VDD.n5197 VDD.n4600 0.04025
R36787 VDD.n5193 VDD.n4600 0.04025
R36788 VDD.n5193 VDD.n5192 0.04025
R36789 VDD.n5192 VDD.n5191 0.04025
R36790 VDD.n5191 VDD.n4602 0.04025
R36791 VDD.n5187 VDD.n4602 0.04025
R36792 VDD.n5187 VDD.n5186 0.04025
R36793 VDD.n5186 VDD.n5185 0.04025
R36794 VDD.n5185 VDD.n4604 0.04025
R36795 VDD.n5181 VDD.n4604 0.04025
R36796 VDD.n5181 VDD.n5180 0.04025
R36797 VDD.n5180 VDD.n5179 0.04025
R36798 VDD.n5179 VDD.n4606 0.04025
R36799 VDD.n5175 VDD.n4606 0.04025
R36800 VDD.n5175 VDD.n5174 0.04025
R36801 VDD.n5174 VDD.n5173 0.04025
R36802 VDD.n5173 VDD.n4608 0.04025
R36803 VDD.n5169 VDD.n4608 0.04025
R36804 VDD.n5169 VDD.n5168 0.04025
R36805 VDD.n5168 VDD.n5167 0.04025
R36806 VDD.n5167 VDD.n4610 0.04025
R36807 VDD.n5163 VDD.n4610 0.04025
R36808 VDD.n5163 VDD.n5162 0.04025
R36809 VDD.n5162 VDD.n5161 0.04025
R36810 VDD.n5161 VDD.n4612 0.04025
R36811 VDD.n5157 VDD.n4612 0.04025
R36812 VDD.n5157 VDD.n5156 0.04025
R36813 VDD.n5156 VDD.n5155 0.04025
R36814 VDD.n5155 VDD.n4614 0.04025
R36815 VDD.n5151 VDD.n4614 0.04025
R36816 VDD.n5151 VDD.n5150 0.04025
R36817 VDD.n5150 VDD.n5149 0.04025
R36818 VDD.n5149 VDD.n4616 0.04025
R36819 VDD.n5145 VDD.n4616 0.04025
R36820 VDD.n5145 VDD.n5144 0.04025
R36821 VDD.n5144 VDD.n5143 0.04025
R36822 VDD.n5143 VDD.n4618 0.04025
R36823 VDD.n5139 VDD.n4618 0.04025
R36824 VDD.n5139 VDD.n5138 0.04025
R36825 VDD.n5138 VDD.n5137 0.04025
R36826 VDD.n5137 VDD.n4620 0.04025
R36827 VDD.n5133 VDD.n4620 0.04025
R36828 VDD.n5133 VDD.n5132 0.04025
R36829 VDD.n5132 VDD.n5131 0.04025
R36830 VDD.n5131 VDD.n4622 0.04025
R36831 VDD.n5127 VDD.n4622 0.04025
R36832 VDD.n5127 VDD.n5126 0.04025
R36833 VDD.n5126 VDD.n5125 0.04025
R36834 VDD.n5125 VDD.n4624 0.04025
R36835 VDD.n5121 VDD.n4624 0.04025
R36836 VDD.n5121 VDD.n5120 0.04025
R36837 VDD.n5120 VDD.n5119 0.04025
R36838 VDD.n5119 VDD.n4626 0.04025
R36839 VDD.n5115 VDD.n4626 0.04025
R36840 VDD.n5115 VDD.n5114 0.04025
R36841 VDD.n5114 VDD.n5113 0.04025
R36842 VDD.n5113 VDD.n4628 0.04025
R36843 VDD.n5109 VDD.n4628 0.04025
R36844 VDD.n5109 VDD.n5108 0.04025
R36845 VDD.n5108 VDD.n5107 0.04025
R36846 VDD.n5107 VDD.n4630 0.04025
R36847 VDD.n5103 VDD.n4630 0.04025
R36848 VDD.n5103 VDD.n5102 0.04025
R36849 VDD.n5102 VDD.n5101 0.04025
R36850 VDD.n5101 VDD.n4632 0.04025
R36851 VDD.n5097 VDD.n4632 0.04025
R36852 VDD.n5097 VDD.n5096 0.04025
R36853 VDD.n5096 VDD.n5095 0.04025
R36854 VDD.n5095 VDD.n4634 0.04025
R36855 VDD.n5091 VDD.n4634 0.04025
R36856 VDD.n5091 VDD.n5090 0.04025
R36857 VDD.n5090 VDD.n5089 0.04025
R36858 VDD.n5089 VDD.n4636 0.04025
R36859 VDD.n5085 VDD.n4636 0.04025
R36860 VDD.n5085 VDD.n5084 0.04025
R36861 VDD.n5084 VDD.n5083 0.04025
R36862 VDD.n5083 VDD.n4638 0.04025
R36863 VDD.n5079 VDD.n4638 0.04025
R36864 VDD.n5079 VDD.n5078 0.04025
R36865 VDD.n5078 VDD.n5077 0.04025
R36866 VDD.n5077 VDD.n4640 0.04025
R36867 VDD.n5073 VDD.n4640 0.04025
R36868 VDD.n5073 VDD.n5072 0.04025
R36869 VDD.n5072 VDD.n5071 0.04025
R36870 VDD.n5071 VDD.n4642 0.04025
R36871 VDD.n5067 VDD.n4642 0.04025
R36872 VDD.n5067 VDD.n5066 0.04025
R36873 VDD.n5066 VDD.n5065 0.04025
R36874 VDD.n5065 VDD.n4644 0.04025
R36875 VDD.n5061 VDD.n4644 0.04025
R36876 VDD.n5061 VDD.n5060 0.04025
R36877 VDD.n5060 VDD.n5059 0.04025
R36878 VDD.n5059 VDD.n4646 0.04025
R36879 VDD.n5055 VDD.n4646 0.04025
R36880 VDD.n5055 VDD.n5054 0.04025
R36881 VDD.n5054 VDD.n5053 0.04025
R36882 VDD.n5053 VDD.n4648 0.04025
R36883 VDD.n5049 VDD.n4648 0.04025
R36884 VDD.n5049 VDD.n5048 0.04025
R36885 VDD.n5048 VDD.n5047 0.04025
R36886 VDD.n5047 VDD.n4650 0.04025
R36887 VDD.n5043 VDD.n4650 0.04025
R36888 VDD.n5043 VDD.n5042 0.04025
R36889 VDD.n5042 VDD.n5041 0.04025
R36890 VDD.n5041 VDD.n4652 0.04025
R36891 VDD.n5037 VDD.n4652 0.04025
R36892 VDD.n5037 VDD.n5036 0.04025
R36893 VDD.n5036 VDD.n5035 0.04025
R36894 VDD.n5035 VDD.n4654 0.04025
R36895 VDD.n5031 VDD.n4654 0.04025
R36896 VDD.n5031 VDD.n5030 0.04025
R36897 VDD.n5030 VDD.n5029 0.04025
R36898 VDD.n5029 VDD.n4656 0.04025
R36899 VDD.n5025 VDD.n4656 0.04025
R36900 VDD.n5025 VDD.n5024 0.04025
R36901 VDD.n5024 VDD.n5023 0.04025
R36902 VDD.n5023 VDD.n4658 0.04025
R36903 VDD.n5019 VDD.n4658 0.04025
R36904 VDD.n5019 VDD.n5018 0.04025
R36905 VDD.n5018 VDD.n5017 0.04025
R36906 VDD.n5017 VDD.n4660 0.04025
R36907 VDD.n5013 VDD.n4660 0.04025
R36908 VDD.n5013 VDD.n5012 0.04025
R36909 VDD.n5012 VDD.n5011 0.04025
R36910 VDD.n5011 VDD.n4662 0.04025
R36911 VDD.n5007 VDD.n4662 0.04025
R36912 VDD.n5007 VDD.n5006 0.04025
R36913 VDD.n5006 VDD.n5005 0.04025
R36914 VDD.n5005 VDD.n4664 0.04025
R36915 VDD.n5001 VDD.n4664 0.04025
R36916 VDD.n5001 VDD.n5000 0.04025
R36917 VDD.n5000 VDD.n4999 0.04025
R36918 VDD.n4999 VDD.n4666 0.04025
R36919 VDD.n4995 VDD.n4666 0.04025
R36920 VDD.n4995 VDD.n4994 0.04025
R36921 VDD.n4994 VDD.n4993 0.04025
R36922 VDD.n4993 VDD.n4668 0.04025
R36923 VDD.n4989 VDD.n4668 0.04025
R36924 VDD.n4989 VDD.n4988 0.04025
R36925 VDD.n4988 VDD.n4987 0.04025
R36926 VDD.n4987 VDD.n4670 0.04025
R36927 VDD.n4983 VDD.n4670 0.04025
R36928 VDD.n4983 VDD.n4982 0.04025
R36929 VDD.n4982 VDD.n4981 0.04025
R36930 VDD.n4981 VDD.n4672 0.04025
R36931 VDD.n4977 VDD.n4672 0.04025
R36932 VDD.n4977 VDD.n4976 0.04025
R36933 VDD.n4976 VDD.n4975 0.04025
R36934 VDD.n4975 VDD.n4674 0.04025
R36935 VDD.n4971 VDD.n4674 0.04025
R36936 VDD.n4971 VDD.n4970 0.04025
R36937 VDD.n4970 VDD.n4969 0.04025
R36938 VDD.n4969 VDD.n4676 0.04025
R36939 VDD.n4965 VDD.n4676 0.04025
R36940 VDD.n4965 VDD.n4964 0.04025
R36941 VDD.n4964 VDD.n4963 0.04025
R36942 VDD.n4963 VDD.n4678 0.04025
R36943 VDD.n4959 VDD.n4678 0.04025
R36944 VDD.n4959 VDD.n4958 0.04025
R36945 VDD.n4958 VDD.n4957 0.04025
R36946 VDD.n4957 VDD.n4680 0.04025
R36947 VDD.n4953 VDD.n4680 0.04025
R36948 VDD.n4953 VDD.n4952 0.04025
R36949 VDD.n4952 VDD.n4951 0.04025
R36950 VDD.n4951 VDD.n4682 0.04025
R36951 VDD.n4947 VDD.n4682 0.04025
R36952 VDD.n4947 VDD.n4946 0.04025
R36953 VDD.n4946 VDD.n4945 0.04025
R36954 VDD.n4945 VDD.n4684 0.04025
R36955 VDD.n4941 VDD.n4684 0.04025
R36956 VDD.n4941 VDD.n4940 0.04025
R36957 VDD.n4940 VDD.n4939 0.04025
R36958 VDD.n4939 VDD.n4686 0.04025
R36959 VDD.n4935 VDD.n4686 0.04025
R36960 VDD.n4935 VDD.n4934 0.04025
R36961 VDD.n4934 VDD.n4933 0.04025
R36962 VDD.n4933 VDD.n4688 0.04025
R36963 VDD.n4929 VDD.n4688 0.04025
R36964 VDD.n4929 VDD.n4928 0.04025
R36965 VDD.n4928 VDD.n4927 0.04025
R36966 VDD.n4927 VDD.n4690 0.04025
R36967 VDD.n4923 VDD.n4690 0.04025
R36968 VDD.n4923 VDD.n4922 0.04025
R36969 VDD.n4922 VDD.n4921 0.04025
R36970 VDD.n4921 VDD.n4692 0.04025
R36971 VDD.n4917 VDD.n4692 0.04025
R36972 VDD.n4917 VDD.n4916 0.04025
R36973 VDD.n4916 VDD.n4915 0.04025
R36974 VDD.n4915 VDD.n4694 0.04025
R36975 VDD.n4911 VDD.n4694 0.04025
R36976 VDD.n4911 VDD.n4910 0.04025
R36977 VDD.n4910 VDD.n4909 0.04025
R36978 VDD.n4909 VDD.n4696 0.04025
R36979 VDD.n4905 VDD.n4696 0.04025
R36980 VDD.n3628 VDD.n3627 0.04025
R36981 VDD.n3627 VDD.n3626 0.04025
R36982 VDD.n3626 VDD.n2747 0.04025
R36983 VDD.n3622 VDD.n2747 0.04025
R36984 VDD.n3622 VDD.n3621 0.04025
R36985 VDD.n3621 VDD.n3620 0.04025
R36986 VDD.n3620 VDD.n2749 0.04025
R36987 VDD.n3616 VDD.n2749 0.04025
R36988 VDD.n3616 VDD.n3615 0.04025
R36989 VDD.n3615 VDD.n3614 0.04025
R36990 VDD.n3614 VDD.n2751 0.04025
R36991 VDD.n3610 VDD.n2751 0.04025
R36992 VDD.n3610 VDD.n3609 0.04025
R36993 VDD.n3609 VDD.n3608 0.04025
R36994 VDD.n3608 VDD.n2753 0.04025
R36995 VDD.n3604 VDD.n2753 0.04025
R36996 VDD.n3604 VDD.n3603 0.04025
R36997 VDD.n3603 VDD.n3602 0.04025
R36998 VDD.n3602 VDD.n2755 0.04025
R36999 VDD.n3598 VDD.n2755 0.04025
R37000 VDD.n3598 VDD.n3597 0.04025
R37001 VDD.n3597 VDD.n3596 0.04025
R37002 VDD.n3596 VDD.n2757 0.04025
R37003 VDD.n3592 VDD.n2757 0.04025
R37004 VDD.n3592 VDD.n3591 0.04025
R37005 VDD.n3591 VDD.n3590 0.04025
R37006 VDD.n3590 VDD.n2759 0.04025
R37007 VDD.n3586 VDD.n2759 0.04025
R37008 VDD.n3586 VDD.n3585 0.04025
R37009 VDD.n3585 VDD.n3584 0.04025
R37010 VDD.n3584 VDD.n2761 0.04025
R37011 VDD.n3580 VDD.n2761 0.04025
R37012 VDD.n3580 VDD.n3579 0.04025
R37013 VDD.n3579 VDD.n3578 0.04025
R37014 VDD.n3578 VDD.n2763 0.04025
R37015 VDD.n3574 VDD.n2763 0.04025
R37016 VDD.n3574 VDD.n3573 0.04025
R37017 VDD.n3573 VDD.n3572 0.04025
R37018 VDD.n3572 VDD.n2765 0.04025
R37019 VDD.n3568 VDD.n2765 0.04025
R37020 VDD.n3568 VDD.n3567 0.04025
R37021 VDD.n3567 VDD.n3566 0.04025
R37022 VDD.n3566 VDD.n2767 0.04025
R37023 VDD.n3562 VDD.n2767 0.04025
R37024 VDD.n3562 VDD.n3561 0.04025
R37025 VDD.n3561 VDD.n3560 0.04025
R37026 VDD.n3560 VDD.n2769 0.04025
R37027 VDD.n3556 VDD.n2769 0.04025
R37028 VDD.n3556 VDD.n3555 0.04025
R37029 VDD.n3555 VDD.n3554 0.04025
R37030 VDD.n3554 VDD.n2771 0.04025
R37031 VDD.n3550 VDD.n2771 0.04025
R37032 VDD.n3550 VDD.n3549 0.04025
R37033 VDD.n3549 VDD.n3548 0.04025
R37034 VDD.n3548 VDD.n2773 0.04025
R37035 VDD.n3544 VDD.n2773 0.04025
R37036 VDD.n3544 VDD.n3543 0.04025
R37037 VDD.n3543 VDD.n3542 0.04025
R37038 VDD.n3542 VDD.n2775 0.04025
R37039 VDD.n3538 VDD.n2775 0.04025
R37040 VDD.n3538 VDD.n3537 0.04025
R37041 VDD.n3537 VDD.n3536 0.04025
R37042 VDD.n3536 VDD.n2777 0.04025
R37043 VDD.n3532 VDD.n2777 0.04025
R37044 VDD.n3532 VDD.n3531 0.04025
R37045 VDD.n3531 VDD.n3530 0.04025
R37046 VDD.n3530 VDD.n2779 0.04025
R37047 VDD.n3526 VDD.n2779 0.04025
R37048 VDD.n3526 VDD.n3525 0.04025
R37049 VDD.n3525 VDD.n3524 0.04025
R37050 VDD.n3524 VDD.n2781 0.04025
R37051 VDD.n3520 VDD.n2781 0.04025
R37052 VDD.n3520 VDD.n3519 0.04025
R37053 VDD.n3519 VDD.n3518 0.04025
R37054 VDD.n3518 VDD.n2783 0.04025
R37055 VDD.n3514 VDD.n2783 0.04025
R37056 VDD.n3514 VDD.n3513 0.04025
R37057 VDD.n3513 VDD.n3512 0.04025
R37058 VDD.n3512 VDD.n2785 0.04025
R37059 VDD.n3508 VDD.n2785 0.04025
R37060 VDD.n3508 VDD.n3507 0.04025
R37061 VDD.n3507 VDD.n3506 0.04025
R37062 VDD.n3506 VDD.n2787 0.04025
R37063 VDD.n3502 VDD.n2787 0.04025
R37064 VDD.n3502 VDD.n3501 0.04025
R37065 VDD.n3501 VDD.n3500 0.04025
R37066 VDD.n3500 VDD.n2789 0.04025
R37067 VDD.n3496 VDD.n2789 0.04025
R37068 VDD.n3496 VDD.n3495 0.04025
R37069 VDD.n3495 VDD.n3494 0.04025
R37070 VDD.n3494 VDD.n2791 0.04025
R37071 VDD.n3490 VDD.n2791 0.04025
R37072 VDD.n3490 VDD.n3489 0.04025
R37073 VDD.n3489 VDD.n3488 0.04025
R37074 VDD.n3488 VDD.n2793 0.04025
R37075 VDD.n3484 VDD.n2793 0.04025
R37076 VDD.n3484 VDD.n3483 0.04025
R37077 VDD.n3483 VDD.n3482 0.04025
R37078 VDD.n3482 VDD.n2795 0.04025
R37079 VDD.n3478 VDD.n2795 0.04025
R37080 VDD.n3478 VDD.n3477 0.04025
R37081 VDD.n3477 VDD.n3476 0.04025
R37082 VDD.n3476 VDD.n2797 0.04025
R37083 VDD.n3472 VDD.n2797 0.04025
R37084 VDD.n3472 VDD.n3471 0.04025
R37085 VDD.n3471 VDD.n3470 0.04025
R37086 VDD.n3470 VDD.n2799 0.04025
R37087 VDD.n3466 VDD.n2799 0.04025
R37088 VDD.n3466 VDD.n3465 0.04025
R37089 VDD.n3465 VDD.n3464 0.04025
R37090 VDD.n3464 VDD.n2801 0.04025
R37091 VDD.n3460 VDD.n2801 0.04025
R37092 VDD.n3460 VDD.n3459 0.04025
R37093 VDD.n3459 VDD.n3458 0.04025
R37094 VDD.n3458 VDD.n2803 0.04025
R37095 VDD.n3454 VDD.n2803 0.04025
R37096 VDD.n3454 VDD.n3453 0.04025
R37097 VDD.n3453 VDD.n3452 0.04025
R37098 VDD.n3452 VDD.n2805 0.04025
R37099 VDD.n3448 VDD.n2805 0.04025
R37100 VDD.n3448 VDD.n3447 0.04025
R37101 VDD.n3447 VDD.n3446 0.04025
R37102 VDD.n3446 VDD.n2807 0.04025
R37103 VDD.n3442 VDD.n2807 0.04025
R37104 VDD.n3442 VDD.n3441 0.04025
R37105 VDD.n3441 VDD.n3440 0.04025
R37106 VDD.n3440 VDD.n2809 0.04025
R37107 VDD.n3436 VDD.n2809 0.04025
R37108 VDD.n3436 VDD.n3435 0.04025
R37109 VDD.n3435 VDD.n3434 0.04025
R37110 VDD.n3434 VDD.n2811 0.04025
R37111 VDD.n3430 VDD.n2811 0.04025
R37112 VDD.n3430 VDD.n3429 0.04025
R37113 VDD.n3429 VDD.n3428 0.04025
R37114 VDD.n3428 VDD.n2813 0.04025
R37115 VDD.n3424 VDD.n2813 0.04025
R37116 VDD.n3424 VDD.n3423 0.04025
R37117 VDD.n3423 VDD.n3422 0.04025
R37118 VDD.n3422 VDD.n2815 0.04025
R37119 VDD.n3418 VDD.n2815 0.04025
R37120 VDD.n3418 VDD.n3417 0.04025
R37121 VDD.n3417 VDD.n3416 0.04025
R37122 VDD.n3416 VDD.n2817 0.04025
R37123 VDD.n3412 VDD.n2817 0.04025
R37124 VDD.n3412 VDD.n3411 0.04025
R37125 VDD.n3411 VDD.n3410 0.04025
R37126 VDD.n3410 VDD.n2819 0.04025
R37127 VDD.n3406 VDD.n2819 0.04025
R37128 VDD.n3406 VDD.n3405 0.04025
R37129 VDD.n3405 VDD.n3404 0.04025
R37130 VDD.n3404 VDD.n2821 0.04025
R37131 VDD.n3400 VDD.n2821 0.04025
R37132 VDD.n3400 VDD.n3399 0.04025
R37133 VDD.n3399 VDD.n3398 0.04025
R37134 VDD.n3398 VDD.n2823 0.04025
R37135 VDD.n3394 VDD.n2823 0.04025
R37136 VDD.n3394 VDD.n3393 0.04025
R37137 VDD.n3393 VDD.n3392 0.04025
R37138 VDD.n3392 VDD.n2825 0.04025
R37139 VDD.n3388 VDD.n2825 0.04025
R37140 VDD.n3388 VDD.n3387 0.04025
R37141 VDD.n3387 VDD.n3386 0.04025
R37142 VDD.n3386 VDD.n2827 0.04025
R37143 VDD.n3382 VDD.n2827 0.04025
R37144 VDD.n3382 VDD.n3381 0.04025
R37145 VDD.n3381 VDD.n3380 0.04025
R37146 VDD.n3380 VDD.n2829 0.04025
R37147 VDD.n3376 VDD.n2829 0.04025
R37148 VDD.n3376 VDD.n3375 0.04025
R37149 VDD.n3375 VDD.n3374 0.04025
R37150 VDD.n3374 VDD.n2831 0.04025
R37151 VDD.n3370 VDD.n2831 0.04025
R37152 VDD.n3370 VDD.n3369 0.04025
R37153 VDD.n3369 VDD.n3368 0.04025
R37154 VDD.n3368 VDD.n2833 0.04025
R37155 VDD.n3364 VDD.n2833 0.04025
R37156 VDD.n3364 VDD.n3363 0.04025
R37157 VDD.n3363 VDD.n3362 0.04025
R37158 VDD.n3362 VDD.n2835 0.04025
R37159 VDD.n3358 VDD.n2835 0.04025
R37160 VDD.n3358 VDD.n3357 0.04025
R37161 VDD.n3357 VDD.n3356 0.04025
R37162 VDD.n3356 VDD.n2837 0.04025
R37163 VDD.n3352 VDD.n2837 0.04025
R37164 VDD.n3352 VDD.n3351 0.04025
R37165 VDD.n3351 VDD.n3350 0.04025
R37166 VDD.n3350 VDD.n2839 0.04025
R37167 VDD.n3346 VDD.n2839 0.04025
R37168 VDD.n3346 VDD.n3345 0.04025
R37169 VDD.n3345 VDD.n3344 0.04025
R37170 VDD.n3344 VDD.n2841 0.04025
R37171 VDD.n3340 VDD.n2841 0.04025
R37172 VDD.n3340 VDD.n3339 0.04025
R37173 VDD.n3339 VDD.n3338 0.04025
R37174 VDD.n3338 VDD.n2843 0.04025
R37175 VDD.n3334 VDD.n2843 0.04025
R37176 VDD.n3334 VDD.n3333 0.04025
R37177 VDD.n3333 VDD.n3332 0.04025
R37178 VDD.n3332 VDD.n2845 0.04025
R37179 VDD.n3328 VDD.n2845 0.04025
R37180 VDD.n3328 VDD.n3327 0.04025
R37181 VDD.n3327 VDD.n3326 0.04025
R37182 VDD.n3326 VDD.n2847 0.04025
R37183 VDD.n3322 VDD.n2847 0.04025
R37184 VDD.n3322 VDD.n3321 0.04025
R37185 VDD.n3321 VDD.n3320 0.04025
R37186 VDD.n3320 VDD.n2849 0.04025
R37187 VDD.n3316 VDD.n2849 0.04025
R37188 VDD.n3316 VDD.n3315 0.04025
R37189 VDD.n3315 VDD.n3314 0.04025
R37190 VDD.n3314 VDD.n2851 0.04025
R37191 VDD.n3310 VDD.n2851 0.04025
R37192 VDD.n3310 VDD.n3309 0.04025
R37193 VDD.n3309 VDD.n3308 0.04025
R37194 VDD.n3308 VDD.n2853 0.04025
R37195 VDD.n3304 VDD.n2853 0.04025
R37196 VDD.n3304 VDD.n3303 0.04025
R37197 VDD.n3303 VDD.n3302 0.04025
R37198 VDD.n3302 VDD.n2855 0.04025
R37199 VDD.n3298 VDD.n2855 0.04025
R37200 VDD.n3298 VDD.n3297 0.04025
R37201 VDD.n3297 VDD.n3296 0.04025
R37202 VDD.n3296 VDD.n2857 0.04025
R37203 VDD.n3292 VDD.n2857 0.04025
R37204 VDD.n3292 VDD.n3291 0.04025
R37205 VDD.n3291 VDD.n3290 0.04025
R37206 VDD.n3290 VDD.n2859 0.04025
R37207 VDD.n3286 VDD.n2859 0.04025
R37208 VDD.n3286 VDD.n3285 0.04025
R37209 VDD.n3285 VDD.n3284 0.04025
R37210 VDD.n3284 VDD.n2861 0.04025
R37211 VDD.n3280 VDD.n2861 0.04025
R37212 VDD.n3280 VDD.n3279 0.04025
R37213 VDD.n3279 VDD.n3278 0.04025
R37214 VDD.n3278 VDD.n2863 0.04025
R37215 VDD.n3274 VDD.n2863 0.04025
R37216 VDD.n3274 VDD.n3273 0.04025
R37217 VDD.n3273 VDD.n3272 0.04025
R37218 VDD.n3272 VDD.n2865 0.04025
R37219 VDD.n3268 VDD.n2865 0.04025
R37220 VDD.n3268 VDD.n3267 0.04025
R37221 VDD.n3267 VDD.n3266 0.04025
R37222 VDD.n3266 VDD.n2867 0.04025
R37223 VDD.n3262 VDD.n2867 0.04025
R37224 VDD.n3262 VDD.n3261 0.04025
R37225 VDD.n3261 VDD.n3260 0.04025
R37226 VDD.n3260 VDD.n2869 0.04025
R37227 VDD.n3256 VDD.n2869 0.04025
R37228 VDD.n3256 VDD.n3255 0.04025
R37229 VDD.n3255 VDD.n3254 0.04025
R37230 VDD.n3254 VDD.n2871 0.04025
R37231 VDD.n3250 VDD.n2871 0.04025
R37232 VDD.n3250 VDD.n3249 0.04025
R37233 VDD.n3249 VDD.n3248 0.04025
R37234 VDD.n3248 VDD.n2873 0.04025
R37235 VDD.n3244 VDD.n2873 0.04025
R37236 VDD.n3244 VDD.n3243 0.04025
R37237 VDD.n3243 VDD.n3242 0.04025
R37238 VDD.n3242 VDD.n2875 0.04025
R37239 VDD.n3238 VDD.n2875 0.04025
R37240 VDD.n3238 VDD.n3237 0.04025
R37241 VDD.n3237 VDD.n3236 0.04025
R37242 VDD.n3236 VDD.n2877 0.04025
R37243 VDD.n3232 VDD.n2877 0.04025
R37244 VDD.n3232 VDD.n3231 0.04025
R37245 VDD.n3231 VDD.n3230 0.04025
R37246 VDD.n3230 VDD.n2879 0.04025
R37247 VDD.n3226 VDD.n2879 0.04025
R37248 VDD.n3226 VDD.n3225 0.04025
R37249 VDD.n3225 VDD.n3224 0.04025
R37250 VDD.n3224 VDD.n2881 0.04025
R37251 VDD.n3220 VDD.n2881 0.04025
R37252 VDD.n3220 VDD.n3219 0.04025
R37253 VDD.n3219 VDD.n3218 0.04025
R37254 VDD.n3218 VDD.n2883 0.04025
R37255 VDD.n3214 VDD.n2883 0.04025
R37256 VDD.n3214 VDD.n3213 0.04025
R37257 VDD.n3213 VDD.n3212 0.04025
R37258 VDD.n3212 VDD.n2885 0.04025
R37259 VDD.n3208 VDD.n2885 0.04025
R37260 VDD.n3208 VDD.n3207 0.04025
R37261 VDD.n3207 VDD.n3206 0.04025
R37262 VDD.n3206 VDD.n2887 0.04025
R37263 VDD.n3202 VDD.n2887 0.04025
R37264 VDD.n3202 VDD.n3201 0.04025
R37265 VDD.n3201 VDD.n3200 0.04025
R37266 VDD.n3200 VDD.n2889 0.04025
R37267 VDD.n3196 VDD.n2889 0.04025
R37268 VDD.n3196 VDD.n3195 0.04025
R37269 VDD.n3195 VDD.n3194 0.04025
R37270 VDD.n3194 VDD.n2891 0.04025
R37271 VDD.n3190 VDD.n2891 0.04025
R37272 VDD.n3190 VDD.n3189 0.04025
R37273 VDD.n3189 VDD.n3188 0.04025
R37274 VDD.n3188 VDD.n2893 0.04025
R37275 VDD.n3184 VDD.n2893 0.04025
R37276 VDD.n3184 VDD.n3183 0.04025
R37277 VDD.n3183 VDD.n3182 0.04025
R37278 VDD.n3182 VDD.n2895 0.04025
R37279 VDD.n3178 VDD.n2895 0.04025
R37280 VDD.n3178 VDD.n3177 0.04025
R37281 VDD.n3177 VDD.n3176 0.04025
R37282 VDD.n3176 VDD.n2897 0.04025
R37283 VDD.n3172 VDD.n2897 0.04025
R37284 VDD.n3172 VDD.n3171 0.04025
R37285 VDD.n3171 VDD.n3170 0.04025
R37286 VDD.n3170 VDD.n2899 0.04025
R37287 VDD.n3166 VDD.n2899 0.04025
R37288 VDD.n3166 VDD.n3165 0.04025
R37289 VDD.n3165 VDD.n3164 0.04025
R37290 VDD.n3164 VDD.n2901 0.04025
R37291 VDD.n3160 VDD.n2901 0.04025
R37292 VDD.n3160 VDD.n3159 0.04025
R37293 VDD.n3159 VDD.n3158 0.04025
R37294 VDD.n3158 VDD.n2903 0.04025
R37295 VDD.n3154 VDD.n2903 0.04025
R37296 VDD.n3154 VDD.n3153 0.04025
R37297 VDD.n3153 VDD.n3152 0.04025
R37298 VDD.n3152 VDD.n2905 0.04025
R37299 VDD.n3148 VDD.n2905 0.04025
R37300 VDD.n3148 VDD.n3147 0.04025
R37301 VDD.n3147 VDD.n3146 0.04025
R37302 VDD.n3146 VDD.n2907 0.04025
R37303 VDD.n3142 VDD.n2907 0.04025
R37304 VDD.n3142 VDD.n3141 0.04025
R37305 VDD.n3141 VDD.n3140 0.04025
R37306 VDD.n3140 VDD.n2909 0.04025
R37307 VDD.n3136 VDD.n2909 0.04025
R37308 VDD.n3136 VDD.n3135 0.04025
R37309 VDD.n3135 VDD.n3134 0.04025
R37310 VDD.n3134 VDD.n2911 0.04025
R37311 VDD.n3130 VDD.n2911 0.04025
R37312 VDD.n3130 VDD.n3129 0.04025
R37313 VDD.n3129 VDD.n3128 0.04025
R37314 VDD.n3128 VDD.n2913 0.04025
R37315 VDD.n3124 VDD.n2913 0.04025
R37316 VDD.n3124 VDD.n3123 0.04025
R37317 VDD.n3123 VDD.n3122 0.04025
R37318 VDD.n3122 VDD.n2915 0.04025
R37319 VDD.n3118 VDD.n2915 0.04025
R37320 VDD.n3118 VDD.n3117 0.04025
R37321 VDD.n3117 VDD.n3116 0.04025
R37322 VDD.n3116 VDD.n2917 0.04025
R37323 VDD.n3112 VDD.n2917 0.04025
R37324 VDD.n3112 VDD.n3111 0.04025
R37325 VDD.n3111 VDD.n3110 0.04025
R37326 VDD.n3110 VDD.n2919 0.04025
R37327 VDD.n3106 VDD.n2919 0.04025
R37328 VDD.n3106 VDD.n3105 0.04025
R37329 VDD.n3105 VDD.n3104 0.04025
R37330 VDD.n3104 VDD.n2921 0.04025
R37331 VDD.n3100 VDD.n2921 0.04025
R37332 VDD.n3100 VDD.n3099 0.04025
R37333 VDD.n3099 VDD.n3098 0.04025
R37334 VDD.n3098 VDD.n2923 0.04025
R37335 VDD.n3094 VDD.n2923 0.04025
R37336 VDD.n3094 VDD.n3093 0.04025
R37337 VDD.n3093 VDD.n3092 0.04025
R37338 VDD.n3092 VDD.n2925 0.04025
R37339 VDD.n3088 VDD.n2925 0.04025
R37340 VDD.n3088 VDD.n3087 0.04025
R37341 VDD.n3087 VDD.n3086 0.04025
R37342 VDD.n3086 VDD.n2927 0.04025
R37343 VDD.n3082 VDD.n2927 0.04025
R37344 VDD.n3082 VDD.n3081 0.04025
R37345 VDD.n3081 VDD.n3080 0.04025
R37346 VDD.n3080 VDD.n2929 0.04025
R37347 VDD.n3076 VDD.n2929 0.04025
R37348 VDD.n3076 VDD.n3075 0.04025
R37349 VDD.n3075 VDD.n3074 0.04025
R37350 VDD.n3074 VDD.n2931 0.04025
R37351 VDD.n3070 VDD.n2931 0.04025
R37352 VDD.n3070 VDD.n3069 0.04025
R37353 VDD.n3069 VDD.n3068 0.04025
R37354 VDD.n3068 VDD.n2933 0.04025
R37355 VDD.n3064 VDD.n2933 0.04025
R37356 VDD.n3064 VDD.n3063 0.04025
R37357 VDD.n3063 VDD.n3062 0.04025
R37358 VDD.n3062 VDD.n2935 0.04025
R37359 VDD.n3058 VDD.n2935 0.04025
R37360 VDD.n3058 VDD.n3057 0.04025
R37361 VDD.n3057 VDD.n3056 0.04025
R37362 VDD.n3056 VDD.n2937 0.04025
R37363 VDD.n3052 VDD.n2937 0.04025
R37364 VDD.n3052 VDD.n3051 0.04025
R37365 VDD.n3051 VDD.n3050 0.04025
R37366 VDD.n3050 VDD.n2939 0.04025
R37367 VDD.n3046 VDD.n2939 0.04025
R37368 VDD.n3046 VDD.n3045 0.04025
R37369 VDD.n3045 VDD.n3044 0.04025
R37370 VDD.n3044 VDD.n2941 0.04025
R37371 VDD.n3040 VDD.n2941 0.04025
R37372 VDD.n3040 VDD.n3039 0.04025
R37373 VDD.n3039 VDD.n3038 0.04025
R37374 VDD.n3038 VDD.n2943 0.04025
R37375 VDD.n3034 VDD.n2943 0.04025
R37376 VDD.n3034 VDD.n3033 0.04025
R37377 VDD.n3033 VDD.n3032 0.04025
R37378 VDD.n3032 VDD.n2945 0.04025
R37379 VDD.n3028 VDD.n2945 0.04025
R37380 VDD.n3028 VDD.n3027 0.04025
R37381 VDD.n3027 VDD.n3026 0.04025
R37382 VDD.n3026 VDD.n2947 0.04025
R37383 VDD.n3022 VDD.n2947 0.04025
R37384 VDD.n3022 VDD.n3021 0.04025
R37385 VDD.n3021 VDD.n3020 0.04025
R37386 VDD.n3020 VDD.n2949 0.04025
R37387 VDD.n3016 VDD.n2949 0.04025
R37388 VDD.n3016 VDD.n3015 0.04025
R37389 VDD.n3015 VDD.n3014 0.04025
R37390 VDD.n3014 VDD.n2951 0.04025
R37391 VDD.n3010 VDD.n2951 0.04025
R37392 VDD.n3010 VDD.n3009 0.04025
R37393 VDD.n3009 VDD.n3008 0.04025
R37394 VDD.n3008 VDD.n2953 0.04025
R37395 VDD.n3004 VDD.n2953 0.04025
R37396 VDD.n3004 VDD.n3003 0.04025
R37397 VDD.n3003 VDD.n3002 0.04025
R37398 VDD.n3002 VDD.n2955 0.04025
R37399 VDD.n2998 VDD.n2955 0.04025
R37400 VDD.n2998 VDD.n2997 0.04025
R37401 VDD.n2997 VDD.n2996 0.04025
R37402 VDD.n2996 VDD.n2957 0.04025
R37403 VDD.n2992 VDD.n2957 0.04025
R37404 VDD.n2992 VDD.n2991 0.04025
R37405 VDD.n2991 VDD.n2990 0.04025
R37406 VDD.n2990 VDD.n2959 0.04025
R37407 VDD.n2986 VDD.n2959 0.04025
R37408 VDD.n2986 VDD.n2985 0.04025
R37409 VDD.n2985 VDD.n2984 0.04025
R37410 VDD.n2984 VDD.n2961 0.04025
R37411 VDD.n2980 VDD.n2961 0.04025
R37412 VDD.n2980 VDD.n2979 0.04025
R37413 VDD.n2979 VDD.n2978 0.04025
R37414 VDD.n2978 VDD.n2963 0.04025
R37415 VDD.n2974 VDD.n2963 0.04025
R37416 VDD.n2974 VDD.n2973 0.04025
R37417 VDD.n2973 VDD.n2972 0.04025
R37418 VDD.n2972 VDD.n2965 0.04025
R37419 VDD.n2968 VDD.n2965 0.04025
R37420 VDD.n2968 VDD.n2967 0.04025
R37421 VDD.n2967 VDD.n1767 0.04025
R37422 VDD.n11039 VDD.n1767 0.04025
R37423 VDD.n11042 VDD.n11039 0.04025
R37424 VDD.n11042 VDD.n11041 0.04025
R37425 VDD.n11041 VDD.n11040 0.04025
R37426 VDD.n11040 VDD.n668 0.04025
R37427 VDD.n11051 VDD.n668 0.04025
R37428 VDD.n11052 VDD.n11051 0.04025
R37429 VDD.n11053 VDD.n11052 0.04025
R37430 VDD.n11053 VDD.n666 0.04025
R37431 VDD.n11059 VDD.n666 0.04025
R37432 VDD.n11060 VDD.n11059 0.04025
R37433 VDD.n11061 VDD.n11060 0.04025
R37434 VDD.n11061 VDD.n664 0.04025
R37435 VDD.n11066 VDD.n664 0.04025
R37436 VDD.n11067 VDD.n11066 0.04025
R37437 VDD.n11068 VDD.n11067 0.04025
R37438 VDD.n11068 VDD.n662 0.04025
R37439 VDD.n11072 VDD.n662 0.04025
R37440 VDD.n11073 VDD.n11072 0.04025
R37441 VDD.n11073 VDD.n660 0.04025
R37442 VDD.n11079 VDD.n660 0.04025
R37443 VDD.n11080 VDD.n11079 0.04025
R37444 VDD.n11081 VDD.n11080 0.04025
R37445 VDD.n11081 VDD.n658 0.04025
R37446 VDD.n11085 VDD.n658 0.04025
R37447 VDD.n11086 VDD.n11085 0.04025
R37448 VDD.n11086 VDD.n656 0.04025
R37449 VDD.n11092 VDD.n656 0.04025
R37450 VDD.n11093 VDD.n11092 0.04025
R37451 VDD.n11094 VDD.n11093 0.04025
R37452 VDD.n11094 VDD.n654 0.04025
R37453 VDD.n11099 VDD.n654 0.04025
R37454 VDD.n11100 VDD.n11099 0.04025
R37455 VDD.n11101 VDD.n11100 0.04025
R37456 VDD.n11101 VDD.n652 0.04025
R37457 VDD.n11105 VDD.n652 0.04025
R37458 VDD.n11106 VDD.n11105 0.04025
R37459 VDD.n11106 VDD.n650 0.04025
R37460 VDD.n11110 VDD.n650 0.04025
R37461 VDD.n11111 VDD.n11110 0.04025
R37462 VDD.n11111 VDD.n647 0.04025
R37463 VDD.n11115 VDD.n647 0.04025
R37464 VDD.n11116 VDD.n11115 0.04025
R37465 VDD.n11117 VDD.n11116 0.04025
R37466 VDD.n11117 VDD.n645 0.04025
R37467 VDD.n11122 VDD.n645 0.04025
R37468 VDD.n11124 VDD.n11122 0.04025
R37469 VDD.n11125 VDD.n11124 0.04025
R37470 VDD.n11125 VDD.n632 0.04025
R37471 VDD.n11132 VDD.n632 0.04025
R37472 VDD.n11133 VDD.n11132 0.04025
R37473 VDD.n11134 VDD.n11133 0.04025
R37474 VDD.n11134 VDD.n630 0.04025
R37475 VDD.n11138 VDD.n630 0.04025
R37476 VDD.n11139 VDD.n11138 0.04025
R37477 VDD.n11140 VDD.n11139 0.04025
R37478 VDD.n11140 VDD.n628 0.04025
R37479 VDD.n11144 VDD.n628 0.04025
R37480 VDD.n11145 VDD.n11144 0.04025
R37481 VDD.n11146 VDD.n11145 0.04025
R37482 VDD.n11146 VDD.n626 0.04025
R37483 VDD.n11150 VDD.n626 0.04025
R37484 VDD.n11151 VDD.n11150 0.04025
R37485 VDD.n11152 VDD.n11151 0.04025
R37486 VDD.n11152 VDD.n624 0.04025
R37487 VDD.n11156 VDD.n624 0.04025
R37488 VDD.n11157 VDD.n11156 0.04025
R37489 VDD.n11158 VDD.n11157 0.04025
R37490 VDD.n11158 VDD.n622 0.04025
R37491 VDD.n11162 VDD.n622 0.04025
R37492 VDD.n11163 VDD.n11162 0.04025
R37493 VDD.n11164 VDD.n11163 0.04025
R37494 VDD.n11164 VDD.n620 0.04025
R37495 VDD.n11168 VDD.n620 0.04025
R37496 VDD.n11169 VDD.n11168 0.04025
R37497 VDD.n11170 VDD.n11169 0.04025
R37498 VDD.n11170 VDD.n618 0.04025
R37499 VDD.n11174 VDD.n618 0.04025
R37500 VDD.n11175 VDD.n11174 0.04025
R37501 VDD.n11176 VDD.n11175 0.04025
R37502 VDD.n11176 VDD.n616 0.04025
R37503 VDD.n11180 VDD.n616 0.04025
R37504 VDD.n11181 VDD.n11180 0.04025
R37505 VDD.n11182 VDD.n11181 0.04025
R37506 VDD.n11182 VDD.n614 0.04025
R37507 VDD.n11186 VDD.n614 0.04025
R37508 VDD.n11187 VDD.n11186 0.04025
R37509 VDD.n11188 VDD.n11187 0.04025
R37510 VDD.n11188 VDD.n612 0.04025
R37511 VDD.n11192 VDD.n612 0.04025
R37512 VDD.n11193 VDD.n11192 0.04025
R37513 VDD.n11194 VDD.n11193 0.04025
R37514 VDD.n11194 VDD.n610 0.04025
R37515 VDD.n11198 VDD.n610 0.04025
R37516 VDD.n11199 VDD.n11198 0.04025
R37517 VDD.n11200 VDD.n11199 0.04025
R37518 VDD.n11200 VDD.n608 0.04025
R37519 VDD.n11204 VDD.n608 0.04025
R37520 VDD.n11205 VDD.n11204 0.04025
R37521 VDD.n11206 VDD.n11205 0.04025
R37522 VDD.n11206 VDD.n606 0.04025
R37523 VDD.n11210 VDD.n606 0.04025
R37524 VDD.n11211 VDD.n11210 0.04025
R37525 VDD.n11212 VDD.n11211 0.04025
R37526 VDD.n11212 VDD.n604 0.04025
R37527 VDD.n11216 VDD.n604 0.04025
R37528 VDD.n11217 VDD.n11216 0.04025
R37529 VDD.n11218 VDD.n11217 0.04025
R37530 VDD.n11218 VDD.n602 0.04025
R37531 VDD.n11222 VDD.n602 0.04025
R37532 VDD.n11223 VDD.n11222 0.04025
R37533 VDD.n11224 VDD.n11223 0.04025
R37534 VDD.n11224 VDD.n600 0.04025
R37535 VDD.n11228 VDD.n600 0.04025
R37536 VDD.n11229 VDD.n11228 0.04025
R37537 VDD.n11230 VDD.n11229 0.04025
R37538 VDD.n11230 VDD.n598 0.04025
R37539 VDD.n11234 VDD.n598 0.04025
R37540 VDD.n11235 VDD.n11234 0.04025
R37541 VDD.n11236 VDD.n11235 0.04025
R37542 VDD.n11236 VDD.n596 0.04025
R37543 VDD.n11240 VDD.n596 0.04025
R37544 VDD.n11241 VDD.n11240 0.04025
R37545 VDD.n11242 VDD.n11241 0.04025
R37546 VDD.n11242 VDD.n594 0.04025
R37547 VDD.n11246 VDD.n594 0.04025
R37548 VDD.n11247 VDD.n11246 0.04025
R37549 VDD.n11248 VDD.n11247 0.04025
R37550 VDD.n11248 VDD.n592 0.04025
R37551 VDD.n11252 VDD.n592 0.04025
R37552 VDD.n11253 VDD.n11252 0.04025
R37553 VDD.n11254 VDD.n11253 0.04025
R37554 VDD.n11254 VDD.n590 0.04025
R37555 VDD.n11258 VDD.n590 0.04025
R37556 VDD.n11259 VDD.n11258 0.04025
R37557 VDD.n11260 VDD.n11259 0.04025
R37558 VDD.n11260 VDD.n588 0.04025
R37559 VDD.n11264 VDD.n588 0.04025
R37560 VDD.n11265 VDD.n11264 0.04025
R37561 VDD.n11266 VDD.n11265 0.04025
R37562 VDD.n11266 VDD.n586 0.04025
R37563 VDD.n11270 VDD.n586 0.04025
R37564 VDD.n11271 VDD.n11270 0.04025
R37565 VDD.n11272 VDD.n11271 0.04025
R37566 VDD.n11272 VDD.n584 0.04025
R37567 VDD.n11276 VDD.n584 0.04025
R37568 VDD.n11277 VDD.n11276 0.04025
R37569 VDD.n11278 VDD.n11277 0.04025
R37570 VDD.n11278 VDD.n582 0.04025
R37571 VDD.n11282 VDD.n582 0.04025
R37572 VDD.n11283 VDD.n11282 0.04025
R37573 VDD.n11284 VDD.n11283 0.04025
R37574 VDD.n11284 VDD.n580 0.04025
R37575 VDD.n11288 VDD.n580 0.04025
R37576 VDD.n11289 VDD.n11288 0.04025
R37577 VDD.n11290 VDD.n11289 0.04025
R37578 VDD.n11290 VDD.n578 0.04025
R37579 VDD.n11294 VDD.n578 0.04025
R37580 VDD.n11295 VDD.n11294 0.04025
R37581 VDD.n11296 VDD.n11295 0.04025
R37582 VDD.n11296 VDD.n576 0.04025
R37583 VDD.n11300 VDD.n576 0.04025
R37584 VDD.n11301 VDD.n11300 0.04025
R37585 VDD.n11302 VDD.n11301 0.04025
R37586 VDD.n11302 VDD.n574 0.04025
R37587 VDD.n11306 VDD.n574 0.04025
R37588 VDD.n11307 VDD.n11306 0.04025
R37589 VDD.n11308 VDD.n11307 0.04025
R37590 VDD.n11308 VDD.n572 0.04025
R37591 VDD.n11312 VDD.n572 0.04025
R37592 VDD.n11313 VDD.n11312 0.04025
R37593 VDD.n11314 VDD.n11313 0.04025
R37594 VDD.n11314 VDD.n570 0.04025
R37595 VDD.n11318 VDD.n570 0.04025
R37596 VDD.n11319 VDD.n11318 0.04025
R37597 VDD.n11320 VDD.n11319 0.04025
R37598 VDD.n11320 VDD.n568 0.04025
R37599 VDD.n11324 VDD.n568 0.04025
R37600 VDD.n11325 VDD.n11324 0.04025
R37601 VDD.n11326 VDD.n11325 0.04025
R37602 VDD.n11326 VDD.n566 0.04025
R37603 VDD.n11330 VDD.n566 0.04025
R37604 VDD.n11331 VDD.n11330 0.04025
R37605 VDD.n11332 VDD.n11331 0.04025
R37606 VDD.n11332 VDD.n564 0.04025
R37607 VDD.n11336 VDD.n564 0.04025
R37608 VDD.n11337 VDD.n11336 0.04025
R37609 VDD.n11338 VDD.n11337 0.04025
R37610 VDD.n11338 VDD.n562 0.04025
R37611 VDD.n11342 VDD.n562 0.04025
R37612 VDD.n11343 VDD.n11342 0.04025
R37613 VDD.n11344 VDD.n11343 0.04025
R37614 VDD.n11344 VDD.n560 0.04025
R37615 VDD.n11348 VDD.n560 0.04025
R37616 VDD.n11349 VDD.n11348 0.04025
R37617 VDD.n11350 VDD.n11349 0.04025
R37618 VDD.n11350 VDD.n558 0.04025
R37619 VDD.n11354 VDD.n558 0.04025
R37620 VDD.n11355 VDD.n11354 0.04025
R37621 VDD.n11356 VDD.n11355 0.04025
R37622 VDD.n11356 VDD.n556 0.04025
R37623 VDD.n11360 VDD.n556 0.04025
R37624 VDD.n11361 VDD.n11360 0.04025
R37625 VDD.n11362 VDD.n11361 0.04025
R37626 VDD.n11362 VDD.n554 0.04025
R37627 VDD.n11366 VDD.n554 0.04025
R37628 VDD.n11367 VDD.n11366 0.04025
R37629 VDD.n11368 VDD.n11367 0.04025
R37630 VDD.n11368 VDD.n552 0.04025
R37631 VDD.n11372 VDD.n552 0.04025
R37632 VDD.n11373 VDD.n11372 0.04025
R37633 VDD.n11374 VDD.n11373 0.04025
R37634 VDD.n11374 VDD.n550 0.04025
R37635 VDD.n11378 VDD.n550 0.04025
R37636 VDD.n11379 VDD.n11378 0.04025
R37637 VDD.n11380 VDD.n11379 0.04025
R37638 VDD.n11380 VDD.n548 0.04025
R37639 VDD.n11384 VDD.n548 0.04025
R37640 VDD.n11385 VDD.n11384 0.04025
R37641 VDD.n11386 VDD.n11385 0.04025
R37642 VDD.n11386 VDD.n546 0.04025
R37643 VDD.n11390 VDD.n546 0.04025
R37644 VDD.n11391 VDD.n11390 0.04025
R37645 VDD.n11392 VDD.n11391 0.04025
R37646 VDD.n11392 VDD.n544 0.04025
R37647 VDD.n11396 VDD.n544 0.04025
R37648 VDD.n11397 VDD.n11396 0.04025
R37649 VDD.n11398 VDD.n11397 0.04025
R37650 VDD.n11398 VDD.n542 0.04025
R37651 VDD.n11402 VDD.n542 0.04025
R37652 VDD.n11403 VDD.n11402 0.04025
R37653 VDD.n11404 VDD.n11403 0.04025
R37654 VDD.n11404 VDD.n540 0.04025
R37655 VDD.n11408 VDD.n540 0.04025
R37656 VDD.n11409 VDD.n11408 0.04025
R37657 VDD.n11410 VDD.n11409 0.04025
R37658 VDD.n11410 VDD.n538 0.04025
R37659 VDD.n11414 VDD.n538 0.04025
R37660 VDD.n11415 VDD.n11414 0.04025
R37661 VDD.n11416 VDD.n11415 0.04025
R37662 VDD.n11416 VDD.n536 0.04025
R37663 VDD.n11420 VDD.n536 0.04025
R37664 VDD.n11421 VDD.n11420 0.04025
R37665 VDD.n11422 VDD.n11421 0.04025
R37666 VDD.n11422 VDD.n534 0.04025
R37667 VDD.n11426 VDD.n534 0.04025
R37668 VDD.n11427 VDD.n11426 0.04025
R37669 VDD.n11428 VDD.n11427 0.04025
R37670 VDD.n11428 VDD.n532 0.04025
R37671 VDD.n11432 VDD.n532 0.04025
R37672 VDD.n11433 VDD.n11432 0.04025
R37673 VDD.n11434 VDD.n11433 0.04025
R37674 VDD.n11434 VDD.n530 0.04025
R37675 VDD.n11438 VDD.n530 0.04025
R37676 VDD.n11439 VDD.n11438 0.04025
R37677 VDD.n11440 VDD.n11439 0.04025
R37678 VDD.n11440 VDD.n528 0.04025
R37679 VDD.n11444 VDD.n528 0.04025
R37680 VDD.n11445 VDD.n11444 0.04025
R37681 VDD.n11446 VDD.n11445 0.04025
R37682 VDD.n11446 VDD.n526 0.04025
R37683 VDD.n11450 VDD.n526 0.04025
R37684 VDD.n11451 VDD.n11450 0.04025
R37685 VDD.n11452 VDD.n11451 0.04025
R37686 VDD.n11452 VDD.n524 0.04025
R37687 VDD.n11456 VDD.n524 0.04025
R37688 VDD.n11457 VDD.n11456 0.04025
R37689 VDD.n11458 VDD.n11457 0.04025
R37690 VDD.n11458 VDD.n522 0.04025
R37691 VDD.n11462 VDD.n522 0.04025
R37692 VDD.n11463 VDD.n11462 0.04025
R37693 VDD.n11464 VDD.n11463 0.04025
R37694 VDD.n11464 VDD.n520 0.04025
R37695 VDD.n11468 VDD.n520 0.04025
R37696 VDD.n11469 VDD.n11468 0.04025
R37697 VDD.n11470 VDD.n11469 0.04025
R37698 VDD.n11470 VDD.n518 0.04025
R37699 VDD.n11474 VDD.n518 0.04025
R37700 VDD.n11475 VDD.n11474 0.04025
R37701 VDD.n11476 VDD.n11475 0.04025
R37702 VDD.n11476 VDD.n516 0.04025
R37703 VDD.n11480 VDD.n516 0.04025
R37704 VDD.n11481 VDD.n11480 0.04025
R37705 VDD.n11482 VDD.n11481 0.04025
R37706 VDD.n11482 VDD.n514 0.04025
R37707 VDD.n11486 VDD.n514 0.04025
R37708 VDD.n11487 VDD.n11486 0.04025
R37709 VDD.n11488 VDD.n11487 0.04025
R37710 VDD.n11488 VDD.n512 0.04025
R37711 VDD.n11492 VDD.n512 0.04025
R37712 VDD.n11493 VDD.n11492 0.04025
R37713 VDD.n11494 VDD.n11493 0.04025
R37714 VDD.n11494 VDD.n510 0.04025
R37715 VDD.n11498 VDD.n510 0.04025
R37716 VDD.n11499 VDD.n11498 0.04025
R37717 VDD.n11500 VDD.n11499 0.04025
R37718 VDD.n11500 VDD.n508 0.04025
R37719 VDD.n11504 VDD.n508 0.04025
R37720 VDD.n11505 VDD.n11504 0.04025
R37721 VDD.n11506 VDD.n11505 0.04025
R37722 VDD.n11506 VDD.n506 0.04025
R37723 VDD.n11510 VDD.n506 0.04025
R37724 VDD.n11511 VDD.n11510 0.04025
R37725 VDD.n11512 VDD.n11511 0.04025
R37726 VDD.n11512 VDD.n504 0.04025
R37727 VDD.n11516 VDD.n504 0.04025
R37728 VDD.n11517 VDD.n11516 0.04025
R37729 VDD.n11518 VDD.n11517 0.04025
R37730 VDD.n11518 VDD.n502 0.04025
R37731 VDD.n11522 VDD.n502 0.04025
R37732 VDD.n11523 VDD.n11522 0.04025
R37733 VDD.n11524 VDD.n11523 0.04025
R37734 VDD.n11524 VDD.n500 0.04025
R37735 VDD.n11528 VDD.n500 0.04025
R37736 VDD.n11529 VDD.n11528 0.04025
R37737 VDD.n11530 VDD.n11529 0.04025
R37738 VDD.n11530 VDD.n498 0.04025
R37739 VDD.n11534 VDD.n498 0.04025
R37740 VDD.n11535 VDD.n11534 0.04025
R37741 VDD.n11536 VDD.n11535 0.04025
R37742 VDD.n11536 VDD.n496 0.04025
R37743 VDD.n11540 VDD.n496 0.04025
R37744 VDD.n11541 VDD.n11540 0.04025
R37745 VDD.n11542 VDD.n11541 0.04025
R37746 VDD.n11542 VDD.n494 0.04025
R37747 VDD.n11546 VDD.n494 0.04025
R37748 VDD.n11547 VDD.n11546 0.04025
R37749 VDD.n11548 VDD.n11547 0.04025
R37750 VDD.n11548 VDD.n492 0.04025
R37751 VDD.n11552 VDD.n492 0.04025
R37752 VDD.n11553 VDD.n11552 0.04025
R37753 VDD.n11554 VDD.n11553 0.04025
R37754 VDD.n11554 VDD.n490 0.04025
R37755 VDD.n11558 VDD.n490 0.04025
R37756 VDD.n11559 VDD.n11558 0.04025
R37757 VDD.n11560 VDD.n11559 0.04025
R37758 VDD.n11560 VDD.n488 0.04025
R37759 VDD.n11564 VDD.n488 0.04025
R37760 VDD.n11565 VDD.n11564 0.04025
R37761 VDD.n11566 VDD.n11565 0.04025
R37762 VDD.n11566 VDD.n486 0.04025
R37763 VDD.n11570 VDD.n486 0.04025
R37764 VDD.n11571 VDD.n11570 0.04025
R37765 VDD.n11572 VDD.n11571 0.04025
R37766 VDD.n11572 VDD.n484 0.04025
R37767 VDD.n11576 VDD.n484 0.04025
R37768 VDD.n11577 VDD.n11576 0.04025
R37769 VDD.n11578 VDD.n11577 0.04025
R37770 VDD.n11578 VDD.n482 0.04025
R37771 VDD.n11582 VDD.n482 0.04025
R37772 VDD.n11583 VDD.n11582 0.04025
R37773 VDD.n11584 VDD.n11583 0.04025
R37774 VDD.n11584 VDD.n480 0.04025
R37775 VDD.n11588 VDD.n480 0.04025
R37776 VDD.n11589 VDD.n11588 0.04025
R37777 VDD.n11590 VDD.n11589 0.04025
R37778 VDD.n11590 VDD.n478 0.04025
R37779 VDD.n11594 VDD.n478 0.04025
R37780 VDD.n11595 VDD.n11594 0.04025
R37781 VDD.n11596 VDD.n11595 0.04025
R37782 VDD.n11596 VDD.n476 0.04025
R37783 VDD.n11600 VDD.n476 0.04025
R37784 VDD.n11601 VDD.n11600 0.04025
R37785 VDD.n11602 VDD.n11601 0.04025
R37786 VDD.n11602 VDD.n474 0.04025
R37787 VDD.n11606 VDD.n474 0.04025
R37788 VDD.n11607 VDD.n11606 0.04025
R37789 VDD.n11608 VDD.n11607 0.04025
R37790 VDD.n11608 VDD.n472 0.04025
R37791 VDD.n11612 VDD.n472 0.04025
R37792 VDD.n11613 VDD.n11612 0.04025
R37793 VDD.n11614 VDD.n11613 0.04025
R37794 VDD.n11614 VDD.n470 0.04025
R37795 VDD.n11618 VDD.n470 0.04025
R37796 VDD.n11619 VDD.n11618 0.04025
R37797 VDD.n11620 VDD.n11619 0.04025
R37798 VDD.n11620 VDD.n468 0.04025
R37799 VDD.n11624 VDD.n468 0.04025
R37800 VDD.n11625 VDD.n11624 0.04025
R37801 VDD.n11626 VDD.n11625 0.04025
R37802 VDD.n11626 VDD.n466 0.04025
R37803 VDD.n11630 VDD.n466 0.04025
R37804 VDD.n11631 VDD.n11630 0.04025
R37805 VDD.n11632 VDD.n11631 0.04025
R37806 VDD.n11632 VDD.n464 0.04025
R37807 VDD.n11636 VDD.n464 0.04025
R37808 VDD.n11637 VDD.n11636 0.04025
R37809 VDD.n11638 VDD.n11637 0.04025
R37810 VDD.n11638 VDD.n462 0.04025
R37811 VDD.n11642 VDD.n462 0.04025
R37812 VDD.n11643 VDD.n11642 0.04025
R37813 VDD.n11644 VDD.n11643 0.04025
R37814 VDD.n11644 VDD.n460 0.04025
R37815 VDD.n11648 VDD.n460 0.04025
R37816 VDD.n11649 VDD.n11648 0.04025
R37817 VDD.n11650 VDD.n11649 0.04025
R37818 VDD.n11650 VDD.n458 0.04025
R37819 VDD.n11654 VDD.n458 0.04025
R37820 VDD.n11655 VDD.n11654 0.04025
R37821 VDD.n11656 VDD.n11655 0.04025
R37822 VDD.n11656 VDD.n456 0.04025
R37823 VDD.n11660 VDD.n456 0.04025
R37824 VDD.n11661 VDD.n11660 0.04025
R37825 VDD.n11662 VDD.n11661 0.04025
R37826 VDD.n11662 VDD.n454 0.04025
R37827 VDD.n11666 VDD.n454 0.04025
R37828 VDD.n11667 VDD.n11666 0.04025
R37829 VDD.n11668 VDD.n11667 0.04025
R37830 VDD.n11668 VDD.n452 0.04025
R37831 VDD.n11672 VDD.n452 0.04025
R37832 VDD.n11673 VDD.n11672 0.04025
R37833 VDD.n11674 VDD.n11673 0.04025
R37834 VDD.n11674 VDD.n450 0.04025
R37835 VDD.n11678 VDD.n450 0.04025
R37836 VDD.n11679 VDD.n11678 0.04025
R37837 VDD.n11680 VDD.n11679 0.04025
R37838 VDD.n11680 VDD.n448 0.04025
R37839 VDD.n11684 VDD.n448 0.04025
R37840 VDD.n11685 VDD.n11684 0.04025
R37841 VDD.n11686 VDD.n11685 0.04025
R37842 VDD.n11686 VDD.n446 0.04025
R37843 VDD.n11690 VDD.n446 0.04025
R37844 VDD.n11691 VDD.n11690 0.04025
R37845 VDD.n11692 VDD.n11691 0.04025
R37846 VDD.n11692 VDD.n444 0.04025
R37847 VDD.n11696 VDD.n444 0.04025
R37848 VDD.n11697 VDD.n11696 0.04025
R37849 VDD.n11698 VDD.n11697 0.04025
R37850 VDD.n11698 VDD.n442 0.04025
R37851 VDD.n11702 VDD.n442 0.04025
R37852 VDD.n11703 VDD.n11702 0.04025
R37853 VDD.n11704 VDD.n11703 0.04025
R37854 VDD.n11704 VDD.n440 0.04025
R37855 VDD.n11708 VDD.n440 0.04025
R37856 VDD.n11709 VDD.n11708 0.04025
R37857 VDD.n11710 VDD.n11709 0.04025
R37858 VDD.n11710 VDD.n438 0.04025
R37859 VDD.n11714 VDD.n438 0.04025
R37860 VDD.n11715 VDD.n11714 0.04025
R37861 VDD.n11716 VDD.n11715 0.04025
R37862 VDD.n11716 VDD.n436 0.04025
R37863 VDD.n11720 VDD.n436 0.04025
R37864 VDD.n11721 VDD.n11720 0.04025
R37865 VDD.n11722 VDD.n11721 0.04025
R37866 VDD.n11722 VDD.n434 0.04025
R37867 VDD.n11726 VDD.n434 0.04025
R37868 VDD.n11727 VDD.n11726 0.04025
R37869 VDD.n11728 VDD.n11727 0.04025
R37870 VDD.n11728 VDD.n432 0.04025
R37871 VDD.n11732 VDD.n432 0.04025
R37872 VDD.n11733 VDD.n11732 0.04025
R37873 VDD.n11734 VDD.n11733 0.04025
R37874 VDD.n11734 VDD.n430 0.04025
R37875 VDD.n11738 VDD.n430 0.04025
R37876 VDD.n11739 VDD.n11738 0.04025
R37877 VDD.n11740 VDD.n11739 0.04025
R37878 VDD.n11740 VDD.n428 0.04025
R37879 VDD.n11744 VDD.n428 0.04025
R37880 VDD.n11745 VDD.n11744 0.04025
R37881 VDD.n11746 VDD.n11745 0.04025
R37882 VDD.n11746 VDD.n426 0.04025
R37883 VDD.n11750 VDD.n426 0.04025
R37884 VDD.n11751 VDD.n11750 0.04025
R37885 VDD.n11752 VDD.n11751 0.04025
R37886 VDD.n11752 VDD.n424 0.04025
R37887 VDD.n11756 VDD.n424 0.04025
R37888 VDD.n11757 VDD.n11756 0.04025
R37889 VDD.n11758 VDD.n11757 0.04025
R37890 VDD.n11758 VDD.n422 0.04025
R37891 VDD.n11762 VDD.n422 0.04025
R37892 VDD.n11763 VDD.n11762 0.04025
R37893 VDD.n11764 VDD.n11763 0.04025
R37894 VDD.n11764 VDD.n420 0.04025
R37895 VDD.n11768 VDD.n420 0.04025
R37896 VDD.n11769 VDD.n11768 0.04025
R37897 VDD.n11770 VDD.n11769 0.04025
R37898 VDD.n11770 VDD.n418 0.04025
R37899 VDD.n11774 VDD.n418 0.04025
R37900 VDD.n11775 VDD.n11774 0.04025
R37901 VDD.n11776 VDD.n11775 0.04025
R37902 VDD.n11776 VDD.n416 0.04025
R37903 VDD.n11780 VDD.n416 0.04025
R37904 VDD.n11781 VDD.n11780 0.04025
R37905 VDD.n11782 VDD.n11781 0.04025
R37906 VDD.n11782 VDD.n414 0.04025
R37907 VDD.n11786 VDD.n414 0.04025
R37908 VDD.n11787 VDD.n11786 0.04025
R37909 VDD.n11788 VDD.n11787 0.04025
R37910 VDD.n11788 VDD.n412 0.04025
R37911 VDD.n11792 VDD.n412 0.04025
R37912 VDD.n11793 VDD.n11792 0.04025
R37913 VDD.n11794 VDD.n11793 0.04025
R37914 VDD.n11794 VDD.n410 0.04025
R37915 VDD.n11798 VDD.n410 0.04025
R37916 VDD.n11799 VDD.n11798 0.04025
R37917 VDD.n11800 VDD.n11799 0.04025
R37918 VDD.n11800 VDD.n408 0.04025
R37919 VDD.n11804 VDD.n408 0.04025
R37920 VDD.n11805 VDD.n11804 0.04025
R37921 VDD.n11806 VDD.n11805 0.04025
R37922 VDD.n11806 VDD.n406 0.04025
R37923 VDD.n11810 VDD.n406 0.04025
R37924 VDD.n11811 VDD.n11810 0.04025
R37925 VDD.n11812 VDD.n404 0.04025
R37926 VDD.n11816 VDD.n404 0.04025
R37927 VDD.n11817 VDD.n11816 0.04025
R37928 VDD.n11818 VDD.n11817 0.04025
R37929 VDD.n11818 VDD.n402 0.04025
R37930 VDD.n11822 VDD.n402 0.04025
R37931 VDD.n11823 VDD.n11822 0.04025
R37932 VDD.n11824 VDD.n11823 0.04025
R37933 VDD.n11824 VDD.n400 0.04025
R37934 VDD.n11828 VDD.n400 0.04025
R37935 VDD.n11829 VDD.n11828 0.04025
R37936 VDD.n11830 VDD.n11829 0.04025
R37937 VDD.n11830 VDD.n398 0.04025
R37938 VDD.n11834 VDD.n398 0.04025
R37939 VDD.n11835 VDD.n11834 0.04025
R37940 VDD.n11836 VDD.n11835 0.04025
R37941 VDD.n11836 VDD.n396 0.04025
R37942 VDD.n11840 VDD.n396 0.04025
R37943 VDD.n11841 VDD.n11840 0.04025
R37944 VDD.n11842 VDD.n11841 0.04025
R37945 VDD.n11842 VDD.n394 0.04025
R37946 VDD.n11846 VDD.n394 0.04025
R37947 VDD.n11847 VDD.n11846 0.04025
R37948 VDD.n11848 VDD.n11847 0.04025
R37949 VDD.n11848 VDD.n392 0.04025
R37950 VDD.n11852 VDD.n392 0.04025
R37951 VDD.n11853 VDD.n11852 0.04025
R37952 VDD.n11854 VDD.n11853 0.04025
R37953 VDD.n11854 VDD.n390 0.04025
R37954 VDD.n11858 VDD.n390 0.04025
R37955 VDD.n11859 VDD.n11858 0.04025
R37956 VDD.n11860 VDD.n11859 0.04025
R37957 VDD.n11860 VDD.n388 0.04025
R37958 VDD.n11864 VDD.n388 0.04025
R37959 VDD.n11865 VDD.n11864 0.04025
R37960 VDD.n11866 VDD.n11865 0.04025
R37961 VDD.n11866 VDD.n386 0.04025
R37962 VDD.n11870 VDD.n386 0.04025
R37963 VDD.n11871 VDD.n11870 0.04025
R37964 VDD.n11873 VDD.n11871 0.04025
R37965 VDD.n11877 VDD.n384 0.04025
R37966 VDD.n11878 VDD.n11877 0.04025
R37967 VDD.n11879 VDD.n11878 0.04025
R37968 VDD.n11879 VDD.n382 0.04025
R37969 VDD.n11883 VDD.n382 0.04025
R37970 VDD.n11884 VDD.n11883 0.04025
R37971 VDD.n11885 VDD.n11884 0.04025
R37972 VDD.n11885 VDD.n380 0.04025
R37973 VDD.n11889 VDD.n380 0.04025
R37974 VDD.n11890 VDD.n11889 0.04025
R37975 VDD.n11891 VDD.n11890 0.04025
R37976 VDD.n11891 VDD.n378 0.04025
R37977 VDD.n11895 VDD.n378 0.04025
R37978 VDD.n11896 VDD.n11895 0.04025
R37979 VDD.n11897 VDD.n11896 0.04025
R37980 VDD.n11897 VDD.n376 0.04025
R37981 VDD.n11901 VDD.n376 0.04025
R37982 VDD.n11902 VDD.n11901 0.04025
R37983 VDD.n11903 VDD.n11902 0.04025
R37984 VDD.n11903 VDD.n374 0.04025
R37985 VDD.n11907 VDD.n374 0.04025
R37986 VDD.n11908 VDD.n11907 0.04025
R37987 VDD.n11909 VDD.n11908 0.04025
R37988 VDD.n11909 VDD.n372 0.04025
R37989 VDD.n11913 VDD.n372 0.04025
R37990 VDD.n11914 VDD.n11913 0.04025
R37991 VDD.n11915 VDD.n11914 0.04025
R37992 VDD.n11915 VDD.n370 0.04025
R37993 VDD.n11919 VDD.n370 0.04025
R37994 VDD.n11920 VDD.n11919 0.04025
R37995 VDD.n11921 VDD.n11920 0.04025
R37996 VDD.n11921 VDD.n368 0.04025
R37997 VDD.n11925 VDD.n368 0.04025
R37998 VDD.n11926 VDD.n11925 0.04025
R37999 VDD.n11927 VDD.n11926 0.04025
R38000 VDD.n11927 VDD.n366 0.04025
R38001 VDD.n11931 VDD.n366 0.04025
R38002 VDD.n11932 VDD.n11931 0.04025
R38003 VDD.n11933 VDD.n11932 0.04025
R38004 VDD.n11933 VDD.n364 0.04025
R38005 VDD.n11937 VDD.n364 0.04025
R38006 VDD.n11938 VDD.n11937 0.04025
R38007 VDD.n11939 VDD.n11938 0.04025
R38008 VDD.n11939 VDD.n362 0.04025
R38009 VDD.n11943 VDD.n362 0.04025
R38010 VDD.n11944 VDD.n11943 0.04025
R38011 VDD.n11945 VDD.n11944 0.04025
R38012 VDD.n11945 VDD.n360 0.04025
R38013 VDD.n11949 VDD.n360 0.04025
R38014 VDD.n11950 VDD.n11949 0.04025
R38015 VDD.n11951 VDD.n11950 0.04025
R38016 VDD.n11951 VDD.n358 0.04025
R38017 VDD.n11955 VDD.n358 0.04025
R38018 VDD.n11956 VDD.n11955 0.04025
R38019 VDD.n11957 VDD.n11956 0.04025
R38020 VDD.n11957 VDD.n356 0.04025
R38021 VDD.n11961 VDD.n356 0.04025
R38022 VDD.n11962 VDD.n11961 0.04025
R38023 VDD.n11963 VDD.n11962 0.04025
R38024 VDD.n11963 VDD.n354 0.04025
R38025 VDD.n11967 VDD.n354 0.04025
R38026 VDD.n11968 VDD.n11967 0.04025
R38027 VDD.n11969 VDD.n11968 0.04025
R38028 VDD.n11969 VDD.n352 0.04025
R38029 VDD.n11973 VDD.n352 0.04025
R38030 VDD.n11974 VDD.n11973 0.04025
R38031 VDD.n11975 VDD.n11974 0.04025
R38032 VDD.n11975 VDD.n350 0.04025
R38033 VDD.n11979 VDD.n350 0.04025
R38034 VDD.n11980 VDD.n11979 0.04025
R38035 VDD.n11981 VDD.n11980 0.04025
R38036 VDD.n11981 VDD.n348 0.04025
R38037 VDD.n11985 VDD.n348 0.04025
R38038 VDD.n11986 VDD.n11985 0.04025
R38039 VDD.n11987 VDD.n11986 0.04025
R38040 VDD.n11987 VDD.n346 0.04025
R38041 VDD.n11991 VDD.n346 0.04025
R38042 VDD.n11992 VDD.n11991 0.04025
R38043 VDD.n11993 VDD.n11992 0.04025
R38044 VDD.n11993 VDD.n344 0.04025
R38045 VDD.n11997 VDD.n344 0.04025
R38046 VDD.n11998 VDD.n11997 0.04025
R38047 VDD.n11999 VDD.n11998 0.04025
R38048 VDD.n11999 VDD.n342 0.04025
R38049 VDD.n12003 VDD.n342 0.04025
R38050 VDD.n12004 VDD.n12003 0.04025
R38051 VDD.n12005 VDD.n12004 0.04025
R38052 VDD.n12005 VDD.n340 0.04025
R38053 VDD.n12009 VDD.n340 0.04025
R38054 VDD.n12010 VDD.n12009 0.04025
R38055 VDD.n12011 VDD.n12010 0.04025
R38056 VDD.n12011 VDD.n338 0.04025
R38057 VDD.n12015 VDD.n338 0.04025
R38058 VDD.n12016 VDD.n12015 0.04025
R38059 VDD.n12017 VDD.n12016 0.04025
R38060 VDD.n12017 VDD.n336 0.04025
R38061 VDD.n12021 VDD.n336 0.04025
R38062 VDD.n12022 VDD.n12021 0.04025
R38063 VDD.n12023 VDD.n12022 0.04025
R38064 VDD.n12023 VDD.n334 0.04025
R38065 VDD.n12027 VDD.n334 0.04025
R38066 VDD.n12028 VDD.n12027 0.04025
R38067 VDD.n12029 VDD.n12028 0.04025
R38068 VDD.n12029 VDD.n332 0.04025
R38069 VDD.n12033 VDD.n332 0.04025
R38070 VDD.n12034 VDD.n12033 0.04025
R38071 VDD.n12035 VDD.n12034 0.04025
R38072 VDD.n12035 VDD.n330 0.04025
R38073 VDD.n12039 VDD.n330 0.04025
R38074 VDD.n12040 VDD.n12039 0.04025
R38075 VDD.n12041 VDD.n12040 0.04025
R38076 VDD.n12041 VDD.n328 0.04025
R38077 VDD.n12045 VDD.n328 0.04025
R38078 VDD.n12046 VDD.n12045 0.04025
R38079 VDD.n12047 VDD.n12046 0.04025
R38080 VDD.n12047 VDD.n326 0.04025
R38081 VDD.n12051 VDD.n326 0.04025
R38082 VDD.n12052 VDD.n12051 0.04025
R38083 VDD.n12053 VDD.n12052 0.04025
R38084 VDD.n12053 VDD.n324 0.04025
R38085 VDD.n12057 VDD.n324 0.04025
R38086 VDD.n12058 VDD.n12057 0.04025
R38087 VDD.n12059 VDD.n12058 0.04025
R38088 VDD.n12059 VDD.n322 0.04025
R38089 VDD.n12063 VDD.n322 0.04025
R38090 VDD.n12064 VDD.n12063 0.04025
R38091 VDD.n12065 VDD.n12064 0.04025
R38092 VDD.n12065 VDD.n320 0.04025
R38093 VDD.n12069 VDD.n320 0.04025
R38094 VDD.n12070 VDD.n12069 0.04025
R38095 VDD.n12071 VDD.n12070 0.04025
R38096 VDD.n12071 VDD.n318 0.04025
R38097 VDD.n12075 VDD.n318 0.04025
R38098 VDD.n12076 VDD.n12075 0.04025
R38099 VDD.n12077 VDD.n12076 0.04025
R38100 VDD.n12077 VDD.n316 0.04025
R38101 VDD.n12081 VDD.n316 0.04025
R38102 VDD.n12082 VDD.n12081 0.04025
R38103 VDD.n12083 VDD.n12082 0.04025
R38104 VDD.n12083 VDD.n314 0.04025
R38105 VDD.n12087 VDD.n314 0.04025
R38106 VDD.n12088 VDD.n12087 0.04025
R38107 VDD.n12089 VDD.n12088 0.04025
R38108 VDD.n12089 VDD.n312 0.04025
R38109 VDD.n12093 VDD.n312 0.04025
R38110 VDD.n12094 VDD.n12093 0.04025
R38111 VDD.n12095 VDD.n12094 0.04025
R38112 VDD.n12095 VDD.n310 0.04025
R38113 VDD.n12099 VDD.n310 0.04025
R38114 VDD.n12100 VDD.n12099 0.04025
R38115 VDD.n12101 VDD.n12100 0.04025
R38116 VDD.n12101 VDD.n308 0.04025
R38117 VDD.n12105 VDD.n308 0.04025
R38118 VDD.n12106 VDD.n12105 0.04025
R38119 VDD.n12107 VDD.n12106 0.04025
R38120 VDD.n12107 VDD.n306 0.04025
R38121 VDD.n12111 VDD.n306 0.04025
R38122 VDD.n12112 VDD.n12111 0.04025
R38123 VDD.n12113 VDD.n12112 0.04025
R38124 VDD.n12113 VDD.n304 0.04025
R38125 VDD.n12117 VDD.n304 0.04025
R38126 VDD.n12118 VDD.n12117 0.04025
R38127 VDD.n12119 VDD.n12118 0.04025
R38128 VDD.n12119 VDD.n302 0.04025
R38129 VDD.n12123 VDD.n302 0.04025
R38130 VDD.n12124 VDD.n12123 0.04025
R38131 VDD.n12125 VDD.n12124 0.04025
R38132 VDD.n12125 VDD.n300 0.04025
R38133 VDD.n12129 VDD.n300 0.04025
R38134 VDD.n12130 VDD.n12129 0.04025
R38135 VDD.n12131 VDD.n12130 0.04025
R38136 VDD.n12131 VDD.n298 0.04025
R38137 VDD.n12135 VDD.n298 0.04025
R38138 VDD.n12136 VDD.n12135 0.04025
R38139 VDD.n12137 VDD.n12136 0.04025
R38140 VDD.n12137 VDD.n296 0.04025
R38141 VDD.n12141 VDD.n296 0.04025
R38142 VDD.n12142 VDD.n12141 0.04025
R38143 VDD.n12143 VDD.n12142 0.04025
R38144 VDD.n12143 VDD.n294 0.04025
R38145 VDD.n12147 VDD.n294 0.04025
R38146 VDD.n12148 VDD.n12147 0.04025
R38147 VDD.n12149 VDD.n12148 0.04025
R38148 VDD.n12149 VDD.n292 0.04025
R38149 VDD.n12153 VDD.n292 0.04025
R38150 VDD.n12154 VDD.n12153 0.04025
R38151 VDD.n12155 VDD.n12154 0.04025
R38152 VDD.n12155 VDD.n290 0.04025
R38153 VDD.n12159 VDD.n290 0.04025
R38154 VDD.n12160 VDD.n12159 0.04025
R38155 VDD.n12161 VDD.n12160 0.04025
R38156 VDD.n12161 VDD.n288 0.04025
R38157 VDD.n12165 VDD.n288 0.04025
R38158 VDD.n12166 VDD.n12165 0.04025
R38159 VDD.n12167 VDD.n12166 0.04025
R38160 VDD.n12167 VDD.n286 0.04025
R38161 VDD.n12171 VDD.n286 0.04025
R38162 VDD.n12172 VDD.n12171 0.04025
R38163 VDD.n12173 VDD.n12172 0.04025
R38164 VDD.n12173 VDD.n284 0.04025
R38165 VDD.n12177 VDD.n284 0.04025
R38166 VDD.n12178 VDD.n12177 0.04025
R38167 VDD.n12179 VDD.n12178 0.04025
R38168 VDD.n12179 VDD.n282 0.04025
R38169 VDD.n12183 VDD.n282 0.04025
R38170 VDD.n12184 VDD.n12183 0.04025
R38171 VDD.n12185 VDD.n12184 0.04025
R38172 VDD.n12185 VDD.n280 0.04025
R38173 VDD.n12189 VDD.n280 0.04025
R38174 VDD.n12190 VDD.n12189 0.04025
R38175 VDD.n12191 VDD.n12190 0.04025
R38176 VDD.n12191 VDD.n278 0.04025
R38177 VDD.n12195 VDD.n278 0.04025
R38178 VDD.n12196 VDD.n12195 0.04025
R38179 VDD.n12197 VDD.n12196 0.04025
R38180 VDD.n12197 VDD.n276 0.04025
R38181 VDD.n12201 VDD.n276 0.04025
R38182 VDD.n12202 VDD.n12201 0.04025
R38183 VDD.n12203 VDD.n12202 0.04025
R38184 VDD.n12203 VDD.n274 0.04025
R38185 VDD.n12207 VDD.n274 0.04025
R38186 VDD.n12208 VDD.n12207 0.04025
R38187 VDD.n12209 VDD.n12208 0.04025
R38188 VDD.n12209 VDD.n272 0.04025
R38189 VDD.n12213 VDD.n272 0.04025
R38190 VDD.n12214 VDD.n12213 0.04025
R38191 VDD.n12215 VDD.n12214 0.04025
R38192 VDD.n12215 VDD.n270 0.04025
R38193 VDD.n12219 VDD.n270 0.04025
R38194 VDD.n12220 VDD.n12219 0.04025
R38195 VDD.n12221 VDD.n12220 0.04025
R38196 VDD.n12221 VDD.n268 0.04025
R38197 VDD.n12225 VDD.n268 0.04025
R38198 VDD.n12226 VDD.n12225 0.04025
R38199 VDD.n12227 VDD.n12226 0.04025
R38200 VDD.n12227 VDD.n266 0.04025
R38201 VDD.n12231 VDD.n266 0.04025
R38202 VDD.n12232 VDD.n12231 0.04025
R38203 VDD.n12233 VDD.n12232 0.04025
R38204 VDD.n12233 VDD.n264 0.04025
R38205 VDD.n12237 VDD.n264 0.04025
R38206 VDD.n12238 VDD.n12237 0.04025
R38207 VDD.n12239 VDD.n12238 0.04025
R38208 VDD.n12239 VDD.n262 0.04025
R38209 VDD.n12243 VDD.n262 0.04025
R38210 VDD.n12244 VDD.n12243 0.04025
R38211 VDD.n12245 VDD.n12244 0.04025
R38212 VDD.n12245 VDD.n260 0.04025
R38213 VDD.n12249 VDD.n260 0.04025
R38214 VDD.n12250 VDD.n12249 0.04025
R38215 VDD.n12251 VDD.n12250 0.04025
R38216 VDD.n12251 VDD.n258 0.04025
R38217 VDD.n12255 VDD.n258 0.04025
R38218 VDD.n12256 VDD.n12255 0.04025
R38219 VDD.n12257 VDD.n12256 0.04025
R38220 VDD.n12257 VDD.n256 0.04025
R38221 VDD.n12261 VDD.n256 0.04025
R38222 VDD.n12262 VDD.n12261 0.04025
R38223 VDD.n12263 VDD.n12262 0.04025
R38224 VDD.n12263 VDD.n254 0.04025
R38225 VDD.n12267 VDD.n254 0.04025
R38226 VDD.n12268 VDD.n12267 0.04025
R38227 VDD.n12269 VDD.n12268 0.04025
R38228 VDD.n12269 VDD.n252 0.04025
R38229 VDD.n12273 VDD.n252 0.04025
R38230 VDD.n12274 VDD.n12273 0.04025
R38231 VDD.n12275 VDD.n12274 0.04025
R38232 VDD.n12275 VDD.n250 0.04025
R38233 VDD.n12279 VDD.n250 0.04025
R38234 VDD.n12280 VDD.n12279 0.04025
R38235 VDD.n12281 VDD.n12280 0.04025
R38236 VDD.n12281 VDD.n248 0.04025
R38237 VDD.n12285 VDD.n248 0.04025
R38238 VDD.n12286 VDD.n12285 0.04025
R38239 VDD.n12287 VDD.n12286 0.04025
R38240 VDD.n12287 VDD.n246 0.04025
R38241 VDD.n12291 VDD.n246 0.04025
R38242 VDD.n12292 VDD.n12291 0.04025
R38243 VDD.n12293 VDD.n12292 0.04025
R38244 VDD.n12293 VDD.n244 0.04025
R38245 VDD.n12297 VDD.n244 0.04025
R38246 VDD.n12298 VDD.n12297 0.04025
R38247 VDD.n12299 VDD.n12298 0.04025
R38248 VDD.n12299 VDD.n242 0.04025
R38249 VDD.n12303 VDD.n242 0.04025
R38250 VDD.n12304 VDD.n12303 0.04025
R38251 VDD.n12305 VDD.n12304 0.04025
R38252 VDD.n12305 VDD.n240 0.04025
R38253 VDD.n12309 VDD.n240 0.04025
R38254 VDD.n12310 VDD.n12309 0.04025
R38255 VDD.n12311 VDD.n12310 0.04025
R38256 VDD.n12311 VDD.n238 0.04025
R38257 VDD.n12315 VDD.n238 0.04025
R38258 VDD.n12316 VDD.n12315 0.04025
R38259 VDD.n12317 VDD.n12316 0.04025
R38260 VDD.n12317 VDD.n236 0.04025
R38261 VDD.n12321 VDD.n236 0.04025
R38262 VDD.n12322 VDD.n12321 0.04025
R38263 VDD.n12323 VDD.n12322 0.04025
R38264 VDD.n12323 VDD.n234 0.04025
R38265 VDD.n12327 VDD.n234 0.04025
R38266 VDD.n12328 VDD.n12327 0.04025
R38267 VDD.n12329 VDD.n12328 0.04025
R38268 VDD.n12329 VDD.n232 0.04025
R38269 VDD.n12333 VDD.n232 0.04025
R38270 VDD.n12334 VDD.n12333 0.04025
R38271 VDD.n12335 VDD.n12334 0.04025
R38272 VDD.n12335 VDD.n230 0.04025
R38273 VDD.n12339 VDD.n230 0.04025
R38274 VDD.n12340 VDD.n12339 0.04025
R38275 VDD.n12341 VDD.n12340 0.04025
R38276 VDD.n12341 VDD.n228 0.04025
R38277 VDD.n12345 VDD.n228 0.04025
R38278 VDD.n12346 VDD.n12345 0.04025
R38279 VDD.n12347 VDD.n12346 0.04025
R38280 VDD.n12347 VDD.n226 0.04025
R38281 VDD.n12351 VDD.n226 0.04025
R38282 VDD.n12352 VDD.n12351 0.04025
R38283 VDD.n12353 VDD.n12352 0.04025
R38284 VDD.n12353 VDD.n224 0.04025
R38285 VDD.n12357 VDD.n224 0.04025
R38286 VDD.n12358 VDD.n12357 0.04025
R38287 VDD.n12359 VDD.n12358 0.04025
R38288 VDD.n12359 VDD.n222 0.04025
R38289 VDD.n12363 VDD.n222 0.04025
R38290 VDD.n12364 VDD.n12363 0.04025
R38291 VDD.n12365 VDD.n12364 0.04025
R38292 VDD.n12365 VDD.n220 0.04025
R38293 VDD.n12369 VDD.n220 0.04025
R38294 VDD.n12370 VDD.n12369 0.04025
R38295 VDD.n12371 VDD.n12370 0.04025
R38296 VDD.n12371 VDD.n218 0.04025
R38297 VDD.n12375 VDD.n218 0.04025
R38298 VDD.n12376 VDD.n12375 0.04025
R38299 VDD.n12377 VDD.n12376 0.04025
R38300 VDD.n12377 VDD.n216 0.04025
R38301 VDD.n12381 VDD.n216 0.04025
R38302 VDD.n12382 VDD.n12381 0.04025
R38303 VDD.n12383 VDD.n12382 0.04025
R38304 VDD.n12383 VDD.n214 0.04025
R38305 VDD.n12387 VDD.n214 0.04025
R38306 VDD.n12388 VDD.n12387 0.04025
R38307 VDD.n12389 VDD.n12388 0.04025
R38308 VDD.n12389 VDD.n212 0.04025
R38309 VDD.n12393 VDD.n212 0.04025
R38310 VDD.n12394 VDD.n12393 0.04025
R38311 VDD.n12395 VDD.n12394 0.04025
R38312 VDD.n12395 VDD.n210 0.04025
R38313 VDD.n12399 VDD.n210 0.04025
R38314 VDD.n12400 VDD.n12399 0.04025
R38315 VDD.n12401 VDD.n12400 0.04025
R38316 VDD.n12401 VDD.n208 0.04025
R38317 VDD.n12405 VDD.n208 0.04025
R38318 VDD.n12406 VDD.n12405 0.04025
R38319 VDD.n12407 VDD.n12406 0.04025
R38320 VDD.n12407 VDD.n206 0.04025
R38321 VDD.n12411 VDD.n206 0.04025
R38322 VDD.n12412 VDD.n12411 0.04025
R38323 VDD.n12413 VDD.n12412 0.04025
R38324 VDD.n12413 VDD.n204 0.04025
R38325 VDD.n12417 VDD.n204 0.04025
R38326 VDD.n12418 VDD.n12417 0.04025
R38327 VDD.n12419 VDD.n12418 0.04025
R38328 VDD.n12419 VDD.n202 0.04025
R38329 VDD.n12423 VDD.n202 0.04025
R38330 VDD.n12424 VDD.n12423 0.04025
R38331 VDD.n12425 VDD.n12424 0.04025
R38332 VDD.n12425 VDD.n200 0.04025
R38333 VDD.n12429 VDD.n200 0.04025
R38334 VDD.n12430 VDD.n12429 0.04025
R38335 VDD.n12431 VDD.n12430 0.04025
R38336 VDD.n12431 VDD.n198 0.04025
R38337 VDD.n12435 VDD.n198 0.04025
R38338 VDD.n12436 VDD.n12435 0.04025
R38339 VDD.n12437 VDD.n12436 0.04025
R38340 VDD.n12437 VDD.n196 0.04025
R38341 VDD.n12441 VDD.n196 0.04025
R38342 VDD.n12447 VDD.n12441 0.04025
R38343 VDD.n9437 VDD.n194 0.04025
R38344 VDD.n9438 VDD.n9437 0.04025
R38345 VDD.n9438 VDD.n9435 0.04025
R38346 VDD.n9442 VDD.n9435 0.04025
R38347 VDD.n9443 VDD.n9442 0.04025
R38348 VDD.n9444 VDD.n9443 0.04025
R38349 VDD.n9444 VDD.n9433 0.04025
R38350 VDD.n9448 VDD.n9433 0.04025
R38351 VDD.n9449 VDD.n9448 0.04025
R38352 VDD.n9450 VDD.n9449 0.04025
R38353 VDD.n9450 VDD.n9431 0.04025
R38354 VDD.n9454 VDD.n9431 0.04025
R38355 VDD.n9455 VDD.n9454 0.04025
R38356 VDD.n9456 VDD.n9455 0.04025
R38357 VDD.n9456 VDD.n9429 0.04025
R38358 VDD.n9460 VDD.n9429 0.04025
R38359 VDD.n9461 VDD.n9460 0.04025
R38360 VDD.n9462 VDD.n9461 0.04025
R38361 VDD.n9462 VDD.n9427 0.04025
R38362 VDD.n9466 VDD.n9427 0.04025
R38363 VDD.n9467 VDD.n9466 0.04025
R38364 VDD.n9468 VDD.n9467 0.04025
R38365 VDD.n9468 VDD.n9425 0.04025
R38366 VDD.n9472 VDD.n9425 0.04025
R38367 VDD.n9473 VDD.n9472 0.04025
R38368 VDD.n9474 VDD.n9473 0.04025
R38369 VDD.n9474 VDD.n9423 0.04025
R38370 VDD.n9478 VDD.n9423 0.04025
R38371 VDD.n9479 VDD.n9478 0.04025
R38372 VDD.n9480 VDD.n9479 0.04025
R38373 VDD.n9480 VDD.n9421 0.04025
R38374 VDD.n9484 VDD.n9421 0.04025
R38375 VDD.n9485 VDD.n9484 0.04025
R38376 VDD.n9486 VDD.n9485 0.04025
R38377 VDD.n9486 VDD.n9419 0.04025
R38378 VDD.n9490 VDD.n9419 0.04025
R38379 VDD.n9491 VDD.n9490 0.04025
R38380 VDD.n9492 VDD.n9491 0.04025
R38381 VDD.n9492 VDD.n9417 0.04025
R38382 VDD.n9496 VDD.n9417 0.04025
R38383 VDD.n9497 VDD.n9496 0.04025
R38384 VDD.n9498 VDD.n9497 0.04025
R38385 VDD.n9498 VDD.n9415 0.04025
R38386 VDD.n9502 VDD.n9415 0.04025
R38387 VDD.n9503 VDD.n9502 0.04025
R38388 VDD.n9504 VDD.n9503 0.04025
R38389 VDD.n9504 VDD.n9413 0.04025
R38390 VDD.n9508 VDD.n9413 0.04025
R38391 VDD.n9509 VDD.n9508 0.04025
R38392 VDD.n9510 VDD.n9509 0.04025
R38393 VDD.n9510 VDD.n9411 0.04025
R38394 VDD.n9514 VDD.n9411 0.04025
R38395 VDD.n9515 VDD.n9514 0.04025
R38396 VDD.n9516 VDD.n9515 0.04025
R38397 VDD.n9516 VDD.n9409 0.04025
R38398 VDD.n9520 VDD.n9409 0.04025
R38399 VDD.n9521 VDD.n9520 0.04025
R38400 VDD.n9522 VDD.n9521 0.04025
R38401 VDD.n9522 VDD.n9407 0.04025
R38402 VDD.n9526 VDD.n9407 0.04025
R38403 VDD.n9527 VDD.n9526 0.04025
R38404 VDD.n9528 VDD.n9527 0.04025
R38405 VDD.n9528 VDD.n9405 0.04025
R38406 VDD.n9532 VDD.n9405 0.04025
R38407 VDD.n9533 VDD.n9532 0.04025
R38408 VDD.n9534 VDD.n9533 0.04025
R38409 VDD.n9534 VDD.n9403 0.04025
R38410 VDD.n9538 VDD.n9403 0.04025
R38411 VDD.n9539 VDD.n9538 0.04025
R38412 VDD.n9540 VDD.n9539 0.04025
R38413 VDD.n9540 VDD.n9401 0.04025
R38414 VDD.n9544 VDD.n9401 0.04025
R38415 VDD.n9545 VDD.n9544 0.04025
R38416 VDD.n9546 VDD.n9545 0.04025
R38417 VDD.n9546 VDD.n9399 0.04025
R38418 VDD.n9550 VDD.n9399 0.04025
R38419 VDD.n9551 VDD.n9550 0.04025
R38420 VDD.n9552 VDD.n9551 0.04025
R38421 VDD.n9552 VDD.n9397 0.04025
R38422 VDD.n9556 VDD.n9397 0.04025
R38423 VDD.n9557 VDD.n9556 0.04025
R38424 VDD.n9558 VDD.n9557 0.04025
R38425 VDD.n9558 VDD.n9395 0.04025
R38426 VDD.n9562 VDD.n9395 0.04025
R38427 VDD.n9563 VDD.n9562 0.04025
R38428 VDD.n9564 VDD.n9563 0.04025
R38429 VDD.n9564 VDD.n9393 0.04025
R38430 VDD.n9568 VDD.n9393 0.04025
R38431 VDD.n9569 VDD.n9568 0.04025
R38432 VDD.n9570 VDD.n9569 0.04025
R38433 VDD.n9570 VDD.n9391 0.04025
R38434 VDD.n9574 VDD.n9391 0.04025
R38435 VDD.n9575 VDD.n9574 0.04025
R38436 VDD.n9576 VDD.n9575 0.04025
R38437 VDD.n9576 VDD.n9389 0.04025
R38438 VDD.n9580 VDD.n9389 0.04025
R38439 VDD.n9581 VDD.n9580 0.04025
R38440 VDD.n9582 VDD.n9581 0.04025
R38441 VDD.n9582 VDD.n9387 0.04025
R38442 VDD.n9586 VDD.n9387 0.04025
R38443 VDD.n9587 VDD.n9586 0.04025
R38444 VDD.n9588 VDD.n9587 0.04025
R38445 VDD.n9588 VDD.n9385 0.04025
R38446 VDD.n9592 VDD.n9385 0.04025
R38447 VDD.n9593 VDD.n9592 0.04025
R38448 VDD.n9594 VDD.n9593 0.04025
R38449 VDD.n9594 VDD.n9383 0.04025
R38450 VDD.n9598 VDD.n9383 0.04025
R38451 VDD.n9599 VDD.n9598 0.04025
R38452 VDD.n9600 VDD.n9599 0.04025
R38453 VDD.n9600 VDD.n9381 0.04025
R38454 VDD.n9604 VDD.n9381 0.04025
R38455 VDD.n9605 VDD.n9604 0.04025
R38456 VDD.n9606 VDD.n9605 0.04025
R38457 VDD.n9606 VDD.n9379 0.04025
R38458 VDD.n9610 VDD.n9379 0.04025
R38459 VDD.n9611 VDD.n9610 0.04025
R38460 VDD.n9612 VDD.n9611 0.04025
R38461 VDD.n9612 VDD.n9377 0.04025
R38462 VDD.n9616 VDD.n9377 0.04025
R38463 VDD.n9617 VDD.n9616 0.04025
R38464 VDD.n9618 VDD.n9617 0.04025
R38465 VDD.n9618 VDD.n9375 0.04025
R38466 VDD.n9622 VDD.n9375 0.04025
R38467 VDD.n9623 VDD.n9622 0.04025
R38468 VDD.n9624 VDD.n9623 0.04025
R38469 VDD.n9624 VDD.n9373 0.04025
R38470 VDD.n9628 VDD.n9373 0.04025
R38471 VDD.n9629 VDD.n9628 0.04025
R38472 VDD.n9630 VDD.n9629 0.04025
R38473 VDD.n9630 VDD.n9371 0.04025
R38474 VDD.n9634 VDD.n9371 0.04025
R38475 VDD.n9635 VDD.n9634 0.04025
R38476 VDD.n9636 VDD.n9635 0.04025
R38477 VDD.n9636 VDD.n9369 0.04025
R38478 VDD.n9640 VDD.n9369 0.04025
R38479 VDD.n9641 VDD.n9640 0.04025
R38480 VDD.n9642 VDD.n9641 0.04025
R38481 VDD.n9642 VDD.n9367 0.04025
R38482 VDD.n9646 VDD.n9367 0.04025
R38483 VDD.n9647 VDD.n9646 0.04025
R38484 VDD.n9648 VDD.n9647 0.04025
R38485 VDD.n9648 VDD.n9365 0.04025
R38486 VDD.n9652 VDD.n9365 0.04025
R38487 VDD.n9653 VDD.n9652 0.04025
R38488 VDD.n9654 VDD.n9653 0.04025
R38489 VDD.n9654 VDD.n9363 0.04025
R38490 VDD.n9658 VDD.n9363 0.04025
R38491 VDD.n9659 VDD.n9658 0.04025
R38492 VDD.n9660 VDD.n9659 0.04025
R38493 VDD.n9660 VDD.n9361 0.04025
R38494 VDD.n9664 VDD.n9361 0.04025
R38495 VDD.n9665 VDD.n9664 0.04025
R38496 VDD.n9666 VDD.n9665 0.04025
R38497 VDD.n9666 VDD.n9359 0.04025
R38498 VDD.n9670 VDD.n9359 0.04025
R38499 VDD.n9671 VDD.n9670 0.04025
R38500 VDD.n9672 VDD.n9671 0.04025
R38501 VDD.n9672 VDD.n9357 0.04025
R38502 VDD.n9676 VDD.n9357 0.04025
R38503 VDD.n9677 VDD.n9676 0.04025
R38504 VDD.n9678 VDD.n9677 0.04025
R38505 VDD.n9678 VDD.n9355 0.04025
R38506 VDD.n9682 VDD.n9355 0.04025
R38507 VDD.n9683 VDD.n9682 0.04025
R38508 VDD.n9684 VDD.n9683 0.04025
R38509 VDD.n9684 VDD.n9353 0.04025
R38510 VDD.n9688 VDD.n9353 0.04025
R38511 VDD.n9689 VDD.n9688 0.04025
R38512 VDD.n9690 VDD.n9689 0.04025
R38513 VDD.n9690 VDD.n9351 0.04025
R38514 VDD.n9694 VDD.n9351 0.04025
R38515 VDD.n9695 VDD.n9694 0.04025
R38516 VDD.n9696 VDD.n9695 0.04025
R38517 VDD.n9696 VDD.n9349 0.04025
R38518 VDD.n9700 VDD.n9349 0.04025
R38519 VDD.n9701 VDD.n9700 0.04025
R38520 VDD.n9702 VDD.n9701 0.04025
R38521 VDD.n9702 VDD.n9347 0.04025
R38522 VDD.n9706 VDD.n9347 0.04025
R38523 VDD.n9707 VDD.n9706 0.04025
R38524 VDD.n9708 VDD.n9707 0.04025
R38525 VDD.n9708 VDD.n9345 0.04025
R38526 VDD.n9712 VDD.n9345 0.04025
R38527 VDD.n9713 VDD.n9712 0.04025
R38528 VDD.n9714 VDD.n9713 0.04025
R38529 VDD.n9714 VDD.n9343 0.04025
R38530 VDD.n9718 VDD.n9343 0.04025
R38531 VDD.n9719 VDD.n9718 0.04025
R38532 VDD.n9720 VDD.n9719 0.04025
R38533 VDD.n9720 VDD.n9341 0.04025
R38534 VDD.n9724 VDD.n9341 0.04025
R38535 VDD.n9725 VDD.n9724 0.04025
R38536 VDD.n9726 VDD.n9725 0.04025
R38537 VDD.n9726 VDD.n9339 0.04025
R38538 VDD.n9730 VDD.n9339 0.04025
R38539 VDD.n9731 VDD.n9730 0.04025
R38540 VDD.n9732 VDD.n9731 0.04025
R38541 VDD.n9732 VDD.n9337 0.04025
R38542 VDD.n9736 VDD.n9337 0.04025
R38543 VDD.n9737 VDD.n9736 0.04025
R38544 VDD.n9738 VDD.n9737 0.04025
R38545 VDD.n9738 VDD.n9335 0.04025
R38546 VDD.n9742 VDD.n9335 0.04025
R38547 VDD.n9743 VDD.n9742 0.04025
R38548 VDD.n9744 VDD.n9743 0.04025
R38549 VDD.n9744 VDD.n9333 0.04025
R38550 VDD.n9748 VDD.n9333 0.04025
R38551 VDD.n9749 VDD.n9748 0.04025
R38552 VDD.n9750 VDD.n9749 0.04025
R38553 VDD.n9750 VDD.n9331 0.04025
R38554 VDD.n9754 VDD.n9331 0.04025
R38555 VDD.n9755 VDD.n9754 0.04025
R38556 VDD.n9756 VDD.n9755 0.04025
R38557 VDD.n9756 VDD.n9329 0.04025
R38558 VDD.n9760 VDD.n9329 0.04025
R38559 VDD.n9761 VDD.n9760 0.04025
R38560 VDD.n9762 VDD.n9761 0.04025
R38561 VDD.n9762 VDD.n9327 0.04025
R38562 VDD.n9766 VDD.n9327 0.04025
R38563 VDD.n9767 VDD.n9766 0.04025
R38564 VDD.n9768 VDD.n9767 0.04025
R38565 VDD.n9768 VDD.n9325 0.04025
R38566 VDD.n9772 VDD.n9325 0.04025
R38567 VDD.n9773 VDD.n9772 0.04025
R38568 VDD.n9774 VDD.n9773 0.04025
R38569 VDD.n9774 VDD.n9323 0.04025
R38570 VDD.n9778 VDD.n9323 0.04025
R38571 VDD.n9779 VDD.n9778 0.04025
R38572 VDD.n9780 VDD.n9779 0.04025
R38573 VDD.n9780 VDD.n9321 0.04025
R38574 VDD.n9784 VDD.n9321 0.04025
R38575 VDD.n9785 VDD.n9784 0.04025
R38576 VDD.n9786 VDD.n9785 0.04025
R38577 VDD.n9786 VDD.n9319 0.04025
R38578 VDD.n9790 VDD.n9319 0.04025
R38579 VDD.n9791 VDD.n9790 0.04025
R38580 VDD.n9792 VDD.n9791 0.04025
R38581 VDD.n9792 VDD.n9317 0.04025
R38582 VDD.n9796 VDD.n9317 0.04025
R38583 VDD.n9797 VDD.n9796 0.04025
R38584 VDD.n9798 VDD.n9797 0.04025
R38585 VDD.n9798 VDD.n9315 0.04025
R38586 VDD.n9802 VDD.n9315 0.04025
R38587 VDD.n9803 VDD.n9802 0.04025
R38588 VDD.n9804 VDD.n9803 0.04025
R38589 VDD.n9804 VDD.n9313 0.04025
R38590 VDD.n9808 VDD.n9313 0.04025
R38591 VDD.n9809 VDD.n9808 0.04025
R38592 VDD.n9810 VDD.n9809 0.04025
R38593 VDD.n9810 VDD.n9311 0.04025
R38594 VDD.n9814 VDD.n9311 0.04025
R38595 VDD.n9815 VDD.n9814 0.04025
R38596 VDD.n9816 VDD.n9815 0.04025
R38597 VDD.n9816 VDD.n9309 0.04025
R38598 VDD.n9820 VDD.n9309 0.04025
R38599 VDD.n9821 VDD.n9820 0.04025
R38600 VDD.n9822 VDD.n9821 0.04025
R38601 VDD.n9822 VDD.n9307 0.04025
R38602 VDD.n9826 VDD.n9307 0.04025
R38603 VDD.n9827 VDD.n9826 0.04025
R38604 VDD.n9828 VDD.n9827 0.04025
R38605 VDD.n9828 VDD.n9305 0.04025
R38606 VDD.n9832 VDD.n9305 0.04025
R38607 VDD.n9833 VDD.n9832 0.04025
R38608 VDD.n9834 VDD.n9833 0.04025
R38609 VDD.n9834 VDD.n9303 0.04025
R38610 VDD.n9838 VDD.n9303 0.04025
R38611 VDD.n9839 VDD.n9838 0.04025
R38612 VDD.n9840 VDD.n9839 0.04025
R38613 VDD.n9840 VDD.n9301 0.04025
R38614 VDD.n9844 VDD.n9301 0.04025
R38615 VDD.n9845 VDD.n9844 0.04025
R38616 VDD.n9846 VDD.n9845 0.04025
R38617 VDD.n9846 VDD.n9299 0.04025
R38618 VDD.n9850 VDD.n9299 0.04025
R38619 VDD.n9851 VDD.n9850 0.04025
R38620 VDD.n9852 VDD.n9851 0.04025
R38621 VDD.n9852 VDD.n9297 0.04025
R38622 VDD.n9856 VDD.n9297 0.04025
R38623 VDD.n9857 VDD.n9856 0.04025
R38624 VDD.n9858 VDD.n9857 0.04025
R38625 VDD.n9858 VDD.n9295 0.04025
R38626 VDD.n9862 VDD.n9295 0.04025
R38627 VDD.n9863 VDD.n9862 0.04025
R38628 VDD.n9864 VDD.n9863 0.04025
R38629 VDD.n9864 VDD.n9293 0.04025
R38630 VDD.n9868 VDD.n9293 0.04025
R38631 VDD.n9869 VDD.n9868 0.04025
R38632 VDD.n9870 VDD.n9869 0.04025
R38633 VDD.n9870 VDD.n9291 0.04025
R38634 VDD.n9874 VDD.n9291 0.04025
R38635 VDD.n9875 VDD.n9874 0.04025
R38636 VDD.n9876 VDD.n9875 0.04025
R38637 VDD.n9876 VDD.n9289 0.04025
R38638 VDD.n9880 VDD.n9289 0.04025
R38639 VDD.n9881 VDD.n9880 0.04025
R38640 VDD.n9882 VDD.n9881 0.04025
R38641 VDD.n9882 VDD.n9287 0.04025
R38642 VDD.n9886 VDD.n9287 0.04025
R38643 VDD.n9887 VDD.n9886 0.04025
R38644 VDD.n9888 VDD.n9887 0.04025
R38645 VDD.n9888 VDD.n9285 0.04025
R38646 VDD.n9892 VDD.n9285 0.04025
R38647 VDD.n9893 VDD.n9892 0.04025
R38648 VDD.n9894 VDD.n9893 0.04025
R38649 VDD.n9894 VDD.n9283 0.04025
R38650 VDD.n9898 VDD.n9283 0.04025
R38651 VDD.n9899 VDD.n9898 0.04025
R38652 VDD.n9900 VDD.n9899 0.04025
R38653 VDD.n9900 VDD.n9281 0.04025
R38654 VDD.n9904 VDD.n9281 0.04025
R38655 VDD.n9905 VDD.n9904 0.04025
R38656 VDD.n9906 VDD.n9905 0.04025
R38657 VDD.n9906 VDD.n9279 0.04025
R38658 VDD.n9910 VDD.n9279 0.04025
R38659 VDD.n9911 VDD.n9910 0.04025
R38660 VDD.n9912 VDD.n9911 0.04025
R38661 VDD.n9912 VDD.n9277 0.04025
R38662 VDD.n9916 VDD.n9277 0.04025
R38663 VDD.n9917 VDD.n9916 0.04025
R38664 VDD.n9918 VDD.n9917 0.04025
R38665 VDD.n9918 VDD.n9275 0.04025
R38666 VDD.n9922 VDD.n9275 0.04025
R38667 VDD.n9923 VDD.n9922 0.04025
R38668 VDD.n9924 VDD.n9923 0.04025
R38669 VDD.n9924 VDD.n9273 0.04025
R38670 VDD.n9928 VDD.n9273 0.04025
R38671 VDD.n9929 VDD.n9928 0.04025
R38672 VDD.n9930 VDD.n9929 0.04025
R38673 VDD.n9930 VDD.n9271 0.04025
R38674 VDD.n9934 VDD.n9271 0.04025
R38675 VDD.n9935 VDD.n9934 0.04025
R38676 VDD.n9936 VDD.n9935 0.04025
R38677 VDD.n9936 VDD.n9269 0.04025
R38678 VDD.n9940 VDD.n9269 0.04025
R38679 VDD.n9941 VDD.n9940 0.04025
R38680 VDD.n9942 VDD.n9941 0.04025
R38681 VDD.n9942 VDD.n9267 0.04025
R38682 VDD.n9946 VDD.n9267 0.04025
R38683 VDD.n9947 VDD.n9946 0.04025
R38684 VDD.n9948 VDD.n9947 0.04025
R38685 VDD.n9948 VDD.n9265 0.04025
R38686 VDD.n9952 VDD.n9265 0.04025
R38687 VDD.n9953 VDD.n9952 0.04025
R38688 VDD.n9954 VDD.n9953 0.04025
R38689 VDD.n9954 VDD.n9263 0.04025
R38690 VDD.n9958 VDD.n9263 0.04025
R38691 VDD.n9959 VDD.n9958 0.04025
R38692 VDD.n9960 VDD.n9959 0.04025
R38693 VDD.n9960 VDD.n9261 0.04025
R38694 VDD.n9964 VDD.n9261 0.04025
R38695 VDD.n9965 VDD.n9964 0.04025
R38696 VDD.n9966 VDD.n9965 0.04025
R38697 VDD.n9966 VDD.n9259 0.04025
R38698 VDD.n9970 VDD.n9259 0.04025
R38699 VDD.n9971 VDD.n9970 0.04025
R38700 VDD.n9972 VDD.n9971 0.04025
R38701 VDD.n9972 VDD.n9257 0.04025
R38702 VDD.n9976 VDD.n9257 0.04025
R38703 VDD.n9977 VDD.n9976 0.04025
R38704 VDD.n9978 VDD.n9977 0.04025
R38705 VDD.n9978 VDD.n9255 0.04025
R38706 VDD.n9982 VDD.n9255 0.04025
R38707 VDD.n9983 VDD.n9982 0.04025
R38708 VDD.n9984 VDD.n9983 0.04025
R38709 VDD.n9984 VDD.n9253 0.04025
R38710 VDD.n9988 VDD.n9253 0.04025
R38711 VDD.n9989 VDD.n9988 0.04025
R38712 VDD.n9990 VDD.n9989 0.04025
R38713 VDD.n9990 VDD.n9251 0.04025
R38714 VDD.n9994 VDD.n9251 0.04025
R38715 VDD.n9995 VDD.n9994 0.04025
R38716 VDD.n9996 VDD.n9995 0.04025
R38717 VDD.n9996 VDD.n9249 0.04025
R38718 VDD.n10000 VDD.n9249 0.04025
R38719 VDD.n10001 VDD.n10000 0.04025
R38720 VDD.n10002 VDD.n10001 0.04025
R38721 VDD.n10002 VDD.n9247 0.04025
R38722 VDD.n10006 VDD.n9247 0.04025
R38723 VDD.n10007 VDD.n10006 0.04025
R38724 VDD.n10008 VDD.n10007 0.04025
R38725 VDD.n10008 VDD.n9245 0.04025
R38726 VDD.n10012 VDD.n9245 0.04025
R38727 VDD.n10013 VDD.n10012 0.04025
R38728 VDD.n10014 VDD.n10013 0.04025
R38729 VDD.n10014 VDD.n9243 0.04025
R38730 VDD.n10018 VDD.n9243 0.04025
R38731 VDD.n10019 VDD.n10018 0.04025
R38732 VDD.n10020 VDD.n10019 0.04025
R38733 VDD.n10020 VDD.n9241 0.04025
R38734 VDD.n10024 VDD.n9241 0.04025
R38735 VDD.n10025 VDD.n10024 0.04025
R38736 VDD.n10026 VDD.n10025 0.04025
R38737 VDD.n10026 VDD.n9239 0.04025
R38738 VDD.n10030 VDD.n9239 0.04025
R38739 VDD.n10031 VDD.n10030 0.04025
R38740 VDD.n10032 VDD.n10031 0.04025
R38741 VDD.n10032 VDD.n9237 0.04025
R38742 VDD.n10036 VDD.n9237 0.04025
R38743 VDD.n10037 VDD.n10036 0.04025
R38744 VDD.n10038 VDD.n10037 0.04025
R38745 VDD.n10038 VDD.n9235 0.04025
R38746 VDD.n10042 VDD.n9235 0.04025
R38747 VDD.n10043 VDD.n10042 0.04025
R38748 VDD.n10044 VDD.n10043 0.04025
R38749 VDD.n10044 VDD.n9233 0.04025
R38750 VDD.n10048 VDD.n9233 0.04025
R38751 VDD.n10049 VDD.n10048 0.04025
R38752 VDD.n10050 VDD.n10049 0.04025
R38753 VDD.n10050 VDD.n9231 0.04025
R38754 VDD.n10054 VDD.n9231 0.04025
R38755 VDD.n10055 VDD.n10054 0.04025
R38756 VDD.n10056 VDD.n10055 0.04025
R38757 VDD.n10056 VDD.n9229 0.04025
R38758 VDD.n10060 VDD.n9229 0.04025
R38759 VDD.n10061 VDD.n10060 0.04025
R38760 VDD.n10062 VDD.n10061 0.04025
R38761 VDD.n10062 VDD.n9227 0.04025
R38762 VDD.n10066 VDD.n9227 0.04025
R38763 VDD.n10067 VDD.n10066 0.04025
R38764 VDD.n10068 VDD.n10067 0.04025
R38765 VDD.n10068 VDD.n9225 0.04025
R38766 VDD.n10072 VDD.n9225 0.04025
R38767 VDD.n10073 VDD.n10072 0.04025
R38768 VDD.n10074 VDD.n10073 0.04025
R38769 VDD.n10074 VDD.n9223 0.04025
R38770 VDD.n10078 VDD.n9223 0.04025
R38771 VDD.n10079 VDD.n10078 0.04025
R38772 VDD.n10080 VDD.n10079 0.04025
R38773 VDD.n10080 VDD.n9221 0.04025
R38774 VDD.n10084 VDD.n9221 0.04025
R38775 VDD.n10085 VDD.n10084 0.04025
R38776 VDD.n10086 VDD.n10085 0.04025
R38777 VDD.n10086 VDD.n9219 0.04025
R38778 VDD.n10090 VDD.n9219 0.04025
R38779 VDD.n10091 VDD.n10090 0.04025
R38780 VDD.n10092 VDD.n10091 0.04025
R38781 VDD.n10092 VDD.n9217 0.04025
R38782 VDD.n10096 VDD.n9217 0.04025
R38783 VDD.n10097 VDD.n10096 0.04025
R38784 VDD.n10098 VDD.n10097 0.04025
R38785 VDD.n10098 VDD.n9215 0.04025
R38786 VDD.n10102 VDD.n9215 0.04025
R38787 VDD.n4904 VDD.n4903 0.04025
R38788 VDD.n4903 VDD.n4698 0.04025
R38789 VDD.n4899 VDD.n4698 0.04025
R38790 VDD.n4899 VDD.n4898 0.04025
R38791 VDD.n4898 VDD.n4897 0.04025
R38792 VDD.n4897 VDD.n4700 0.04025
R38793 VDD.n4893 VDD.n4700 0.04025
R38794 VDD.n4893 VDD.n4892 0.04025
R38795 VDD.n4892 VDD.n4891 0.04025
R38796 VDD.n4891 VDD.n4702 0.04025
R38797 VDD.n4887 VDD.n4702 0.04025
R38798 VDD.n4887 VDD.n4886 0.04025
R38799 VDD.n4886 VDD.n4885 0.04025
R38800 VDD.n4885 VDD.n4704 0.04025
R38801 VDD.n4881 VDD.n4704 0.04025
R38802 VDD.n4881 VDD.n4880 0.04025
R38803 VDD.n4880 VDD.n4879 0.04025
R38804 VDD.n4879 VDD.n4706 0.04025
R38805 VDD.n4875 VDD.n4706 0.04025
R38806 VDD.n4875 VDD.n4874 0.04025
R38807 VDD.n4874 VDD.n4873 0.04025
R38808 VDD.n4873 VDD.n4708 0.04025
R38809 VDD.n4869 VDD.n4708 0.04025
R38810 VDD.n4869 VDD.n4868 0.04025
R38811 VDD.n4868 VDD.n4867 0.04025
R38812 VDD.n4867 VDD.n4710 0.04025
R38813 VDD.n4863 VDD.n4710 0.04025
R38814 VDD.n4863 VDD.n4862 0.04025
R38815 VDD.n4862 VDD.n4861 0.04025
R38816 VDD.n4861 VDD.n4712 0.04025
R38817 VDD.n4857 VDD.n4712 0.04025
R38818 VDD.n4857 VDD.n4856 0.04025
R38819 VDD.n4856 VDD.n4855 0.04025
R38820 VDD.n4855 VDD.n4714 0.04025
R38821 VDD.n4851 VDD.n4714 0.04025
R38822 VDD.n4851 VDD.n4850 0.04025
R38823 VDD.n4850 VDD.n4849 0.04025
R38824 VDD.n4849 VDD.n4716 0.04025
R38825 VDD.n4845 VDD.n4716 0.04025
R38826 VDD.n4845 VDD.n4844 0.04025
R38827 VDD.n4844 VDD.n4843 0.04025
R38828 VDD.n4843 VDD.n4718 0.04025
R38829 VDD.n4839 VDD.n4718 0.04025
R38830 VDD.n4839 VDD.n4838 0.04025
R38831 VDD.n4838 VDD.n4837 0.04025
R38832 VDD.n4837 VDD.n4720 0.04025
R38833 VDD.n4833 VDD.n4720 0.04025
R38834 VDD.n4833 VDD.n4832 0.04025
R38835 VDD.n4832 VDD.n4831 0.04025
R38836 VDD.n4831 VDD.n4722 0.04025
R38837 VDD.n4827 VDD.n4722 0.04025
R38838 VDD.n4827 VDD.n4826 0.04025
R38839 VDD.n4826 VDD.n4825 0.04025
R38840 VDD.n4825 VDD.n4724 0.04025
R38841 VDD.n4821 VDD.n4724 0.04025
R38842 VDD.n4821 VDD.n4820 0.04025
R38843 VDD.n4820 VDD.n4819 0.04025
R38844 VDD.n4819 VDD.n4726 0.04025
R38845 VDD.n4815 VDD.n4726 0.04025
R38846 VDD.n4815 VDD.n4814 0.04025
R38847 VDD.n4814 VDD.n4813 0.04025
R38848 VDD.n4813 VDD.n4728 0.04025
R38849 VDD.n4809 VDD.n4728 0.04025
R38850 VDD.n4809 VDD.n4808 0.04025
R38851 VDD.n4808 VDD.n4807 0.04025
R38852 VDD.n4807 VDD.n4730 0.04025
R38853 VDD.n4803 VDD.n4730 0.04025
R38854 VDD.n4803 VDD.n4802 0.04025
R38855 VDD.n4802 VDD.n4801 0.04025
R38856 VDD.n4801 VDD.n4732 0.04025
R38857 VDD.n4797 VDD.n4732 0.04025
R38858 VDD.n4797 VDD.n4796 0.04025
R38859 VDD.n4796 VDD.n4795 0.04025
R38860 VDD.n4795 VDD.n4734 0.04025
R38861 VDD.n4791 VDD.n4734 0.04025
R38862 VDD.n4791 VDD.n4790 0.04025
R38863 VDD.n4790 VDD.n4789 0.04025
R38864 VDD.n4789 VDD.n4736 0.04025
R38865 VDD.n4785 VDD.n4736 0.04025
R38866 VDD.n4785 VDD.n4784 0.04025
R38867 VDD.n4784 VDD.n4783 0.04025
R38868 VDD.n4783 VDD.n4738 0.04025
R38869 VDD.n4779 VDD.n4738 0.04025
R38870 VDD.n4779 VDD.n4778 0.04025
R38871 VDD.n4778 VDD.n4777 0.04025
R38872 VDD.n4777 VDD.n4740 0.04025
R38873 VDD.n4773 VDD.n4740 0.04025
R38874 VDD.n4773 VDD.n4772 0.04025
R38875 VDD.n4772 VDD.n4771 0.04025
R38876 VDD.n4771 VDD.n4742 0.04025
R38877 VDD.n4767 VDD.n4742 0.04025
R38878 VDD.n4767 VDD.n4766 0.04025
R38879 VDD.n4766 VDD.n4765 0.04025
R38880 VDD.n4765 VDD.n4744 0.04025
R38881 VDD.n4761 VDD.n4744 0.04025
R38882 VDD.n4761 VDD.n4760 0.04025
R38883 VDD.n4760 VDD.n4759 0.04025
R38884 VDD.n4759 VDD.n4746 0.04025
R38885 VDD.n4755 VDD.n4746 0.04025
R38886 VDD.n4755 VDD.n4754 0.04025
R38887 VDD.n4754 VDD.n4753 0.04025
R38888 VDD.n4753 VDD.n4748 0.04025
R38889 VDD.n4749 VDD.n4748 0.04025
R38890 VDD.n4749 VDD.n2244 0.04025
R38891 VDD.n7819 VDD.n2244 0.04025
R38892 VDD.n7819 VDD.n7818 0.04025
R38893 VDD.n7818 VDD.n7817 0.04025
R38894 VDD.n7817 VDD.n2245 0.04025
R38895 VDD.n7813 VDD.n2245 0.04025
R38896 VDD.n7813 VDD.n7812 0.04025
R38897 VDD.n7812 VDD.n7811 0.04025
R38898 VDD.n7811 VDD.n2247 0.04025
R38899 VDD.n7806 VDD.n2247 0.04025
R38900 VDD.n7806 VDD.n7805 0.04025
R38901 VDD.n7805 VDD.n7804 0.04025
R38902 VDD.n7804 VDD.n2249 0.04025
R38903 VDD.n7800 VDD.n2249 0.04025
R38904 VDD.n7800 VDD.n7799 0.04025
R38905 VDD.n7799 VDD.n2251 0.04025
R38906 VDD.n7795 VDD.n2251 0.04025
R38907 VDD.n7795 VDD.n7794 0.04025
R38908 VDD.n7794 VDD.n2253 0.04025
R38909 VDD.n7790 VDD.n2253 0.04025
R38910 VDD.n7790 VDD.n7789 0.04025
R38911 VDD.n7789 VDD.n7788 0.04025
R38912 VDD.n7788 VDD.n2255 0.04025
R38913 VDD.n7784 VDD.n2255 0.04025
R38914 VDD.n7784 VDD.n7783 0.04025
R38915 VDD.n7783 VDD.n7782 0.04025
R38916 VDD.n7782 VDD.n2257 0.04025
R38917 VDD.n7777 VDD.n2257 0.04025
R38918 VDD.n7777 VDD.n7776 0.04025
R38919 VDD.n7776 VDD.n7775 0.04025
R38920 VDD.n7775 VDD.n2259 0.04025
R38921 VDD.n7771 VDD.n2259 0.04025
R38922 VDD.n7771 VDD.n7770 0.04025
R38923 VDD.n7770 VDD.n7769 0.04025
R38924 VDD.n7769 VDD.n2262 0.04025
R38925 VDD.n7765 VDD.n2262 0.04025
R38926 VDD.n7765 VDD.n7764 0.04025
R38927 VDD.n7764 VDD.n7763 0.04025
R38928 VDD.n7763 VDD.n2264 0.04025
R38929 VDD.n7758 VDD.n2264 0.04025
R38930 VDD.n7758 VDD.n7757 0.04025
R38931 VDD.n7757 VDD.n7756 0.04025
R38932 VDD.n7756 VDD.n2267 0.04025
R38933 VDD.n7752 VDD.n2267 0.04025
R38934 VDD.n7752 VDD.n7751 0.04025
R38935 VDD.n7751 VDD.n7750 0.04025
R38936 VDD.n7750 VDD.n2269 0.04025
R38937 VDD.n7746 VDD.n2269 0.04025
R38938 VDD.n7746 VDD.n7745 0.04025
R38939 VDD.n7745 VDD.n2271 0.04025
R38940 VDD.n7741 VDD.n2271 0.04025
R38941 VDD.n7741 VDD.n7740 0.04025
R38942 VDD.n7740 VDD.n2273 0.04025
R38943 VDD.n7736 VDD.n2273 0.04025
R38944 VDD.n7736 VDD.n7735 0.04025
R38945 VDD.n7735 VDD.n7734 0.04025
R38946 VDD.n7734 VDD.n2275 0.04025
R38947 VDD.n7730 VDD.n2275 0.04025
R38948 VDD.n7730 VDD.n7729 0.04025
R38949 VDD.n7729 VDD.n7728 0.04025
R38950 VDD.n7728 VDD.n2277 0.04025
R38951 VDD.n7723 VDD.n2277 0.04025
R38952 VDD.n7723 VDD.n7722 0.04025
R38953 VDD.n7722 VDD.n7721 0.04025
R38954 VDD.n7721 VDD.n2279 0.04025
R38955 VDD.n7716 VDD.n2279 0.04025
R38956 VDD.n7716 VDD.n7715 0.04025
R38957 VDD.n7715 VDD.n7714 0.04025
R38958 VDD.n7714 VDD.n2281 0.04025
R38959 VDD.n7710 VDD.n2281 0.04025
R38960 VDD.n7710 VDD.n7709 0.04025
R38961 VDD.n7709 VDD.n2284 0.04025
R38962 VDD.n7705 VDD.n2284 0.04025
R38963 VDD.n7705 VDD.n7704 0.04025
R38964 VDD.n7704 VDD.n7703 0.04025
R38965 VDD.n7703 VDD.n2286 0.04025
R38966 VDD.n7698 VDD.n2286 0.04025
R38967 VDD.n7698 VDD.n7697 0.04025
R38968 VDD.n7697 VDD.n7696 0.04025
R38969 VDD.n7696 VDD.n2288 0.04025
R38970 VDD.n7692 VDD.n2288 0.04025
R38971 VDD.n7692 VDD.n7691 0.04025
R38972 VDD.n7691 VDD.n7690 0.04025
R38973 VDD.n7690 VDD.n2290 0.04025
R38974 VDD.n7686 VDD.n2290 0.04025
R38975 VDD.n7686 VDD.n7685 0.04025
R38976 VDD.n7685 VDD.n2293 0.04025
R38977 VDD.n7680 VDD.n2293 0.04025
R38978 VDD.n7680 VDD.n7679 0.04025
R38979 VDD.n7679 VDD.n7678 0.04025
R38980 VDD.n7678 VDD.n7179 0.04025
R38981 VDD.n7674 VDD.n7179 0.04025
R38982 VDD.n7674 VDD.n7673 0.04025
R38983 VDD.n7673 VDD.n7672 0.04025
R38984 VDD.n7672 VDD.n7181 0.04025
R38985 VDD.n7668 VDD.n7181 0.04025
R38986 VDD.n7668 VDD.n7667 0.04025
R38987 VDD.n7667 VDD.n7666 0.04025
R38988 VDD.n7666 VDD.n7183 0.04025
R38989 VDD.n7662 VDD.n7183 0.04025
R38990 VDD.n7662 VDD.n7661 0.04025
R38991 VDD.n7661 VDD.n7660 0.04025
R38992 VDD.n7660 VDD.n7185 0.04025
R38993 VDD.n7656 VDD.n7185 0.04025
R38994 VDD.n7656 VDD.n7655 0.04025
R38995 VDD.n7655 VDD.n7654 0.04025
R38996 VDD.n7654 VDD.n7187 0.04025
R38997 VDD.n7650 VDD.n7187 0.04025
R38998 VDD.n7650 VDD.n7649 0.04025
R38999 VDD.n7649 VDD.n7648 0.04025
R39000 VDD.n7648 VDD.n7189 0.04025
R39001 VDD.n7644 VDD.n7189 0.04025
R39002 VDD.n7644 VDD.n7643 0.04025
R39003 VDD.n7643 VDD.n7642 0.04025
R39004 VDD.n7642 VDD.n7191 0.04025
R39005 VDD.n7638 VDD.n7191 0.04025
R39006 VDD.n7638 VDD.n7637 0.04025
R39007 VDD.n7637 VDD.n7636 0.04025
R39008 VDD.n7636 VDD.n7193 0.04025
R39009 VDD.n7632 VDD.n7193 0.04025
R39010 VDD.n7632 VDD.n7631 0.04025
R39011 VDD.n7631 VDD.n7630 0.04025
R39012 VDD.n7630 VDD.n7195 0.04025
R39013 VDD.n7626 VDD.n7195 0.04025
R39014 VDD.n7626 VDD.n7625 0.04025
R39015 VDD.n7625 VDD.n7624 0.04025
R39016 VDD.n7624 VDD.n7197 0.04025
R39017 VDD.n7620 VDD.n7197 0.04025
R39018 VDD.n7620 VDD.n7619 0.04025
R39019 VDD.n7619 VDD.n7618 0.04025
R39020 VDD.n7618 VDD.n7199 0.04025
R39021 VDD.n7614 VDD.n7199 0.04025
R39022 VDD.n7614 VDD.n7613 0.04025
R39023 VDD.n7613 VDD.n7612 0.04025
R39024 VDD.n7612 VDD.n7201 0.04025
R39025 VDD.n7608 VDD.n7201 0.04025
R39026 VDD.n7608 VDD.n7607 0.04025
R39027 VDD.n7607 VDD.n7606 0.04025
R39028 VDD.n7606 VDD.n7203 0.04025
R39029 VDD.n7602 VDD.n7203 0.04025
R39030 VDD.n7602 VDD.n7601 0.04025
R39031 VDD.n7601 VDD.n7600 0.04025
R39032 VDD.n7600 VDD.n7205 0.04025
R39033 VDD.n7596 VDD.n7205 0.04025
R39034 VDD.n7596 VDD.n7595 0.04025
R39035 VDD.n7595 VDD.n7594 0.04025
R39036 VDD.n7594 VDD.n7207 0.04025
R39037 VDD.n7590 VDD.n7207 0.04025
R39038 VDD.n7590 VDD.n7589 0.04025
R39039 VDD.n7589 VDD.n7588 0.04025
R39040 VDD.n7588 VDD.n7209 0.04025
R39041 VDD.n7584 VDD.n7209 0.04025
R39042 VDD.n7584 VDD.n7583 0.04025
R39043 VDD.n7583 VDD.n7582 0.04025
R39044 VDD.n7582 VDD.n7211 0.04025
R39045 VDD.n7578 VDD.n7211 0.04025
R39046 VDD.n7578 VDD.n7577 0.04025
R39047 VDD.n7577 VDD.n7576 0.04025
R39048 VDD.n7576 VDD.n7213 0.04025
R39049 VDD.n7572 VDD.n7213 0.04025
R39050 VDD.n7572 VDD.n7571 0.04025
R39051 VDD.n7571 VDD.n7570 0.04025
R39052 VDD.n7570 VDD.n7215 0.04025
R39053 VDD.n7566 VDD.n7215 0.04025
R39054 VDD.n7566 VDD.n7565 0.04025
R39055 VDD.n7565 VDD.n7564 0.04025
R39056 VDD.n7564 VDD.n7217 0.04025
R39057 VDD.n7560 VDD.n7217 0.04025
R39058 VDD.n7560 VDD.n7559 0.04025
R39059 VDD.n7559 VDD.n7558 0.04025
R39060 VDD.n7558 VDD.n7219 0.04025
R39061 VDD.n7554 VDD.n7219 0.04025
R39062 VDD.n7554 VDD.n7553 0.04025
R39063 VDD.n7553 VDD.n7552 0.04025
R39064 VDD.n7552 VDD.n7221 0.04025
R39065 VDD.n7548 VDD.n7221 0.04025
R39066 VDD.n7548 VDD.n7547 0.04025
R39067 VDD.n7547 VDD.n7546 0.04025
R39068 VDD.n7546 VDD.n7223 0.04025
R39069 VDD.n7542 VDD.n7223 0.04025
R39070 VDD.n7542 VDD.n7541 0.04025
R39071 VDD.n7541 VDD.n7540 0.04025
R39072 VDD.n7540 VDD.n7225 0.04025
R39073 VDD.n7536 VDD.n7225 0.04025
R39074 VDD.n7536 VDD.n7535 0.04025
R39075 VDD.n7535 VDD.n7534 0.04025
R39076 VDD.n7534 VDD.n7227 0.04025
R39077 VDD.n7530 VDD.n7227 0.04025
R39078 VDD.n7530 VDD.n7529 0.04025
R39079 VDD.n7529 VDD.n7528 0.04025
R39080 VDD.n7528 VDD.n7229 0.04025
R39081 VDD.n7524 VDD.n7229 0.04025
R39082 VDD.n7524 VDD.n7523 0.04025
R39083 VDD.n7523 VDD.n7522 0.04025
R39084 VDD.n7522 VDD.n7231 0.04025
R39085 VDD.n7518 VDD.n7231 0.04025
R39086 VDD.n7518 VDD.n7517 0.04025
R39087 VDD.n7517 VDD.n7516 0.04025
R39088 VDD.n7516 VDD.n7233 0.04025
R39089 VDD.n7512 VDD.n7233 0.04025
R39090 VDD.n7512 VDD.n7511 0.04025
R39091 VDD.n7511 VDD.n7510 0.04025
R39092 VDD.n7510 VDD.n7235 0.04025
R39093 VDD.n7506 VDD.n7235 0.04025
R39094 VDD.n7506 VDD.n7505 0.04025
R39095 VDD.n7505 VDD.n7504 0.04025
R39096 VDD.n7504 VDD.n7237 0.04025
R39097 VDD.n7500 VDD.n7237 0.04025
R39098 VDD.n7500 VDD.n7499 0.04025
R39099 VDD.n7499 VDD.n7498 0.04025
R39100 VDD.n7498 VDD.n7239 0.04025
R39101 VDD.n7494 VDD.n7239 0.04025
R39102 VDD.n7494 VDD.n7493 0.04025
R39103 VDD.n7493 VDD.n7492 0.04025
R39104 VDD.n7492 VDD.n7241 0.04025
R39105 VDD.n7488 VDD.n7241 0.04025
R39106 VDD.n7488 VDD.n7487 0.04025
R39107 VDD.n7487 VDD.n7486 0.04025
R39108 VDD.n7486 VDD.n7243 0.04025
R39109 VDD.n7482 VDD.n7243 0.04025
R39110 VDD.n7482 VDD.n7481 0.04025
R39111 VDD.n7481 VDD.n7480 0.04025
R39112 VDD.n7480 VDD.n7245 0.04025
R39113 VDD.n7476 VDD.n7245 0.04025
R39114 VDD.n7476 VDD.n7475 0.04025
R39115 VDD.n7475 VDD.n7474 0.04025
R39116 VDD.n7474 VDD.n7247 0.04025
R39117 VDD.n7470 VDD.n7247 0.04025
R39118 VDD.n7470 VDD.n7469 0.04025
R39119 VDD.n7469 VDD.n7468 0.04025
R39120 VDD.n7468 VDD.n7249 0.04025
R39121 VDD.n7464 VDD.n7249 0.04025
R39122 VDD.n7464 VDD.n7463 0.04025
R39123 VDD.n7463 VDD.n7462 0.04025
R39124 VDD.n7462 VDD.n7251 0.04025
R39125 VDD.n7458 VDD.n7251 0.04025
R39126 VDD.n7458 VDD.n7457 0.04025
R39127 VDD.n7457 VDD.n7456 0.04025
R39128 VDD.n7456 VDD.n7253 0.04025
R39129 VDD.n7452 VDD.n7253 0.04025
R39130 VDD.n7452 VDD.n7451 0.04025
R39131 VDD.n7451 VDD.n7450 0.04025
R39132 VDD.n7450 VDD.n7255 0.04025
R39133 VDD.n7446 VDD.n7255 0.04025
R39134 VDD.n7446 VDD.n7445 0.04025
R39135 VDD.n7445 VDD.n7444 0.04025
R39136 VDD.n7444 VDD.n7257 0.04025
R39137 VDD.n7440 VDD.n7257 0.04025
R39138 VDD.n7440 VDD.n7439 0.04025
R39139 VDD.n7439 VDD.n7438 0.04025
R39140 VDD.n7438 VDD.n7259 0.04025
R39141 VDD.n7434 VDD.n7259 0.04025
R39142 VDD.n7434 VDD.n7433 0.04025
R39143 VDD.n7433 VDD.n7432 0.04025
R39144 VDD.n7432 VDD.n7261 0.04025
R39145 VDD.n7428 VDD.n7261 0.04025
R39146 VDD.n7428 VDD.n7427 0.04025
R39147 VDD.n7427 VDD.n7426 0.04025
R39148 VDD.n7426 VDD.n7263 0.04025
R39149 VDD.n7422 VDD.n7263 0.04025
R39150 VDD.n7422 VDD.n7421 0.04025
R39151 VDD.n7421 VDD.n7420 0.04025
R39152 VDD.n7420 VDD.n7265 0.04025
R39153 VDD.n7416 VDD.n7265 0.04025
R39154 VDD.n7416 VDD.n7415 0.04025
R39155 VDD.n7415 VDD.n7414 0.04025
R39156 VDD.n7414 VDD.n7267 0.04025
R39157 VDD.n7410 VDD.n7267 0.04025
R39158 VDD.n7410 VDD.n7409 0.04025
R39159 VDD.n7409 VDD.n7408 0.04025
R39160 VDD.n7408 VDD.n7269 0.04025
R39161 VDD.n7404 VDD.n7269 0.04025
R39162 VDD.n7404 VDD.n7403 0.04025
R39163 VDD.n7403 VDD.n7402 0.04025
R39164 VDD.n7402 VDD.n7271 0.04025
R39165 VDD.n7398 VDD.n7271 0.04025
R39166 VDD.n7398 VDD.n7397 0.04025
R39167 VDD.n7397 VDD.n7396 0.04025
R39168 VDD.n7396 VDD.n7273 0.04025
R39169 VDD.n7392 VDD.n7273 0.04025
R39170 VDD.n7392 VDD.n7391 0.04025
R39171 VDD.n7391 VDD.n7390 0.04025
R39172 VDD.n7390 VDD.n7275 0.04025
R39173 VDD.n7386 VDD.n7275 0.04025
R39174 VDD.n7386 VDD.n7385 0.04025
R39175 VDD.n7385 VDD.n7384 0.04025
R39176 VDD.n7384 VDD.n7277 0.04025
R39177 VDD.n7380 VDD.n7277 0.04025
R39178 VDD.n7380 VDD.n7379 0.04025
R39179 VDD.n7379 VDD.n7378 0.04025
R39180 VDD.n7378 VDD.n7279 0.04025
R39181 VDD.n7374 VDD.n7279 0.04025
R39182 VDD.n7374 VDD.n7373 0.04025
R39183 VDD.n7373 VDD.n7372 0.04025
R39184 VDD.n7372 VDD.n7281 0.04025
R39185 VDD.n7368 VDD.n7281 0.04025
R39186 VDD.n7368 VDD.n7367 0.04025
R39187 VDD.n7367 VDD.n7366 0.04025
R39188 VDD.n7366 VDD.n7283 0.04025
R39189 VDD.n7362 VDD.n7283 0.04025
R39190 VDD.n7362 VDD.n7361 0.04025
R39191 VDD.n7361 VDD.n7360 0.04025
R39192 VDD.n7360 VDD.n7285 0.04025
R39193 VDD.n7356 VDD.n7285 0.04025
R39194 VDD.n7356 VDD.n7355 0.04025
R39195 VDD.n7355 VDD.n7354 0.04025
R39196 VDD.n7354 VDD.n7287 0.04025
R39197 VDD.n7350 VDD.n7287 0.04025
R39198 VDD.n7350 VDD.n7349 0.04025
R39199 VDD.n7349 VDD.n7348 0.04025
R39200 VDD.n7348 VDD.n7289 0.04025
R39201 VDD.n7344 VDD.n7289 0.04025
R39202 VDD.n7344 VDD.n7343 0.04025
R39203 VDD.n7343 VDD.n7342 0.04025
R39204 VDD.n7342 VDD.n7291 0.04025
R39205 VDD.n7338 VDD.n7291 0.04025
R39206 VDD.n7338 VDD.n7337 0.04025
R39207 VDD.n7337 VDD.n7336 0.04025
R39208 VDD.n7336 VDD.n7293 0.04025
R39209 VDD.n7332 VDD.n7293 0.04025
R39210 VDD.n7332 VDD.n7331 0.04025
R39211 VDD.n7331 VDD.n7330 0.04025
R39212 VDD.n7330 VDD.n7295 0.04025
R39213 VDD.n7326 VDD.n7295 0.04025
R39214 VDD.n7326 VDD.n7325 0.04025
R39215 VDD.n7325 VDD.n7324 0.04025
R39216 VDD.n7324 VDD.n7297 0.04025
R39217 VDD.n7320 VDD.n7297 0.04025
R39218 VDD.n7320 VDD.n7319 0.04025
R39219 VDD.n7319 VDD.n7318 0.04025
R39220 VDD.n7318 VDD.n7299 0.04025
R39221 VDD.n7314 VDD.n7299 0.04025
R39222 VDD.n7314 VDD.n7313 0.04025
R39223 VDD.n7313 VDD.n7312 0.04025
R39224 VDD.n7312 VDD.n7301 0.04025
R39225 VDD.n7308 VDD.n7301 0.04025
R39226 VDD.n7308 VDD.n7307 0.04025
R39227 VDD.n7307 VDD.n7306 0.04025
R39228 VDD.n7306 VDD.n7303 0.04025
R39229 VDD.n7303 VDD.n2087 0.04025
R39230 VDD.n8169 VDD.n2087 0.04025
R39231 VDD.n8170 VDD.n8169 0.04025
R39232 VDD.n8171 VDD.n8170 0.04025
R39233 VDD.n8171 VDD.n2085 0.04025
R39234 VDD.n8176 VDD.n2085 0.04025
R39235 VDD.n8177 VDD.n8176 0.04025
R39236 VDD.n8178 VDD.n8177 0.04025
R39237 VDD.n8178 VDD.n2083 0.04025
R39238 VDD.n8184 VDD.n2083 0.04025
R39239 VDD.n8185 VDD.n8184 0.04025
R39240 VDD.n8186 VDD.n8185 0.04025
R39241 VDD.n8186 VDD.n2081 0.04025
R39242 VDD.n8191 VDD.n2081 0.04025
R39243 VDD.n8192 VDD.n8191 0.04025
R39244 VDD.n8193 VDD.n8192 0.04025
R39245 VDD.n8193 VDD.n2079 0.04025
R39246 VDD.n8197 VDD.n2079 0.04025
R39247 VDD.n8198 VDD.n8197 0.04025
R39248 VDD.n8198 VDD.n2077 0.04025
R39249 VDD.n8204 VDD.n2077 0.04025
R39250 VDD.n8205 VDD.n8204 0.04025
R39251 VDD.n8206 VDD.n8205 0.04025
R39252 VDD.n8206 VDD.n2075 0.04025
R39253 VDD.n8210 VDD.n2075 0.04025
R39254 VDD.n8211 VDD.n8210 0.04025
R39255 VDD.n8211 VDD.n2073 0.04025
R39256 VDD.n8217 VDD.n2073 0.04025
R39257 VDD.n8218 VDD.n8217 0.04025
R39258 VDD.n8219 VDD.n8218 0.04025
R39259 VDD.n8219 VDD.n2071 0.04025
R39260 VDD.n8224 VDD.n2071 0.04025
R39261 VDD.n8225 VDD.n8224 0.04025
R39262 VDD.n8226 VDD.n8225 0.04025
R39263 VDD.n8226 VDD.n2069 0.04025
R39264 VDD.n8231 VDD.n2069 0.04025
R39265 VDD.n8232 VDD.n8231 0.04025
R39266 VDD.n8233 VDD.n8232 0.04025
R39267 VDD.n8233 VDD.n2067 0.04025
R39268 VDD.n8239 VDD.n2067 0.04025
R39269 VDD.n8240 VDD.n8239 0.04025
R39270 VDD.n8241 VDD.n8240 0.04025
R39271 VDD.n8241 VDD.n2065 0.04025
R39272 VDD.n8245 VDD.n2065 0.04025
R39273 VDD.n8246 VDD.n8245 0.04025
R39274 VDD.n8246 VDD.n2063 0.04025
R39275 VDD.n8252 VDD.n2063 0.04025
R39276 VDD.n8253 VDD.n8252 0.04025
R39277 VDD.n10764 VDD.n8253 0.04025
R39278 VDD.n10764 VDD.n10763 0.04025
R39279 VDD.n10763 VDD.n10762 0.04025
R39280 VDD.n10762 VDD.n8254 0.04025
R39281 VDD.n10758 VDD.n8254 0.04025
R39282 VDD.n10758 VDD.n10757 0.04025
R39283 VDD.n10757 VDD.n10756 0.04025
R39284 VDD.n10756 VDD.n8256 0.04025
R39285 VDD.n10752 VDD.n8256 0.04025
R39286 VDD.n10752 VDD.n10751 0.04025
R39287 VDD.n10751 VDD.n10750 0.04025
R39288 VDD.n10750 VDD.n8258 0.04025
R39289 VDD.n10746 VDD.n8258 0.04025
R39290 VDD.n10746 VDD.n10745 0.04025
R39291 VDD.n10745 VDD.n10744 0.04025
R39292 VDD.n10744 VDD.n8260 0.04025
R39293 VDD.n10740 VDD.n8260 0.04025
R39294 VDD.n10740 VDD.n10739 0.04025
R39295 VDD.n10739 VDD.n10738 0.04025
R39296 VDD.n10738 VDD.n8262 0.04025
R39297 VDD.n10734 VDD.n8262 0.04025
R39298 VDD.n10734 VDD.n10733 0.04025
R39299 VDD.n10733 VDD.n10732 0.04025
R39300 VDD.n10732 VDD.n8264 0.04025
R39301 VDD.n10728 VDD.n8264 0.04025
R39302 VDD.n10728 VDD.n10727 0.04025
R39303 VDD.n10727 VDD.n10726 0.04025
R39304 VDD.n10726 VDD.n8266 0.04025
R39305 VDD.n10722 VDD.n8266 0.04025
R39306 VDD.n10722 VDD.n10721 0.04025
R39307 VDD.n10721 VDD.n10720 0.04025
R39308 VDD.n10720 VDD.n8268 0.04025
R39309 VDD.n10716 VDD.n8268 0.04025
R39310 VDD.n10716 VDD.n10715 0.04025
R39311 VDD.n10715 VDD.n10714 0.04025
R39312 VDD.n10714 VDD.n8270 0.04025
R39313 VDD.n10710 VDD.n8270 0.04025
R39314 VDD.n10710 VDD.n10709 0.04025
R39315 VDD.n10709 VDD.n10708 0.04025
R39316 VDD.n10708 VDD.n8272 0.04025
R39317 VDD.n10704 VDD.n8272 0.04025
R39318 VDD.n10704 VDD.n10703 0.04025
R39319 VDD.n10703 VDD.n10702 0.04025
R39320 VDD.n10702 VDD.n8274 0.04025
R39321 VDD.n10698 VDD.n8274 0.04025
R39322 VDD.n10698 VDD.n10697 0.04025
R39323 VDD.n10697 VDD.n10696 0.04025
R39324 VDD.n10696 VDD.n8276 0.04025
R39325 VDD.n10692 VDD.n8276 0.04025
R39326 VDD.n10692 VDD.n10691 0.04025
R39327 VDD.n10691 VDD.n10690 0.04025
R39328 VDD.n10690 VDD.n8278 0.04025
R39329 VDD.n10686 VDD.n8278 0.04025
R39330 VDD.n10686 VDD.n10685 0.04025
R39331 VDD.n10685 VDD.n10684 0.04025
R39332 VDD.n10684 VDD.n8280 0.04025
R39333 VDD.n10680 VDD.n8280 0.04025
R39334 VDD.n10680 VDD.n10679 0.04025
R39335 VDD.n10679 VDD.n10678 0.04025
R39336 VDD.n10678 VDD.n8282 0.04025
R39337 VDD.n10674 VDD.n8282 0.04025
R39338 VDD.n10674 VDD.n10673 0.04025
R39339 VDD.n10673 VDD.n10672 0.04025
R39340 VDD.n10672 VDD.n8284 0.04025
R39341 VDD.n10668 VDD.n8284 0.04025
R39342 VDD.n10668 VDD.n10667 0.04025
R39343 VDD.n10667 VDD.n10666 0.04025
R39344 VDD.n10666 VDD.n8286 0.04025
R39345 VDD.n10662 VDD.n8286 0.04025
R39346 VDD.n10662 VDD.n10661 0.04025
R39347 VDD.n10661 VDD.n10660 0.04025
R39348 VDD.n10660 VDD.n8288 0.04025
R39349 VDD.n10656 VDD.n8288 0.04025
R39350 VDD.n10656 VDD.n10655 0.04025
R39351 VDD.n10655 VDD.n10654 0.04025
R39352 VDD.n10654 VDD.n8290 0.04025
R39353 VDD.n10650 VDD.n8290 0.04025
R39354 VDD.n10650 VDD.n10649 0.04025
R39355 VDD.n10649 VDD.n10648 0.04025
R39356 VDD.n10648 VDD.n8292 0.04025
R39357 VDD.n10644 VDD.n8292 0.04025
R39358 VDD.n10644 VDD.n10643 0.04025
R39359 VDD.n10643 VDD.n10642 0.04025
R39360 VDD.n10642 VDD.n8294 0.04025
R39361 VDD.n10638 VDD.n8294 0.04025
R39362 VDD.n10638 VDD.n10637 0.04025
R39363 VDD.n10637 VDD.n10636 0.04025
R39364 VDD.n10636 VDD.n8296 0.04025
R39365 VDD.n10632 VDD.n8296 0.04025
R39366 VDD.n10632 VDD.n10631 0.04025
R39367 VDD.n10631 VDD.n10630 0.04025
R39368 VDD.n10630 VDD.n8298 0.04025
R39369 VDD.n10626 VDD.n8298 0.04025
R39370 VDD.n10626 VDD.n10625 0.04025
R39371 VDD.n10625 VDD.n10624 0.04025
R39372 VDD.n10624 VDD.n8300 0.04025
R39373 VDD.n10620 VDD.n8300 0.04025
R39374 VDD.n10620 VDD.n10619 0.04025
R39375 VDD.n10619 VDD.n10618 0.04025
R39376 VDD.n10618 VDD.n8302 0.04025
R39377 VDD.n10614 VDD.n8302 0.04025
R39378 VDD.n10614 VDD.n10613 0.04025
R39379 VDD.n10613 VDD.n10612 0.04025
R39380 VDD.n10612 VDD.n8304 0.04025
R39381 VDD.n10608 VDD.n8304 0.04025
R39382 VDD.n10608 VDD.n10607 0.04025
R39383 VDD.n10607 VDD.n10606 0.04025
R39384 VDD.n10606 VDD.n8306 0.04025
R39385 VDD.n10602 VDD.n8306 0.04025
R39386 VDD.n10602 VDD.n10601 0.04025
R39387 VDD.n10601 VDD.n10600 0.04025
R39388 VDD.n10600 VDD.n8308 0.04025
R39389 VDD.n10596 VDD.n8308 0.04025
R39390 VDD.n10596 VDD.n10595 0.04025
R39391 VDD.n10595 VDD.n10594 0.04025
R39392 VDD.n10594 VDD.n8310 0.04025
R39393 VDD.n10590 VDD.n8310 0.04025
R39394 VDD.n10590 VDD.n10589 0.04025
R39395 VDD.n10589 VDD.n10588 0.04025
R39396 VDD.n10588 VDD.n8312 0.04025
R39397 VDD.n10584 VDD.n8312 0.04025
R39398 VDD.n10584 VDD.n10583 0.04025
R39399 VDD.n10583 VDD.n10582 0.04025
R39400 VDD.n10582 VDD.n8314 0.04025
R39401 VDD.n10578 VDD.n8314 0.04025
R39402 VDD.n10578 VDD.n10577 0.04025
R39403 VDD.n10577 VDD.n10576 0.04025
R39404 VDD.n10576 VDD.n8316 0.04025
R39405 VDD.n10572 VDD.n8316 0.04025
R39406 VDD.n10572 VDD.n10571 0.04025
R39407 VDD.n10571 VDD.n10570 0.04025
R39408 VDD.n10570 VDD.n8318 0.04025
R39409 VDD.n10566 VDD.n8318 0.04025
R39410 VDD.n10566 VDD.n10565 0.04025
R39411 VDD.n10565 VDD.n10564 0.04025
R39412 VDD.n10564 VDD.n8320 0.04025
R39413 VDD.n10560 VDD.n8320 0.04025
R39414 VDD.n10560 VDD.n10559 0.04025
R39415 VDD.n10559 VDD.n10558 0.04025
R39416 VDD.n10558 VDD.n8322 0.04025
R39417 VDD.n10554 VDD.n8322 0.04025
R39418 VDD.n10554 VDD.n10553 0.04025
R39419 VDD.n10553 VDD.n10552 0.04025
R39420 VDD.n10552 VDD.n8324 0.04025
R39421 VDD.n10548 VDD.n8324 0.04025
R39422 VDD.n10548 VDD.n10547 0.04025
R39423 VDD.n10547 VDD.n10546 0.04025
R39424 VDD.n10546 VDD.n8326 0.04025
R39425 VDD.n10542 VDD.n8326 0.04025
R39426 VDD.n10542 VDD.n10541 0.04025
R39427 VDD.n10541 VDD.n10540 0.04025
R39428 VDD.n10540 VDD.n8328 0.04025
R39429 VDD.n10536 VDD.n8328 0.04025
R39430 VDD.n10536 VDD.n10535 0.04025
R39431 VDD.n10535 VDD.n10534 0.04025
R39432 VDD.n10534 VDD.n8330 0.04025
R39433 VDD.n10530 VDD.n8330 0.04025
R39434 VDD.n10530 VDD.n10529 0.04025
R39435 VDD.n10529 VDD.n10528 0.04025
R39436 VDD.n10528 VDD.n8332 0.04025
R39437 VDD.n10524 VDD.n8332 0.04025
R39438 VDD.n10524 VDD.n10523 0.04025
R39439 VDD.n10523 VDD.n10522 0.04025
R39440 VDD.n10522 VDD.n8334 0.04025
R39441 VDD.n10518 VDD.n8334 0.04025
R39442 VDD.n10518 VDD.n10517 0.04025
R39443 VDD.n10517 VDD.n10516 0.04025
R39444 VDD.n10516 VDD.n8336 0.04025
R39445 VDD.n10512 VDD.n8336 0.04025
R39446 VDD.n10512 VDD.n10511 0.04025
R39447 VDD.n10511 VDD.n10510 0.04025
R39448 VDD.n10510 VDD.n8338 0.04025
R39449 VDD.n10506 VDD.n8338 0.04025
R39450 VDD.n10506 VDD.n10505 0.04025
R39451 VDD.n10505 VDD.n10504 0.04025
R39452 VDD.n10504 VDD.n8340 0.04025
R39453 VDD.n10500 VDD.n8340 0.04025
R39454 VDD.n10500 VDD.n10499 0.04025
R39455 VDD.n10499 VDD.n10498 0.04025
R39456 VDD.n10498 VDD.n8342 0.04025
R39457 VDD.n10494 VDD.n8342 0.04025
R39458 VDD.n10494 VDD.n10493 0.04025
R39459 VDD.n10493 VDD.n10492 0.04025
R39460 VDD.n10492 VDD.n8344 0.04025
R39461 VDD.n10488 VDD.n8344 0.04025
R39462 VDD.n10488 VDD.n10487 0.04025
R39463 VDD.n10487 VDD.n10486 0.04025
R39464 VDD.n10486 VDD.n8346 0.04025
R39465 VDD.n10482 VDD.n8346 0.04025
R39466 VDD.n10482 VDD.n10481 0.04025
R39467 VDD.n10481 VDD.n10480 0.04025
R39468 VDD.n10480 VDD.n8348 0.04025
R39469 VDD.n10476 VDD.n8348 0.04025
R39470 VDD.n10476 VDD.n10475 0.04025
R39471 VDD.n10475 VDD.n10474 0.04025
R39472 VDD.n10474 VDD.n8350 0.04025
R39473 VDD.n10470 VDD.n8350 0.04025
R39474 VDD.n10470 VDD.n10469 0.04025
R39475 VDD.n10469 VDD.n10468 0.04025
R39476 VDD.n10468 VDD.n8352 0.04025
R39477 VDD.n10464 VDD.n8352 0.04025
R39478 VDD.n10464 VDD.n10463 0.04025
R39479 VDD.n10463 VDD.n10462 0.04025
R39480 VDD.n10462 VDD.n8354 0.04025
R39481 VDD.n10458 VDD.n8354 0.04025
R39482 VDD.n10458 VDD.n10457 0.04025
R39483 VDD.n10457 VDD.n10456 0.04025
R39484 VDD.n10456 VDD.n8356 0.04025
R39485 VDD.n10452 VDD.n8356 0.04025
R39486 VDD.n10452 VDD.n10451 0.04025
R39487 VDD.n10451 VDD.n10450 0.04025
R39488 VDD.n10450 VDD.n8358 0.04025
R39489 VDD.n10446 VDD.n8358 0.04025
R39490 VDD.n10446 VDD.n10445 0.04025
R39491 VDD.n10445 VDD.n10444 0.04025
R39492 VDD.n10444 VDD.n8360 0.04025
R39493 VDD.n10440 VDD.n8360 0.04025
R39494 VDD.n10440 VDD.n10439 0.04025
R39495 VDD.n10439 VDD.n10438 0.04025
R39496 VDD.n10438 VDD.n8362 0.04025
R39497 VDD.n10434 VDD.n8362 0.04025
R39498 VDD.n10434 VDD.n10433 0.04025
R39499 VDD.n10433 VDD.n10432 0.04025
R39500 VDD.n10432 VDD.n8364 0.04025
R39501 VDD.n10428 VDD.n8364 0.04025
R39502 VDD.n10428 VDD.n10427 0.04025
R39503 VDD.n10427 VDD.n10426 0.04025
R39504 VDD.n10426 VDD.n8366 0.04025
R39505 VDD.n10422 VDD.n8366 0.04025
R39506 VDD.n10422 VDD.n10421 0.04025
R39507 VDD.n10421 VDD.n10420 0.04025
R39508 VDD.n10420 VDD.n8368 0.04025
R39509 VDD.n10416 VDD.n8368 0.04025
R39510 VDD.n10416 VDD.n10415 0.04025
R39511 VDD.n10415 VDD.n10414 0.04025
R39512 VDD.n10414 VDD.n8370 0.04025
R39513 VDD.n10410 VDD.n8370 0.04025
R39514 VDD.n10410 VDD.n10409 0.04025
R39515 VDD.n10409 VDD.n10408 0.04025
R39516 VDD.n10408 VDD.n8372 0.04025
R39517 VDD.n10404 VDD.n8372 0.04025
R39518 VDD.n10404 VDD.n10403 0.04025
R39519 VDD.n10403 VDD.n10402 0.04025
R39520 VDD.n10402 VDD.n8374 0.04025
R39521 VDD.n10398 VDD.n8374 0.04025
R39522 VDD.n10398 VDD.n10397 0.04025
R39523 VDD.n10397 VDD.n10396 0.04025
R39524 VDD.n10396 VDD.n8376 0.04025
R39525 VDD.n10392 VDD.n8376 0.04025
R39526 VDD.n10392 VDD.n10391 0.04025
R39527 VDD.n10391 VDD.n10390 0.04025
R39528 VDD.n10390 VDD.n8378 0.04025
R39529 VDD.n10386 VDD.n8378 0.04025
R39530 VDD.n10386 VDD.n10385 0.04025
R39531 VDD.n10385 VDD.n10384 0.04025
R39532 VDD.n10384 VDD.n8380 0.04025
R39533 VDD.n10380 VDD.n8380 0.04025
R39534 VDD.n10380 VDD.n10379 0.04025
R39535 VDD.n10379 VDD.n10378 0.04025
R39536 VDD.n10378 VDD.n8382 0.04025
R39537 VDD.n10374 VDD.n8382 0.04025
R39538 VDD.n10374 VDD.n10373 0.04025
R39539 VDD.n10373 VDD.n10372 0.04025
R39540 VDD.n10372 VDD.n8384 0.04025
R39541 VDD.n10368 VDD.n8384 0.04025
R39542 VDD.n10368 VDD.n10367 0.04025
R39543 VDD.n10367 VDD.n10366 0.04025
R39544 VDD.n10366 VDD.n8386 0.04025
R39545 VDD.n10362 VDD.n8386 0.04025
R39546 VDD.n10362 VDD.n10361 0.04025
R39547 VDD.n10361 VDD.n10360 0.04025
R39548 VDD.n10360 VDD.n8388 0.04025
R39549 VDD.n10356 VDD.n8388 0.04025
R39550 VDD.n10356 VDD.n10355 0.04025
R39551 VDD.n10355 VDD.n10354 0.04025
R39552 VDD.n10354 VDD.n8390 0.04025
R39553 VDD.n10350 VDD.n8390 0.04025
R39554 VDD.n10350 VDD.n10349 0.04025
R39555 VDD.n10349 VDD.n10348 0.04025
R39556 VDD.n10348 VDD.n8392 0.04025
R39557 VDD.n10344 VDD.n8392 0.04025
R39558 VDD.n10344 VDD.n10343 0.04025
R39559 VDD.n10343 VDD.n10342 0.04025
R39560 VDD.n10342 VDD.n8394 0.04025
R39561 VDD.n10338 VDD.n8394 0.04025
R39562 VDD.n10338 VDD.n10337 0.04025
R39563 VDD.n10337 VDD.n10336 0.04025
R39564 VDD.n10336 VDD.n8396 0.04025
R39565 VDD.n10332 VDD.n8396 0.04025
R39566 VDD.n10332 VDD.n10331 0.04025
R39567 VDD.n10331 VDD.n10330 0.04025
R39568 VDD.n10330 VDD.n8398 0.04025
R39569 VDD.n10326 VDD.n8398 0.04025
R39570 VDD.n10326 VDD.n10325 0.04025
R39571 VDD.n10325 VDD.n10324 0.04025
R39572 VDD.n10324 VDD.n8400 0.04025
R39573 VDD.n10320 VDD.n8400 0.04025
R39574 VDD.n10320 VDD.n10319 0.04025
R39575 VDD.n10319 VDD.n10318 0.04025
R39576 VDD.n10318 VDD.n8402 0.04025
R39577 VDD.n10314 VDD.n8402 0.04025
R39578 VDD.n10314 VDD.n10313 0.04025
R39579 VDD.n10313 VDD.n10312 0.04025
R39580 VDD.n10312 VDD.n8404 0.04025
R39581 VDD.n10308 VDD.n8404 0.04025
R39582 VDD.n10308 VDD.n10307 0.04025
R39583 VDD.n10307 VDD.n10306 0.04025
R39584 VDD.n10306 VDD.n8406 0.04025
R39585 VDD.n10302 VDD.n8406 0.04025
R39586 VDD.n10302 VDD.n10301 0.04025
R39587 VDD.n10301 VDD.n10300 0.04025
R39588 VDD.n10300 VDD.n8408 0.04025
R39589 VDD.n10296 VDD.n8408 0.04025
R39590 VDD.n10296 VDD.n10295 0.04025
R39591 VDD.n10295 VDD.n10294 0.04025
R39592 VDD.n10294 VDD.n8410 0.04025
R39593 VDD.n10290 VDD.n8410 0.04025
R39594 VDD.n10290 VDD.n10289 0.04025
R39595 VDD.n10289 VDD.n10288 0.04025
R39596 VDD.n10288 VDD.n8412 0.04025
R39597 VDD.n10284 VDD.n8412 0.04025
R39598 VDD.n10284 VDD.n10283 0.04025
R39599 VDD.n10283 VDD.n10282 0.04025
R39600 VDD.n10282 VDD.n8414 0.04025
R39601 VDD.n10278 VDD.n8414 0.04025
R39602 VDD.n10278 VDD.n10277 0.04025
R39603 VDD.n10277 VDD.n10276 0.04025
R39604 VDD.n10276 VDD.n8416 0.04025
R39605 VDD.n10272 VDD.n8416 0.04025
R39606 VDD.n10272 VDD.n10271 0.04025
R39607 VDD.n10271 VDD.n10270 0.04025
R39608 VDD.n10270 VDD.n8418 0.04025
R39609 VDD.n10266 VDD.n8418 0.04025
R39610 VDD.n10266 VDD.n10265 0.04025
R39611 VDD.n10265 VDD.n10264 0.04025
R39612 VDD.n10264 VDD.n8420 0.04025
R39613 VDD.n10260 VDD.n8420 0.04025
R39614 VDD.n10260 VDD.n10259 0.04025
R39615 VDD.n10259 VDD.n10258 0.04025
R39616 VDD.n10258 VDD.n8422 0.04025
R39617 VDD.n10254 VDD.n8422 0.04025
R39618 VDD.n10254 VDD.n10253 0.04025
R39619 VDD.n10253 VDD.n10252 0.04025
R39620 VDD.n10252 VDD.n8424 0.04025
R39621 VDD.n10248 VDD.n8424 0.04025
R39622 VDD.n10248 VDD.n10247 0.04025
R39623 VDD.n10247 VDD.n10246 0.04025
R39624 VDD.n10246 VDD.n8426 0.04025
R39625 VDD.n10242 VDD.n8426 0.04025
R39626 VDD.n10242 VDD.n10241 0.04025
R39627 VDD.n10241 VDD.n10240 0.04025
R39628 VDD.n10240 VDD.n8428 0.04025
R39629 VDD.n10236 VDD.n8428 0.04025
R39630 VDD.n10236 VDD.n10235 0.04025
R39631 VDD.n10235 VDD.n10234 0.04025
R39632 VDD.n10234 VDD.n8430 0.04025
R39633 VDD.n10230 VDD.n8430 0.04025
R39634 VDD.n10230 VDD.n10229 0.04025
R39635 VDD.n10229 VDD.n10228 0.04025
R39636 VDD.n10228 VDD.n8432 0.04025
R39637 VDD.n10224 VDD.n8432 0.04025
R39638 VDD.n10224 VDD.n10223 0.04025
R39639 VDD.n10223 VDD.n10222 0.04025
R39640 VDD.n10222 VDD.n8434 0.04025
R39641 VDD.n10218 VDD.n8434 0.04025
R39642 VDD.n10218 VDD.n10217 0.04025
R39643 VDD.n10217 VDD.n10216 0.04025
R39644 VDD.n10216 VDD.n8436 0.04025
R39645 VDD.n10212 VDD.n8436 0.04025
R39646 VDD.n10212 VDD.n10211 0.04025
R39647 VDD.n10211 VDD.n10210 0.04025
R39648 VDD.n10210 VDD.n8438 0.04025
R39649 VDD.n10206 VDD.n8438 0.04025
R39650 VDD.n10206 VDD.n10205 0.04025
R39651 VDD.n10205 VDD.n10204 0.04025
R39652 VDD.n10204 VDD.n8440 0.04025
R39653 VDD.n10200 VDD.n8440 0.04025
R39654 VDD.n10200 VDD.n10199 0.04025
R39655 VDD.n10199 VDD.n10198 0.04025
R39656 VDD.n10198 VDD.n8442 0.04025
R39657 VDD.n10194 VDD.n8442 0.04025
R39658 VDD.n10194 VDD.n10193 0.04025
R39659 VDD.n10193 VDD.n10192 0.04025
R39660 VDD.n10192 VDD.n8444 0.04025
R39661 VDD.n10188 VDD.n8444 0.04025
R39662 VDD.n10188 VDD.n10187 0.04025
R39663 VDD.n10187 VDD.n10186 0.04025
R39664 VDD.n10186 VDD.n8446 0.04025
R39665 VDD.n10182 VDD.n8446 0.04025
R39666 VDD.n10182 VDD.n10181 0.04025
R39667 VDD.n10181 VDD.n10180 0.04025
R39668 VDD.n10180 VDD.n8448 0.04025
R39669 VDD.n10176 VDD.n8448 0.04025
R39670 VDD.n10176 VDD.n10175 0.04025
R39671 VDD.n10175 VDD.n10174 0.04025
R39672 VDD.n10174 VDD.n8450 0.04025
R39673 VDD.n10170 VDD.n8450 0.04025
R39674 VDD.n10170 VDD.n10169 0.04025
R39675 VDD.n10169 VDD.n10168 0.04025
R39676 VDD.n10168 VDD.n8452 0.04025
R39677 VDD.n10164 VDD.n8452 0.04025
R39678 VDD.n10164 VDD.n10163 0.04025
R39679 VDD.n10163 VDD.n10162 0.04025
R39680 VDD.n10162 VDD.n8454 0.04025
R39681 VDD.n10158 VDD.n8454 0.04025
R39682 VDD.n10158 VDD.n10157 0.04025
R39683 VDD.n10157 VDD.n10156 0.04025
R39684 VDD.n10156 VDD.n8456 0.04025
R39685 VDD.n10152 VDD.n8456 0.04025
R39686 VDD.n10152 VDD.n10151 0.04025
R39687 VDD.n10151 VDD.n10150 0.04025
R39688 VDD.n10150 VDD.n8458 0.04025
R39689 VDD.n10146 VDD.n9200 0.04025
R39690 VDD.n10146 VDD.n10145 0.04025
R39691 VDD.n10145 VDD.n10144 0.04025
R39692 VDD.n10144 VDD.n9201 0.04025
R39693 VDD.n10140 VDD.n9201 0.04025
R39694 VDD.n10140 VDD.n10139 0.04025
R39695 VDD.n10139 VDD.n10138 0.04025
R39696 VDD.n10138 VDD.n9203 0.04025
R39697 VDD.n10134 VDD.n9203 0.04025
R39698 VDD.n10134 VDD.n10133 0.04025
R39699 VDD.n10133 VDD.n10132 0.04025
R39700 VDD.n10132 VDD.n9205 0.04025
R39701 VDD.n10128 VDD.n9205 0.04025
R39702 VDD.n10128 VDD.n10127 0.04025
R39703 VDD.n10127 VDD.n10126 0.04025
R39704 VDD.n10126 VDD.n9207 0.04025
R39705 VDD.n10122 VDD.n9207 0.04025
R39706 VDD.n10122 VDD.n10121 0.04025
R39707 VDD.n10121 VDD.n10120 0.04025
R39708 VDD.n10120 VDD.n9209 0.04025
R39709 VDD.n10116 VDD.n9209 0.04025
R39710 VDD.n10116 VDD.n10115 0.04025
R39711 VDD.n10115 VDD.n10114 0.04025
R39712 VDD.n10114 VDD.n9211 0.04025
R39713 VDD.n10110 VDD.n9211 0.04025
R39714 VDD.n10110 VDD.n10109 0.04025
R39715 VDD.n10109 VDD.n10108 0.04025
R39716 VDD.n10108 VDD.n9213 0.04025
R39717 VDD.n10104 VDD.n9213 0.04025
R39718 VDD.n10104 VDD.n10103 0.04025
R39719 VDD.n10147 VDD.n9186 0.04025
R39720 VDD.n10143 VDD.n9186 0.04025
R39721 VDD.n10143 VDD.n10142 0.04025
R39722 VDD.n10142 VDD.n10141 0.04025
R39723 VDD.n10141 VDD.n9202 0.04025
R39724 VDD.n10137 VDD.n9202 0.04025
R39725 VDD.n10137 VDD.n10136 0.04025
R39726 VDD.n10136 VDD.n10135 0.04025
R39727 VDD.n10135 VDD.n9204 0.04025
R39728 VDD.n10131 VDD.n9204 0.04025
R39729 VDD.n10131 VDD.n10130 0.04025
R39730 VDD.n10130 VDD.n10129 0.04025
R39731 VDD.n10129 VDD.n9206 0.04025
R39732 VDD.n10125 VDD.n9206 0.04025
R39733 VDD.n10125 VDD.n10124 0.04025
R39734 VDD.n10124 VDD.n10123 0.04025
R39735 VDD.n10123 VDD.n9208 0.04025
R39736 VDD.n10119 VDD.n9208 0.04025
R39737 VDD.n10119 VDD.n10118 0.04025
R39738 VDD.n10118 VDD.n10117 0.04025
R39739 VDD.n10117 VDD.n9210 0.04025
R39740 VDD.n10113 VDD.n9210 0.04025
R39741 VDD.n10113 VDD.n10112 0.04025
R39742 VDD.n10112 VDD.n10111 0.04025
R39743 VDD.n10111 VDD.n9212 0.04025
R39744 VDD.n10107 VDD.n9212 0.04025
R39745 VDD.n10107 VDD.n10106 0.04025
R39746 VDD.n10106 VDD.n10105 0.04025
R39747 VDD.n10105 VDD.n9214 0.04025
R39748 VDD.n9439 VDD.n9436 0.04025
R39749 VDD.n9440 VDD.n9439 0.04025
R39750 VDD.n9441 VDD.n9440 0.04025
R39751 VDD.n9441 VDD.n9434 0.04025
R39752 VDD.n9445 VDD.n9434 0.04025
R39753 VDD.n9446 VDD.n9445 0.04025
R39754 VDD.n9447 VDD.n9446 0.04025
R39755 VDD.n9447 VDD.n9432 0.04025
R39756 VDD.n9451 VDD.n9432 0.04025
R39757 VDD.n9452 VDD.n9451 0.04025
R39758 VDD.n9453 VDD.n9452 0.04025
R39759 VDD.n9453 VDD.n9430 0.04025
R39760 VDD.n9457 VDD.n9430 0.04025
R39761 VDD.n9458 VDD.n9457 0.04025
R39762 VDD.n9459 VDD.n9458 0.04025
R39763 VDD.n9459 VDD.n9428 0.04025
R39764 VDD.n9463 VDD.n9428 0.04025
R39765 VDD.n9464 VDD.n9463 0.04025
R39766 VDD.n9465 VDD.n9464 0.04025
R39767 VDD.n9465 VDD.n9426 0.04025
R39768 VDD.n9469 VDD.n9426 0.04025
R39769 VDD.n9470 VDD.n9469 0.04025
R39770 VDD.n9471 VDD.n9470 0.04025
R39771 VDD.n9471 VDD.n9424 0.04025
R39772 VDD.n9475 VDD.n9424 0.04025
R39773 VDD.n9476 VDD.n9475 0.04025
R39774 VDD.n9477 VDD.n9476 0.04025
R39775 VDD.n9477 VDD.n9422 0.04025
R39776 VDD.n9481 VDD.n9422 0.04025
R39777 VDD.n9482 VDD.n9481 0.04025
R39778 VDD.n9483 VDD.n9482 0.04025
R39779 VDD.n9483 VDD.n9420 0.04025
R39780 VDD.n9487 VDD.n9420 0.04025
R39781 VDD.n9488 VDD.n9487 0.04025
R39782 VDD.n9489 VDD.n9488 0.04025
R39783 VDD.n9489 VDD.n9418 0.04025
R39784 VDD.n9493 VDD.n9418 0.04025
R39785 VDD.n9494 VDD.n9493 0.04025
R39786 VDD.n9495 VDD.n9494 0.04025
R39787 VDD.n9495 VDD.n9416 0.04025
R39788 VDD.n9499 VDD.n9416 0.04025
R39789 VDD.n9500 VDD.n9499 0.04025
R39790 VDD.n9501 VDD.n9500 0.04025
R39791 VDD.n9501 VDD.n9414 0.04025
R39792 VDD.n9505 VDD.n9414 0.04025
R39793 VDD.n9506 VDD.n9505 0.04025
R39794 VDD.n9507 VDD.n9506 0.04025
R39795 VDD.n9507 VDD.n9412 0.04025
R39796 VDD.n9511 VDD.n9412 0.04025
R39797 VDD.n9512 VDD.n9511 0.04025
R39798 VDD.n9513 VDD.n9512 0.04025
R39799 VDD.n9513 VDD.n9410 0.04025
R39800 VDD.n9517 VDD.n9410 0.04025
R39801 VDD.n9518 VDD.n9517 0.04025
R39802 VDD.n9519 VDD.n9518 0.04025
R39803 VDD.n9519 VDD.n9408 0.04025
R39804 VDD.n9523 VDD.n9408 0.04025
R39805 VDD.n9524 VDD.n9523 0.04025
R39806 VDD.n9525 VDD.n9524 0.04025
R39807 VDD.n9525 VDD.n9406 0.04025
R39808 VDD.n9529 VDD.n9406 0.04025
R39809 VDD.n9530 VDD.n9529 0.04025
R39810 VDD.n9531 VDD.n9530 0.04025
R39811 VDD.n9531 VDD.n9404 0.04025
R39812 VDD.n9535 VDD.n9404 0.04025
R39813 VDD.n9536 VDD.n9535 0.04025
R39814 VDD.n9537 VDD.n9536 0.04025
R39815 VDD.n9537 VDD.n9402 0.04025
R39816 VDD.n9541 VDD.n9402 0.04025
R39817 VDD.n9542 VDD.n9541 0.04025
R39818 VDD.n9543 VDD.n9542 0.04025
R39819 VDD.n9543 VDD.n9400 0.04025
R39820 VDD.n9547 VDD.n9400 0.04025
R39821 VDD.n9548 VDD.n9547 0.04025
R39822 VDD.n9549 VDD.n9548 0.04025
R39823 VDD.n9549 VDD.n9398 0.04025
R39824 VDD.n9553 VDD.n9398 0.04025
R39825 VDD.n9554 VDD.n9553 0.04025
R39826 VDD.n9555 VDD.n9554 0.04025
R39827 VDD.n9555 VDD.n9396 0.04025
R39828 VDD.n9559 VDD.n9396 0.04025
R39829 VDD.n9560 VDD.n9559 0.04025
R39830 VDD.n9561 VDD.n9560 0.04025
R39831 VDD.n9561 VDD.n9394 0.04025
R39832 VDD.n9565 VDD.n9394 0.04025
R39833 VDD.n9566 VDD.n9565 0.04025
R39834 VDD.n9567 VDD.n9566 0.04025
R39835 VDD.n9567 VDD.n9392 0.04025
R39836 VDD.n9571 VDD.n9392 0.04025
R39837 VDD.n9572 VDD.n9571 0.04025
R39838 VDD.n9573 VDD.n9572 0.04025
R39839 VDD.n9573 VDD.n9390 0.04025
R39840 VDD.n9577 VDD.n9390 0.04025
R39841 VDD.n9578 VDD.n9577 0.04025
R39842 VDD.n9579 VDD.n9578 0.04025
R39843 VDD.n9579 VDD.n9388 0.04025
R39844 VDD.n9583 VDD.n9388 0.04025
R39845 VDD.n9584 VDD.n9583 0.04025
R39846 VDD.n9585 VDD.n9584 0.04025
R39847 VDD.n9585 VDD.n9386 0.04025
R39848 VDD.n9589 VDD.n9386 0.04025
R39849 VDD.n9590 VDD.n9589 0.04025
R39850 VDD.n9591 VDD.n9590 0.04025
R39851 VDD.n9591 VDD.n9384 0.04025
R39852 VDD.n9595 VDD.n9384 0.04025
R39853 VDD.n9596 VDD.n9595 0.04025
R39854 VDD.n9597 VDD.n9596 0.04025
R39855 VDD.n9597 VDD.n9382 0.04025
R39856 VDD.n9601 VDD.n9382 0.04025
R39857 VDD.n9602 VDD.n9601 0.04025
R39858 VDD.n9603 VDD.n9602 0.04025
R39859 VDD.n9603 VDD.n9380 0.04025
R39860 VDD.n9607 VDD.n9380 0.04025
R39861 VDD.n9608 VDD.n9607 0.04025
R39862 VDD.n9609 VDD.n9608 0.04025
R39863 VDD.n9609 VDD.n9378 0.04025
R39864 VDD.n9613 VDD.n9378 0.04025
R39865 VDD.n9614 VDD.n9613 0.04025
R39866 VDD.n9615 VDD.n9614 0.04025
R39867 VDD.n9615 VDD.n9376 0.04025
R39868 VDD.n9619 VDD.n9376 0.04025
R39869 VDD.n9620 VDD.n9619 0.04025
R39870 VDD.n9621 VDD.n9620 0.04025
R39871 VDD.n9621 VDD.n9374 0.04025
R39872 VDD.n9625 VDD.n9374 0.04025
R39873 VDD.n9626 VDD.n9625 0.04025
R39874 VDD.n9627 VDD.n9626 0.04025
R39875 VDD.n9627 VDD.n9372 0.04025
R39876 VDD.n9631 VDD.n9372 0.04025
R39877 VDD.n9632 VDD.n9631 0.04025
R39878 VDD.n9633 VDD.n9632 0.04025
R39879 VDD.n9633 VDD.n9370 0.04025
R39880 VDD.n9637 VDD.n9370 0.04025
R39881 VDD.n9638 VDD.n9637 0.04025
R39882 VDD.n9639 VDD.n9638 0.04025
R39883 VDD.n9639 VDD.n9368 0.04025
R39884 VDD.n9643 VDD.n9368 0.04025
R39885 VDD.n9644 VDD.n9643 0.04025
R39886 VDD.n9645 VDD.n9644 0.04025
R39887 VDD.n9645 VDD.n9366 0.04025
R39888 VDD.n9649 VDD.n9366 0.04025
R39889 VDD.n9650 VDD.n9649 0.04025
R39890 VDD.n9651 VDD.n9650 0.04025
R39891 VDD.n9651 VDD.n9364 0.04025
R39892 VDD.n9655 VDD.n9364 0.04025
R39893 VDD.n9656 VDD.n9655 0.04025
R39894 VDD.n9657 VDD.n9656 0.04025
R39895 VDD.n9657 VDD.n9362 0.04025
R39896 VDD.n9661 VDD.n9362 0.04025
R39897 VDD.n9662 VDD.n9661 0.04025
R39898 VDD.n9663 VDD.n9662 0.04025
R39899 VDD.n9663 VDD.n9360 0.04025
R39900 VDD.n9667 VDD.n9360 0.04025
R39901 VDD.n9668 VDD.n9667 0.04025
R39902 VDD.n9669 VDD.n9668 0.04025
R39903 VDD.n9669 VDD.n9358 0.04025
R39904 VDD.n9673 VDD.n9358 0.04025
R39905 VDD.n9674 VDD.n9673 0.04025
R39906 VDD.n9675 VDD.n9674 0.04025
R39907 VDD.n9675 VDD.n9356 0.04025
R39908 VDD.n9679 VDD.n9356 0.04025
R39909 VDD.n9680 VDD.n9679 0.04025
R39910 VDD.n9681 VDD.n9680 0.04025
R39911 VDD.n9681 VDD.n9354 0.04025
R39912 VDD.n9685 VDD.n9354 0.04025
R39913 VDD.n9686 VDD.n9685 0.04025
R39914 VDD.n9687 VDD.n9686 0.04025
R39915 VDD.n9687 VDD.n9352 0.04025
R39916 VDD.n9691 VDD.n9352 0.04025
R39917 VDD.n9692 VDD.n9691 0.04025
R39918 VDD.n9693 VDD.n9692 0.04025
R39919 VDD.n9693 VDD.n9350 0.04025
R39920 VDD.n9697 VDD.n9350 0.04025
R39921 VDD.n9698 VDD.n9697 0.04025
R39922 VDD.n9699 VDD.n9698 0.04025
R39923 VDD.n9699 VDD.n9348 0.04025
R39924 VDD.n9703 VDD.n9348 0.04025
R39925 VDD.n9704 VDD.n9703 0.04025
R39926 VDD.n9705 VDD.n9704 0.04025
R39927 VDD.n9705 VDD.n9346 0.04025
R39928 VDD.n9709 VDD.n9346 0.04025
R39929 VDD.n9710 VDD.n9709 0.04025
R39930 VDD.n9711 VDD.n9710 0.04025
R39931 VDD.n9711 VDD.n9344 0.04025
R39932 VDD.n9715 VDD.n9344 0.04025
R39933 VDD.n9716 VDD.n9715 0.04025
R39934 VDD.n9717 VDD.n9716 0.04025
R39935 VDD.n9717 VDD.n9342 0.04025
R39936 VDD.n9721 VDD.n9342 0.04025
R39937 VDD.n9722 VDD.n9721 0.04025
R39938 VDD.n9723 VDD.n9722 0.04025
R39939 VDD.n9723 VDD.n9340 0.04025
R39940 VDD.n9727 VDD.n9340 0.04025
R39941 VDD.n9728 VDD.n9727 0.04025
R39942 VDD.n9729 VDD.n9728 0.04025
R39943 VDD.n9729 VDD.n9338 0.04025
R39944 VDD.n9733 VDD.n9338 0.04025
R39945 VDD.n9734 VDD.n9733 0.04025
R39946 VDD.n9735 VDD.n9734 0.04025
R39947 VDD.n9735 VDD.n9336 0.04025
R39948 VDD.n9739 VDD.n9336 0.04025
R39949 VDD.n9740 VDD.n9739 0.04025
R39950 VDD.n9741 VDD.n9740 0.04025
R39951 VDD.n9741 VDD.n9334 0.04025
R39952 VDD.n9745 VDD.n9334 0.04025
R39953 VDD.n9746 VDD.n9745 0.04025
R39954 VDD.n9747 VDD.n9746 0.04025
R39955 VDD.n9747 VDD.n9332 0.04025
R39956 VDD.n9751 VDD.n9332 0.04025
R39957 VDD.n9752 VDD.n9751 0.04025
R39958 VDD.n9753 VDD.n9752 0.04025
R39959 VDD.n9753 VDD.n9330 0.04025
R39960 VDD.n9757 VDD.n9330 0.04025
R39961 VDD.n9758 VDD.n9757 0.04025
R39962 VDD.n9759 VDD.n9758 0.04025
R39963 VDD.n9759 VDD.n9328 0.04025
R39964 VDD.n9763 VDD.n9328 0.04025
R39965 VDD.n9764 VDD.n9763 0.04025
R39966 VDD.n9765 VDD.n9764 0.04025
R39967 VDD.n9765 VDD.n9326 0.04025
R39968 VDD.n9769 VDD.n9326 0.04025
R39969 VDD.n9770 VDD.n9769 0.04025
R39970 VDD.n9771 VDD.n9770 0.04025
R39971 VDD.n9771 VDD.n9324 0.04025
R39972 VDD.n9775 VDD.n9324 0.04025
R39973 VDD.n9776 VDD.n9775 0.04025
R39974 VDD.n9777 VDD.n9776 0.04025
R39975 VDD.n9777 VDD.n9322 0.04025
R39976 VDD.n9781 VDD.n9322 0.04025
R39977 VDD.n9782 VDD.n9781 0.04025
R39978 VDD.n9783 VDD.n9782 0.04025
R39979 VDD.n9783 VDD.n9320 0.04025
R39980 VDD.n9787 VDD.n9320 0.04025
R39981 VDD.n9788 VDD.n9787 0.04025
R39982 VDD.n9789 VDD.n9788 0.04025
R39983 VDD.n9789 VDD.n9318 0.04025
R39984 VDD.n9793 VDD.n9318 0.04025
R39985 VDD.n9794 VDD.n9793 0.04025
R39986 VDD.n9795 VDD.n9794 0.04025
R39987 VDD.n9795 VDD.n9316 0.04025
R39988 VDD.n9799 VDD.n9316 0.04025
R39989 VDD.n9800 VDD.n9799 0.04025
R39990 VDD.n9801 VDD.n9800 0.04025
R39991 VDD.n9801 VDD.n9314 0.04025
R39992 VDD.n9805 VDD.n9314 0.04025
R39993 VDD.n9806 VDD.n9805 0.04025
R39994 VDD.n9807 VDD.n9806 0.04025
R39995 VDD.n9807 VDD.n9312 0.04025
R39996 VDD.n9811 VDD.n9312 0.04025
R39997 VDD.n9812 VDD.n9811 0.04025
R39998 VDD.n9813 VDD.n9812 0.04025
R39999 VDD.n9813 VDD.n9310 0.04025
R40000 VDD.n9817 VDD.n9310 0.04025
R40001 VDD.n9818 VDD.n9817 0.04025
R40002 VDD.n9819 VDD.n9818 0.04025
R40003 VDD.n9819 VDD.n9308 0.04025
R40004 VDD.n9823 VDD.n9308 0.04025
R40005 VDD.n9824 VDD.n9823 0.04025
R40006 VDD.n9825 VDD.n9824 0.04025
R40007 VDD.n9825 VDD.n9306 0.04025
R40008 VDD.n9829 VDD.n9306 0.04025
R40009 VDD.n9830 VDD.n9829 0.04025
R40010 VDD.n9831 VDD.n9830 0.04025
R40011 VDD.n9831 VDD.n9304 0.04025
R40012 VDD.n9835 VDD.n9304 0.04025
R40013 VDD.n9836 VDD.n9835 0.04025
R40014 VDD.n9837 VDD.n9836 0.04025
R40015 VDD.n9837 VDD.n9302 0.04025
R40016 VDD.n9841 VDD.n9302 0.04025
R40017 VDD.n9842 VDD.n9841 0.04025
R40018 VDD.n9843 VDD.n9842 0.04025
R40019 VDD.n9843 VDD.n9300 0.04025
R40020 VDD.n9847 VDD.n9300 0.04025
R40021 VDD.n9848 VDD.n9847 0.04025
R40022 VDD.n9849 VDD.n9848 0.04025
R40023 VDD.n9849 VDD.n9298 0.04025
R40024 VDD.n9853 VDD.n9298 0.04025
R40025 VDD.n9854 VDD.n9853 0.04025
R40026 VDD.n9855 VDD.n9854 0.04025
R40027 VDD.n9855 VDD.n9296 0.04025
R40028 VDD.n9859 VDD.n9296 0.04025
R40029 VDD.n9860 VDD.n9859 0.04025
R40030 VDD.n9861 VDD.n9860 0.04025
R40031 VDD.n9861 VDD.n9294 0.04025
R40032 VDD.n9865 VDD.n9294 0.04025
R40033 VDD.n9866 VDD.n9865 0.04025
R40034 VDD.n9867 VDD.n9866 0.04025
R40035 VDD.n9867 VDD.n9292 0.04025
R40036 VDD.n9871 VDD.n9292 0.04025
R40037 VDD.n9872 VDD.n9871 0.04025
R40038 VDD.n9873 VDD.n9872 0.04025
R40039 VDD.n9873 VDD.n9290 0.04025
R40040 VDD.n9877 VDD.n9290 0.04025
R40041 VDD.n9878 VDD.n9877 0.04025
R40042 VDD.n9879 VDD.n9878 0.04025
R40043 VDD.n9879 VDD.n9288 0.04025
R40044 VDD.n9883 VDD.n9288 0.04025
R40045 VDD.n9884 VDD.n9883 0.04025
R40046 VDD.n9885 VDD.n9884 0.04025
R40047 VDD.n9885 VDD.n9286 0.04025
R40048 VDD.n9889 VDD.n9286 0.04025
R40049 VDD.n9890 VDD.n9889 0.04025
R40050 VDD.n9891 VDD.n9890 0.04025
R40051 VDD.n9891 VDD.n9284 0.04025
R40052 VDD.n9895 VDD.n9284 0.04025
R40053 VDD.n9896 VDD.n9895 0.04025
R40054 VDD.n9897 VDD.n9896 0.04025
R40055 VDD.n9897 VDD.n9282 0.04025
R40056 VDD.n9901 VDD.n9282 0.04025
R40057 VDD.n9902 VDD.n9901 0.04025
R40058 VDD.n9903 VDD.n9902 0.04025
R40059 VDD.n9903 VDD.n9280 0.04025
R40060 VDD.n9907 VDD.n9280 0.04025
R40061 VDD.n9908 VDD.n9907 0.04025
R40062 VDD.n9909 VDD.n9908 0.04025
R40063 VDD.n9909 VDD.n9278 0.04025
R40064 VDD.n9913 VDD.n9278 0.04025
R40065 VDD.n9914 VDD.n9913 0.04025
R40066 VDD.n9915 VDD.n9914 0.04025
R40067 VDD.n9915 VDD.n9276 0.04025
R40068 VDD.n9919 VDD.n9276 0.04025
R40069 VDD.n9920 VDD.n9919 0.04025
R40070 VDD.n9921 VDD.n9920 0.04025
R40071 VDD.n9921 VDD.n9274 0.04025
R40072 VDD.n9925 VDD.n9274 0.04025
R40073 VDD.n9926 VDD.n9925 0.04025
R40074 VDD.n9927 VDD.n9926 0.04025
R40075 VDD.n9927 VDD.n9272 0.04025
R40076 VDD.n9931 VDD.n9272 0.04025
R40077 VDD.n9932 VDD.n9931 0.04025
R40078 VDD.n9933 VDD.n9932 0.04025
R40079 VDD.n9933 VDD.n9270 0.04025
R40080 VDD.n9937 VDD.n9270 0.04025
R40081 VDD.n9938 VDD.n9937 0.04025
R40082 VDD.n9939 VDD.n9938 0.04025
R40083 VDD.n9939 VDD.n9268 0.04025
R40084 VDD.n9943 VDD.n9268 0.04025
R40085 VDD.n9944 VDD.n9943 0.04025
R40086 VDD.n9945 VDD.n9944 0.04025
R40087 VDD.n9945 VDD.n9266 0.04025
R40088 VDD.n9949 VDD.n9266 0.04025
R40089 VDD.n9950 VDD.n9949 0.04025
R40090 VDD.n9951 VDD.n9950 0.04025
R40091 VDD.n9951 VDD.n9264 0.04025
R40092 VDD.n9955 VDD.n9264 0.04025
R40093 VDD.n9956 VDD.n9955 0.04025
R40094 VDD.n9957 VDD.n9956 0.04025
R40095 VDD.n9957 VDD.n9262 0.04025
R40096 VDD.n9961 VDD.n9262 0.04025
R40097 VDD.n9962 VDD.n9961 0.04025
R40098 VDD.n9963 VDD.n9962 0.04025
R40099 VDD.n9963 VDD.n9260 0.04025
R40100 VDD.n9967 VDD.n9260 0.04025
R40101 VDD.n9968 VDD.n9967 0.04025
R40102 VDD.n9969 VDD.n9968 0.04025
R40103 VDD.n9969 VDD.n9258 0.04025
R40104 VDD.n9973 VDD.n9258 0.04025
R40105 VDD.n9974 VDD.n9973 0.04025
R40106 VDD.n9975 VDD.n9974 0.04025
R40107 VDD.n9975 VDD.n9256 0.04025
R40108 VDD.n9979 VDD.n9256 0.04025
R40109 VDD.n9980 VDD.n9979 0.04025
R40110 VDD.n9981 VDD.n9980 0.04025
R40111 VDD.n9981 VDD.n9254 0.04025
R40112 VDD.n9985 VDD.n9254 0.04025
R40113 VDD.n9986 VDD.n9985 0.04025
R40114 VDD.n9987 VDD.n9986 0.04025
R40115 VDD.n9987 VDD.n9252 0.04025
R40116 VDD.n9991 VDD.n9252 0.04025
R40117 VDD.n9992 VDD.n9991 0.04025
R40118 VDD.n9993 VDD.n9992 0.04025
R40119 VDD.n9993 VDD.n9250 0.04025
R40120 VDD.n9997 VDD.n9250 0.04025
R40121 VDD.n9998 VDD.n9997 0.04025
R40122 VDD.n9999 VDD.n9998 0.04025
R40123 VDD.n9999 VDD.n9248 0.04025
R40124 VDD.n10003 VDD.n9248 0.04025
R40125 VDD.n10004 VDD.n10003 0.04025
R40126 VDD.n10005 VDD.n10004 0.04025
R40127 VDD.n10005 VDD.n9246 0.04025
R40128 VDD.n10009 VDD.n9246 0.04025
R40129 VDD.n10010 VDD.n10009 0.04025
R40130 VDD.n10011 VDD.n10010 0.04025
R40131 VDD.n10011 VDD.n9244 0.04025
R40132 VDD.n10015 VDD.n9244 0.04025
R40133 VDD.n10016 VDD.n10015 0.04025
R40134 VDD.n10017 VDD.n10016 0.04025
R40135 VDD.n10017 VDD.n9242 0.04025
R40136 VDD.n10021 VDD.n9242 0.04025
R40137 VDD.n10022 VDD.n10021 0.04025
R40138 VDD.n10023 VDD.n10022 0.04025
R40139 VDD.n10023 VDD.n9240 0.04025
R40140 VDD.n10027 VDD.n9240 0.04025
R40141 VDD.n10028 VDD.n10027 0.04025
R40142 VDD.n10029 VDD.n10028 0.04025
R40143 VDD.n10029 VDD.n9238 0.04025
R40144 VDD.n10033 VDD.n9238 0.04025
R40145 VDD.n10034 VDD.n10033 0.04025
R40146 VDD.n10035 VDD.n10034 0.04025
R40147 VDD.n10035 VDD.n9236 0.04025
R40148 VDD.n10039 VDD.n9236 0.04025
R40149 VDD.n10040 VDD.n10039 0.04025
R40150 VDD.n10041 VDD.n10040 0.04025
R40151 VDD.n10041 VDD.n9234 0.04025
R40152 VDD.n10045 VDD.n9234 0.04025
R40153 VDD.n10046 VDD.n10045 0.04025
R40154 VDD.n10047 VDD.n10046 0.04025
R40155 VDD.n10047 VDD.n9232 0.04025
R40156 VDD.n10051 VDD.n9232 0.04025
R40157 VDD.n10052 VDD.n10051 0.04025
R40158 VDD.n10053 VDD.n10052 0.04025
R40159 VDD.n10053 VDD.n9230 0.04025
R40160 VDD.n10057 VDD.n9230 0.04025
R40161 VDD.n10058 VDD.n10057 0.04025
R40162 VDD.n10059 VDD.n10058 0.04025
R40163 VDD.n10059 VDD.n9228 0.04025
R40164 VDD.n10063 VDD.n9228 0.04025
R40165 VDD.n10064 VDD.n10063 0.04025
R40166 VDD.n10065 VDD.n10064 0.04025
R40167 VDD.n10065 VDD.n9226 0.04025
R40168 VDD.n10069 VDD.n9226 0.04025
R40169 VDD.n10070 VDD.n10069 0.04025
R40170 VDD.n10071 VDD.n10070 0.04025
R40171 VDD.n10071 VDD.n9224 0.04025
R40172 VDD.n10075 VDD.n9224 0.04025
R40173 VDD.n10076 VDD.n10075 0.04025
R40174 VDD.n10077 VDD.n10076 0.04025
R40175 VDD.n10077 VDD.n9222 0.04025
R40176 VDD.n10081 VDD.n9222 0.04025
R40177 VDD.n10082 VDD.n10081 0.04025
R40178 VDD.n10083 VDD.n10082 0.04025
R40179 VDD.n10083 VDD.n9220 0.04025
R40180 VDD.n10087 VDD.n9220 0.04025
R40181 VDD.n10088 VDD.n10087 0.04025
R40182 VDD.n10089 VDD.n10088 0.04025
R40183 VDD.n10089 VDD.n9218 0.04025
R40184 VDD.n10093 VDD.n9218 0.04025
R40185 VDD.n10094 VDD.n10093 0.04025
R40186 VDD.n10095 VDD.n10094 0.04025
R40187 VDD.n10095 VDD.n9216 0.04025
R40188 VDD.n10099 VDD.n9216 0.04025
R40189 VDD.n10100 VDD.n10099 0.04025
R40190 VDD.n10101 VDD.n10100 0.04025
R40191 VDD.n11814 VDD.n11813 0.04025
R40192 VDD.n11815 VDD.n11814 0.04025
R40193 VDD.n11815 VDD.n403 0.04025
R40194 VDD.n11819 VDD.n403 0.04025
R40195 VDD.n11820 VDD.n11819 0.04025
R40196 VDD.n11821 VDD.n11820 0.04025
R40197 VDD.n11821 VDD.n401 0.04025
R40198 VDD.n11825 VDD.n401 0.04025
R40199 VDD.n11826 VDD.n11825 0.04025
R40200 VDD.n11827 VDD.n11826 0.04025
R40201 VDD.n11827 VDD.n399 0.04025
R40202 VDD.n11831 VDD.n399 0.04025
R40203 VDD.n11832 VDD.n11831 0.04025
R40204 VDD.n11833 VDD.n11832 0.04025
R40205 VDD.n11833 VDD.n397 0.04025
R40206 VDD.n11837 VDD.n397 0.04025
R40207 VDD.n11838 VDD.n11837 0.04025
R40208 VDD.n11839 VDD.n11838 0.04025
R40209 VDD.n11839 VDD.n395 0.04025
R40210 VDD.n11843 VDD.n395 0.04025
R40211 VDD.n11844 VDD.n11843 0.04025
R40212 VDD.n11845 VDD.n11844 0.04025
R40213 VDD.n11845 VDD.n393 0.04025
R40214 VDD.n11849 VDD.n393 0.04025
R40215 VDD.n11850 VDD.n11849 0.04025
R40216 VDD.n11851 VDD.n11850 0.04025
R40217 VDD.n11851 VDD.n391 0.04025
R40218 VDD.n11855 VDD.n391 0.04025
R40219 VDD.n11856 VDD.n11855 0.04025
R40220 VDD.n11857 VDD.n11856 0.04025
R40221 VDD.n11857 VDD.n389 0.04025
R40222 VDD.n11861 VDD.n389 0.04025
R40223 VDD.n11862 VDD.n11861 0.04025
R40224 VDD.n11863 VDD.n11862 0.04025
R40225 VDD.n11863 VDD.n387 0.04025
R40226 VDD.n11867 VDD.n387 0.04025
R40227 VDD.n11868 VDD.n11867 0.04025
R40228 VDD.n11869 VDD.n11868 0.04025
R40229 VDD.n11869 VDD.n385 0.04025
R40230 VDD.n11874 VDD.n385 0.04025
R40231 VDD.n11875 VDD.n11874 0.04025
R40232 VDD.n11876 VDD.n11875 0.04025
R40233 VDD.n11876 VDD.n383 0.04025
R40234 VDD.n11880 VDD.n383 0.04025
R40235 VDD.n11881 VDD.n11880 0.04025
R40236 VDD.n11882 VDD.n11881 0.04025
R40237 VDD.n11882 VDD.n381 0.04025
R40238 VDD.n11886 VDD.n381 0.04025
R40239 VDD.n11887 VDD.n11886 0.04025
R40240 VDD.n11888 VDD.n11887 0.04025
R40241 VDD.n11888 VDD.n379 0.04025
R40242 VDD.n11892 VDD.n379 0.04025
R40243 VDD.n11893 VDD.n11892 0.04025
R40244 VDD.n11894 VDD.n11893 0.04025
R40245 VDD.n11894 VDD.n377 0.04025
R40246 VDD.n11898 VDD.n377 0.04025
R40247 VDD.n11899 VDD.n11898 0.04025
R40248 VDD.n11900 VDD.n11899 0.04025
R40249 VDD.n11900 VDD.n375 0.04025
R40250 VDD.n11904 VDD.n375 0.04025
R40251 VDD.n11905 VDD.n11904 0.04025
R40252 VDD.n11906 VDD.n11905 0.04025
R40253 VDD.n11906 VDD.n373 0.04025
R40254 VDD.n11910 VDD.n373 0.04025
R40255 VDD.n11911 VDD.n11910 0.04025
R40256 VDD.n11912 VDD.n11911 0.04025
R40257 VDD.n11912 VDD.n371 0.04025
R40258 VDD.n11916 VDD.n371 0.04025
R40259 VDD.n11917 VDD.n11916 0.04025
R40260 VDD.n11918 VDD.n11917 0.04025
R40261 VDD.n11918 VDD.n369 0.04025
R40262 VDD.n11922 VDD.n369 0.04025
R40263 VDD.n11923 VDD.n11922 0.04025
R40264 VDD.n11924 VDD.n11923 0.04025
R40265 VDD.n11924 VDD.n367 0.04025
R40266 VDD.n11928 VDD.n367 0.04025
R40267 VDD.n11929 VDD.n11928 0.04025
R40268 VDD.n11930 VDD.n11929 0.04025
R40269 VDD.n11930 VDD.n365 0.04025
R40270 VDD.n11934 VDD.n365 0.04025
R40271 VDD.n11935 VDD.n11934 0.04025
R40272 VDD.n11936 VDD.n11935 0.04025
R40273 VDD.n11936 VDD.n363 0.04025
R40274 VDD.n11940 VDD.n363 0.04025
R40275 VDD.n11941 VDD.n11940 0.04025
R40276 VDD.n11942 VDD.n11941 0.04025
R40277 VDD.n11942 VDD.n361 0.04025
R40278 VDD.n11946 VDD.n361 0.04025
R40279 VDD.n11947 VDD.n11946 0.04025
R40280 VDD.n11948 VDD.n11947 0.04025
R40281 VDD.n11948 VDD.n359 0.04025
R40282 VDD.n11952 VDD.n359 0.04025
R40283 VDD.n11953 VDD.n11952 0.04025
R40284 VDD.n11954 VDD.n11953 0.04025
R40285 VDD.n11954 VDD.n357 0.04025
R40286 VDD.n11958 VDD.n357 0.04025
R40287 VDD.n11959 VDD.n11958 0.04025
R40288 VDD.n11960 VDD.n11959 0.04025
R40289 VDD.n11960 VDD.n355 0.04025
R40290 VDD.n11964 VDD.n355 0.04025
R40291 VDD.n11965 VDD.n11964 0.04025
R40292 VDD.n11966 VDD.n11965 0.04025
R40293 VDD.n11966 VDD.n353 0.04025
R40294 VDD.n11970 VDD.n353 0.04025
R40295 VDD.n11971 VDD.n11970 0.04025
R40296 VDD.n11972 VDD.n11971 0.04025
R40297 VDD.n11972 VDD.n351 0.04025
R40298 VDD.n11976 VDD.n351 0.04025
R40299 VDD.n11977 VDD.n11976 0.04025
R40300 VDD.n11978 VDD.n11977 0.04025
R40301 VDD.n11978 VDD.n349 0.04025
R40302 VDD.n11982 VDD.n349 0.04025
R40303 VDD.n11983 VDD.n11982 0.04025
R40304 VDD.n11984 VDD.n11983 0.04025
R40305 VDD.n11984 VDD.n347 0.04025
R40306 VDD.n11988 VDD.n347 0.04025
R40307 VDD.n11989 VDD.n11988 0.04025
R40308 VDD.n11990 VDD.n11989 0.04025
R40309 VDD.n11990 VDD.n345 0.04025
R40310 VDD.n11994 VDD.n345 0.04025
R40311 VDD.n11995 VDD.n11994 0.04025
R40312 VDD.n11996 VDD.n11995 0.04025
R40313 VDD.n11996 VDD.n343 0.04025
R40314 VDD.n12000 VDD.n343 0.04025
R40315 VDD.n12001 VDD.n12000 0.04025
R40316 VDD.n12002 VDD.n12001 0.04025
R40317 VDD.n12002 VDD.n341 0.04025
R40318 VDD.n12006 VDD.n341 0.04025
R40319 VDD.n12007 VDD.n12006 0.04025
R40320 VDD.n12008 VDD.n12007 0.04025
R40321 VDD.n12008 VDD.n339 0.04025
R40322 VDD.n12012 VDD.n339 0.04025
R40323 VDD.n12013 VDD.n12012 0.04025
R40324 VDD.n12014 VDD.n12013 0.04025
R40325 VDD.n12014 VDD.n337 0.04025
R40326 VDD.n12018 VDD.n337 0.04025
R40327 VDD.n12019 VDD.n12018 0.04025
R40328 VDD.n12020 VDD.n12019 0.04025
R40329 VDD.n12020 VDD.n335 0.04025
R40330 VDD.n12024 VDD.n335 0.04025
R40331 VDD.n12025 VDD.n12024 0.04025
R40332 VDD.n12026 VDD.n12025 0.04025
R40333 VDD.n12026 VDD.n333 0.04025
R40334 VDD.n12030 VDD.n333 0.04025
R40335 VDD.n12031 VDD.n12030 0.04025
R40336 VDD.n12032 VDD.n12031 0.04025
R40337 VDD.n12032 VDD.n331 0.04025
R40338 VDD.n12036 VDD.n331 0.04025
R40339 VDD.n12037 VDD.n12036 0.04025
R40340 VDD.n12038 VDD.n12037 0.04025
R40341 VDD.n12038 VDD.n329 0.04025
R40342 VDD.n12042 VDD.n329 0.04025
R40343 VDD.n12043 VDD.n12042 0.04025
R40344 VDD.n12044 VDD.n12043 0.04025
R40345 VDD.n12044 VDD.n327 0.04025
R40346 VDD.n12048 VDD.n327 0.04025
R40347 VDD.n12049 VDD.n12048 0.04025
R40348 VDD.n12050 VDD.n12049 0.04025
R40349 VDD.n12050 VDD.n325 0.04025
R40350 VDD.n12054 VDD.n325 0.04025
R40351 VDD.n12055 VDD.n12054 0.04025
R40352 VDD.n12056 VDD.n12055 0.04025
R40353 VDD.n12056 VDD.n323 0.04025
R40354 VDD.n12060 VDD.n323 0.04025
R40355 VDD.n12061 VDD.n12060 0.04025
R40356 VDD.n12062 VDD.n12061 0.04025
R40357 VDD.n12062 VDD.n321 0.04025
R40358 VDD.n12066 VDD.n321 0.04025
R40359 VDD.n12067 VDD.n12066 0.04025
R40360 VDD.n12068 VDD.n12067 0.04025
R40361 VDD.n12068 VDD.n319 0.04025
R40362 VDD.n12072 VDD.n319 0.04025
R40363 VDD.n12073 VDD.n12072 0.04025
R40364 VDD.n12074 VDD.n12073 0.04025
R40365 VDD.n12074 VDD.n317 0.04025
R40366 VDD.n12078 VDD.n317 0.04025
R40367 VDD.n12079 VDD.n12078 0.04025
R40368 VDD.n12080 VDD.n12079 0.04025
R40369 VDD.n12080 VDD.n315 0.04025
R40370 VDD.n12084 VDD.n315 0.04025
R40371 VDD.n12085 VDD.n12084 0.04025
R40372 VDD.n12086 VDD.n12085 0.04025
R40373 VDD.n12086 VDD.n313 0.04025
R40374 VDD.n12090 VDD.n313 0.04025
R40375 VDD.n12091 VDD.n12090 0.04025
R40376 VDD.n12092 VDD.n12091 0.04025
R40377 VDD.n12092 VDD.n311 0.04025
R40378 VDD.n12096 VDD.n311 0.04025
R40379 VDD.n12097 VDD.n12096 0.04025
R40380 VDD.n12098 VDD.n12097 0.04025
R40381 VDD.n12098 VDD.n309 0.04025
R40382 VDD.n12102 VDD.n309 0.04025
R40383 VDD.n12103 VDD.n12102 0.04025
R40384 VDD.n12104 VDD.n12103 0.04025
R40385 VDD.n12104 VDD.n307 0.04025
R40386 VDD.n12108 VDD.n307 0.04025
R40387 VDD.n12109 VDD.n12108 0.04025
R40388 VDD.n12110 VDD.n12109 0.04025
R40389 VDD.n12110 VDD.n305 0.04025
R40390 VDD.n12114 VDD.n305 0.04025
R40391 VDD.n12115 VDD.n12114 0.04025
R40392 VDD.n12116 VDD.n12115 0.04025
R40393 VDD.n12116 VDD.n303 0.04025
R40394 VDD.n12120 VDD.n303 0.04025
R40395 VDD.n12121 VDD.n12120 0.04025
R40396 VDD.n12122 VDD.n12121 0.04025
R40397 VDD.n12122 VDD.n301 0.04025
R40398 VDD.n12126 VDD.n301 0.04025
R40399 VDD.n12127 VDD.n12126 0.04025
R40400 VDD.n12128 VDD.n12127 0.04025
R40401 VDD.n12128 VDD.n299 0.04025
R40402 VDD.n12132 VDD.n299 0.04025
R40403 VDD.n12133 VDD.n12132 0.04025
R40404 VDD.n12134 VDD.n12133 0.04025
R40405 VDD.n12134 VDD.n297 0.04025
R40406 VDD.n12138 VDD.n297 0.04025
R40407 VDD.n12139 VDD.n12138 0.04025
R40408 VDD.n12140 VDD.n12139 0.04025
R40409 VDD.n12140 VDD.n295 0.04025
R40410 VDD.n12144 VDD.n295 0.04025
R40411 VDD.n12145 VDD.n12144 0.04025
R40412 VDD.n12146 VDD.n12145 0.04025
R40413 VDD.n12146 VDD.n293 0.04025
R40414 VDD.n12150 VDD.n293 0.04025
R40415 VDD.n12151 VDD.n12150 0.04025
R40416 VDD.n12152 VDD.n12151 0.04025
R40417 VDD.n12152 VDD.n291 0.04025
R40418 VDD.n12156 VDD.n291 0.04025
R40419 VDD.n12157 VDD.n12156 0.04025
R40420 VDD.n12158 VDD.n12157 0.04025
R40421 VDD.n12158 VDD.n289 0.04025
R40422 VDD.n12162 VDD.n289 0.04025
R40423 VDD.n12163 VDD.n12162 0.04025
R40424 VDD.n12164 VDD.n12163 0.04025
R40425 VDD.n12164 VDD.n287 0.04025
R40426 VDD.n12168 VDD.n287 0.04025
R40427 VDD.n12169 VDD.n12168 0.04025
R40428 VDD.n12170 VDD.n12169 0.04025
R40429 VDD.n12170 VDD.n285 0.04025
R40430 VDD.n12174 VDD.n285 0.04025
R40431 VDD.n12175 VDD.n12174 0.04025
R40432 VDD.n12176 VDD.n12175 0.04025
R40433 VDD.n12176 VDD.n283 0.04025
R40434 VDD.n12180 VDD.n283 0.04025
R40435 VDD.n12181 VDD.n12180 0.04025
R40436 VDD.n12182 VDD.n12181 0.04025
R40437 VDD.n12182 VDD.n281 0.04025
R40438 VDD.n12186 VDD.n281 0.04025
R40439 VDD.n12187 VDD.n12186 0.04025
R40440 VDD.n12188 VDD.n12187 0.04025
R40441 VDD.n12188 VDD.n279 0.04025
R40442 VDD.n12192 VDD.n279 0.04025
R40443 VDD.n12193 VDD.n12192 0.04025
R40444 VDD.n12194 VDD.n12193 0.04025
R40445 VDD.n12194 VDD.n277 0.04025
R40446 VDD.n12198 VDD.n277 0.04025
R40447 VDD.n12199 VDD.n12198 0.04025
R40448 VDD.n12200 VDD.n12199 0.04025
R40449 VDD.n12200 VDD.n275 0.04025
R40450 VDD.n12204 VDD.n275 0.04025
R40451 VDD.n12205 VDD.n12204 0.04025
R40452 VDD.n12206 VDD.n12205 0.04025
R40453 VDD.n12206 VDD.n273 0.04025
R40454 VDD.n12210 VDD.n273 0.04025
R40455 VDD.n12211 VDD.n12210 0.04025
R40456 VDD.n12212 VDD.n12211 0.04025
R40457 VDD.n12212 VDD.n271 0.04025
R40458 VDD.n12216 VDD.n271 0.04025
R40459 VDD.n12217 VDD.n12216 0.04025
R40460 VDD.n12218 VDD.n12217 0.04025
R40461 VDD.n12218 VDD.n269 0.04025
R40462 VDD.n12222 VDD.n269 0.04025
R40463 VDD.n12223 VDD.n12222 0.04025
R40464 VDD.n12224 VDD.n12223 0.04025
R40465 VDD.n12224 VDD.n267 0.04025
R40466 VDD.n12228 VDD.n267 0.04025
R40467 VDD.n12229 VDD.n12228 0.04025
R40468 VDD.n12230 VDD.n12229 0.04025
R40469 VDD.n12230 VDD.n265 0.04025
R40470 VDD.n12234 VDD.n265 0.04025
R40471 VDD.n12235 VDD.n12234 0.04025
R40472 VDD.n12236 VDD.n12235 0.04025
R40473 VDD.n12236 VDD.n263 0.04025
R40474 VDD.n12240 VDD.n263 0.04025
R40475 VDD.n12241 VDD.n12240 0.04025
R40476 VDD.n12242 VDD.n12241 0.04025
R40477 VDD.n12242 VDD.n261 0.04025
R40478 VDD.n12246 VDD.n261 0.04025
R40479 VDD.n12247 VDD.n12246 0.04025
R40480 VDD.n12248 VDD.n12247 0.04025
R40481 VDD.n12248 VDD.n259 0.04025
R40482 VDD.n12252 VDD.n259 0.04025
R40483 VDD.n12253 VDD.n12252 0.04025
R40484 VDD.n12254 VDD.n12253 0.04025
R40485 VDD.n12254 VDD.n257 0.04025
R40486 VDD.n12258 VDD.n257 0.04025
R40487 VDD.n12259 VDD.n12258 0.04025
R40488 VDD.n12260 VDD.n12259 0.04025
R40489 VDD.n12260 VDD.n255 0.04025
R40490 VDD.n12264 VDD.n255 0.04025
R40491 VDD.n12265 VDD.n12264 0.04025
R40492 VDD.n12266 VDD.n12265 0.04025
R40493 VDD.n12266 VDD.n253 0.04025
R40494 VDD.n12270 VDD.n253 0.04025
R40495 VDD.n12271 VDD.n12270 0.04025
R40496 VDD.n12272 VDD.n12271 0.04025
R40497 VDD.n12272 VDD.n251 0.04025
R40498 VDD.n12276 VDD.n251 0.04025
R40499 VDD.n12277 VDD.n12276 0.04025
R40500 VDD.n12278 VDD.n12277 0.04025
R40501 VDD.n12278 VDD.n249 0.04025
R40502 VDD.n12282 VDD.n249 0.04025
R40503 VDD.n12283 VDD.n12282 0.04025
R40504 VDD.n12284 VDD.n12283 0.04025
R40505 VDD.n12284 VDD.n247 0.04025
R40506 VDD.n12288 VDD.n247 0.04025
R40507 VDD.n12289 VDD.n12288 0.04025
R40508 VDD.n12290 VDD.n12289 0.04025
R40509 VDD.n12290 VDD.n245 0.04025
R40510 VDD.n12294 VDD.n245 0.04025
R40511 VDD.n12295 VDD.n12294 0.04025
R40512 VDD.n12296 VDD.n12295 0.04025
R40513 VDD.n12296 VDD.n243 0.04025
R40514 VDD.n12300 VDD.n243 0.04025
R40515 VDD.n12301 VDD.n12300 0.04025
R40516 VDD.n12302 VDD.n12301 0.04025
R40517 VDD.n12302 VDD.n241 0.04025
R40518 VDD.n12306 VDD.n241 0.04025
R40519 VDD.n12307 VDD.n12306 0.04025
R40520 VDD.n12308 VDD.n12307 0.04025
R40521 VDD.n12308 VDD.n239 0.04025
R40522 VDD.n12312 VDD.n239 0.04025
R40523 VDD.n12313 VDD.n12312 0.04025
R40524 VDD.n12314 VDD.n12313 0.04025
R40525 VDD.n12314 VDD.n237 0.04025
R40526 VDD.n12318 VDD.n237 0.04025
R40527 VDD.n12319 VDD.n12318 0.04025
R40528 VDD.n12320 VDD.n12319 0.04025
R40529 VDD.n12320 VDD.n235 0.04025
R40530 VDD.n12324 VDD.n235 0.04025
R40531 VDD.n12325 VDD.n12324 0.04025
R40532 VDD.n12326 VDD.n12325 0.04025
R40533 VDD.n12326 VDD.n233 0.04025
R40534 VDD.n12330 VDD.n233 0.04025
R40535 VDD.n12331 VDD.n12330 0.04025
R40536 VDD.n12332 VDD.n12331 0.04025
R40537 VDD.n12332 VDD.n231 0.04025
R40538 VDD.n12336 VDD.n231 0.04025
R40539 VDD.n12337 VDD.n12336 0.04025
R40540 VDD.n12338 VDD.n12337 0.04025
R40541 VDD.n12338 VDD.n229 0.04025
R40542 VDD.n12342 VDD.n229 0.04025
R40543 VDD.n12343 VDD.n12342 0.04025
R40544 VDD.n12344 VDD.n12343 0.04025
R40545 VDD.n12344 VDD.n227 0.04025
R40546 VDD.n12348 VDD.n227 0.04025
R40547 VDD.n12349 VDD.n12348 0.04025
R40548 VDD.n12350 VDD.n12349 0.04025
R40549 VDD.n12350 VDD.n225 0.04025
R40550 VDD.n12354 VDD.n225 0.04025
R40551 VDD.n12355 VDD.n12354 0.04025
R40552 VDD.n12356 VDD.n12355 0.04025
R40553 VDD.n12356 VDD.n223 0.04025
R40554 VDD.n12360 VDD.n223 0.04025
R40555 VDD.n12361 VDD.n12360 0.04025
R40556 VDD.n12362 VDD.n12361 0.04025
R40557 VDD.n12362 VDD.n221 0.04025
R40558 VDD.n12366 VDD.n221 0.04025
R40559 VDD.n12367 VDD.n12366 0.04025
R40560 VDD.n12368 VDD.n12367 0.04025
R40561 VDD.n12368 VDD.n219 0.04025
R40562 VDD.n12372 VDD.n219 0.04025
R40563 VDD.n12373 VDD.n12372 0.04025
R40564 VDD.n12374 VDD.n12373 0.04025
R40565 VDD.n12374 VDD.n217 0.04025
R40566 VDD.n12378 VDD.n217 0.04025
R40567 VDD.n12379 VDD.n12378 0.04025
R40568 VDD.n12380 VDD.n12379 0.04025
R40569 VDD.n12380 VDD.n215 0.04025
R40570 VDD.n12384 VDD.n215 0.04025
R40571 VDD.n12385 VDD.n12384 0.04025
R40572 VDD.n12386 VDD.n12385 0.04025
R40573 VDD.n12386 VDD.n213 0.04025
R40574 VDD.n12390 VDD.n213 0.04025
R40575 VDD.n12391 VDD.n12390 0.04025
R40576 VDD.n12392 VDD.n12391 0.04025
R40577 VDD.n12392 VDD.n211 0.04025
R40578 VDD.n12396 VDD.n211 0.04025
R40579 VDD.n12397 VDD.n12396 0.04025
R40580 VDD.n12398 VDD.n12397 0.04025
R40581 VDD.n12398 VDD.n209 0.04025
R40582 VDD.n12402 VDD.n209 0.04025
R40583 VDD.n12403 VDD.n12402 0.04025
R40584 VDD.n12404 VDD.n12403 0.04025
R40585 VDD.n12404 VDD.n207 0.04025
R40586 VDD.n12408 VDD.n207 0.04025
R40587 VDD.n12409 VDD.n12408 0.04025
R40588 VDD.n12410 VDD.n12409 0.04025
R40589 VDD.n12410 VDD.n205 0.04025
R40590 VDD.n12414 VDD.n205 0.04025
R40591 VDD.n12415 VDD.n12414 0.04025
R40592 VDD.n12416 VDD.n12415 0.04025
R40593 VDD.n12416 VDD.n203 0.04025
R40594 VDD.n12420 VDD.n203 0.04025
R40595 VDD.n12421 VDD.n12420 0.04025
R40596 VDD.n12422 VDD.n12421 0.04025
R40597 VDD.n12422 VDD.n201 0.04025
R40598 VDD.n12426 VDD.n201 0.04025
R40599 VDD.n12427 VDD.n12426 0.04025
R40600 VDD.n12428 VDD.n12427 0.04025
R40601 VDD.n12428 VDD.n199 0.04025
R40602 VDD.n12432 VDD.n199 0.04025
R40603 VDD.n12433 VDD.n12432 0.04025
R40604 VDD.n12434 VDD.n12433 0.04025
R40605 VDD.n12434 VDD.n197 0.04025
R40606 VDD.n12438 VDD.n197 0.04025
R40607 VDD.n12439 VDD.n12438 0.04025
R40608 VDD.n12440 VDD.n12439 0.04025
R40609 VDD.n7843 VDD.n7842 0.0395167
R40610 VDD.n2173 VDD.n2172 0.0394276
R40611 VDD.n6875 VDD.n2390 0.0392688
R40612 VDD.n8052 VDD.n8051 0.0387235
R40613 VDD.n8048 VDD.n8047 0.0383
R40614 VDD.n9137 VDD.n9136 0.0382419
R40615 VDD.n9126 VDD.n9125 0.0382419
R40616 VDD.n12565 VDD.n12563 0.0382419
R40617 VDD.n12577 VDD.n12576 0.0382419
R40618 VDD.n10148 VDD.n10147 0.037625
R40619 VDD.n8052 VDD.n2148 0.0373471
R40620 VDD.n7942 VDD.n7854 0.0371353
R40621 VDD.n1564 VDD.n1563 0.0370902
R40622 VDD.n1542 VDD.n1541 0.0370902
R40623 VDD.n1640 VDD.n771 0.0370902
R40624 VDD.n1529 VDD.n1528 0.0370902
R40625 VDD.n7912 VDD.n7911 0.0369637
R40626 VDD.n7943 VDD.n7942 0.0369235
R40627 VDD.n7912 VDD.n7863 0.0367529
R40628 VDD.n12567 VDD.n12566 0.0364748
R40629 VDD.n12574 VDD.n12573 0.0364748
R40630 VDD.n9184 VDD.n9183 0.0363759
R40631 VDD.n5369 VDD.n5368 0.0360345
R40632 VDD.n6372 VDD.n5375 0.0360345
R40633 VDD.n6368 VDD.n6367 0.0360345
R40634 VDD.n5944 VDD.n5943 0.0360345
R40635 VDD.n2366 VDD.n2365 0.0360345
R40636 VDD.n7135 VDD.n2316 0.0360345
R40637 VDD.n7131 VDD.n7130 0.0360345
R40638 VDD.n7044 VDD.n7043 0.0360345
R40639 VDD.n7864 VDD.n2146 0.0359624
R40640 VDD.n12641 VDD.n12638 0.0359286
R40641 VDD.n1003 VDD.n957 0.0359286
R40642 VDD.n1755 VDD.n1754 0.0359286
R40643 VDD.n9135 VDD.n9134 0.0357174
R40644 VDD.n6024 VDD.n5299 0.0347688
R40645 VDD.n6174 VDD.n6171 0.0347688
R40646 VDD.n6412 VDD.n5299 0.0347688
R40647 VDD.n8011 VDD.n8010 0.0347688
R40648 VDD.n2403 VDD.n2402 0.0347688
R40649 VDD.n2402 VDD.n2396 0.0347688
R40650 VDD.n8133 VDD.n8132 0.0346711
R40651 VDD.n8134 VDD.n8133 0.0346711
R40652 VDD.n8134 VDD.n2090 0.0346711
R40653 VDD.n8136 VDD.n2090 0.0346711
R40654 VDD.n8139 VDD.n8138 0.0346711
R40655 VDD.n8162 VDD.n8139 0.0346711
R40656 VDD.n8112 VDD.n8111 0.0346711
R40657 VDD.n8113 VDD.n8112 0.0346711
R40658 VDD.n8113 VDD.n2092 0.0346711
R40659 VDD.n8115 VDD.n2092 0.0346711
R40660 VDD.n8118 VDD.n8117 0.0346711
R40661 VDD.n8119 VDD.n8118 0.0346711
R40662 VDD.n8119 VDD.n2091 0.0346711
R40663 VDD.n8121 VDD.n2091 0.0346711
R40664 VDD.n8100 VDD.n8099 0.0346711
R40665 VDD.n8101 VDD.n8100 0.0346711
R40666 VDD.n8101 VDD.n2103 0.0346711
R40667 VDD.n8103 VDD.n2103 0.0346711
R40668 VDD.n8106 VDD.n8105 0.0346711
R40669 VDD.n8107 VDD.n8106 0.0346711
R40670 VDD.n8107 VDD.n2102 0.0346711
R40671 VDD.n8109 VDD.n2102 0.0346711
R40672 VDD.n5584 VDD.n5551 0.0346711
R40673 VDD.n5582 VDD.n5551 0.0346711
R40674 VDD.n5582 VDD.n5581 0.0346711
R40675 VDD.n5581 VDD.n5580 0.0346711
R40676 VDD.n5578 VDD.n5552 0.0346711
R40677 VDD.n5576 VDD.n5552 0.0346711
R40678 VDD.n5605 VDD.n5549 0.0346711
R40679 VDD.n5603 VDD.n5549 0.0346711
R40680 VDD.n5603 VDD.n5602 0.0346711
R40681 VDD.n5602 VDD.n5601 0.0346711
R40682 VDD.n5599 VDD.n5550 0.0346711
R40683 VDD.n5597 VDD.n5550 0.0346711
R40684 VDD.n5597 VDD.n5596 0.0346711
R40685 VDD.n5596 VDD.n5595 0.0346711
R40686 VDD.n5626 VDD.n5547 0.0346711
R40687 VDD.n5624 VDD.n5547 0.0346711
R40688 VDD.n5624 VDD.n5623 0.0346711
R40689 VDD.n5623 VDD.n5622 0.0346711
R40690 VDD.n5620 VDD.n5548 0.0346711
R40691 VDD.n5618 VDD.n5548 0.0346711
R40692 VDD.n5618 VDD.n5617 0.0346711
R40693 VDD.n5617 VDD.n5616 0.0346711
R40694 VDD.n5666 VDD.n5542 0.0346711
R40695 VDD.n5664 VDD.n5542 0.0346711
R40696 VDD.n5664 VDD.n5663 0.0346711
R40697 VDD.n5663 VDD.n5662 0.0346711
R40698 VDD.n5660 VDD.n5543 0.0346711
R40699 VDD.n5658 VDD.n5543 0.0346711
R40700 VDD.n5867 VDD.n5866 0.0346711
R40701 VDD.n5868 VDD.n5867 0.0346711
R40702 VDD.n5868 VDD.n5668 0.0346711
R40703 VDD.n5870 VDD.n5668 0.0346711
R40704 VDD.n5873 VDD.n5872 0.0346711
R40705 VDD.n5874 VDD.n5873 0.0346711
R40706 VDD.n5874 VDD.n5667 0.0346711
R40707 VDD.n5876 VDD.n5667 0.0346711
R40708 VDD.n5855 VDD.n5854 0.0346711
R40709 VDD.n5856 VDD.n5855 0.0346711
R40710 VDD.n5856 VDD.n5679 0.0346711
R40711 VDD.n5858 VDD.n5679 0.0346711
R40712 VDD.n5861 VDD.n5860 0.0346711
R40713 VDD.n5862 VDD.n5861 0.0346711
R40714 VDD.n5862 VDD.n5678 0.0346711
R40715 VDD.n5864 VDD.n5678 0.0346711
R40716 VDD.n5812 VDD.n5811 0.0346711
R40717 VDD.n5813 VDD.n5812 0.0346711
R40718 VDD.n5813 VDD.n5681 0.0346711
R40719 VDD.n5815 VDD.n5681 0.0346711
R40720 VDD.n5818 VDD.n5817 0.0346711
R40721 VDD.n5841 VDD.n5818 0.0346711
R40722 VDD.n5800 VDD.n5799 0.0346711
R40723 VDD.n5801 VDD.n5800 0.0346711
R40724 VDD.n5801 VDD.n5692 0.0346711
R40725 VDD.n5803 VDD.n5692 0.0346711
R40726 VDD.n5806 VDD.n5805 0.0346711
R40727 VDD.n5807 VDD.n5806 0.0346711
R40728 VDD.n5807 VDD.n5691 0.0346711
R40729 VDD.n5809 VDD.n5691 0.0346711
R40730 VDD.n5779 VDD.n5778 0.0346711
R40731 VDD.n5780 VDD.n5779 0.0346711
R40732 VDD.n5780 VDD.n5694 0.0346711
R40733 VDD.n5782 VDD.n5694 0.0346711
R40734 VDD.n5785 VDD.n5784 0.0346711
R40735 VDD.n5786 VDD.n5785 0.0346711
R40736 VDD.n5786 VDD.n5693 0.0346711
R40737 VDD.n5788 VDD.n5693 0.0346711
R40738 VDD.n5745 VDD.n5744 0.0346711
R40739 VDD.n5746 VDD.n5745 0.0346711
R40740 VDD.n5746 VDD.n5705 0.0346711
R40741 VDD.n5748 VDD.n5705 0.0346711
R40742 VDD.n5751 VDD.n5750 0.0346711
R40743 VDD.n5774 VDD.n5751 0.0346711
R40744 VDD.n5724 VDD.n5723 0.0346711
R40745 VDD.n5725 VDD.n5724 0.0346711
R40746 VDD.n5725 VDD.n5707 0.0346711
R40747 VDD.n5727 VDD.n5707 0.0346711
R40748 VDD.n5730 VDD.n5729 0.0346711
R40749 VDD.n5731 VDD.n5730 0.0346711
R40750 VDD.n5731 VDD.n5706 0.0346711
R40751 VDD.n5733 VDD.n5706 0.0346711
R40752 VDD.n11036 VDD.n1769 0.0346711
R40753 VDD.n11034 VDD.n1769 0.0346711
R40754 VDD.n11034 VDD.n11033 0.0346711
R40755 VDD.n11033 VDD.n11032 0.0346711
R40756 VDD.n5718 VDD.n1770 0.0346711
R40757 VDD.n5719 VDD.n5718 0.0346711
R40758 VDD.n5719 VDD.n5717 0.0346711
R40759 VDD.n5721 VDD.n5717 0.0346711
R40760 VDD.n8975 VDD.n8971 0.0346711
R40761 VDD.n8973 VDD.n8971 0.0346711
R40762 VDD.n8973 VDD.n8972 0.0346711
R40763 VDD.n8972 VDD.n8490 0.0346711
R40764 VDD.n9039 VDD.n9038 0.0346711
R40765 VDD.n9040 VDD.n9039 0.0346711
R40766 VDD.n9040 VDD.n8489 0.0346711
R40767 VDD.n9042 VDD.n8489 0.0346711
R40768 VDD.n8948 VDD.n8947 0.0346711
R40769 VDD.n8949 VDD.n8948 0.0346711
R40770 VDD.n8949 VDD.n8502 0.0346711
R40771 VDD.n8951 VDD.n8502 0.0346711
R40772 VDD.n9007 VDD.n8952 0.0346711
R40773 VDD.n9005 VDD.n8952 0.0346711
R40774 VDD.n8848 VDD.n8844 0.0346711
R40775 VDD.n8846 VDD.n8844 0.0346711
R40776 VDD.n8846 VDD.n8845 0.0346711
R40777 VDD.n8845 VDD.n8507 0.0346711
R40778 VDD.n8942 VDD.n8941 0.0346711
R40779 VDD.n8943 VDD.n8942 0.0346711
R40780 VDD.n8943 VDD.n8506 0.0346711
R40781 VDD.n8945 VDD.n8506 0.0346711
R40782 VDD.n8839 VDD.n8838 0.0346711
R40783 VDD.n8840 VDD.n8839 0.0346711
R40784 VDD.n8840 VDD.n8521 0.0346711
R40785 VDD.n8842 VDD.n8521 0.0346711
R40786 VDD.n8876 VDD.n8843 0.0346711
R40787 VDD.n8874 VDD.n8843 0.0346711
R40788 VDD.n8874 VDD.n8873 0.0346711
R40789 VDD.n8873 VDD.n8872 0.0346711
R40790 VDD.n8547 VDD.n8543 0.0346711
R40791 VDD.n8545 VDD.n8543 0.0346711
R40792 VDD.n8545 VDD.n8544 0.0346711
R40793 VDD.n8544 VDD.n8526 0.0346711
R40794 VDD.n8811 VDD.n8810 0.0346711
R40795 VDD.n8834 VDD.n8811 0.0346711
R40796 VDD.n8550 VDD.n184 0.0346711
R40797 VDD.n8551 VDD.n8550 0.0346711
R40798 VDD.n8551 VDD.n8549 0.0346711
R40799 VDD.n8553 VDD.n8549 0.0346711
R40800 VDD.n8556 VDD.n8555 0.0346711
R40801 VDD.n8557 VDD.n8556 0.0346711
R40802 VDD.n8557 VDD.n8548 0.0346711
R40803 VDD.n8559 VDD.n8548 0.0346711
R40804 VDD.n171 VDD.n170 0.0346711
R40805 VDD.n172 VDD.n171 0.0346711
R40806 VDD.n172 VDD.n125 0.0346711
R40807 VDD.n174 VDD.n125 0.0346711
R40808 VDD.n187 VDD.n186 0.0346711
R40809 VDD.n188 VDD.n187 0.0346711
R40810 VDD.n188 VDD.n185 0.0346711
R40811 VDD.n190 VDD.n185 0.0346711
R40812 VDD.n9092 VDD.n8470 0.0346711
R40813 VDD.n9093 VDD.n9092 0.0346711
R40814 VDD.n9093 VDD.n9091 0.0346711
R40815 VDD.n9095 VDD.n9091 0.0346711
R40816 VDD.n9098 VDD.n9097 0.0346711
R40817 VDD.n9121 VDD.n9098 0.0346711
R40818 VDD.n8488 VDD.n8484 0.0346711
R40819 VDD.n8486 VDD.n8484 0.0346711
R40820 VDD.n8486 VDD.n8485 0.0346711
R40821 VDD.n8485 VDD.n8472 0.0346711
R40822 VDD.n9163 VDD.n9162 0.0346711
R40823 VDD.n9164 VDD.n9163 0.0346711
R40824 VDD.n9164 VDD.n8471 0.0346711
R40825 VDD.n9166 VDD.n8471 0.0346711
R40826 VDD.n137 VDD.n106 0.0346711
R40827 VDD.n138 VDD.n137 0.0346711
R40828 VDD.n138 VDD.n136 0.0346711
R40829 VDD.n140 VDD.n136 0.0346711
R40830 VDD.n143 VDD.n142 0.0346711
R40831 VDD.n166 VDD.n143 0.0346711
R40832 VDD.n12498 VDD.n104 0.0346711
R40833 VDD.n12496 VDD.n104 0.0346711
R40834 VDD.n12496 VDD.n12495 0.0346711
R40835 VDD.n12495 VDD.n12494 0.0346711
R40836 VDD.n12492 VDD.n105 0.0346711
R40837 VDD.n12490 VDD.n105 0.0346711
R40838 VDD.n12490 VDD.n12489 0.0346711
R40839 VDD.n12489 VDD.n12488 0.0346711
R40840 VDD.n91 VDD.n90 0.0346711
R40841 VDD.n92 VDD.n91 0.0346711
R40842 VDD.n92 VDD.n45 0.0346711
R40843 VDD.n94 VDD.n45 0.0346711
R40844 VDD.n12501 VDD.n12500 0.0346711
R40845 VDD.n12502 VDD.n12501 0.0346711
R40846 VDD.n12502 VDD.n12499 0.0346711
R40847 VDD.n12504 VDD.n12499 0.0346711
R40848 VDD.n48 VDD.n26 0.0346711
R40849 VDD.n49 VDD.n48 0.0346711
R40850 VDD.n49 VDD.n47 0.0346711
R40851 VDD.n51 VDD.n47 0.0346711
R40852 VDD.n54 VDD.n53 0.0346711
R40853 VDD.n77 VDD.n54 0.0346711
R40854 VDD.n12554 VDD.n24 0.0346711
R40855 VDD.n12552 VDD.n24 0.0346711
R40856 VDD.n12552 VDD.n12551 0.0346711
R40857 VDD.n12551 VDD.n12550 0.0346711
R40858 VDD.n12548 VDD.n25 0.0346711
R40859 VDD.n12546 VDD.n25 0.0346711
R40860 VDD.n12546 VDD.n12545 0.0346711
R40861 VDD.n12545 VDD.n12544 0.0346711
R40862 VDD.n12588 VDD.n12587 0.0346711
R40863 VDD.n12589 VDD.n12588 0.0346711
R40864 VDD.n12589 VDD.n12556 0.0346711
R40865 VDD.n12591 VDD.n12556 0.0346711
R40866 VDD.n12595 VDD.n12594 0.0346711
R40867 VDD.n12596 VDD.n12595 0.0346711
R40868 VDD.n12596 VDD.n12555 0.0346711
R40869 VDD.n12598 VDD.n12555 0.0346711
R40870 VDD.n12580 VDD.n12579 0.0345
R40871 VDD.n11129 VDD.n638 0.0345
R40872 VDD.n1763 VDD.n674 0.0345
R40873 VDD.n6325 VDD.n6324 0.0345
R40874 VDD.n6014 VDD.n6011 0.0345
R40875 VDD.n5538 VDD.n5537 0.0345
R40876 VDD.n5886 VDD.n5880 0.0345
R40877 VDD.n5911 VDD.n5910 0.0345
R40878 VDD.n8088 VDD.n1996 0.0345
R40879 VDD.n8090 VDD.n2118 0.0345
R40880 VDD.n12632 VDD.n12631 0.0345
R40881 VDD.n12635 VDD.n3 0.0345
R40882 VDD.n1000 VDD.n953 0.0345
R40883 VDD.n1760 VDD.n1759 0.0345
R40884 VDD.n6024 VDD.n6022 0.0341759
R40885 VDD.n6036 VDD.n6023 0.0341759
R40886 VDD.n6033 VDD.n6023 0.0341759
R40887 VDD.n6033 VDD.n6032 0.0341759
R40888 VDD.n6032 VDD.n6031 0.0341759
R40889 VDD.n6031 VDD.n6025 0.0341759
R40890 VDD.n6029 VDD.n6025 0.0341759
R40891 VDD.n6028 VDD.n6026 0.0341759
R40892 VDD.n6026 VDD.n5283 0.0341759
R40893 VDD.n6574 VDD.n6573 0.0341759
R40894 VDD.n6573 VDD.n5284 0.0341759
R40895 VDD.n6571 VDD.n5284 0.0341759
R40896 VDD.n6570 VDD.n5285 0.0341759
R40897 VDD.n6568 VDD.n5285 0.0341759
R40898 VDD.n6568 VDD.n6567 0.0341759
R40899 VDD.n6567 VDD.n6566 0.0341759
R40900 VDD.n6566 VDD.n5286 0.0341759
R40901 VDD.n6563 VDD.n5286 0.0341759
R40902 VDD.n6171 VDD.n6018 0.0341759
R40903 VDD.n6169 VDD.n6168 0.0341759
R40904 VDD.n6168 VDD.n6167 0.0341759
R40905 VDD.n6167 VDD.n6158 0.0341759
R40906 VDD.n6164 VDD.n6158 0.0341759
R40907 VDD.n6164 VDD.n6163 0.0341759
R40908 VDD.n6163 VDD.n6162 0.0341759
R40909 VDD.n6161 VDD.n6159 0.0341759
R40910 VDD.n6159 VDD.n5302 0.0341759
R40911 VDD.n6400 VDD.n6399 0.0341759
R40912 VDD.n6400 VDD.n5301 0.0341759
R40913 VDD.n6402 VDD.n5301 0.0341759
R40914 VDD.n6404 VDD.n6403 0.0341759
R40915 VDD.n6405 VDD.n6404 0.0341759
R40916 VDD.n6405 VDD.n5300 0.0341759
R40917 VDD.n6408 VDD.n5300 0.0341759
R40918 VDD.n6409 VDD.n6408 0.0341759
R40919 VDD.n6410 VDD.n6409 0.0341759
R40920 VDD.n8010 VDD.n2166 0.0341759
R40921 VDD.n8008 VDD.n2166 0.0341759
R40922 VDD.n8008 VDD.n8007 0.0341759
R40923 VDD.n8007 VDD.n8006 0.0341759
R40924 VDD.n8006 VDD.n2167 0.0341759
R40925 VDD.n8003 VDD.n2167 0.0341759
R40926 VDD.n8003 VDD.n8002 0.0341759
R40927 VDD.n8002 VDD.n8001 0.0341759
R40928 VDD.n8000 VDD.n2168 0.0341759
R40929 VDD.n7998 VDD.n2168 0.0341759
R40930 VDD.n2186 VDD.n2185 0.0341759
R40931 VDD.n2185 VDD.n2169 0.0341759
R40932 VDD.n2183 VDD.n2169 0.0341759
R40933 VDD.n2182 VDD.n2170 0.0341759
R40934 VDD.n2180 VDD.n2170 0.0341759
R40935 VDD.n2180 VDD.n2179 0.0341759
R40936 VDD.n2179 VDD.n2178 0.0341759
R40937 VDD.n2178 VDD.n2171 0.0341759
R40938 VDD.n2175 VDD.n2171 0.0341759
R40939 VDD.n2175 VDD.n2174 0.0341759
R40940 VDD.n2174 VDD.n2173 0.0341759
R40941 VDD.n2404 VDD.n2403 0.0341759
R40942 VDD.n6850 VDD.n2395 0.0341759
R40943 VDD.n6853 VDD.n2395 0.0341759
R40944 VDD.n6854 VDD.n6853 0.0341759
R40945 VDD.n6855 VDD.n6854 0.0341759
R40946 VDD.n6855 VDD.n2394 0.0341759
R40947 VDD.n6857 VDD.n2394 0.0341759
R40948 VDD.n6858 VDD.n2393 0.0341759
R40949 VDD.n6860 VDD.n2393 0.0341759
R40950 VDD.n6863 VDD.n6862 0.0341759
R40951 VDD.n6863 VDD.n2392 0.0341759
R40952 VDD.n6865 VDD.n2392 0.0341759
R40953 VDD.n6867 VDD.n6866 0.0341759
R40954 VDD.n6868 VDD.n6867 0.0341759
R40955 VDD.n6868 VDD.n2391 0.0341759
R40956 VDD.n6871 VDD.n2391 0.0341759
R40957 VDD.n6872 VDD.n6871 0.0341759
R40958 VDD.n6873 VDD.n6872 0.0341759
R40959 VDD.n6726 VDD.n2407 0.0341759
R40960 VDD.n6723 VDD.n2407 0.0341759
R40961 VDD.n6723 VDD.n6722 0.0341759
R40962 VDD.n6722 VDD.n6721 0.0341759
R40963 VDD.n6721 VDD.n6715 0.0341759
R40964 VDD.n6719 VDD.n6715 0.0341759
R40965 VDD.n6718 VDD.n6716 0.0341759
R40966 VDD.n6716 VDD.n2370 0.0341759
R40967 VDD.n7037 VDD.n7036 0.0341759
R40968 VDD.n7036 VDD.n2371 0.0341759
R40969 VDD.n7034 VDD.n2371 0.0341759
R40970 VDD.n7033 VDD.n2372 0.0341759
R40971 VDD.n7031 VDD.n2372 0.0341759
R40972 VDD.n7031 VDD.n7030 0.0341759
R40973 VDD.n7030 VDD.n7029 0.0341759
R40974 VDD.n7029 VDD.n2373 0.0341759
R40975 VDD.n7026 VDD.n2373 0.0341759
R40976 VDD.n5950 VDD.n5936 0.0337609
R40977 VDD.n6624 VDD.n6593 0.0337609
R40978 VDD.n5980 VDD.n5978 0.0337609
R40979 VDD.n5951 VDD.n5950 0.0337609
R40980 VDD.n6624 VDD.n6623 0.0337609
R40981 VDD.n5936 VDD.n5922 0.0331854
R40982 VDD.n5934 VDD.n5922 0.0331854
R40983 VDD.n5934 VDD.n5933 0.0331854
R40984 VDD.n5933 VDD.n5932 0.0331854
R40985 VDD.n5932 VDD.n5923 0.0331854
R40986 VDD.n5929 VDD.n5923 0.0331854
R40987 VDD.n5929 VDD.n5928 0.0331854
R40988 VDD.n5928 VDD.n5927 0.0331854
R40989 VDD.n5926 VDD.n5924 0.0331854
R40990 VDD.n5924 VDD.n5274 0.0331854
R40991 VDD.n6581 VDD.n6580 0.0331854
R40992 VDD.n6581 VDD.n5273 0.0331854
R40993 VDD.n6583 VDD.n5273 0.0331854
R40994 VDD.n6585 VDD.n6584 0.0331854
R40995 VDD.n6586 VDD.n6585 0.0331854
R40996 VDD.n6586 VDD.n5272 0.0331854
R40997 VDD.n6589 VDD.n5272 0.0331854
R40998 VDD.n6590 VDD.n6589 0.0331854
R40999 VDD.n6591 VDD.n6590 0.0331854
R41000 VDD.n6591 VDD.n5271 0.0331854
R41001 VDD.n6593 VDD.n5271 0.0331854
R41002 VDD.n5978 VDD.n5916 0.0331854
R41003 VDD.n5976 VDD.n5916 0.0331854
R41004 VDD.n5976 VDD.n5975 0.0331854
R41005 VDD.n5975 VDD.n5974 0.0331854
R41006 VDD.n5974 VDD.n5917 0.0331854
R41007 VDD.n5971 VDD.n5917 0.0331854
R41008 VDD.n5971 VDD.n5970 0.0331854
R41009 VDD.n5970 VDD.n5969 0.0331854
R41010 VDD.n5968 VDD.n5918 0.0331854
R41011 VDD.n5966 VDD.n5918 0.0331854
R41012 VDD.n5964 VDD.n5963 0.0331854
R41013 VDD.n5963 VDD.n5919 0.0331854
R41014 VDD.n5961 VDD.n5919 0.0331854
R41015 VDD.n5960 VDD.n5920 0.0331854
R41016 VDD.n5958 VDD.n5920 0.0331854
R41017 VDD.n5958 VDD.n5957 0.0331854
R41018 VDD.n5957 VDD.n5956 0.0331854
R41019 VDD.n5956 VDD.n5921 0.0331854
R41020 VDD.n5953 VDD.n5921 0.0331854
R41021 VDD.n5953 VDD.n5952 0.0331854
R41022 VDD.n5952 VDD.n5951 0.0331854
R41023 VDD.n6623 VDD.n6594 0.0331854
R41024 VDD.n6621 VDD.n6594 0.0331854
R41025 VDD.n6621 VDD.n6620 0.0331854
R41026 VDD.n6620 VDD.n6619 0.0331854
R41027 VDD.n6619 VDD.n6595 0.0331854
R41028 VDD.n6616 VDD.n6595 0.0331854
R41029 VDD.n6616 VDD.n6615 0.0331854
R41030 VDD.n6615 VDD.n6614 0.0331854
R41031 VDD.n6613 VDD.n6596 0.0331854
R41032 VDD.n6611 VDD.n6596 0.0331854
R41033 VDD.n6609 VDD.n6608 0.0331854
R41034 VDD.n6608 VDD.n6597 0.0331854
R41035 VDD.n6606 VDD.n6597 0.0331854
R41036 VDD.n6605 VDD.n6598 0.0331854
R41037 VDD.n6603 VDD.n6598 0.0331854
R41038 VDD.n6603 VDD.n6602 0.0331854
R41039 VDD.n6602 VDD.n6601 0.0331854
R41040 VDD.n7845 VDD.n2208 0.0331854
R41041 VDD.n7845 VDD.n7844 0.0331854
R41042 VDD.n7844 VDD.n7843 0.0331854
R41043 VDD.n1664 VDD.n1663 0.0331792
R41044 VDD.n1571 VDD.n1570 0.0331792
R41045 VDD.n1573 VDD.n1572 0.0331792
R41046 VDD.n1575 VDD.n1574 0.0331792
R41047 VDD.n1590 VDD.n1589 0.0331792
R41048 VDD.n1588 VDD.n1587 0.0331792
R41049 VDD.n1586 VDD.n1585 0.0331792
R41050 VDD.n1584 VDD.n1583 0.0331792
R41051 VDD.n1670 VDD.n1669 0.0331792
R41052 VDD.n1668 VDD.n1667 0.0331792
R41053 VDD.n1666 VDD.n1665 0.0331792
R41054 VDD.n7683 VDD.n7177 0.0328372
R41055 VDD.n6303 VDD.n6302 0.0325255
R41056 VDD.n6307 VDD.n6306 0.0325255
R41057 VDD.n5986 VDD.n5985 0.0325255
R41058 VDD.n6316 VDD.n6315 0.0325255
R41059 VDD.n6193 VDD.n6192 0.0325255
R41060 VDD.n6198 VDD.n6197 0.0325255
R41061 VDD.n6183 VDD.n6182 0.0325255
R41062 VDD.n6188 VDD.n6187 0.0325255
R41063 VDD.n6029 VDD.n6028 0.0325158
R41064 VDD.n6571 VDD.n6570 0.0325158
R41065 VDD.n6162 VDD.n6161 0.0325158
R41066 VDD.n6403 VDD.n6402 0.0325158
R41067 VDD.n8001 VDD.n8000 0.0325158
R41068 VDD.n2183 VDD.n2182 0.0325158
R41069 VDD.n6858 VDD.n6857 0.0325158
R41070 VDD.n6866 VDD.n6865 0.0325158
R41071 VDD.n6719 VDD.n6718 0.0325158
R41072 VDD.n7034 VDD.n7033 0.0325158
R41073 VDD.n1660 VDD.n1659 0.0324891
R41074 VDD.n1645 VDD.n1644 0.0324891
R41075 VDD.n7946 VDD.n7945 0.0320529
R41076 VDD.n7944 VDD.n7943 0.0320529
R41077 VDD.n7887 VDD.n7854 0.0320529
R41078 VDD.n7888 VDD.n2148 0.0320529
R41079 VDD.n8051 VDD.n8050 0.0320529
R41080 VDD.n8049 VDD.n8048 0.0320529
R41081 VDD.n2172 VDD.n2149 0.0320529
R41082 VDD.n1663 VDD.n753 0.0320159
R41083 VDD.n1662 VDD.n753 0.0320159
R41084 VDD.n1569 VDD.n1509 0.0320159
R41085 VDD.n1570 VDD.n1509 0.0320159
R41086 VDD.n1571 VDD.n1508 0.0320159
R41087 VDD.n1572 VDD.n1508 0.0320159
R41088 VDD.n1575 VDD.n1505 0.0320159
R41089 VDD.n1576 VDD.n1505 0.0320159
R41090 VDD.n1591 VDD.n1577 0.0320159
R41091 VDD.n1590 VDD.n1577 0.0320159
R41092 VDD.n1589 VDD.n1578 0.0320159
R41093 VDD.n1588 VDD.n1578 0.0320159
R41094 VDD.n1587 VDD.n1579 0.0320159
R41095 VDD.n1586 VDD.n1579 0.0320159
R41096 VDD.n1585 VDD.n1580 0.0320159
R41097 VDD.n1584 VDD.n1580 0.0320159
R41098 VDD.n1583 VDD.n1581 0.0320159
R41099 VDD.n1582 VDD.n1581 0.0320159
R41100 VDD.n1671 VDD.n748 0.0320159
R41101 VDD.n1670 VDD.n748 0.0320159
R41102 VDD.n1669 VDD.n749 0.0320159
R41103 VDD.n1668 VDD.n749 0.0320159
R41104 VDD.n1667 VDD.n750 0.0320159
R41105 VDD.n1666 VDD.n750 0.0320159
R41106 VDD.n6686 VDD.n6685 0.0319413
R41107 VDD.n6685 VDD.n6641 0.0319104
R41108 VDD.n7861 VDD.n2204 0.0319052
R41109 VDD.n7863 VDD.n7862 0.0319052
R41110 VDD.n7911 VDD.n7910 0.0319052
R41111 VDD.n7177 VDD.n7176 0.031686
R41112 VDD.n2296 VDD.n2295 0.031686
R41113 VDD.n2294 VDD.n2209 0.031686
R41114 VDD.n7838 VDD.n7837 0.031686
R41115 VDD.n7840 VDD.n7839 0.031686
R41116 VDD.n7842 VDD.n7841 0.031686
R41117 VDD.n2390 VDD.n2389 0.031686
R41118 VDD.n2388 VDD.n2387 0.031686
R41119 VDD.n2386 VDD.n2239 0.031686
R41120 VDD.n7831 VDD.n7830 0.031686
R41121 VDD.n7829 VDD.n7828 0.031686
R41122 VDD.n7826 VDD.n7825 0.031686
R41123 VDD.n7824 VDD.n7823 0.031686
R41124 VDD.n9134 VDD.n9127 0.0316781
R41125 VDD.n5927 VDD.n5926 0.0315742
R41126 VDD.n6584 VDD.n6583 0.0315742
R41127 VDD.n5969 VDD.n5968 0.0315742
R41128 VDD.n5961 VDD.n5960 0.0315742
R41129 VDD.n6614 VDD.n6613 0.0315742
R41130 VDD.n6606 VDD.n6605 0.0315742
R41131 VDD.n6711 VDD.n6710 0.0315707
R41132 VDD.n6702 VDD.n6701 0.0315707
R41133 VDD.n6697 VDD.n6696 0.0315707
R41134 VDD.n6688 VDD.n6687 0.0315707
R41135 VDD.n6640 VDD.n6639 0.0315707
R41136 VDD.n5437 VDD.n5436 0.0315707
R41137 VDD.n5442 VDD.n5441 0.0315707
R41138 VDD.n6627 VDD.n6626 0.0315707
R41139 VDD.n5368 VDD.n5367 0.0313793
R41140 VDD.n6373 VDD.n6372 0.0313793
R41141 VDD.n6368 VDD.n5377 0.0313793
R41142 VDD.n5943 VDD.n5941 0.0313793
R41143 VDD.n2366 VDD.n2360 0.0313793
R41144 VDD.n7136 VDD.n7135 0.0313793
R41145 VDD.n7131 VDD.n2320 0.0313793
R41146 VDD.n7043 VDD.n2347 0.0313793
R41147 VDD.n7309 VDD.n7302 0.0312734
R41148 VDD.n2208 VDD.n2206 0.0311937
R41149 VDD.n9124 VDD.n9123 0.0308128
R41150 VDD.n9139 VDD.n9138 0.0307932
R41151 VDD.n2970 VDD.n2969 0.0305815
R41152 VDD.n6575 VDD.n5283 0.0303814
R41153 VDD.n6398 VDD.n5302 0.0303814
R41154 VDD.n6861 VDD.n6860 0.0303814
R41155 VDD.n7038 VDD.n2370 0.0303814
R41156 VDD.n5288 VDD.n2410 0.0302628
R41157 VDD.n6413 VDD.n6412 0.0302628
R41158 VDD.n6876 VDD.n6875 0.0302628
R41159 VDD.n2396 VDD.n2375 0.0302628
R41160 VDD.n8162 VDD.n8161 0.0302193
R41161 VDD.n5576 VDD.n5575 0.0302193
R41162 VDD.n5658 VDD.n5657 0.0302193
R41163 VDD.n5841 VDD.n5840 0.0302193
R41164 VDD.n5774 VDD.n5773 0.0302193
R41165 VDD.n9005 VDD.n9004 0.0302193
R41166 VDD.n8834 VDD.n8833 0.0302193
R41167 VDD.n9121 VDD.n9120 0.0302193
R41168 VDD.n166 VDD.n165 0.0302193
R41169 VDD.n77 VDD.n76 0.0302193
R41170 VDD.n7998 VDD.n7997 0.0295514
R41171 VDD.n6579 VDD.n5274 0.0295026
R41172 VDD.n5966 VDD.n5965 0.0295026
R41173 VDD.n6611 VDD.n6610 0.0295026
R41174 VDD.n2056 VDD.n2055 0.0293162
R41175 VDD.n2057 VDD.n2056 0.0293162
R41176 VDD.n2057 VDD.n2026 0.0293162
R41177 VDD.n2059 VDD.n2026 0.0293162
R41178 VDD.n10771 VDD.n2060 0.0293162
R41179 VDD.n10769 VDD.n2060 0.0293162
R41180 VDD.n10769 VDD.n10768 0.0293162
R41181 VDD.n10768 VDD.n10767 0.0293162
R41182 VDD.n2045 VDD.n2044 0.0293162
R41183 VDD.n2045 VDD.n2037 0.0293162
R41184 VDD.n2047 VDD.n2037 0.0293162
R41185 VDD.n2050 VDD.n2049 0.0293162
R41186 VDD.n2051 VDD.n2050 0.0293162
R41187 VDD.n2051 VDD.n2036 0.0293162
R41188 VDD.n2053 VDD.n2036 0.0293162
R41189 VDD.n10808 VDD.n2005 0.0293162
R41190 VDD.n10806 VDD.n2005 0.0293162
R41191 VDD.n10806 VDD.n10805 0.0293162
R41192 VDD.n10805 VDD.n10804 0.0293162
R41193 VDD.n10802 VDD.n2006 0.0293162
R41194 VDD.n10800 VDD.n2006 0.0293162
R41195 VDD.n10800 VDD.n10799 0.0293162
R41196 VDD.n10799 VDD.n10798 0.0293162
R41197 VDD.n1983 VDD.n1982 0.0293162
R41198 VDD.n1984 VDD.n1983 0.0293162
R41199 VDD.n1984 VDD.n1953 0.0293162
R41200 VDD.n1986 VDD.n1953 0.0293162
R41201 VDD.n10811 VDD.n10810 0.0293162
R41202 VDD.n10812 VDD.n10811 0.0293162
R41203 VDD.n10812 VDD.n10809 0.0293162
R41204 VDD.n10814 VDD.n10809 0.0293162
R41205 VDD.n1963 VDD.n1962 0.0293162
R41206 VDD.n1963 VDD.n1955 0.0293162
R41207 VDD.n1965 VDD.n1955 0.0293162
R41208 VDD.n1968 VDD.n1967 0.0293162
R41209 VDD.n1969 VDD.n1968 0.0293162
R41210 VDD.n1969 VDD.n1954 0.0293162
R41211 VDD.n1971 VDD.n1954 0.0293162
R41212 VDD.n10866 VDD.n1932 0.0293162
R41213 VDD.n10864 VDD.n1932 0.0293162
R41214 VDD.n10864 VDD.n10863 0.0293162
R41215 VDD.n10863 VDD.n10862 0.0293162
R41216 VDD.n10860 VDD.n1933 0.0293162
R41217 VDD.n10858 VDD.n1933 0.0293162
R41218 VDD.n10858 VDD.n10857 0.0293162
R41219 VDD.n10857 VDD.n10856 0.0293162
R41220 VDD.n5509 VDD.n5504 0.0293162
R41221 VDD.n5507 VDD.n5504 0.0293162
R41222 VDD.n5507 VDD.n5506 0.0293162
R41223 VDD.n5506 VDD.n5505 0.0293162
R41224 VDD.n10869 VDD.n10868 0.0293162
R41225 VDD.n10870 VDD.n10869 0.0293162
R41226 VDD.n10870 VDD.n10867 0.0293162
R41227 VDD.n10872 VDD.n10867 0.0293162
R41228 VDD.n5519 VDD.n5518 0.0293162
R41229 VDD.n5519 VDD.n5511 0.0293162
R41230 VDD.n5521 VDD.n5511 0.0293162
R41231 VDD.n5524 VDD.n5523 0.0293162
R41232 VDD.n5525 VDD.n5524 0.0293162
R41233 VDD.n5525 VDD.n5510 0.0293162
R41234 VDD.n5527 VDD.n5510 0.0293162
R41235 VDD.n10921 VDD.n1905 0.0293162
R41236 VDD.n10919 VDD.n1905 0.0293162
R41237 VDD.n10919 VDD.n10918 0.0293162
R41238 VDD.n10918 VDD.n10917 0.0293162
R41239 VDD.n10915 VDD.n1906 0.0293162
R41240 VDD.n10913 VDD.n1906 0.0293162
R41241 VDD.n10913 VDD.n10912 0.0293162
R41242 VDD.n10912 VDD.n10911 0.0293162
R41243 VDD.n1891 VDD.n1890 0.0293162
R41244 VDD.n1892 VDD.n1891 0.0293162
R41245 VDD.n1892 VDD.n1861 0.0293162
R41246 VDD.n1894 VDD.n1861 0.0293162
R41247 VDD.n10924 VDD.n10923 0.0293162
R41248 VDD.n10925 VDD.n10924 0.0293162
R41249 VDD.n10925 VDD.n10922 0.0293162
R41250 VDD.n10927 VDD.n10922 0.0293162
R41251 VDD.n1871 VDD.n1870 0.0293162
R41252 VDD.n1871 VDD.n1863 0.0293162
R41253 VDD.n1873 VDD.n1863 0.0293162
R41254 VDD.n1876 VDD.n1875 0.0293162
R41255 VDD.n1877 VDD.n1876 0.0293162
R41256 VDD.n1877 VDD.n1862 0.0293162
R41257 VDD.n1879 VDD.n1862 0.0293162
R41258 VDD.n10976 VDD.n1840 0.0293162
R41259 VDD.n10974 VDD.n1840 0.0293162
R41260 VDD.n10974 VDD.n10973 0.0293162
R41261 VDD.n10973 VDD.n10972 0.0293162
R41262 VDD.n10970 VDD.n1841 0.0293162
R41263 VDD.n10968 VDD.n1841 0.0293162
R41264 VDD.n10968 VDD.n10967 0.0293162
R41265 VDD.n10967 VDD.n10966 0.0293162
R41266 VDD.n1826 VDD.n1825 0.0293162
R41267 VDD.n1827 VDD.n1826 0.0293162
R41268 VDD.n1827 VDD.n1796 0.0293162
R41269 VDD.n1829 VDD.n1796 0.0293162
R41270 VDD.n10979 VDD.n10978 0.0293162
R41271 VDD.n10980 VDD.n10979 0.0293162
R41272 VDD.n10980 VDD.n10977 0.0293162
R41273 VDD.n10982 VDD.n10977 0.0293162
R41274 VDD.n1815 VDD.n1814 0.0293162
R41275 VDD.n1815 VDD.n1807 0.0293162
R41276 VDD.n1817 VDD.n1807 0.0293162
R41277 VDD.n1820 VDD.n1819 0.0293162
R41278 VDD.n1821 VDD.n1820 0.0293162
R41279 VDD.n1821 VDD.n1806 0.0293162
R41280 VDD.n1823 VDD.n1806 0.0293162
R41281 VDD.n1775 VDD.n1774 0.0293162
R41282 VDD.n1776 VDD.n1775 0.0293162
R41283 VDD.n1776 VDD.n1773 0.0293162
R41284 VDD.n1778 VDD.n1773 0.0293162
R41285 VDD.n11025 VDD.n1779 0.0293162
R41286 VDD.n11023 VDD.n1779 0.0293162
R41287 VDD.n11023 VDD.n11022 0.0293162
R41288 VDD.n11022 VDD.n11021 0.0293162
R41289 VDD.n9071 VDD.n9070 0.0293162
R41290 VDD.n9071 VDD.n8474 0.0293162
R41291 VDD.n9073 VDD.n8474 0.0293162
R41292 VDD.n9155 VDD.n9074 0.0293162
R41293 VDD.n9153 VDD.n9074 0.0293162
R41294 VDD.n9153 VDD.n9152 0.0293162
R41295 VDD.n9152 VDD.n9151 0.0293162
R41296 VDD.n9023 VDD.n9022 0.0293162
R41297 VDD.n9024 VDD.n9023 0.0293162
R41298 VDD.n9024 VDD.n8494 0.0293162
R41299 VDD.n9026 VDD.n8494 0.0293162
R41300 VDD.n9031 VDD.n9027 0.0293162
R41301 VDD.n9029 VDD.n9027 0.0293162
R41302 VDD.n9029 VDD.n9028 0.0293162
R41303 VDD.n9028 VDD.n8476 0.0293162
R41304 VDD.n8906 VDD.n8902 0.0293162
R41305 VDD.n8904 VDD.n8902 0.0293162
R41306 VDD.n8904 VDD.n8903 0.0293162
R41307 VDD.n8903 VDD.n8499 0.0293162
R41308 VDD.n9017 VDD.n9016 0.0293162
R41309 VDD.n9018 VDD.n9017 0.0293162
R41310 VDD.n9018 VDD.n8498 0.0293162
R41311 VDD.n9020 VDD.n8498 0.0293162
R41312 VDD.n8898 VDD.n8897 0.0293162
R41313 VDD.n8898 VDD.n8512 0.0293162
R41314 VDD.n8900 VDD.n8512 0.0293162
R41315 VDD.n8934 VDD.n8901 0.0293162
R41316 VDD.n8932 VDD.n8901 0.0293162
R41317 VDD.n8932 VDD.n8931 0.0293162
R41318 VDD.n8931 VDD.n8930 0.0293162
R41319 VDD.n8775 VDD.n8771 0.0293162
R41320 VDD.n8773 VDD.n8771 0.0293162
R41321 VDD.n8773 VDD.n8772 0.0293162
R41322 VDD.n8772 VDD.n8518 0.0293162
R41323 VDD.n8886 VDD.n8885 0.0293162
R41324 VDD.n8887 VDD.n8886 0.0293162
R41325 VDD.n8887 VDD.n8517 0.0293162
R41326 VDD.n8889 VDD.n8517 0.0293162
R41327 VDD.n8766 VDD.n8765 0.0293162
R41328 VDD.n8767 VDD.n8766 0.0293162
R41329 VDD.n8767 VDD.n8531 0.0293162
R41330 VDD.n8769 VDD.n8531 0.0293162
R41331 VDD.n8803 VDD.n8770 0.0293162
R41332 VDD.n8801 VDD.n8770 0.0293162
R41333 VDD.n8801 VDD.n8800 0.0293162
R41334 VDD.n8800 VDD.n8799 0.0293162
R41335 VDD.n8755 VDD.n8754 0.0293162
R41336 VDD.n8755 VDD.n8581 0.0293162
R41337 VDD.n8757 VDD.n8581 0.0293162
R41338 VDD.n8760 VDD.n8759 0.0293162
R41339 VDD.n8761 VDD.n8760 0.0293162
R41340 VDD.n8761 VDD.n8580 0.0293162
R41341 VDD.n8763 VDD.n8580 0.0293162
R41342 VDD.n9149 VDD.n9084 0.0293162
R41343 VDD.n9147 VDD.n9084 0.0293162
R41344 VDD.n9147 VDD.n9146 0.0293162
R41345 VDD.n9146 VDD.n9145 0.0293162
R41346 VDD.n9143 VDD.n9085 0.0293162
R41347 VDD.n9141 VDD.n9085 0.0293162
R41348 VDD.n9141 VDD.n9140 0.0293162
R41349 VDD.n9140 VDD.n9139 0.0293162
R41350 VDD.n8737 VDD.n8736 0.0293162
R41351 VDD.n8738 VDD.n8737 0.0293162
R41352 VDD.n8738 VDD.n8593 0.0293162
R41353 VDD.n8740 VDD.n8593 0.0293162
R41354 VDD.n8743 VDD.n8742 0.0293162
R41355 VDD.n8744 VDD.n8743 0.0293162
R41356 VDD.n8744 VDD.n8592 0.0293162
R41357 VDD.n8746 VDD.n8592 0.0293162
R41358 VDD.n8716 VDD.n8715 0.0293162
R41359 VDD.n8717 VDD.n8716 0.0293162
R41360 VDD.n8717 VDD.n8595 0.0293162
R41361 VDD.n8719 VDD.n8595 0.0293162
R41362 VDD.n8722 VDD.n8721 0.0293162
R41363 VDD.n8723 VDD.n8722 0.0293162
R41364 VDD.n8723 VDD.n8594 0.0293162
R41365 VDD.n8725 VDD.n8594 0.0293162
R41366 VDD.n8705 VDD.n8704 0.0293162
R41367 VDD.n8705 VDD.n8606 0.0293162
R41368 VDD.n8707 VDD.n8606 0.0293162
R41369 VDD.n8710 VDD.n8709 0.0293162
R41370 VDD.n8711 VDD.n8710 0.0293162
R41371 VDD.n8711 VDD.n8605 0.0293162
R41372 VDD.n8713 VDD.n8605 0.0293162
R41373 VDD.n8678 VDD.n8677 0.0293162
R41374 VDD.n8679 VDD.n8678 0.0293162
R41375 VDD.n8679 VDD.n8609 0.0293162
R41376 VDD.n8681 VDD.n8609 0.0293162
R41377 VDD.n8684 VDD.n8683 0.0293162
R41378 VDD.n8685 VDD.n8684 0.0293162
R41379 VDD.n8685 VDD.n8608 0.0293162
R41380 VDD.n8687 VDD.n8608 0.0293162
R41381 VDD.n8666 VDD.n8665 0.0293162
R41382 VDD.n8667 VDD.n8666 0.0293162
R41383 VDD.n8667 VDD.n8620 0.0293162
R41384 VDD.n8669 VDD.n8620 0.0293162
R41385 VDD.n8672 VDD.n8671 0.0293162
R41386 VDD.n8673 VDD.n8672 0.0293162
R41387 VDD.n8673 VDD.n8619 0.0293162
R41388 VDD.n8675 VDD.n8619 0.0293162
R41389 VDD.n8646 VDD.n8645 0.0293162
R41390 VDD.n8646 VDD.n8622 0.0293162
R41391 VDD.n8648 VDD.n8622 0.0293162
R41392 VDD.n8651 VDD.n8650 0.0293162
R41393 VDD.n8652 VDD.n8651 0.0293162
R41394 VDD.n8652 VDD.n8621 0.0293162
R41395 VDD.n8654 VDD.n8621 0.0293162
R41396 VDD.n12620 VDD.n11 0.0293162
R41397 VDD.n12618 VDD.n11 0.0293162
R41398 VDD.n12618 VDD.n12617 0.0293162
R41399 VDD.n12617 VDD.n12616 0.0293162
R41400 VDD.n8634 VDD.n12 0.0293162
R41401 VDD.n8635 VDD.n8634 0.0293162
R41402 VDD.n8635 VDD.n8633 0.0293162
R41403 VDD.n8637 VDD.n8633 0.0293162
R41404 VDD.n7683 VDD.n7682 0.029
R41405 VDD.n2139 VDD.n2138 0.0289485
R41406 VDD.n1177 VDD.n1176 0.0287717
R41407 VDD.n1206 VDD.n1188 0.0287717
R41408 VDD.n1164 VDD.n1163 0.0287717
R41409 VDD.n1176 VDD.n1175 0.0287717
R41410 VDD.n1336 VDD.n1318 0.0287717
R41411 VDD.n1305 VDD.n1304 0.0287717
R41412 VDD.n1337 VDD.n1336 0.0287717
R41413 VDD.n1383 VDD.n1364 0.0287717
R41414 VDD.n1304 VDD.n1286 0.0287717
R41415 VDD.n1073 VDD.n1072 0.0287717
R41416 VDD.n1384 VDD.n1383 0.0287717
R41417 VDD.n1269 VDD.n1250 0.0287717
R41418 VDD.n1237 VDD.n1236 0.0287717
R41419 VDD.n1270 VDD.n1269 0.0287717
R41420 VDD.n1207 VDD.n1206 0.0287717
R41421 VDD.n1236 VDD.n1218 0.0287717
R41422 VDD.n1060 VDD.n1059 0.0287717
R41423 VDD.n1072 VDD.n1071 0.0287717
R41424 VDD.n905 VDD.n0 0.0287717
R41425 VDD.n1059 VDD.n916 0.0287717
R41426 VDD.n1751 VDD.n1750 0.0287717
R41427 VDD.n1163 VDD.n1162 0.0287717
R41428 VDD.n8132 VDD.n8131 0.0284144
R41429 VDD.n8165 VDD.n8164 0.0284144
R41430 VDD.n8111 VDD.n8110 0.0284144
R41431 VDD.n8131 VDD.n8121 0.0284144
R41432 VDD.n8099 VDD.n8098 0.0284144
R41433 VDD.n8110 VDD.n8109 0.0284144
R41434 VDD.n5594 VDD.n5584 0.0284144
R41435 VDD.n8098 VDD.n2104 0.0284144
R41436 VDD.n5615 VDD.n5605 0.0284144
R41437 VDD.n5595 VDD.n5594 0.0284144
R41438 VDD.n5636 VDD.n5626 0.0284144
R41439 VDD.n5616 VDD.n5615 0.0284144
R41440 VDD.n5900 VDD.n5666 0.0284144
R41441 VDD.n5637 VDD.n5636 0.0284144
R41442 VDD.n5866 VDD.n5865 0.0284144
R41443 VDD.n5900 VDD.n5876 0.0284144
R41444 VDD.n5854 VDD.n5853 0.0284144
R41445 VDD.n5865 VDD.n5864 0.0284144
R41446 VDD.n5811 VDD.n5810 0.0284144
R41447 VDD.n5853 VDD.n5843 0.0284144
R41448 VDD.n5799 VDD.n5798 0.0284144
R41449 VDD.n5810 VDD.n5809 0.0284144
R41450 VDD.n5778 VDD.n5777 0.0284144
R41451 VDD.n5798 VDD.n5788 0.0284144
R41452 VDD.n5744 VDD.n5743 0.0284144
R41453 VDD.n5777 VDD.n5776 0.0284144
R41454 VDD.n5723 VDD.n5722 0.0284144
R41455 VDD.n5743 VDD.n5733 0.0284144
R41456 VDD.n11037 VDD.n11036 0.0284144
R41457 VDD.n5722 VDD.n5721 0.0284144
R41458 VDD.n8998 VDD.n8975 0.0284144
R41459 VDD.n9043 VDD.n9042 0.0284144
R41460 VDD.n8947 VDD.n8946 0.0284144
R41461 VDD.n8999 VDD.n8998 0.0284144
R41462 VDD.n8871 VDD.n8848 0.0284144
R41463 VDD.n8946 VDD.n8945 0.0284144
R41464 VDD.n8838 VDD.n8837 0.0284144
R41465 VDD.n8872 VDD.n8871 0.0284144
R41466 VDD.n8560 VDD.n8547 0.0284144
R41467 VDD.n8837 VDD.n8836 0.0284144
R41468 VDD.n12449 VDD.n184 0.0284144
R41469 VDD.n8560 VDD.n8559 0.0284144
R41470 VDD.n170 VDD.n169 0.0284144
R41471 VDD.n12449 VDD.n190 0.0284144
R41472 VDD.n9167 VDD.n8470 0.0284144
R41473 VDD.n9043 VDD.n8488 0.0284144
R41474 VDD.n9167 VDD.n9166 0.0284144
R41475 VDD.n12487 VDD.n106 0.0284144
R41476 VDD.n169 VDD.n168 0.0284144
R41477 VDD.n12505 VDD.n12498 0.0284144
R41478 VDD.n12488 VDD.n12487 0.0284144
R41479 VDD.n90 VDD.n89 0.0284144
R41480 VDD.n12505 VDD.n12504 0.0284144
R41481 VDD.n12543 VDD.n26 0.0284144
R41482 VDD.n89 VDD.n79 0.0284144
R41483 VDD.n12599 VDD.n12554 0.0284144
R41484 VDD.n12544 VDD.n12543 0.0284144
R41485 VDD.n12587 VDD.n12586 0.0284144
R41486 VDD.n12599 VDD.n12598 0.0284144
R41487 VDD.n6713 VDD.n5220 0.0282968
R41488 VDD.n1177 VDD.n1117 0.0282826
R41489 VDD.n1178 VDD.n1117 0.0282826
R41490 VDD.n1179 VDD.n1116 0.0282826
R41491 VDD.n1181 VDD.n1116 0.0282826
R41492 VDD.n1182 VDD.n1181 0.0282826
R41493 VDD.n1184 VDD.n1115 0.0282826
R41494 VDD.n1186 VDD.n1115 0.0282826
R41495 VDD.n1187 VDD.n1114 0.0282826
R41496 VDD.n1188 VDD.n1114 0.0282826
R41497 VDD.n1164 VDD.n1138 0.0282826
R41498 VDD.n1165 VDD.n1138 0.0282826
R41499 VDD.n1166 VDD.n1137 0.0282826
R41500 VDD.n1168 VDD.n1137 0.0282826
R41501 VDD.n1169 VDD.n1168 0.0282826
R41502 VDD.n1171 VDD.n1136 0.0282826
R41503 VDD.n1173 VDD.n1136 0.0282826
R41504 VDD.n1174 VDD.n1135 0.0282826
R41505 VDD.n1175 VDD.n1135 0.0282826
R41506 VDD.n1318 VDD.n1312 0.0282826
R41507 VDD.n1317 VDD.n1312 0.0282826
R41508 VDD.n1316 VDD.n1313 0.0282826
R41509 VDD.n1314 VDD.n1313 0.0282826
R41510 VDD.n1314 VDD.n757 0.0282826
R41511 VDD.n1655 VDD.n756 0.0282826
R41512 VDD.n1657 VDD.n756 0.0282826
R41513 VDD.n1658 VDD.n755 0.0282826
R41514 VDD.n1659 VDD.n755 0.0282826
R41515 VDD.n1660 VDD.n754 0.0282826
R41516 VDD.n1305 VDD.n1280 0.0282826
R41517 VDD.n1306 VDD.n1280 0.0282826
R41518 VDD.n1308 VDD.n1307 0.0282826
R41519 VDD.n1309 VDD.n1308 0.0282826
R41520 VDD.n1309 VDD.n1278 0.0282826
R41521 VDD.n1341 VDD.n1279 0.0282826
R41522 VDD.n1339 VDD.n1279 0.0282826
R41523 VDD.n1338 VDD.n1311 0.0282826
R41524 VDD.n1337 VDD.n1311 0.0282826
R41525 VDD.n1364 VDD.n1080 0.0282826
R41526 VDD.n1363 VDD.n1080 0.0282826
R41527 VDD.n1362 VDD.n1081 0.0282826
R41528 VDD.n1360 VDD.n1081 0.0282826
R41529 VDD.n1360 VDD.n1359 0.0282826
R41530 VDD.n1282 VDD.n1082 0.0282826
R41531 VDD.n1284 VDD.n1282 0.0282826
R41532 VDD.n1285 VDD.n1281 0.0282826
R41533 VDD.n1286 VDD.n1281 0.0282826
R41534 VDD.n1073 VDD.n878 0.0282826
R41535 VDD.n1074 VDD.n878 0.0282826
R41536 VDD.n1076 VDD.n1075 0.0282826
R41537 VDD.n1077 VDD.n1076 0.0282826
R41538 VDD.n1077 VDD.n876 0.0282826
R41539 VDD.n1388 VDD.n877 0.0282826
R41540 VDD.n1386 VDD.n877 0.0282826
R41541 VDD.n1385 VDD.n1079 0.0282826
R41542 VDD.n1384 VDD.n1079 0.0282826
R41543 VDD.n1250 VDD.n1244 0.0282826
R41544 VDD.n1249 VDD.n1244 0.0282826
R41545 VDD.n1248 VDD.n1245 0.0282826
R41546 VDD.n1246 VDD.n1245 0.0282826
R41547 VDD.n1246 VDD.n765 0.0282826
R41548 VDD.n1649 VDD.n766 0.0282826
R41549 VDD.n1647 VDD.n766 0.0282826
R41550 VDD.n1646 VDD.n767 0.0282826
R41551 VDD.n1645 VDD.n767 0.0282826
R41552 VDD.n1644 VDD.n768 0.0282826
R41553 VDD.n1237 VDD.n1109 0.0282826
R41554 VDD.n1238 VDD.n1109 0.0282826
R41555 VDD.n1240 VDD.n1239 0.0282826
R41556 VDD.n1241 VDD.n1240 0.0282826
R41557 VDD.n1241 VDD.n1107 0.0282826
R41558 VDD.n1274 VDD.n1108 0.0282826
R41559 VDD.n1272 VDD.n1108 0.0282826
R41560 VDD.n1271 VDD.n1243 0.0282826
R41561 VDD.n1270 VDD.n1243 0.0282826
R41562 VDD.n1207 VDD.n1113 0.0282826
R41563 VDD.n1208 VDD.n1113 0.0282826
R41564 VDD.n1209 VDD.n1112 0.0282826
R41565 VDD.n1211 VDD.n1112 0.0282826
R41566 VDD.n1212 VDD.n1211 0.0282826
R41567 VDD.n1214 VDD.n1111 0.0282826
R41568 VDD.n1216 VDD.n1111 0.0282826
R41569 VDD.n1217 VDD.n1110 0.0282826
R41570 VDD.n1218 VDD.n1110 0.0282826
R41571 VDD.n1060 VDD.n900 0.0282826
R41572 VDD.n1061 VDD.n900 0.0282826
R41573 VDD.n1062 VDD.n899 0.0282826
R41574 VDD.n1064 VDD.n899 0.0282826
R41575 VDD.n1065 VDD.n1064 0.0282826
R41576 VDD.n1067 VDD.n898 0.0282826
R41577 VDD.n1069 VDD.n898 0.0282826
R41578 VDD.n1070 VDD.n897 0.0282826
R41579 VDD.n1071 VDD.n897 0.0282826
R41580 VDD.n905 VDD.n904 0.0282826
R41581 VDD.n906 VDD.n904 0.0282826
R41582 VDD.n907 VDD.n903 0.0282826
R41583 VDD.n909 VDD.n903 0.0282826
R41584 VDD.n910 VDD.n909 0.0282826
R41585 VDD.n912 VDD.n902 0.0282826
R41586 VDD.n914 VDD.n902 0.0282826
R41587 VDD.n915 VDD.n901 0.0282826
R41588 VDD.n916 VDD.n901 0.0282826
R41589 VDD.n1750 VDD.n683 0.0282826
R41590 VDD.n1749 VDD.n683 0.0282826
R41591 VDD.n1748 VDD.n684 0.0282826
R41592 VDD.n1746 VDD.n684 0.0282826
R41593 VDD.n1746 VDD.n1745 0.0282826
R41594 VDD.n1158 VDD.n685 0.0282826
R41595 VDD.n1160 VDD.n1158 0.0282826
R41596 VDD.n1161 VDD.n1157 0.0282826
R41597 VDD.n1162 VDD.n1157 0.0282826
R41598 VDD.n11873 VDD.n11872 0.027875
R41599 VDD.n8086 VDD.n2120 0.027874
R41600 VDD.n72 VDD.n56 0.0271036
R41601 VDD.n161 VDD.n145 0.0271036
R41602 VDD.n5771 VDD.n5755 0.0271036
R41603 VDD.n5838 VDD.n5822 0.0271036
R41604 VDD.n5655 VDD.n5639 0.0271036
R41605 VDD.n5573 VDD.n5557 0.0271036
R41606 VDD.n8159 VDD.n8143 0.0271036
R41607 VDD.n9116 VDD.n9100 0.0271036
R41608 VDD.n8829 VDD.n8813 0.0271036
R41609 VDD.n9000 VDD.n8969 0.0271036
R41610 VDD.n12572 VDD.n12570 0.0270708
R41611 VDD.n1179 VDD.n1178 0.026913
R41612 VDD.n1184 VDD.n1183 0.026913
R41613 VDD.n1187 VDD.n1186 0.026913
R41614 VDD.n1166 VDD.n1165 0.026913
R41615 VDD.n1171 VDD.n1170 0.026913
R41616 VDD.n1174 VDD.n1173 0.026913
R41617 VDD.n1317 VDD.n1316 0.026913
R41618 VDD.n1655 VDD.n1654 0.026913
R41619 VDD.n1658 VDD.n1657 0.026913
R41620 VDD.n1307 VDD.n1306 0.026913
R41621 VDD.n1342 VDD.n1341 0.026913
R41622 VDD.n1339 VDD.n1338 0.026913
R41623 VDD.n1363 VDD.n1362 0.026913
R41624 VDD.n1358 VDD.n1082 0.026913
R41625 VDD.n1285 VDD.n1284 0.026913
R41626 VDD.n1075 VDD.n1074 0.026913
R41627 VDD.n1389 VDD.n1388 0.026913
R41628 VDD.n1386 VDD.n1385 0.026913
R41629 VDD.n1249 VDD.n1248 0.026913
R41630 VDD.n1650 VDD.n1649 0.026913
R41631 VDD.n1647 VDD.n1646 0.026913
R41632 VDD.n1239 VDD.n1238 0.026913
R41633 VDD.n1275 VDD.n1274 0.026913
R41634 VDD.n1272 VDD.n1271 0.026913
R41635 VDD.n1209 VDD.n1208 0.026913
R41636 VDD.n1214 VDD.n1213 0.026913
R41637 VDD.n1217 VDD.n1216 0.026913
R41638 VDD.n1062 VDD.n1061 0.026913
R41639 VDD.n1067 VDD.n1066 0.026913
R41640 VDD.n1070 VDD.n1069 0.026913
R41641 VDD.n907 VDD.n906 0.026913
R41642 VDD.n912 VDD.n911 0.026913
R41643 VDD.n915 VDD.n914 0.026913
R41644 VDD.n1749 VDD.n1748 0.026913
R41645 VDD.n1744 VDD.n685 0.026913
R41646 VDD.n1161 VDD.n1160 0.026913
R41647 VDD.n1531 VDD.n1530 0.0266202
R41648 VDD.n1544 VDD.n1543 0.0266202
R41649 VDD.n8079 VDD.n2122 0.0261926
R41650 VDD.n9436 VDD.n195 0.026
R41651 VDD.n8075 VDD.n2125 0.0259774
R41652 VDD.n5201 VDD.n5200 0.025625
R41653 VDD.n6302 VDD.n6301 0.0249708
R41654 VDD.n6304 VDD.n6303 0.0249708
R41655 VDD.n6308 VDD.n6307 0.0249708
R41656 VDD.n6306 VDD.n6305 0.0249708
R41657 VDD.n5985 VDD.n5984 0.0249708
R41658 VDD.n5987 VDD.n5986 0.0249708
R41659 VDD.n6315 VDD.n6314 0.0249708
R41660 VDD.n6317 VDD.n6316 0.0249708
R41661 VDD.n6192 VDD.n6191 0.0249708
R41662 VDD.n6194 VDD.n6193 0.0249708
R41663 VDD.n6197 VDD.n6196 0.0249708
R41664 VDD.n6199 VDD.n6198 0.0249708
R41665 VDD.n6182 VDD.n6181 0.0249708
R41666 VDD.n6184 VDD.n6183 0.0249708
R41667 VDD.n6187 VDD.n6186 0.0249708
R41668 VDD.n6189 VDD.n6188 0.0249708
R41669 VDD.n8080 VDD.n2119 0.0242213
R41670 VDD.n8164 VDD.n2089 0.0240829
R41671 VDD.n5556 VDD.n2104 0.0240829
R41672 VDD.n5638 VDD.n5637 0.0240829
R41673 VDD.n5843 VDD.n5680 0.0240829
R41674 VDD.n5776 VDD.n5704 0.0240829
R41675 VDD.n9001 VDD.n8999 0.0240829
R41676 VDD.n8836 VDD.n8525 0.0240829
R41677 VDD.n9123 VDD.n9090 0.0240829
R41678 VDD.n168 VDD.n135 0.0240829
R41679 VDD.n79 VDD.n46 0.0240829
R41680 VDD.n2055 VDD.n2054 0.02404
R41681 VDD.n10767 VDD.n10766 0.02404
R41682 VDD.n2054 VDD.n2053 0.02404
R41683 VDD.n10815 VDD.n10808 0.02404
R41684 VDD.n10798 VDD.n10797 0.02404
R41685 VDD.n1982 VDD.n1981 0.02404
R41686 VDD.n10815 VDD.n10814 0.02404
R41687 VDD.n1981 VDD.n1971 0.02404
R41688 VDD.n10873 VDD.n10866 0.02404
R41689 VDD.n10856 VDD.n10855 0.02404
R41690 VDD.n5528 VDD.n5509 0.02404
R41691 VDD.n10873 VDD.n10872 0.02404
R41692 VDD.n5528 VDD.n5527 0.02404
R41693 VDD.n10928 VDD.n10921 0.02404
R41694 VDD.n10911 VDD.n10910 0.02404
R41695 VDD.n1890 VDD.n1889 0.02404
R41696 VDD.n10928 VDD.n10927 0.02404
R41697 VDD.n1889 VDD.n1879 0.02404
R41698 VDD.n10983 VDD.n10976 0.02404
R41699 VDD.n10966 VDD.n10965 0.02404
R41700 VDD.n1825 VDD.n1824 0.02404
R41701 VDD.n10983 VDD.n10982 0.02404
R41702 VDD.n1824 VDD.n1823 0.02404
R41703 VDD.n1774 VDD.n644 0.02404
R41704 VDD.n11021 VDD.n11020 0.02404
R41705 VDD.n9151 VDD.n9150 0.02404
R41706 VDD.n9022 VDD.n9021 0.02404
R41707 VDD.n9063 VDD.n8476 0.02404
R41708 VDD.n8929 VDD.n8906 0.02404
R41709 VDD.n9021 VDD.n9020 0.02404
R41710 VDD.n8930 VDD.n8929 0.02404
R41711 VDD.n8798 VDD.n8775 0.02404
R41712 VDD.n8890 VDD.n8889 0.02404
R41713 VDD.n8765 VDD.n8764 0.02404
R41714 VDD.n8799 VDD.n8798 0.02404
R41715 VDD.n8764 VDD.n8763 0.02404
R41716 VDD.n9150 VDD.n9149 0.02404
R41717 VDD.n8736 VDD.n8735 0.02404
R41718 VDD.n8747 VDD.n8746 0.02404
R41719 VDD.n8715 VDD.n8714 0.02404
R41720 VDD.n8735 VDD.n8725 0.02404
R41721 VDD.n8714 VDD.n8713 0.02404
R41722 VDD.n8677 VDD.n8676 0.02404
R41723 VDD.n8697 VDD.n8687 0.02404
R41724 VDD.n8665 VDD.n8664 0.02404
R41725 VDD.n8676 VDD.n8675 0.02404
R41726 VDD.n8664 VDD.n8654 0.02404
R41727 VDD.n12621 VDD.n12620 0.02404
R41728 VDD.n8638 VDD.n8637 0.02404
R41729 VDD.n2142 VDD.n2141 0.0234742
R41730 VDD.n2140 VDD.n2139 0.0234742
R41731 VDD.n6713 VDD.n6712 0.0232316
R41732 VDD.n2044 VDD.n2043 0.0232283
R41733 VDD.n1962 VDD.n1961 0.0232283
R41734 VDD.n5518 VDD.n5517 0.0232283
R41735 VDD.n1870 VDD.n1869 0.0232283
R41736 VDD.n1814 VDD.n1813 0.0232283
R41737 VDD.n9070 VDD.n9069 0.0232283
R41738 VDD.n8897 VDD.n8896 0.0232283
R41739 VDD.n8754 VDD.n8753 0.0232283
R41740 VDD.n8704 VDD.n8703 0.0232283
R41741 VDD.n8645 VDD.n8644 0.0232283
R41742 VDD.n6379 VDD.n5374 0.0228966
R41743 VDD.n6362 VDD.n6361 0.0228966
R41744 VDD.n7142 VDD.n2311 0.0228966
R41745 VDD.n7125 VDD.n7124 0.0228966
R41746 VDD.n6379 VDD.n6378 0.0228448
R41747 VDD.n6361 VDD.n5473 0.0228448
R41748 VDD.n7142 VDD.n7141 0.0228448
R41749 VDD.n7124 VDD.n2323 0.0228448
R41750 VDD.n1204 VDD.n1203 0.0225862
R41751 VDD.n1133 VDD.n1132 0.0225862
R41752 VDD.n1334 VDD.n1333 0.0225862
R41753 VDD.n1381 VDD.n1380 0.0225862
R41754 VDD.n1267 VDD.n1266 0.0225862
R41755 VDD.n1234 VDD.n1233 0.0225862
R41756 VDD.n1302 VDD.n1301 0.0225862
R41757 VDD.n895 VDD.n894 0.0225862
R41758 VDD.n1057 VDD.n1056 0.0225862
R41759 VDD.n1155 VDD.n1154 0.0225862
R41760 VDD.n2132 VDD.n2131 0.0224615
R41761 VDD.n12570 VDD.n12569 0.0222742
R41762 VDD.n1642 VDD.n769 0.0221383
R41763 VDD.n6706 VDD.n6705 0.0217183
R41764 VDD.n6692 VDD.n6691 0.0217183
R41765 VDD.n6635 VDD.n5267 0.0217183
R41766 VDD.n6631 VDD.n6630 0.0217183
R41767 VDD.n2120 VDD.n2119 0.021485
R41768 VDD.n4591 VDD.n4590 0.0214211
R41769 VDD.n4590 VDD.n2409 0.0214211
R41770 VDD.n2425 VDD.n2424 0.0207876
R41771 VDD.n5217 VDD.n4593 0.0207876
R41772 VDD.n5204 VDD.n5203 0.0207876
R41773 VDD.n4592 VDD.n2424 0.0207876
R41774 VDD.n5205 VDD.n4594 0.0207876
R41775 VDD.n4599 VDD.n4597 0.0207876
R41776 VDD.n12444 VDD.n194 0.0207876
R41777 VDD.n9200 VDD.n9199 0.0207876
R41778 VDD.n9187 VDD.n8458 0.0207876
R41779 VDD.n12447 VDD.n12446 0.0207876
R41780 VDD.n5366 VDD.n5365 0.0206724
R41781 VDD.n5371 VDD.n5370 0.0206724
R41782 VDD.n6375 VDD.n6374 0.0206724
R41783 VDD.n6217 VDD.n6216 0.0206724
R41784 VDD.n6264 VDD.n6263 0.0206724
R41785 VDD.n6366 VDD.n6365 0.0206724
R41786 VDD.n5940 VDD.n5939 0.0206724
R41787 VDD.n5946 VDD.n5945 0.0206724
R41788 VDD.n2359 VDD.n2358 0.0206724
R41789 VDD.n2364 VDD.n2363 0.0206724
R41790 VDD.n7138 VDD.n7137 0.0206724
R41791 VDD.n2315 VDD.n2314 0.0206724
R41792 VDD.n2398 VDD.n2397 0.0206724
R41793 VDD.n7129 VDD.n7128 0.0206724
R41794 VDD.n2346 VDD.n2345 0.0206724
R41795 VDD.n7046 VDD.n7045 0.0206724
R41796 VDD.n1708 VDD.n728 0.0206207
R41797 VDD.n1610 VDD.n802 0.0206207
R41798 VDD.n1442 VDD.n839 0.0206207
R41799 VDD.n1480 VDD.n1476 0.0206207
R41800 VDD.n1708 VDD.n1707 0.0206207
R41801 VDD.n1732 VDD.n699 0.0206207
R41802 VDD.n1732 VDD.n1731 0.0206207
R41803 VDD.n6563 VDD.n6562 0.0204161
R41804 VDD.n6410 VDD.n5297 0.0204161
R41805 VDD.n6873 VDD.n2384 0.0204161
R41806 VDD.n7026 VDD.n7025 0.0204161
R41807 VDD.n1533 VDD.n1532 0.0203361
R41808 VDD.n1546 VDD.n1545 0.0203361
R41809 VDD.n75 VDD.n72 0.0199738
R41810 VDD.n164 VDD.n161 0.0199738
R41811 VDD.n5772 VDD.n5771 0.0199738
R41812 VDD.n5839 VDD.n5838 0.0199738
R41813 VDD.n5656 VDD.n5655 0.0199738
R41814 VDD.n5574 VDD.n5573 0.0199738
R41815 VDD.n8160 VDD.n8159 0.0199738
R41816 VDD.n9119 VDD.n9116 0.0199738
R41817 VDD.n8832 VDD.n8829 0.0199738
R41818 VDD.n9003 VDD.n8969 0.0199738
R41819 VDD.n6037 VDD.n6022 0.019782
R41820 VDD.n6157 VDD.n6018 0.019782
R41821 VDD.n6849 VDD.n2404 0.019782
R41822 VDD.n6727 VDD.n2406 0.019782
R41823 VDD.n6009 VDD.n6007 0.0196477
R41824 VDD.n6331 VDD.n6330 0.0196477
R41825 VDD.n7173 VDD.n7172 0.0196477
R41826 VDD.n7096 VDD.n7095 0.0196477
R41827 VDD.n9138 VDD.n9137 0.0193079
R41828 VDD.n9136 VDD.n9135 0.0193079
R41829 VDD.n9127 VDD.n9126 0.0193079
R41830 VDD.n9125 VDD.n9124 0.0193079
R41831 VDD.n12566 VDD.n12565 0.0193079
R41832 VDD.n12569 VDD.n12567 0.0193079
R41833 VDD.n12573 VDD.n12572 0.0193079
R41834 VDD.n12576 VDD.n12574 0.0193079
R41835 VDD.n8128 VDD.n8127 0.0192265
R41836 VDD.n2032 VDD.n2031 0.0192265
R41837 VDD.n2099 VDD.n2098 0.0192265
R41838 VDD.n10793 VDD.n10792 0.0192265
R41839 VDD.n5591 VDD.n5590 0.0192265
R41840 VDD.n1977 VDD.n1976 0.0192265
R41841 VDD.n5612 VDD.n5611 0.0192265
R41842 VDD.n10851 VDD.n10850 0.0192265
R41843 VDD.n5897 VDD.n5896 0.0192265
R41844 VDD.n5499 VDD.n5498 0.0192265
R41845 VDD.n5675 VDD.n5674 0.0192265
R41846 VDD.n10906 VDD.n10905 0.0192265
R41847 VDD.n5688 VDD.n5687 0.0192265
R41848 VDD.n1885 VDD.n1884 0.0192265
R41849 VDD.n5795 VDD.n5794 0.0192265
R41850 VDD.n10961 VDD.n10960 0.0192265
R41851 VDD.n5740 VDD.n5739 0.0192265
R41852 VDD.n1802 VDD.n1801 0.0192265
R41853 VDD.n5714 VDD.n5713 0.0192265
R41854 VDD.n11016 VDD.n11015 0.0192265
R41855 VDD.n9060 VDD.n9059 0.0192265
R41856 VDD.n9048 VDD.n9046 0.0192265
R41857 VDD.n8926 VDD.n8925 0.0192265
R41858 VDD.n8914 VDD.n8912 0.0192265
R41859 VDD.n8852 VDD.n8849 0.0192265
R41860 VDD.n8867 VDD.n8866 0.0192265
R41861 VDD.n8577 VDD.n8576 0.0192265
R41862 VDD.n8565 VDD.n8563 0.0192265
R41863 VDD.n9081 VDD.n9080 0.0192265
R41864 VDD.n9172 VDD.n9170 0.0192265
R41865 VDD.n8589 VDD.n8588 0.0192265
R41866 VDD.n12454 VDD.n12452 0.0192265
R41867 VDD.n8602 VDD.n8601 0.0192265
R41868 VDD.n12483 VDD.n12482 0.0192265
R41869 VDD.n8694 VDD.n8693 0.0192265
R41870 VDD.n12510 VDD.n12508 0.0192265
R41871 VDD.n8661 VDD.n8660 0.0192265
R41872 VDD.n12539 VDD.n12538 0.0192265
R41873 VDD.n8630 VDD.n8629 0.0192265
R41874 VDD.n12604 VDD.n12602 0.0192265
R41875 VDD.n8086 VDD.n8085 0.019179
R41876 VDD.n2116 VDD.n2115 0.0190522
R41877 VDD.n10823 VDD.n10821 0.0190522
R41878 VDD.n5633 VDD.n5632 0.0190522
R41879 VDD.n10878 VDD.n10876 0.0190522
R41880 VDD.n5850 VDD.n5849 0.0190522
R41881 VDD.n10933 VDD.n10931 0.0190522
R41882 VDD.n5701 VDD.n5700 0.0190522
R41883 VDD.n10988 VDD.n10986 0.0190522
R41884 VDD.n8979 VDD.n8976 0.0190522
R41885 VDD.n8994 VDD.n8993 0.0190522
R41886 VDD.n8795 VDD.n8794 0.0190522
R41887 VDD.n8783 VDD.n8781 0.0190522
R41888 VDD.n8732 VDD.n8731 0.0190522
R41889 VDD.n131 VDD.n130 0.0190522
R41890 VDD.n8616 VDD.n8615 0.0190522
R41891 VDD.n85 VDD.n84 0.0190522
R41892 VDD.n6707 VDD.n6706 0.0189386
R41893 VDD.n6693 VDD.n6692 0.0189386
R41894 VDD.n6636 VDD.n6635 0.0189386
R41895 VDD.n6631 VDD.n5269 0.0189386
R41896 VDD.n12562 VDD.n12559 0.0186448
R41897 VDD.n12578 VDD.n12559 0.0186448
R41898 VDD.n643 VDD.n637 0.0186448
R41899 VDD.n639 VDD.n637 0.0186448
R41900 VDD.n11128 VDD.n636 0.0186448
R41901 VDD.n675 VDD.n672 0.0186448
R41902 VDD.n675 VDD.n671 0.0186448
R41903 VDD.n674 VDD.n670 0.0186448
R41904 VDD.n6322 VDD.n6321 0.0186448
R41905 VDD.n5982 VDD.n5913 0.0186448
R41906 VDD.n6324 VDD.n5915 0.0186448
R41907 VDD.n6321 VDD.n5983 0.0186448
R41908 VDD.n5983 VDD.n5982 0.0186448
R41909 VDD.n5981 VDD.n5915 0.0186448
R41910 VDD.n6176 VDD.n6015 0.0186448
R41911 VDD.n6178 VDD.n6017 0.0186448
R41912 VDD.n6172 VDD.n6012 0.0186448
R41913 VDD.n6176 VDD.n6012 0.0186448
R41914 VDD.n6017 VDD.n6011 0.0186448
R41915 VDD.n5532 VDD.n5531 0.0186448
R41916 VDD.n5531 VDD.n5530 0.0186448
R41917 VDD.n5536 VDD.n5535 0.0186448
R41918 VDD.n5882 VDD.n5881 0.0186448
R41919 VDD.n5887 VDD.n5881 0.0186448
R41920 VDD.n5885 VDD.n5884 0.0186448
R41921 VDD.n5906 VDD.n5904 0.0186448
R41922 VDD.n5903 VDD.n5540 0.0186448
R41923 VDD.n5909 VDD.n5908 0.0186448
R41924 VDD.n10816 VDD.n1997 0.0186448
R41925 VDD.n2003 VDD.n1997 0.0186448
R41926 VDD.n10818 VDD.n1996 0.0186448
R41927 VDD.n8093 VDD.n2110 0.0186448
R41928 VDD.n2110 VDD.n2107 0.0186448
R41929 VDD.n2118 VDD.n2117 0.0186448
R41930 VDD.n10816 VDD.n2001 0.0186448
R41931 VDD.n10819 VDD.n10818 0.0186448
R41932 VDD.n8094 VDD.n8093 0.0186448
R41933 VDD.n8091 VDD.n2107 0.0186448
R41934 VDD.n2117 VDD.n2109 0.0186448
R41935 VDD.n2003 VDD.n2002 0.0186448
R41936 VDD.n5533 VDD.n5532 0.0186448
R41937 VDD.n5883 VDD.n5882 0.0186448
R41938 VDD.n5904 VDD.n5903 0.0186448
R41939 VDD.n5530 VDD.n5489 0.0186448
R41940 VDD.n5910 VDD.n5909 0.0186448
R41941 VDD.n5884 VDD.n5880 0.0186448
R41942 VDD.n5888 VDD.n5887 0.0186448
R41943 VDD.n5537 VDD.n5536 0.0186448
R41944 VDD.n1764 VDD.n671 0.0186448
R41945 VDD.n11045 VDD.n670 0.0186448
R41946 VDD.n11047 VDD.n672 0.0186448
R41947 VDD.n11129 VDD.n11128 0.0186448
R41948 VDD.n639 VDD.n634 0.0186448
R41949 VDD.n643 VDD.n635 0.0186448
R41950 VDD.n12578 VDD.n12561 0.0186448
R41951 VDD.n12580 VDD.n12560 0.0186448
R41952 VDD.n12584 VDD.n12562 0.0186448
R41953 VDD.n12628 VDD.n12627 0.0186448
R41954 VDD.n12622 VDD.n8 0.0186448
R41955 VDD.n12631 VDD.n10 0.0186448
R41956 VDD.n12629 VDD.n10 0.0186448
R41957 VDD.n12627 VDD.n12623 0.0186448
R41958 VDD.n12623 VDD.n12622 0.0186448
R41959 VDD.n12638 VDD.n12637 0.0186448
R41960 VDD.n4 VDD.n3 0.0186448
R41961 VDD.n1001 VDD.n955 0.0186448
R41962 VDD.n999 VDD.n953 0.0186448
R41963 VDD.n1754 VDD.n1753 0.0186448
R41964 VDD.n1758 VDD.n1757 0.0186448
R41965 VDD.n1753 VDD.n677 0.0186448
R41966 VDD.n1759 VDD.n1758 0.0186448
R41967 VDD.n999 VDD.n954 0.0186448
R41968 VDD.n957 VDD.n955 0.0186448
R41969 VDD.n5 VDD.n4 0.0186448
R41970 VDD.n12637 VDD.n12636 0.0186448
R41971 VDD.n10772 VDD.n2059 0.0185609
R41972 VDD.n2048 VDD.n2047 0.0185609
R41973 VDD.n10804 VDD.n10803 0.0185609
R41974 VDD.n1987 VDD.n1986 0.0185609
R41975 VDD.n1966 VDD.n1965 0.0185609
R41976 VDD.n10862 VDD.n10861 0.0185609
R41977 VDD.n5505 VDD.n1922 0.0185609
R41978 VDD.n5522 VDD.n5521 0.0185609
R41979 VDD.n10917 VDD.n10916 0.0185609
R41980 VDD.n1895 VDD.n1894 0.0185609
R41981 VDD.n1874 VDD.n1873 0.0185609
R41982 VDD.n10972 VDD.n10971 0.0185609
R41983 VDD.n1830 VDD.n1829 0.0185609
R41984 VDD.n1818 VDD.n1817 0.0185609
R41985 VDD.n11026 VDD.n1778 0.0185609
R41986 VDD.n9156 VDD.n9073 0.0185609
R41987 VDD.n9032 VDD.n9026 0.0185609
R41988 VDD.n9015 VDD.n8499 0.0185609
R41989 VDD.n8935 VDD.n8900 0.0185609
R41990 VDD.n8884 VDD.n8518 0.0185609
R41991 VDD.n8804 VDD.n8769 0.0185609
R41992 VDD.n8758 VDD.n8757 0.0185609
R41993 VDD.n9145 VDD.n9144 0.0185609
R41994 VDD.n8741 VDD.n8740 0.0185609
R41995 VDD.n8720 VDD.n8719 0.0185609
R41996 VDD.n8708 VDD.n8707 0.0185609
R41997 VDD.n8682 VDD.n8681 0.0185609
R41998 VDD.n8670 VDD.n8669 0.0185609
R41999 VDD.n8649 VDD.n8648 0.0185609
R42000 VDD.n12616 VDD.n12615 0.0185609
R42001 VDD.n8065 VDD.n8064 0.0185
R42002 VDD.n8125 VDD.n8124 0.0183497
R42003 VDD.n2028 VDD.n2027 0.0183497
R42004 VDD.n2096 VDD.n2095 0.0183497
R42005 VDD.n10789 VDD.n10788 0.0183497
R42006 VDD.n5588 VDD.n5587 0.0183497
R42007 VDD.n1973 VDD.n1972 0.0183497
R42008 VDD.n5609 VDD.n5608 0.0183497
R42009 VDD.n10847 VDD.n10846 0.0183497
R42010 VDD.n5894 VDD.n5893 0.0183497
R42011 VDD.n5495 VDD.n5494 0.0183497
R42012 VDD.n5672 VDD.n5671 0.0183497
R42013 VDD.n10902 VDD.n10901 0.0183497
R42014 VDD.n5685 VDD.n5684 0.0183497
R42015 VDD.n1881 VDD.n1880 0.0183497
R42016 VDD.n5792 VDD.n5791 0.0183497
R42017 VDD.n10957 VDD.n10956 0.0183497
R42018 VDD.n5737 VDD.n5736 0.0183497
R42019 VDD.n1798 VDD.n1797 0.0183497
R42020 VDD.n5711 VDD.n5710 0.0183497
R42021 VDD.n11012 VDD.n11011 0.0183497
R42022 VDD.n9057 VDD.n9056 0.0183497
R42023 VDD.n9050 VDD.n9049 0.0183497
R42024 VDD.n8923 VDD.n8922 0.0183497
R42025 VDD.n8916 VDD.n8915 0.0183497
R42026 VDD.n8854 VDD.n8853 0.0183497
R42027 VDD.n8863 VDD.n8862 0.0183497
R42028 VDD.n8574 VDD.n8573 0.0183497
R42029 VDD.n8567 VDD.n8566 0.0183497
R42030 VDD.n9078 VDD.n9077 0.0183497
R42031 VDD.n9174 VDD.n9173 0.0183497
R42032 VDD.n8586 VDD.n8585 0.0183497
R42033 VDD.n12456 VDD.n12455 0.0183497
R42034 VDD.n8599 VDD.n8598 0.0183497
R42035 VDD.n12479 VDD.n12478 0.0183497
R42036 VDD.n8691 VDD.n8690 0.0183497
R42037 VDD.n12512 VDD.n12511 0.0183497
R42038 VDD.n8658 VDD.n8657 0.0183497
R42039 VDD.n12535 VDD.n12534 0.0183497
R42040 VDD.n8627 VDD.n8626 0.0183497
R42041 VDD.n12606 VDD.n12605 0.0183497
R42042 VDD.n2113 VDD.n2112 0.0181836
R42043 VDD.n10825 VDD.n10824 0.0181836
R42044 VDD.n5630 VDD.n5629 0.0181836
R42045 VDD.n10880 VDD.n10879 0.0181836
R42046 VDD.n5847 VDD.n5846 0.0181836
R42047 VDD.n10935 VDD.n10934 0.0181836
R42048 VDD.n5698 VDD.n5697 0.0181836
R42049 VDD.n10990 VDD.n10989 0.0181836
R42050 VDD.n8981 VDD.n8980 0.0181836
R42051 VDD.n8990 VDD.n8989 0.0181836
R42052 VDD.n8792 VDD.n8791 0.0181836
R42053 VDD.n8785 VDD.n8784 0.0181836
R42054 VDD.n8729 VDD.n8728 0.0181836
R42055 VDD.n127 VDD.n126 0.0181836
R42056 VDD.n8613 VDD.n8612 0.0181836
R42057 VDD.n81 VDD.n80 0.0181836
R42058 VDD.n9130 VDD.n9128 0.0181276
R42059 VDD.n9132 VDD.n9128 0.0181276
R42060 VDD.n9133 VDD.n8459 0.0181276
R42061 VDD.n8081 VDD.n8079 0.0179831
R42062 VDD.n8075 VDD.n8074 0.0178367
R42063 VDD.n6037 VDD.n6036 0.0177463
R42064 VDD.n6169 VDD.n6157 0.0177463
R42065 VDD.n6850 VDD.n6849 0.0177463
R42066 VDD.n6727 VDD.n6726 0.0177463
R42067 VDD.n12563 VDD.n9 0.0176669
R42068 VDD.n8138 VDD.n8137 0.0175856
R42069 VDD.n8117 VDD.n8116 0.0175856
R42070 VDD.n8105 VDD.n8104 0.0175856
R42071 VDD.n5579 VDD.n5578 0.0175856
R42072 VDD.n5600 VDD.n5599 0.0175856
R42073 VDD.n5621 VDD.n5620 0.0175856
R42074 VDD.n5661 VDD.n5660 0.0175856
R42075 VDD.n5872 VDD.n5871 0.0175856
R42076 VDD.n5860 VDD.n5859 0.0175856
R42077 VDD.n5817 VDD.n5816 0.0175856
R42078 VDD.n5805 VDD.n5804 0.0175856
R42079 VDD.n5784 VDD.n5783 0.0175856
R42080 VDD.n5750 VDD.n5749 0.0175856
R42081 VDD.n5729 VDD.n5728 0.0175856
R42082 VDD.n11031 VDD.n1770 0.0175856
R42083 VDD.n9038 VDD.n9037 0.0175856
R42084 VDD.n9008 VDD.n9007 0.0175856
R42085 VDD.n8941 VDD.n8940 0.0175856
R42086 VDD.n8877 VDD.n8876 0.0175856
R42087 VDD.n8810 VDD.n8809 0.0175856
R42088 VDD.n8555 VDD.n8554 0.0175856
R42089 VDD.n186 VDD.n175 0.0175856
R42090 VDD.n9097 VDD.n9096 0.0175856
R42091 VDD.n9162 VDD.n9161 0.0175856
R42092 VDD.n142 VDD.n141 0.0175856
R42093 VDD.n12493 VDD.n12492 0.0175856
R42094 VDD.n12500 VDD.n95 0.0175856
R42095 VDD.n53 VDD.n52 0.0175856
R42096 VDD.n12549 VDD.n12548 0.0175856
R42097 VDD.n12594 VDD.n12593 0.0175856
R42098 VDD.n10797 VDD.n2007 0.0175462
R42099 VDD.n10855 VDD.n1934 0.0175462
R42100 VDD.n10910 VDD.n1907 0.0175462
R42101 VDD.n10965 VDD.n1842 0.0175462
R42102 VDD.n11020 VDD.n1780 0.0175462
R42103 VDD.n9064 VDD.n9063 0.0175462
R42104 VDD.n8891 VDD.n8890 0.0175462
R42105 VDD.n8748 VDD.n8747 0.0175462
R42106 VDD.n8698 VDD.n8697 0.0175462
R42107 VDD.n8639 VDD.n8638 0.0175462
R42108 VDD.n6699 VDD.n5262 0.0174226
R42109 VDD.n7124 VDD.n2322 0.0174226
R42110 VDD.n6361 VDD.n5472 0.0174226
R42111 VDD.n5445 VDD.n5444 0.0174226
R42112 VDD.n6379 VDD.n5361 0.0174226
R42113 VDD.n6699 VDD.n5263 0.0174226
R42114 VDD.n6380 VDD.n6379 0.0174226
R42115 VDD.n6361 VDD.n6360 0.0174226
R42116 VDD.n7143 VDD.n7142 0.0174226
R42117 VDD.n5444 VDD.n5433 0.0174226
R42118 VDD.n7142 VDD.n2310 0.0174226
R42119 VDD.n7124 VDD.n7123 0.0174226
R42120 VDD.n12440 VDD.n195 0.017375
R42121 VDD.n1664 VDD.n752 0.0172098
R42122 VDD.n1573 VDD.n1507 0.0172098
R42123 VDD.n1574 VDD.n1507 0.0172098
R42124 VDD.n1665 VDD.n752 0.0172098
R42125 VDD.n5262 VDD.n5222 0.0171298
R42126 VDD.n5260 VDD.n5222 0.0171298
R42127 VDD.n5260 VDD.n5259 0.0171298
R42128 VDD.n5259 VDD.n5258 0.0171298
R42129 VDD.n5258 VDD.n5225 0.0171298
R42130 VDD.n5255 VDD.n5225 0.0171298
R42131 VDD.n5255 VDD.n5254 0.0171298
R42132 VDD.n5254 VDD.n5253 0.0171298
R42133 VDD.n5252 VDD.n5227 0.0171298
R42134 VDD.n5250 VDD.n5227 0.0171298
R42135 VDD.n5248 VDD.n5247 0.0171298
R42136 VDD.n5247 VDD.n5230 0.0171298
R42137 VDD.n5245 VDD.n5230 0.0171298
R42138 VDD.n5244 VDD.n5231 0.0171298
R42139 VDD.n5242 VDD.n5231 0.0171298
R42140 VDD.n5242 VDD.n5241 0.0171298
R42141 VDD.n5241 VDD.n5240 0.0171298
R42142 VDD.n5240 VDD.n5234 0.0171298
R42143 VDD.n5237 VDD.n5234 0.0171298
R42144 VDD.n5237 VDD.n5236 0.0171298
R42145 VDD.n5236 VDD.n2322 0.0171298
R42146 VDD.n5472 VDD.n5379 0.0171298
R42147 VDD.n5470 VDD.n5379 0.0171298
R42148 VDD.n5470 VDD.n5469 0.0171298
R42149 VDD.n5469 VDD.n5468 0.0171298
R42150 VDD.n5468 VDD.n5382 0.0171298
R42151 VDD.n5465 VDD.n5382 0.0171298
R42152 VDD.n5465 VDD.n5464 0.0171298
R42153 VDD.n5464 VDD.n5463 0.0171298
R42154 VDD.n5462 VDD.n5384 0.0171298
R42155 VDD.n5460 VDD.n5384 0.0171298
R42156 VDD.n5458 VDD.n5457 0.0171298
R42157 VDD.n5457 VDD.n5387 0.0171298
R42158 VDD.n5455 VDD.n5387 0.0171298
R42159 VDD.n5454 VDD.n5388 0.0171298
R42160 VDD.n5452 VDD.n5388 0.0171298
R42161 VDD.n5452 VDD.n5451 0.0171298
R42162 VDD.n5451 VDD.n5450 0.0171298
R42163 VDD.n5450 VDD.n5391 0.0171298
R42164 VDD.n5447 VDD.n5391 0.0171298
R42165 VDD.n5447 VDD.n5446 0.0171298
R42166 VDD.n5446 VDD.n5445 0.0171298
R42167 VDD.n5361 VDD.n5321 0.0171298
R42168 VDD.n5359 VDD.n5321 0.0171298
R42169 VDD.n5359 VDD.n5358 0.0171298
R42170 VDD.n5358 VDD.n5357 0.0171298
R42171 VDD.n5357 VDD.n5324 0.0171298
R42172 VDD.n5354 VDD.n5324 0.0171298
R42173 VDD.n5354 VDD.n5353 0.0171298
R42174 VDD.n5353 VDD.n5352 0.0171298
R42175 VDD.n5351 VDD.n5326 0.0171298
R42176 VDD.n5349 VDD.n5326 0.0171298
R42177 VDD.n5347 VDD.n5346 0.0171298
R42178 VDD.n5346 VDD.n5329 0.0171298
R42179 VDD.n5344 VDD.n5329 0.0171298
R42180 VDD.n5343 VDD.n5330 0.0171298
R42181 VDD.n5341 VDD.n5330 0.0171298
R42182 VDD.n5341 VDD.n5340 0.0171298
R42183 VDD.n5340 VDD.n5339 0.0171298
R42184 VDD.n5339 VDD.n5333 0.0171298
R42185 VDD.n5336 VDD.n5333 0.0171298
R42186 VDD.n5336 VDD.n5335 0.0171298
R42187 VDD.n5335 VDD.n5263 0.0171298
R42188 VDD.n6010 VDD.n6009 0.0171298
R42189 VDD.n6007 VDD.n5989 0.0171298
R42190 VDD.n6005 VDD.n5989 0.0171298
R42191 VDD.n6005 VDD.n6004 0.0171298
R42192 VDD.n6004 VDD.n6003 0.0171298
R42193 VDD.n6003 VDD.n5992 0.0171298
R42194 VDD.n6000 VDD.n5992 0.0171298
R42195 VDD.n6000 VDD.n5999 0.0171298
R42196 VDD.n5999 VDD.n5998 0.0171298
R42197 VDD.n5997 VDD.n5995 0.0171298
R42198 VDD.n5995 VDD.n5313 0.0171298
R42199 VDD.n6393 VDD.n6392 0.0171298
R42200 VDD.n6392 VDD.n5315 0.0171298
R42201 VDD.n6390 VDD.n5315 0.0171298
R42202 VDD.n6389 VDD.n5316 0.0171298
R42203 VDD.n6387 VDD.n5316 0.0171298
R42204 VDD.n6387 VDD.n6386 0.0171298
R42205 VDD.n6386 VDD.n6385 0.0171298
R42206 VDD.n6385 VDD.n5319 0.0171298
R42207 VDD.n6382 VDD.n5319 0.0171298
R42208 VDD.n6382 VDD.n6381 0.0171298
R42209 VDD.n6381 VDD.n6380 0.0171298
R42210 VDD.n6330 VDD.n5486 0.0171298
R42211 VDD.n6331 VDD.n5485 0.0171298
R42212 VDD.n6333 VDD.n5485 0.0171298
R42213 VDD.n6333 VDD.n5484 0.0171298
R42214 VDD.n6336 VDD.n5484 0.0171298
R42215 VDD.n6336 VDD.n5483 0.0171298
R42216 VDD.n6339 VDD.n5483 0.0171298
R42217 VDD.n6339 VDD.n5482 0.0171298
R42218 VDD.n6341 VDD.n5482 0.0171298
R42219 VDD.n6342 VDD.n5480 0.0171298
R42220 VDD.n6344 VDD.n5480 0.0171298
R42221 VDD.n6347 VDD.n5479 0.0171298
R42222 VDD.n6347 VDD.n5478 0.0171298
R42223 VDD.n6349 VDD.n5478 0.0171298
R42224 VDD.n6350 VDD.n5477 0.0171298
R42225 VDD.n6352 VDD.n5477 0.0171298
R42226 VDD.n6352 VDD.n5476 0.0171298
R42227 VDD.n6355 VDD.n5476 0.0171298
R42228 VDD.n6355 VDD.n5475 0.0171298
R42229 VDD.n6358 VDD.n5475 0.0171298
R42230 VDD.n6358 VDD.n5474 0.0171298
R42231 VDD.n6360 VDD.n5474 0.0171298
R42232 VDD.n7143 VDD.n2309 0.0171298
R42233 VDD.n7145 VDD.n2309 0.0171298
R42234 VDD.n7145 VDD.n2308 0.0171298
R42235 VDD.n7148 VDD.n2308 0.0171298
R42236 VDD.n7148 VDD.n2307 0.0171298
R42237 VDD.n7151 VDD.n2307 0.0171298
R42238 VDD.n7151 VDD.n2306 0.0171298
R42239 VDD.n7153 VDD.n2306 0.0171298
R42240 VDD.n7154 VDD.n2304 0.0171298
R42241 VDD.n7156 VDD.n2304 0.0171298
R42242 VDD.n7159 VDD.n2303 0.0171298
R42243 VDD.n7159 VDD.n2302 0.0171298
R42244 VDD.n7161 VDD.n2302 0.0171298
R42245 VDD.n7162 VDD.n2301 0.0171298
R42246 VDD.n7164 VDD.n2301 0.0171298
R42247 VDD.n7164 VDD.n2300 0.0171298
R42248 VDD.n7167 VDD.n2300 0.0171298
R42249 VDD.n7167 VDD.n2299 0.0171298
R42250 VDD.n7170 VDD.n2299 0.0171298
R42251 VDD.n7170 VDD.n2298 0.0171298
R42252 VDD.n7172 VDD.n2298 0.0171298
R42253 VDD.n7173 VDD.n2297 0.0171298
R42254 VDD.n5433 VDD.n5393 0.0171298
R42255 VDD.n5431 VDD.n5393 0.0171298
R42256 VDD.n5431 VDD.n5430 0.0171298
R42257 VDD.n5430 VDD.n5429 0.0171298
R42258 VDD.n5429 VDD.n5396 0.0171298
R42259 VDD.n5426 VDD.n5396 0.0171298
R42260 VDD.n5426 VDD.n5425 0.0171298
R42261 VDD.n5425 VDD.n5424 0.0171298
R42262 VDD.n5423 VDD.n5398 0.0171298
R42263 VDD.n5421 VDD.n5398 0.0171298
R42264 VDD.n5419 VDD.n5418 0.0171298
R42265 VDD.n5418 VDD.n5401 0.0171298
R42266 VDD.n5416 VDD.n5401 0.0171298
R42267 VDD.n5415 VDD.n5402 0.0171298
R42268 VDD.n5413 VDD.n5402 0.0171298
R42269 VDD.n5413 VDD.n5412 0.0171298
R42270 VDD.n5412 VDD.n5411 0.0171298
R42271 VDD.n5411 VDD.n5405 0.0171298
R42272 VDD.n5408 VDD.n5405 0.0171298
R42273 VDD.n5408 VDD.n5407 0.0171298
R42274 VDD.n5407 VDD.n2310 0.0171298
R42275 VDD.n7123 VDD.n2324 0.0171298
R42276 VDD.n7121 VDD.n2324 0.0171298
R42277 VDD.n7121 VDD.n7120 0.0171298
R42278 VDD.n7120 VDD.n7119 0.0171298
R42279 VDD.n7119 VDD.n2327 0.0171298
R42280 VDD.n7116 VDD.n2327 0.0171298
R42281 VDD.n7116 VDD.n7115 0.0171298
R42282 VDD.n7115 VDD.n7114 0.0171298
R42283 VDD.n7113 VDD.n2329 0.0171298
R42284 VDD.n7111 VDD.n2329 0.0171298
R42285 VDD.n7109 VDD.n7108 0.0171298
R42286 VDD.n7108 VDD.n7089 0.0171298
R42287 VDD.n7106 VDD.n7089 0.0171298
R42288 VDD.n7105 VDD.n7090 0.0171298
R42289 VDD.n7103 VDD.n7090 0.0171298
R42290 VDD.n7103 VDD.n7102 0.0171298
R42291 VDD.n7102 VDD.n7101 0.0171298
R42292 VDD.n7101 VDD.n7093 0.0171298
R42293 VDD.n7098 VDD.n7093 0.0171298
R42294 VDD.n7098 VDD.n7097 0.0171298
R42295 VDD.n7097 VDD.n7096 0.0171298
R42296 VDD.n7095 VDD.n2240 0.0171298
R42297 VDD.n1530 VDD.n1523 0.0167842
R42298 VDD.n1531 VDD.n1522 0.0167842
R42299 VDD.n1532 VDD.n1522 0.0167842
R42300 VDD.n1547 VDD.n1546 0.0167842
R42301 VDD.n1545 VDD.n1534 0.0167842
R42302 VDD.n1544 VDD.n1534 0.0167842
R42303 VDD.n1543 VDD.n1535 0.0167842
R42304 VDD.n1672 VDD.n1671 0.016681
R42305 VDD.n4590 VDD.n4589 0.016625
R42306 VDD.n1582 VDD.n747 0.0165752
R42307 VDD.n1202 VDD.n1201 0.0164828
R42308 VDD.n1200 VDD.n1199 0.0164828
R42309 VDD.n1198 VDD.n1197 0.0164828
R42310 VDD.n1196 VDD.n1195 0.0164828
R42311 VDD.n1434 VDD.n1433 0.0164828
R42312 VDD.n1436 VDD.n1435 0.0164828
R42313 VDD.n1438 VDD.n1437 0.0164828
R42314 VDD.n1440 VDD.n1439 0.0164828
R42315 VDD.n1131 VDD.n1130 0.0164828
R42316 VDD.n1129 VDD.n1128 0.0164828
R42317 VDD.n1127 VDD.n1126 0.0164828
R42318 VDD.n1125 VDD.n1124 0.0164828
R42319 VDD.n872 VDD.n871 0.0164828
R42320 VDD.n870 VDD.n869 0.0164828
R42321 VDD.n868 VDD.n867 0.0164828
R42322 VDD.n866 VDD.n865 0.0164828
R42323 VDD.n801 VDD.n800 0.0164828
R42324 VDD.n799 VDD.n798 0.0164828
R42325 VDD.n797 VDD.n796 0.0164828
R42326 VDD.n795 VDD.n794 0.0164828
R42327 VDD.n1326 VDD.n1325 0.0164828
R42328 VDD.n1328 VDD.n1327 0.0164828
R42329 VDD.n1330 VDD.n1329 0.0164828
R42330 VDD.n1332 VDD.n1331 0.0164828
R42331 VDD.n838 VDD.n837 0.0164828
R42332 VDD.n836 VDD.n835 0.0164828
R42333 VDD.n834 VDD.n833 0.0164828
R42334 VDD.n832 VDD.n831 0.0164828
R42335 VDD.n1373 VDD.n1372 0.0164828
R42336 VDD.n1375 VDD.n1374 0.0164828
R42337 VDD.n1377 VDD.n1376 0.0164828
R42338 VDD.n1379 VDD.n1378 0.0164828
R42339 VDD.n1265 VDD.n1264 0.0164828
R42340 VDD.n1263 VDD.n1262 0.0164828
R42341 VDD.n1261 VDD.n1260 0.0164828
R42342 VDD.n1259 VDD.n1258 0.0164828
R42343 VDD.n1617 VDD.n1616 0.0164828
R42344 VDD.n1615 VDD.n1614 0.0164828
R42345 VDD.n1613 VDD.n1612 0.0164828
R42346 VDD.n1232 VDD.n1231 0.0164828
R42347 VDD.n1230 VDD.n1229 0.0164828
R42348 VDD.n1228 VDD.n1227 0.0164828
R42349 VDD.n1226 VDD.n1225 0.0164828
R42350 VDD.n1099 VDD.n1098 0.0164828
R42351 VDD.n1097 VDD.n1096 0.0164828
R42352 VDD.n1095 VDD.n813 0.0164828
R42353 VDD.n1475 VDD.n1474 0.0164828
R42354 VDD.n1473 VDD.n1472 0.0164828
R42355 VDD.n1471 VDD.n1470 0.0164828
R42356 VDD.n1469 VDD.n1468 0.0164828
R42357 VDD.n1294 VDD.n1293 0.0164828
R42358 VDD.n1296 VDD.n1295 0.0164828
R42359 VDD.n1298 VDD.n1297 0.0164828
R42360 VDD.n1300 VDD.n1299 0.0164828
R42361 VDD.n1706 VDD.n1705 0.0164828
R42362 VDD.n1704 VDD.n1703 0.0164828
R42363 VDD.n1702 VDD.n1701 0.0164828
R42364 VDD.n1700 VDD.n1699 0.0164828
R42365 VDD.n887 VDD.n886 0.0164828
R42366 VDD.n889 VDD.n888 0.0164828
R42367 VDD.n891 VDD.n890 0.0164828
R42368 VDD.n893 VDD.n892 0.0164828
R42369 VDD.n929 VDD.n928 0.0164828
R42370 VDD.n931 VDD.n930 0.0164828
R42371 VDD.n933 VDD.n932 0.0164828
R42372 VDD.n935 VDD.n934 0.0164828
R42373 VDD.n1049 VDD.n1048 0.0164828
R42374 VDD.n1051 VDD.n1050 0.0164828
R42375 VDD.n1053 VDD.n1052 0.0164828
R42376 VDD.n1055 VDD.n1054 0.0164828
R42377 VDD.n1153 VDD.n1152 0.0164828
R42378 VDD.n1151 VDD.n1150 0.0164828
R42379 VDD.n1149 VDD.n1148 0.0164828
R42380 VDD.n1147 VDD.n1146 0.0164828
R42381 VDD.n1724 VDD.n1723 0.0164828
R42382 VDD.n1726 VDD.n1725 0.0164828
R42383 VDD.n1728 VDD.n1727 0.0164828
R42384 VDD.n1730 VDD.n1729 0.0164828
R42385 VDD.n2136 VDD.n2135 0.0163144
R42386 VDD.n5253 VDD.n5252 0.01631
R42387 VDD.n5245 VDD.n5244 0.01631
R42388 VDD.n5463 VDD.n5462 0.01631
R42389 VDD.n5455 VDD.n5454 0.01631
R42390 VDD.n5352 VDD.n5351 0.01631
R42391 VDD.n5344 VDD.n5343 0.01631
R42392 VDD.n5998 VDD.n5997 0.01631
R42393 VDD.n6390 VDD.n6389 0.01631
R42394 VDD.n6342 VDD.n6341 0.01631
R42395 VDD.n6350 VDD.n6349 0.01631
R42396 VDD.n7154 VDD.n7153 0.01631
R42397 VDD.n7162 VDD.n7161 0.01631
R42398 VDD.n5424 VDD.n5423 0.01631
R42399 VDD.n5416 VDD.n5415 0.01631
R42400 VDD.n7114 VDD.n7113 0.01631
R42401 VDD.n7106 VDD.n7105 0.01631
R42402 VDD.n6562 VDD.n5287 0.0162238
R42403 VDD.n5298 VDD.n5297 0.0162238
R42404 VDD.n2385 VDD.n2384 0.0162238
R42405 VDD.n7025 VDD.n2374 0.0162238
R42406 VDD.n5363 VDD.n5362 0.0159138
R42407 VDD.n5365 VDD.n5364 0.0159138
R42408 VDD.n5367 VDD.n5366 0.0159138
R42409 VDD.n5370 VDD.n5369 0.0159138
R42410 VDD.n5372 VDD.n5371 0.0159138
R42411 VDD.n5374 VDD.n5373 0.0159138
R42412 VDD.n6378 VDD.n6377 0.0159138
R42413 VDD.n6376 VDD.n6375 0.0159138
R42414 VDD.n6374 VDD.n6373 0.0159138
R42415 VDD.n6216 VDD.n5375 0.0159138
R42416 VDD.n6218 VDD.n6217 0.0159138
R42417 VDD.n6265 VDD.n6264 0.0159138
R42418 VDD.n6263 VDD.n5377 0.0159138
R42419 VDD.n6367 VDD.n6366 0.0159138
R42420 VDD.n6365 VDD.n6364 0.0159138
R42421 VDD.n6363 VDD.n6362 0.0159138
R42422 VDD.n5937 VDD.n5473 0.0159138
R42423 VDD.n5939 VDD.n5938 0.0159138
R42424 VDD.n5941 VDD.n5940 0.0159138
R42425 VDD.n5945 VDD.n5944 0.0159138
R42426 VDD.n5947 VDD.n5946 0.0159138
R42427 VDD.n5949 VDD.n5948 0.0159138
R42428 VDD.n2358 VDD.n2341 0.0159138
R42429 VDD.n2360 VDD.n2359 0.0159138
R42430 VDD.n2365 VDD.n2364 0.0159138
R42431 VDD.n2363 VDD.n2362 0.0159138
R42432 VDD.n2361 VDD.n2311 0.0159138
R42433 VDD.n7141 VDD.n7140 0.0159138
R42434 VDD.n7139 VDD.n7138 0.0159138
R42435 VDD.n7137 VDD.n7136 0.0159138
R42436 VDD.n2316 VDD.n2315 0.0159138
R42437 VDD.n2314 VDD.n2313 0.0159138
R42438 VDD.n2401 VDD.n2400 0.0159138
R42439 VDD.n2399 VDD.n2398 0.0159138
R42440 VDD.n2397 VDD.n2320 0.0159138
R42441 VDD.n7130 VDD.n7129 0.0159138
R42442 VDD.n7128 VDD.n7127 0.0159138
R42443 VDD.n7126 VDD.n7125 0.0159138
R42444 VDD.n2343 VDD.n2323 0.0159138
R42445 VDD.n2345 VDD.n2344 0.0159138
R42446 VDD.n2347 VDD.n2346 0.0159138
R42447 VDD.n7045 VDD.n7044 0.0159138
R42448 VDD.n7047 VDD.n7046 0.0159138
R42449 VDD.n1205 VDD.n1204 0.0159138
R42450 VDD.n1203 VDD.n1190 0.0159138
R42451 VDD.n1202 VDD.n1190 0.0159138
R42452 VDD.n1201 VDD.n1191 0.0159138
R42453 VDD.n1200 VDD.n1191 0.0159138
R42454 VDD.n1199 VDD.n1192 0.0159138
R42455 VDD.n1198 VDD.n1192 0.0159138
R42456 VDD.n1197 VDD.n1193 0.0159138
R42457 VDD.n1196 VDD.n1193 0.0159138
R42458 VDD.n1195 VDD.n1194 0.0159138
R42459 VDD.n1194 VDD.n851 0.0159138
R42460 VDD.n1432 VDD.n843 0.0159138
R42461 VDD.n1433 VDD.n843 0.0159138
R42462 VDD.n1434 VDD.n842 0.0159138
R42463 VDD.n1435 VDD.n842 0.0159138
R42464 VDD.n1436 VDD.n841 0.0159138
R42465 VDD.n1437 VDD.n841 0.0159138
R42466 VDD.n1438 VDD.n840 0.0159138
R42467 VDD.n1439 VDD.n840 0.0159138
R42468 VDD.n1134 VDD.n1133 0.0159138
R42469 VDD.n1132 VDD.n1119 0.0159138
R42470 VDD.n1131 VDD.n1119 0.0159138
R42471 VDD.n1130 VDD.n1120 0.0159138
R42472 VDD.n1129 VDD.n1120 0.0159138
R42473 VDD.n1128 VDD.n1121 0.0159138
R42474 VDD.n1127 VDD.n1121 0.0159138
R42475 VDD.n1126 VDD.n1122 0.0159138
R42476 VDD.n1125 VDD.n1122 0.0159138
R42477 VDD.n1124 VDD.n1123 0.0159138
R42478 VDD.n1123 VDD.n852 0.0159138
R42479 VDD.n873 VDD.n860 0.0159138
R42480 VDD.n872 VDD.n860 0.0159138
R42481 VDD.n871 VDD.n861 0.0159138
R42482 VDD.n870 VDD.n861 0.0159138
R42483 VDD.n869 VDD.n862 0.0159138
R42484 VDD.n868 VDD.n862 0.0159138
R42485 VDD.n867 VDD.n863 0.0159138
R42486 VDD.n866 VDD.n863 0.0159138
R42487 VDD.n865 VDD.n864 0.0159138
R42488 VDD.n864 VDD.n728 0.0159138
R42489 VDD.n802 VDD.n788 0.0159138
R42490 VDD.n801 VDD.n788 0.0159138
R42491 VDD.n800 VDD.n789 0.0159138
R42492 VDD.n799 VDD.n789 0.0159138
R42493 VDD.n798 VDD.n790 0.0159138
R42494 VDD.n797 VDD.n790 0.0159138
R42495 VDD.n796 VDD.n791 0.0159138
R42496 VDD.n795 VDD.n791 0.0159138
R42497 VDD.n794 VDD.n792 0.0159138
R42498 VDD.n793 VDD.n792 0.0159138
R42499 VDD.n1324 VDD.n745 0.0159138
R42500 VDD.n1325 VDD.n1324 0.0159138
R42501 VDD.n1326 VDD.n1323 0.0159138
R42502 VDD.n1327 VDD.n1323 0.0159138
R42503 VDD.n1328 VDD.n1322 0.0159138
R42504 VDD.n1329 VDD.n1322 0.0159138
R42505 VDD.n1330 VDD.n1321 0.0159138
R42506 VDD.n1331 VDD.n1321 0.0159138
R42507 VDD.n1332 VDD.n1320 0.0159138
R42508 VDD.n1333 VDD.n1320 0.0159138
R42509 VDD.n1334 VDD.n1319 0.0159138
R42510 VDD.n839 VDD.n825 0.0159138
R42511 VDD.n838 VDD.n825 0.0159138
R42512 VDD.n837 VDD.n826 0.0159138
R42513 VDD.n836 VDD.n826 0.0159138
R42514 VDD.n835 VDD.n827 0.0159138
R42515 VDD.n834 VDD.n827 0.0159138
R42516 VDD.n833 VDD.n828 0.0159138
R42517 VDD.n832 VDD.n828 0.0159138
R42518 VDD.n831 VDD.n829 0.0159138
R42519 VDD.n830 VDD.n829 0.0159138
R42520 VDD.n1371 VDD.n1370 0.0159138
R42521 VDD.n1372 VDD.n1370 0.0159138
R42522 VDD.n1373 VDD.n1369 0.0159138
R42523 VDD.n1374 VDD.n1369 0.0159138
R42524 VDD.n1375 VDD.n1368 0.0159138
R42525 VDD.n1376 VDD.n1368 0.0159138
R42526 VDD.n1377 VDD.n1367 0.0159138
R42527 VDD.n1378 VDD.n1367 0.0159138
R42528 VDD.n1379 VDD.n1366 0.0159138
R42529 VDD.n1380 VDD.n1366 0.0159138
R42530 VDD.n1381 VDD.n1365 0.0159138
R42531 VDD.n1268 VDD.n1267 0.0159138
R42532 VDD.n1266 VDD.n1252 0.0159138
R42533 VDD.n1265 VDD.n1252 0.0159138
R42534 VDD.n1264 VDD.n1253 0.0159138
R42535 VDD.n1263 VDD.n1253 0.0159138
R42536 VDD.n1262 VDD.n1254 0.0159138
R42537 VDD.n1261 VDD.n1254 0.0159138
R42538 VDD.n1260 VDD.n1255 0.0159138
R42539 VDD.n1259 VDD.n1255 0.0159138
R42540 VDD.n1258 VDD.n1256 0.0159138
R42541 VDD.n1257 VDD.n1256 0.0159138
R42542 VDD.n1618 VDD.n785 0.0159138
R42543 VDD.n1617 VDD.n785 0.0159138
R42544 VDD.n1616 VDD.n786 0.0159138
R42545 VDD.n1615 VDD.n786 0.0159138
R42546 VDD.n1614 VDD.n787 0.0159138
R42547 VDD.n1613 VDD.n787 0.0159138
R42548 VDD.n1235 VDD.n1234 0.0159138
R42549 VDD.n1233 VDD.n1220 0.0159138
R42550 VDD.n1232 VDD.n1220 0.0159138
R42551 VDD.n1231 VDD.n1221 0.0159138
R42552 VDD.n1230 VDD.n1221 0.0159138
R42553 VDD.n1229 VDD.n1222 0.0159138
R42554 VDD.n1228 VDD.n1222 0.0159138
R42555 VDD.n1227 VDD.n1223 0.0159138
R42556 VDD.n1226 VDD.n1223 0.0159138
R42557 VDD.n1225 VDD.n1224 0.0159138
R42558 VDD.n1224 VDD.n1085 0.0159138
R42559 VDD.n1100 VDD.n1092 0.0159138
R42560 VDD.n1099 VDD.n1092 0.0159138
R42561 VDD.n1098 VDD.n1093 0.0159138
R42562 VDD.n1097 VDD.n1093 0.0159138
R42563 VDD.n1096 VDD.n1094 0.0159138
R42564 VDD.n1095 VDD.n1094 0.0159138
R42565 VDD.n1476 VDD.n1462 0.0159138
R42566 VDD.n1475 VDD.n1462 0.0159138
R42567 VDD.n1474 VDD.n1463 0.0159138
R42568 VDD.n1473 VDD.n1463 0.0159138
R42569 VDD.n1472 VDD.n1464 0.0159138
R42570 VDD.n1471 VDD.n1464 0.0159138
R42571 VDD.n1470 VDD.n1465 0.0159138
R42572 VDD.n1469 VDD.n1465 0.0159138
R42573 VDD.n1468 VDD.n1466 0.0159138
R42574 VDD.n1467 VDD.n1466 0.0159138
R42575 VDD.n1292 VDD.n742 0.0159138
R42576 VDD.n1293 VDD.n1292 0.0159138
R42577 VDD.n1294 VDD.n1291 0.0159138
R42578 VDD.n1295 VDD.n1291 0.0159138
R42579 VDD.n1296 VDD.n1290 0.0159138
R42580 VDD.n1297 VDD.n1290 0.0159138
R42581 VDD.n1298 VDD.n1289 0.0159138
R42582 VDD.n1299 VDD.n1289 0.0159138
R42583 VDD.n1300 VDD.n1288 0.0159138
R42584 VDD.n1301 VDD.n1288 0.0159138
R42585 VDD.n1302 VDD.n1287 0.0159138
R42586 VDD.n1707 VDD.n730 0.0159138
R42587 VDD.n1706 VDD.n730 0.0159138
R42588 VDD.n1705 VDD.n731 0.0159138
R42589 VDD.n1704 VDD.n731 0.0159138
R42590 VDD.n1703 VDD.n732 0.0159138
R42591 VDD.n1702 VDD.n732 0.0159138
R42592 VDD.n1701 VDD.n733 0.0159138
R42593 VDD.n1700 VDD.n733 0.0159138
R42594 VDD.n1699 VDD.n734 0.0159138
R42595 VDD.n1698 VDD.n734 0.0159138
R42596 VDD.n885 VDD.n884 0.0159138
R42597 VDD.n886 VDD.n884 0.0159138
R42598 VDD.n887 VDD.n883 0.0159138
R42599 VDD.n888 VDD.n883 0.0159138
R42600 VDD.n889 VDD.n882 0.0159138
R42601 VDD.n890 VDD.n882 0.0159138
R42602 VDD.n891 VDD.n881 0.0159138
R42603 VDD.n892 VDD.n881 0.0159138
R42604 VDD.n893 VDD.n880 0.0159138
R42605 VDD.n894 VDD.n880 0.0159138
R42606 VDD.n895 VDD.n879 0.0159138
R42607 VDD.n927 VDD.n699 0.0159138
R42608 VDD.n928 VDD.n927 0.0159138
R42609 VDD.n929 VDD.n926 0.0159138
R42610 VDD.n930 VDD.n926 0.0159138
R42611 VDD.n931 VDD.n925 0.0159138
R42612 VDD.n932 VDD.n925 0.0159138
R42613 VDD.n933 VDD.n924 0.0159138
R42614 VDD.n934 VDD.n924 0.0159138
R42615 VDD.n935 VDD.n923 0.0159138
R42616 VDD.n936 VDD.n923 0.0159138
R42617 VDD.n1047 VDD.n922 0.0159138
R42618 VDD.n1048 VDD.n922 0.0159138
R42619 VDD.n1049 VDD.n921 0.0159138
R42620 VDD.n1050 VDD.n921 0.0159138
R42621 VDD.n1051 VDD.n920 0.0159138
R42622 VDD.n1052 VDD.n920 0.0159138
R42623 VDD.n1053 VDD.n919 0.0159138
R42624 VDD.n1054 VDD.n919 0.0159138
R42625 VDD.n1055 VDD.n918 0.0159138
R42626 VDD.n1056 VDD.n918 0.0159138
R42627 VDD.n1057 VDD.n917 0.0159138
R42628 VDD.n1156 VDD.n1155 0.0159138
R42629 VDD.n1154 VDD.n1140 0.0159138
R42630 VDD.n1153 VDD.n1140 0.0159138
R42631 VDD.n1152 VDD.n1141 0.0159138
R42632 VDD.n1151 VDD.n1141 0.0159138
R42633 VDD.n1150 VDD.n1142 0.0159138
R42634 VDD.n1149 VDD.n1142 0.0159138
R42635 VDD.n1148 VDD.n1143 0.0159138
R42636 VDD.n1147 VDD.n1143 0.0159138
R42637 VDD.n1146 VDD.n1144 0.0159138
R42638 VDD.n1145 VDD.n1144 0.0159138
R42639 VDD.n1722 VDD.n705 0.0159138
R42640 VDD.n1723 VDD.n705 0.0159138
R42641 VDD.n1724 VDD.n704 0.0159138
R42642 VDD.n1725 VDD.n704 0.0159138
R42643 VDD.n1726 VDD.n703 0.0159138
R42644 VDD.n1727 VDD.n703 0.0159138
R42645 VDD.n1728 VDD.n702 0.0159138
R42646 VDD.n1729 VDD.n702 0.0159138
R42647 VDD.n1730 VDD.n701 0.0159138
R42648 VDD.n1731 VDD.n701 0.0159138
R42649 VDD.n8137 VDD.n8136 0.0159011
R42650 VDD.n8116 VDD.n8115 0.0159011
R42651 VDD.n8104 VDD.n8103 0.0159011
R42652 VDD.n5580 VDD.n5579 0.0159011
R42653 VDD.n5601 VDD.n5600 0.0159011
R42654 VDD.n5622 VDD.n5621 0.0159011
R42655 VDD.n5662 VDD.n5661 0.0159011
R42656 VDD.n5871 VDD.n5870 0.0159011
R42657 VDD.n5859 VDD.n5858 0.0159011
R42658 VDD.n5816 VDD.n5815 0.0159011
R42659 VDD.n5804 VDD.n5803 0.0159011
R42660 VDD.n5783 VDD.n5782 0.0159011
R42661 VDD.n5749 VDD.n5748 0.0159011
R42662 VDD.n5728 VDD.n5727 0.0159011
R42663 VDD.n11032 VDD.n11031 0.0159011
R42664 VDD.n9037 VDD.n8490 0.0159011
R42665 VDD.n9008 VDD.n8951 0.0159011
R42666 VDD.n8940 VDD.n8507 0.0159011
R42667 VDD.n8877 VDD.n8842 0.0159011
R42668 VDD.n8809 VDD.n8526 0.0159011
R42669 VDD.n8554 VDD.n8553 0.0159011
R42670 VDD.n175 VDD.n174 0.0159011
R42671 VDD.n9096 VDD.n9095 0.0159011
R42672 VDD.n9161 VDD.n8472 0.0159011
R42673 VDD.n141 VDD.n140 0.0159011
R42674 VDD.n12494 VDD.n12493 0.0159011
R42675 VDD.n95 VDD.n94 0.0159011
R42676 VDD.n52 VDD.n51 0.0159011
R42677 VDD.n12550 VDD.n12549 0.0159011
R42678 VDD.n12593 VDD.n12591 0.0159011
R42679 VDD.n10149 VDD.n10148 0.015875
R42680 VDD.n2134 VDD.n2133 0.0156839
R42681 VDD.n2137 VDD.n2136 0.0154737
R42682 VDD.n6180 VDD.n6179 0.0154453
R42683 VDD.n6320 VDD.n6318 0.0153631
R42684 VDD.n5250 VDD.n5249 0.015256
R42685 VDD.n5460 VDD.n5459 0.015256
R42686 VDD.n5349 VDD.n5348 0.015256
R42687 VDD.n6394 VDD.n5313 0.015256
R42688 VDD.n6344 VDD.n5481 0.015256
R42689 VDD.n7156 VDD.n2305 0.015256
R42690 VDD.n5421 VDD.n5420 0.015256
R42691 VDD.n7111 VDD.n7110 0.015256
R42692 VDD.n2163 VDD.n2162 0.0148793
R42693 VDD.n1548 VDD.n1533 0.014653
R42694 VDD.n1495 VDD.n1494 0.0142459
R42695 VDD.n1607 VDD.n1606 0.0142459
R42696 VDD.n1595 VDD.n1594 0.0142459
R42697 VDD.n1711 VDD.n1710 0.0142459
R42698 VDD.n1398 VDD.n1397 0.0142459
R42699 VDD.n1407 VDD.n1406 0.0142459
R42700 VDD.n1445 VDD.n1444 0.0142459
R42701 VDD.n1460 VDD.n1459 0.0142459
R42702 VDD.n1483 VDD.n1482 0.0142459
R42703 VDD.n1735 VDD.n1734 0.0142459
R42704 VDD.n720 VDD.n719 0.0142459
R42705 VDD.n2161 VDD.n2160 0.0142069
R42706 VDD.n6714 VDD.n2406 0.0141364
R42707 VDD.n6700 VDD.n6699 0.0138734
R42708 VDD.n5444 VDD.n5438 0.0138734
R42709 VDD.n8015 VDD.n8014 0.0138448
R42710 VDD.n6699 VDD.n6698 0.0138425
R42711 VDD.n5444 VDD.n5443 0.0138425
R42712 VDD.n1559 VDD.n1558 0.0137787
R42713 VDD.n1554 VDD.n1517 0.0137787
R42714 VDD.n6190 VDD.n6010 0.0137336
R42715 VDD.n5487 VDD.n5486 0.0137336
R42716 VDD.n10777 VDD.n2020 0.0136837
R42717 VDD.n10784 VDD.n2010 0.0136837
R42718 VDD.n10835 VDD.n1947 0.0136837
R42719 VDD.n10842 VDD.n1937 0.0136837
R42720 VDD.n10897 VDD.n1910 0.0136837
R42721 VDD.n10945 VDD.n1855 0.0136837
R42722 VDD.n10952 VDD.n1845 0.0136837
R42723 VDD.n11000 VDD.n1790 0.0136837
R42724 VDD.n11007 VDD.n1783 0.0136837
R42725 VDD.n9053 VDD.n9052 0.0136837
R42726 VDD.n8919 VDD.n8918 0.0136837
R42727 VDD.n8861 VDD.n8858 0.0136837
R42728 VDD.n8570 VDD.n8569 0.0136837
R42729 VDD.n9177 VDD.n9176 0.0136837
R42730 VDD.n12459 VDD.n12458 0.0136837
R42731 VDD.n12477 VDD.n12474 0.0136837
R42732 VDD.n12515 VDD.n12514 0.0136837
R42733 VDD.n12533 VDD.n12530 0.0136837
R42734 VDD.n12609 VDD.n12608 0.0136837
R42735 VDD.n10828 VDD.n1993 0.013561
R42736 VDD.n10883 VDD.n1928 0.013561
R42737 VDD.n10938 VDD.n1901 0.013561
R42738 VDD.n10993 VDD.n1836 0.013561
R42739 VDD.n8988 VDD.n8985 0.013561
R42740 VDD.n8788 VDD.n8787 0.013561
R42741 VDD.n12467 VDD.n122 0.013561
R42742 VDD.n12523 VDD.n42 0.013561
R42743 VDD.n1537 VDD.n1512 0.0133852
R42744 VDD.n1553 VDD.n1518 0.0133852
R42745 VDD.n1752 VDD.n682 0.0131331
R42746 VDD.n996 VDD.n995 0.0131331
R42747 VDD.n1007 VDD.n1006 0.0131331
R42748 VDD.n7822 VDD.n2242 0.012875
R42749 VDD.n11872 VDD.n384 0.012875
R42750 VDD.n6601 VDD.n6599 0.012725
R42751 VDD.n952 VDD.n951 0.0126485
R42752 VDD.n6709 VDD.n6708 0.0125453
R42753 VDD.n6704 VDD.n6703 0.0125453
R42754 VDD.n6695 VDD.n6694 0.0125453
R42755 VDD.n6690 VDD.n6689 0.0125453
R42756 VDD.n6638 VDD.n6637 0.0125453
R42757 VDD.n5435 VDD.n5434 0.0125453
R42758 VDD.n5440 VDD.n5439 0.0125453
R42759 VDD.n6629 VDD.n6628 0.0125453
R42760 VDD.n1495 VDD.n805 0.0124383
R42761 VDD.n1496 VDD.n805 0.0124383
R42762 VDD.n1608 VDD.n1497 0.0124383
R42763 VDD.n1607 VDD.n1497 0.0124383
R42764 VDD.n1606 VDD.n1498 0.0124383
R42765 VDD.n1605 VDD.n1498 0.0124383
R42766 VDD.n1604 VDD.n1499 0.0124383
R42767 VDD.n1602 VDD.n1499 0.0124383
R42768 VDD.n1602 VDD.n1601 0.0124383
R42769 VDD.n1599 VDD.n1502 0.0124383
R42770 VDD.n1597 VDD.n1502 0.0124383
R42771 VDD.n1596 VDD.n1503 0.0124383
R42772 VDD.n1595 VDD.n1503 0.0124383
R42773 VDD.n1594 VDD.n1504 0.0124383
R42774 VDD.n1710 VDD.n727 0.0124383
R42775 VDD.n1709 VDD.n727 0.0124383
R42776 VDD.n1396 VDD.n729 0.0124383
R42777 VDD.n1397 VDD.n1396 0.0124383
R42778 VDD.n1398 VDD.n1395 0.0124383
R42779 VDD.n1399 VDD.n1395 0.0124383
R42780 VDD.n1400 VDD.n1394 0.0124383
R42781 VDD.n1402 VDD.n1394 0.0124383
R42782 VDD.n1402 VDD.n1391 0.0124383
R42783 VDD.n1411 VDD.n1393 0.0124383
R42784 VDD.n1409 VDD.n1393 0.0124383
R42785 VDD.n1408 VDD.n1404 0.0124383
R42786 VDD.n1407 VDD.n1404 0.0124383
R42787 VDD.n1406 VDD.n1405 0.0124383
R42788 VDD.n1405 VDD.n824 0.0124383
R42789 VDD.n1443 VDD.n822 0.0124383
R42790 VDD.n1444 VDD.n822 0.0124383
R42791 VDD.n1446 VDD.n1445 0.0124383
R42792 VDD.n1450 VDD.n819 0.0124383
R42793 VDD.n1452 VDD.n819 0.0124383
R42794 VDD.n1452 VDD.n820 0.0124383
R42795 VDD.n1455 VDD.n817 0.0124383
R42796 VDD.n1457 VDD.n817 0.0124383
R42797 VDD.n1458 VDD.n816 0.0124383
R42798 VDD.n1459 VDD.n816 0.0124383
R42799 VDD.n1460 VDD.n815 0.0124383
R42800 VDD.n1461 VDD.n815 0.0124383
R42801 VDD.n1481 VDD.n812 0.0124383
R42802 VDD.n1482 VDD.n812 0.0124383
R42803 VDD.n1483 VDD.n811 0.0124383
R42804 VDD.n1484 VDD.n811 0.0124383
R42805 VDD.n1485 VDD.n809 0.0124383
R42806 VDD.n1487 VDD.n809 0.0124383
R42807 VDD.n1487 VDD.n810 0.0124383
R42808 VDD.n1490 VDD.n807 0.0124383
R42809 VDD.n1492 VDD.n807 0.0124383
R42810 VDD.n1493 VDD.n806 0.0124383
R42811 VDD.n1494 VDD.n806 0.0124383
R42812 VDD.n951 VDD.n943 0.0124383
R42813 VDD.n950 VDD.n943 0.0124383
R42814 VDD.n948 VDD.n944 0.0124383
R42815 VDD.n946 VDD.n944 0.0124383
R42816 VDD.n946 VDD.n693 0.0124383
R42817 VDD.n1739 VDD.n695 0.0124383
R42818 VDD.n1737 VDD.n695 0.0124383
R42819 VDD.n1735 VDD.n697 0.0124383
R42820 VDD.n1734 VDD.n698 0.0124383
R42821 VDD.n1733 VDD.n698 0.0124383
R42822 VDD.n718 VDD.n700 0.0124383
R42823 VDD.n719 VDD.n718 0.0124383
R42824 VDD.n720 VDD.n717 0.0124383
R42825 VDD.n721 VDD.n717 0.0124383
R42826 VDD.n722 VDD.n716 0.0124383
R42827 VDD.n724 VDD.n716 0.0124383
R42828 VDD.n724 VDD.n713 0.0124383
R42829 VDD.n1715 VDD.n715 0.0124383
R42830 VDD.n1713 VDD.n715 0.0124383
R42831 VDD.n1712 VDD.n726 0.0124383
R42832 VDD.n1711 VDD.n726 0.0124383
R42833 VDD.n9183 VDD.n8459 0.0123552
R42834 VDD.n1005 VDD.n1004 0.0120089
R42835 VDD.n2138 VDD.n2137 0.0119536
R42836 VDD.n2135 VDD.n2134 0.0119536
R42837 VDD.n2133 VDD.n2132 0.0119536
R42838 VDD.n1605 VDD.n1604 0.0118498
R42839 VDD.n1600 VDD.n1599 0.0118498
R42840 VDD.n1597 VDD.n1596 0.0118498
R42841 VDD.n1400 VDD.n1399 0.0118498
R42842 VDD.n1412 VDD.n1411 0.0118498
R42843 VDD.n1409 VDD.n1408 0.0118498
R42844 VDD.n1455 VDD.n818 0.0118498
R42845 VDD.n1458 VDD.n1457 0.0118498
R42846 VDD.n1485 VDD.n1484 0.0118498
R42847 VDD.n1490 VDD.n808 0.0118498
R42848 VDD.n1493 VDD.n1492 0.0118498
R42849 VDD.n1740 VDD.n1739 0.0118498
R42850 VDD.n1737 VDD.n1736 0.0118498
R42851 VDD.n722 VDD.n721 0.0118498
R42852 VDD.n1716 VDD.n1715 0.0118498
R42853 VDD.n1713 VDD.n1712 0.0118498
R42854 VDD.n8067 VDD.n8066 0.0117759
R42855 VDD.n2156 VDD.n2147 0.0117759
R42856 VDD.n2165 VDD.n2164 0.0117759
R42857 VDD.n8016 VDD.n8015 0.0117759
R42858 VDD.n2130 VDD.n2129 0.0116909
R42859 VDD.n1610 VDD.n1496 0.0115976
R42860 VDD.n1610 VDD.n1608 0.0115976
R42861 VDD.n1709 VDD.n1708 0.0115976
R42862 VDD.n1708 VDD.n729 0.0115976
R42863 VDD.n1442 VDD.n824 0.0115976
R42864 VDD.n1443 VDD.n1442 0.0115976
R42865 VDD.n1480 VDD.n1461 0.0115976
R42866 VDD.n1481 VDD.n1480 0.0115976
R42867 VDD.n1733 VDD.n1732 0.0115976
R42868 VDD.n1732 VDD.n700 0.0115976
R42869 VDD.n9134 VDD.n9133 0.0114862
R42870 VDD.n1022 VDD.n1 0.0114467
R42871 VDD.n6297 VDD.n6296 0.0113718
R42872 VDD.n6269 VDD.n6268 0.0113718
R42873 VDD.n6261 VDD.n6260 0.0113718
R42874 VDD.n6657 VDD.n6656 0.0113718
R42875 VDD.n7051 VDD.n7050 0.0113718
R42876 VDD.n10777 VDD.n2023 0.0113038
R42877 VDD.n10787 VDD.n10784 0.0113038
R42878 VDD.n10835 VDD.n1950 0.0113038
R42879 VDD.n10845 VDD.n10842 0.0113038
R42880 VDD.n10900 VDD.n10897 0.0113038
R42881 VDD.n10945 VDD.n1858 0.0113038
R42882 VDD.n10955 VDD.n10952 0.0113038
R42883 VDD.n11000 VDD.n1793 0.0113038
R42884 VDD.n11010 VDD.n11007 0.0113038
R42885 VDD.n9055 VDD.n9053 0.0113038
R42886 VDD.n8921 VDD.n8919 0.0113038
R42887 VDD.n8858 VDD.n8857 0.0113038
R42888 VDD.n8572 VDD.n8570 0.0113038
R42889 VDD.n9177 VDD.n8465 0.0113038
R42890 VDD.n12459 VDD.n180 0.0113038
R42891 VDD.n12474 VDD.n109 0.0113038
R42892 VDD.n12515 VDD.n100 0.0113038
R42893 VDD.n12530 VDD.n29 0.0113038
R42894 VDD.n12609 VDD.n20 0.0113038
R42895 VDD.n10828 VDD.n10827 0.0112032
R42896 VDD.n10883 VDD.n10882 0.0112032
R42897 VDD.n10938 VDD.n10937 0.0112032
R42898 VDD.n10993 VDD.n10992 0.0112032
R42899 VDD.n8985 VDD.n8984 0.0112032
R42900 VDD.n8790 VDD.n8788 0.0112032
R42901 VDD.n12467 VDD.n119 0.0112032
R42902 VDD.n12523 VDD.n39 0.0112032
R42903 VDD.n2158 VDD.n2157 0.0111034
R42904 VDD.n8142 VDD.n8141 0.0109679
R42905 VDD.n5555 VDD.n5554 0.0109679
R42906 VDD.n5546 VDD.n5545 0.0109679
R42907 VDD.n5821 VDD.n5820 0.0109679
R42908 VDD.n5754 VDD.n5753 0.0109679
R42909 VDD.n9002 VDD.n8970 0.0109679
R42910 VDD.n8831 VDD.n8830 0.0109679
R42911 VDD.n9118 VDD.n9117 0.0109679
R42912 VDD.n163 VDD.n162 0.0109679
R42913 VDD.n74 VDD.n73 0.0109679
R42914 VDD.n5202 VDD.n5201 0.0109148
R42915 VDD.n5201 VDD.n2408 0.0109148
R42916 VDD.n1569 VDD.n1568 0.0108543
R42917 VDD.n7175 VDD.n7174 0.0108058
R42918 VDD.n7827 VDD.n2241 0.0108058
R42919 VDD.n1661 VDD.n754 0.0106739
R42920 VDD.n1643 VDD.n768 0.0106739
R42921 VDD.n1447 VDD.n1446 0.0102524
R42922 VDD.n6685 VDD.n5265 0.0101084
R42923 VDD.n6685 VDD.n6684 0.0101084
R42924 VDD.n7760 VDD.n2265 0.0101084
R42925 VDD.n6297 VDD.n6200 0.00994219
R42926 VDD.n6296 VDD.n6201 0.00994219
R42927 VDD.n6294 VDD.n6201 0.00994219
R42928 VDD.n6294 VDD.n6293 0.00994219
R42929 VDD.n6293 VDD.n6292 0.00994219
R42930 VDD.n6292 VDD.n6204 0.00994219
R42931 VDD.n6289 VDD.n6204 0.00994219
R42932 VDD.n6289 VDD.n6288 0.00994219
R42933 VDD.n6288 VDD.n6287 0.00994219
R42934 VDD.n6286 VDD.n6206 0.00994219
R42935 VDD.n6284 VDD.n6206 0.00994219
R42936 VDD.n6282 VDD.n6281 0.00994219
R42937 VDD.n6281 VDD.n6209 0.00994219
R42938 VDD.n6279 VDD.n6209 0.00994219
R42939 VDD.n6278 VDD.n6210 0.00994219
R42940 VDD.n6276 VDD.n6210 0.00994219
R42941 VDD.n6276 VDD.n6275 0.00994219
R42942 VDD.n6275 VDD.n6274 0.00994219
R42943 VDD.n6274 VDD.n6213 0.00994219
R42944 VDD.n6271 VDD.n6213 0.00994219
R42945 VDD.n6271 VDD.n6270 0.00994219
R42946 VDD.n6270 VDD.n6269 0.00994219
R42947 VDD.n6268 VDD.n6215 0.00994219
R42948 VDD.n6267 VDD.n6215 0.00994219
R42949 VDD.n6262 VDD.n6219 0.00994219
R42950 VDD.n6261 VDD.n6219 0.00994219
R42951 VDD.n6260 VDD.n6220 0.00994219
R42952 VDD.n6258 VDD.n6220 0.00994219
R42953 VDD.n6258 VDD.n6257 0.00994219
R42954 VDD.n6257 VDD.n6256 0.00994219
R42955 VDD.n6256 VDD.n6223 0.00994219
R42956 VDD.n6253 VDD.n6223 0.00994219
R42957 VDD.n6253 VDD.n6252 0.00994219
R42958 VDD.n6252 VDD.n6251 0.00994219
R42959 VDD.n6250 VDD.n6225 0.00994219
R42960 VDD.n6248 VDD.n6225 0.00994219
R42961 VDD.n6246 VDD.n6245 0.00994219
R42962 VDD.n6245 VDD.n6228 0.00994219
R42963 VDD.n6243 VDD.n6228 0.00994219
R42964 VDD.n6242 VDD.n6229 0.00994219
R42965 VDD.n6240 VDD.n6229 0.00994219
R42966 VDD.n6240 VDD.n6239 0.00994219
R42967 VDD.n6239 VDD.n6238 0.00994219
R42968 VDD.n6238 VDD.n6232 0.00994219
R42969 VDD.n6235 VDD.n6232 0.00994219
R42970 VDD.n6235 VDD.n6234 0.00994219
R42971 VDD.n6234 VDD.n5265 0.00994219
R42972 VDD.n6684 VDD.n6642 0.00994219
R42973 VDD.n6682 VDD.n6642 0.00994219
R42974 VDD.n6682 VDD.n6681 0.00994219
R42975 VDD.n6681 VDD.n6680 0.00994219
R42976 VDD.n6680 VDD.n6645 0.00994219
R42977 VDD.n6677 VDD.n6645 0.00994219
R42978 VDD.n6677 VDD.n6676 0.00994219
R42979 VDD.n6676 VDD.n6675 0.00994219
R42980 VDD.n6674 VDD.n6647 0.00994219
R42981 VDD.n6672 VDD.n6647 0.00994219
R42982 VDD.n6669 VDD.n6648 0.00994219
R42983 VDD.n6669 VDD.n6649 0.00994219
R42984 VDD.n6667 VDD.n6649 0.00994219
R42985 VDD.n6666 VDD.n6650 0.00994219
R42986 VDD.n6664 VDD.n6650 0.00994219
R42987 VDD.n6664 VDD.n6663 0.00994219
R42988 VDD.n6663 VDD.n6662 0.00994219
R42989 VDD.n6662 VDD.n6653 0.00994219
R42990 VDD.n6659 VDD.n6653 0.00994219
R42991 VDD.n6659 VDD.n6658 0.00994219
R42992 VDD.n6658 VDD.n6657 0.00994219
R42993 VDD.n6656 VDD.n6655 0.00994219
R42994 VDD.n6655 VDD.n2342 0.00994219
R42995 VDD.n7049 VDD.n2340 0.00994219
R42996 VDD.n7050 VDD.n2340 0.00994219
R42997 VDD.n7051 VDD.n2339 0.00994219
R42998 VDD.n7053 VDD.n2339 0.00994219
R42999 VDD.n7053 VDD.n2338 0.00994219
R43000 VDD.n7056 VDD.n2338 0.00994219
R43001 VDD.n7056 VDD.n2337 0.00994219
R43002 VDD.n7059 VDD.n2337 0.00994219
R43003 VDD.n7059 VDD.n2336 0.00994219
R43004 VDD.n7061 VDD.n2336 0.00994219
R43005 VDD.n7064 VDD.n7063 0.00994219
R43006 VDD.n7063 VDD.n2333 0.00994219
R43007 VDD.n7083 VDD.n7082 0.00994219
R43008 VDD.n7082 VDD.n2335 0.00994219
R43009 VDD.n7080 VDD.n2335 0.00994219
R43010 VDD.n7079 VDD.n7066 0.00994219
R43011 VDD.n7077 VDD.n7066 0.00994219
R43012 VDD.n7077 VDD.n7076 0.00994219
R43013 VDD.n7076 VDD.n7075 0.00994219
R43014 VDD.n7075 VDD.n7069 0.00994219
R43015 VDD.n7072 VDD.n7069 0.00994219
R43016 VDD.n7072 VDD.n7071 0.00994219
R43017 VDD.n7071 VDD.n2265 0.00994219
R43018 VDD.n10772 VDD.n10771 0.00983484
R43019 VDD.n2049 VDD.n2048 0.00983484
R43020 VDD.n10803 VDD.n10802 0.00983484
R43021 VDD.n10810 VDD.n1987 0.00983484
R43022 VDD.n1967 VDD.n1966 0.00983484
R43023 VDD.n10861 VDD.n10860 0.00983484
R43024 VDD.n10868 VDD.n1922 0.00983484
R43025 VDD.n5523 VDD.n5522 0.00983484
R43026 VDD.n10916 VDD.n10915 0.00983484
R43027 VDD.n10923 VDD.n1895 0.00983484
R43028 VDD.n1875 VDD.n1874 0.00983484
R43029 VDD.n10971 VDD.n10970 0.00983484
R43030 VDD.n10978 VDD.n1830 0.00983484
R43031 VDD.n1819 VDD.n1818 0.00983484
R43032 VDD.n11026 VDD.n11025 0.00983484
R43033 VDD.n9156 VDD.n9155 0.00983484
R43034 VDD.n9032 VDD.n9031 0.00983484
R43035 VDD.n9016 VDD.n9015 0.00983484
R43036 VDD.n8935 VDD.n8934 0.00983484
R43037 VDD.n8885 VDD.n8884 0.00983484
R43038 VDD.n8804 VDD.n8803 0.00983484
R43039 VDD.n8759 VDD.n8758 0.00983484
R43040 VDD.n9144 VDD.n9143 0.00983484
R43041 VDD.n8742 VDD.n8741 0.00983484
R43042 VDD.n8721 VDD.n8720 0.00983484
R43043 VDD.n8709 VDD.n8708 0.00983484
R43044 VDD.n8683 VDD.n8682 0.00983484
R43045 VDD.n8671 VDD.n8670 0.00983484
R43046 VDD.n8650 VDD.n8649 0.00983484
R43047 VDD.n12615 VDD.n12 0.00983484
R43048 VDD.n8130 VDD.n8128 0.00983194
R43049 VDD.n8127 VDD.n8125 0.00983194
R43050 VDD.n8124 VDD.n2020 0.00983194
R43051 VDD.n2027 VDD.n2023 0.00983194
R43052 VDD.n2031 VDD.n2028 0.00983194
R43053 VDD.n2035 VDD.n2032 0.00983194
R43054 VDD.n2101 VDD.n2099 0.00983194
R43055 VDD.n2098 VDD.n2096 0.00983194
R43056 VDD.n2095 VDD.n2010 0.00983194
R43057 VDD.n10788 VDD.n10787 0.00983194
R43058 VDD.n10792 VDD.n10789 0.00983194
R43059 VDD.n10796 VDD.n10793 0.00983194
R43060 VDD.n5593 VDD.n5591 0.00983194
R43061 VDD.n5590 VDD.n5588 0.00983194
R43062 VDD.n5587 VDD.n1947 0.00983194
R43063 VDD.n1972 VDD.n1950 0.00983194
R43064 VDD.n1976 VDD.n1973 0.00983194
R43065 VDD.n1980 VDD.n1977 0.00983194
R43066 VDD.n5614 VDD.n5612 0.00983194
R43067 VDD.n5611 VDD.n5609 0.00983194
R43068 VDD.n5608 VDD.n1937 0.00983194
R43069 VDD.n10846 VDD.n10845 0.00983194
R43070 VDD.n10850 VDD.n10847 0.00983194
R43071 VDD.n10854 VDD.n10851 0.00983194
R43072 VDD.n5899 VDD.n5897 0.00983194
R43073 VDD.n5896 VDD.n5894 0.00983194
R43074 VDD.n5893 VDD.n5892 0.00983194
R43075 VDD.n5494 VDD.n5493 0.00983194
R43076 VDD.n5498 VDD.n5495 0.00983194
R43077 VDD.n5502 VDD.n5499 0.00983194
R43078 VDD.n5677 VDD.n5675 0.00983194
R43079 VDD.n5674 VDD.n5672 0.00983194
R43080 VDD.n5671 VDD.n1910 0.00983194
R43081 VDD.n10901 VDD.n10900 0.00983194
R43082 VDD.n10905 VDD.n10902 0.00983194
R43083 VDD.n10909 VDD.n10906 0.00983194
R43084 VDD.n5690 VDD.n5688 0.00983194
R43085 VDD.n5687 VDD.n5685 0.00983194
R43086 VDD.n5684 VDD.n1855 0.00983194
R43087 VDD.n1880 VDD.n1858 0.00983194
R43088 VDD.n1884 VDD.n1881 0.00983194
R43089 VDD.n1888 VDD.n1885 0.00983194
R43090 VDD.n5797 VDD.n5795 0.00983194
R43091 VDD.n5794 VDD.n5792 0.00983194
R43092 VDD.n5791 VDD.n1845 0.00983194
R43093 VDD.n10956 VDD.n10955 0.00983194
R43094 VDD.n10960 VDD.n10957 0.00983194
R43095 VDD.n10964 VDD.n10961 0.00983194
R43096 VDD.n5742 VDD.n5740 0.00983194
R43097 VDD.n5739 VDD.n5737 0.00983194
R43098 VDD.n5736 VDD.n1790 0.00983194
R43099 VDD.n1797 VDD.n1793 0.00983194
R43100 VDD.n1801 VDD.n1798 0.00983194
R43101 VDD.n1805 VDD.n1802 0.00983194
R43102 VDD.n5716 VDD.n5714 0.00983194
R43103 VDD.n5713 VDD.n5711 0.00983194
R43104 VDD.n5710 VDD.n1783 0.00983194
R43105 VDD.n11011 VDD.n11010 0.00983194
R43106 VDD.n11015 VDD.n11012 0.00983194
R43107 VDD.n11019 VDD.n11016 0.00983194
R43108 VDD.n9062 VDD.n9060 0.00983194
R43109 VDD.n9059 VDD.n9057 0.00983194
R43110 VDD.n9056 VDD.n9055 0.00983194
R43111 VDD.n9052 VDD.n9050 0.00983194
R43112 VDD.n9049 VDD.n9048 0.00983194
R43113 VDD.n9046 VDD.n9045 0.00983194
R43114 VDD.n8928 VDD.n8926 0.00983194
R43115 VDD.n8925 VDD.n8923 0.00983194
R43116 VDD.n8922 VDD.n8921 0.00983194
R43117 VDD.n8918 VDD.n8916 0.00983194
R43118 VDD.n8915 VDD.n8914 0.00983194
R43119 VDD.n8912 VDD.n8505 0.00983194
R43120 VDD.n8849 VDD.n8516 0.00983194
R43121 VDD.n8853 VDD.n8852 0.00983194
R43122 VDD.n8857 VDD.n8854 0.00983194
R43123 VDD.n8862 VDD.n8861 0.00983194
R43124 VDD.n8866 VDD.n8863 0.00983194
R43125 VDD.n8870 VDD.n8867 0.00983194
R43126 VDD.n8579 VDD.n8577 0.00983194
R43127 VDD.n8576 VDD.n8574 0.00983194
R43128 VDD.n8573 VDD.n8572 0.00983194
R43129 VDD.n8569 VDD.n8567 0.00983194
R43130 VDD.n8566 VDD.n8565 0.00983194
R43131 VDD.n8563 VDD.n8562 0.00983194
R43132 VDD.n9083 VDD.n9081 0.00983194
R43133 VDD.n9080 VDD.n9078 0.00983194
R43134 VDD.n9077 VDD.n8465 0.00983194
R43135 VDD.n9176 VDD.n9174 0.00983194
R43136 VDD.n9173 VDD.n9172 0.00983194
R43137 VDD.n9170 VDD.n9169 0.00983194
R43138 VDD.n8591 VDD.n8589 0.00983194
R43139 VDD.n8588 VDD.n8586 0.00983194
R43140 VDD.n8585 VDD.n180 0.00983194
R43141 VDD.n12458 VDD.n12456 0.00983194
R43142 VDD.n12455 VDD.n12454 0.00983194
R43143 VDD.n12452 VDD.n12451 0.00983194
R43144 VDD.n8604 VDD.n8602 0.00983194
R43145 VDD.n8601 VDD.n8599 0.00983194
R43146 VDD.n8598 VDD.n109 0.00983194
R43147 VDD.n12478 VDD.n12477 0.00983194
R43148 VDD.n12482 VDD.n12479 0.00983194
R43149 VDD.n12486 VDD.n12483 0.00983194
R43150 VDD.n8696 VDD.n8694 0.00983194
R43151 VDD.n8693 VDD.n8691 0.00983194
R43152 VDD.n8690 VDD.n100 0.00983194
R43153 VDD.n12514 VDD.n12512 0.00983194
R43154 VDD.n12511 VDD.n12510 0.00983194
R43155 VDD.n12508 VDD.n12507 0.00983194
R43156 VDD.n8663 VDD.n8661 0.00983194
R43157 VDD.n8660 VDD.n8658 0.00983194
R43158 VDD.n8657 VDD.n29 0.00983194
R43159 VDD.n12534 VDD.n12533 0.00983194
R43160 VDD.n12538 VDD.n12535 0.00983194
R43161 VDD.n12542 VDD.n12539 0.00983194
R43162 VDD.n8632 VDD.n8630 0.00983194
R43163 VDD.n8629 VDD.n8627 0.00983194
R43164 VDD.n8626 VDD.n20 0.00983194
R43165 VDD.n12608 VDD.n12606 0.00983194
R43166 VDD.n12605 VDD.n12604 0.00983194
R43167 VDD.n12602 VDD.n12601 0.00983194
R43168 VDD.n2115 VDD.n2113 0.00974509
R43169 VDD.n2112 VDD.n1993 0.00974509
R43170 VDD.n10827 VDD.n10825 0.00974509
R43171 VDD.n10824 VDD.n10823 0.00974509
R43172 VDD.n5635 VDD.n5633 0.00974509
R43173 VDD.n5632 VDD.n5630 0.00974509
R43174 VDD.n5629 VDD.n1928 0.00974509
R43175 VDD.n10882 VDD.n10880 0.00974509
R43176 VDD.n10879 VDD.n10878 0.00974509
R43177 VDD.n10876 VDD.n10875 0.00974509
R43178 VDD.n5852 VDD.n5850 0.00974509
R43179 VDD.n5849 VDD.n5847 0.00974509
R43180 VDD.n5846 VDD.n1901 0.00974509
R43181 VDD.n10937 VDD.n10935 0.00974509
R43182 VDD.n10934 VDD.n10933 0.00974509
R43183 VDD.n10931 VDD.n10930 0.00974509
R43184 VDD.n5703 VDD.n5701 0.00974509
R43185 VDD.n5700 VDD.n5698 0.00974509
R43186 VDD.n5697 VDD.n1836 0.00974509
R43187 VDD.n10992 VDD.n10990 0.00974509
R43188 VDD.n10989 VDD.n10988 0.00974509
R43189 VDD.n10986 VDD.n10985 0.00974509
R43190 VDD.n8976 VDD.n8497 0.00974509
R43191 VDD.n8980 VDD.n8979 0.00974509
R43192 VDD.n8984 VDD.n8981 0.00974509
R43193 VDD.n8989 VDD.n8988 0.00974509
R43194 VDD.n8993 VDD.n8990 0.00974509
R43195 VDD.n8997 VDD.n8994 0.00974509
R43196 VDD.n8797 VDD.n8795 0.00974509
R43197 VDD.n8794 VDD.n8792 0.00974509
R43198 VDD.n8791 VDD.n8790 0.00974509
R43199 VDD.n8787 VDD.n8785 0.00974509
R43200 VDD.n8784 VDD.n8783 0.00974509
R43201 VDD.n8781 VDD.n8524 0.00974509
R43202 VDD.n8734 VDD.n8732 0.00974509
R43203 VDD.n8731 VDD.n8729 0.00974509
R43204 VDD.n8728 VDD.n119 0.00974509
R43205 VDD.n126 VDD.n122 0.00974509
R43206 VDD.n130 VDD.n127 0.00974509
R43207 VDD.n134 VDD.n131 0.00974509
R43208 VDD.n8618 VDD.n8616 0.00974509
R43209 VDD.n8615 VDD.n8613 0.00974509
R43210 VDD.n8612 VDD.n39 0.00974509
R43211 VDD.n80 VDD.n42 0.00974509
R43212 VDD.n84 VDD.n81 0.00974509
R43213 VDD.n88 VDD.n85 0.00974509
R43214 VDD.n6712 VDD.n6711 0.00970384
R43215 VDD.n6710 VDD.n6709 0.00970384
R43216 VDD.n6708 VDD.n6707 0.00970384
R43217 VDD.n6705 VDD.n6704 0.00970384
R43218 VDD.n6703 VDD.n6702 0.00970384
R43219 VDD.n6701 VDD.n6700 0.00970384
R43220 VDD.n6698 VDD.n6697 0.00970384
R43221 VDD.n6696 VDD.n6695 0.00970384
R43222 VDD.n6694 VDD.n6693 0.00970384
R43223 VDD.n6691 VDD.n6690 0.00970384
R43224 VDD.n6689 VDD.n6688 0.00970384
R43225 VDD.n6687 VDD.n6686 0.00970384
R43226 VDD.n6641 VDD.n6640 0.00970384
R43227 VDD.n6639 VDD.n6638 0.00970384
R43228 VDD.n6637 VDD.n6636 0.00970384
R43229 VDD.n5434 VDD.n5267 0.00970384
R43230 VDD.n5436 VDD.n5435 0.00970384
R43231 VDD.n5438 VDD.n5437 0.00970384
R43232 VDD.n5443 VDD.n5442 0.00970384
R43233 VDD.n5441 VDD.n5440 0.00970384
R43234 VDD.n5439 VDD.n5269 0.00970384
R43235 VDD.n6630 VDD.n6629 0.00970384
R43236 VDD.n6628 VDD.n6627 0.00970384
R43237 VDD.n6626 VDD.n6625 0.00970384
R43238 VDD.n950 VDD.n949 0.00969752
R43239 VDD.n970 VDD.n969 0.00964201
R43240 VDD.n972 VDD.n971 0.00964201
R43241 VDD.n974 VDD.n973 0.00964201
R43242 VDD.n976 VDD.n975 0.00964201
R43243 VDD.n988 VDD.n987 0.00964201
R43244 VDD.n990 VDD.n989 0.00964201
R43245 VDD.n992 VDD.n991 0.00964201
R43246 VDD.n994 VDD.n993 0.00964201
R43247 VDD.n1009 VDD.n1008 0.00964201
R43248 VDD.n1011 VDD.n1010 0.00964201
R43249 VDD.n1013 VDD.n1012 0.00964201
R43250 VDD.n1015 VDD.n1014 0.00964201
R43251 VDD.n1030 VDD.n1029 0.00964201
R43252 VDD.n1028 VDD.n1027 0.00964201
R43253 VDD.n1026 VDD.n1025 0.00964201
R43254 VDD.n1024 VDD.n1023 0.00964201
R43255 VDD.n1206 VDD.n1189 0.0095
R43256 VDD.n1176 VDD.n1118 0.0095
R43257 VDD.n1336 VDD.n1335 0.0095
R43258 VDD.n1383 VDD.n1382 0.0095
R43259 VDD.n1269 VDD.n1251 0.0095
R43260 VDD.n1236 VDD.n1219 0.0095
R43261 VDD.n1304 VDD.n1303 0.0095
R43262 VDD.n1072 VDD.n896 0.0095
R43263 VDD.n1059 VDD.n1058 0.0095
R43264 VDD.n1163 VDD.n1139 0.0095
R43265 VDD.n6287 VDD.n6286 0.00947673
R43266 VDD.n6279 VDD.n6278 0.00947673
R43267 VDD.n6251 VDD.n6250 0.00947673
R43268 VDD.n6243 VDD.n6242 0.00947673
R43269 VDD.n6675 VDD.n6674 0.00947673
R43270 VDD.n6667 VDD.n6666 0.00947673
R43271 VDD.n7064 VDD.n7061 0.00947673
R43272 VDD.n7080 VDD.n7079 0.00947673
R43273 VDD.n5892 VDD.n5890 0.00945616
R43274 VDD.n8017 VDD.n8016 0.00944828
R43275 VDD.n968 VDD.n682 0.00931657
R43276 VDD.n969 VDD.n968 0.00931657
R43277 VDD.n970 VDD.n967 0.00931657
R43278 VDD.n971 VDD.n967 0.00931657
R43279 VDD.n972 VDD.n966 0.00931657
R43280 VDD.n973 VDD.n966 0.00931657
R43281 VDD.n974 VDD.n965 0.00931657
R43282 VDD.n975 VDD.n965 0.00931657
R43283 VDD.n976 VDD.n964 0.00931657
R43284 VDD.n977 VDD.n964 0.00931657
R43285 VDD.n986 VDD.n963 0.00931657
R43286 VDD.n987 VDD.n963 0.00931657
R43287 VDD.n988 VDD.n962 0.00931657
R43288 VDD.n989 VDD.n962 0.00931657
R43289 VDD.n990 VDD.n961 0.00931657
R43290 VDD.n991 VDD.n961 0.00931657
R43291 VDD.n992 VDD.n960 0.00931657
R43292 VDD.n993 VDD.n960 0.00931657
R43293 VDD.n994 VDD.n959 0.00931657
R43294 VDD.n995 VDD.n959 0.00931657
R43295 VDD.n996 VDD.n958 0.00931657
R43296 VDD.n997 VDD.n958 0.00931657
R43297 VDD.n1005 VDD.n942 0.00931657
R43298 VDD.n1006 VDD.n942 0.00931657
R43299 VDD.n1007 VDD.n941 0.00931657
R43300 VDD.n1008 VDD.n941 0.00931657
R43301 VDD.n1009 VDD.n940 0.00931657
R43302 VDD.n1010 VDD.n940 0.00931657
R43303 VDD.n1011 VDD.n939 0.00931657
R43304 VDD.n1012 VDD.n939 0.00931657
R43305 VDD.n1013 VDD.n938 0.00931657
R43306 VDD.n1014 VDD.n938 0.00931657
R43307 VDD.n1015 VDD.n937 0.00931657
R43308 VDD.n1016 VDD.n937 0.00931657
R43309 VDD.n1031 VDD.n1017 0.00931657
R43310 VDD.n1030 VDD.n1017 0.00931657
R43311 VDD.n1029 VDD.n1018 0.00931657
R43312 VDD.n1028 VDD.n1018 0.00931657
R43313 VDD.n1027 VDD.n1019 0.00931657
R43314 VDD.n1026 VDD.n1019 0.00931657
R43315 VDD.n1025 VDD.n1020 0.00931657
R43316 VDD.n1024 VDD.n1020 0.00931657
R43317 VDD.n1023 VDD.n1021 0.00931657
R43318 VDD.n1022 VDD.n1021 0.00931657
R43319 VDD.n6267 VDD.n6266 0.00927724
R43320 VDD.n6266 VDD.n6262 0.00927724
R43321 VDD.n7048 VDD.n2342 0.00927724
R43322 VDD.n7049 VDD.n7048 0.00927724
R43323 VDD.n6284 VDD.n6283 0.00887828
R43324 VDD.n6248 VDD.n6247 0.00887828
R43325 VDD.n6672 VDD.n2350 0.00887828
R43326 VDD.n7084 VDD.n2333 0.00887828
R43327 VDD.n1450 VDD.n1449 0.00882321
R43328 VDD.n8014 VDD.n8013 0.00877586
R43329 VDD.n1612 VDD.n1610 0.00867241
R43330 VDD.n1480 VDD.n813 0.00867241
R43331 VDD.n5493 VDD.n1919 0.00864196
R43332 VDD.n1418 VDD.n852 0.00841379
R43333 VDD.n1678 VDD.n745 0.00841379
R43334 VDD.n1619 VDD.n1618 0.00841379
R43335 VDD.n1106 VDD.n1100 0.00841379
R43336 VDD.n1684 VDD.n742 0.00841379
R43337 VDD.n1698 VDD.n1697 0.00841379
R43338 VDD.n1045 VDD.n936 0.00841379
R43339 VDD.n1145 VDD.n706 0.00841379
R43340 VDD.n12583 VDD.n12577 0.0083892
R43341 VDD.n1426 VDD.n851 0.00836207
R43342 VDD.n1432 VDD.n1431 0.00836207
R43343 VDD.n1417 VDD.n873 0.00836207
R43344 VDD.n793 VDD.n744 0.00836207
R43345 VDD.n830 VDD.n738 0.00836207
R43346 VDD.n1371 VDD.n739 0.00836207
R43347 VDD.n1257 VDD.n783 0.00836207
R43348 VDD.n1352 VDD.n1085 0.00836207
R43349 VDD.n1467 VDD.n741 0.00836207
R43350 VDD.n885 VDD.n736 0.00836207
R43351 VDD.n1047 VDD.n1046 0.00836207
R43352 VDD.n1722 VDD.n1721 0.00836207
R43353 VDD.n1002 VDD.n997 0.00831065
R43354 VDD.n1637 VDD.n773 0.00808484
R43355 VDD.n1593 VDD.n1592 0.00806656
R43356 VDD.n6300 VDD.n6200 0.00801385
R43357 VDD.n1567 VDD.n1566 0.00800848
R43358 VDD.n697 VDD.n696 0.00797611
R43359 VDD.n7890 VDD.n7889 0.00791176
R43360 VDD.n7909 VDD.n7864 0.00787705
R43361 VDD.n8013 VDD.n8012 0.00763793
R43362 VDD.n1636 VDD.n774 0.0076267
R43363 VDD.n776 VDD.n775 0.0076267
R43364 VDD.n1635 VDD.n1634 0.0076267
R43365 VDD.n7983 VDD.n7982 0.0073513
R43366 VDD.n2196 VDD.n2195 0.0073513
R43367 VDD.n2191 VDD.n2190 0.0073513
R43368 VDD.n7989 VDD.n2192 0.0073513
R43369 VDD.n7988 VDD.n7987 0.0073513
R43370 VDD.n2221 VDD.n2220 0.0073513
R43371 VDD.n2224 VDD.n2223 0.0073513
R43372 VDD.n2231 VDD.n2212 0.0073513
R43373 VDD.n2214 VDD.n2213 0.0073513
R43374 VDD.n2228 VDD.n2227 0.0073513
R43375 VDD.n1542 VDD.n1535 0.00716667
R43376 VDD.n9134 VDD.n9132 0.00714138
R43377 VDD.n7986 VDD.n2193 0.00713029
R43378 VDD.n2219 VDD.n2218 0.00713029
R43379 VDD.n1529 VDD.n1523 0.00711202
R43380 VDD.n7980 VDD.n2197 0.0070075
R43381 VDD.n7979 VDD.n2194 0.0070075
R43382 VDD.n2217 VDD.n2216 0.0070075
R43383 VDD.n2215 VDD.n2207 0.0070075
R43384 VDD.n2038 VDD.n2007 0.0069938
R43385 VDD.n1956 VDD.n1934 0.0069938
R43386 VDD.n5512 VDD.n1907 0.0069938
R43387 VDD.n1864 VDD.n1842 0.0069938
R43388 VDD.n1808 VDD.n1780 0.0069938
R43389 VDD.n9064 VDD.n8475 0.0069938
R43390 VDD.n8891 VDD.n8513 0.0069938
R43391 VDD.n8748 VDD.n8582 0.0069938
R43392 VDD.n8698 VDD.n8607 0.0069938
R43393 VDD.n8639 VDD.n8623 0.0069938
R43394 VDD.n2160 VDD.n2159 0.00696552
R43395 VDD.n7962 VDD.n7961 0.00693383
R43396 VDD.n7965 VDD.n2202 0.00693383
R43397 VDD.n7968 VDD.n7966 0.00693383
R43398 VDD.n7967 VDD.n2200 0.00693383
R43399 VDD.n7970 VDD.n7969 0.00693383
R43400 VDD.n1206 VDD.n1205 0.00691379
R43401 VDD.n1176 VDD.n1134 0.00691379
R43402 VDD.n1336 VDD.n1319 0.00691379
R43403 VDD.n1383 VDD.n1365 0.00691379
R43404 VDD.n1269 VDD.n1268 0.00691379
R43405 VDD.n1236 VDD.n1235 0.00691379
R43406 VDD.n1304 VDD.n1287 0.00691379
R43407 VDD.n1072 VDD.n879 0.00691379
R43408 VDD.n1059 VDD.n917 0.00691379
R43409 VDD.n1163 VDD.n1156 0.00691379
R43410 VDD.n7175 VDD.n2297 0.00682401
R43411 VDD.n7827 VDD.n2240 0.00682401
R43412 VDD.n10821 VDD.n10820 0.00664271
R43413 VDD.n2043 VDD.n2038 0.00658794
R43414 VDD.n1961 VDD.n1956 0.00658794
R43415 VDD.n5517 VDD.n5512 0.00658794
R43416 VDD.n1869 VDD.n1864 0.00658794
R43417 VDD.n1813 VDD.n1808 0.00658794
R43418 VDD.n9069 VDD.n8475 0.00658794
R43419 VDD.n8896 VDD.n8513 0.00658794
R43420 VDD.n8753 VDD.n8582 0.00658794
R43421 VDD.n8703 VDD.n8607 0.00658794
R43422 VDD.n8644 VDD.n8623 0.00658794
R43423 VDD.n2233 VDD.n2211 0.00656548
R43424 VDD.n7993 VDD.n2189 0.00651637
R43425 VDD.n8017 VDD.n2165 0.0065
R43426 VDD.n2201 VDD.n2199 0.0064427
R43427 VDD.n10760 VDD.n10759 0.00633837
R43428 VDD.n1633 VDD.n777 0.00625226
R43429 VDD.n1519 VDD.n778 0.00625226
R43430 VDD.n1632 VDD.n1631 0.00625226
R43431 VDD.n8092 VDD.n2116 0.00617735
R43432 VDD.n12448 VDD.n195 0.00617182
R43433 VDD.n12445 VDD.n195 0.00617182
R43434 VDD.n12626 VDD.n12621 0.00599088
R43435 VDD.n1736 VDD.n696 0.00595628
R43436 VDD.n7975 VDD.n7973 0.00595157
R43437 VDD.n7974 VDD.n2198 0.00595157
R43438 VDD.n7977 VDD.n7976 0.00595157
R43439 VDD.n7850 VDD.n7849 0.00595157
R43440 VDD.n7851 VDD.n2206 0.00595157
R43441 VDD.n12630 VDD.n12625 0.00580154
R43442 VDD.n6320 VDD.n6319 0.00551189
R43443 VDD.n6319 VDD.n5914 0.00551189
R43444 VDD.n6177 VDD.n6016 0.00551189
R43445 VDD.n6179 VDD.n6016 0.00551189
R43446 VDD.n6174 VDD.n6173 0.00550912
R43447 VDD.n2159 VDD.n2158 0.00531034
R43448 VDD.n5768 VDD.n5763 0.00523684
R43449 VDD.n5759 VDD.n5758 0.00523684
R43450 VDD.n5835 VDD.n5830 0.00523684
R43451 VDD.n5826 VDD.n5825 0.00523684
R43452 VDD.n5652 VDD.n5647 0.00523684
R43453 VDD.n5643 VDD.n5642 0.00523684
R43454 VDD.n5570 VDD.n5565 0.00523684
R43455 VDD.n5561 VDD.n5560 0.00523684
R43456 VDD.n8156 VDD.n8151 0.00523684
R43457 VDD.n8147 VDD.n8146 0.00523684
R43458 VDD.n7997 VDD.n2186 0.00512451
R43459 VDD.n1442 VDD.n823 0.00510675
R43460 VDD.n1440 VDD.n823 0.00506157
R43461 VDD.n1756 VDD.n1752 0.00505621
R43462 VDD.n984 VDD.n977 0.00502663
R43463 VDD.n1033 VDD.n1016 0.00502663
R43464 VDD.n5980 VDD.n5979 0.00501642
R43465 VDD.n7305 VDD.n7302 0.00500851
R43466 VDD.n7305 VDD.n7304 0.00500851
R43467 VDD.n7304 VDD.n2088 0.00500851
R43468 VDD.n8168 VDD.n2086 0.00500851
R43469 VDD.n8172 VDD.n2086 0.00500851
R43470 VDD.n8175 VDD.n8174 0.00500851
R43471 VDD.n8175 VDD.n2084 0.00500851
R43472 VDD.n8179 VDD.n2084 0.00500851
R43473 VDD.n8180 VDD.n8179 0.00500851
R43474 VDD.n8183 VDD.n8180 0.00500851
R43475 VDD.n8187 VDD.n2082 0.00500851
R43476 VDD.n8190 VDD.n8189 0.00500851
R43477 VDD.n8190 VDD.n2080 0.00500851
R43478 VDD.n8194 VDD.n2080 0.00500851
R43479 VDD.n8195 VDD.n8194 0.00500851
R43480 VDD.n8196 VDD.n8195 0.00500851
R43481 VDD.n8200 VDD.n8199 0.00500851
R43482 VDD.n8203 VDD.n8200 0.00500851
R43483 VDD.n8207 VDD.n2076 0.00500851
R43484 VDD.n8208 VDD.n8207 0.00500851
R43485 VDD.n8209 VDD.n8208 0.00500851
R43486 VDD.n8213 VDD.n8212 0.00500851
R43487 VDD.n8216 VDD.n8213 0.00500851
R43488 VDD.n8220 VDD.n2072 0.00500851
R43489 VDD.n8221 VDD.n8220 0.00500851
R43490 VDD.n8223 VDD.n2070 0.00500851
R43491 VDD.n8227 VDD.n2070 0.00500851
R43492 VDD.n8228 VDD.n8227 0.00500851
R43493 VDD.n8230 VDD.n8228 0.00500851
R43494 VDD.n8234 VDD.n2068 0.00500851
R43495 VDD.n8235 VDD.n8234 0.00500851
R43496 VDD.n8238 VDD.n2066 0.00500851
R43497 VDD.n8242 VDD.n2066 0.00500851
R43498 VDD.n8243 VDD.n8242 0.00500851
R43499 VDD.n8244 VDD.n8243 0.00500851
R43500 VDD.n8248 VDD.n8247 0.00500851
R43501 VDD.n8251 VDD.n8248 0.00500851
R43502 VDD.n10765 VDD.n2062 0.00500851
R43503 VDD.n10761 VDD.n2062 0.00500851
R43504 VDD.n10761 VDD.n10760 0.00500851
R43505 VDD.n986 VDD.n985 0.00499704
R43506 VDD.n1032 VDD.n1031 0.00499704
R43507 VDD.n1564 VDD.n1510 0.00497964
R43508 VDD.n7960 VDD.n2203 0.00489563
R43509 VDD.n1630 VDD.n779 0.00487783
R43510 VDD.n781 VDD.n780 0.00487783
R43511 VDD.n1629 VDD.n1628 0.00487783
R43512 VDD.n1592 VDD.n1504 0.00487179
R43513 VDD.n2157 VDD.n2156 0.00484483
R43514 VDD.n8141 VDD.n8140 0.00483155
R43515 VDD.n5554 VDD.n5553 0.00483155
R43516 VDD.n5545 VDD.n5544 0.00483155
R43517 VDD.n5820 VDD.n5819 0.00483155
R43518 VDD.n5753 VDD.n5752 0.00483155
R43519 VDD.n8970 VDD.n8953 0.00483155
R43520 VDD.n8830 VDD.n8812 0.00483155
R43521 VDD.n9117 VDD.n9099 0.00483155
R43522 VDD.n162 VDD.n144 0.00483155
R43523 VDD.n73 VDD.n55 0.00483155
R43524 VDD.n8244 VDD.n2064 0.00479584
R43525 VDD.n8212 VDD.n2074 0.00475331
R43526 VDD.n8182 VDD.n2082 0.00462571
R43527 VDD.n8202 VDD.n2076 0.00462571
R43528 VDD.n8188 VDD.n8187 0.00454064
R43529 VDD.n770 VDD.n769 0.00452149
R43530 VDD.n12640 VDD.n12639 0.00449408
R43531 VDD.n12581 VDD.n12558 0.00447616
R43532 VDD.n12582 VDD.n12581 0.00446857
R43533 VDD.n12583 VDD.n12582 0.00446857
R43534 VDD VDD.n0 0.0044645
R43535 VDD.n8223 VDD.n8222 0.00445558
R43536 VDD.n6323 VDD.n5980 0.00444161
R43537 VDD.n5288 VDD.n5287 0.00441304
R43538 VDD.n6413 VDD.n5298 0.00441304
R43539 VDD.n6876 VDD.n2385 0.00441304
R43540 VDD.n2375 VDD.n2374 0.00441304
R43541 VDD.n1628 VDD.n1627 0.00436878
R43542 VDD.n1639 VDD.n1638 0.00434333
R43543 VDD.n773 VDD.n772 0.00434333
R43544 VDD.n1626 VDD.n782 0.00431787
R43545 VDD.n6575 VDD.n6574 0.00429447
R43546 VDD.n6399 VDD.n6398 0.00429447
R43547 VDD.n6862 VDD.n6861 0.00429447
R43548 VDD.n7038 VDD.n7037 0.00429447
R43549 VDD.n1638 VDD.n772 0.00424152
R43550 VDD.n6580 VDD.n6579 0.00418286
R43551 VDD.n5965 VDD.n5964 0.00418286
R43552 VDD.n6610 VDD.n6609 0.00418286
R43553 VDD.n12639 VDD.n0 0.00416864
R43554 VDD.n1641 VDD.n770 0.00406335
R43555 VDD.n60 VDD.n59 0.00405263
R43556 VDD.n69 VDD.n68 0.00405263
R43557 VDD.n149 VDD.n148 0.00405263
R43558 VDD.n158 VDD.n157 0.00405263
R43559 VDD.n9104 VDD.n9103 0.00405263
R43560 VDD.n9113 VDD.n9112 0.00405263
R43561 VDD.n8817 VDD.n8816 0.00405263
R43562 VDD.n8826 VDD.n8825 0.00405263
R43563 VDD.n8957 VDD.n8956 0.00405263
R43564 VDD.n8966 VDD.n8965 0.00405263
R43565 VDD.n6175 VDD.n6174 0.00403102
R43566 VDD.n10766 VDD.n2061 0.00403025
R43567 VDD.n1631 VDD.n1630 0.00398699
R43568 VDD.n8251 VDD.n8250 0.00394518
R43569 VDD.n2054 VDD.n2035 0.00388205
R43570 VDD.n10797 VDD.n10796 0.00388205
R43571 VDD.n1981 VDD.n1980 0.00388205
R43572 VDD.n10855 VDD.n10854 0.00388205
R43573 VDD.n10910 VDD.n10909 0.00388205
R43574 VDD.n1889 VDD.n1888 0.00388205
R43575 VDD.n10965 VDD.n10964 0.00388205
R43576 VDD.n1824 VDD.n1805 0.00388205
R43577 VDD.n11020 VDD.n11019 0.00388205
R43578 VDD.n9063 VDD.n9062 0.00385073
R43579 VDD.n8929 VDD.n8928 0.00385073
R43580 VDD.n8890 VDD.n8516 0.00385073
R43581 VDD.n8764 VDD.n8579 0.00385073
R43582 VDD.n9150 VDD.n9083 0.00385073
R43583 VDD.n8747 VDD.n8591 0.00385073
R43584 VDD.n8714 VDD.n8604 0.00385073
R43585 VDD.n8697 VDD.n8696 0.00385073
R43586 VDD.n8664 VDD.n8663 0.00385073
R43587 VDD.n8638 VDD.n8632 0.00385073
R43588 VDD.n10875 VDD.n10873 0.00385057
R43589 VDD.n10930 VDD.n10928 0.00385057
R43590 VDD.n10985 VDD.n10983 0.00385057
R43591 VDD.n9021 VDD.n8497 0.00381954
R43592 VDD.n8798 VDD.n8797 0.00381954
R43593 VDD.n8735 VDD.n8734 0.00381954
R43594 VDD.n8676 VDD.n8618 0.00381954
R43595 VDD.n10148 VDD.n9184 0.00378966
R43596 VDD.n10148 VDD.n9185 0.00378966
R43597 VDD.n8199 VDD.n2078 0.00377505
R43598 VDD.n11136 VDD.n11135 0.00372459
R43599 VDD.n6190 VDD.n5988 0.0037107
R43600 VDD.n6328 VDD.n5487 0.00371011
R43601 VDD.n780 VDD.n779 0.00370701
R43602 VDD.n1629 VDD.n781 0.00370701
R43603 VDD.n949 VDD.n948 0.00364636
R43604 VDD.n8215 VDD.n2072 0.00360491
R43605 VDD.n8238 VDD.n8237 0.00360491
R43606 VDD.n10820 VDD.n2000 0.00360238
R43607 VDD.n1640 VDD.n1639 0.00357975
R43608 VDD.n8064 VDD.n2147 0.00355172
R43609 VDD.n10815 VDD.n2004 0.00354033
R43610 VDD.n1565 VDD.n1564 0.00352885
R43611 VDD.n1449 VDD.n821 0.00352662
R43612 VDD.n7853 VDD.n7852 0.00342224
R43613 VDD.n5950 VDD.n5949 0.00334483
R43614 VDD.n10890 VDD.n1919 0.0031618
R43615 VDD.n7853 VDD.n2205 0.00302933
R43616 VDD.n8174 VDD.n8173 0.00300945
R43617 VDD.n12586 VDD.n12558 0.00289832
R43618 VDD.n8012 VDD.n8011 0.00277586
R43619 VDD.n8230 VDD.n8229 0.00275425
R43620 VDD.n8229 VDD.n2068 0.00275425
R43621 VDD.n680 VDD.n679 0.00274852
R43622 VDD.n5362 VDD.n5299 0.00272414
R43623 VDD.n2402 VDD.n2401 0.00272414
R43624 VDD.n5902 VDD.n5541 0.00272168
R43625 VDD.n5905 VDD.n5901 0.00272168
R43626 VDD.n5889 VDD.n1918 0.00272168
R43627 VDD.n5534 VDD.n5490 0.00272168
R43628 VDD.n5907 VDD.n5541 0.00272168
R43629 VDD.n5905 VDD.n5902 0.00272168
R43630 VDD.n5529 VDD.n5490 0.00272168
R43631 VDD.n5890 VDD.n5889 0.00272168
R43632 VDD.n8092 VDD.n2108 0.00270566
R43633 VDD.n8095 VDD.n2108 0.00270566
R43634 VDD.n1447 VDD.n821 0.00268589
R43635 VDD.n8068 VDD.n8067 0.00267241
R43636 VDD.n5529 VDD.n5528 0.00266075
R43637 VDD.n5220 VDD.n2411 0.00263633
R43638 VDD.n5218 VDD.n2411 0.00263633
R43639 VDD.n1548 VDD.n1547 0.00263115
R43640 VDD.n1756 VDD.n681 0.00262663
R43641 VDD.n998 VDD.n956 0.00262663
R43642 VDD.n12640 VDD.n2 0.00262663
R43643 VDD.n681 VDD.n678 0.00262663
R43644 VDD.n1002 VDD.n998 0.00262663
R43645 VDD.n12642 VDD.n2 0.00262663
R43646 VDD.n1634 VDD.n1633 0.00261256
R43647 VDD.n5503 VDD.n5502 0.00259812
R43648 VDD.n8098 VDD.n2105 0.00257859
R43649 VDD.n6300 VDD.n6299 0.00254425
R43650 VDD.n7963 VDD.n7960 0.0025382
R43651 VDD.n8173 VDD.n8172 0.00249905
R43652 VDD.n5249 VDD.n5248 0.00237378
R43653 VDD.n5459 VDD.n5458 0.00237378
R43654 VDD.n5348 VDD.n5347 0.00237378
R43655 VDD.n6394 VDD.n6393 0.00237378
R43656 VDD.n5481 VDD.n5479 0.00237378
R43657 VDD.n2305 VDD.n2303 0.00237378
R43658 VDD.n5420 VDD.n5419 0.00237378
R43659 VDD.n7110 VDD.n7109 0.00237378
R43660 VDD.n956 VDD.n952 0.00236391
R43661 VDD.n8011 VDD.n2121 0.00236207
R43662 VDD.n7820 VDD.n2243 0.00235027
R43663 VDD.n7816 VDD.n2243 0.00235027
R43664 VDD.n7816 VDD.n7815 0.00235027
R43665 VDD.n7815 VDD.n7814 0.00235027
R43666 VDD.n7814 VDD.n2246 0.00235027
R43667 VDD.n7810 VDD.n2246 0.00235027
R43668 VDD.n7808 VDD.n7807 0.00235027
R43669 VDD.n7807 VDD.n2248 0.00235027
R43670 VDD.n7803 VDD.n2248 0.00235027
R43671 VDD.n7803 VDD.n7802 0.00235027
R43672 VDD.n7802 VDD.n7801 0.00235027
R43673 VDD.n7798 VDD.n7797 0.00235027
R43674 VDD.n7797 VDD.n7796 0.00235027
R43675 VDD.n7793 VDD.n7792 0.00235027
R43676 VDD.n7792 VDD.n7791 0.00235027
R43677 VDD.n7791 VDD.n2254 0.00235027
R43678 VDD.n7787 VDD.n2254 0.00235027
R43679 VDD.n7787 VDD.n7786 0.00235027
R43680 VDD.n7786 VDD.n7785 0.00235027
R43681 VDD.n7785 VDD.n2256 0.00235027
R43682 VDD.n7781 VDD.n2256 0.00235027
R43683 VDD.n7779 VDD.n7778 0.00235027
R43684 VDD.n7778 VDD.n2258 0.00235027
R43685 VDD.n7774 VDD.n7773 0.00235027
R43686 VDD.n7773 VDD.n7772 0.00235027
R43687 VDD.n7772 VDD.n2261 0.00235027
R43688 VDD.n7768 VDD.n2261 0.00235027
R43689 VDD.n7768 VDD.n7767 0.00235027
R43690 VDD.n7767 VDD.n7766 0.00235027
R43691 VDD.n7766 VDD.n2263 0.00235027
R43692 VDD.n7762 VDD.n2263 0.00235027
R43693 VDD.n7762 VDD.n7761 0.00235027
R43694 VDD.n7759 VDD.n2266 0.00235027
R43695 VDD.n7755 VDD.n2266 0.00235027
R43696 VDD.n7755 VDD.n7754 0.00235027
R43697 VDD.n7754 VDD.n7753 0.00235027
R43698 VDD.n7753 VDD.n2268 0.00235027
R43699 VDD.n7749 VDD.n2268 0.00235027
R43700 VDD.n7749 VDD.n7748 0.00235027
R43701 VDD.n7748 VDD.n7747 0.00235027
R43702 VDD.n7744 VDD.n7743 0.00235027
R43703 VDD.n7743 VDD.n7742 0.00235027
R43704 VDD.n7739 VDD.n7738 0.00235027
R43705 VDD.n7738 VDD.n7737 0.00235027
R43706 VDD.n7737 VDD.n2274 0.00235027
R43707 VDD.n7733 VDD.n2274 0.00235027
R43708 VDD.n7733 VDD.n7732 0.00235027
R43709 VDD.n7732 VDD.n7731 0.00235027
R43710 VDD.n7731 VDD.n2276 0.00235027
R43711 VDD.n7727 VDD.n2276 0.00235027
R43712 VDD.n7727 VDD.n7726 0.00235027
R43713 VDD.n7724 VDD.n2278 0.00235027
R43714 VDD.n7720 VDD.n2278 0.00235027
R43715 VDD.n7718 VDD.n7717 0.00235027
R43716 VDD.n7717 VDD.n2280 0.00235027
R43717 VDD.n7713 VDD.n7712 0.00235027
R43718 VDD.n7712 VDD.n7711 0.00235027
R43719 VDD.n7708 VDD.n7707 0.00235027
R43720 VDD.n7707 VDD.n7706 0.00235027
R43721 VDD.n7706 VDD.n2285 0.00235027
R43722 VDD.n7702 VDD.n2285 0.00235027
R43723 VDD.n7702 VDD.n7701 0.00235027
R43724 VDD.n7699 VDD.n2287 0.00235027
R43725 VDD.n7695 VDD.n2287 0.00235027
R43726 VDD.n7695 VDD.n7694 0.00235027
R43727 VDD.n7694 VDD.n7693 0.00235027
R43728 VDD.n7693 VDD.n2289 0.00235027
R43729 VDD.n7689 VDD.n7688 0.00235027
R43730 VDD.n7688 VDD.n7687 0.00235027
R43731 VDD.n7747 VDD.n2270 0.00233282
R43732 VDD.n1632 VDD.n778 0.00233258
R43733 VDD.n7781 VDD.n7780 0.00231536
R43734 VDD.n2969 VDD.n2966 0.00229222
R43735 VDD.n2966 VDD.n1768 0.00229222
R43736 VDD.n11038 VDD.n1768 0.00229222
R43737 VDD.n11050 VDD.n11049 0.00229222
R43738 VDD.n11050 VDD.n667 0.00229222
R43739 VDD.n11054 VDD.n667 0.00229222
R43740 VDD.n11055 VDD.n11054 0.00229222
R43741 VDD.n11058 VDD.n11055 0.00229222
R43742 VDD.n11062 VDD.n665 0.00229222
R43743 VDD.n11065 VDD.n11064 0.00229222
R43744 VDD.n11065 VDD.n663 0.00229222
R43745 VDD.n11069 VDD.n663 0.00229222
R43746 VDD.n11070 VDD.n11069 0.00229222
R43747 VDD.n11071 VDD.n11070 0.00229222
R43748 VDD.n11075 VDD.n11074 0.00229222
R43749 VDD.n11078 VDD.n11075 0.00229222
R43750 VDD.n11082 VDD.n659 0.00229222
R43751 VDD.n11083 VDD.n11082 0.00229222
R43752 VDD.n11084 VDD.n11083 0.00229222
R43753 VDD.n11088 VDD.n11087 0.00229222
R43754 VDD.n11091 VDD.n11088 0.00229222
R43755 VDD.n11095 VDD.n655 0.00229222
R43756 VDD.n11096 VDD.n11095 0.00229222
R43757 VDD.n11098 VDD.n653 0.00229222
R43758 VDD.n11102 VDD.n653 0.00229222
R43759 VDD.n11103 VDD.n11102 0.00229222
R43760 VDD.n11104 VDD.n11103 0.00229222
R43761 VDD.n11108 VDD.n11107 0.00229222
R43762 VDD.n11109 VDD.n11108 0.00229222
R43763 VDD.n11113 VDD.n11112 0.00229222
R43764 VDD.n11114 VDD.n11113 0.00229222
R43765 VDD.n11114 VDD.n646 0.00229222
R43766 VDD.n11118 VDD.n646 0.00229222
R43767 VDD.n11121 VDD.n11120 0.00229222
R43768 VDD.n11131 VDD.n631 0.00229222
R43769 VDD.n11135 VDD.n631 0.00229222
R43770 VDD.n11131 VDD.n11130 0.00225841
R43771 VDD.n11119 VDD.n11118 0.00220768
R43772 VDD.n6625 VDD.n6624 0.0021987
R43773 VDD.n11087 VDD.n657 0.00219078
R43774 VDD.n11121 VDD.n640 0.00219078
R43775 VDD.n12643 VDD.n1 0.00218639
R43776 VDD.n8168 VDD.n8167 0.00215879
R43777 VDD.n7719 VDD.n7718 0.00215826
R43778 VDD.n12625 VDD.n9 0.00214095
R43779 VDD.n11057 VDD.n665 0.00214005
R43780 VDD.n11077 VDD.n659 0.00214005
R43781 VDD.n8167 VDD.n8165 0.00211626
R43782 VDD.n11063 VDD.n11062 0.00210624
R43783 VDD.n7966 VDD.n7965 0.00209618
R43784 VDD.n11098 VDD.n11097 0.00207242
R43785 VDD.n12643 VDD.n12642 0.00206805
R43786 VDD.n7975 VDD.n7974 0.00202251
R43787 VDD.n7977 VDD.n2198 0.00202251
R43788 VDD.n7976 VDD.n2197 0.00202251
R43789 VDD.n7850 VDD.n2207 0.00202251
R43790 VDD.n7849 VDD.n2205 0.00202251
R43791 VDD.n7852 VDD.n7851 0.00202251
R43792 VDD.n7809 VDD.n7808 0.00200116
R43793 VDD.n7742 VDD.n2272 0.00198371
R43794 VDD.n5901 VDD.n5900 0.00197182
R43795 VDD.n2260 VDD.n2258 0.00196625
R43796 VDD.n12630 VDD.n12621 0.00195161
R43797 VDD.n2282 VDD.n2280 0.0019488
R43798 VDD.n7700 VDD.n7699 0.00193134
R43799 VDD.n12579 VDD.n12561 0.00192857
R43800 VDD.n638 VDD.n634 0.00192857
R43801 VDD.n1764 VDD.n1763 0.00192857
R43802 VDD.n6325 VDD.n5913 0.00192857
R43803 VDD.n6015 VDD.n6014 0.00192857
R43804 VDD.n5538 VDD.n5489 0.00192857
R43805 VDD.n5888 VDD.n5886 0.00192857
R43806 VDD.n5911 VDD.n5540 0.00192857
R43807 VDD.n8088 VDD.n2002 0.00192857
R43808 VDD.n8091 VDD.n8090 0.00192857
R43809 VDD.n12632 VDD.n8 0.00192857
R43810 VDD.n12636 VDD.n12635 0.00192857
R43811 VDD.n1001 VDD.n1000 0.00192857
R43812 VDD.n1760 VDD.n677 0.00192857
R43813 VDD.n1751 VDD.n680 0.00192012
R43814 VDD.n8216 VDD.n8215 0.00190359
R43815 VDD.n8237 VDD.n8235 0.00190359
R43816 VDD.n11126 VDD.n644 0.00190334
R43817 VDD.n8068 VDD.n2146 0.00189655
R43818 VDD.n1004 VDD.n952 0.00189053
R43819 VDD.n1183 VDD.n1182 0.00186957
R43820 VDD.n1170 VDD.n1169 0.00186957
R43821 VDD.n1654 VDD.n757 0.00186957
R43822 VDD.n1342 VDD.n1278 0.00186957
R43823 VDD.n1359 VDD.n1358 0.00186957
R43824 VDD.n1389 VDD.n876 0.00186957
R43825 VDD.n1650 VDD.n765 0.00186957
R43826 VDD.n1275 VDD.n1107 0.00186957
R43827 VDD.n1213 VDD.n1212 0.00186957
R43828 VDD.n1066 VDD.n1065 0.00186957
R43829 VDD.n911 VDD.n910 0.00186957
R43830 VDD.n1745 VDD.n1744 0.00186957
R43831 VDD.n11123 VDD.n642 0.00186953
R43832 VDD.n7725 VDD.n7724 0.00180915
R43833 VDD.n2291 VDD.n2289 0.00180915
R43834 VDD.n11074 VDD.n661 0.0018019
R43835 VDD.n5528 VDD.n5503 0.00178392
R43836 VDD.n7801 VDD.n2250 0.00175679
R43837 VDD.n11090 VDD.n655 0.00173427
R43838 VDD.n11112 VDD.n649 0.00173427
R43839 VDD.n8165 VDD.n2088 0.00173346
R43840 VDD.n8196 VDD.n2078 0.00173346
R43841 VDD.n8131 VDD.n8130 0.00168998
R43842 VDD.n8110 VDD.n2101 0.00168998
R43843 VDD.n5594 VDD.n5593 0.00168998
R43844 VDD.n5615 VDD.n5614 0.00168998
R43845 VDD.n5900 VDD.n5899 0.00168998
R43846 VDD.n5865 VDD.n5677 0.00168998
R43847 VDD.n5810 VDD.n5690 0.00168998
R43848 VDD.n5798 VDD.n5797 0.00168998
R43849 VDD.n5743 VDD.n5742 0.00168998
R43850 VDD.n5722 VDD.n5716 0.00168998
R43851 VDD.n9045 VDD.n9043 0.00168998
R43852 VDD.n8946 VDD.n8505 0.00168998
R43853 VDD.n8871 VDD.n8870 0.00168998
R43854 VDD.n8562 VDD.n8560 0.00168998
R43855 VDD.n9169 VDD.n9167 0.00168998
R43856 VDD.n12451 VDD.n12449 0.00168998
R43857 VDD.n12487 VDD.n12486 0.00168998
R43858 VDD.n12507 VDD.n12505 0.00168998
R43859 VDD.n12543 VDD.n12542 0.00168998
R43860 VDD.n12601 VDD.n12599 0.00168998
R43861 VDD.n2164 VDD.n2163 0.00168966
R43862 VDD.n6744 VDD.n6741 0.00168421
R43863 VDD.n6753 VDD.n6751 0.00168421
R43864 VDD.n6756 VDD.n6748 0.00168421
R43865 VDD.n6997 VDD.n6996 0.00168421
R43866 VDD.n6992 VDD.n6991 0.00168421
R43867 VDD.n6987 VDD.n6986 0.00168421
R43868 VDD.n6982 VDD.n6981 0.00168421
R43869 VDD.n6900 VDD.n6899 0.00168421
R43870 VDD.n6895 VDD.n6894 0.00168421
R43871 VDD.n6890 VDD.n6889 0.00168421
R43872 VDD.n6949 VDD.n6948 0.00168421
R43873 VDD.n6944 VDD.n6943 0.00168421
R43874 VDD.n6939 VDD.n6938 0.00168421
R43875 VDD.n6934 VDD.n6933 0.00168421
R43876 VDD.n6919 VDD.n6918 0.00168421
R43877 VDD.n6914 VDD.n6913 0.00168421
R43878 VDD.n6909 VDD.n6908 0.00168421
R43879 VDD.n6524 VDD.n6446 0.00168421
R43880 VDD.n6527 VDD.n6443 0.00168421
R43881 VDD.n6530 VDD.n6440 0.00168421
R43882 VDD.n6533 VDD.n6437 0.00168421
R43883 VDD.n6433 VDD.n6432 0.00168421
R43884 VDD.n6428 VDD.n6427 0.00168421
R43885 VDD.n6423 VDD.n6422 0.00168421
R43886 VDD.n6484 VDD.n6483 0.00168421
R43887 VDD.n6487 VDD.n6480 0.00168421
R43888 VDD.n6490 VDD.n6477 0.00168421
R43889 VDD.n6493 VDD.n6474 0.00168421
R43890 VDD.n6470 VDD.n6469 0.00168421
R43891 VDD.n6465 VDD.n6464 0.00168421
R43892 VDD.n6460 VDD.n6459 0.00168421
R43893 VDD.n6071 VDD.n6068 0.00168421
R43894 VDD.n6065 VDD.n6064 0.00168421
R43895 VDD.n6060 VDD.n6059 0.00168421
R43896 VDD.n6114 VDD.n6111 0.00168421
R43897 VDD.n6108 VDD.n6107 0.00168421
R43898 VDD.n6103 VDD.n6102 0.00168421
R43899 VDD.n7940 VDD.n7939 0.00168421
R43900 VDD.n7935 VDD.n7934 0.00168421
R43901 VDD.n7930 VDD.n7929 0.00168421
R43902 VDD.n7925 VDD.n7924 0.00168421
R43903 VDD.n7921 VDD.n7920 0.00168421
R43904 VDD.n7916 VDD.n7915 0.00168421
R43905 VDD.n7892 VDD.n7885 0.00168421
R43906 VDD.n7895 VDD.n7881 0.00168421
R43907 VDD.n7898 VDD.n7877 0.00168421
R43908 VDD.n7901 VDD.n7874 0.00168421
R43909 VDD.n7904 VDD.n7871 0.00168421
R43910 VDD.n7907 VDD.n7867 0.00168421
R43911 VDD.n8045 VDD.n8044 0.00168421
R43912 VDD.n8040 VDD.n8039 0.00168421
R43913 VDD.n8035 VDD.n8034 0.00168421
R43914 VDD.n8030 VDD.n8029 0.00168421
R43915 VDD.n8026 VDD.n8025 0.00168421
R43916 VDD.n8021 VDD.n8020 0.00168421
R43917 VDD.n6738 VDD.n6735 0.00168421
R43918 VDD.n6802 VDD.n6733 0.00168421
R43919 VDD.n6805 VDD.n6730 0.00168421
R43920 VDD.n6329 VDD.n6328 0.00168023
R43921 VDD.n6008 VDD.n5988 0.00167963
R43922 VDD.n8098 VDD.n8097 0.0016789
R43923 VDD.n5636 VDD.n5635 0.0016789
R43924 VDD.n5853 VDD.n5852 0.0016789
R43925 VDD.n5777 VDD.n5703 0.0016789
R43926 VDD.n8998 VDD.n8997 0.0016789
R43927 VDD.n8837 VDD.n8524 0.0016789
R43928 VDD.n169 VDD.n134 0.0016789
R43929 VDD.n89 VDD.n88 0.0016789
R43930 VDD.n7760 VDD.n7759 0.00161715
R43931 VDD.n7711 VDD.n2283 0.00159969
R43932 VDD.n6283 VDD.n6282 0.00156391
R43933 VDD.n6247 VDD.n6246 0.00156391
R43934 VDD.n6648 VDD.n2350 0.00156391
R43935 VDD.n7084 VDD.n7083 0.00156391
R43936 VDD.n8250 VDD.n2061 0.00156333
R43937 VDD.n2162 VDD.n2161 0.00153448
R43938 VDD.n7973 VDD.n2199 0.00153138
R43939 VDD.n11044 VDD.n673 0.00153137
R43940 VDD.n679 VDD.n678 0.00150592
R43941 VDD.n1520 VDD.n1519 0.00149265
R43942 VDD.n10766 VDD.n10765 0.00147826
R43943 VDD.n11046 VDD.n676 0.00146374
R43944 VDD.n7687 VDD.n2292 0.00146005
R43945 VDD.n7793 VDD.n2252 0.00144259
R43946 VDD.n1641 VDD.n1640 0.00144174
R43947 VDD.n7796 VDD.n2252 0.00140768
R43948 VDD.n11049 VDD.n11048 0.00139611
R43949 VDD.n11104 VDD.n651 0.00139611
R43950 VDD.n11107 VDD.n651 0.00139611
R43951 VDD.n7684 VDD.n2292 0.00139023
R43952 VDD.n6299 VDD.n6298 0.00138218
R43953 VDD.n1520 VDD.n777 0.00133993
R43954 VDD.n7993 VDD.n7992 0.00133493
R43955 VDD.n11046 VDD.n673 0.00132848
R43956 VDD.n676 VDD.n669 0.00129466
R43957 VDD.n2233 VDD.n2232 0.00128581
R43958 VDD.n10890 VDD.n1918 0.00128288
R43959 VDD.n11044 VDD.n11043 0.00126085
R43960 VDD.n7708 VDD.n2283 0.00125058
R43961 VDD.n1637 VDD.n1636 0.00123812
R43962 VDD.n7822 VDD.n7821 0.00123313
R43963 VDD.n7761 VDD.n7760 0.00123313
R43964 VDD.n11043 VDD.n1766 0.0011594
R43965 VDD.n11037 VDD.n1766 0.0011425
R43966 VDD.n7798 VDD.n2250 0.00109348
R43967 VDD.n1601 VDD.n1600 0.00108851
R43968 VDD.n1412 VDD.n1391 0.00108851
R43969 VDD.n820 VDD.n818 0.00108851
R43970 VDD.n810 VDD.n808 0.00108851
R43971 VDD.n1740 VDD.n693 0.00108851
R43972 VDD.n1716 VDD.n713 0.00108851
R43973 VDD.n5979 VDD.n5914 0.00107482
R43974 VDD.n8066 VDD.n8065 0.00106897
R43975 VDD.n12586 VDD.n12585 0.00106802
R43976 VDD.n11091 VDD.n11090 0.00105796
R43977 VDD.n11109 VDD.n649 0.00105796
R43978 VDD.n8222 VDD.n8221 0.00105293
R43979 VDD.n7821 VDD.n7820 0.00104112
R43980 VDD.n7726 VDD.n7725 0.00104112
R43981 VDD.n7689 VDD.n2291 0.00104112
R43982 VDD.n6599 VDD.n2203 0.00104025
R43983 VDD.n7963 VDD.n7962 0.00104025
R43984 VDD.n7961 VDD.n2202 0.00104025
R43985 VDD.n7968 VDD.n7967 0.00104025
R43986 VDD.n7970 VDD.n2200 0.00104025
R43987 VDD.n7969 VDD.n2201 0.00104025
R43988 VDD.n7684 VDD.n7683 0.00102366
R43989 VDD.n6177 VDD.n6175 0.000992701
R43990 VDD.n11038 VDD.n11037 0.000990325
R43991 VDD.n11071 VDD.n661 0.000990325
R43992 VDD.n8189 VDD.n8188 0.000967864
R43993 VDD.n7980 VDD.n7979 0.000966576
R43994 VDD.n2216 VDD.n2215 0.000966576
R43995 VDD.n775 VDD.n774 0.000958145
R43996 VDD.n1635 VDD.n776 0.000958145
R43997 VDD.n1672 VDD.n747 0.000923032
R43998 VDD.n7701 VDD.n7700 0.000918929
R43999 VDD.n7713 VDD.n2282 0.000901474
R44000 VDD.n1558 VDD.n1512 0.000893443
R44001 VDD.n1554 VDD.n1553 0.000893443
R44002 VDD.n11127 VDD.n642 0.000888878
R44003 VDD.n644 VDD.n633 0.000888878
R44004 VDD.n7774 VDD.n2260 0.000884019
R44005 VDD.n8183 VDD.n8182 0.000882798
R44006 VDD.n8203 VDD.n8202 0.000882798
R44007 VDD.n10817 VDD.n10815 0.000872285
R44008 VDD.n7739 VDD.n2272 0.000866563
R44009 VDD.n7810 VDD.n7809 0.000849108
R44010 VDD.n2004 VDD.n2000 0.000810238
R44011 VDD.n2131 VDD.n2130 0.000762697
R44012 VDD.n8209 VDD.n2074 0.000755198
R44013 VDD.n2218 VDD.n2193 0.00072101
R44014 VDD.n11097 VDD.n11096 0.000719801
R44015 VDD.n8247 VDD.n2064 0.000712665
R44016 VDD.n1418 VDD.n1417 0.000706897
R44017 VDD.n1678 VDD.n744 0.000706897
R44018 VDD.n1619 VDD.n783 0.000706897
R44019 VDD.n1352 VDD.n1106 0.000706897
R44020 VDD.n1684 VDD.n741 0.000706897
R44021 VDD.n1697 VDD.n736 0.000706897
R44022 VDD.n1046 VDD.n1045 0.000706897
R44023 VDD.n1721 VDD.n706 0.000706897
R44024 VDD.n7720 VDD.n7719 0.000692009
R44025 VDD.n11064 VDD.n11063 0.000685985
R44026 VDD.n1425 VDD.n844 0.000655172
R44027 VDD.n1691 VDD.n1690 0.000655172
R44028 VDD.n8097 VDD.n8095 0.000655119
R44029 VDD.n11058 VDD.n11057 0.00065217
R44030 VDD.n11078 VDD.n11077 0.00065217
R44031 VDD.n7983 VDD.n2194 0.000622783
R44032 VDD.n7982 VDD.n2196 0.000622783
R44033 VDD.n2195 VDD.n2189 0.000622783
R44034 VDD.n7992 VDD.n2190 0.000622783
R44035 VDD.n2192 VDD.n2191 0.000622783
R44036 VDD.n7989 VDD.n7988 0.000622783
R44037 VDD.n7987 VDD.n7986 0.000622783
R44038 VDD.n2220 VDD.n2219 0.000622783
R44039 VDD.n2223 VDD.n2221 0.000622783
R44040 VDD.n2224 VDD.n2211 0.000622783
R44041 VDD.n2232 VDD.n2231 0.000622783
R44042 VDD.n2213 VDD.n2212 0.000622783
R44043 VDD.n2228 VDD.n2214 0.000622783
R44044 VDD.n2227 VDD.n2217 0.000622783
R44045 VDD.n8161 VDD.n8140 0.000620321
R44046 VDD.n8142 VDD.n2089 0.000620321
R44047 VDD.n5575 VDD.n5553 0.000620321
R44048 VDD.n5556 VDD.n5555 0.000620321
R44049 VDD.n5657 VDD.n5544 0.000620321
R44050 VDD.n5638 VDD.n5546 0.000620321
R44051 VDD.n5840 VDD.n5819 0.000620321
R44052 VDD.n5821 VDD.n5680 0.000620321
R44053 VDD.n5773 VDD.n5752 0.000620321
R44054 VDD.n5754 VDD.n5704 0.000620321
R44055 VDD.n9004 VDD.n8953 0.000620321
R44056 VDD.n9002 VDD.n9001 0.000620321
R44057 VDD.n8833 VDD.n8812 0.000620321
R44058 VDD.n8831 VDD.n8525 0.000620321
R44059 VDD.n9120 VDD.n9099 0.000620321
R44060 VDD.n9118 VDD.n9090 0.000620321
R44061 VDD.n165 VDD.n144 0.000620321
R44062 VDD.n163 VDD.n135 0.000620321
R44063 VDD.n76 VDD.n55 0.000620321
R44064 VDD.n74 VDD.n46 0.000620321
R44065 VDD.n985 VDD.n984 0.000618343
R44066 VDD.n1033 VDD.n1032 0.000618343
R44067 VDD.n1627 VDD.n1626 0.00060181
R44068 VDD.n11048 VDD.n669 0.000601447
R44069 VDD.n11084 VDD.n657 0.000601447
R44070 VDD.n11123 VDD.n640 0.000601447
R44071 VDD.n11120 VDD.n11119 0.000584539
R44072 VDD.n1567 VDD.n782 0.000576357
R44073 VDD.n1566 VDD.n1565 0.000576357
R44074 VDD.n1568 VDD.n1510 0.000576357
R44075 VDD.n1426 VDD.n1425 0.000551724
R44076 VDD.n1431 VDD.n844 0.000551724
R44077 VDD.n1691 VDD.n738 0.000551724
R44078 VDD.n1690 VDD.n739 0.000551724
R44079 VDD.n7780 VDD.n7779 0.000534911
R44080 VDD.n11127 VDD.n11126 0.000533816
R44081 VDD.n11130 VDD.n633 0.000533816
R44082 VDD.n7744 VDD.n2270 0.000517455
R44083 a_52635_49681.n19 a_52635_49681.n17 7.94229
R44084 a_52635_49681.n193 a_52635_49681.n190 7.94229
R44085 a_52635_49681.n147 a_52635_49681.t81 6.58663
R44086 a_52635_49681.n103 a_52635_49681.t2 6.58663
R44087 a_52635_49681.n148 a_52635_49681.n145 5.95439
R44088 a_52635_49681.n104 a_52635_49681.n101 5.95439
R44089 a_52635_49681.n16 a_52635_49681.t111 5.69423
R44090 a_52635_49681.n20 a_52635_49681.t175 5.69423
R44091 a_52635_49681.n192 a_52635_49681.t151 5.69423
R44092 a_52635_49681.n188 a_52635_49681.t120 5.69423
R44093 a_52635_49681.n16 a_52635_49681.n15 5.49558
R44094 a_52635_49681.n192 a_52635_49681.n191 5.49558
R44095 a_52635_49681.n145 a_52635_49681.t9 5.31528
R44096 a_52635_49681.n101 a_52635_49681.t17 5.31528
R44097 a_52635_49681.n0 a_52635_49681.n12 4.22068
R44098 a_52635_49681.n1 a_52635_49681.t126 5.69068
R44099 a_52635_49681.n2 a_52635_49681.n57 4.22068
R44100 a_52635_49681.n3 a_52635_49681.t100 5.69068
R44101 a_52635_49681.n4 a_52635_49681.n56 4.22068
R44102 a_52635_49681.n6 a_52635_49681.n64 3.84173
R44103 a_52635_49681.n9 a_52635_49681.n60 3.84173
R44104 a_52635_49681.n11 a_52635_49681.n197 4.22067
R44105 a_52635_49681.n5 a_52635_49681.t31 5.31173
R44106 a_52635_49681.n7 a_52635_49681.t57 5.31173
R44107 a_52635_49681.n8 a_52635_49681.t27 5.31173
R44108 a_52635_49681.n10 a_52635_49681.t46 5.31173
R44109 a_52635_49681.n144 a_52635_49681.n142 4.50663
R44110 a_52635_49681.n100 a_52635_49681.n59 4.50663
R44111 a_52635_49681.n65 a_52635_49681.n7 4.46113
R44112 a_52635_49681.n19 a_52635_49681.n18 4.22423
R44113 a_52635_49681.n190 a_52635_49681.n189 4.22423
R44114 a_52635_49681.n26 a_52635_49681.t156 4.05054
R44115 a_52635_49681.n31 a_52635_49681.t150 4.05054
R44116 a_52635_49681.n33 a_52635_49681.t147 4.05054
R44117 a_52635_49681.n40 a_52635_49681.t138 4.05054
R44118 a_52635_49681.n42 a_52635_49681.t144 4.05054
R44119 a_52635_49681.n48 a_52635_49681.t142 4.05054
R44120 a_52635_49681.n50 a_52635_49681.t116 4.05054
R44121 a_52635_49681.n21 a_52635_49681.t140 4.05054
R44122 a_52635_49681.n159 a_52635_49681.t131 4.05054
R44123 a_52635_49681.n164 a_52635_49681.t127 4.05054
R44124 a_52635_49681.n166 a_52635_49681.t123 4.05054
R44125 a_52635_49681.n173 a_52635_49681.t105 4.05054
R44126 a_52635_49681.n175 a_52635_49681.t117 4.05054
R44127 a_52635_49681.n181 a_52635_49681.t114 4.05054
R44128 a_52635_49681.n183 a_52635_49681.t94 4.05054
R44129 a_52635_49681.n154 a_52635_49681.t107 4.05054
R44130 a_52635_49681.n150 a_52635_49681.n55 3.97558
R44131 a_52635_49681.n26 a_52635_49681.t135 3.87765
R44132 a_52635_49681.n31 a_52635_49681.t133 3.87765
R44133 a_52635_49681.n33 a_52635_49681.t129 3.87765
R44134 a_52635_49681.n40 a_52635_49681.t109 3.87765
R44135 a_52635_49681.n42 a_52635_49681.t124 3.87765
R44136 a_52635_49681.n48 a_52635_49681.t119 3.87765
R44137 a_52635_49681.n50 a_52635_49681.t98 3.87765
R44138 a_52635_49681.n21 a_52635_49681.t113 3.87765
R44139 a_52635_49681.n159 a_52635_49681.t173 3.87765
R44140 a_52635_49681.n164 a_52635_49681.t169 3.87765
R44141 a_52635_49681.n166 a_52635_49681.t168 3.87765
R44142 a_52635_49681.n173 a_52635_49681.t149 3.87765
R44143 a_52635_49681.n175 a_52635_49681.t164 3.87765
R44144 a_52635_49681.n181 a_52635_49681.t162 3.87765
R44145 a_52635_49681.n183 a_52635_49681.t137 3.87765
R44146 a_52635_49681.n154 a_52635_49681.t154 3.87765
R44147 a_52635_49681.n147 a_52635_49681.n146 3.84528
R44148 a_52635_49681.n144 a_52635_49681.n143 3.84528
R44149 a_52635_49681.n103 a_52635_49681.n102 3.84528
R44150 a_52635_49681.n100 a_52635_49681.n99 3.84528
R44151 a_52635_49681.n136 a_52635_49681.n132 3.79678
R44152 a_52635_49681.n119 a_52635_49681.n115 3.79678
R44153 a_52635_49681.n77 a_52635_49681.n73 3.79678
R44154 a_52635_49681.n92 a_52635_49681.n88 3.79678
R44155 a_52635_49681.n108 a_52635_49681.n10 3.87644
R44156 a_52635_49681.n128 a_52635_49681.n124 3.73034
R44157 a_52635_49681.n97 a_52635_49681.n81 3.73034
R44158 a_52635_49681.n53 a_52635_49681.n20 3.25667
R44159 a_52635_49681.n153 a_52635_49681.n4 3.15553
R44160 a_52635_49681.n54 a_52635_49681.n11 3.15589
R44161 a_52635_49681.n148 a_52635_49681.n147 3.00663
R44162 a_52635_49681.n104 a_52635_49681.n103 3.00663
R44163 a_52635_49681.n111 a_52635_49681.n109 2.7866
R44164 a_52635_49681.n114 a_52635_49681.n112 2.7866
R44165 a_52635_49681.n118 a_52635_49681.n116 2.7866
R44166 a_52635_49681.n122 a_52635_49681.n120 2.7866
R44167 a_52635_49681.n127 a_52635_49681.n125 2.7866
R44168 a_52635_49681.n131 a_52635_49681.n129 2.7866
R44169 a_52635_49681.n135 a_52635_49681.n133 2.7866
R44170 a_52635_49681.n139 a_52635_49681.n137 2.7866
R44171 a_52635_49681.n84 a_52635_49681.n82 2.7866
R44172 a_52635_49681.n87 a_52635_49681.n85 2.7866
R44173 a_52635_49681.n91 a_52635_49681.n89 2.7866
R44174 a_52635_49681.n95 a_52635_49681.n93 2.7866
R44175 a_52635_49681.n80 a_52635_49681.n78 2.7866
R44176 a_52635_49681.n76 a_52635_49681.n74 2.7866
R44177 a_52635_49681.n72 a_52635_49681.n70 2.7866
R44178 a_52635_49681.n68 a_52635_49681.n66 2.7866
R44179 a_52635_49681.n25 a_52635_49681.n21 2.73714
R44180 a_52635_49681.n158 a_52635_49681.n154 2.73714
R44181 a_52635_49681.n30 a_52635_49681.n26 2.73672
R44182 a_52635_49681.n163 a_52635_49681.n159 2.73672
R44183 a_52635_49681.n115 a_52635_49681.n111 2.73672
R44184 a_52635_49681.n88 a_52635_49681.n84 2.73672
R44185 a_52635_49681.n43 a_52635_49681.n41 2.60203
R44186 a_52635_49681.n176 a_52635_49681.n174 2.60203
R44187 a_52635_49681.n29 a_52635_49681.n28 2.58054
R44188 a_52635_49681.n38 a_52635_49681.n37 2.58054
R44189 a_52635_49681.n46 a_52635_49681.n45 2.58054
R44190 a_52635_49681.n24 a_52635_49681.n23 2.58054
R44191 a_52635_49681.n162 a_52635_49681.n161 2.58054
R44192 a_52635_49681.n171 a_52635_49681.n170 2.58054
R44193 a_52635_49681.n179 a_52635_49681.n178 2.58054
R44194 a_52635_49681.n157 a_52635_49681.n156 2.58054
R44195 a_52635_49681.n51 a_52635_49681.n49 2.53418
R44196 a_52635_49681.n34 a_52635_49681.n32 2.53418
R44197 a_52635_49681.n184 a_52635_49681.n182 2.53418
R44198 a_52635_49681.n167 a_52635_49681.n165 2.53418
R44199 a_52635_49681.n188 a_52635_49681.n187 2.51873
R44200 a_52635_49681.n29 a_52635_49681.n27 2.40765
R44201 a_52635_49681.n38 a_52635_49681.n36 2.40765
R44202 a_52635_49681.n46 a_52635_49681.n44 2.40765
R44203 a_52635_49681.n24 a_52635_49681.n22 2.40765
R44204 a_52635_49681.n162 a_52635_49681.n160 2.40765
R44205 a_52635_49681.n171 a_52635_49681.n169 2.40765
R44206 a_52635_49681.n179 a_52635_49681.n177 2.40765
R44207 a_52635_49681.n157 a_52635_49681.n155 2.40765
R44208 a_52635_49681.n107 a_52635_49681.n8 2.37644
R44209 a_52635_49681.n63 a_52635_49681.n5 2.37644
R44210 a_52635_49681.n17 a_52635_49681.n13 2.23844
R44211 a_52635_49681.n111 a_52635_49681.n110 2.2016
R44212 a_52635_49681.n114 a_52635_49681.n113 2.2016
R44213 a_52635_49681.n118 a_52635_49681.n117 2.2016
R44214 a_52635_49681.n122 a_52635_49681.n121 2.2016
R44215 a_52635_49681.n127 a_52635_49681.n126 2.2016
R44216 a_52635_49681.n131 a_52635_49681.n130 2.2016
R44217 a_52635_49681.n135 a_52635_49681.n134 2.2016
R44218 a_52635_49681.n139 a_52635_49681.n138 2.2016
R44219 a_52635_49681.n84 a_52635_49681.n83 2.2016
R44220 a_52635_49681.n87 a_52635_49681.n86 2.2016
R44221 a_52635_49681.n91 a_52635_49681.n90 2.2016
R44222 a_52635_49681.n95 a_52635_49681.n94 2.2016
R44223 a_52635_49681.n80 a_52635_49681.n79 2.2016
R44224 a_52635_49681.n76 a_52635_49681.n75 2.2016
R44225 a_52635_49681.n72 a_52635_49681.n71 2.2016
R44226 a_52635_49681.n68 a_52635_49681.n67 2.2016
R44227 a_52635_49681.n98 a_52635_49681.n63 2.0852
R44228 a_52635_49681.n142 a_52635_49681.n55 1.85726
R44229 a_52635_49681.n151 a_52635_49681.n150 1.83738
R44230 a_52635_49681.n141 a_52635_49681.n140 1.65018
R44231 a_52635_49681.n69 a_52635_49681.n65 1.65018
R44232 a_52635_49681.n152 a_52635_49681.n2 1.65553
R44233 a_52635_49681.n196 a_52635_49681.n0 1.65553
R44234 a_52635_49681.n186 a_52635_49681.n185 1.5005
R44235 a_52635_49681.n53 a_52635_49681.n52 1.5005
R44236 a_52635_49681.n105 a_52635_49681.n104 1.5005
R44237 a_52635_49681.n107 a_52635_49681.n106 1.5005
R44238 a_52635_49681.n149 a_52635_49681.n148 1.5005
R44239 a_52635_49681.n98 a_52635_49681.n97 1.5005
R44240 a_52635_49681.n124 a_52635_49681.n58 1.5005
R44241 a_52635_49681.n152 a_52635_49681.n151 1.5005
R44242 a_52635_49681.n168 a_52635_49681.n14 1.5005
R44243 a_52635_49681.n194 a_52635_49681.n193 1.5005
R44244 a_52635_49681.n35 a_52635_49681.n13 1.5005
R44245 a_52635_49681.n196 a_52635_49681.n195 1.5005
R44246 a_52635_49681.n12 a_52635_49681.t121 1.4705
R44247 a_52635_49681.n12 a_52635_49681.t93 1.4705
R44248 a_52635_49681.n15 a_52635_49681.t88 1.4705
R44249 a_52635_49681.n15 a_52635_49681.t128 1.4705
R44250 a_52635_49681.n18 a_52635_49681.t170 1.4705
R44251 a_52635_49681.n18 a_52635_49681.t115 1.4705
R44252 a_52635_49681.n27 a_52635_49681.t91 1.4705
R44253 a_52635_49681.n27 a_52635_49681.t166 1.4705
R44254 a_52635_49681.n28 a_52635_49681.t108 1.4705
R44255 a_52635_49681.n28 a_52635_49681.t97 1.4705
R44256 a_52635_49681.n36 a_52635_49681.t155 1.4705
R44257 a_52635_49681.n36 a_52635_49681.t125 1.4705
R44258 a_52635_49681.n37 a_52635_49681.t89 1.4705
R44259 a_52635_49681.n37 a_52635_49681.t145 1.4705
R44260 a_52635_49681.n44 a_52635_49681.t163 1.4705
R44261 a_52635_49681.n44 a_52635_49681.t134 1.4705
R44262 a_52635_49681.n45 a_52635_49681.t96 1.4705
R44263 a_52635_49681.n45 a_52635_49681.t153 1.4705
R44264 a_52635_49681.n22 a_52635_49681.t143 1.4705
R44265 a_52635_49681.n22 a_52635_49681.t112 1.4705
R44266 a_52635_49681.n23 a_52635_49681.t171 1.4705
R44267 a_52635_49681.n23 a_52635_49681.t139 1.4705
R44268 a_52635_49681.n191 a_52635_49681.t122 1.4705
R44269 a_52635_49681.n191 a_52635_49681.t167 1.4705
R44270 a_52635_49681.n189 a_52635_49681.t110 1.4705
R44271 a_52635_49681.n189 a_52635_49681.t157 1.4705
R44272 a_52635_49681.n160 a_52635_49681.t132 1.4705
R44273 a_52635_49681.n160 a_52635_49681.t104 1.4705
R44274 a_52635_49681.n161 a_52635_49681.t90 1.4705
R44275 a_52635_49681.n161 a_52635_49681.t161 1.4705
R44276 a_52635_49681.n169 a_52635_49681.t101 1.4705
R44277 a_52635_49681.n169 a_52635_49681.t165 1.4705
R44278 a_52635_49681.n170 a_52635_49681.t148 1.4705
R44279 a_52635_49681.n170 a_52635_49681.t118 1.4705
R44280 a_52635_49681.n177 a_52635_49681.t103 1.4705
R44281 a_52635_49681.n177 a_52635_49681.t172 1.4705
R44282 a_52635_49681.n178 a_52635_49681.t160 1.4705
R44283 a_52635_49681.n178 a_52635_49681.t130 1.4705
R44284 a_52635_49681.n155 a_52635_49681.t95 1.4705
R44285 a_52635_49681.n155 a_52635_49681.t152 1.4705
R44286 a_52635_49681.n156 a_52635_49681.t141 1.4705
R44287 a_52635_49681.n156 a_52635_49681.t106 1.4705
R44288 a_52635_49681.n57 a_52635_49681.t99 1.4705
R44289 a_52635_49681.n57 a_52635_49681.t159 1.4705
R44290 a_52635_49681.n56 a_52635_49681.t158 1.4705
R44291 a_52635_49681.n56 a_52635_49681.t146 1.4705
R44292 a_52635_49681.n62 a_52635_49681.t55 1.4705
R44293 a_52635_49681.n62 a_52635_49681.t26 1.4705
R44294 a_52635_49681.n64 a_52635_49681.t62 1.4705
R44295 a_52635_49681.n64 a_52635_49681.t29 1.4705
R44296 a_52635_49681.n109 a_52635_49681.t48 1.4705
R44297 a_52635_49681.n109 a_52635_49681.t70 1.4705
R44298 a_52635_49681.n110 a_52635_49681.t43 1.4705
R44299 a_52635_49681.n110 a_52635_49681.t66 1.4705
R44300 a_52635_49681.n112 a_52635_49681.t74 1.4705
R44301 a_52635_49681.n112 a_52635_49681.t35 1.4705
R44302 a_52635_49681.n113 a_52635_49681.t68 1.4705
R44303 a_52635_49681.n113 a_52635_49681.t30 1.4705
R44304 a_52635_49681.n116 a_52635_49681.t84 1.4705
R44305 a_52635_49681.n116 a_52635_49681.t78 1.4705
R44306 a_52635_49681.n117 a_52635_49681.t72 1.4705
R44307 a_52635_49681.n117 a_52635_49681.t69 1.4705
R44308 a_52635_49681.n120 a_52635_49681.t16 1.4705
R44309 a_52635_49681.n120 a_52635_49681.t58 1.4705
R44310 a_52635_49681.n121 a_52635_49681.t7 1.4705
R44311 a_52635_49681.n121 a_52635_49681.t50 1.4705
R44312 a_52635_49681.n125 a_52635_49681.t71 1.4705
R44313 a_52635_49681.n125 a_52635_49681.t85 1.4705
R44314 a_52635_49681.n126 a_52635_49681.t67 1.4705
R44315 a_52635_49681.n126 a_52635_49681.t73 1.4705
R44316 a_52635_49681.n129 a_52635_49681.t3 1.4705
R44317 a_52635_49681.n129 a_52635_49681.t49 1.4705
R44318 a_52635_49681.n130 a_52635_49681.t80 1.4705
R44319 a_52635_49681.n130 a_52635_49681.t44 1.4705
R44320 a_52635_49681.n133 a_52635_49681.t13 1.4705
R44321 a_52635_49681.n133 a_52635_49681.t32 1.4705
R44322 a_52635_49681.n134 a_52635_49681.t1 1.4705
R44323 a_52635_49681.n134 a_52635_49681.t28 1.4705
R44324 a_52635_49681.n137 a_52635_49681.t12 1.4705
R44325 a_52635_49681.n137 a_52635_49681.t63 1.4705
R44326 a_52635_49681.n138 a_52635_49681.t0 1.4705
R44327 a_52635_49681.n138 a_52635_49681.t59 1.4705
R44328 a_52635_49681.n82 a_52635_49681.t54 1.4705
R44329 a_52635_49681.n82 a_52635_49681.t77 1.4705
R44330 a_52635_49681.n83 a_52635_49681.t51 1.4705
R44331 a_52635_49681.n83 a_52635_49681.t75 1.4705
R44332 a_52635_49681.n85 a_52635_49681.t83 1.4705
R44333 a_52635_49681.n85 a_52635_49681.t37 1.4705
R44334 a_52635_49681.n86 a_52635_49681.t82 1.4705
R44335 a_52635_49681.n86 a_52635_49681.t36 1.4705
R44336 a_52635_49681.n89 a_52635_49681.t6 1.4705
R44337 a_52635_49681.n89 a_52635_49681.t87 1.4705
R44338 a_52635_49681.n90 a_52635_49681.t4 1.4705
R44339 a_52635_49681.n90 a_52635_49681.t86 1.4705
R44340 a_52635_49681.n93 a_52635_49681.t24 1.4705
R44341 a_52635_49681.n93 a_52635_49681.t61 1.4705
R44342 a_52635_49681.n94 a_52635_49681.t23 1.4705
R44343 a_52635_49681.n94 a_52635_49681.t60 1.4705
R44344 a_52635_49681.n78 a_52635_49681.t79 1.4705
R44345 a_52635_49681.n78 a_52635_49681.t8 1.4705
R44346 a_52635_49681.n79 a_52635_49681.t76 1.4705
R44347 a_52635_49681.n79 a_52635_49681.t5 1.4705
R44348 a_52635_49681.n74 a_52635_49681.t11 1.4705
R44349 a_52635_49681.n74 a_52635_49681.t56 1.4705
R44350 a_52635_49681.n75 a_52635_49681.t10 1.4705
R44351 a_52635_49681.n75 a_52635_49681.t53 1.4705
R44352 a_52635_49681.n70 a_52635_49681.t21 1.4705
R44353 a_52635_49681.n70 a_52635_49681.t34 1.4705
R44354 a_52635_49681.n71 a_52635_49681.t19 1.4705
R44355 a_52635_49681.n71 a_52635_49681.t33 1.4705
R44356 a_52635_49681.n66 a_52635_49681.t20 1.4705
R44357 a_52635_49681.n66 a_52635_49681.t65 1.4705
R44358 a_52635_49681.n67 a_52635_49681.t18 1.4705
R44359 a_52635_49681.n67 a_52635_49681.t64 1.4705
R44360 a_52635_49681.n146 a_52635_49681.t14 1.4705
R44361 a_52635_49681.n146 a_52635_49681.t38 1.4705
R44362 a_52635_49681.n143 a_52635_49681.t39 1.4705
R44363 a_52635_49681.n143 a_52635_49681.t42 1.4705
R44364 a_52635_49681.n61 a_52635_49681.t45 1.4705
R44365 a_52635_49681.n61 a_52635_49681.t15 1.4705
R44366 a_52635_49681.n60 a_52635_49681.t52 1.4705
R44367 a_52635_49681.n60 a_52635_49681.t25 1.4705
R44368 a_52635_49681.n102 a_52635_49681.t22 1.4705
R44369 a_52635_49681.n102 a_52635_49681.t40 1.4705
R44370 a_52635_49681.n99 a_52635_49681.t41 1.4705
R44371 a_52635_49681.n99 a_52635_49681.t47 1.4705
R44372 a_52635_49681.n197 a_52635_49681.t92 1.4705
R44373 a_52635_49681.t174 a_52635_49681.n197 1.4705
R44374 a_52635_49681.n30 a_52635_49681.n29 1.46537
R44375 a_52635_49681.n32 a_52635_49681.n31 1.46537
R44376 a_52635_49681.n39 a_52635_49681.n38 1.46537
R44377 a_52635_49681.n41 a_52635_49681.n40 1.46537
R44378 a_52635_49681.n43 a_52635_49681.n42 1.46537
R44379 a_52635_49681.n47 a_52635_49681.n46 1.46537
R44380 a_52635_49681.n49 a_52635_49681.n48 1.46537
R44381 a_52635_49681.n25 a_52635_49681.n24 1.46537
R44382 a_52635_49681.n163 a_52635_49681.n162 1.46537
R44383 a_52635_49681.n165 a_52635_49681.n164 1.46537
R44384 a_52635_49681.n172 a_52635_49681.n171 1.46537
R44385 a_52635_49681.n174 a_52635_49681.n173 1.46537
R44386 a_52635_49681.n176 a_52635_49681.n175 1.46537
R44387 a_52635_49681.n180 a_52635_49681.n179 1.46537
R44388 a_52635_49681.n182 a_52635_49681.n181 1.46537
R44389 a_52635_49681.n158 a_52635_49681.n157 1.46537
R44390 a_52635_49681.n115 a_52635_49681.n114 1.46537
R44391 a_52635_49681.n119 a_52635_49681.n118 1.46537
R44392 a_52635_49681.n123 a_52635_49681.n122 1.46537
R44393 a_52635_49681.n128 a_52635_49681.n127 1.46537
R44394 a_52635_49681.n132 a_52635_49681.n131 1.46537
R44395 a_52635_49681.n136 a_52635_49681.n135 1.46537
R44396 a_52635_49681.n140 a_52635_49681.n139 1.46537
R44397 a_52635_49681.n88 a_52635_49681.n87 1.46537
R44398 a_52635_49681.n92 a_52635_49681.n91 1.46537
R44399 a_52635_49681.n96 a_52635_49681.n95 1.46537
R44400 a_52635_49681.n81 a_52635_49681.n80 1.46537
R44401 a_52635_49681.n77 a_52635_49681.n76 1.46537
R44402 a_52635_49681.n73 a_52635_49681.n72 1.46537
R44403 a_52635_49681.n69 a_52635_49681.n68 1.46537
R44404 a_52635_49681.n34 a_52635_49681.n33 1.46535
R44405 a_52635_49681.n51 a_52635_49681.n50 1.46535
R44406 a_52635_49681.n167 a_52635_49681.n166 1.46535
R44407 a_52635_49681.n184 a_52635_49681.n183 1.46535
R44408 a_52635_49681.n20 a_52635_49681.n19 1.27228
R44409 a_52635_49681.n49 a_52635_49681.n47 1.27228
R44410 a_52635_49681.n47 a_52635_49681.n43 1.27228
R44411 a_52635_49681.n41 a_52635_49681.n39 1.27228
R44412 a_52635_49681.n32 a_52635_49681.n30 1.27228
R44413 a_52635_49681.n190 a_52635_49681.n188 1.27228
R44414 a_52635_49681.n182 a_52635_49681.n180 1.27228
R44415 a_52635_49681.n180 a_52635_49681.n176 1.27228
R44416 a_52635_49681.n174 a_52635_49681.n172 1.27228
R44417 a_52635_49681.n165 a_52635_49681.n163 1.27228
R44418 a_52635_49681.n140 a_52635_49681.n136 1.27228
R44419 a_52635_49681.n132 a_52635_49681.n128 1.27228
R44420 a_52635_49681.n123 a_52635_49681.n119 1.27228
R44421 a_52635_49681.n73 a_52635_49681.n69 1.27228
R44422 a_52635_49681.n81 a_52635_49681.n77 1.27228
R44423 a_52635_49681.n96 a_52635_49681.n92 1.27228
R44424 a_52635_49681.n145 a_52635_49681.n144 1.27228
R44425 a_52635_49681.n101 a_52635_49681.n100 1.27228
R44426 a_52635_49681.n150 a_52635_49681.n149 1.25341
R44427 a_52635_49681.n153 a_52635_49681.n55 1.23151
R44428 a_52635_49681.n17 a_52635_49681.n16 1.01873
R44429 a_52635_49681.n193 a_52635_49681.n192 1.01873
R44430 a_52635_49681.n54 a_52635_49681.n53 0.778574
R44431 a_52635_49681.n186 a_52635_49681.n153 0.778574
R44432 a_52635_49681.n195 a_52635_49681.n13 0.778574
R44433 a_52635_49681.n151 a_52635_49681.n14 0.778574
R44434 a_52635_49681.n187 a_52635_49681.n186 0.738439
R44435 a_52635_49681.n194 a_52635_49681.n14 0.738439
R44436 a_52635_49681.n142 a_52635_49681.n141 0.737223
R44437 a_52635_49681.n65 a_52635_49681.n59 0.737223
R44438 a_52635_49681.n149 a_52635_49681.n58 0.737223
R44439 a_52635_49681.n105 a_52635_49681.n98 0.737223
R44440 a_52635_49681.n108 a_52635_49681.n59 0.725061
R44441 a_52635_49681.n106 a_52635_49681.n105 0.725061
R44442 a_52635_49681.n52 a_52635_49681.n51 0.699581
R44443 a_52635_49681.n35 a_52635_49681.n34 0.699581
R44444 a_52635_49681.n185 a_52635_49681.n184 0.699581
R44445 a_52635_49681.n168 a_52635_49681.n167 0.699581
R44446 a_52635_49681.n141 a_52635_49681.n108 0.585196
R44447 a_52635_49681.n106 a_52635_49681.n58 0.585196
R44448 a_52635_49681.n52 a_52635_49681.n25 0.557791
R44449 a_52635_49681.n39 a_52635_49681.n35 0.557791
R44450 a_52635_49681.n185 a_52635_49681.n158 0.557791
R44451 a_52635_49681.n172 a_52635_49681.n168 0.557791
R44452 a_52635_49681.n187 a_52635_49681.n54 0.530466
R44453 a_52635_49681.n195 a_52635_49681.n194 0.530466
R44454 a_52635_49681.n124 a_52635_49681.n123 0.150184
R44455 a_52635_49681.n97 a_52635_49681.n96 0.150184
R44456 a_52635_49681.n3 a_52635_49681.n4 1.27228
R44457 a_52635_49681.n152 a_52635_49681.n3 7.30549
R44458 a_52635_49681.t102 a_52635_49681.n2 6.96214
R44459 a_52635_49681.n9 a_52635_49681.n10 1.26457
R44460 a_52635_49681.n107 a_52635_49681.n9 6.59229
R44461 a_52635_49681.n61 a_52635_49681.n8 5.10549
R44462 a_52635_49681.n6 a_52635_49681.n7 1.26457
R44463 a_52635_49681.n63 a_52635_49681.n6 6.59229
R44464 a_52635_49681.n62 a_52635_49681.n5 5.10549
R44465 a_52635_49681.n11 a_52635_49681.n1 1.27192
R44466 a_52635_49681.n196 a_52635_49681.n1 7.30549
R44467 a_52635_49681.t136 a_52635_49681.n0 6.96214
R44468 a_57977_n12421.t0 a_57977_n12421.t1 93.1589
R44469 a_57977_n12421.t0 a_57977_n12421.t2 24.9014
R44470 a_100820_11614.n2 a_100820_11614.t19 12.8637
R44471 a_100820_11614.n1 a_100820_11614.t1 10.7018
R44472 a_100820_11614.n1 a_100820_11614.t7 10.1659
R44473 a_100820_11614.n1 a_100820_11614.t6 9.64387
R44474 a_100820_11614.t0 a_100820_11614.n1 9.27665
R44475 a_100820_11614.n1 a_100820_11614.n2 8.75198
R44476 a_100820_11614.n2 a_100820_11614.t14 8.14051
R44477 a_100820_11614.n2 a_100820_11614.t10 8.14051
R44478 a_100820_11614.n2 a_100820_11614.t8 8.14051
R44479 a_100820_11614.n2 a_100820_11614.t17 8.14051
R44480 a_100820_11614.n2 a_100820_11614.t21 8.06917
R44481 a_100820_11614.n2 a_100820_11614.t18 8.06917
R44482 a_100820_11614.n2 a_100820_11614.t11 8.06917
R44483 a_100820_11614.n2 a_100820_11614.t15 8.06917
R44484 a_100820_11614.n2 a_100820_11614.t13 8.06917
R44485 a_100820_11614.n2 a_100820_11614.t23 8.06917
R44486 a_100820_11614.n2 a_100820_11614.t9 8.06917
R44487 a_100820_11614.n0 a_100820_11614.t4 7.94068
R44488 a_100820_11614.n1 a_100820_11614.t2 7.72524
R44489 a_100820_11614.n0 a_100820_11614.t5 7.22855
R44490 a_100820_11614.n1 a_100820_11614.t3 7.17942
R44491 a_100820_11614.t16 a_100820_11614.n2 8.33649
R44492 a_100820_11614.n2 a_100820_11614.t20 8.33649
R44493 a_100820_11614.t22 a_100820_11614.n2 8.33556
R44494 a_100820_11614.n2 a_100820_11614.t12 8.33556
R44495 a_100820_11614.n1 a_100820_11614.n0 7.46075
R44496 a_30324_4421.t2 a_30324_4421.t0 21.6693
R44497 a_30324_4421.t1 a_30324_4421.t0 15.3476
R44498 a_31284_4481.t0 a_31284_4481.t2 41.3314
R44499 a_31284_4481.t2 a_31284_4481.t1 15.0742
R44500 a_100820_10448.t0 a_100820_10448.t7 12.7127
R44501 a_100820_10448.t0 a_100820_10448.t10 10.2828
R44502 a_100820_10448.t0 a_100820_10448.t8 10.2828
R44503 a_100820_10448.t0 a_100820_10448.t18 10.2828
R44504 a_100820_10448.t0 a_100820_10448.t14 10.2828
R44505 a_100820_10448.t0 a_100820_10448.t21 10.1333
R44506 a_100820_10448.t0 a_100820_10448.t22 10.1333
R44507 a_100820_10448.t0 a_100820_10448.t6 10.1333
R44508 a_100820_10448.t0 a_100820_10448.t4 10.1333
R44509 a_100820_10448.t0 a_100820_10448.t3 9.72545
R44510 a_100820_10448.t0 a_100820_10448.t17 9.57156
R44511 a_100820_10448.t0 a_100820_10448.t15 9.57156
R44512 a_100820_10448.t0 a_100820_10448.t16 9.57156
R44513 a_100820_10448.t0 a_100820_10448.t12 9.57156
R44514 a_100820_10448.t0 a_100820_10448.t23 9.57156
R44515 a_100820_10448.t0 a_100820_10448.t19 9.57156
R44516 a_100820_10448.t0 a_100820_10448.t20 9.57156
R44517 a_100820_10448.t0 a_100820_10448.t13 9.57156
R44518 a_100820_10448.t3 a_100820_10448.t2 8.02945
R44519 a_100820_10448.t0 a_100820_10448.t1 8.02708
R44520 a_100820_10448.t0 a_100820_10448.t9 7.90829
R44521 a_100820_10448.t0 a_100820_10448.t11 7.90829
R44522 a_100820_10448.t5 a_100820_10448.t0 7.41776
R44523 a_53829_n36382.n5 a_53829_n36382.n1 10.2377
R44524 a_53829_n36382.n4 a_53829_n36382.t0 10.2105
R44525 a_53829_n36382.n4 a_53829_n36382.t1 9.99998
R44526 a_53829_n36382.n5 a_53829_n36382.t7 9.80532
R44527 a_53829_n36382.n5 a_53829_n36382.t5 9.55206
R44528 a_53829_n36382.n0 a_53829_n36382.t9 8.17385
R44529 a_53829_n36382.n3 a_53829_n36382.t21 8.17299
R44530 a_53829_n36382.n3 a_53829_n36382.t10 8.17134
R44531 a_53829_n36382.n0 a_53829_n36382.t23 8.16754
R44532 a_53829_n36382.n1 a_53829_n36382.t17 8.10567
R44533 a_53829_n36382.n1 a_53829_n36382.t20 8.10567
R44534 a_53829_n36382.n3 a_53829_n36382.t16 8.10567
R44535 a_53829_n36382.n3 a_53829_n36382.t11 8.10567
R44536 a_53829_n36382.n1 a_53829_n36382.t18 8.10567
R44537 a_53829_n36382.n1 a_53829_n36382.t19 8.10567
R44538 a_53829_n36382.n0 a_53829_n36382.t15 8.10567
R44539 a_53829_n36382.n0 a_53829_n36382.t14 8.10567
R44540 a_53829_n36382.n6 a_53829_n36382.t3 7.74888
R44541 a_53829_n36382.n7 a_53829_n36382.t6 7.73141
R44542 a_53829_n36382.n6 a_53829_n36382.t2 7.46359
R44543 a_53829_n36382.t4 a_53829_n36382.n7 7.13081
R44544 a_53829_n36382.n4 a_53829_n36382.n6 2.2505
R44545 a_53829_n36382.n7 a_53829_n36382.n5 2.2505
R44546 a_53829_n36382.t8 a_53829_n36382.n1 8.35729
R44547 a_53829_n36382.n1 a_53829_n36382.t22 8.37586
R44548 a_53829_n36382.n0 a_53829_n36382.t12 8.38104
R44549 a_53829_n36382.n1 a_53829_n36382.n0 4.35658
R44550 a_53829_n36382.n5 a_53829_n36382.n4 2.96863
R44551 a_53829_n36382.n2 a_53829_n36382.n1 1.08819
R44552 a_53829_n36382.n2 a_53829_n36382.n3 1.08408
R44553 a_53829_n36382.n2 a_53829_n36382.t13 8.6675
R44554 a_36032_n36322.n1 a_36032_n36322.n0 26.5241
R44555 a_36032_n36322.n1 a_36032_n36322.t1 11.5094
R44556 a_36032_n36322.n0 a_36032_n36322.t2 10.937
R44557 a_36032_n36322.n0 a_36032_n36322.t3 9.33982
R44558 a_36032_n36322.t0 a_36032_n36322.n1 9.24966
R44559 a_35502_25545.n345 a_35502_25545.t22 10.621
R44560 a_35502_25545.n349 a_35502_25545.t71 10.621
R44561 a_35502_25545.n342 a_35502_25545.n326 10.3121
R44562 a_35502_25545.n347 a_35502_25545.t91 10.3044
R44563 a_35502_25545.n351 a_35502_25545.t20 10.3044
R44564 a_35502_25545.n346 a_35502_25545.t48 9.9994
R44565 a_35502_25545.n350 a_35502_25545.t26 9.9994
R44566 a_35502_25545.n345 a_35502_25545.t24 9.999
R44567 a_35502_25545.n349 a_35502_25545.t62 9.999
R44568 a_35502_25545.n224 a_35502_25545.t39 8.33806
R44569 a_35502_25545.n319 a_35502_25545.t64 8.3366
R44570 a_35502_25545.n278 a_35502_25545.t35 8.26493
R44571 a_35502_25545.n96 a_35502_25545.t69 8.35715
R44572 a_35502_25545.n43 a_35502_25545.t81 8.06917
R44573 a_35502_25545.n55 a_35502_25545.t77 8.06917
R44574 a_35502_25545.n122 a_35502_25545.t102 8.06917
R44575 a_35502_25545.n31 a_35502_25545.t85 8.06917
R44576 a_35502_25545.n132 a_35502_25545.t30 8.06917
R44577 a_35502_25545.n50 a_35502_25545.t47 8.06917
R44578 a_35502_25545.n57 a_35502_25545.t51 8.06917
R44579 a_35502_25545.n17 a_35502_25545.t80 8.06917
R44580 a_35502_25545.n78 a_35502_25545.t100 8.06917
R44581 a_35502_25545.n28 a_35502_25545.t45 8.06917
R44582 a_35502_25545.n133 a_35502_25545.t72 8.06917
R44583 a_35502_25545.n9 a_35502_25545.t29 8.06917
R44584 a_35502_25545.n8 a_35502_25545.t59 8.06917
R44585 a_35502_25545.n170 a_35502_25545.t56 8.06917
R44586 a_35502_25545.n6 a_35502_25545.t57 8.06917
R44587 a_35502_25545.n5 a_35502_25545.t86 8.06917
R44588 a_35502_25545.n175 a_35502_25545.t83 8.06917
R44589 a_35502_25545.n40 a_35502_25545.t76 8.06917
R44590 a_35502_25545.n93 a_35502_25545.t44 8.06917
R44591 a_35502_25545.n75 a_35502_25545.t78 8.06917
R44592 a_35502_25545.n61 a_35502_25545.t103 8.06917
R44593 a_35502_25545.n34 a_35502_25545.t41 8.06917
R44594 a_35502_25545.n90 a_35502_25545.t49 8.06917
R44595 a_35502_25545.n2 a_35502_25545.t75 8.06917
R44596 a_35502_25545.n86 a_35502_25545.t95 8.06917
R44597 a_35502_25545.n71 a_35502_25545.t40 8.06917
R44598 a_35502_25545.n65 a_35502_25545.t68 8.06917
R44599 a_35502_25545.n125 a_35502_25545.t28 8.06917
R44600 a_35502_25545.n23 a_35502_25545.t54 8.06917
R44601 a_35502_25545.n163 a_35502_25545.t52 8.06917
R44602 a_35502_25545.n128 a_35502_25545.t53 8.06917
R44603 a_35502_25545.n20 a_35502_25545.t82 8.06917
R44604 a_35502_25545.n152 a_35502_25545.t79 8.06917
R44605 a_35502_25545.n82 a_35502_25545.t73 8.06917
R44606 a_35502_25545.n68 a_35502_25545.t96 8.06917
R44607 a_35502_25545.n108 a_35502_25545.t66 8.06917
R44608 a_35502_25545.n97 a_35502_25545.t74 8.06917
R44609 a_35502_25545.n259 a_35502_25545.t97 8.06917
R44610 a_35502_25545.n248 a_35502_25545.t36 8.06917
R44611 a_35502_25545.n247 a_35502_25545.t42 8.06917
R44612 a_35502_25545.n246 a_35502_25545.t88 8.06917
R44613 a_35502_25545.n95 a_35502_25545.t101 8.06917
R44614 a_35502_25545.n239 a_35502_25545.t46 8.06917
R44615 a_35502_25545.n112 a_35502_25545.t98 8.06917
R44616 a_35502_25545.n225 a_35502_25545.t94 8.06917
R44617 a_35502_25545.n231 a_35502_25545.t63 8.06917
R44618 a_35502_25545.n232 a_35502_25545.t67 8.06917
R44619 a_35502_25545.n233 a_35502_25545.t38 8.06917
R44620 a_35502_25545.n109 a_35502_25545.t37 8.06917
R44621 a_35502_25545.n100 a_35502_25545.t65 8.06917
R44622 a_35502_25545.n267 a_35502_25545.t89 8.06917
R44623 a_35502_25545.n318 a_35502_25545.t99 8.06917
R44624 a_35502_25545.n118 a_35502_25545.t43 8.06917
R44625 a_35502_25545.n316 a_35502_25545.t84 8.06917
R44626 a_35502_25545.n315 a_35502_25545.t33 8.06917
R44627 a_35502_25545.n314 a_35502_25545.t31 8.06917
R44628 a_35502_25545.n312 a_35502_25545.t61 8.06917
R44629 a_35502_25545.n305 a_35502_25545.t70 8.06917
R44630 a_35502_25545.n115 a_35502_25545.t92 8.06917
R44631 a_35502_25545.n300 a_35502_25545.t34 8.06917
R44632 a_35502_25545.n101 a_35502_25545.t60 8.06917
R44633 a_35502_25545.n119 a_35502_25545.t87 8.06917
R44634 a_35502_25545.n289 a_35502_25545.t32 8.06917
R44635 a_35502_25545.n288 a_35502_25545.t58 8.06917
R44636 a_35502_25545.n287 a_35502_25545.t55 8.06917
R44637 a_35502_25545.n274 a_35502_25545.t93 8.06917
R44638 a_35502_25545.n277 a_35502_25545.t90 8.06917
R44639 a_35502_25545.n330 a_35502_25545.t5 6.49245
R44640 a_35502_25545.n327 a_35502_25545.t17 6.49245
R44641 a_35502_25545.n138 a_35502_25545.t2 6.50349
R44642 a_35502_25545.n343 a_35502_25545.t23 5.70664
R44643 a_35502_25545.n353 a_35502_25545.t21 5.23357
R44644 a_35502_25545.n328 a_35502_25545.t19 5.22068
R44645 a_35502_25545.t27 a_35502_25545.n353 5.15077
R44646 a_35502_25545.n343 a_35502_25545.t25 4.6582
R44647 a_35502_25545.n84 a_35502_25545.n69 2.0194
R44648 a_35502_25545.n178 a_35502_25545.n123 2.42484
R44649 a_35502_25545.n123 a_35502_25545.n177 2.4256
R44650 a_35502_25545.n110 a_35502_25545.n109 2.25048
R44651 a_35502_25545.n115 a_35502_25545.n113 2.25048
R44652 a_35502_25545.n134 a_35502_25545.t4 5.23239
R44653 a_35502_25545.n135 a_35502_25545.t12 5.23239
R44654 a_35502_25545.n339 a_35502_25545.n338 4.60825
R44655 a_35502_25545.t8 a_35502_25545.n138 5.23239
R44656 a_35502_25545.n10 a_35502_25545.n9 1.44552
R44657 a_35502_25545.n7 a_35502_25545.n6 1.44552
R44658 a_35502_25545.n126 a_35502_25545.n125 2.22591
R44659 a_35502_25545.n129 a_35502_25545.n128 2.22591
R44660 a_35502_25545.n85 a_35502_25545.n159 4.51491
R44661 a_35502_25545.n216 a_35502_25545.n215 4.51075
R44662 a_35502_25545.n62 a_35502_25545.n61 2.21906
R44663 a_35502_25545.n66 a_35502_25545.n65 2.21906
R44664 a_35502_25545.n34 a_35502_25545.n35 2.21826
R44665 a_35502_25545.n40 a_35502_25545.n39 2.21826
R44666 a_35502_25545.n338 a_35502_25545.n334 4.50168
R44667 a_35502_25545.n12 a_35502_25545.n5 2.21666
R44668 a_35502_25545.n11 a_35502_25545.n174 4.5005
R44669 a_35502_25545.n184 a_35502_25545.n183 4.5005
R44670 a_35502_25545.n14 a_35502_25545.n8 2.21666
R44671 a_35502_25545.n13 a_35502_25545.n169 4.5005
R44672 a_35502_25545.n202 a_35502_25545.n201 4.5005
R44673 a_35502_25545.n194 a_35502_25545.n193 4.5005
R44674 a_35502_25545.n78 a_35502_25545.n79 2.21666
R44675 a_35502_25545.n191 a_35502_25545.n27 4.5005
R44676 a_35502_25545.n28 a_35502_25545.n25 2.21666
R44677 a_35502_25545.n26 a_35502_25545.n190 4.5005
R44678 a_35502_25545.n189 a_35502_25545.n133 4.5005
R44679 a_35502_25545.n188 a_35502_25545.n187 4.5005
R44680 a_35502_25545.n51 a_35502_25545.n50 2.21666
R44681 a_35502_25545.n196 a_35502_25545.n49 4.5005
R44682 a_35502_25545.n198 a_35502_25545.n197 4.5005
R44683 a_35502_25545.n58 a_35502_25545.n57 2.21666
R44684 a_35502_25545.n16 a_35502_25545.n171 4.5005
R44685 a_35502_25545.n18 a_35502_25545.n17 2.21666
R44686 a_35502_25545.n0 a_35502_25545.n1 0.0657695
R44687 a_35502_25545.n30 a_35502_25545.n206 4.5005
R44688 a_35502_25545.n32 a_35502_25545.n31 2.21666
R44689 a_35502_25545.n131 a_35502_25545.n205 4.5005
R44690 a_35502_25545.n132 a_35502_25545.n204 4.5005
R44691 a_35502_25545.n208 a_35502_25545.n203 4.5005
R44692 a_35502_25545.n44 a_35502_25545.n43 2.21666
R44693 a_35502_25545.n42 a_35502_25545.n181 4.5005
R44694 a_35502_25545.n180 a_35502_25545.n54 4.5005
R44695 a_35502_25545.n55 a_35502_25545.n52 2.21666
R44696 a_35502_25545.n53 a_35502_25545.n178 4.5005
R44697 a_35502_25545.n123 a_35502_25545.n122 0.0107891
R44698 a_35502_25545.n127 a_35502_25545.n158 4.5005
R44699 a_35502_25545.n21 a_35502_25545.n20 2.21666
R44700 a_35502_25545.n19 a_35502_25545.n151 4.5005
R44701 a_35502_25545.n157 a_35502_25545.n156 4.5005
R44702 a_35502_25545.n124 a_35502_25545.n166 4.5005
R44703 a_35502_25545.n24 a_35502_25545.n23 2.21666
R44704 a_35502_25545.n22 a_35502_25545.n162 4.5005
R44705 a_35502_25545.n165 a_35502_25545.n164 4.5005
R44706 a_35502_25545.n65 a_35502_25545.n67 2.21666
R44707 a_35502_25545.n64 a_35502_25545.n107 4.5005
R44708 a_35502_25545.n71 a_35502_25545.n73 2.21666
R44709 a_35502_25545.n70 a_35502_25545.n105 4.5005
R44710 a_35502_25545.n86 a_35502_25545.n88 2.21666
R44711 a_35502_25545.n215 a_35502_25545.n214 4.5005
R44712 a_35502_25545.n2 a_35502_25545.n3 2.21666
R44713 a_35502_25545.n90 a_35502_25545.n92 2.21666
R44714 a_35502_25545.n89 a_35502_25545.n102 4.5005
R44715 a_35502_25545.n160 a_35502_25545.n120 4.5005
R44716 a_35502_25545.n36 a_35502_25545.n34 2.21666
R44717 a_35502_25545.n61 a_35502_25545.n63 2.21666
R44718 a_35502_25545.n60 a_35502_25545.n106 4.5005
R44719 a_35502_25545.n75 a_35502_25545.n77 2.21666
R44720 a_35502_25545.n74 a_35502_25545.n104 4.5005
R44721 a_35502_25545.n68 a_35502_25545.n69 0.0231698
R44722 a_35502_25545.n82 a_35502_25545.n84 2.21666
R44723 a_35502_25545.n153 a_35502_25545.n81 4.5005
R44724 a_35502_25545.n121 a_35502_25545.n154 4.5005
R44725 a_35502_25545.n41 a_35502_25545.n40 2.21666
R44726 a_35502_25545.n83 a_35502_25545.n82 2.21666
R44727 a_35502_25545.n81 a_35502_25545.n103 4.5005
R44728 a_35502_25545.n38 a_35502_25545.n121 4.5005
R44729 a_35502_25545.n64 a_35502_25545.n219 4.5005
R44730 a_35502_25545.n72 a_35502_25545.n71 2.21666
R44731 a_35502_25545.n70 a_35502_25545.n218 4.5005
R44732 a_35502_25545.n87 a_35502_25545.n86 2.21666
R44733 a_35502_25545.n85 a_35502_25545.n217 4.5005
R44734 a_35502_25545.n2 a_35502_25545.n4 2.21666
R44735 a_35502_25545.n91 a_35502_25545.n90 2.21666
R44736 a_35502_25545.n89 a_35502_25545.n213 4.5005
R44737 a_35502_25545.n212 a_35502_25545.n120 4.5005
R44738 a_35502_25545.n60 a_35502_25545.n168 4.5005
R44739 a_35502_25545.n76 a_35502_25545.n75 2.21666
R44740 a_35502_25545.n74 a_35502_25545.n167 4.5005
R44741 a_35502_25545.n94 a_35502_25545.n93 0.023589
R44742 a_35502_25545.n56 a_35502_25545.n55 2.21666
R44743 a_35502_25545.n179 a_35502_25545.n54 4.5005
R44744 a_35502_25545.n42 a_35502_25545.n176 4.5005
R44745 a_35502_25545.n43 a_35502_25545.n45 2.21666
R44746 a_35502_25545.n53 a_35502_25545.n177 4.5005
R44747 a_35502_25545.n80 a_35502_25545.n78 2.21666
R44748 a_35502_25545.n193 a_35502_25545.n192 4.5005
R44749 a_35502_25545.n187 a_35502_25545.n186 4.5005
R44750 a_35502_25545.n185 a_35502_25545.n133 4.5005
R44751 a_35502_25545.n26 a_35502_25545.n173 4.5005
R44752 a_35502_25545.n29 a_35502_25545.n28 2.21666
R44753 a_35502_25545.n27 a_35502_25545.n172 4.5005
R44754 a_35502_25545.n57 a_35502_25545.n59 2.21666
R44755 a_35502_25545.n199 a_35502_25545.n198 4.5005
R44756 a_35502_25545.n47 a_35502_25545.n49 4.5005
R44757 a_35502_25545.n50 a_35502_25545.n48 2.21666
R44758 a_35502_25545.n17 a_35502_25545.n15 2.21666
R44759 a_35502_25545.n195 a_35502_25545.n16 4.5005
R44760 a_35502_25545.n209 a_35502_25545.n208 4.5005
R44761 a_35502_25545.n132 a_35502_25545.n130 4.5005
R44762 a_35502_25545.n131 a_35502_25545.n207 4.5005
R44763 a_35502_25545.n33 a_35502_25545.n31 2.21666
R44764 a_35502_25545.n30 a_35502_25545.n0 0.0743189
R44765 a_35502_25545.n299 a_35502_25545.n148 4.5005
R44766 a_35502_25545.n279 a_35502_25545.n276 4.5005
R44767 a_35502_25545.n281 a_35502_25545.n280 4.5005
R44768 a_35502_25545.n282 a_35502_25545.n275 4.5005
R44769 a_35502_25545.n284 a_35502_25545.n283 4.5005
R44770 a_35502_25545.n286 a_35502_25545.n285 4.5005
R44771 a_35502_25545.n291 a_35502_25545.n290 4.5005
R44772 a_35502_25545.n119 a_35502_25545.n292 4.5005
R44773 a_35502_25545.n293 a_35502_25545.n149 4.5005
R44774 a_35502_25545.n295 a_35502_25545.n294 4.5005
R44775 a_35502_25545.n296 a_35502_25545.n101 4.5005
R44776 a_35502_25545.n298 a_35502_25545.n297 4.5005
R44777 a_35502_25545.n302 a_35502_25545.n114 4.5005
R44778 a_35502_25545.n304 a_35502_25545.n303 4.5005
R44779 a_35502_25545.n306 a_35502_25545.n147 4.5005
R44780 a_35502_25545.n308 a_35502_25545.n307 4.5005
R44781 a_35502_25545.n309 a_35502_25545.n146 4.5005
R44782 a_35502_25545.n311 a_35502_25545.n310 4.5005
R44783 a_35502_25545.n313 a_35502_25545.n145 4.5005
R44784 a_35502_25545.n323 a_35502_25545.n322 4.5005
R44785 a_35502_25545.n118 a_35502_25545.n116 4.5005
R44786 a_35502_25545.n117 a_35502_25545.n321 4.5005
R44787 a_35502_25545.n320 a_35502_25545.n317 4.5005
R44788 a_35502_25545.n230 a_35502_25545.n222 4.5005
R44789 a_35502_25545.n112 a_35502_25545.n229 4.5005
R44790 a_35502_25545.n228 a_35502_25545.n111 4.5005
R44791 a_35502_25545.n227 a_35502_25545.n226 4.5005
R44792 a_35502_25545.n270 a_35502_25545.n269 4.5005
R44793 a_35502_25545.n268 a_35502_25545.n223 4.5005
R44794 a_35502_25545.n266 a_35502_25545.n265 4.5005
R44795 a_35502_25545.n264 a_35502_25545.n98 4.5005
R44796 a_35502_25545.n263 a_35502_25545.n100 4.5005
R44797 a_35502_25545.n99 a_35502_25545.n234 4.5005
R44798 a_35502_25545.n262 a_35502_25545.n261 4.5005
R44799 a_35502_25545.n250 a_35502_25545.n249 4.5005
R44800 a_35502_25545.n108 a_35502_25545.n251 4.5005
R44801 a_35502_25545.n252 a_35502_25545.n236 4.5005
R44802 a_35502_25545.n254 a_35502_25545.n253 4.5005
R44803 a_35502_25545.n255 a_35502_25545.n97 4.5005
R44804 a_35502_25545.n257 a_35502_25545.n256 4.5005
R44805 a_35502_25545.n258 a_35502_25545.n235 4.5005
R44806 a_35502_25545.n245 a_35502_25545.n244 4.5005
R44807 a_35502_25545.n243 a_35502_25545.n237 4.5005
R44808 a_35502_25545.n242 a_35502_25545.n241 4.5005
R44809 a_35502_25545.n240 a_35502_25545.n238 4.5005
R44810 a_35502_25545.n337 a_35502_25545.n336 4.5005
R44811 a_35502_25545.n137 a_35502_25545.n136 2.24327
R44812 a_35502_25545.n141 a_35502_25545.n139 4.5005
R44813 a_35502_25545.n142 a_35502_25545.n140 2.24296
R44814 a_35502_25545.n338 a_35502_25545.t3 3.83265
R44815 a_35502_25545.n335 a_35502_25545.t10 3.82765
R44816 a_35502_25545.n142 a_35502_25545.t14 3.82673
R44817 a_35502_25545.n332 a_35502_25545.t1 3.78255
R44818 a_35502_25545.n136 a_35502_25545.t6 3.76633
R44819 a_35502_25545.n330 a_35502_25545.t13 3.75068
R44820 a_35502_25545.n327 a_35502_25545.t0 3.75068
R44821 a_35502_25545.n329 a_35502_25545.t7 3.74975
R44822 a_35502_25545.n221 a_35502_25545.n143 3.37223
R44823 a_35502_25545.n113 a_35502_25545.n301 3.02216
R44824 a_35502_25545.n217 a_35502_25545.n216 2.89625
R44825 a_35502_25545.n18 a_35502_25545.n194 2.95081
R44826 a_35502_25545.n214 a_35502_25545.n159 2.88162
R44827 a_35502_25545.n192 a_35502_25545.n15 2.95081
R44828 a_35502_25545.n344 a_35502_25545.n342 2.76066
R44829 a_35502_25545.n344 a_35502_25545.n343 2.57313
R44830 a_35502_25545.n69 a_35502_25545.n83 2.00991
R44831 a_35502_25545.n272 a_35502_25545.n271 2.30989
R44832 a_35502_25545.n325 a_35502_25545.n144 2.30989
R44833 a_35502_25545.n301 a_35502_25545.n300 2.29659
R44834 a_35502_25545.n260 a_35502_25545.n259 2.2812
R44835 a_35502_25545.n331 a_35502_25545.n329 2.24389
R44836 a_35502_25545.n200 a_35502_25545.n170 2.23529
R44837 a_35502_25545.n182 a_35502_25545.n175 2.23529
R44838 a_35502_25545.n163 a_35502_25545.n161 2.23423
R44839 a_35502_25545.n155 a_35502_25545.n152 2.23423
R44840 a_35502_25545.n285 a_35502_25545.n273 2.18975
R44841 a_35502_25545.n324 a_35502_25545.n145 2.18975
R44842 a_35502_25545.n271 a_35502_25545.n222 2.16725
R44843 a_35502_25545.n250 a_35502_25545.n144 2.16725
R44844 a_35502_25545.n221 a_35502_25545.n220 2.11247
R44845 a_35502_25545.n186 a_35502_25545.n150 2.102
R44846 a_35502_25545.n46 a_35502_25545.n209 2.102
R44847 a_35502_25545.n341 a_35502_25545.n333 2.07395
R44848 a_35502_25545.n220 a_35502_25545.n150 2.07182
R44849 a_35502_25545.n210 a_35502_25545.n46 2.07182
R44850 a_35502_25545.n37 a_35502_25545.n66 2.13751
R44851 a_35502_25545.n211 a_35502_25545.n62 2.13751
R44852 a_35502_25545.n342 a_35502_25545.n341 1.90955
R44853 a_35502_25545.n353 a_35502_25545.n352 1.71486
R44854 a_35502_25545.n210 a_35502_25545.n143 1.50911
R44855 a_35502_25545.n220 a_35502_25545.n37 1.5005
R44856 a_35502_25545.n211 a_35502_25545.n210 1.5005
R44857 a_35502_25545.n273 a_35502_25545.n272 1.5005
R44858 a_35502_25545.n325 a_35502_25545.n324 1.5005
R44859 a_35502_25545.n341 a_35502_25545.n340 1.5005
R44860 a_35502_25545.n352 a_35502_25545.n351 1.5005
R44861 a_35502_25545.n348 a_35502_25545.n347 1.5005
R44862 a_35502_25545.t10 a_35502_25545.t15 1.4705
R44863 a_35502_25545.t13 a_35502_25545.t18 1.4705
R44864 a_35502_25545.t1 a_35502_25545.t9 1.4705
R44865 a_35502_25545.t0 a_35502_25545.t16 1.4705
R44866 a_35502_25545.n279 a_35502_25545.n278 1.39514
R44867 a_35502_25545.n272 a_35502_25545.n221 1.39023
R44868 a_35502_25545.n326 a_35502_25545.n325 1.39023
R44869 a_35502_25545.n328 a_35502_25545.n327 1.27228
R44870 a_35502_25545.n314 a_35502_25545.n313 1.26997
R44871 a_35502_25545.n287 a_35502_25545.n286 1.26997
R44872 a_35502_25545.n322 a_35502_25545.n316 1.24392
R44873 a_35502_25545.n290 a_35502_25545.n289 1.24392
R44874 a_35502_25545.n249 a_35502_25545.n248 1.24204
R44875 a_35502_25545.n231 a_35502_25545.n230 1.24204
R44876 a_35502_25545.n331 a_35502_25545.n330 1.20682
R44877 a_35502_25545.n246 a_35502_25545.n245 1.20414
R44878 a_35502_25545.n269 a_35502_25545.n233 1.20414
R44879 a_35502_25545.n320 a_35502_25545.n319 1.14132
R44880 a_35502_25545.n332 a_35502_25545.n140 1.20835
R44881 a_35502_25545.n227 a_35502_25545.n224 1.13598
R44882 a_35502_25545.n339 a_35502_25545.n335 1.13573
R44883 a_35502_25545.n346 a_35502_25545.n345 0.90675
R44884 a_35502_25545.n350 a_35502_25545.n349 0.90675
R44885 a_35502_25545.n335 a_35502_25545.n135 0.939226
R44886 a_35502_25545.n291 a_35502_25545.n273 0.752
R44887 a_35502_25545.n324 a_35502_25545.n323 0.752
R44888 a_35502_25545.n271 a_35502_25545.n270 0.71825
R44889 a_35502_25545.n244 a_35502_25545.n144 0.71825
R44890 a_35502_25545.n315 a_35502_25545.n314 0.663658
R44891 a_35502_25545.n316 a_35502_25545.n315 0.663658
R44892 a_35502_25545.n288 a_35502_25545.n287 0.663658
R44893 a_35502_25545.n289 a_35502_25545.n288 0.663658
R44894 a_35502_25545.n247 a_35502_25545.n246 0.655156
R44895 a_35502_25545.n248 a_35502_25545.n247 0.655156
R44896 a_35502_25545.n233 a_35502_25545.n232 0.655156
R44897 a_35502_25545.n232 a_35502_25545.n231 0.655156
R44898 a_35502_25545.n326 a_35502_25545.n143 0.603852
R44899 a_35502_25545.n333 a_35502_25545.n332 0.596867
R44900 a_35502_25545.n96 a_35502_25545.n95 0.313126
R44901 a_35502_25545.n278 a_35502_25545.n277 0.432797
R44902 a_35502_25545.n304 a_35502_25545.n114 0.394842
R44903 a_35502_25545.n299 a_35502_25545.n298 0.394842
R44904 a_35502_25545.n117 a_35502_25545.n317 0.381816
R44905 a_35502_25545.n294 a_35502_25545.n293 0.381816
R44906 a_35502_25545.n241 a_35502_25545.n240 0.379447
R44907 a_35502_25545.n258 a_35502_25545.n257 0.379447
R44908 a_35502_25545.n253 a_35502_25545.n252 0.379447
R44909 a_35502_25545.n266 a_35502_25545.n98 0.379447
R44910 a_35502_25545.n99 a_35502_25545.n262 0.379447
R44911 a_35502_25545.n226 a_35502_25545.n111 0.379447
R44912 a_35502_25545.n178 a_35502_25545.n52 0.44431
R44913 a_35502_25545.n79 a_35502_25545.n191 0.44431
R44914 a_35502_25545.n58 a_35502_25545.n171 0.44431
R44915 a_35502_25545.n1 a_35502_25545.n206 1.94004
R44916 a_35502_25545.n88 a_35502_25545.n105 0.44431
R44917 a_35502_25545.n94 a_35502_25545.n104 1.95665
R44918 a_35502_25545.n56 a_35502_25545.n177 0.44431
R44919 a_35502_25545.n80 a_35502_25545.n172 0.44431
R44920 a_35502_25545.n59 a_35502_25545.n195 0.44431
R44921 a_35502_25545.n297 a_35502_25545.n148 0.375125
R44922 a_35502_25545.n303 a_35502_25545.n302 0.375125
R44923 a_35502_25545.n190 a_35502_25545.n25 0.431935
R44924 a_35502_25545.n32 a_35502_25545.n205 0.431935
R44925 a_35502_25545.n73 a_35502_25545.n107 0.431935
R44926 a_35502_25545.n77 a_35502_25545.n106 0.431935
R44927 a_35502_25545.n29 a_35502_25545.n173 0.431935
R44928 a_35502_25545.n207 a_35502_25545.n33 0.431935
R44929 a_35502_25545.n295 a_35502_25545.n149 0.36275
R44930 a_35502_25545.n321 a_35502_25545.n320 0.36275
R44931 a_35502_25545.n183 a_35502_25545.n174 0.3605
R44932 a_35502_25545.n201 a_35502_25545.n169 0.3605
R44933 a_35502_25545.n156 a_35502_25545.n151 0.3605
R44934 a_35502_25545.n164 a_35502_25545.n162 0.3605
R44935 a_35502_25545.n38 a_35502_25545.n103 0.3605
R44936 a_35502_25545.n219 a_35502_25545.n72 0.429685
R44937 a_35502_25545.n218 a_35502_25545.n87 0.429685
R44938 a_35502_25545.n213 a_35502_25545.n212 0.3605
R44939 a_35502_25545.n168 a_35502_25545.n76 0.429685
R44940 a_35502_25545.n167 a_35502_25545.n94 1.93517
R44941 a_35502_25545.n228 a_35502_25545.n227 0.3605
R44942 a_35502_25545.n265 a_35502_25545.n264 0.3605
R44943 a_35502_25545.n261 a_35502_25545.n234 0.3605
R44944 a_35502_25545.n256 a_35502_25545.n235 0.3605
R44945 a_35502_25545.n254 a_35502_25545.n236 0.3605
R44946 a_35502_25545.n242 a_35502_25545.n238 0.3605
R44947 a_35502_25545.n333 a_35502_25545.n328 0.339591
R44948 a_35502_25545.n319 a_35502_25545.n318 0.335806
R44949 a_35502_25545.n225 a_35502_25545.n224 0.33475
R44950 a_35502_25545.n347 a_35502_25545.n346 0.320048
R44951 a_35502_25545.n351 a_35502_25545.n350 0.320048
R44952 a_35502_25545.n307 a_35502_25545.n146 0.302474
R44953 a_35502_25545.n282 a_35502_25545.n281 0.302474
R44954 a_35502_25545.n181 a_35502_25545.n180 0.287375
R44955 a_35502_25545.n197 a_35502_25545.n196 0.287375
R44956 a_35502_25545.n154 a_35502_25545.n153 0.287375
R44957 a_35502_25545.n160 a_35502_25545.n102 0.287375
R44958 a_35502_25545.n179 a_35502_25545.n176 0.287375
R44959 a_35502_25545.n47 a_35502_25545.n199 0.287375
R44960 a_35502_25545.n280 a_35502_25545.n275 0.287375
R44961 a_35502_25545.n309 a_35502_25545.n308 0.287375
R44962 a_35502_25545.n348 a_35502_25545.n344 0.212426
R44963 a_35502_25545.n156 a_35502_25545.n155 0.208888
R44964 a_35502_25545.n164 a_35502_25545.n161 0.208888
R44965 a_35502_25545.n183 a_35502_25545.n182 0.20887
R44966 a_35502_25545.n201 a_35502_25545.n200 0.20887
R44967 a_35502_25545.n139 a_35502_25545.n331 0.208385
R44968 a_35502_25545.n301 a_35502_25545.n148 0.208099
R44969 a_35502_25545.n260 a_35502_25545.n235 0.208099
R44970 a_35502_25545.n245 a_35502_25545.n237 0.147342
R44971 a_35502_25545.n257 a_35502_25545.n97 0.147342
R44972 a_35502_25545.n252 a_35502_25545.n108 0.147342
R44973 a_35502_25545.n269 a_35502_25545.n268 0.147342
R44974 a_35502_25545.n100 a_35502_25545.n98 0.147342
R44975 a_35502_25545.n112 a_35502_25545.n111 0.147342
R44976 a_35502_25545.n307 a_35502_25545.n306 0.147342
R44977 a_35502_25545.n311 a_35502_25545.n146 0.147342
R44978 a_35502_25545.n118 a_35502_25545.n117 0.147342
R44979 a_35502_25545.n281 a_35502_25545.n276 0.147342
R44980 a_35502_25545.n283 a_35502_25545.n282 0.147342
R44981 a_35502_25545.n293 a_35502_25545.n119 0.147342
R44982 a_35502_25545.n298 a_35502_25545.n101 0.147342
R44983 a_35502_25545.n180 a_35502_25545.n52 0.209185
R44984 a_35502_25545.n181 a_35502_25545.n44 0.209185
R44985 a_35502_25545.n182 a_35502_25545.n44 0.825446
R44986 a_35502_25545.n12 a_35502_25545.n174 0.209185
R44987 a_35502_25545.n7 a_35502_25545.n12 0.565419
R44988 a_35502_25545.n188 a_35502_25545.n7 0.834884
R44989 a_35502_25545.n189 a_35502_25545.n188 0.14
R44990 a_35502_25545.n190 a_35502_25545.n189 0.14
R44991 a_35502_25545.n191 a_35502_25545.n25 0.209185
R44992 a_35502_25545.n194 a_35502_25545.n79 0.209185
R44993 a_35502_25545.n18 a_35502_25545.n171 0.209185
R44994 a_35502_25545.n197 a_35502_25545.n58 0.209185
R44995 a_35502_25545.n196 a_35502_25545.n51 0.209185
R44996 a_35502_25545.n200 a_35502_25545.n51 0.825446
R44997 a_35502_25545.n14 a_35502_25545.n169 0.209185
R44998 a_35502_25545.n10 a_35502_25545.n14 0.565419
R44999 a_35502_25545.n203 a_35502_25545.n10 0.834884
R45000 a_35502_25545.n204 a_35502_25545.n203 0.14
R45001 a_35502_25545.n205 a_35502_25545.n204 0.14
R45002 a_35502_25545.n206 a_35502_25545.n32 0.209185
R45003 a_35502_25545.n153 a_35502_25545.n84 0.209185
R45004 a_35502_25545.n154 a_35502_25545.n41 0.209185
R45005 a_35502_25545.n155 a_35502_25545.n41 0.825427
R45006 a_35502_25545.n21 a_35502_25545.n151 0.209185
R45007 a_35502_25545.n158 a_35502_25545.n21 0.429685
R45008 a_35502_25545.n158 a_35502_25545.n129 0.208907
R45009 a_35502_25545.n67 a_35502_25545.n129 0.836657
R45010 a_35502_25545.n67 a_35502_25545.n107 0.209185
R45011 a_35502_25545.n73 a_35502_25545.n105 0.209185
R45012 a_35502_25545.n88 a_35502_25545.n159 0.209185
R45013 a_35502_25545.n214 a_35502_25545.n3 0.209185
R45014 a_35502_25545.n3 a_35502_25545.n92 0.513496
R45015 a_35502_25545.n92 a_35502_25545.n102 0.209185
R45016 a_35502_25545.n36 a_35502_25545.n160 0.209185
R45017 a_35502_25545.n36 a_35502_25545.n161 0.825427
R45018 a_35502_25545.n24 a_35502_25545.n162 0.209185
R45019 a_35502_25545.n166 a_35502_25545.n24 0.429685
R45020 a_35502_25545.n166 a_35502_25545.n126 0.208907
R45021 a_35502_25545.n63 a_35502_25545.n126 0.836657
R45022 a_35502_25545.n63 a_35502_25545.n106 0.209185
R45023 a_35502_25545.n77 a_35502_25545.n104 0.209185
R45024 a_35502_25545.n83 a_35502_25545.n103 0.209185
R45025 a_35502_25545.n39 a_35502_25545.n38 0.209137
R45026 a_35502_25545.n39 a_35502_25545.n37 0.886485
R45027 a_35502_25545.n219 a_35502_25545.n66 0.209113
R45028 a_35502_25545.n218 a_35502_25545.n72 0.209185
R45029 a_35502_25545.n217 a_35502_25545.n87 0.209185
R45030 a_35502_25545.n216 a_35502_25545.n4 0.209185
R45031 a_35502_25545.n91 a_35502_25545.n4 0.498871
R45032 a_35502_25545.n213 a_35502_25545.n91 0.209185
R45033 a_35502_25545.n212 a_35502_25545.n35 0.209137
R45034 a_35502_25545.n211 a_35502_25545.n35 0.886485
R45035 a_35502_25545.n168 a_35502_25545.n62 0.209113
R45036 a_35502_25545.n167 a_35502_25545.n76 0.209185
R45037 a_35502_25545.n56 a_35502_25545.n179 0.209185
R45038 a_35502_25545.n45 a_35502_25545.n176 0.209185
R45039 a_35502_25545.n150 a_35502_25545.n45 0.908935
R45040 a_35502_25545.n186 a_35502_25545.n185 0.14
R45041 a_35502_25545.n185 a_35502_25545.n173 0.14
R45042 a_35502_25545.n29 a_35502_25545.n172 0.209185
R45043 a_35502_25545.n192 a_35502_25545.n80 0.209185
R45044 a_35502_25545.n195 a_35502_25545.n15 0.209185
R45045 a_35502_25545.n199 a_35502_25545.n59 0.209185
R45046 a_35502_25545.n48 a_35502_25545.n47 0.209185
R45047 a_35502_25545.n48 a_35502_25545.n46 0.908935
R45048 a_35502_25545.n209 a_35502_25545.n130 0.14
R45049 a_35502_25545.n207 a_35502_25545.n130 0.14
R45050 a_35502_25545.n33 a_35502_25545.n0 1.54288
R45051 a_35502_25545.n280 a_35502_25545.n279 0.14
R45052 a_35502_25545.n284 a_35502_25545.n275 0.14
R45053 a_35502_25545.n285 a_35502_25545.n284 0.14
R45054 a_35502_25545.n292 a_35502_25545.n291 0.14
R45055 a_35502_25545.n292 a_35502_25545.n149 0.14
R45056 a_35502_25545.n296 a_35502_25545.n295 0.14
R45057 a_35502_25545.n297 a_35502_25545.n296 0.14
R45058 a_35502_25545.n302 a_35502_25545.n113 0.208168
R45059 a_35502_25545.n303 a_35502_25545.n147 0.14
R45060 a_35502_25545.n308 a_35502_25545.n147 0.14
R45061 a_35502_25545.n310 a_35502_25545.n309 0.14
R45062 a_35502_25545.n310 a_35502_25545.n145 0.14
R45063 a_35502_25545.n323 a_35502_25545.n116 0.14
R45064 a_35502_25545.n321 a_35502_25545.n116 0.14
R45065 a_35502_25545.n229 a_35502_25545.n228 0.14
R45066 a_35502_25545.n229 a_35502_25545.n222 0.14
R45067 a_35502_25545.n270 a_35502_25545.n223 0.14
R45068 a_35502_25545.n265 a_35502_25545.n223 0.14
R45069 a_35502_25545.n264 a_35502_25545.n263 0.14
R45070 a_35502_25545.n263 a_35502_25545.n234 0.14
R45071 a_35502_25545.n261 a_35502_25545.n110 0.208168
R45072 a_35502_25545.n110 a_35502_25545.n260 3.03679
R45073 a_35502_25545.n256 a_35502_25545.n255 0.14
R45074 a_35502_25545.n255 a_35502_25545.n254 0.14
R45075 a_35502_25545.n251 a_35502_25545.n236 0.14
R45076 a_35502_25545.n251 a_35502_25545.n250 0.14
R45077 a_35502_25545.n244 a_35502_25545.n243 0.14
R45078 a_35502_25545.n243 a_35502_25545.n242 0.14
R45079 a_35502_25545.n96 a_35502_25545.n238 1.12911
R45080 a_35502_25545.n137 a_35502_25545.n138 1.2061
R45081 a_35502_25545.n336 a_35502_25545.n137 0.230885
R45082 a_35502_25545.n336 a_35502_25545.n334 0.14
R45083 a_35502_25545.n134 a_35502_25545.n135 1.27228
R45084 a_35502_25545.t11 a_35502_25545.n134 6.50385
R45085 a_35502_25545.n140 a_35502_25545.n139 0.230894
R45086 a_35502_25545.n142 a_35502_25545.n141 0.138586
R45087 a_35502_25545.n337 a_35502_25545.n136 0.137318
R45088 a_35502_25545.n226 a_35502_25545.n225 0.128395
R45089 a_35502_25545.n318 a_35502_25545.n317 0.128395
R45090 a_35502_25545.n241 a_35502_25545.n239 0.118921
R45091 a_35502_25545.n259 a_35502_25545.n258 0.118921
R45092 a_35502_25545.n267 a_35502_25545.n266 0.118921
R45093 a_35502_25545.n313 a_35502_25545.n312 0.114184
R45094 a_35502_25545.n286 a_35502_25545.n274 0.114184
R45095 a_35502_25545.n305 a_35502_25545.n304 0.113
R45096 a_35502_25545.n338 a_35502_25545.n337 0.110782
R45097 a_35502_25545.n141 a_35502_25545.n329 0.109514
R45098 a_35502_25545.n13 a_35502_25545.n202 0.109179
R45099 a_35502_25545.n11 a_35502_25545.n184 0.109179
R45100 a_35502_25545.n57 a_35502_25545.n16 0.107155
R45101 a_35502_25545.n78 a_35502_25545.n27 0.107155
R45102 a_35502_25545.n55 a_35502_25545.n53 0.107155
R45103 a_35502_25545.n352 a_35502_25545.n348 0.105095
R45104 a_35502_25545.n131 a_35502_25545.n31 0.103632
R45105 a_35502_25545.n28 a_35502_25545.n26 0.103632
R45106 a_35502_25545.n300 a_35502_25545.n299 0.103526
R45107 a_35502_25545.n22 a_35502_25545.n165 0.102991
R45108 a_35502_25545.n124 a_35502_25545.n23 0.102991
R45109 a_35502_25545.n19 a_35502_25545.n157 0.102991
R45110 a_35502_25545.n127 a_35502_25545.n20 0.102991
R45111 a_35502_25545.n340 a_35502_25545.n339 0.0995
R45112 a_35502_25545.n75 a_35502_25545.n60 0.0933826
R45113 a_35502_25545.n71 a_35502_25545.n64 0.0933826
R45114 a_35502_25545.n93 a_35502_25545.n74 0.092742
R45115 a_35502_25545.n90 a_35502_25545.n2 0.092742
R45116 a_35502_25545.n86 a_35502_25545.n70 0.092742
R45117 a_35502_25545.n82 a_35502_25545.n68 0.092742
R45118 a_35502_25545.n198 a_35502_25545.n49 0.0821726
R45119 a_35502_25545.n42 a_35502_25545.n54 0.0821726
R45120 a_35502_25545.n120 a_35502_25545.n89 0.0821726
R45121 a_35502_25545.n121 a_35502_25545.n81 0.0821726
R45122 a_35502_25545.n128 a_35502_25545.n127 0.0427776
R45123 a_35502_25545.n125 a_35502_25545.n124 0.0427776
R45124 a_35502_25545.n340 a_35502_25545.n334 0.041
R45125 a_35502_25545.n132 a_35502_25545.n131 0.0402153
R45126 a_35502_25545.n26 a_35502_25545.n133 0.0402153
R45127 a_35502_25545.n53 a_35502_25545.n122 0.0402153
R45128 a_35502_25545.n187 a_35502_25545.n133 0.0402153
R45129 a_35502_25545.n208 a_35502_25545.n132 0.0402153
R45130 a_35502_25545.n306 a_35502_25545.n305 0.0348421
R45131 a_35502_25545.n277 a_35502_25545.n276 0.0348421
R45132 a_35502_25545.n202 a_35502_25545.n170 0.0344623
R45133 a_35502_25545.n184 a_35502_25545.n175 0.0344623
R45134 a_35502_25545.n312 a_35502_25545.n311 0.0336579
R45135 a_35502_25545.n283 a_35502_25545.n274 0.0336579
R45136 a_35502_25545.n165 a_35502_25545.n163 0.0325285
R45137 a_35502_25545.n157 a_35502_25545.n152 0.0325285
R45138 a_35502_25545.n239 a_35502_25545.n237 0.0289211
R45139 a_35502_25545.n268 a_35502_25545.n267 0.0289211
R45140 a_35502_25545.n240 a_35502_25545.n95 0.166289
R45141 a_35502_25545.n115 a_35502_25545.n114 0.156816
R45142 a_35502_25545.n262 a_35502_25545.n109 0.156816
R45143 a_35502_25545.n9 a_35502_25545.n8 0.154009
R45144 a_35502_25545.n6 a_35502_25545.n5 0.154009
R45145 a_35502_25545.n290 a_35502_25545.n119 0.147342
R45146 a_35502_25545.n322 a_35502_25545.n118 0.147342
R45147 a_35502_25545.n230 a_35502_25545.n112 0.147342
R45148 a_35502_25545.n249 a_35502_25545.n108 0.147342
R45149 a_35502_25545.n294 a_35502_25545.n101 0.147342
R45150 a_35502_25545.n100 a_35502_25545.n99 0.147342
R45151 a_35502_25545.n253 a_35502_25545.n97 0.147342
R45152 a_35502_25545.n90 a_35502_25545.n89 0.0943434
R45153 a_35502_25545.n82 a_35502_25545.n81 0.0943434
R45154 a_35502_25545.n75 a_35502_25545.n74 0.0901797
R45155 a_35502_25545.n71 a_35502_25545.n70 0.0901797
R45156 a_35502_25545.n8 a_35502_25545.n13 0.0847264
R45157 a_35502_25545.n5 a_35502_25545.n11 0.0847264
R45158 a_35502_25545.n86 a_35502_25545.n85 0.0799306
R45159 a_35502_25545.n193 a_35502_25545.n78 0.0799306
R45160 a_35502_25545.n65 a_35502_25545.n64 0.0799306
R45161 a_35502_25545.n61 a_35502_25545.n60 0.0799306
R45162 a_35502_25545.n198 a_35502_25545.n57 0.0799306
R45163 a_35502_25545.n55 a_35502_25545.n54 0.0799306
R45164 a_35502_25545.n50 a_35502_25545.n49 0.0799306
R45165 a_35502_25545.n43 a_35502_25545.n42 0.0799306
R45166 a_35502_25545.n121 a_35502_25545.n40 0.0799306
R45167 a_35502_25545.n120 a_35502_25545.n34 0.0799306
R45168 a_35502_25545.n31 a_35502_25545.n30 0.0799306
R45169 a_35502_25545.n28 a_35502_25545.n27 0.0799306
R45170 a_35502_25545.n23 a_35502_25545.n22 0.0799306
R45171 a_35502_25545.n20 a_35502_25545.n19 0.0799306
R45172 a_35502_25545.n17 a_35502_25545.n16 0.0799306
R45173 a_35502_25545.n215 a_35502_25545.n2 0.0799306
R45174 a_35502_25545.n1 a_35502_25545.t50 8.08727
R45175 a_33249_35053.n109 a_33249_35053.n106 9.23995
R45176 a_33249_35053.n35 a_33249_35053.n33 7.94229
R45177 a_33249_35053.n80 a_33249_35053.n77 7.94229
R45178 a_33249_35053.n108 a_33249_35053.t92 6.72766
R45179 a_33249_35053.n129 a_33249_35053.n127 6.58329
R45180 a_33249_35053.n106 a_33249_35053.n14 6.01251
R45181 a_33249_35053.n126 a_33249_35053.t130 5.85326
R45182 a_33249_35053.n130 a_33249_35053.t117 5.85326
R45183 a_33249_35053.n126 a_33249_35053.n125 5.84661
R45184 a_33249_35053.n32 a_33249_35053.t51 5.69423
R45185 a_33249_35053.n36 a_33249_35053.t61 5.69423
R45186 a_33249_35053.n79 a_33249_35053.t58 5.69423
R45187 a_33249_35053.n75 a_33249_35053.t64 5.69423
R45188 a_33249_35053.n32 a_33249_35053.n31 5.49558
R45189 a_33249_35053.n79 a_33249_35053.n78 5.49558
R45190 a_33249_35053.n157 a_33249_35053.n0 4.58971
R45191 a_33249_35053.n1 a_33249_35053.t126 5.84971
R45192 a_33249_35053.n2 a_33249_35053.n132 4.58971
R45193 a_33249_35053.n3 a_33249_35053.n103 4.22068
R45194 a_33249_35053.n4 a_33249_35053.t65 5.69068
R45195 a_33249_35053.n5 a_33249_35053.n102 4.22068
R45196 a_33249_35053.n6 a_33249_35053.n72 4.22068
R45197 a_33249_35053.t62 a_33249_35053.n7 5.69068
R45198 a_33249_35053.n71 a_33249_35053.n8 4.22068
R45199 a_33249_35053.n9 a_33249_35053.t103 5.47076
R45200 a_33249_35053.n129 a_33249_35053.n128 4.59326
R45201 a_33249_35053.n109 a_33249_35053.n108 4.52463
R45202 a_33249_35053.n110 a_33249_35053.t91 4.41563
R45203 a_33249_35053.n119 a_33249_35053.t0 4.41563
R45204 a_33249_35053.n35 a_33249_35053.n34 4.22423
R45205 a_33249_35053.n77 a_33249_35053.n76 4.22423
R45206 a_33249_35053.n108 a_33249_35053.n107 4.21432
R45207 a_33249_35053.n150 a_33249_35053.t139 4.21195
R45208 a_33249_35053.n152 a_33249_35053.t134 4.21195
R45209 a_33249_35053.n137 a_33249_35053.t123 4.21195
R45210 a_33249_35053.n135 a_33249_35053.t115 4.21195
R45211 a_33249_35053.n42 a_33249_35053.t30 4.05054
R45212 a_33249_35053.n47 a_33249_35053.t8 4.05054
R45213 a_33249_35053.n49 a_33249_35053.t39 4.05054
R45214 a_33249_35053.n56 a_33249_35053.t43 4.05054
R45215 a_33249_35053.n58 a_33249_35053.t33 4.05054
R45216 a_33249_35053.n64 a_33249_35053.t37 4.05054
R45217 a_33249_35053.n66 a_33249_35053.t69 4.05054
R45218 a_33249_35053.n37 a_33249_35053.t85 4.05054
R45219 a_33249_35053.n21 a_33249_35053.t34 4.05054
R45220 a_33249_35053.n26 a_33249_35053.t19 4.05054
R45221 a_33249_35053.n28 a_33249_35053.t53 4.05054
R45222 a_33249_35053.n88 a_33249_35053.t59 4.05054
R45223 a_33249_35053.n90 a_33249_35053.t42 4.05054
R45224 a_33249_35053.n96 a_33249_35053.t47 4.05054
R45225 a_33249_35053.n98 a_33249_35053.t79 4.05054
R45226 a_33249_35053.n16 a_33249_35053.t4 4.05054
R45227 a_33249_35053.n150 a_33249_35053.t106 4.03668
R45228 a_33249_35053.n152 a_33249_35053.t137 4.03668
R45229 a_33249_35053.n137 a_33249_35053.t124 4.03668
R45230 a_33249_35053.n135 a_33249_35053.t120 4.03668
R45231 a_33249_35053.n42 a_33249_35053.t32 3.87765
R45232 a_33249_35053.n47 a_33249_35053.t13 3.87765
R45233 a_33249_35053.n49 a_33249_35053.t48 3.87765
R45234 a_33249_35053.n56 a_33249_35053.t52 3.87765
R45235 a_33249_35053.n58 a_33249_35053.t38 3.87765
R45236 a_33249_35053.n64 a_33249_35053.t41 3.87765
R45237 a_33249_35053.n66 a_33249_35053.t73 3.87765
R45238 a_33249_35053.n37 a_33249_35053.t2 3.87765
R45239 a_33249_35053.n21 a_33249_35053.t36 3.87765
R45240 a_33249_35053.n26 a_33249_35053.t21 3.87765
R45241 a_33249_35053.n28 a_33249_35053.t56 3.87765
R45242 a_33249_35053.n88 a_33249_35053.t60 3.87765
R45243 a_33249_35053.n90 a_33249_35053.t44 3.87765
R45244 a_33249_35053.n96 a_33249_35053.t49 3.87765
R45245 a_33249_35053.n98 a_33249_35053.t80 3.87765
R45246 a_33249_35053.n16 a_33249_35053.t5 3.87765
R45247 a_33249_35053.n110 a_33249_35053.t105 3.833
R45248 a_33249_35053.n119 a_33249_35053.t96 3.833
R45249 a_33249_35053.n146 a_33249_35053.n142 3.81703
R45250 a_33249_35053.n133 a_33249_35053.n2 3.95161
R45251 a_33249_35053.n118 a_33249_35053.n114 3.80578
R45252 a_33249_35053.n123 a_33249_35053.n9 3.90344
R45253 a_33249_35053.n124 a_33249_35053.n10 3.69568
R45254 a_33249_35053.n69 a_33249_35053.n36 3.25667
R45255 a_33249_35053.n113 a_33249_35053.n111 3.15563
R45256 a_33249_35053.n117 a_33249_35053.n115 3.15563
R45257 a_33249_35053.n8 a_33249_35053.n70 3.15553
R45258 a_33249_35053.n105 a_33249_35053.n5 3.15553
R45259 a_33249_35053.n149 a_33249_35053.n148 2.95195
R45260 a_33249_35053.n145 a_33249_35053.n144 2.95195
R45261 a_33249_35053.n141 a_33249_35053.n140 2.95195
R45262 a_33249_35053.n13 a_33249_35053.n12 2.95195
R45263 a_33249_35053.n149 a_33249_35053.n147 2.77668
R45264 a_33249_35053.n145 a_33249_35053.n143 2.77668
R45265 a_33249_35053.n141 a_33249_35053.n139 2.77668
R45266 a_33249_35053.n13 a_33249_35053.n11 2.77668
R45267 a_33249_35053.n41 a_33249_35053.n37 2.73714
R45268 a_33249_35053.n20 a_33249_35053.n16 2.73714
R45269 a_33249_35053.n46 a_33249_35053.n42 2.73672
R45270 a_33249_35053.n25 a_33249_35053.n21 2.73672
R45271 a_33249_35053.n151 a_33249_35053.n149 2.71872
R45272 a_33249_35053.n114 a_33249_35053.n110 2.71872
R45273 a_33249_35053.n59 a_33249_35053.n57 2.60203
R45274 a_33249_35053.n91 a_33249_35053.n89 2.60203
R45275 a_33249_35053.n131 a_33249_35053.n124 2.5825
R45276 a_33249_35053.n45 a_33249_35053.n44 2.58054
R45277 a_33249_35053.n54 a_33249_35053.n53 2.58054
R45278 a_33249_35053.n62 a_33249_35053.n61 2.58054
R45279 a_33249_35053.n40 a_33249_35053.n39 2.58054
R45280 a_33249_35053.n24 a_33249_35053.n23 2.58054
R45281 a_33249_35053.n86 a_33249_35053.n85 2.58054
R45282 a_33249_35053.n94 a_33249_35053.n93 2.58054
R45283 a_33249_35053.n19 a_33249_35053.n18 2.58054
R45284 a_33249_35053.n113 a_33249_35053.n112 2.573
R45285 a_33249_35053.n117 a_33249_35053.n116 2.573
R45286 a_33249_35053.n138 a_33249_35053.n136 2.56118
R45287 a_33249_35053.n153 a_33249_35053.n151 2.56118
R45288 a_33249_35053.n131 a_33249_35053.n130 2.54573
R45289 a_33249_35053.n67 a_33249_35053.n65 2.53418
R45290 a_33249_35053.n50 a_33249_35053.n48 2.53418
R45291 a_33249_35053.n99 a_33249_35053.n97 2.53418
R45292 a_33249_35053.n29 a_33249_35053.n27 2.53418
R45293 a_33249_35053.n75 a_33249_35053.n15 2.51873
R45294 a_33249_35053.n45 a_33249_35053.n43 2.40765
R45295 a_33249_35053.n54 a_33249_35053.n52 2.40765
R45296 a_33249_35053.n62 a_33249_35053.n60 2.40765
R45297 a_33249_35053.n40 a_33249_35053.n38 2.40765
R45298 a_33249_35053.n24 a_33249_35053.n22 2.40765
R45299 a_33249_35053.n86 a_33249_35053.n84 2.40765
R45300 a_33249_35053.n94 a_33249_35053.n92 2.40765
R45301 a_33249_35053.n19 a_33249_35053.n17 2.40765
R45302 a_33249_35053.n156 a_33249_35053.n155 2.27857
R45303 a_33249_35053.n33 a_33249_35053.n30 2.23844
R45304 a_33249_35053.n134 a_33249_35053.n13 2.00466
R45305 a_33249_35053.n121 a_33249_35053.n120 1.67718
R45306 a_33249_35053.n0 a_33249_35053.n156 1.67353
R45307 a_33249_35053.n73 a_33249_35053.n6 1.65553
R45308 a_33249_35053.n104 a_33249_35053.n3 1.65553
R45309 a_33249_35053.n101 a_33249_35053.n100 1.5005
R45310 a_33249_35053.n69 a_33249_35053.n68 1.5005
R45311 a_33249_35053.n104 a_33249_35053.n14 1.5005
R45312 a_33249_35053.n83 a_33249_35053.n82 1.5005
R45313 a_33249_35053.n81 a_33249_35053.n80 1.5005
R45314 a_33249_35053.n74 a_33249_35053.n73 1.5005
R45315 a_33249_35053.n51 a_33249_35053.n30 1.5005
R45316 a_33249_35053.n134 a_33249_35053.n133 1.5005
R45317 a_33249_35053.n155 a_33249_35053.n154 1.5005
R45318 a_33249_35053.n127 a_33249_35053.n10 1.5005
R45319 a_33249_35053.n103 a_33249_35053.t68 1.4705
R45320 a_33249_35053.n103 a_33249_35053.t10 1.4705
R45321 a_33249_35053.n102 a_33249_35053.t74 1.4705
R45322 a_33249_35053.n102 a_33249_35053.t18 1.4705
R45323 a_33249_35053.n31 a_33249_35053.t78 1.4705
R45324 a_33249_35053.n31 a_33249_35053.t29 1.4705
R45325 a_33249_35053.n34 a_33249_35053.t88 1.4705
R45326 a_33249_35053.n34 a_33249_35053.t46 1.4705
R45327 a_33249_35053.n43 a_33249_35053.t71 1.4705
R45328 a_33249_35053.n43 a_33249_35053.t14 1.4705
R45329 a_33249_35053.n44 a_33249_35053.t67 1.4705
R45330 a_33249_35053.n44 a_33249_35053.t9 1.4705
R45331 a_33249_35053.n52 a_33249_35053.t77 1.4705
R45332 a_33249_35053.n52 a_33249_35053.t23 1.4705
R45333 a_33249_35053.n53 a_33249_35053.t70 1.4705
R45334 a_33249_35053.n53 a_33249_35053.t12 1.4705
R45335 a_33249_35053.n60 a_33249_35053.t81 1.4705
R45336 a_33249_35053.n60 a_33249_35053.t11 1.4705
R45337 a_33249_35053.n61 a_33249_35053.t72 1.4705
R45338 a_33249_35053.n61 a_33249_35053.t6 1.4705
R45339 a_33249_35053.n38 a_33249_35053.t24 1.4705
R45340 a_33249_35053.n38 a_33249_35053.t50 1.4705
R45341 a_33249_35053.n39 a_33249_35053.t15 1.4705
R45342 a_33249_35053.n39 a_33249_35053.t40 1.4705
R45343 a_33249_35053.n72 a_33249_35053.t63 1.4705
R45344 a_33249_35053.n72 a_33249_35053.t1 1.4705
R45345 a_33249_35053.n71 a_33249_35053.t66 1.4705
R45346 a_33249_35053.n71 a_33249_35053.t7 1.4705
R45347 a_33249_35053.n78 a_33249_35053.t84 1.4705
R45348 a_33249_35053.n78 a_33249_35053.t31 1.4705
R45349 a_33249_35053.n76 a_33249_35053.t3 1.4705
R45350 a_33249_35053.n76 a_33249_35053.t54 1.4705
R45351 a_33249_35053.n22 a_33249_35053.t76 1.4705
R45352 a_33249_35053.n22 a_33249_35053.t22 1.4705
R45353 a_33249_35053.n23 a_33249_35053.t75 1.4705
R45354 a_33249_35053.n23 a_33249_35053.t20 1.4705
R45355 a_33249_35053.n84 a_33249_35053.t83 1.4705
R45356 a_33249_35053.n84 a_33249_35053.t27 1.4705
R45357 a_33249_35053.n85 a_33249_35053.t82 1.4705
R45358 a_33249_35053.n85 a_33249_35053.t25 1.4705
R45359 a_33249_35053.n92 a_33249_35053.t87 1.4705
R45360 a_33249_35053.n92 a_33249_35053.t17 1.4705
R45361 a_33249_35053.n93 a_33249_35053.t86 1.4705
R45362 a_33249_35053.n93 a_33249_35053.t16 1.4705
R45363 a_33249_35053.n17 a_33249_35053.t28 1.4705
R45364 a_33249_35053.n17 a_33249_35053.t57 1.4705
R45365 a_33249_35053.n18 a_33249_35053.t26 1.4705
R45366 a_33249_35053.n18 a_33249_35053.t55 1.4705
R45367 a_33249_35053.n151 a_33249_35053.n150 1.46537
R45368 a_33249_35053.n146 a_33249_35053.n145 1.46537
R45369 a_33249_35053.n142 a_33249_35053.n141 1.46537
R45370 a_33249_35053.n138 a_33249_35053.n137 1.46537
R45371 a_33249_35053.n46 a_33249_35053.n45 1.46537
R45372 a_33249_35053.n48 a_33249_35053.n47 1.46537
R45373 a_33249_35053.n55 a_33249_35053.n54 1.46537
R45374 a_33249_35053.n57 a_33249_35053.n56 1.46537
R45375 a_33249_35053.n59 a_33249_35053.n58 1.46537
R45376 a_33249_35053.n63 a_33249_35053.n62 1.46537
R45377 a_33249_35053.n65 a_33249_35053.n64 1.46537
R45378 a_33249_35053.n41 a_33249_35053.n40 1.46537
R45379 a_33249_35053.n25 a_33249_35053.n24 1.46537
R45380 a_33249_35053.n27 a_33249_35053.n26 1.46537
R45381 a_33249_35053.n87 a_33249_35053.n86 1.46537
R45382 a_33249_35053.n89 a_33249_35053.n88 1.46537
R45383 a_33249_35053.n91 a_33249_35053.n90 1.46537
R45384 a_33249_35053.n95 a_33249_35053.n94 1.46537
R45385 a_33249_35053.n97 a_33249_35053.n96 1.46537
R45386 a_33249_35053.n20 a_33249_35053.n19 1.46537
R45387 a_33249_35053.n114 a_33249_35053.n113 1.46537
R45388 a_33249_35053.n118 a_33249_35053.n117 1.46537
R45389 a_33249_35053.n120 a_33249_35053.n119 1.46537
R45390 a_33249_35053.n153 a_33249_35053.n152 1.46535
R45391 a_33249_35053.n136 a_33249_35053.n135 1.46535
R45392 a_33249_35053.n50 a_33249_35053.n49 1.46535
R45393 a_33249_35053.n67 a_33249_35053.n66 1.46535
R45394 a_33249_35053.n29 a_33249_35053.n28 1.46535
R45395 a_33249_35053.n99 a_33249_35053.n98 1.46535
R45396 a_33249_35053.n106 a_33249_35053.n105 1.43535
R45397 a_33249_35053.n124 a_33249_35053.n123 1.31908
R45398 a_33249_35053.n36 a_33249_35053.n35 1.27228
R45399 a_33249_35053.n65 a_33249_35053.n63 1.27228
R45400 a_33249_35053.n63 a_33249_35053.n59 1.27228
R45401 a_33249_35053.n57 a_33249_35053.n55 1.27228
R45402 a_33249_35053.n48 a_33249_35053.n46 1.27228
R45403 a_33249_35053.n77 a_33249_35053.n75 1.27228
R45404 a_33249_35053.n97 a_33249_35053.n95 1.27228
R45405 a_33249_35053.n95 a_33249_35053.n91 1.27228
R45406 a_33249_35053.n89 a_33249_35053.n87 1.27228
R45407 a_33249_35053.n27 a_33249_35053.n25 1.27228
R45408 a_33249_35053.n157 a_33249_35053.t127 1.2605
R45409 a_33249_35053.n157 a_33249_35053.t125 1.2605
R45410 a_33249_35053.n132 a_33249_35053.t113 1.2605
R45411 a_33249_35053.n132 a_33249_35053.t111 1.2605
R45412 a_33249_35053.n147 a_33249_35053.t118 1.2605
R45413 a_33249_35053.n147 a_33249_35053.t136 1.2605
R45414 a_33249_35053.n148 a_33249_35053.t112 1.2605
R45415 a_33249_35053.n148 a_33249_35053.t132 1.2605
R45416 a_33249_35053.n143 a_33249_35053.t121 1.2605
R45417 a_33249_35053.n143 a_33249_35053.t133 1.2605
R45418 a_33249_35053.n144 a_33249_35053.t116 1.2605
R45419 a_33249_35053.n144 a_33249_35053.t131 1.2605
R45420 a_33249_35053.n139 a_33249_35053.t138 1.2605
R45421 a_33249_35053.n139 a_33249_35053.t110 1.2605
R45422 a_33249_35053.n140 a_33249_35053.t135 1.2605
R45423 a_33249_35053.n140 a_33249_35053.t108 1.2605
R45424 a_33249_35053.n11 a_33249_35053.t109 1.2605
R45425 a_33249_35053.n11 a_33249_35053.t122 1.2605
R45426 a_33249_35053.n12 a_33249_35053.t107 1.2605
R45427 a_33249_35053.n12 a_33249_35053.t119 1.2605
R45428 a_33249_35053.n111 a_33249_35053.t100 1.2605
R45429 a_33249_35053.n111 a_33249_35053.t97 1.2605
R45430 a_33249_35053.n112 a_33249_35053.t98 1.2605
R45431 a_33249_35053.n112 a_33249_35053.t93 1.2605
R45432 a_33249_35053.n115 a_33249_35053.t101 1.2605
R45433 a_33249_35053.n115 a_33249_35053.t104 1.2605
R45434 a_33249_35053.n116 a_33249_35053.t90 1.2605
R45435 a_33249_35053.n116 a_33249_35053.t94 1.2605
R45436 a_33249_35053.n107 a_33249_35053.t89 1.2605
R45437 a_33249_35053.n107 a_33249_35053.t95 1.2605
R45438 a_33249_35053.n122 a_33249_35053.t99 1.2605
R45439 a_33249_35053.n122 a_33249_35053.t102 1.2605
R45440 a_33249_35053.n125 a_33249_35053.t128 1.2605
R45441 a_33249_35053.n125 a_33249_35053.t141 1.2605
R45442 a_33249_35053.n128 a_33249_35053.t114 1.2605
R45443 a_33249_35053.n128 a_33249_35053.t129 1.2605
R45444 a_33249_35053.n130 a_33249_35053.n129 1.25428
R45445 a_33249_35053.n142 a_33249_35053.n138 1.25428
R45446 a_33249_35053.n120 a_33249_35053.n118 1.25428
R45447 a_33249_35053.n127 a_33249_35053.n126 1.04573
R45448 a_33249_35053.n33 a_33249_35053.n32 1.01873
R45449 a_33249_35053.n80 a_33249_35053.n79 1.01873
R45450 a_33249_35053.n70 a_33249_35053.n69 0.778574
R45451 a_33249_35053.n105 a_33249_35053.n101 0.778574
R45452 a_33249_35053.n74 a_33249_35053.n30 0.778574
R45453 a_33249_35053.n82 a_33249_35053.n14 0.778574
R45454 a_33249_35053.n101 a_33249_35053.n15 0.738439
R45455 a_33249_35053.n82 a_33249_35053.n81 0.738439
R45456 a_33249_35053.n133 a_33249_35053.n131 0.738439
R45457 a_33249_35053.n155 a_33249_35053.n10 0.738439
R45458 a_33249_35053.n121 a_33249_35053.n109 0.737223
R45459 a_33249_35053.n68 a_33249_35053.n67 0.699581
R45460 a_33249_35053.n51 a_33249_35053.n50 0.699581
R45461 a_33249_35053.n100 a_33249_35053.n99 0.699581
R45462 a_33249_35053.n83 a_33249_35053.n29 0.699581
R45463 a_33249_35053.n136 a_33249_35053.n134 0.699581
R45464 a_33249_35053.n154 a_33249_35053.n153 0.699581
R45465 a_33249_35053.n123 a_33249_35053.n121 0.585196
R45466 a_33249_35053.n68 a_33249_35053.n41 0.557791
R45467 a_33249_35053.n55 a_33249_35053.n51 0.557791
R45468 a_33249_35053.n100 a_33249_35053.n20 0.557791
R45469 a_33249_35053.n87 a_33249_35053.n83 0.557791
R45470 a_33249_35053.n154 a_33249_35053.n146 0.539791
R45471 a_33249_35053.n70 a_33249_35053.n15 0.530466
R45472 a_33249_35053.n81 a_33249_35053.n74 0.530466
R45473 a_33249_35053.n7 a_33249_35053.n8 1.27228
R45474 a_33249_35053.n73 a_33249_35053.n7 7.30549
R45475 a_33249_35053.t35 a_33249_35053.n6 6.96214
R45476 a_33249_35053.n4 a_33249_35053.n5 1.27228
R45477 a_33249_35053.n104 a_33249_35053.n4 7.30549
R45478 a_33249_35053.t45 a_33249_35053.n3 6.96214
R45479 a_33249_35053.n122 a_33249_35053.n9 5.45652
R45480 a_33249_35053.n1 a_33249_35053.n2 1.25428
R45481 a_33249_35053.n1 a_33249_35053.n156 5.95549
R45482 a_33249_35053.t140 a_33249_35053.n0 7.10317
R45483 a_31953_n19727.n226 a_31953_n19727.n321 15.3954
R45484 a_31953_n19727.n321 a_31953_n19727.t72 13.6649
R45485 a_31953_n19727.n233 a_31953_n19727.t99 10.1674
R45486 a_31953_n19727.t174 a_31953_n19727.n238 10.1674
R45487 a_31953_n19727.n239 a_31953_n19727.t174 10.1674
R45488 a_31953_n19727.t159 a_31953_n19727.n242 10.1674
R45489 a_31953_n19727.n243 a_31953_n19727.t159 10.1674
R45490 a_31953_n19727.n255 a_31953_n19727.t238 10.1674
R45491 a_31953_n19727.t238 a_31953_n19727.n254 10.1674
R45492 a_31953_n19727.n251 a_31953_n19727.t311 10.1674
R45493 a_31953_n19727.t311 a_31953_n19727.n250 10.1674
R45494 a_31953_n19727.n247 a_31953_n19727.t299 10.1674
R45495 a_31953_n19727.t299 a_31953_n19727.n246 10.1674
R45496 a_31953_n19727.t78 a_31953_n19727.n263 10.1674
R45497 a_31953_n19727.n264 a_31953_n19727.t78 10.1674
R45498 a_31953_n19727.t146 a_31953_n19727.n267 10.1674
R45499 a_31953_n19727.n268 a_31953_n19727.t146 10.1674
R45500 a_31953_n19727.t128 a_31953_n19727.n271 10.1674
R45501 a_31953_n19727.n272 a_31953_n19727.t128 10.1674
R45502 a_31953_n19727.n466 a_31953_n19727.t246 10.1674
R45503 a_31953_n19727.t317 a_31953_n19727.n471 10.1674
R45504 a_31953_n19727.n472 a_31953_n19727.t317 10.1674
R45505 a_31953_n19727.t98 a_31953_n19727.n475 10.1674
R45506 a_31953_n19727.n476 a_31953_n19727.t98 10.1674
R45507 a_31953_n19727.t86 a_31953_n19727.n483 10.1674
R45508 a_31953_n19727.n484 a_31953_n19727.t86 10.1674
R45509 a_31953_n19727.t158 a_31953_n19727.n487 10.1674
R45510 a_31953_n19727.n488 a_31953_n19727.t158 10.1674
R45511 a_31953_n19727.t222 a_31953_n19727.n491 10.1674
R45512 a_31953_n19727.n492 a_31953_n19727.t222 10.1674
R45513 a_31953_n19727.n505 a_31953_n19727.t296 10.1674
R45514 a_31953_n19727.t296 a_31953_n19727.n504 10.1674
R45515 a_31953_n19727.n501 a_31953_n19727.t354 10.1674
R45516 a_31953_n19727.t354 a_31953_n19727.n500 10.1674
R45517 a_31953_n19727.n499 a_31953_n19727.t137 10.1674
R45518 a_31953_n19727.t137 a_31953_n19727.n498 10.1674
R45519 a_31953_n19727.n279 a_31953_n19727.t180 10.1674
R45520 a_31953_n19727.t255 a_31953_n19727.n284 10.1674
R45521 a_31953_n19727.n285 a_31953_n19727.t255 10.1674
R45522 a_31953_n19727.t240 a_31953_n19727.n288 10.1674
R45523 a_31953_n19727.n289 a_31953_n19727.t240 10.1674
R45524 a_31953_n19727.n301 a_31953_n19727.t312 10.1674
R45525 a_31953_n19727.t312 a_31953_n19727.n300 10.1674
R45526 a_31953_n19727.n297 a_31953_n19727.t91 10.1674
R45527 a_31953_n19727.t91 a_31953_n19727.n296 10.1674
R45528 a_31953_n19727.n293 a_31953_n19727.t81 10.1674
R45529 a_31953_n19727.t81 a_31953_n19727.n292 10.1674
R45530 a_31953_n19727.t151 a_31953_n19727.n309 10.1674
R45531 a_31953_n19727.n310 a_31953_n19727.t151 10.1674
R45532 a_31953_n19727.t231 a_31953_n19727.n313 10.1674
R45533 a_31953_n19727.n314 a_31953_n19727.t231 10.1674
R45534 a_31953_n19727.t210 a_31953_n19727.n317 10.1674
R45535 a_31953_n19727.n318 a_31953_n19727.t210 10.1674
R45536 a_31953_n19727.n364 a_31953_n19727.t126 10.1674
R45537 a_31953_n19727.n360 a_31953_n19727.t203 10.1674
R45538 a_31953_n19727.t203 a_31953_n19727.n359 10.1674
R45539 a_31953_n19727.n356 a_31953_n19727.t279 10.1674
R45540 a_31953_n19727.t279 a_31953_n19727.n355 10.1674
R45541 a_31953_n19727.t266 a_31953_n19727.n325 10.1674
R45542 a_31953_n19727.n326 a_31953_n19727.t266 10.1674
R45543 a_31953_n19727.t336 a_31953_n19727.n329 10.1674
R45544 a_31953_n19727.n330 a_31953_n19727.t336 10.1674
R45545 a_31953_n19727.t103 a_31953_n19727.n333 10.1674
R45546 a_31953_n19727.n334 a_31953_n19727.t103 10.1674
R45547 a_31953_n19727.n347 a_31953_n19727.t179 10.1674
R45548 a_31953_n19727.t179 a_31953_n19727.n346 10.1674
R45549 a_31953_n19727.n343 a_31953_n19727.t235 10.1674
R45550 a_31953_n19727.t235 a_31953_n19727.n342 10.1674
R45551 a_31953_n19727.n341 a_31953_n19727.t309 10.1674
R45552 a_31953_n19727.t309 a_31953_n19727.n340 10.1674
R45553 a_31953_n19727.n373 a_31953_n19727.t293 10.1674
R45554 a_31953_n19727.t74 a_31953_n19727.n378 10.1674
R45555 a_31953_n19727.n379 a_31953_n19727.t74 10.1674
R45556 a_31953_n19727.t356 a_31953_n19727.n382 10.1674
R45557 a_31953_n19727.n383 a_31953_n19727.t356 10.1674
R45558 a_31953_n19727.n395 a_31953_n19727.t138 10.1674
R45559 a_31953_n19727.t138 a_31953_n19727.n394 10.1674
R45560 a_31953_n19727.n391 a_31953_n19727.t215 10.1674
R45561 a_31953_n19727.t215 a_31953_n19727.n390 10.1674
R45562 a_31953_n19727.n387 a_31953_n19727.t200 10.1674
R45563 a_31953_n19727.t200 a_31953_n19727.n386 10.1674
R45564 a_31953_n19727.t278 a_31953_n19727.n403 10.1674
R45565 a_31953_n19727.n404 a_31953_n19727.t278 10.1674
R45566 a_31953_n19727.t351 a_31953_n19727.n407 10.1674
R45567 a_31953_n19727.n408 a_31953_n19727.t351 10.1674
R45568 a_31953_n19727.t318 a_31953_n19727.n411 10.1674
R45569 a_31953_n19727.n412 a_31953_n19727.t318 10.1674
R45570 a_31953_n19727.n457 a_31953_n19727.t90 10.1674
R45571 a_31953_n19727.n453 a_31953_n19727.t166 10.1674
R45572 a_31953_n19727.t166 a_31953_n19727.n452 10.1674
R45573 a_31953_n19727.n449 a_31953_n19727.t245 10.1674
R45574 a_31953_n19727.t245 a_31953_n19727.n448 10.1674
R45575 a_31953_n19727.t230 a_31953_n19727.n418 10.1674
R45576 a_31953_n19727.n419 a_31953_n19727.t230 10.1674
R45577 a_31953_n19727.t304 a_31953_n19727.n422 10.1674
R45578 a_31953_n19727.n423 a_31953_n19727.t304 10.1674
R45579 a_31953_n19727.t360 a_31953_n19727.n426 10.1674
R45580 a_31953_n19727.n427 a_31953_n19727.t360 10.1674
R45581 a_31953_n19727.n440 a_31953_n19727.t142 10.1674
R45582 a_31953_n19727.t142 a_31953_n19727.n439 10.1674
R45583 a_31953_n19727.n436 a_31953_n19727.t209 10.1674
R45584 a_31953_n19727.t209 a_31953_n19727.n435 10.1674
R45585 a_31953_n19727.n434 a_31953_n19727.t282 10.1674
R45586 a_31953_n19727.t282 a_31953_n19727.n433 10.1674
R45587 a_31953_n19727.n235 a_31953_n19727.t197 10.1674
R45588 a_31953_n19727.t276 a_31953_n19727.n240 10.1674
R45589 a_31953_n19727.n241 a_31953_n19727.t276 10.1674
R45590 a_31953_n19727.t262 a_31953_n19727.n244 10.1674
R45591 a_31953_n19727.n245 a_31953_n19727.t262 10.1674
R45592 a_31953_n19727.n257 a_31953_n19727.t333 10.1674
R45593 a_31953_n19727.t333 a_31953_n19727.n256 10.1674
R45594 a_31953_n19727.n253 a_31953_n19727.t117 10.1674
R45595 a_31953_n19727.t117 a_31953_n19727.n252 10.1674
R45596 a_31953_n19727.n249 a_31953_n19727.t102 10.1674
R45597 a_31953_n19727.t102 a_31953_n19727.n248 10.1674
R45598 a_31953_n19727.t177 a_31953_n19727.n265 10.1674
R45599 a_31953_n19727.n266 a_31953_n19727.t177 10.1674
R45600 a_31953_n19727.t253 a_31953_n19727.n269 10.1674
R45601 a_31953_n19727.n270 a_31953_n19727.t253 10.1674
R45602 a_31953_n19727.t224 a_31953_n19727.n273 10.1674
R45603 a_31953_n19727.n274 a_31953_n19727.t224 10.1674
R45604 a_31953_n19727.n468 a_31953_n19727.t290 10.1674
R45605 a_31953_n19727.t361 a_31953_n19727.n473 10.1674
R45606 a_31953_n19727.n474 a_31953_n19727.t361 10.1674
R45607 a_31953_n19727.t143 a_31953_n19727.n477 10.1674
R45608 a_31953_n19727.n478 a_31953_n19727.t143 10.1674
R45609 a_31953_n19727.t135 a_31953_n19727.n485 10.1674
R45610 a_31953_n19727.n486 a_31953_n19727.t135 10.1674
R45611 a_31953_n19727.t214 a_31953_n19727.n489 10.1674
R45612 a_31953_n19727.n490 a_31953_n19727.t214 10.1674
R45613 a_31953_n19727.t274 a_31953_n19727.n493 10.1674
R45614 a_31953_n19727.n494 a_31953_n19727.t274 10.1674
R45615 a_31953_n19727.n507 a_31953_n19727.t346 10.1674
R45616 a_31953_n19727.t346 a_31953_n19727.n506 10.1674
R45617 a_31953_n19727.n503 a_31953_n19727.t110 10.1674
R45618 a_31953_n19727.t110 a_31953_n19727.n502 10.1674
R45619 a_31953_n19727.t184 a_31953_n19727.n496 10.1674
R45620 a_31953_n19727.n497 a_31953_n19727.t184 10.1674
R45621 a_31953_n19727.n281 a_31953_n19727.t114 10.1674
R45622 a_31953_n19727.t189 a_31953_n19727.n286 10.1674
R45623 a_31953_n19727.n287 a_31953_n19727.t189 10.1674
R45624 a_31953_n19727.t172 a_31953_n19727.n290 10.1674
R45625 a_31953_n19727.n291 a_31953_n19727.t172 10.1674
R45626 a_31953_n19727.n303 a_31953_n19727.t251 10.1674
R45627 a_31953_n19727.t251 a_31953_n19727.n302 10.1674
R45628 a_31953_n19727.n299 a_31953_n19727.t320 10.1674
R45629 a_31953_n19727.t320 a_31953_n19727.n298 10.1674
R45630 a_31953_n19727.n295 a_31953_n19727.t310 10.1674
R45631 a_31953_n19727.t310 a_31953_n19727.n294 10.1674
R45632 a_31953_n19727.t89 a_31953_n19727.n311 10.1674
R45633 a_31953_n19727.n312 a_31953_n19727.t89 10.1674
R45634 a_31953_n19727.t164 a_31953_n19727.n315 10.1674
R45635 a_31953_n19727.n316 a_31953_n19727.t164 10.1674
R45636 a_31953_n19727.t139 a_31953_n19727.n319 10.1674
R45637 a_31953_n19727.n320 a_31953_n19727.t139 10.1674
R45638 a_31953_n19727.n366 a_31953_n19727.t305 10.1674
R45639 a_31953_n19727.n362 a_31953_n19727.t87 10.1674
R45640 a_31953_n19727.t87 a_31953_n19727.n361 10.1674
R45641 a_31953_n19727.n358 a_31953_n19727.t161 10.1674
R45642 a_31953_n19727.t161 a_31953_n19727.n357 10.1674
R45643 a_31953_n19727.t145 a_31953_n19727.n327 10.1674
R45644 a_31953_n19727.n328 a_31953_n19727.t145 10.1674
R45645 a_31953_n19727.t226 a_31953_n19727.n331 10.1674
R45646 a_31953_n19727.n332 a_31953_n19727.t226 10.1674
R45647 a_31953_n19727.t288 a_31953_n19727.n335 10.1674
R45648 a_31953_n19727.n336 a_31953_n19727.t288 10.1674
R45649 a_31953_n19727.n349 a_31953_n19727.t359 10.1674
R45650 a_31953_n19727.t359 a_31953_n19727.n348 10.1674
R45651 a_31953_n19727.n345 a_31953_n19727.t125 10.1674
R45652 a_31953_n19727.t125 a_31953_n19727.n344 10.1674
R45653 a_31953_n19727.t202 a_31953_n19727.n338 10.1674
R45654 a_31953_n19727.n339 a_31953_n19727.t202 10.1674
R45655 a_31953_n19727.n375 a_31953_n19727.t258 10.1674
R45656 a_31953_n19727.t326 a_31953_n19727.n380 10.1674
R45657 a_31953_n19727.n381 a_31953_n19727.t326 10.1674
R45658 a_31953_n19727.t314 a_31953_n19727.n384 10.1674
R45659 a_31953_n19727.n385 a_31953_n19727.t314 10.1674
R45660 a_31953_n19727.n397 a_31953_n19727.t94 10.1674
R45661 a_31953_n19727.t94 a_31953_n19727.n396 10.1674
R45662 a_31953_n19727.n393 a_31953_n19727.t168 10.1674
R45663 a_31953_n19727.t168 a_31953_n19727.n392 10.1674
R45664 a_31953_n19727.n389 a_31953_n19727.t155 10.1674
R45665 a_31953_n19727.t155 a_31953_n19727.n388 10.1674
R45666 a_31953_n19727.t234 a_31953_n19727.n405 10.1674
R45667 a_31953_n19727.n406 a_31953_n19727.t234 10.1674
R45668 a_31953_n19727.t308 a_31953_n19727.n409 10.1674
R45669 a_31953_n19727.n410 a_31953_n19727.t308 10.1674
R45670 a_31953_n19727.t285 a_31953_n19727.n413 10.1674
R45671 a_31953_n19727.n414 a_31953_n19727.t285 10.1674
R45672 a_31953_n19727.n459 a_31953_n19727.t193 10.1674
R45673 a_31953_n19727.n455 a_31953_n19727.t268 10.1674
R45674 a_31953_n19727.t268 a_31953_n19727.n454 10.1674
R45675 a_31953_n19727.n451 a_31953_n19727.t340 10.1674
R45676 a_31953_n19727.t340 a_31953_n19727.n450 10.1674
R45677 a_31953_n19727.t323 a_31953_n19727.n420 10.1674
R45678 a_31953_n19727.n421 a_31953_n19727.t323 10.1674
R45679 a_31953_n19727.t108 a_31953_n19727.n424 10.1674
R45680 a_31953_n19727.n425 a_31953_n19727.t108 10.1674
R45681 a_31953_n19727.t165 a_31953_n19727.n428 10.1674
R45682 a_31953_n19727.n429 a_31953_n19727.t165 10.1674
R45683 a_31953_n19727.n442 a_31953_n19727.t244 10.1674
R45684 a_31953_n19727.t244 a_31953_n19727.n441 10.1674
R45685 a_31953_n19727.n438 a_31953_n19727.t300 10.1674
R45686 a_31953_n19727.t300 a_31953_n19727.n437 10.1674
R45687 a_31953_n19727.t80 a_31953_n19727.n431 10.1674
R45688 a_31953_n19727.n432 a_31953_n19727.t80 10.1674
R45689 a_31953_n19727.t99 a_31953_n19727.n232 10.1409
R45690 a_31953_n19727.t246 a_31953_n19727.n465 10.1409
R45691 a_31953_n19727.t180 a_31953_n19727.n278 10.1409
R45692 a_31953_n19727.t126 a_31953_n19727.n363 10.1409
R45693 a_31953_n19727.t293 a_31953_n19727.n372 10.1409
R45694 a_31953_n19727.t90 a_31953_n19727.n456 10.1409
R45695 a_31953_n19727.t197 a_31953_n19727.n234 10.1409
R45696 a_31953_n19727.t290 a_31953_n19727.n467 10.1409
R45697 a_31953_n19727.t114 a_31953_n19727.n280 10.1409
R45698 a_31953_n19727.t305 a_31953_n19727.n365 10.1409
R45699 a_31953_n19727.t258 a_31953_n19727.n374 10.1409
R45700 a_31953_n19727.t193 a_31953_n19727.n458 10.1409
R45701 a_31953_n19727.t195 a_31953_n19727.n232 9.54631
R45702 a_31953_n19727.n214 a_31953_n19727.t273 9.54631
R45703 a_31953_n19727.t100 a_31953_n19727.n213 9.54631
R45704 a_31953_n19727.n234 a_31953_n19727.t208 9.54631
R45705 a_31953_n19727.t141 a_31953_n19727.n465 9.54631
R45706 a_31953_n19727.n216 a_31953_n19727.t330 9.54631
R45707 a_31953_n19727.t104 a_31953_n19727.n215 9.54631
R45708 a_31953_n19727.n467 a_31953_n19727.t358 9.54631
R45709 a_31953_n19727.t275 a_31953_n19727.n278 9.54631
R45710 a_31953_n19727.n218 a_31953_n19727.t187 9.54631
R45711 a_31953_n19727.t181 a_31953_n19727.n217 9.54631
R45712 a_31953_n19727.n280 a_31953_n19727.t286 9.54631
R45713 a_31953_n19727.t315 a_31953_n19727.n363 9.54631
R45714 a_31953_n19727.n220 a_31953_n19727.t350 9.54631
R45715 a_31953_n19727.t283 a_31953_n19727.n219 9.54631
R45716 a_31953_n19727.n365 a_31953_n19727.t243 9.54631
R45717 a_31953_n19727.t316 a_31953_n19727.n372 9.54631
R45718 a_31953_n19727.n222 a_31953_n19727.t130 9.54631
R45719 a_31953_n19727.t348 a_31953_n19727.n221 9.54631
R45720 a_31953_n19727.n374 a_31953_n19727.t132 9.54631
R45721 a_31953_n19727.t196 a_31953_n19727.n456 9.54631
R45722 a_31953_n19727.n224 a_31953_n19727.t148 9.54631
R45723 a_31953_n19727.t227 a_31953_n19727.n223 9.54631
R45724 a_31953_n19727.n458 a_31953_n19727.t123 9.54631
R45725 a_31953_n19727.n233 a_31953_n19727.t195 9.54355
R45726 a_31953_n19727.t273 a_31953_n19727.n237 9.54355
R45727 a_31953_n19727.n236 a_31953_n19727.t100 9.54355
R45728 a_31953_n19727.n235 a_31953_n19727.t208 9.54355
R45729 a_31953_n19727.n239 a_31953_n19727.t271 9.54355
R45730 a_31953_n19727.t271 a_31953_n19727.n238 9.54355
R45731 a_31953_n19727.t345 a_31953_n19727.n4 9.54355
R45732 a_31953_n19727.n1 a_31953_n19727.t345 9.54355
R45733 a_31953_n19727.n2 a_31953_n19727.t175 9.54355
R45734 a_31953_n19727.t175 a_31953_n19727.n0 9.54355
R45735 a_31953_n19727.n241 a_31953_n19727.t281 9.54355
R45736 a_31953_n19727.n240 a_31953_n19727.t281 9.54355
R45737 a_31953_n19727.n243 a_31953_n19727.t259 9.54355
R45738 a_31953_n19727.t259 a_31953_n19727.n242 9.54355
R45739 a_31953_n19727.t329 a_31953_n19727.n8 9.54355
R45740 a_31953_n19727.n6 a_31953_n19727.t329 9.54355
R45741 a_31953_n19727.n7 a_31953_n19727.t160 9.54355
R45742 a_31953_n19727.t160 a_31953_n19727.n5 9.54355
R45743 a_31953_n19727.n245 a_31953_n19727.t270 9.54355
R45744 a_31953_n19727.n244 a_31953_n19727.t270 9.54355
R45745 a_31953_n19727.t327 a_31953_n19727.n254 9.54355
R45746 a_31953_n19727.n255 a_31953_n19727.t327 9.54355
R45747 a_31953_n19727.n13 a_31953_n19727.t60 9.54355
R45748 a_31953_n19727.t60 a_31953_n19727.n11 9.54355
R45749 a_31953_n19727.t38 a_31953_n19727.n12 9.54355
R45750 a_31953_n19727.n9 a_31953_n19727.t38 9.54355
R45751 a_31953_n19727.n256 a_31953_n19727.t342 9.54355
R45752 a_31953_n19727.n257 a_31953_n19727.t342 9.54355
R45753 a_31953_n19727.t112 a_31953_n19727.n250 9.54355
R45754 a_31953_n19727.n251 a_31953_n19727.t112 9.54355
R45755 a_31953_n19727.n17 a_31953_n19727.t48 9.54355
R45756 a_31953_n19727.t48 a_31953_n19727.n15 9.54355
R45757 a_31953_n19727.t16 a_31953_n19727.n16 9.54355
R45758 a_31953_n19727.n14 a_31953_n19727.t16 9.54355
R45759 a_31953_n19727.n252 a_31953_n19727.t121 9.54355
R45760 a_31953_n19727.n253 a_31953_n19727.t121 9.54355
R45761 a_31953_n19727.t95 a_31953_n19727.n246 9.54355
R45762 a_31953_n19727.n247 a_31953_n19727.t95 9.54355
R45763 a_31953_n19727.n22 a_31953_n19727.t52 9.54355
R45764 a_31953_n19727.t52 a_31953_n19727.n20 9.54355
R45765 a_31953_n19727.t20 a_31953_n19727.n21 9.54355
R45766 a_31953_n19727.n18 a_31953_n19727.t20 9.54355
R45767 a_31953_n19727.n248 a_31953_n19727.t111 9.54355
R45768 a_31953_n19727.n249 a_31953_n19727.t111 9.54355
R45769 a_31953_n19727.n264 a_31953_n19727.t170 9.54355
R45770 a_31953_n19727.t170 a_31953_n19727.n263 9.54355
R45771 a_31953_n19727.t250 a_31953_n19727.n26 9.54355
R45772 a_31953_n19727.n24 a_31953_n19727.t250 9.54355
R45773 a_31953_n19727.n25 a_31953_n19727.t79 9.54355
R45774 a_31953_n19727.t79 a_31953_n19727.n23 9.54355
R45775 a_31953_n19727.n266 a_31953_n19727.t186 9.54355
R45776 a_31953_n19727.n265 a_31953_n19727.t186 9.54355
R45777 a_31953_n19727.n268 a_31953_n19727.t248 9.54355
R45778 a_31953_n19727.t248 a_31953_n19727.n267 9.54355
R45779 a_31953_n19727.t319 a_31953_n19727.n31 9.54355
R45780 a_31953_n19727.n28 a_31953_n19727.t319 9.54355
R45781 a_31953_n19727.n29 a_31953_n19727.t149 9.54355
R45782 a_31953_n19727.t149 a_31953_n19727.n27 9.54355
R45783 a_31953_n19727.n270 a_31953_n19727.t261 9.54355
R45784 a_31953_n19727.n269 a_31953_n19727.t261 9.54355
R45785 a_31953_n19727.n272 a_31953_n19727.t221 9.54355
R45786 a_31953_n19727.t221 a_31953_n19727.n271 9.54355
R45787 a_31953_n19727.t295 a_31953_n19727.n35 9.54355
R45788 a_31953_n19727.n33 a_31953_n19727.t295 9.54355
R45789 a_31953_n19727.n34 a_31953_n19727.t129 9.54355
R45790 a_31953_n19727.t129 a_31953_n19727.n32 9.54355
R45791 a_31953_n19727.n274 a_31953_n19727.t229 9.54355
R45792 a_31953_n19727.n273 a_31953_n19727.t229 9.54355
R45793 a_31953_n19727.n466 a_31953_n19727.t141 9.54355
R45794 a_31953_n19727.t330 a_31953_n19727.n470 9.54355
R45795 a_31953_n19727.n469 a_31953_n19727.t104 9.54355
R45796 a_31953_n19727.n468 a_31953_n19727.t358 9.54355
R45797 a_31953_n19727.n472 a_31953_n19727.t220 9.54355
R45798 a_31953_n19727.t220 a_31953_n19727.n471 9.54355
R45799 a_31953_n19727.t115 a_31953_n19727.n40 9.54355
R45800 a_31953_n19727.n37 a_31953_n19727.t115 9.54355
R45801 a_31953_n19727.n38 a_31953_n19727.t182 9.54355
R45802 a_31953_n19727.t182 a_31953_n19727.n36 9.54355
R45803 a_31953_n19727.n474 a_31953_n19727.t140 9.54355
R45804 a_31953_n19727.n473 a_31953_n19727.t140 9.54355
R45805 a_31953_n19727.n476 a_31953_n19727.t292 9.54355
R45806 a_31953_n19727.t292 a_31953_n19727.n475 9.54355
R45807 a_31953_n19727.t190 a_31953_n19727.n44 9.54355
R45808 a_31953_n19727.n42 a_31953_n19727.t190 9.54355
R45809 a_31953_n19727.n43 a_31953_n19727.t260 9.54355
R45810 a_31953_n19727.t260 a_31953_n19727.n41 9.54355
R45811 a_31953_n19727.n478 a_31953_n19727.t217 9.54355
R45812 a_31953_n19727.n477 a_31953_n19727.t217 9.54355
R45813 a_31953_n19727.n484 a_31953_n19727.t284 9.54355
R45814 a_31953_n19727.t284 a_31953_n19727.n483 9.54355
R45815 a_31953_n19727.t50 a_31953_n19727.n49 9.54355
R45816 a_31953_n19727.n46 a_31953_n19727.t50 9.54355
R45817 a_31953_n19727.n47 a_31953_n19727.t36 9.54355
R45818 a_31953_n19727.t36 a_31953_n19727.n45 9.54355
R45819 a_31953_n19727.n486 a_31953_n19727.t204 9.54355
R45820 a_31953_n19727.n485 a_31953_n19727.t204 9.54355
R45821 a_31953_n19727.n488 a_31953_n19727.t355 9.54355
R45822 a_31953_n19727.t355 a_31953_n19727.n487 9.54355
R45823 a_31953_n19727.t34 a_31953_n19727.n54 9.54355
R45824 a_31953_n19727.n51 a_31953_n19727.t34 9.54355
R45825 a_31953_n19727.n52 a_31953_n19727.t12 9.54355
R45826 a_31953_n19727.t12 a_31953_n19727.n50 9.54355
R45827 a_31953_n19727.n490 a_31953_n19727.t280 9.54355
R45828 a_31953_n19727.n489 a_31953_n19727.t280 9.54355
R45829 a_31953_n19727.n492 a_31953_n19727.t122 9.54355
R45830 a_31953_n19727.t122 a_31953_n19727.n491 9.54355
R45831 a_31953_n19727.t18 a_31953_n19727.n58 9.54355
R45832 a_31953_n19727.n56 a_31953_n19727.t18 9.54355
R45833 a_31953_n19727.n57 a_31953_n19727.t70 9.54355
R45834 a_31953_n19727.t70 a_31953_n19727.n55 9.54355
R45835 a_31953_n19727.n494 a_31953_n19727.t337 9.54355
R45836 a_31953_n19727.n493 a_31953_n19727.t337 9.54355
R45837 a_31953_n19727.t198 a_31953_n19727.n504 9.54355
R45838 a_31953_n19727.n505 a_31953_n19727.t198 9.54355
R45839 a_31953_n19727.n63 a_31953_n19727.t88 9.54355
R45840 a_31953_n19727.t88 a_31953_n19727.n61 9.54355
R45841 a_31953_n19727.t152 a_31953_n19727.n62 9.54355
R45842 a_31953_n19727.n59 a_31953_n19727.t152 9.54355
R45843 a_31953_n19727.n506 a_31953_n19727.t119 9.54355
R45844 a_31953_n19727.n507 a_31953_n19727.t119 9.54355
R45845 a_31953_n19727.t257 a_31953_n19727.n500 9.54355
R45846 a_31953_n19727.n501 a_31953_n19727.t257 9.54355
R45847 a_31953_n19727.n67 a_31953_n19727.t144 9.54355
R45848 a_31953_n19727.t144 a_31953_n19727.n65 9.54355
R45849 a_31953_n19727.t218 a_31953_n19727.n66 9.54355
R45850 a_31953_n19727.n64 a_31953_n19727.t218 9.54355
R45851 a_31953_n19727.n502 a_31953_n19727.t178 9.54355
R45852 a_31953_n19727.n503 a_31953_n19727.t178 9.54355
R45853 a_31953_n19727.t325 a_31953_n19727.n498 9.54355
R45854 a_31953_n19727.n499 a_31953_n19727.t325 9.54355
R45855 a_31953_n19727.n70 a_31953_n19727.t223 9.54355
R45856 a_31953_n19727.t223 a_31953_n19727.n68 9.54355
R45857 a_31953_n19727.n69 a_31953_n19727.t289 9.54355
R45858 a_31953_n19727.n495 a_31953_n19727.t289 9.54355
R45859 a_31953_n19727.n497 a_31953_n19727.t254 9.54355
R45860 a_31953_n19727.n496 a_31953_n19727.t254 9.54355
R45861 a_31953_n19727.n279 a_31953_n19727.t275 9.54355
R45862 a_31953_n19727.t187 a_31953_n19727.n283 9.54355
R45863 a_31953_n19727.n282 a_31953_n19727.t181 9.54355
R45864 a_31953_n19727.n281 a_31953_n19727.t286 9.54355
R45865 a_31953_n19727.n285 a_31953_n19727.t347 9.54355
R45866 a_31953_n19727.t347 a_31953_n19727.n284 9.54355
R45867 a_31953_n19727.t264 a_31953_n19727.n75 9.54355
R45868 a_31953_n19727.n72 a_31953_n19727.t264 9.54355
R45869 a_31953_n19727.n73 a_31953_n19727.t256 9.54355
R45870 a_31953_n19727.t256 a_31953_n19727.n71 9.54355
R45871 a_31953_n19727.n287 a_31953_n19727.t357 9.54355
R45872 a_31953_n19727.n286 a_31953_n19727.t357 9.54355
R45873 a_31953_n19727.n289 a_31953_n19727.t331 9.54355
R45874 a_31953_n19727.t331 a_31953_n19727.n288 9.54355
R45875 a_31953_n19727.t249 a_31953_n19727.n79 9.54355
R45876 a_31953_n19727.n77 a_31953_n19727.t249 9.54355
R45877 a_31953_n19727.n78 a_31953_n19727.t242 9.54355
R45878 a_31953_n19727.t242 a_31953_n19727.n76 9.54355
R45879 a_31953_n19727.n291 a_31953_n19727.t343 9.54355
R45880 a_31953_n19727.n290 a_31953_n19727.t343 9.54355
R45881 a_31953_n19727.t116 a_31953_n19727.n300 9.54355
R45882 a_31953_n19727.n301 a_31953_n19727.t116 9.54355
R45883 a_31953_n19727.n84 a_31953_n19727.t10 9.54355
R45884 a_31953_n19727.t10 a_31953_n19727.n82 9.54355
R45885 a_31953_n19727.t14 a_31953_n19727.n83 9.54355
R45886 a_31953_n19727.n80 a_31953_n19727.t14 9.54355
R45887 a_31953_n19727.n302 a_31953_n19727.t124 9.54355
R45888 a_31953_n19727.n303 a_31953_n19727.t124 9.54355
R45889 a_31953_n19727.t191 a_31953_n19727.n296 9.54355
R45890 a_31953_n19727.n297 a_31953_n19727.t191 9.54355
R45891 a_31953_n19727.n88 a_31953_n19727.t62 9.54355
R45892 a_31953_n19727.t62 a_31953_n19727.n86 9.54355
R45893 a_31953_n19727.t64 a_31953_n19727.n87 9.54355
R45894 a_31953_n19727.n85 a_31953_n19727.t64 9.54355
R45895 a_31953_n19727.n298 a_31953_n19727.t201 9.54355
R45896 a_31953_n19727.n299 a_31953_n19727.t201 9.54355
R45897 a_31953_n19727.t173 a_31953_n19727.n292 9.54355
R45898 a_31953_n19727.n293 a_31953_n19727.t173 9.54355
R45899 a_31953_n19727.n93 a_31953_n19727.t66 9.54355
R45900 a_31953_n19727.t66 a_31953_n19727.n91 9.54355
R45901 a_31953_n19727.t68 a_31953_n19727.n92 9.54355
R45902 a_31953_n19727.n89 a_31953_n19727.t68 9.54355
R45903 a_31953_n19727.n294 a_31953_n19727.t188 9.54355
R45904 a_31953_n19727.n295 a_31953_n19727.t188 9.54355
R45905 a_31953_n19727.n310 a_31953_n19727.t252 9.54355
R45906 a_31953_n19727.t252 a_31953_n19727.n309 9.54355
R45907 a_31953_n19727.t163 a_31953_n19727.n97 9.54355
R45908 a_31953_n19727.n95 a_31953_n19727.t163 9.54355
R45909 a_31953_n19727.n96 a_31953_n19727.t153 9.54355
R45910 a_31953_n19727.t153 a_31953_n19727.n94 9.54355
R45911 a_31953_n19727.n312 a_31953_n19727.t265 9.54355
R45912 a_31953_n19727.n311 a_31953_n19727.t265 9.54355
R45913 a_31953_n19727.n314 a_31953_n19727.t321 9.54355
R45914 a_31953_n19727.t321 a_31953_n19727.n313 9.54355
R45915 a_31953_n19727.t241 a_31953_n19727.n102 9.54355
R45916 a_31953_n19727.n99 a_31953_n19727.t241 9.54355
R45917 a_31953_n19727.n100 a_31953_n19727.t232 9.54355
R45918 a_31953_n19727.t232 a_31953_n19727.n98 9.54355
R45919 a_31953_n19727.n316 a_31953_n19727.t335 9.54355
R45920 a_31953_n19727.n315 a_31953_n19727.t335 9.54355
R45921 a_31953_n19727.n318 a_31953_n19727.t297 9.54355
R45922 a_31953_n19727.t297 a_31953_n19727.n317 9.54355
R45923 a_31953_n19727.t216 a_31953_n19727.n106 9.54355
R45924 a_31953_n19727.n104 a_31953_n19727.t216 9.54355
R45925 a_31953_n19727.n105 a_31953_n19727.t211 9.54355
R45926 a_31953_n19727.t211 a_31953_n19727.n103 9.54355
R45927 a_31953_n19727.n320 a_31953_n19727.t306 9.54355
R45928 a_31953_n19727.n319 a_31953_n19727.t306 9.54355
R45929 a_31953_n19727.n364 a_31953_n19727.t315 9.54355
R45930 a_31953_n19727.t350 a_31953_n19727.n368 9.54355
R45931 a_31953_n19727.n367 a_31953_n19727.t283 9.54355
R45932 a_31953_n19727.n366 a_31953_n19727.t243 9.54355
R45933 a_31953_n19727.t96 a_31953_n19727.n359 9.54355
R45934 a_31953_n19727.n360 a_31953_n19727.t96 9.54355
R45935 a_31953_n19727.n111 a_31953_n19727.t131 9.54355
R45936 a_31953_n19727.t131 a_31953_n19727.n109 9.54355
R45937 a_31953_n19727.t353 a_31953_n19727.n110 9.54355
R45938 a_31953_n19727.n107 a_31953_n19727.t353 9.54355
R45939 a_31953_n19727.n361 a_31953_n19727.t313 9.54355
R45940 a_31953_n19727.n362 a_31953_n19727.t313 9.54355
R45941 a_31953_n19727.t171 a_31953_n19727.n355 9.54355
R45942 a_31953_n19727.n356 a_31953_n19727.t171 9.54355
R45943 a_31953_n19727.n116 a_31953_n19727.t206 9.54355
R45944 a_31953_n19727.t206 a_31953_n19727.n114 9.54355
R45945 a_31953_n19727.t136 a_31953_n19727.n115 9.54355
R45946 a_31953_n19727.n112 a_31953_n19727.t136 9.54355
R45947 a_31953_n19727.n357 a_31953_n19727.t92 9.54355
R45948 a_31953_n19727.n358 a_31953_n19727.t92 9.54355
R45949 a_31953_n19727.n326 a_31953_n19727.t156 9.54355
R45950 a_31953_n19727.t156 a_31953_n19727.n325 9.54355
R45951 a_31953_n19727.t44 a_31953_n19727.n120 9.54355
R45952 a_31953_n19727.n118 a_31953_n19727.t44 9.54355
R45953 a_31953_n19727.n119 a_31953_n19727.t58 9.54355
R45954 a_31953_n19727.t58 a_31953_n19727.n117 9.54355
R45955 a_31953_n19727.n328 a_31953_n19727.t82 9.54355
R45956 a_31953_n19727.n327 a_31953_n19727.t82 9.54355
R45957 a_31953_n19727.n330 a_31953_n19727.t236 9.54355
R45958 a_31953_n19727.t236 a_31953_n19727.n329 9.54355
R45959 a_31953_n19727.t24 a_31953_n19727.n125 9.54355
R45960 a_31953_n19727.n122 a_31953_n19727.t24 9.54355
R45961 a_31953_n19727.n123 a_31953_n19727.t42 9.54355
R45962 a_31953_n19727.t42 a_31953_n19727.n121 9.54355
R45963 a_31953_n19727.n332 a_31953_n19727.t154 9.54355
R45964 a_31953_n19727.n331 a_31953_n19727.t154 9.54355
R45965 a_31953_n19727.n334 a_31953_n19727.t294 9.54355
R45966 a_31953_n19727.t294 a_31953_n19727.n333 9.54355
R45967 a_31953_n19727.t8 a_31953_n19727.n129 9.54355
R45968 a_31953_n19727.n127 a_31953_n19727.t8 9.54355
R45969 a_31953_n19727.n128 a_31953_n19727.t30 9.54355
R45970 a_31953_n19727.t30 a_31953_n19727.n126 9.54355
R45971 a_31953_n19727.n336 a_31953_n19727.t219 9.54355
R45972 a_31953_n19727.n335 a_31953_n19727.t219 9.54355
R45973 a_31953_n19727.t75 a_31953_n19727.n346 9.54355
R45974 a_31953_n19727.n347 a_31953_n19727.t75 9.54355
R45975 a_31953_n19727.n134 a_31953_n19727.t105 9.54355
R45976 a_31953_n19727.t105 a_31953_n19727.n132 9.54355
R45977 a_31953_n19727.t332 a_31953_n19727.n133 9.54355
R45978 a_31953_n19727.n130 a_31953_n19727.t332 9.54355
R45979 a_31953_n19727.n348 a_31953_n19727.t291 9.54355
R45980 a_31953_n19727.n349 a_31953_n19727.t291 9.54355
R45981 a_31953_n19727.t134 a_31953_n19727.n342 9.54355
R45982 a_31953_n19727.n343 a_31953_n19727.t134 9.54355
R45983 a_31953_n19727.n138 a_31953_n19727.t162 9.54355
R45984 a_31953_n19727.t162 a_31953_n19727.n136 9.54355
R45985 a_31953_n19727.t93 a_31953_n19727.n137 9.54355
R45986 a_31953_n19727.n135 a_31953_n19727.t93 9.54355
R45987 a_31953_n19727.n344 a_31953_n19727.t352 9.54355
R45988 a_31953_n19727.n345 a_31953_n19727.t352 9.54355
R45989 a_31953_n19727.t213 a_31953_n19727.n340 9.54355
R45990 a_31953_n19727.n341 a_31953_n19727.t213 9.54355
R45991 a_31953_n19727.n141 a_31953_n19727.t239 9.54355
R45992 a_31953_n19727.t239 a_31953_n19727.n139 9.54355
R45993 a_31953_n19727.n140 a_31953_n19727.t167 9.54355
R45994 a_31953_n19727.n337 a_31953_n19727.t167 9.54355
R45995 a_31953_n19727.n339 a_31953_n19727.t133 9.54355
R45996 a_31953_n19727.n338 a_31953_n19727.t133 9.54355
R45997 a_31953_n19727.n373 a_31953_n19727.t316 9.54355
R45998 a_31953_n19727.t130 a_31953_n19727.n377 9.54355
R45999 a_31953_n19727.n376 a_31953_n19727.t348 9.54355
R46000 a_31953_n19727.n375 a_31953_n19727.t132 9.54355
R46001 a_31953_n19727.n379 a_31953_n19727.t97 9.54355
R46002 a_31953_n19727.t97 a_31953_n19727.n378 9.54355
R46003 a_31953_n19727.t205 a_31953_n19727.n146 9.54355
R46004 a_31953_n19727.n143 a_31953_n19727.t205 9.54355
R46005 a_31953_n19727.n144 a_31953_n19727.t127 9.54355
R46006 a_31953_n19727.t127 a_31953_n19727.n142 9.54355
R46007 a_31953_n19727.n381 a_31953_n19727.t207 9.54355
R46008 a_31953_n19727.n380 a_31953_n19727.t207 9.54355
R46009 a_31953_n19727.n383 a_31953_n19727.t85 9.54355
R46010 a_31953_n19727.t85 a_31953_n19727.n382 9.54355
R46011 a_31953_n19727.t192 a_31953_n19727.n150 9.54355
R46012 a_31953_n19727.n148 a_31953_n19727.t192 9.54355
R46013 a_31953_n19727.n149 a_31953_n19727.t118 9.54355
R46014 a_31953_n19727.t118 a_31953_n19727.n147 9.54355
R46015 a_31953_n19727.n385 a_31953_n19727.t194 9.54355
R46016 a_31953_n19727.n384 a_31953_n19727.t194 9.54355
R46017 a_31953_n19727.t157 a_31953_n19727.n394 9.54355
R46018 a_31953_n19727.n395 a_31953_n19727.t157 9.54355
R46019 a_31953_n19727.n155 a_31953_n19727.t26 9.54355
R46020 a_31953_n19727.t26 a_31953_n19727.n153 9.54355
R46021 a_31953_n19727.t46 a_31953_n19727.n154 9.54355
R46022 a_31953_n19727.n151 a_31953_n19727.t46 9.54355
R46023 a_31953_n19727.n396 a_31953_n19727.t269 9.54355
R46024 a_31953_n19727.n397 a_31953_n19727.t269 9.54355
R46025 a_31953_n19727.t237 a_31953_n19727.n390 9.54355
R46026 a_31953_n19727.n391 a_31953_n19727.t237 9.54355
R46027 a_31953_n19727.n159 a_31953_n19727.t4 9.54355
R46028 a_31953_n19727.t4 a_31953_n19727.n157 9.54355
R46029 a_31953_n19727.t28 a_31953_n19727.n158 9.54355
R46030 a_31953_n19727.n156 a_31953_n19727.t28 9.54355
R46031 a_31953_n19727.n392 a_31953_n19727.t341 9.54355
R46032 a_31953_n19727.n393 a_31953_n19727.t341 9.54355
R46033 a_31953_n19727.t225 a_31953_n19727.n386 9.54355
R46034 a_31953_n19727.n387 a_31953_n19727.t225 9.54355
R46035 a_31953_n19727.n164 a_31953_n19727.t6 9.54355
R46036 a_31953_n19727.t6 a_31953_n19727.n162 9.54355
R46037 a_31953_n19727.t32 a_31953_n19727.n163 9.54355
R46038 a_31953_n19727.n160 a_31953_n19727.t32 9.54355
R46039 a_31953_n19727.n388 a_31953_n19727.t324 9.54355
R46040 a_31953_n19727.n389 a_31953_n19727.t324 9.54355
R46041 a_31953_n19727.n404 a_31953_n19727.t298 9.54355
R46042 a_31953_n19727.t298 a_31953_n19727.n403 9.54355
R46043 a_31953_n19727.t107 a_31953_n19727.n168 9.54355
R46044 a_31953_n19727.n166 a_31953_n19727.t107 9.54355
R46045 a_31953_n19727.n167 a_31953_n19727.t322 9.54355
R46046 a_31953_n19727.t322 a_31953_n19727.n165 9.54355
R46047 a_31953_n19727.n406 a_31953_n19727.t109 9.54355
R46048 a_31953_n19727.n405 a_31953_n19727.t109 9.54355
R46049 a_31953_n19727.n408 a_31953_n19727.t77 9.54355
R46050 a_31953_n19727.t77 a_31953_n19727.n407 9.54355
R46051 a_31953_n19727.t183 a_31953_n19727.n173 9.54355
R46052 a_31953_n19727.n170 a_31953_n19727.t183 9.54355
R46053 a_31953_n19727.n171 a_31953_n19727.t106 9.54355
R46054 a_31953_n19727.t106 a_31953_n19727.n169 9.54355
R46055 a_31953_n19727.n410 a_31953_n19727.t185 9.54355
R46056 a_31953_n19727.n409 a_31953_n19727.t185 9.54355
R46057 a_31953_n19727.n412 a_31953_n19727.t349 9.54355
R46058 a_31953_n19727.t349 a_31953_n19727.n411 9.54355
R46059 a_31953_n19727.t147 a_31953_n19727.n177 9.54355
R46060 a_31953_n19727.n175 a_31953_n19727.t147 9.54355
R46061 a_31953_n19727.n176 a_31953_n19727.t76 9.54355
R46062 a_31953_n19727.t76 a_31953_n19727.n174 9.54355
R46063 a_31953_n19727.n414 a_31953_n19727.t150 9.54355
R46064 a_31953_n19727.n413 a_31953_n19727.t150 9.54355
R46065 a_31953_n19727.n457 a_31953_n19727.t196 9.54355
R46066 a_31953_n19727.t148 a_31953_n19727.n461 9.54355
R46067 a_31953_n19727.n460 a_31953_n19727.t227 9.54355
R46068 a_31953_n19727.n459 a_31953_n19727.t123 9.54355
R46069 a_31953_n19727.t272 a_31953_n19727.n452 9.54355
R46070 a_31953_n19727.n453 a_31953_n19727.t272 9.54355
R46071 a_31953_n19727.n182 a_31953_n19727.t228 9.54355
R46072 a_31953_n19727.t228 a_31953_n19727.n180 9.54355
R46073 a_31953_n19727.t301 a_31953_n19727.n181 9.54355
R46074 a_31953_n19727.n178 a_31953_n19727.t301 9.54355
R46075 a_31953_n19727.n454 a_31953_n19727.t199 9.54355
R46076 a_31953_n19727.n455 a_31953_n19727.t199 9.54355
R46077 a_31953_n19727.t344 a_31953_n19727.n448 9.54355
R46078 a_31953_n19727.n449 a_31953_n19727.t344 9.54355
R46079 a_31953_n19727.n187 a_31953_n19727.t302 9.54355
R46080 a_31953_n19727.t302 a_31953_n19727.n185 9.54355
R46081 a_31953_n19727.t83 a_31953_n19727.n186 9.54355
R46082 a_31953_n19727.n183 a_31953_n19727.t83 9.54355
R46083 a_31953_n19727.n450 a_31953_n19727.t277 9.54355
R46084 a_31953_n19727.n451 a_31953_n19727.t277 9.54355
R46085 a_31953_n19727.n419 a_31953_n19727.t328 9.54355
R46086 a_31953_n19727.t328 a_31953_n19727.n418 9.54355
R46087 a_31953_n19727.t22 a_31953_n19727.n191 9.54355
R46088 a_31953_n19727.n189 a_31953_n19727.t22 9.54355
R46089 a_31953_n19727.n190 a_31953_n19727.t2 9.54355
R46090 a_31953_n19727.t2 a_31953_n19727.n188 9.54355
R46091 a_31953_n19727.n421 a_31953_n19727.t263 9.54355
R46092 a_31953_n19727.n420 a_31953_n19727.t263 9.54355
R46093 a_31953_n19727.n423 a_31953_n19727.t113 9.54355
R46094 a_31953_n19727.t113 a_31953_n19727.n422 9.54355
R46095 a_31953_n19727.t0 a_31953_n19727.n196 9.54355
R46096 a_31953_n19727.n193 a_31953_n19727.t0 9.54355
R46097 a_31953_n19727.n194 a_31953_n19727.t54 9.54355
R46098 a_31953_n19727.t54 a_31953_n19727.n192 9.54355
R46099 a_31953_n19727.n425 a_31953_n19727.t334 9.54355
R46100 a_31953_n19727.n424 a_31953_n19727.t334 9.54355
R46101 a_31953_n19727.n427 a_31953_n19727.t169 9.54355
R46102 a_31953_n19727.t169 a_31953_n19727.n426 9.54355
R46103 a_31953_n19727.t56 a_31953_n19727.n200 9.54355
R46104 a_31953_n19727.n198 a_31953_n19727.t56 9.54355
R46105 a_31953_n19727.n199 a_31953_n19727.t40 9.54355
R46106 a_31953_n19727.t40 a_31953_n19727.n197 9.54355
R46107 a_31953_n19727.n429 a_31953_n19727.t101 9.54355
R46108 a_31953_n19727.n428 a_31953_n19727.t101 9.54355
R46109 a_31953_n19727.t247 a_31953_n19727.n439 9.54355
R46110 a_31953_n19727.n440 a_31953_n19727.t247 9.54355
R46111 a_31953_n19727.n205 a_31953_n19727.t212 9.54355
R46112 a_31953_n19727.t212 a_31953_n19727.n203 9.54355
R46113 a_31953_n19727.t287 a_31953_n19727.n204 9.54355
R46114 a_31953_n19727.n201 a_31953_n19727.t287 9.54355
R46115 a_31953_n19727.n441 a_31953_n19727.t176 9.54355
R46116 a_31953_n19727.n442 a_31953_n19727.t176 9.54355
R46117 a_31953_n19727.t303 a_31953_n19727.n435 9.54355
R46118 a_31953_n19727.n436 a_31953_n19727.t303 9.54355
R46119 a_31953_n19727.n209 a_31953_n19727.t267 9.54355
R46120 a_31953_n19727.t267 a_31953_n19727.n207 9.54355
R46121 a_31953_n19727.t338 a_31953_n19727.n208 9.54355
R46122 a_31953_n19727.n206 a_31953_n19727.t338 9.54355
R46123 a_31953_n19727.n437 a_31953_n19727.t233 9.54355
R46124 a_31953_n19727.n438 a_31953_n19727.t233 9.54355
R46125 a_31953_n19727.t84 a_31953_n19727.n433 9.54355
R46126 a_31953_n19727.n434 a_31953_n19727.t84 9.54355
R46127 a_31953_n19727.n212 a_31953_n19727.t339 9.54355
R46128 a_31953_n19727.t339 a_31953_n19727.n210 9.54355
R46129 a_31953_n19727.n211 a_31953_n19727.t120 9.54355
R46130 a_31953_n19727.n430 a_31953_n19727.t120 9.54355
R46131 a_31953_n19727.n432 a_31953_n19727.t307 9.54355
R46132 a_31953_n19727.n431 a_31953_n19727.t307 9.54355
R46133 a_31953_n19727.n321 a_31953_n19727.t73 6.62729
R46134 a_31953_n19727.n464 a_31953_n19727.n463 3.90251
R46135 a_31953_n19727.n463 a_31953_n19727.n225 3.89899
R46136 a_31953_n19727.n479 a_31953_n19727.t37 3.3605
R46137 a_31953_n19727.n227 a_31953_n19727.t13 3.3605
R46138 a_31953_n19727.n231 a_31953_n19727.t39 3.3605
R46139 a_31953_n19727.n230 a_31953_n19727.t17 3.3605
R46140 a_31953_n19727.n229 a_31953_n19727.t21 3.3605
R46141 a_31953_n19727.n259 a_31953_n19727.t61 3.3605
R46142 a_31953_n19727.n260 a_31953_n19727.t49 3.3605
R46143 a_31953_n19727.n261 a_31953_n19727.t53 3.3605
R46144 a_31953_n19727.n277 a_31953_n19727.t15 3.3605
R46145 a_31953_n19727.n276 a_31953_n19727.t65 3.3605
R46146 a_31953_n19727.n275 a_31953_n19727.t69 3.3605
R46147 a_31953_n19727.n305 a_31953_n19727.t11 3.3605
R46148 a_31953_n19727.n306 a_31953_n19727.t63 3.3605
R46149 a_31953_n19727.n307 a_31953_n19727.t67 3.3605
R46150 a_31953_n19727.n322 a_31953_n19727.t59 3.3605
R46151 a_31953_n19727.n323 a_31953_n19727.t43 3.3605
R46152 a_31953_n19727.n324 a_31953_n19727.t31 3.3605
R46153 a_31953_n19727.n353 a_31953_n19727.t45 3.3605
R46154 a_31953_n19727.n352 a_31953_n19727.t25 3.3605
R46155 a_31953_n19727.n351 a_31953_n19727.t9 3.3605
R46156 a_31953_n19727.n371 a_31953_n19727.t47 3.3605
R46157 a_31953_n19727.n370 a_31953_n19727.t29 3.3605
R46158 a_31953_n19727.n369 a_31953_n19727.t33 3.3605
R46159 a_31953_n19727.n399 a_31953_n19727.t27 3.3605
R46160 a_31953_n19727.n400 a_31953_n19727.t5 3.3605
R46161 a_31953_n19727.n401 a_31953_n19727.t7 3.3605
R46162 a_31953_n19727.n415 a_31953_n19727.t3 3.3605
R46163 a_31953_n19727.n416 a_31953_n19727.t55 3.3605
R46164 a_31953_n19727.n417 a_31953_n19727.t41 3.3605
R46165 a_31953_n19727.n446 a_31953_n19727.t23 3.3605
R46166 a_31953_n19727.n445 a_31953_n19727.t1 3.3605
R46167 a_31953_n19727.n444 a_31953_n19727.t57 3.3605
R46168 a_31953_n19727.n481 a_31953_n19727.t51 3.3605
R46169 a_31953_n19727.n480 a_31953_n19727.t35 3.3605
R46170 a_31953_n19727.n228 a_31953_n19727.t19 3.3605
R46171 a_31953_n19727.t71 a_31953_n19727.n509 3.3605
R46172 a_31953_n19727.n258 a_31953_n19727.n231 2.59662
R46173 a_31953_n19727.n304 a_31953_n19727.n277 2.59662
R46174 a_31953_n19727.n354 a_31953_n19727.n322 2.59662
R46175 a_31953_n19727.n398 a_31953_n19727.n371 2.59662
R46176 a_31953_n19727.n447 a_31953_n19727.n415 2.59662
R46177 a_31953_n19727.n482 a_31953_n19727.n479 2.59562
R46178 a_31953_n19727.n262 a_31953_n19727.n229 2.59544
R46179 a_31953_n19727.n308 a_31953_n19727.n275 2.59544
R46180 a_31953_n19727.n350 a_31953_n19727.n324 2.59544
R46181 a_31953_n19727.n402 a_31953_n19727.n369 2.59544
R46182 a_31953_n19727.n443 a_31953_n19727.n417 2.59544
R46183 a_31953_n19727.n509 a_31953_n19727.n508 2.59544
R46184 a_31953_n19727.n259 a_31953_n19727.n258 2.58354
R46185 a_31953_n19727.n305 a_31953_n19727.n304 2.58354
R46186 a_31953_n19727.n354 a_31953_n19727.n353 2.58354
R46187 a_31953_n19727.n399 a_31953_n19727.n398 2.58354
R46188 a_31953_n19727.n447 a_31953_n19727.n446 2.58354
R46189 a_31953_n19727.n482 a_31953_n19727.n481 2.58354
R46190 a_31953_n19727.n262 a_31953_n19727.n261 2.58235
R46191 a_31953_n19727.n308 a_31953_n19727.n307 2.58235
R46192 a_31953_n19727.n351 a_31953_n19727.n350 2.58235
R46193 a_31953_n19727.n402 a_31953_n19727.n401 2.58235
R46194 a_31953_n19727.n444 a_31953_n19727.n443 2.58235
R46195 a_31953_n19727.n508 a_31953_n19727.n228 2.58235
R46196 a_31953_n19727.n225 a_31953_n19727.n226 0.0196917
R46197 a_31953_n19727.n131 a_31953_n19727.n139 1.6805
R46198 a_31953_n19727.n202 a_31953_n19727.n210 1.6805
R46199 a_31953_n19727.n60 a_31953_n19727.n68 1.6805
R46200 a_31953_n19727.n74 a_31953_n19727.n218 1.59324
R46201 a_31953_n19727.n145 a_31953_n19727.n222 1.59324
R46202 a_31953_n19727.n3 a_31953_n19727.n214 1.59324
R46203 a_31953_n19727.n350 a_31953_n19727.n131 1.5005
R46204 a_31953_n19727.n113 a_31953_n19727.n354 1.5005
R46205 a_31953_n19727.n90 a_31953_n19727.n308 1.5005
R46206 a_31953_n19727.n304 a_31953_n19727.n74 1.5005
R46207 a_31953_n19727.n131 a_31953_n19727.n141 1.5005
R46208 a_31953_n19727.n131 a_31953_n19727.n138 1.5005
R46209 a_31953_n19727.n136 a_31953_n19727.n131 1.5005
R46210 a_31953_n19727.n131 a_31953_n19727.n134 1.5005
R46211 a_31953_n19727.n132 a_31953_n19727.n131 1.5005
R46212 a_31953_n19727.n129 a_31953_n19727.n124 1.5005
R46213 a_31953_n19727.n131 a_31953_n19727.n127 1.5005
R46214 a_31953_n19727.n125 a_31953_n19727.n124 1.5005
R46215 a_31953_n19727.n124 a_31953_n19727.n122 1.5005
R46216 a_31953_n19727.n120 a_31953_n19727.n113 1.5005
R46217 a_31953_n19727.n124 a_31953_n19727.n118 1.5005
R46218 a_31953_n19727.n108 a_31953_n19727.n116 1.5005
R46219 a_31953_n19727.n114 a_31953_n19727.n113 1.5005
R46220 a_31953_n19727.n108 a_31953_n19727.n111 1.5005
R46221 a_31953_n19727.n109 a_31953_n19727.n108 1.5005
R46222 a_31953_n19727.n108 a_31953_n19727.n220 1.5005
R46223 a_31953_n19727.n106 a_31953_n19727.n101 1.5005
R46224 a_31953_n19727.n101 a_31953_n19727.n104 1.5005
R46225 a_31953_n19727.n102 a_31953_n19727.n101 1.5005
R46226 a_31953_n19727.n101 a_31953_n19727.n99 1.5005
R46227 a_31953_n19727.n97 a_31953_n19727.n90 1.5005
R46228 a_31953_n19727.n101 a_31953_n19727.n95 1.5005
R46229 a_31953_n19727.n81 a_31953_n19727.n93 1.5005
R46230 a_31953_n19727.n91 a_31953_n19727.n90 1.5005
R46231 a_31953_n19727.n81 a_31953_n19727.n88 1.5005
R46232 a_31953_n19727.n86 a_31953_n19727.n81 1.5005
R46233 a_31953_n19727.n74 a_31953_n19727.n84 1.5005
R46234 a_31953_n19727.n82 a_31953_n19727.n81 1.5005
R46235 a_31953_n19727.n79 a_31953_n19727.n74 1.5005
R46236 a_31953_n19727.n74 a_31953_n19727.n77 1.5005
R46237 a_31953_n19727.n75 a_31953_n19727.n74 1.5005
R46238 a_31953_n19727.n74 a_31953_n19727.n72 1.5005
R46239 a_31953_n19727.n443 a_31953_n19727.n202 1.5005
R46240 a_31953_n19727.n184 a_31953_n19727.n447 1.5005
R46241 a_31953_n19727.n161 a_31953_n19727.n402 1.5005
R46242 a_31953_n19727.n398 a_31953_n19727.n145 1.5005
R46243 a_31953_n19727.n202 a_31953_n19727.n212 1.5005
R46244 a_31953_n19727.n202 a_31953_n19727.n209 1.5005
R46245 a_31953_n19727.n207 a_31953_n19727.n202 1.5005
R46246 a_31953_n19727.n202 a_31953_n19727.n205 1.5005
R46247 a_31953_n19727.n203 a_31953_n19727.n202 1.5005
R46248 a_31953_n19727.n200 a_31953_n19727.n195 1.5005
R46249 a_31953_n19727.n202 a_31953_n19727.n198 1.5005
R46250 a_31953_n19727.n196 a_31953_n19727.n195 1.5005
R46251 a_31953_n19727.n195 a_31953_n19727.n193 1.5005
R46252 a_31953_n19727.n191 a_31953_n19727.n184 1.5005
R46253 a_31953_n19727.n195 a_31953_n19727.n189 1.5005
R46254 a_31953_n19727.n179 a_31953_n19727.n187 1.5005
R46255 a_31953_n19727.n185 a_31953_n19727.n184 1.5005
R46256 a_31953_n19727.n179 a_31953_n19727.n182 1.5005
R46257 a_31953_n19727.n180 a_31953_n19727.n179 1.5005
R46258 a_31953_n19727.n179 a_31953_n19727.n224 1.5005
R46259 a_31953_n19727.n177 a_31953_n19727.n172 1.5005
R46260 a_31953_n19727.n172 a_31953_n19727.n175 1.5005
R46261 a_31953_n19727.n173 a_31953_n19727.n172 1.5005
R46262 a_31953_n19727.n172 a_31953_n19727.n170 1.5005
R46263 a_31953_n19727.n168 a_31953_n19727.n161 1.5005
R46264 a_31953_n19727.n172 a_31953_n19727.n166 1.5005
R46265 a_31953_n19727.n152 a_31953_n19727.n164 1.5005
R46266 a_31953_n19727.n162 a_31953_n19727.n161 1.5005
R46267 a_31953_n19727.n152 a_31953_n19727.n159 1.5005
R46268 a_31953_n19727.n157 a_31953_n19727.n152 1.5005
R46269 a_31953_n19727.n145 a_31953_n19727.n155 1.5005
R46270 a_31953_n19727.n153 a_31953_n19727.n152 1.5005
R46271 a_31953_n19727.n150 a_31953_n19727.n145 1.5005
R46272 a_31953_n19727.n145 a_31953_n19727.n148 1.5005
R46273 a_31953_n19727.n146 a_31953_n19727.n145 1.5005
R46274 a_31953_n19727.n145 a_31953_n19727.n143 1.5005
R46275 a_31953_n19727.n48 a_31953_n19727.n482 1.5005
R46276 a_31953_n19727.n19 a_31953_n19727.n262 1.5005
R46277 a_31953_n19727.n258 a_31953_n19727.n3 1.5005
R46278 a_31953_n19727.n60 a_31953_n19727.n70 1.5005
R46279 a_31953_n19727.n60 a_31953_n19727.n67 1.5005
R46280 a_31953_n19727.n65 a_31953_n19727.n60 1.5005
R46281 a_31953_n19727.n60 a_31953_n19727.n63 1.5005
R46282 a_31953_n19727.n61 a_31953_n19727.n60 1.5005
R46283 a_31953_n19727.n58 a_31953_n19727.n53 1.5005
R46284 a_31953_n19727.n60 a_31953_n19727.n56 1.5005
R46285 a_31953_n19727.n54 a_31953_n19727.n53 1.5005
R46286 a_31953_n19727.n53 a_31953_n19727.n51 1.5005
R46287 a_31953_n19727.n49 a_31953_n19727.n48 1.5005
R46288 a_31953_n19727.n53 a_31953_n19727.n46 1.5005
R46289 a_31953_n19727.n44 a_31953_n19727.n39 1.5005
R46290 a_31953_n19727.n48 a_31953_n19727.n42 1.5005
R46291 a_31953_n19727.n40 a_31953_n19727.n39 1.5005
R46292 a_31953_n19727.n39 a_31953_n19727.n37 1.5005
R46293 a_31953_n19727.n39 a_31953_n19727.n216 1.5005
R46294 a_31953_n19727.n35 a_31953_n19727.n30 1.5005
R46295 a_31953_n19727.n30 a_31953_n19727.n33 1.5005
R46296 a_31953_n19727.n31 a_31953_n19727.n30 1.5005
R46297 a_31953_n19727.n30 a_31953_n19727.n28 1.5005
R46298 a_31953_n19727.n26 a_31953_n19727.n19 1.5005
R46299 a_31953_n19727.n30 a_31953_n19727.n24 1.5005
R46300 a_31953_n19727.n10 a_31953_n19727.n22 1.5005
R46301 a_31953_n19727.n20 a_31953_n19727.n19 1.5005
R46302 a_31953_n19727.n10 a_31953_n19727.n17 1.5005
R46303 a_31953_n19727.n15 a_31953_n19727.n10 1.5005
R46304 a_31953_n19727.n3 a_31953_n19727.n13 1.5005
R46305 a_31953_n19727.n11 a_31953_n19727.n10 1.5005
R46306 a_31953_n19727.n8 a_31953_n19727.n3 1.5005
R46307 a_31953_n19727.n3 a_31953_n19727.n6 1.5005
R46308 a_31953_n19727.n4 a_31953_n19727.n3 1.5005
R46309 a_31953_n19727.n3 a_31953_n19727.n1 1.5005
R46310 a_31953_n19727.n508 a_31953_n19727.n60 1.5005
R46311 a_31953_n19727.n260 a_31953_n19727.n259 1.06274
R46312 a_31953_n19727.n261 a_31953_n19727.n260 1.06274
R46313 a_31953_n19727.n231 a_31953_n19727.n230 1.06274
R46314 a_31953_n19727.n230 a_31953_n19727.n229 1.06274
R46315 a_31953_n19727.n306 a_31953_n19727.n305 1.06274
R46316 a_31953_n19727.n307 a_31953_n19727.n306 1.06274
R46317 a_31953_n19727.n277 a_31953_n19727.n276 1.06274
R46318 a_31953_n19727.n276 a_31953_n19727.n275 1.06274
R46319 a_31953_n19727.n353 a_31953_n19727.n352 1.06274
R46320 a_31953_n19727.n352 a_31953_n19727.n351 1.06274
R46321 a_31953_n19727.n323 a_31953_n19727.n322 1.06274
R46322 a_31953_n19727.n324 a_31953_n19727.n323 1.06274
R46323 a_31953_n19727.n400 a_31953_n19727.n399 1.06274
R46324 a_31953_n19727.n401 a_31953_n19727.n400 1.06274
R46325 a_31953_n19727.n371 a_31953_n19727.n370 1.06274
R46326 a_31953_n19727.n370 a_31953_n19727.n369 1.06274
R46327 a_31953_n19727.n446 a_31953_n19727.n445 1.06274
R46328 a_31953_n19727.n445 a_31953_n19727.n444 1.06274
R46329 a_31953_n19727.n416 a_31953_n19727.n415 1.06274
R46330 a_31953_n19727.n417 a_31953_n19727.n416 1.06274
R46331 a_31953_n19727.n481 a_31953_n19727.n480 1.06274
R46332 a_31953_n19727.n480 a_31953_n19727.n228 1.06274
R46333 a_31953_n19727.n479 a_31953_n19727.n227 1.06274
R46334 a_31953_n19727.n509 a_31953_n19727.n227 1.06274
R46335 a_31953_n19727.n236 a_31953_n19727.n235 0.97759
R46336 a_31953_n19727.n237 a_31953_n19727.n233 0.97759
R46337 a_31953_n19727.n240 a_31953_n19727.n0 0.97759
R46338 a_31953_n19727.n1 a_31953_n19727.n238 0.97759
R46339 a_31953_n19727.n2 a_31953_n19727.n241 0.97759
R46340 a_31953_n19727.n4 a_31953_n19727.n239 0.97759
R46341 a_31953_n19727.n244 a_31953_n19727.n5 0.97759
R46342 a_31953_n19727.n6 a_31953_n19727.n242 0.97759
R46343 a_31953_n19727.n7 a_31953_n19727.n245 0.97759
R46344 a_31953_n19727.n8 a_31953_n19727.n243 0.97759
R46345 a_31953_n19727.n9 a_31953_n19727.n257 0.97759
R46346 a_31953_n19727.n11 a_31953_n19727.n255 0.97759
R46347 a_31953_n19727.n256 a_31953_n19727.n12 0.97759
R46348 a_31953_n19727.n13 a_31953_n19727.n254 0.97759
R46349 a_31953_n19727.n14 a_31953_n19727.n253 0.97759
R46350 a_31953_n19727.n15 a_31953_n19727.n251 0.97759
R46351 a_31953_n19727.n252 a_31953_n19727.n16 0.97759
R46352 a_31953_n19727.n17 a_31953_n19727.n250 0.97759
R46353 a_31953_n19727.n18 a_31953_n19727.n249 0.97759
R46354 a_31953_n19727.n20 a_31953_n19727.n247 0.97759
R46355 a_31953_n19727.n248 a_31953_n19727.n21 0.97759
R46356 a_31953_n19727.n22 a_31953_n19727.n246 0.97759
R46357 a_31953_n19727.n265 a_31953_n19727.n23 0.97759
R46358 a_31953_n19727.n24 a_31953_n19727.n263 0.97759
R46359 a_31953_n19727.n25 a_31953_n19727.n266 0.97759
R46360 a_31953_n19727.n26 a_31953_n19727.n264 0.97759
R46361 a_31953_n19727.n269 a_31953_n19727.n27 0.97759
R46362 a_31953_n19727.n28 a_31953_n19727.n267 0.97759
R46363 a_31953_n19727.n29 a_31953_n19727.n270 0.97759
R46364 a_31953_n19727.n31 a_31953_n19727.n268 0.97759
R46365 a_31953_n19727.n273 a_31953_n19727.n32 0.97759
R46366 a_31953_n19727.n33 a_31953_n19727.n271 0.97759
R46367 a_31953_n19727.n34 a_31953_n19727.n274 0.97759
R46368 a_31953_n19727.n35 a_31953_n19727.n272 0.97759
R46369 a_31953_n19727.n469 a_31953_n19727.n468 0.97759
R46370 a_31953_n19727.n470 a_31953_n19727.n466 0.97759
R46371 a_31953_n19727.n473 a_31953_n19727.n36 0.97759
R46372 a_31953_n19727.n37 a_31953_n19727.n471 0.97759
R46373 a_31953_n19727.n38 a_31953_n19727.n474 0.97759
R46374 a_31953_n19727.n40 a_31953_n19727.n472 0.97759
R46375 a_31953_n19727.n477 a_31953_n19727.n41 0.97759
R46376 a_31953_n19727.n42 a_31953_n19727.n475 0.97759
R46377 a_31953_n19727.n43 a_31953_n19727.n478 0.97759
R46378 a_31953_n19727.n44 a_31953_n19727.n476 0.97759
R46379 a_31953_n19727.n485 a_31953_n19727.n45 0.97759
R46380 a_31953_n19727.n46 a_31953_n19727.n483 0.97759
R46381 a_31953_n19727.n47 a_31953_n19727.n486 0.97759
R46382 a_31953_n19727.n49 a_31953_n19727.n484 0.97759
R46383 a_31953_n19727.n489 a_31953_n19727.n50 0.97759
R46384 a_31953_n19727.n51 a_31953_n19727.n487 0.97759
R46385 a_31953_n19727.n52 a_31953_n19727.n490 0.97759
R46386 a_31953_n19727.n54 a_31953_n19727.n488 0.97759
R46387 a_31953_n19727.n493 a_31953_n19727.n55 0.97759
R46388 a_31953_n19727.n56 a_31953_n19727.n491 0.97759
R46389 a_31953_n19727.n57 a_31953_n19727.n494 0.97759
R46390 a_31953_n19727.n58 a_31953_n19727.n492 0.97759
R46391 a_31953_n19727.n59 a_31953_n19727.n507 0.97759
R46392 a_31953_n19727.n61 a_31953_n19727.n505 0.97759
R46393 a_31953_n19727.n506 a_31953_n19727.n62 0.97759
R46394 a_31953_n19727.n63 a_31953_n19727.n504 0.97759
R46395 a_31953_n19727.n64 a_31953_n19727.n503 0.97759
R46396 a_31953_n19727.n65 a_31953_n19727.n501 0.97759
R46397 a_31953_n19727.n502 a_31953_n19727.n66 0.97759
R46398 a_31953_n19727.n67 a_31953_n19727.n500 0.97759
R46399 a_31953_n19727.n496 a_31953_n19727.n495 0.97759
R46400 a_31953_n19727.n68 a_31953_n19727.n499 0.97759
R46401 a_31953_n19727.n69 a_31953_n19727.n497 0.97759
R46402 a_31953_n19727.n70 a_31953_n19727.n498 0.97759
R46403 a_31953_n19727.n282 a_31953_n19727.n281 0.97759
R46404 a_31953_n19727.n283 a_31953_n19727.n279 0.97759
R46405 a_31953_n19727.n286 a_31953_n19727.n71 0.97759
R46406 a_31953_n19727.n72 a_31953_n19727.n284 0.97759
R46407 a_31953_n19727.n73 a_31953_n19727.n287 0.97759
R46408 a_31953_n19727.n75 a_31953_n19727.n285 0.97759
R46409 a_31953_n19727.n290 a_31953_n19727.n76 0.97759
R46410 a_31953_n19727.n77 a_31953_n19727.n288 0.97759
R46411 a_31953_n19727.n78 a_31953_n19727.n291 0.97759
R46412 a_31953_n19727.n79 a_31953_n19727.n289 0.97759
R46413 a_31953_n19727.n80 a_31953_n19727.n303 0.97759
R46414 a_31953_n19727.n82 a_31953_n19727.n301 0.97759
R46415 a_31953_n19727.n302 a_31953_n19727.n83 0.97759
R46416 a_31953_n19727.n84 a_31953_n19727.n300 0.97759
R46417 a_31953_n19727.n85 a_31953_n19727.n299 0.97759
R46418 a_31953_n19727.n86 a_31953_n19727.n297 0.97759
R46419 a_31953_n19727.n298 a_31953_n19727.n87 0.97759
R46420 a_31953_n19727.n88 a_31953_n19727.n296 0.97759
R46421 a_31953_n19727.n89 a_31953_n19727.n295 0.97759
R46422 a_31953_n19727.n91 a_31953_n19727.n293 0.97759
R46423 a_31953_n19727.n294 a_31953_n19727.n92 0.97759
R46424 a_31953_n19727.n93 a_31953_n19727.n292 0.97759
R46425 a_31953_n19727.n311 a_31953_n19727.n94 0.97759
R46426 a_31953_n19727.n95 a_31953_n19727.n309 0.97759
R46427 a_31953_n19727.n96 a_31953_n19727.n312 0.97759
R46428 a_31953_n19727.n97 a_31953_n19727.n310 0.97759
R46429 a_31953_n19727.n315 a_31953_n19727.n98 0.97759
R46430 a_31953_n19727.n99 a_31953_n19727.n313 0.97759
R46431 a_31953_n19727.n100 a_31953_n19727.n316 0.97759
R46432 a_31953_n19727.n102 a_31953_n19727.n314 0.97759
R46433 a_31953_n19727.n319 a_31953_n19727.n103 0.97759
R46434 a_31953_n19727.n104 a_31953_n19727.n317 0.97759
R46435 a_31953_n19727.n105 a_31953_n19727.n320 0.97759
R46436 a_31953_n19727.n106 a_31953_n19727.n318 0.97759
R46437 a_31953_n19727.n367 a_31953_n19727.n366 0.97759
R46438 a_31953_n19727.n368 a_31953_n19727.n364 0.97759
R46439 a_31953_n19727.n107 a_31953_n19727.n362 0.97759
R46440 a_31953_n19727.n109 a_31953_n19727.n360 0.97759
R46441 a_31953_n19727.n361 a_31953_n19727.n110 0.97759
R46442 a_31953_n19727.n111 a_31953_n19727.n359 0.97759
R46443 a_31953_n19727.n112 a_31953_n19727.n358 0.97759
R46444 a_31953_n19727.n114 a_31953_n19727.n356 0.97759
R46445 a_31953_n19727.n357 a_31953_n19727.n115 0.97759
R46446 a_31953_n19727.n116 a_31953_n19727.n355 0.97759
R46447 a_31953_n19727.n327 a_31953_n19727.n117 0.97759
R46448 a_31953_n19727.n118 a_31953_n19727.n325 0.97759
R46449 a_31953_n19727.n119 a_31953_n19727.n328 0.97759
R46450 a_31953_n19727.n120 a_31953_n19727.n326 0.97759
R46451 a_31953_n19727.n331 a_31953_n19727.n121 0.97759
R46452 a_31953_n19727.n122 a_31953_n19727.n329 0.97759
R46453 a_31953_n19727.n123 a_31953_n19727.n332 0.97759
R46454 a_31953_n19727.n125 a_31953_n19727.n330 0.97759
R46455 a_31953_n19727.n335 a_31953_n19727.n126 0.97759
R46456 a_31953_n19727.n127 a_31953_n19727.n333 0.97759
R46457 a_31953_n19727.n128 a_31953_n19727.n336 0.97759
R46458 a_31953_n19727.n129 a_31953_n19727.n334 0.97759
R46459 a_31953_n19727.n130 a_31953_n19727.n349 0.97759
R46460 a_31953_n19727.n132 a_31953_n19727.n347 0.97759
R46461 a_31953_n19727.n348 a_31953_n19727.n133 0.97759
R46462 a_31953_n19727.n134 a_31953_n19727.n346 0.97759
R46463 a_31953_n19727.n135 a_31953_n19727.n345 0.97759
R46464 a_31953_n19727.n136 a_31953_n19727.n343 0.97759
R46465 a_31953_n19727.n344 a_31953_n19727.n137 0.97759
R46466 a_31953_n19727.n138 a_31953_n19727.n342 0.97759
R46467 a_31953_n19727.n338 a_31953_n19727.n337 0.97759
R46468 a_31953_n19727.n139 a_31953_n19727.n341 0.97759
R46469 a_31953_n19727.n140 a_31953_n19727.n339 0.97759
R46470 a_31953_n19727.n141 a_31953_n19727.n340 0.97759
R46471 a_31953_n19727.n376 a_31953_n19727.n375 0.97759
R46472 a_31953_n19727.n377 a_31953_n19727.n373 0.97759
R46473 a_31953_n19727.n380 a_31953_n19727.n142 0.97759
R46474 a_31953_n19727.n143 a_31953_n19727.n378 0.97759
R46475 a_31953_n19727.n144 a_31953_n19727.n381 0.97759
R46476 a_31953_n19727.n146 a_31953_n19727.n379 0.97759
R46477 a_31953_n19727.n384 a_31953_n19727.n147 0.97759
R46478 a_31953_n19727.n148 a_31953_n19727.n382 0.97759
R46479 a_31953_n19727.n149 a_31953_n19727.n385 0.97759
R46480 a_31953_n19727.n150 a_31953_n19727.n383 0.97759
R46481 a_31953_n19727.n151 a_31953_n19727.n397 0.97759
R46482 a_31953_n19727.n153 a_31953_n19727.n395 0.97759
R46483 a_31953_n19727.n396 a_31953_n19727.n154 0.97759
R46484 a_31953_n19727.n155 a_31953_n19727.n394 0.97759
R46485 a_31953_n19727.n156 a_31953_n19727.n393 0.97759
R46486 a_31953_n19727.n157 a_31953_n19727.n391 0.97759
R46487 a_31953_n19727.n392 a_31953_n19727.n158 0.97759
R46488 a_31953_n19727.n159 a_31953_n19727.n390 0.97759
R46489 a_31953_n19727.n160 a_31953_n19727.n389 0.97759
R46490 a_31953_n19727.n162 a_31953_n19727.n387 0.97759
R46491 a_31953_n19727.n388 a_31953_n19727.n163 0.97759
R46492 a_31953_n19727.n164 a_31953_n19727.n386 0.97759
R46493 a_31953_n19727.n405 a_31953_n19727.n165 0.97759
R46494 a_31953_n19727.n166 a_31953_n19727.n403 0.97759
R46495 a_31953_n19727.n167 a_31953_n19727.n406 0.97759
R46496 a_31953_n19727.n168 a_31953_n19727.n404 0.97759
R46497 a_31953_n19727.n409 a_31953_n19727.n169 0.97759
R46498 a_31953_n19727.n170 a_31953_n19727.n407 0.97759
R46499 a_31953_n19727.n171 a_31953_n19727.n410 0.97759
R46500 a_31953_n19727.n173 a_31953_n19727.n408 0.97759
R46501 a_31953_n19727.n413 a_31953_n19727.n174 0.97759
R46502 a_31953_n19727.n175 a_31953_n19727.n411 0.97759
R46503 a_31953_n19727.n176 a_31953_n19727.n414 0.97759
R46504 a_31953_n19727.n177 a_31953_n19727.n412 0.97759
R46505 a_31953_n19727.n460 a_31953_n19727.n459 0.97759
R46506 a_31953_n19727.n461 a_31953_n19727.n457 0.97759
R46507 a_31953_n19727.n178 a_31953_n19727.n455 0.97759
R46508 a_31953_n19727.n180 a_31953_n19727.n453 0.97759
R46509 a_31953_n19727.n454 a_31953_n19727.n181 0.97759
R46510 a_31953_n19727.n182 a_31953_n19727.n452 0.97759
R46511 a_31953_n19727.n183 a_31953_n19727.n451 0.97759
R46512 a_31953_n19727.n185 a_31953_n19727.n449 0.97759
R46513 a_31953_n19727.n450 a_31953_n19727.n186 0.97759
R46514 a_31953_n19727.n187 a_31953_n19727.n448 0.97759
R46515 a_31953_n19727.n420 a_31953_n19727.n188 0.97759
R46516 a_31953_n19727.n189 a_31953_n19727.n418 0.97759
R46517 a_31953_n19727.n190 a_31953_n19727.n421 0.97759
R46518 a_31953_n19727.n191 a_31953_n19727.n419 0.97759
R46519 a_31953_n19727.n424 a_31953_n19727.n192 0.97759
R46520 a_31953_n19727.n193 a_31953_n19727.n422 0.97759
R46521 a_31953_n19727.n194 a_31953_n19727.n425 0.97759
R46522 a_31953_n19727.n196 a_31953_n19727.n423 0.97759
R46523 a_31953_n19727.n428 a_31953_n19727.n197 0.97759
R46524 a_31953_n19727.n198 a_31953_n19727.n426 0.97759
R46525 a_31953_n19727.n199 a_31953_n19727.n429 0.97759
R46526 a_31953_n19727.n200 a_31953_n19727.n427 0.97759
R46527 a_31953_n19727.n201 a_31953_n19727.n442 0.97759
R46528 a_31953_n19727.n203 a_31953_n19727.n440 0.97759
R46529 a_31953_n19727.n441 a_31953_n19727.n204 0.97759
R46530 a_31953_n19727.n205 a_31953_n19727.n439 0.97759
R46531 a_31953_n19727.n206 a_31953_n19727.n438 0.97759
R46532 a_31953_n19727.n207 a_31953_n19727.n436 0.97759
R46533 a_31953_n19727.n437 a_31953_n19727.n208 0.97759
R46534 a_31953_n19727.n209 a_31953_n19727.n435 0.97759
R46535 a_31953_n19727.n431 a_31953_n19727.n430 0.97759
R46536 a_31953_n19727.n210 a_31953_n19727.n434 0.97759
R46537 a_31953_n19727.n211 a_31953_n19727.n432 0.97759
R46538 a_31953_n19727.n212 a_31953_n19727.n433 0.97759
R46539 a_31953_n19727.n234 a_31953_n19727.n213 0.931516
R46540 a_31953_n19727.n214 a_31953_n19727.n232 0.931516
R46541 a_31953_n19727.n467 a_31953_n19727.n215 0.931516
R46542 a_31953_n19727.n216 a_31953_n19727.n465 0.931516
R46543 a_31953_n19727.n280 a_31953_n19727.n217 0.931516
R46544 a_31953_n19727.n218 a_31953_n19727.n278 0.931516
R46545 a_31953_n19727.n365 a_31953_n19727.n219 0.931516
R46546 a_31953_n19727.n220 a_31953_n19727.n363 0.931516
R46547 a_31953_n19727.n374 a_31953_n19727.n221 0.931516
R46548 a_31953_n19727.n222 a_31953_n19727.n372 0.931516
R46549 a_31953_n19727.n458 a_31953_n19727.n223 0.931516
R46550 a_31953_n19727.n224 a_31953_n19727.n456 0.931516
R46551 a_31953_n19727.n74 a_31953_n19727.n81 0.82023
R46552 a_31953_n19727.n145 a_31953_n19727.n152 0.82023
R46553 a_31953_n19727.n3 a_31953_n19727.n10 0.82023
R46554 a_31953_n19727.n131 a_31953_n19727.n124 0.818405
R46555 a_31953_n19727.n202 a_31953_n19727.n195 0.818405
R46556 a_31953_n19727.n60 a_31953_n19727.n53 0.818405
R46557 a_31953_n19727.n463 a_31953_n19727.n462 0.7505
R46558 a_31953_n19727.n462 a_31953_n19727.n172 0.717155
R46559 a_31953_n19727.n464 a_31953_n19727.n30 0.717155
R46560 a_31953_n19727.n226 a_31953_n19727.n101 0.711725
R46561 a_31953_n19727.n108 a_31953_n19727.n113 0.639622
R46562 a_31953_n19727.n179 a_31953_n19727.n184 0.639622
R46563 a_31953_n19727.n48 a_31953_n19727.n39 0.639622
R46564 a_31953_n19727.n237 a_31953_n19727.n236 0.62434
R46565 a_31953_n19727.n470 a_31953_n19727.n469 0.62434
R46566 a_31953_n19727.n283 a_31953_n19727.n282 0.62434
R46567 a_31953_n19727.n368 a_31953_n19727.n367 0.62434
R46568 a_31953_n19727.n377 a_31953_n19727.n376 0.62434
R46569 a_31953_n19727.n461 a_31953_n19727.n460 0.62434
R46570 a_31953_n19727.n212 a_31953_n19727.n211 0.62434
R46571 a_31953_n19727.n430 a_31953_n19727.n210 0.62434
R46572 a_31953_n19727.n209 a_31953_n19727.n208 0.62434
R46573 a_31953_n19727.n207 a_31953_n19727.n206 0.62434
R46574 a_31953_n19727.n205 a_31953_n19727.n204 0.62434
R46575 a_31953_n19727.n203 a_31953_n19727.n201 0.62434
R46576 a_31953_n19727.n200 a_31953_n19727.n199 0.62434
R46577 a_31953_n19727.n198 a_31953_n19727.n197 0.62434
R46578 a_31953_n19727.n196 a_31953_n19727.n194 0.62434
R46579 a_31953_n19727.n193 a_31953_n19727.n192 0.62434
R46580 a_31953_n19727.n191 a_31953_n19727.n190 0.62434
R46581 a_31953_n19727.n189 a_31953_n19727.n188 0.62434
R46582 a_31953_n19727.n187 a_31953_n19727.n186 0.62434
R46583 a_31953_n19727.n185 a_31953_n19727.n183 0.62434
R46584 a_31953_n19727.n182 a_31953_n19727.n181 0.62434
R46585 a_31953_n19727.n180 a_31953_n19727.n178 0.62434
R46586 a_31953_n19727.n177 a_31953_n19727.n176 0.62434
R46587 a_31953_n19727.n175 a_31953_n19727.n174 0.62434
R46588 a_31953_n19727.n173 a_31953_n19727.n171 0.62434
R46589 a_31953_n19727.n170 a_31953_n19727.n169 0.62434
R46590 a_31953_n19727.n168 a_31953_n19727.n167 0.62434
R46591 a_31953_n19727.n166 a_31953_n19727.n165 0.62434
R46592 a_31953_n19727.n164 a_31953_n19727.n163 0.62434
R46593 a_31953_n19727.n162 a_31953_n19727.n160 0.62434
R46594 a_31953_n19727.n159 a_31953_n19727.n158 0.62434
R46595 a_31953_n19727.n157 a_31953_n19727.n156 0.62434
R46596 a_31953_n19727.n155 a_31953_n19727.n154 0.62434
R46597 a_31953_n19727.n153 a_31953_n19727.n151 0.62434
R46598 a_31953_n19727.n150 a_31953_n19727.n149 0.62434
R46599 a_31953_n19727.n148 a_31953_n19727.n147 0.62434
R46600 a_31953_n19727.n146 a_31953_n19727.n144 0.62434
R46601 a_31953_n19727.n143 a_31953_n19727.n142 0.62434
R46602 a_31953_n19727.n141 a_31953_n19727.n140 0.62434
R46603 a_31953_n19727.n337 a_31953_n19727.n139 0.62434
R46604 a_31953_n19727.n138 a_31953_n19727.n137 0.62434
R46605 a_31953_n19727.n136 a_31953_n19727.n135 0.62434
R46606 a_31953_n19727.n134 a_31953_n19727.n133 0.62434
R46607 a_31953_n19727.n132 a_31953_n19727.n130 0.62434
R46608 a_31953_n19727.n129 a_31953_n19727.n128 0.62434
R46609 a_31953_n19727.n127 a_31953_n19727.n126 0.62434
R46610 a_31953_n19727.n125 a_31953_n19727.n123 0.62434
R46611 a_31953_n19727.n122 a_31953_n19727.n121 0.62434
R46612 a_31953_n19727.n120 a_31953_n19727.n119 0.62434
R46613 a_31953_n19727.n118 a_31953_n19727.n117 0.62434
R46614 a_31953_n19727.n116 a_31953_n19727.n115 0.62434
R46615 a_31953_n19727.n114 a_31953_n19727.n112 0.62434
R46616 a_31953_n19727.n111 a_31953_n19727.n110 0.62434
R46617 a_31953_n19727.n109 a_31953_n19727.n107 0.62434
R46618 a_31953_n19727.n106 a_31953_n19727.n105 0.62434
R46619 a_31953_n19727.n104 a_31953_n19727.n103 0.62434
R46620 a_31953_n19727.n102 a_31953_n19727.n100 0.62434
R46621 a_31953_n19727.n99 a_31953_n19727.n98 0.62434
R46622 a_31953_n19727.n97 a_31953_n19727.n96 0.62434
R46623 a_31953_n19727.n95 a_31953_n19727.n94 0.62434
R46624 a_31953_n19727.n93 a_31953_n19727.n92 0.62434
R46625 a_31953_n19727.n91 a_31953_n19727.n89 0.62434
R46626 a_31953_n19727.n88 a_31953_n19727.n87 0.62434
R46627 a_31953_n19727.n86 a_31953_n19727.n85 0.62434
R46628 a_31953_n19727.n84 a_31953_n19727.n83 0.62434
R46629 a_31953_n19727.n82 a_31953_n19727.n80 0.62434
R46630 a_31953_n19727.n79 a_31953_n19727.n78 0.62434
R46631 a_31953_n19727.n77 a_31953_n19727.n76 0.62434
R46632 a_31953_n19727.n75 a_31953_n19727.n73 0.62434
R46633 a_31953_n19727.n72 a_31953_n19727.n71 0.62434
R46634 a_31953_n19727.n70 a_31953_n19727.n69 0.62434
R46635 a_31953_n19727.n495 a_31953_n19727.n68 0.62434
R46636 a_31953_n19727.n67 a_31953_n19727.n66 0.62434
R46637 a_31953_n19727.n65 a_31953_n19727.n64 0.62434
R46638 a_31953_n19727.n63 a_31953_n19727.n62 0.62434
R46639 a_31953_n19727.n61 a_31953_n19727.n59 0.62434
R46640 a_31953_n19727.n58 a_31953_n19727.n57 0.62434
R46641 a_31953_n19727.n56 a_31953_n19727.n55 0.62434
R46642 a_31953_n19727.n54 a_31953_n19727.n52 0.62434
R46643 a_31953_n19727.n51 a_31953_n19727.n50 0.62434
R46644 a_31953_n19727.n49 a_31953_n19727.n47 0.62434
R46645 a_31953_n19727.n46 a_31953_n19727.n45 0.62434
R46646 a_31953_n19727.n44 a_31953_n19727.n43 0.62434
R46647 a_31953_n19727.n42 a_31953_n19727.n41 0.62434
R46648 a_31953_n19727.n40 a_31953_n19727.n38 0.62434
R46649 a_31953_n19727.n37 a_31953_n19727.n36 0.62434
R46650 a_31953_n19727.n35 a_31953_n19727.n34 0.62434
R46651 a_31953_n19727.n33 a_31953_n19727.n32 0.62434
R46652 a_31953_n19727.n31 a_31953_n19727.n29 0.62434
R46653 a_31953_n19727.n28 a_31953_n19727.n27 0.62434
R46654 a_31953_n19727.n26 a_31953_n19727.n25 0.62434
R46655 a_31953_n19727.n24 a_31953_n19727.n23 0.62434
R46656 a_31953_n19727.n22 a_31953_n19727.n21 0.62434
R46657 a_31953_n19727.n20 a_31953_n19727.n18 0.62434
R46658 a_31953_n19727.n17 a_31953_n19727.n16 0.62434
R46659 a_31953_n19727.n15 a_31953_n19727.n14 0.62434
R46660 a_31953_n19727.n13 a_31953_n19727.n12 0.62434
R46661 a_31953_n19727.n11 a_31953_n19727.n9 0.62434
R46662 a_31953_n19727.n8 a_31953_n19727.n7 0.62434
R46663 a_31953_n19727.n6 a_31953_n19727.n5 0.62434
R46664 a_31953_n19727.n4 a_31953_n19727.n2 0.62434
R46665 a_31953_n19727.n1 a_31953_n19727.n0 0.62434
R46666 a_31953_n19727.n462 a_31953_n19727.n179 0.617426
R46667 a_31953_n19727.n39 a_31953_n19727.n464 0.617426
R46668 a_31953_n19727.n225 a_31953_n19727.n108 0.604351
R46669 a_31953_n19727.n224 a_31953_n19727.n223 0.595087
R46670 a_31953_n19727.n222 a_31953_n19727.n221 0.595087
R46671 a_31953_n19727.n220 a_31953_n19727.n219 0.595087
R46672 a_31953_n19727.n218 a_31953_n19727.n217 0.595087
R46673 a_31953_n19727.n216 a_31953_n19727.n215 0.595087
R46674 a_31953_n19727.n214 a_31953_n19727.n213 0.595087
R46675 a_31953_n19727.n124 a_31953_n19727.n113 0.545973
R46676 a_31953_n19727.n195 a_31953_n19727.n184 0.545973
R46677 a_31953_n19727.n53 a_31953_n19727.n48 0.545973
R46678 a_31953_n19727.n81 a_31953_n19727.n90 0.545365
R46679 a_31953_n19727.n152 a_31953_n19727.n161 0.545365
R46680 a_31953_n19727.n10 a_31953_n19727.n19 0.545365
R46681 a_31953_n19727.n30 a_31953_n19727.n19 0.452324
R46682 a_31953_n19727.n172 a_31953_n19727.n161 0.452324
R46683 a_31953_n19727.n101 a_31953_n19727.n90 0.452324
R46684 a_31699_20742.n388 a_31699_20742.n313 16.7377
R46685 a_31699_20742.n314 a_31699_20742.t1 10.214
R46686 a_31699_20742.n324 a_31699_20742.t131 10.214
R46687 a_31699_20742.n335 a_31699_20742.t220 10.214
R46688 a_31699_20742.n346 a_31699_20742.t60 10.214
R46689 a_31699_20742.n356 a_31699_20742.t141 10.214
R46690 a_31699_20742.n320 a_31699_20742.t27 10.2117
R46691 a_31699_20742.n330 a_31699_20742.t213 10.2117
R46692 a_31699_20742.n341 a_31699_20742.t81 10.2117
R46693 a_31699_20742.n352 a_31699_20742.t143 10.2117
R46694 a_31699_20742.n362 a_31699_20742.t224 10.2117
R46695 a_31699_20742.n317 a_31699_20742.t185 9.58832
R46696 a_31699_20742.n327 a_31699_20742.t52 9.58832
R46697 a_31699_20742.n338 a_31699_20742.t23 9.58832
R46698 a_31699_20742.n370 a_31699_20742.t144 9.58832
R46699 a_31699_20742.n349 a_31699_20742.t17 9.58832
R46700 a_31699_20742.n359 a_31699_20742.t62 9.58832
R46701 a_31699_20742.n319 a_31699_20742.t89 9.58085
R46702 a_31699_20742.n329 a_31699_20742.t172 9.58085
R46703 a_31699_20742.n340 a_31699_20742.t3 9.58085
R46704 a_31699_20742.n372 a_31699_20742.t45 9.58085
R46705 a_31699_20742.n351 a_31699_20742.t29 9.58085
R46706 a_31699_20742.n361 a_31699_20742.t184 9.58085
R46707 a_31699_20742.n318 a_31699_20742.t256 9.58045
R46708 a_31699_20742.n316 a_31699_20742.t37 9.58045
R46709 a_31699_20742.n315 a_31699_20742.t7 9.58045
R46710 a_31699_20742.n328 a_31699_20742.t127 9.58045
R46711 a_31699_20742.n326 a_31699_20742.t153 9.58045
R46712 a_31699_20742.n325 a_31699_20742.t108 9.58045
R46713 a_31699_20742.n339 a_31699_20742.t13 9.58045
R46714 a_31699_20742.n337 a_31699_20742.t244 9.58045
R46715 a_31699_20742.n336 a_31699_20742.t199 9.58045
R46716 a_31699_20742.n371 a_31699_20742.t219 9.58045
R46717 a_31699_20742.n350 a_31699_20742.t39 9.58045
R46718 a_31699_20742.n348 a_31699_20742.t85 9.58045
R46719 a_31699_20742.n347 a_31699_20742.t255 9.58045
R46720 a_31699_20742.n360 a_31699_20742.t134 9.58045
R46721 a_31699_20742.n358 a_31699_20742.t164 9.58045
R46722 a_31699_20742.n357 a_31699_20742.t118 9.58045
R46723 a_31699_20742.n314 a_31699_20742.t33 9.58005
R46724 a_31699_20742.n324 a_31699_20742.t180 9.58005
R46725 a_31699_20742.n335 a_31699_20742.t46 9.58005
R46726 a_31699_20742.n346 a_31699_20742.t111 9.58005
R46727 a_31699_20742.n356 a_31699_20742.t192 9.58005
R46728 a_31699_20742.n320 a_31699_20742.t41 9.57886
R46729 a_31699_20742.n321 a_31699_20742.t15 9.57886
R46730 a_31699_20742.n322 a_31699_20742.t25 9.57886
R46731 a_31699_20742.n330 a_31699_20742.t138 9.57886
R46732 a_31699_20742.n331 a_31699_20742.t72 9.57886
R46733 a_31699_20742.n332 a_31699_20742.t218 9.57886
R46734 a_31699_20742.n341 a_31699_20742.t234 9.57886
R46735 a_31699_20742.n342 a_31699_20742.t163 9.57886
R46736 a_31699_20742.n343 a_31699_20742.t92 9.57886
R46737 a_31699_20742.n352 a_31699_20742.t71 9.57886
R46738 a_31699_20742.n353 a_31699_20742.t226 9.57886
R46739 a_31699_20742.n354 a_31699_20742.t150 9.57886
R46740 a_31699_20742.n362 a_31699_20742.t149 9.57886
R46741 a_31699_20742.n363 a_31699_20742.t82 9.57886
R46742 a_31699_20742.n364 a_31699_20742.t235 9.57886
R46743 a_31699_20742.n376 a_31699_20742.t35 8.38951
R46744 a_31699_20742.n389 a_31699_20742.t0 8.38805
R46745 a_31699_20742.n367 a_31699_20742.t11 8.38752
R46746 a_31699_20742.n268 a_31699_20742.t142 8.38704
R46747 a_31699_20742.n262 a_31699_20742.t207 8.38704
R46748 a_31699_20742.n211 a_31699_20742.t242 8.46135
R46749 a_31699_20742.n213 a_31699_20742.t148 8.46135
R46750 a_31699_20742.n193 a_31699_20742.t69 8.48081
R46751 a_31699_20742.n188 a_31699_20742.t228 8.48081
R46752 a_31699_20742.n168 a_31699_20742.t156 8.10567
R46753 a_31699_20742.n130 a_31699_20742.t51 8.10567
R46754 a_31699_20742.n130 a_31699_20742.t223 8.10567
R46755 a_31699_20742.n131 a_31699_20742.t147 8.10567
R46756 a_31699_20742.n131 a_31699_20742.t222 8.10567
R46757 a_31699_20742.n113 a_31699_20742.t87 8.10567
R46758 a_31699_20742.n113 a_31699_20742.t237 8.10567
R46759 a_31699_20742.n127 a_31699_20742.t162 8.10567
R46760 a_31699_20742.n127 a_31699_20742.t94 8.10567
R46761 a_31699_20742.n110 a_31699_20742.t70 8.10567
R46762 a_31699_20742.n110 a_31699_20742.t217 8.10567
R46763 a_31699_20742.n124 a_31699_20742.t166 8.10567
R46764 a_31699_20742.n124 a_31699_20742.t75 8.10567
R46765 a_31699_20742.n173 a_31699_20742.t73 8.10567
R46766 a_31699_20742.n173 a_31699_20742.t201 8.10567
R46767 a_31699_20742.n219 a_31699_20742.t128 8.10567
R46768 a_31699_20742.n176 a_31699_20742.t124 8.10567
R46769 a_31699_20742.n176 a_31699_20742.t221 8.10567
R46770 a_31699_20742.n175 a_31699_20742.t146 8.10567
R46771 a_31699_20742.n168 a_31699_20742.t90 8.10567
R46772 a_31699_20742.n136 a_31699_20742.t238 8.10567
R46773 a_31699_20742.n136 a_31699_20742.t187 8.10567
R46774 a_31699_20742.n90 a_31699_20742.t145 8.10567
R46775 a_31699_20742.n158 a_31699_20742.t258 8.10567
R46776 a_31699_20742.n158 a_31699_20742.t216 8.10567
R46777 a_31699_20742.n159 a_31699_20742.t139 8.10567
R46778 a_31699_20742.n159 a_31699_20742.t214 8.10567
R46779 a_31699_20742.n83 a_31699_20742.t76 8.10567
R46780 a_31699_20742.n83 a_31699_20742.t227 8.10567
R46781 a_31699_20742.n162 a_31699_20742.t151 8.10567
R46782 a_31699_20742.n162 a_31699_20742.t84 8.10567
R46783 a_31699_20742.n87 a_31699_20742.t59 8.10567
R46784 a_31699_20742.n87 a_31699_20742.t209 8.10567
R46785 a_31699_20742.n86 a_31699_20742.t161 8.10567
R46786 a_31699_20742.n86 a_31699_20742.t66 8.10567
R46787 a_31699_20742.n198 a_31699_20742.t247 8.10567
R46788 a_31699_20742.n198 a_31699_20742.t154 8.10567
R46789 a_31699_20742.n226 a_31699_20742.t78 8.10567
R46790 a_31699_20742.n201 a_31699_20742.t74 8.10567
R46791 a_31699_20742.n201 a_31699_20742.t174 8.10567
R46792 a_31699_20742.n200 a_31699_20742.t100 8.10567
R46793 a_31699_20742.n90 a_31699_20742.t77 8.10567
R46794 a_31699_20742.n90 a_31699_20742.t230 8.10567
R46795 a_31699_20742.n90 a_31699_20742.t181 8.10567
R46796 a_31699_20742.n165 a_31699_20742.t93 8.10567
R46797 a_31699_20742.n120 a_31699_20742.t205 8.10567
R46798 a_31699_20742.n120 a_31699_20742.t159 8.10567
R46799 a_31699_20742.n121 a_31699_20742.t86 8.10567
R46800 a_31699_20742.n121 a_31699_20742.t158 8.10567
R46801 a_31699_20742.n107 a_31699_20742.t243 8.10567
R46802 a_31699_20742.n107 a_31699_20742.t168 8.10567
R46803 a_31699_20742.n106 a_31699_20742.t97 8.10567
R46804 a_31699_20742.n106 a_31699_20742.t249 8.10567
R46805 a_31699_20742.n103 a_31699_20742.t229 8.10567
R46806 a_31699_20742.n103 a_31699_20742.t152 8.10567
R46807 a_31699_20742.n102 a_31699_20742.t106 8.10567
R46808 a_31699_20742.n102 a_31699_20742.t236 8.10567
R46809 a_31699_20742.n179 a_31699_20742.t233 8.10567
R46810 a_31699_20742.n179 a_31699_20742.t136 8.10567
R46811 a_31699_20742.n178 a_31699_20742.t63 8.10567
R46812 a_31699_20742.n182 a_31699_20742.t56 8.10567
R46813 a_31699_20742.n182 a_31699_20742.t157 8.10567
R46814 a_31699_20742.n181 a_31699_20742.t83 8.10567
R46815 a_31699_20742.n165 a_31699_20742.t245 8.10567
R46816 a_31699_20742.n134 a_31699_20742.t170 8.10567
R46817 a_31699_20742.n134 a_31699_20742.t125 8.10567
R46818 a_31699_20742.n100 a_31699_20742.t54 8.10567
R46819 a_31699_20742.n214 a_31699_20742.t167 8.10567
R46820 a_31699_20742.n214 a_31699_20742.t123 8.10567
R46821 a_31699_20742.n153 a_31699_20742.t49 8.10567
R46822 a_31699_20742.n153 a_31699_20742.t122 8.10567
R46823 a_31699_20742.n93 a_31699_20742.t206 8.10567
R46824 a_31699_20742.n93 a_31699_20742.t133 8.10567
R46825 a_31699_20742.n92 a_31699_20742.t57 8.10567
R46826 a_31699_20742.n92 a_31699_20742.t215 8.10567
R46827 a_31699_20742.n97 a_31699_20742.t193 8.10567
R46828 a_31699_20742.n97 a_31699_20742.t117 8.10567
R46829 a_31699_20742.n96 a_31699_20742.t68 8.10567
R46830 a_31699_20742.n96 a_31699_20742.t200 8.10567
R46831 a_31699_20742.n204 a_31699_20742.t155 8.10567
R46832 a_31699_20742.n204 a_31699_20742.t61 8.10567
R46833 a_31699_20742.n203 a_31699_20742.t211 8.10567
R46834 a_31699_20742.n206 a_31699_20742.t203 8.10567
R46835 a_31699_20742.n206 a_31699_20742.t80 8.10567
R46836 a_31699_20742.n230 a_31699_20742.t232 8.10567
R46837 a_31699_20742.n100 a_31699_20742.t210 8.10567
R46838 a_31699_20742.n100 a_31699_20742.t135 8.10567
R46839 a_31699_20742.n100 a_31699_20742.t88 8.10567
R46840 a_31699_20742.n49 a_31699_20742.t107 8.10567
R46841 a_31699_20742.n47 a_31699_20742.t252 8.10567
R46842 a_31699_20742.n45 a_31699_20742.t182 8.10567
R46843 a_31699_20742.n260 a_31699_20742.t113 8.10567
R46844 a_31699_20742.n307 a_31699_20742.t53 8.10567
R46845 a_31699_20742.n306 a_31699_20742.t183 8.10567
R46846 a_31699_20742.n305 a_31699_20742.t110 8.10567
R46847 a_31699_20742.n192 a_31699_20742.t241 8.10567
R46848 a_31699_20742.n43 a_31699_20742.t165 8.10567
R46849 a_31699_20742.n41 a_31699_20742.t240 8.10567
R46850 a_31699_20742.n59 a_31699_20742.t176 8.10567
R46851 a_31699_20742.n57 a_31699_20742.t109 8.10567
R46852 a_31699_20742.n261 a_31699_20742.t253 8.10567
R46853 a_31699_20742.n301 a_31699_20742.t104 8.10567
R46854 a_31699_20742.n300 a_31699_20742.t202 8.10567
R46855 a_31699_20742.n299 a_31699_20742.t130 8.10567
R46856 a_31699_20742.n190 a_31699_20742.t91 8.10567
R46857 a_31699_20742.n55 a_31699_20742.t239 8.10567
R46858 a_31699_20742.n53 a_31699_20742.t188 8.10567
R46859 a_31699_20742.n52 a_31699_20742.t96 8.10567
R46860 a_31699_20742.n0 a_31699_20742.t55 8.10567
R46861 a_31699_20742.n1 a_31699_20742.t204 8.10567
R46862 a_31699_20742.n18 a_31699_20742.t132 8.10567
R46863 a_31699_20742.n144 a_31699_20742.t65 8.10567
R46864 a_31699_20742.n279 a_31699_20742.t264 8.10567
R46865 a_31699_20742.n278 a_31699_20742.t173 8.10567
R46866 a_31699_20742.n277 a_31699_20742.t99 8.10567
R46867 a_31699_20742.n210 a_31699_20742.t198 8.10567
R46868 a_31699_20742.n16 a_31699_20742.t121 8.10567
R46869 a_31699_20742.n28 a_31699_20742.t196 8.10567
R46870 a_31699_20742.n37 a_31699_20742.t129 8.10567
R46871 a_31699_20742.n5 a_31699_20742.t58 8.10567
R46872 a_31699_20742.n141 a_31699_20742.t208 8.10567
R46873 a_31699_20742.n276 a_31699_20742.t95 8.10567
R46874 a_31699_20742.n275 a_31699_20742.t195 8.10567
R46875 a_31699_20742.n274 a_31699_20742.t120 8.10567
R46876 a_31699_20742.n147 a_31699_20742.t260 8.10567
R46877 a_31699_20742.n3 a_31699_20742.t189 8.10567
R46878 a_31699_20742.n20 a_31699_20742.t140 8.10567
R46879 a_31699_20742.n30 a_31699_20742.t47 8.10567
R46880 a_31699_20742.n69 a_31699_20742.t261 8.10567
R46881 a_31699_20742.n67 a_31699_20742.t190 8.10567
R46882 a_31699_20742.n65 a_31699_20742.t115 8.10567
R46883 a_31699_20742.n286 a_31699_20742.t48 8.10567
R46884 a_31699_20742.n282 a_31699_20742.t212 8.10567
R46885 a_31699_20742.n283 a_31699_20742.t119 8.10567
R46886 a_31699_20742.n284 a_31699_20742.t263 8.10567
R46887 a_31699_20742.n189 a_31699_20742.t179 8.10567
R46888 a_31699_20742.n63 a_31699_20742.t105 8.10567
R46889 a_31699_20742.n61 a_31699_20742.t177 8.10567
R46890 a_31699_20742.n79 a_31699_20742.t112 8.10567
R46891 a_31699_20742.n77 a_31699_20742.t262 8.10567
R46892 a_31699_20742.n267 a_31699_20742.t194 8.10567
R46893 a_31699_20742.n272 a_31699_20742.t257 8.10567
R46894 a_31699_20742.n271 a_31699_20742.t137 8.10567
R46895 a_31699_20742.n270 a_31699_20742.t64 8.10567
R46896 a_31699_20742.n186 a_31699_20742.t246 8.10567
R46897 a_31699_20742.n75 a_31699_20742.t171 8.10567
R46898 a_31699_20742.n73 a_31699_20742.t126 8.10567
R46899 a_31699_20742.n71 a_31699_20742.t251 8.10567
R46900 a_31699_20742.n7 a_31699_20742.t186 8.10567
R46901 a_31699_20742.n8 a_31699_20742.t114 8.10567
R46902 a_31699_20742.n24 a_31699_20742.t259 8.10567
R46903 a_31699_20742.n142 a_31699_20742.t197 8.10567
R46904 a_31699_20742.n293 a_31699_20742.t175 8.10567
R46905 a_31699_20742.n294 a_31699_20742.t79 8.10567
R46906 a_31699_20742.n295 a_31699_20742.t231 8.10567
R46907 a_31699_20742.n212 a_31699_20742.t103 8.10567
R46908 a_31699_20742.n22 a_31699_20742.t250 8.10567
R46909 a_31699_20742.n32 a_31699_20742.t102 8.10567
R46910 a_31699_20742.n13 a_31699_20742.t254 8.10567
R46911 a_31699_20742.n14 a_31699_20742.t191 8.10567
R46912 a_31699_20742.n138 a_31699_20742.t116 8.10567
R46913 a_31699_20742.n291 a_31699_20742.t225 8.10567
R46914 a_31699_20742.n290 a_31699_20742.t101 8.10567
R46915 a_31699_20742.n289 a_31699_20742.t248 8.10567
R46916 a_31699_20742.n10 a_31699_20742.t169 8.10567
R46917 a_31699_20742.n11 a_31699_20742.t98 8.10567
R46918 a_31699_20742.n26 a_31699_20742.t50 8.10567
R46919 a_31699_20742.n34 a_31699_20742.t178 8.10567
R46920 a_31699_20742.n377 a_31699_20742.t9 8.10567
R46921 a_31699_20742.n382 a_31699_20742.t21 8.10567
R46922 a_31699_20742.n373 a_31699_20742.t31 8.10567
R46923 a_31699_20742.n184 a_31699_20742.t5 8.10567
R46924 a_31699_20742.n81 a_31699_20742.t19 8.10567
R46925 a_31699_20742.n366 a_31699_20742.t43 8.10567
R46926 a_31699_20742.n244 a_31699_20742.t2 6.61324
R46927 a_31699_20742.n241 a_31699_20742.t12 6.57135
R46928 a_31699_20742.n246 a_31699_20742.t26 5.34147
R46929 a_31699_20742.n245 a_31699_20742.t38 5.34147
R46930 a_31699_20742.n191 a_31699_20742.n190 1.45673
R46931 a_31699_20742.n187 a_31699_20742.n186 1.45673
R46932 a_31699_20742.n185 a_31699_20742.n184 1.45673
R46933 a_31699_20742.n148 a_31699_20742.n147 1.45418
R46934 a_31699_20742.n146 a_31699_20742.n10 1.45418
R46935 a_31699_20742.n145 a_31699_20742.n144 1.45392
R46936 a_31699_20742.n143 a_31699_20742.n142 1.45392
R46937 a_31699_20742.n242 a_31699_20742.n235 3.82989
R46938 a_31699_20742.n241 a_31699_20742.n391 3.82989
R46939 a_31699_20742.n234 a_31699_20742.n235 0.0670308
R46940 a_31699_20742.n233 a_31699_20742.t32 5.29989
R46941 a_31699_20742.n232 a_31699_20742.t6 5.29989
R46942 a_31699_20742.n174 a_31699_20742.n173 0.592804
R46943 a_31699_20742.n177 a_31699_20742.n176 0.592804
R46944 a_31699_20742.n180 a_31699_20742.n179 0.592804
R46945 a_31699_20742.n183 a_31699_20742.n182 0.592804
R46946 a_31699_20742.n199 a_31699_20742.n198 0.592738
R46947 a_31699_20742.n202 a_31699_20742.n201 0.592738
R46948 a_31699_20742.n205 a_31699_20742.n204 0.592738
R46949 a_31699_20742.n206 a_31699_20742.n207 0.592738
R46950 a_31699_20742.n159 a_31699_20742.n161 0.591918
R46951 a_31699_20742.n164 a_31699_20742.n162 0.591918
R46952 a_31699_20742.n157 a_31699_20742.n86 0.591918
R46953 a_31699_20742.n155 a_31699_20742.n153 0.591918
R46954 a_31699_20742.n152 a_31699_20742.n92 0.591918
R46955 a_31699_20742.n96 a_31699_20742.n150 0.591918
R46956 a_31699_20742.n83 a_31699_20742.n84 0.591886
R46957 a_31699_20742.n87 a_31699_20742.n88 0.591826
R46958 a_31699_20742.n90 a_31699_20742.n91 0.067621
R46959 a_31699_20742.n93 a_31699_20742.n94 0.591826
R46960 a_31699_20742.n98 a_31699_20742.n97 0.591886
R46961 a_31699_20742.n101 a_31699_20742.n100 0.0676312
R46962 a_31699_20742.n240 a_31699_20742.n239 1.46537
R46963 a_31699_20742.n110 a_31699_20742.n112 0.604258
R46964 a_31699_20742.n124 a_31699_20742.n125 0.591264
R46965 a_31699_20742.n113 a_31699_20742.n115 0.604258
R46966 a_31699_20742.n128 a_31699_20742.n127 0.591264
R46967 a_31699_20742.n132 a_31699_20742.n131 0.591264
R46968 a_31699_20742.n169 a_31699_20742.n168 0.604258
R46969 a_31699_20742.n136 a_31699_20742.n137 0.031901
R46970 a_31699_20742.n86 a_31699_20742.n156 0.591264
R46971 a_31699_20742.n89 a_31699_20742.n87 0.604195
R46972 a_31699_20742.n162 a_31699_20742.n163 0.591264
R46973 a_31699_20742.n83 a_31699_20742.n85 0.604258
R46974 a_31699_20742.n160 a_31699_20742.n159 0.591264
R46975 a_31699_20742.n216 a_31699_20742.n158 0.0732126
R46976 a_31699_20742.n105 a_31699_20742.n103 0.604258
R46977 a_31699_20742.n102 a_31699_20742.n116 0.591264
R46978 a_31699_20742.n109 a_31699_20742.n107 0.604258
R46979 a_31699_20742.n106 a_31699_20742.n118 0.591264
R46980 a_31699_20742.n121 a_31699_20742.n122 0.591264
R46981 a_31699_20742.n166 a_31699_20742.n165 0.604258
R46982 a_31699_20742.n134 a_31699_20742.n135 0.031901
R46983 a_31699_20742.n165 a_31699_20742.n167 0.604258
R46984 a_31699_20742.n117 a_31699_20742.n102 0.591264
R46985 a_31699_20742.n103 a_31699_20742.n104 0.604258
R46986 a_31699_20742.n119 a_31699_20742.n106 0.591264
R46987 a_31699_20742.n107 a_31699_20742.n108 0.604258
R46988 a_31699_20742.n123 a_31699_20742.n121 0.591264
R46989 a_31699_20742.n120 a_31699_20742.n171 0.0301596
R46990 a_31699_20742.n149 a_31699_20742.n96 0.591264
R46991 a_31699_20742.n97 a_31699_20742.n99 0.604258
R46992 a_31699_20742.n92 a_31699_20742.n151 0.591264
R46993 a_31699_20742.n95 a_31699_20742.n93 0.604195
R46994 a_31699_20742.n153 a_31699_20742.n154 0.591264
R46995 a_31699_20742.n214 a_31699_20742.n215 0.0732126
R46996 a_31699_20742.n168 a_31699_20742.n170 0.604258
R46997 a_31699_20742.n126 a_31699_20742.n124 0.591264
R46998 a_31699_20742.n111 a_31699_20742.n110 0.604258
R46999 a_31699_20742.n127 a_31699_20742.n129 0.591264
R47000 a_31699_20742.n114 a_31699_20742.n113 0.604258
R47001 a_31699_20742.n131 a_31699_20742.n133 0.591264
R47002 a_31699_20742.n130 a_31699_20742.n172 0.0301596
R47003 a_31699_20742.n141 a_31699_20742.n140 0.359454
R47004 a_31699_20742.n5 a_31699_20742.n6 1.44113
R47005 a_31699_20742.n37 a_31699_20742.n38 1.44113
R47006 a_31699_20742.n31 a_31699_20742.n30 1.44113
R47007 a_31699_20742.n21 a_31699_20742.n20 1.44113
R47008 a_31699_20742.n3 a_31699_20742.n4 1.44113
R47009 a_31699_20742.n18 a_31699_20742.n19 1.44113
R47010 a_31699_20742.n1 a_31699_20742.n2 1.44113
R47011 a_31699_20742.n0 a_31699_20742.n36 1.44113
R47012 a_31699_20742.n29 a_31699_20742.n28 1.44113
R47013 a_31699_20742.n17 a_31699_20742.n16 1.44113
R47014 a_31699_20742.n210 a_31699_20742.n211 0.332154
R47015 a_31699_20742.n79 a_31699_20742.n80 1.44113
R47016 a_31699_20742.n78 a_31699_20742.n77 1.44113
R47017 a_31699_20742.n269 a_31699_20742.n266 4.5005
R47018 a_31699_20742.n72 a_31699_20742.n71 1.44113
R47019 a_31699_20742.n73 a_31699_20742.n74 1.44113
R47020 a_31699_20742.n76 a_31699_20742.n75 1.44113
R47021 a_31699_20742.n70 a_31699_20742.n69 1.44113
R47022 a_31699_20742.n68 a_31699_20742.n67 1.44113
R47023 a_31699_20742.n66 a_31699_20742.n65 1.44113
R47024 a_31699_20742.n285 a_31699_20742.n273 4.5005
R47025 a_31699_20742.n61 a_31699_20742.n62 1.44113
R47026 a_31699_20742.n64 a_31699_20742.n63 1.44113
R47027 a_31699_20742.n189 a_31699_20742.n188 0.349872
R47028 a_31699_20742.n139 a_31699_20742.n138 0.359454
R47029 a_31699_20742.n15 a_31699_20742.n14 1.44113
R47030 a_31699_20742.n13 a_31699_20742.n40 1.44113
R47031 a_31699_20742.n35 a_31699_20742.n34 1.44113
R47032 a_31699_20742.n27 a_31699_20742.n26 1.44113
R47033 a_31699_20742.n11 a_31699_20742.n12 1.44113
R47034 a_31699_20742.n25 a_31699_20742.n24 1.44113
R47035 a_31699_20742.n8 a_31699_20742.n9 1.44113
R47036 a_31699_20742.n39 a_31699_20742.n7 1.44113
R47037 a_31699_20742.n32 a_31699_20742.n33 1.44113
R47038 a_31699_20742.n22 a_31699_20742.n23 1.44113
R47039 a_31699_20742.n212 a_31699_20742.n213 0.332154
R47040 a_31699_20742.n59 a_31699_20742.n60 1.44113
R47041 a_31699_20742.n57 a_31699_20742.n58 1.44113
R47042 a_31699_20742.n264 a_31699_20742.n263 4.5005
R47043 a_31699_20742.n52 a_31699_20742.n51 1.44113
R47044 a_31699_20742.n53 a_31699_20742.n54 1.44113
R47045 a_31699_20742.n56 a_31699_20742.n55 1.44113
R47046 a_31699_20742.n49 a_31699_20742.n50 1.44113
R47047 a_31699_20742.n48 a_31699_20742.n47 1.44113
R47048 a_31699_20742.n46 a_31699_20742.n45 1.44113
R47049 a_31699_20742.n304 a_31699_20742.n303 4.5005
R47050 a_31699_20742.n42 a_31699_20742.n41 1.44113
R47051 a_31699_20742.n44 a_31699_20742.n43 1.44113
R47052 a_31699_20742.n192 a_31699_20742.n193 0.349872
R47053 a_31699_20742.n369 a_31699_20742.n368 4.5005
R47054 a_31699_20742.n82 a_31699_20742.n81 1.44113
R47055 a_31699_20742.n385 a_31699_20742.n384 4.5005
R47056 a_31699_20742.n383 a_31699_20742.n374 4.5005
R47057 a_31699_20742.n382 a_31699_20742.n381 4.5005
R47058 a_31699_20742.n380 a_31699_20742.n375 4.5005
R47059 a_31699_20742.n379 a_31699_20742.n378 4.5005
R47060 a_31699_20742.n309 a_31699_20742.n252 3.97759
R47061 a_31699_20742.n244 a_31699_20742.n243 3.87147
R47062 a_31699_20742.n240 a_31699_20742.t4 3.86699
R47063 a_31699_20742.n240 a_31699_20742.t30 3.66212
R47064 a_31699_20742.n251 a_31699_20742.n239 3.08458
R47065 a_31699_20742.n239 a_31699_20742.n250 2.73715
R47066 a_31699_20742.n246 a_31699_20742.n245 2.51878
R47067 a_31699_20742.n251 a_31699_20742.n217 2.44398
R47068 a_31699_20742.n218 a_31699_20742.n247 3.87147
R47069 a_31699_20742.n250 a_31699_20742.n248 2.39895
R47070 a_31699_20742.n288 a_31699_20742.n265 2.30989
R47071 a_31699_20742.n280 a_31699_20742.n197 2.30989
R47072 a_31699_20742.n302 a_31699_20742.n260 2.25752
R47073 a_31699_20742.n287 a_31699_20742.n286 2.25752
R47074 a_31699_20742.n386 a_31699_20742.n373 2.25278
R47075 a_31699_20742.n218 a_31699_20742.n217 0.0670397
R47076 a_31699_20742.n220 a_31699_20742.n219 1.44642
R47077 a_31699_20742.n221 a_31699_20742.n175 1.44642
R47078 a_31699_20742.n222 a_31699_20742.n178 1.44642
R47079 a_31699_20742.n223 a_31699_20742.n181 1.44642
R47080 a_31699_20742.n227 a_31699_20742.n226 1.44612
R47081 a_31699_20742.n228 a_31699_20742.n200 1.44612
R47082 a_31699_20742.n229 a_31699_20742.n203 1.44612
R47083 a_31699_20742.n231 a_31699_20742.n230 1.44612
R47084 a_31699_20742.n250 a_31699_20742.n249 2.19216
R47085 a_31699_20742.n117 a_31699_20742.n255 2.49908
R47086 a_31699_20742.n224 a_31699_20742.n123 2.49908
R47087 a_31699_20742.n225 a_31699_20742.n126 2.49908
R47088 a_31699_20742.n133 a_31699_20742.n311 2.49908
R47089 a_31699_20742.n254 a_31699_20742.n237 2.07182
R47090 a_31699_20742.n256 a_31699_20742.n236 2.07182
R47091 a_31699_20742.n237 a_31699_20742.n157 2.4644
R47092 a_31699_20742.n161 a_31699_20742.n236 2.4644
R47093 a_31699_20742.n150 a_31699_20742.n257 2.4644
R47094 a_31699_20742.n238 a_31699_20742.n155 2.4644
R47095 a_31699_20742.n309 a_31699_20742.n308 2.01366
R47096 a_31699_20742.n334 a_31699_20742.n323 1.61908
R47097 a_31699_20742.n313 a_31699_20742.n312 1.53101
R47098 a_31699_20742.n310 a_31699_20742.n309 1.53101
R47099 a_31699_20742.n257 a_31699_20742.n253 1.5005
R47100 a_31699_20742.n255 a_31699_20742.n254 1.5005
R47101 a_31699_20742.n312 a_31699_20742.n225 1.5005
R47102 a_31699_20742.n311 a_31699_20742.n310 1.5005
R47103 a_31699_20742.n258 a_31699_20742.n238 1.5005
R47104 a_31699_20742.n256 a_31699_20742.n224 1.5005
R47105 a_31699_20742.n296 a_31699_20742.n196 1.5005
R47106 a_31699_20742.n288 a_31699_20742.n194 1.5005
R47107 a_31699_20742.n298 a_31699_20742.n297 1.5005
R47108 a_31699_20742.n308 a_31699_20742.n195 1.5005
R47109 a_31699_20742.n292 a_31699_20742.n259 1.5005
R47110 a_31699_20742.n281 a_31699_20742.n280 1.5005
R47111 a_31699_20742.n209 a_31699_20742.n365 1.5005
R47112 a_31699_20742.n208 a_31699_20742.n355 1.5005
R47113 a_31699_20742.n209 a_31699_20742.n387 1.5005
R47114 a_31699_20742.n345 a_31699_20742.n344 1.5005
R47115 a_31699_20742.n334 a_31699_20742.n333 1.5005
R47116 a_31699_20742.n234 a_31699_20742.n390 1.5005
R47117 a_31699_20742.n254 a_31699_20742.n253 1.47516
R47118 a_31699_20742.n258 a_31699_20742.n256 1.47516
R47119 a_31699_20742.n247 a_31699_20742.t16 1.4705
R47120 a_31699_20742.n247 a_31699_20742.t42 1.4705
R47121 a_31699_20742.n243 a_31699_20742.t34 1.4705
R47122 a_31699_20742.n243 a_31699_20742.t8 1.4705
R47123 a_31699_20742.n248 a_31699_20742.t24 1.4705
R47124 a_31699_20742.n248 a_31699_20742.t14 1.4705
R47125 a_31699_20742.n249 a_31699_20742.t18 1.4705
R47126 a_31699_20742.n249 a_31699_20742.t40 1.4705
R47127 a_31699_20742.n242 a_31699_20742.t22 1.4705
R47128 a_31699_20742.n242 a_31699_20742.t10 1.4705
R47129 a_31699_20742.t44 a_31699_20742.n391 1.4705
R47130 a_31699_20742.n391 a_31699_20742.t20 1.4705
R47131 a_31699_20742.n388 a_31699_20742.n209 1.42915
R47132 a_31699_20742.n297 a_31699_20742.n252 1.41182
R47133 a_31699_20742.n140 a_31699_20742.t160 8.49836
R47134 a_31699_20742.n139 a_31699_20742.t67 8.49836
R47135 a_31699_20742.n245 a_31699_20742.n244 1.27228
R47136 a_31699_20742.n28 a_31699_20742.n279 1.24866
R47137 a_31699_20742.n30 a_31699_20742.n276 1.24866
R47138 a_31699_20742.n293 a_31699_20742.n32 1.24866
R47139 a_31699_20742.n34 a_31699_20742.n291 1.24866
R47140 a_31699_20742.n277 a_31699_20742.n0 1.24629
R47141 a_31699_20742.n274 a_31699_20742.n37 1.24629
R47142 a_31699_20742.n7 a_31699_20742.n295 1.24629
R47143 a_31699_20742.n289 a_31699_20742.n13 1.24629
R47144 a_31699_20742.n296 a_31699_20742.n288 1.23709
R47145 a_31699_20742.n280 a_31699_20742.n259 1.23709
R47146 a_31699_20742.n305 a_31699_20742.n49 1.22261
R47147 a_31699_20742.n299 a_31699_20742.n59 1.22261
R47148 a_31699_20742.n69 a_31699_20742.n284 1.22261
R47149 a_31699_20742.n270 a_31699_20742.n79 1.22261
R47150 a_31699_20742.n41 a_31699_20742.n307 1.21313
R47151 a_31699_20742.n52 a_31699_20742.n301 1.21313
R47152 a_31699_20742.n282 a_31699_20742.n61 1.21313
R47153 a_31699_20742.n71 a_31699_20742.n272 1.21313
R47154 a_31699_20742.n217 a_31699_20742.n246 1.20609
R47155 a_31699_20742.n390 a_31699_20742.n389 1.17709
R47156 a_31699_20742.n269 a_31699_20742.n268 1.12904
R47157 a_31699_20742.n263 a_31699_20742.n262 1.12904
R47158 a_31699_20742.n368 a_31699_20742.n367 1.129
R47159 a_31699_20742.n379 a_31699_20742.n376 1.12765
R47160 a_31699_20742.n317 a_31699_20742.n316 0.915282
R47161 a_31699_20742.n327 a_31699_20742.n326 0.915282
R47162 a_31699_20742.n338 a_31699_20742.n337 0.915282
R47163 a_31699_20742.n349 a_31699_20742.n348 0.915282
R47164 a_31699_20742.n359 a_31699_20742.n358 0.915282
R47165 a_31699_20742.n390 a_31699_20742.n251 0.886209
R47166 a_31699_20742.n297 a_31699_20742.n296 0.809892
R47167 a_31699_20742.n308 a_31699_20742.n259 0.809892
R47168 a_31699_20742.n31 a_31699_20742.n265 0.888471
R47169 a_31699_20742.n197 a_31699_20742.n29 0.888471
R47170 a_31699_20742.n196 a_31699_20742.n35 0.888471
R47171 a_31699_20742.n33 a_31699_20742.n292 0.888471
R47172 a_31699_20742.n389 a_31699_20742.n388 0.741617
R47173 a_31699_20742.n194 a_31699_20742.n72 0.854361
R47174 a_31699_20742.n62 a_31699_20742.n281 0.854361
R47175 a_31699_20742.n298 a_31699_20742.n51 0.854361
R47176 a_31699_20742.n195 a_31699_20742.n42 0.854361
R47177 a_31699_20742.n323 a_31699_20742.n322 0.688348
R47178 a_31699_20742.n333 a_31699_20742.n332 0.688348
R47179 a_31699_20742.n344 a_31699_20742.n343 0.688348
R47180 a_31699_20742.n355 a_31699_20742.n354 0.688348
R47181 a_31699_20742.n365 a_31699_20742.n364 0.688348
R47182 a_31699_20742.n306 a_31699_20742.n305 0.673132
R47183 a_31699_20742.n307 a_31699_20742.n306 0.673132
R47184 a_31699_20742.n300 a_31699_20742.n299 0.673132
R47185 a_31699_20742.n301 a_31699_20742.n300 0.673132
R47186 a_31699_20742.n278 a_31699_20742.n277 0.673132
R47187 a_31699_20742.n279 a_31699_20742.n278 0.673132
R47188 a_31699_20742.n275 a_31699_20742.n274 0.673132
R47189 a_31699_20742.n276 a_31699_20742.n275 0.673132
R47190 a_31699_20742.n284 a_31699_20742.n283 0.673132
R47191 a_31699_20742.n283 a_31699_20742.n282 0.673132
R47192 a_31699_20742.n271 a_31699_20742.n270 0.673132
R47193 a_31699_20742.n272 a_31699_20742.n271 0.673132
R47194 a_31699_20742.n295 a_31699_20742.n294 0.673132
R47195 a_31699_20742.n294 a_31699_20742.n293 0.673132
R47196 a_31699_20742.n290 a_31699_20742.n289 0.673132
R47197 a_31699_20742.n291 a_31699_20742.n290 0.673132
R47198 a_31699_20742.n318 a_31699_20742.n317 0.655148
R47199 a_31699_20742.n328 a_31699_20742.n327 0.655148
R47200 a_31699_20742.n339 a_31699_20742.n338 0.655148
R47201 a_31699_20742.n371 a_31699_20742.n370 0.655148
R47202 a_31699_20742.n350 a_31699_20742.n349 0.655148
R47203 a_31699_20742.n360 a_31699_20742.n359 0.655148
R47204 a_31699_20742.n316 a_31699_20742.n315 0.63334
R47205 a_31699_20742.n322 a_31699_20742.n321 0.63334
R47206 a_31699_20742.n321 a_31699_20742.n320 0.63334
R47207 a_31699_20742.n326 a_31699_20742.n325 0.63334
R47208 a_31699_20742.n332 a_31699_20742.n331 0.63334
R47209 a_31699_20742.n331 a_31699_20742.n330 0.63334
R47210 a_31699_20742.n337 a_31699_20742.n336 0.63334
R47211 a_31699_20742.n343 a_31699_20742.n342 0.63334
R47212 a_31699_20742.n342 a_31699_20742.n341 0.63334
R47213 a_31699_20742.n348 a_31699_20742.n347 0.63334
R47214 a_31699_20742.n354 a_31699_20742.n353 0.63334
R47215 a_31699_20742.n353 a_31699_20742.n352 0.63334
R47216 a_31699_20742.n358 a_31699_20742.n357 0.63334
R47217 a_31699_20742.n364 a_31699_20742.n363 0.63334
R47218 a_31699_20742.n363 a_31699_20742.n362 0.63334
R47219 a_31699_20742.n315 a_31699_20742.n314 0.63225
R47220 a_31699_20742.n319 a_31699_20742.n318 0.63225
R47221 a_31699_20742.n325 a_31699_20742.n324 0.63225
R47222 a_31699_20742.n329 a_31699_20742.n328 0.63225
R47223 a_31699_20742.n336 a_31699_20742.n335 0.63225
R47224 a_31699_20742.n340 a_31699_20742.n339 0.63225
R47225 a_31699_20742.n372 a_31699_20742.n371 0.63225
R47226 a_31699_20742.n347 a_31699_20742.n346 0.63225
R47227 a_31699_20742.n351 a_31699_20742.n350 0.63225
R47228 a_31699_20742.n357 a_31699_20742.n356 0.63225
R47229 a_31699_20742.n361 a_31699_20742.n360 0.63225
R47230 a_31699_20742.n387 a_31699_20742.n386 0.622055
R47231 a_31699_20742.n313 a_31699_20742.n252 0.602344
R47232 a_31699_20742.n312 a_31699_20742.n253 0.571818
R47233 a_31699_20742.n310 a_31699_20742.n258 0.571818
R47234 a_31699_20742.n208 a_31699_20742.n345 0.467527
R47235 a_31699_20742.n63 a_31699_20742.n189 0.379447
R47236 a_31699_20742.n384 a_31699_20742.n383 0.379447
R47237 a_31699_20742.n378 a_31699_20742.n375 0.379447
R47238 a_31699_20742.n112 a_31699_20742.n125 1.14293
R47239 a_31699_20742.n115 a_31699_20742.n128 1.14293
R47240 a_31699_20742.n172 a_31699_20742.n132 1.74606
R47241 a_31699_20742.n105 a_31699_20742.n116 1.14293
R47242 a_31699_20742.n109 a_31699_20742.n118 1.14293
R47243 a_31699_20742.n171 a_31699_20742.n122 1.74606
R47244 a_31699_20742.n104 a_31699_20742.n117 1.14293
R47245 a_31699_20742.n108 a_31699_20742.n119 1.14293
R47246 a_31699_20742.n171 a_31699_20742.n123 1.74702
R47247 a_31699_20742.n111 a_31699_20742.n126 1.14293
R47248 a_31699_20742.n129 a_31699_20742.n114 1.14293
R47249 a_31699_20742.n172 a_31699_20742.n133 1.74702
R47250 a_31699_20742.n21 a_31699_20742.n4 0.647707
R47251 a_31699_20742.n2 a_31699_20742.n19 0.647707
R47252 a_31699_20742.n211 a_31699_20742.n17 1.34142
R47253 a_31699_20742.n12 a_31699_20742.n27 0.647707
R47254 a_31699_20742.n9 a_31699_20742.n25 0.647707
R47255 a_31699_20742.n213 a_31699_20742.n23 1.34142
R47256 a_31699_20742.n21 a_31699_20742.n31 0.635332
R47257 a_31699_20742.n145 a_31699_20742.n19 0.634233
R47258 a_31699_20742.n29 a_31699_20742.n17 0.635332
R47259 a_31699_20742.n35 a_31699_20742.n27 0.635332
R47260 a_31699_20742.n143 a_31699_20742.n25 0.634233
R47261 a_31699_20742.n23 a_31699_20742.n33 0.635332
R47262 a_31699_20742.n221 a_31699_20742.n177 0.891677
R47263 a_31699_20742.n174 a_31699_20742.n220 0.891677
R47264 a_31699_20742.n228 a_31699_20742.n202 0.891728
R47265 a_31699_20742.n199 a_31699_20742.n227 0.891728
R47266 a_31699_20742.n157 a_31699_20742.n88 1.1526
R47267 a_31699_20742.n84 a_31699_20742.n164 1.15248
R47268 a_31699_20742.n161 a_31699_20742.n216 1.74338
R47269 a_31699_20742.n223 a_31699_20742.n183 0.891677
R47270 a_31699_20742.n222 a_31699_20742.n180 0.891677
R47271 a_31699_20742.n207 a_31699_20742.n231 0.891728
R47272 a_31699_20742.n229 a_31699_20742.n205 0.891728
R47273 a_31699_20742.n98 a_31699_20742.n150 1.15284
R47274 a_31699_20742.n94 a_31699_20742.n152 1.1526
R47275 a_31699_20742.n155 a_31699_20742.n215 1.74338
R47276 a_31699_20742.n78 a_31699_20742.n269 0.496611
R47277 a_31699_20742.n66 a_31699_20742.n273 0.496611
R47278 a_31699_20742.n263 a_31699_20742.n58 0.496611
R47279 a_31699_20742.n303 a_31699_20742.n46 0.496611
R47280 a_31699_20742.n385 a_31699_20742.n374 0.3605
R47281 a_31699_20742.n380 a_31699_20742.n379 0.3605
R47282 a_31699_20742.n368 a_31699_20742.n82 0.495486
R47283 a_31699_20742.n262 a_31699_20742.n261 0.327481
R47284 a_31699_20742.n268 a_31699_20742.n267 0.327481
R47285 a_31699_20742.n367 a_31699_20742.n366 0.32675
R47286 a_31699_20742.n377 a_31699_20742.n376 0.324133
R47287 a_31699_20742.n345 a_31699_20742.n334 0.301209
R47288 a_31699_20742.n148 a_31699_20742.n4 0.558475
R47289 a_31699_20742.n36 a_31699_20742.n2 0.559597
R47290 a_31699_20742.n146 a_31699_20742.n12 0.558475
R47291 a_31699_20742.n39 a_31699_20742.n9 0.559597
R47292 a_31699_20742.n323 a_31699_20742.n319 0.254694
R47293 a_31699_20742.n333 a_31699_20742.n329 0.254694
R47294 a_31699_20742.n344 a_31699_20742.n340 0.254694
R47295 a_31699_20742.n387 a_31699_20742.n372 0.254694
R47296 a_31699_20742.n355 a_31699_20742.n351 0.254694
R47297 a_31699_20742.n365 a_31699_20742.n361 0.254694
R47298 a_31699_20742.n287 a_31699_20742.n273 0.208099
R47299 a_31699_20742.n303 a_31699_20742.n302 0.208099
R47300 a_31699_20742.n386 a_31699_20742.n385 0.208099
R47301 a_31699_20742.n384 a_31699_20742.n373 0.147342
R47302 a_31699_20742.n383 a_31699_20742.n382 0.147342
R47303 a_31699_20742.n382 a_31699_20742.n375 0.147342
R47304 a_31699_20742.n378 a_31699_20742.n377 0.147342
R47305 a_31699_20742.n369 a_31699_20742.n366 0.143789
R47306 a_31699_20742.n304 a_31699_20742.n260 0.142605
R47307 a_31699_20742.n264 a_31699_20742.n261 0.142605
R47308 a_31699_20742.n286 a_31699_20742.n285 0.142605
R47309 a_31699_20742.n267 a_31699_20742.n266 0.142605
R47310 a_31699_20742.n137 a_31699_20742.n169 1.73389
R47311 a_31699_20742.n221 a_31699_20742.n169 1.19478
R47312 a_31699_20742.n125 a_31699_20742.n177 1.49218
R47313 a_31699_20742.n128 a_31699_20742.n112 3.79267
R47314 a_31699_20742.n220 a_31699_20742.n115 1.19478
R47315 a_31699_20742.n174 a_31699_20742.n132 1.49218
R47316 a_31699_20742.n228 a_31699_20742.n91 1.6448
R47317 a_31699_20742.n156 a_31699_20742.n202 1.49177
R47318 a_31699_20742.n156 a_31699_20742.n89 1.14306
R47319 a_31699_20742.n89 a_31699_20742.n163 3.79279
R47320 a_31699_20742.n85 a_31699_20742.n163 1.14293
R47321 a_31699_20742.n227 a_31699_20742.n85 1.19475
R47322 a_31699_20742.n199 a_31699_20742.n160 1.49177
R47323 a_31699_20742.n216 a_31699_20742.n160 1.74677
R47324 a_31699_20742.n91 a_31699_20742.n237 1.65371
R47325 a_31699_20742.n164 a_31699_20742.n88 3.7612
R47326 a_31699_20742.n84 a_31699_20742.n236 1.21357
R47327 a_31699_20742.n166 a_31699_20742.n135 1.73389
R47328 a_31699_20742.n223 a_31699_20742.n166 1.19478
R47329 a_31699_20742.n116 a_31699_20742.n183 1.49218
R47330 a_31699_20742.n118 a_31699_20742.n105 3.79267
R47331 a_31699_20742.n222 a_31699_20742.n109 1.19478
R47332 a_31699_20742.n122 a_31699_20742.n180 1.49218
R47333 a_31699_20742.n135 a_31699_20742.n167 1.7332
R47334 a_31699_20742.n255 a_31699_20742.n167 1.21084
R47335 a_31699_20742.n104 a_31699_20742.n119 3.79267
R47336 a_31699_20742.n108 a_31699_20742.n224 1.21084
R47337 a_31699_20742.n231 a_31699_20742.n101 1.64472
R47338 a_31699_20742.n207 a_31699_20742.n149 1.49177
R47339 a_31699_20742.n99 a_31699_20742.n149 1.14329
R47340 a_31699_20742.n151 a_31699_20742.n99 3.79231
R47341 a_31699_20742.n95 a_31699_20742.n151 1.14306
R47342 a_31699_20742.n229 a_31699_20742.n95 1.19488
R47343 a_31699_20742.n154 a_31699_20742.n205 1.49177
R47344 a_31699_20742.n154 a_31699_20742.n215 1.74677
R47345 a_31699_20742.n257 a_31699_20742.n101 1.65364
R47346 a_31699_20742.n152 a_31699_20742.n98 3.76072
R47347 a_31699_20742.n94 a_31699_20742.n238 1.21369
R47348 a_31699_20742.n170 a_31699_20742.n137 1.7332
R47349 a_31699_20742.n170 a_31699_20742.n225 1.21084
R47350 a_31699_20742.n111 a_31699_20742.n129 3.79267
R47351 a_31699_20742.n114 a_31699_20742.n311 1.21084
R47352 a_31699_20742.n140 a_31699_20742.n6 1.34213
R47353 a_31699_20742.n38 a_31699_20742.n6 0.559597
R47354 a_31699_20742.n265 a_31699_20742.n38 2.32622
R47355 a_31699_20742.n145 a_31699_20742.n148 3.29987
R47356 a_31699_20742.n36 a_31699_20742.n197 2.32622
R47357 a_31699_20742.n80 a_31699_20742.n78 0.633082
R47358 a_31699_20742.n80 a_31699_20742.n194 2.30372
R47359 a_31699_20742.n74 a_31699_20742.n72 0.633082
R47360 a_31699_20742.n74 a_31699_20742.n76 0.633082
R47361 a_31699_20742.n76 a_31699_20742.n187 0.631741
R47362 a_31699_20742.n187 a_31699_20742.n287 3.17649
R47363 a_31699_20742.n66 a_31699_20742.n68 0.633082
R47364 a_31699_20742.n68 a_31699_20742.n70 0.633082
R47365 a_31699_20742.n70 a_31699_20742.n281 2.30372
R47366 a_31699_20742.n62 a_31699_20742.n64 0.633082
R47367 a_31699_20742.n64 a_31699_20742.n188 1.32892
R47368 a_31699_20742.n15 a_31699_20742.n139 1.34213
R47369 a_31699_20742.n40 a_31699_20742.n15 0.559597
R47370 a_31699_20742.n40 a_31699_20742.n196 2.32622
R47371 a_31699_20742.n146 a_31699_20742.n143 3.29987
R47372 a_31699_20742.n39 a_31699_20742.n292 2.32622
R47373 a_31699_20742.n60 a_31699_20742.n58 0.633082
R47374 a_31699_20742.n298 a_31699_20742.n60 2.30372
R47375 a_31699_20742.n54 a_31699_20742.n51 0.633082
R47376 a_31699_20742.n56 a_31699_20742.n54 0.633082
R47377 a_31699_20742.n191 a_31699_20742.n56 0.631741
R47378 a_31699_20742.n302 a_31699_20742.n191 3.17649
R47379 a_31699_20742.n48 a_31699_20742.n46 0.633082
R47380 a_31699_20742.n50 a_31699_20742.n48 0.633082
R47381 a_31699_20742.n50 a_31699_20742.n195 2.30372
R47382 a_31699_20742.n44 a_31699_20742.n42 0.633082
R47383 a_31699_20742.n44 a_31699_20742.n193 1.32892
R47384 a_31699_20742.n185 a_31699_20742.n82 0.631741
R47385 a_31699_20742.n370 a_31699_20742.n185 0.917116
R47386 a_31699_20742.n381 a_31699_20742.n374 0.14
R47387 a_31699_20742.n381 a_31699_20742.n380 0.14
R47388 a_31699_20742.n241 a_31699_20742.n232 1.27192
R47389 a_31699_20742.n233 a_31699_20742.n232 2.51878
R47390 a_31699_20742.n234 a_31699_20742.n233 1.2061
R47391 a_31699_20742.t36 a_31699_20742.n235 6.57099
R47392 a_31699_20742.n218 a_31699_20742.t28 6.61288
R47393 a_31699_20742.n71 a_31699_20742.n73 0.966816
R47394 a_31699_20742.n61 a_31699_20742.n63 0.966816
R47395 a_31699_20742.n53 a_31699_20742.n52 0.966816
R47396 a_31699_20742.n8 a_31699_20742.n7 0.889842
R47397 a_31699_20742.n1 a_31699_20742.n0 0.889842
R47398 a_31699_20742.n11 a_31699_20742.n10 0.771421
R47399 a_31699_20742.n147 a_31699_20742.n3 0.771421
R47400 a_31699_20742.n26 a_31699_20742.n11 0.688526
R47401 a_31699_20742.n24 a_31699_20742.n8 0.688526
R47402 a_31699_20742.n22 a_31699_20742.n212 0.688526
R47403 a_31699_20742.n3 a_31699_20742.n20 0.688526
R47404 a_31699_20742.n1 a_31699_20742.n18 0.688526
R47405 a_31699_20742.n16 a_31699_20742.n210 0.688526
R47406 a_31699_20742.n14 a_31699_20742.n138 0.688526
R47407 a_31699_20742.n5 a_31699_20742.n141 0.688526
R47408 a_31699_20742.n34 a_31699_20742.n26 0.6755
R47409 a_31699_20742.n32 a_31699_20742.n22 0.6755
R47410 a_31699_20742.n20 a_31699_20742.n30 0.6755
R47411 a_31699_20742.n28 a_31699_20742.n16 0.6755
R47412 a_31699_20742.n77 a_31699_20742.n79 0.673132
R47413 a_31699_20742.n77 a_31699_20742.n266 0.673132
R47414 a_31699_20742.n73 a_31699_20742.n75 0.673132
R47415 a_31699_20742.n67 a_31699_20742.n69 0.673132
R47416 a_31699_20742.n65 a_31699_20742.n67 0.673132
R47417 a_31699_20742.n285 a_31699_20742.n65 0.673132
R47418 a_31699_20742.n59 a_31699_20742.n57 0.673132
R47419 a_31699_20742.n57 a_31699_20742.n264 0.673132
R47420 a_31699_20742.n55 a_31699_20742.n53 0.673132
R47421 a_31699_20742.n47 a_31699_20742.n49 0.673132
R47422 a_31699_20742.n47 a_31699_20742.n45 0.673132
R47423 a_31699_20742.n45 a_31699_20742.n304 0.673132
R47424 a_31699_20742.n43 a_31699_20742.n192 0.673132
R47425 a_31699_20742.n41 a_31699_20742.n43 0.673132
R47426 a_31699_20742.n81 a_31699_20742.n369 0.671947
R47427 a_31699_20742.n127 a_31699_20742.n113 0.609682
R47428 a_31699_20742.n124 a_31699_20742.n110 0.609682
R47429 a_31699_20742.n107 a_31699_20742.n106 0.609682
R47430 a_31699_20742.n103 a_31699_20742.n102 0.609682
R47431 a_31699_20742.n97 a_31699_20742.n96 0.609682
R47432 a_31699_20742.n93 a_31699_20742.n92 0.609682
R47433 a_31699_20742.n87 a_31699_20742.n86 0.609682
R47434 a_31699_20742.n162 a_31699_20742.n83 0.609682
R47435 a_31699_20742.n14 a_31699_20742.n13 0.596158
R47436 a_31699_20742.n37 a_31699_20742.n5 0.596158
R47437 a_31699_20742.n18 a_31699_20742.n144 0.559447
R47438 a_31699_20742.n142 a_31699_20742.n24 0.559447
R47439 a_31699_20742.n190 a_31699_20742.n55 0.531026
R47440 a_31699_20742.n75 a_31699_20742.n186 0.531026
R47441 a_31699_20742.n184 a_31699_20742.n81 0.531026
R47442 a_31699_20742.n209 a_31699_20742.n208 0.427696
R47443 a_31699_20742.n182 a_31699_20742.n181 0.386311
R47444 a_31699_20742.n179 a_31699_20742.n178 0.386311
R47445 a_31699_20742.n176 a_31699_20742.n175 0.386311
R47446 a_31699_20742.n219 a_31699_20742.n173 0.386311
R47447 a_31699_20742.n131 a_31699_20742.n130 0.369148
R47448 a_31699_20742.n121 a_31699_20742.n120 0.369148
R47449 a_31699_20742.n230 a_31699_20742.n206 0.364343
R47450 a_31699_20742.n204 a_31699_20742.n203 0.364343
R47451 a_31699_20742.n201 a_31699_20742.n200 0.364343
R47452 a_31699_20742.n226 a_31699_20742.n198 0.364343
R47453 a_31699_20742.n159 a_31699_20742.n158 0.354735
R47454 a_31699_20742.n214 a_31699_20742.n153 0.354735
R47455 a_31699_20742.n168 a_31699_20742.n136 0.347689
R47456 a_31699_20742.n165 a_31699_20742.n134 0.347689
R47457 a_35502_24538.n131 a_35502_24538.n130 12.734
R47458 a_35502_24538.n57 a_35502_24538.t36 8.41809
R47459 a_35502_24538.n58 a_35502_24538.t59 8.41809
R47460 a_35502_24538.n57 a_35502_24538.t34 8.37125
R47461 a_35502_24538.n61 a_35502_24538.t41 8.37125
R47462 a_35502_24538.n58 a_35502_24538.t56 8.37125
R47463 a_35502_24538.n104 a_35502_24538.t25 8.33806
R47464 a_35502_24538.n98 a_35502_24538.t61 8.3366
R47465 a_35502_24538.n83 a_35502_24538.t47 8.26493
R47466 a_35502_24538.n117 a_35502_24538.t39 8.2602
R47467 a_35502_24538.n17 a_35502_24538.t42 8.06917
R47468 a_35502_24538.n28 a_35502_24538.t38 8.06917
R47469 a_35502_24538.n13 a_35502_24538.t50 8.06917
R47470 a_35502_24538.n13 a_35502_24538.t48 8.06917
R47471 a_35502_24538.n11 a_35502_24538.t40 8.06917
R47472 a_35502_24538.n11 a_35502_24538.t55 8.06917
R47473 a_35502_24538.n63 a_35502_24538.t26 8.06917
R47474 a_35502_24538.n17 a_35502_24538.t53 8.06917
R47475 a_35502_24538.n30 a_35502_24538.t24 8.06917
R47476 a_35502_24538.n7 a_35502_24538.t64 8.06917
R47477 a_35502_24538.n7 a_35502_24538.t37 8.06917
R47478 a_35502_24538.n32 a_35502_24538.t49 8.06917
R47479 a_35502_24538.n77 a_35502_24538.t62 8.06917
R47480 a_35502_24538.n3 a_35502_24538.t33 8.06917
R47481 a_35502_24538.n3 a_35502_24538.t31 8.06917
R47482 a_35502_24538.n21 a_35502_24538.t60 8.06917
R47483 a_35502_24538.n21 a_35502_24538.t32 8.06917
R47484 a_35502_24538.n71 a_35502_24538.t46 8.06917
R47485 a_35502_24538.n97 a_35502_24538.t29 8.06917
R47486 a_35502_24538.n0 a_35502_24538.t28 8.06917
R47487 a_35502_24538.n95 a_35502_24538.t57 8.06917
R47488 a_35502_24538.n94 a_35502_24538.t30 8.06917
R47489 a_35502_24538.n93 a_35502_24538.t45 8.06917
R47490 a_35502_24538.n91 a_35502_24538.t63 8.06917
R47491 a_35502_24538.n84 a_35502_24538.t35 8.06917
R47492 a_35502_24538.n111 a_35502_24538.t43 8.06917
R47493 a_35502_24538.n105 a_35502_24538.t54 8.06917
R47494 a_35502_24538.n113 a_35502_24538.t27 8.06917
R47495 a_35502_24538.n114 a_35502_24538.t58 8.06917
R47496 a_35502_24538.n115 a_35502_24538.t44 8.06917
R47497 a_35502_24538.n118 a_35502_24538.t52 8.06917
R47498 a_35502_24538.n124 a_35502_24538.t51 8.06917
R47499 a_35502_24538.n60 a_35502_24538.t0 6.65728
R47500 a_35502_24538.n46 a_35502_24538.t7 6.51495
R47501 a_35502_24538.n134 a_35502_24538.t15 6.40828
R47502 a_35502_24538.n43 a_35502_24538.t17 6.37877
R47503 a_35502_24538.n60 a_35502_24538.t1 5.74368
R47504 a_35502_24538.n47 a_35502_24538.t6 5.24318
R47505 a_35502_24538.n65 a_35502_24538.n31 2.4223
R47506 a_35502_24538.n72 a_35502_24538.n33 2.42484
R47507 a_35502_24538.n73 a_35502_24538.n33 2.4256
R47508 a_35502_24538.n39 a_35502_24538.n38 2.24636
R47509 a_35502_24538.t11 a_35502_24538.n35 5.26436
R47510 a_35502_24538.n54 a_35502_24538.n43 4.60825
R47511 a_35502_24538.n34 a_35502_24538.n138 3.79435
R47512 a_35502_24538.n38 a_35502_24538.n134 4.59811
R47513 a_35502_24538.n22 a_35502_24538.n21 0.592766
R47514 a_35502_24538.n12 a_35502_24538.n11 0.592803
R47515 a_35502_24538.n15 a_35502_24538.n13 0.591918
R47516 a_35502_24538.n17 a_35502_24538.n18 0.591826
R47517 a_35502_24538.n37 a_35502_24538.n36 2.24389
R47518 a_35502_24538.n50 a_35502_24538.n44 4.5005
R47519 a_35502_24538.n10 a_35502_24538.n67 4.5005
R47520 a_35502_24538.n13 a_35502_24538.n14 0.591264
R47521 a_35502_24538.n68 a_35502_24538.n24 4.5005
R47522 a_35502_24538.n31 a_35502_24538.n30 0.0133501
R47523 a_35502_24538.n16 a_35502_24538.n65 4.5005
R47524 a_35502_24538.n19 a_35502_24538.n17 0.604195
R47525 a_35502_24538.n29 a_35502_24538.n64 4.5005
R47526 a_35502_24538.n70 a_35502_24538.n69 4.5005
R47527 a_35502_24538.n28 a_35502_24538.n27 0.0143905
R47528 a_35502_24538.n20 a_35502_24538.n75 4.5005
R47529 a_35502_24538.n2 a_35502_24538.n76 4.5005
R47530 a_35502_24538.n3 a_35502_24538.n4 0.591675
R47531 a_35502_24538.n9 a_35502_24538.n7 0.604671
R47532 a_35502_24538.n6 a_35502_24538.n72 4.5005
R47533 a_35502_24538.n32 a_35502_24538.n33 0.0107891
R47534 a_35502_24538.n7 a_35502_24538.n8 0.604671
R47535 a_35502_24538.n73 a_35502_24538.n6 4.5005
R47536 a_35502_24538.n2 a_35502_24538.n23 4.5005
R47537 a_35502_24538.n5 a_35502_24538.n3 0.591675
R47538 a_35502_24538.n85 a_35502_24538.n82 4.5005
R47539 a_35502_24538.n87 a_35502_24538.n86 4.5005
R47540 a_35502_24538.n88 a_35502_24538.n81 4.5005
R47541 a_35502_24538.n90 a_35502_24538.n89 4.5005
R47542 a_35502_24538.n92 a_35502_24538.n80 4.5005
R47543 a_35502_24538.n1 a_35502_24538.n0 1.44113
R47544 a_35502_24538.n99 a_35502_24538.n96 4.5005
R47545 a_35502_24538.n112 a_35502_24538.n101 4.5005
R47546 a_35502_24538.n110 a_35502_24538.n109 4.5005
R47547 a_35502_24538.n108 a_35502_24538.n103 4.5005
R47548 a_35502_24538.n107 a_35502_24538.n106 4.5005
R47549 a_35502_24538.n127 a_35502_24538.n126 4.5005
R47550 a_35502_24538.n125 a_35502_24538.n102 4.5005
R47551 a_35502_24538.n123 a_35502_24538.n122 4.5005
R47552 a_35502_24538.n121 a_35502_24538.n116 4.5005
R47553 a_35502_24538.n120 a_35502_24538.n119 4.5005
R47554 a_35502_24538.n42 a_35502_24538.n41 2.23676
R47555 a_35502_24538.n139 a_35502_24538.n40 4.5005
R47556 a_35502_24538.n36 a_35502_24538.t9 3.79594
R47557 a_35502_24538.n41 a_35502_24538.t3 3.79475
R47558 a_35502_24538.t23 a_35502_24538.n141 3.77936
R47559 a_35502_24538.n51 a_35502_24538.t12 3.77818
R47560 a_35502_24538.n46 a_35502_24538.n45 3.77318
R47561 a_35502_24538.n137 a_35502_24538.n136 3.77081
R47562 a_35502_24538.n49 a_35502_24538.n48 3.75571
R47563 a_35502_24538.n132 a_35502_24538.n56 2.69513
R47564 a_35502_24538.n78 a_35502_24538.n76 2.4256
R47565 a_35502_24538.n23 a_35502_24538.n78 2.42484
R47566 a_35502_24538.n31 a_35502_24538.n64 2.43326
R47567 a_35502_24538.n38 a_35502_24538.n135 2.32949
R47568 a_35502_24538.n129 a_35502_24538.n100 2.30989
R47569 a_35502_24538.n54 a_35502_24538.n53 2.30818
R47570 a_35502_24538.n141 a_35502_24538.n140 2.24481
R47571 a_35502_24538.n55 a_35502_24538.n54 2.2442
R47572 a_35502_24538.n52 a_35502_24538.n51 2.24358
R47573 a_35502_24538.n74 a_35502_24538.n71 2.23529
R47574 a_35502_24538.n66 a_35502_24538.n63 2.23423
R47575 a_35502_24538.n100 a_35502_24538.n80 2.18975
R47576 a_35502_24538.n128 a_35502_24538.n101 2.16725
R47577 a_35502_24538.n26 a_35502_24538.n5 2.4981
R47578 a_35502_24538.n130 a_35502_24538.n79 2.07557
R47579 a_35502_24538.n79 a_35502_24538.n25 2.07182
R47580 a_35502_24538.n25 a_35502_24538.n15 2.4644
R47581 a_35502_24538.n61 a_35502_24538.n60 1.7613
R47582 a_35502_24538.n59 a_35502_24538.n57 1.55888
R47583 a_35502_24538.n79 a_35502_24538.n26 1.5005
R47584 a_35502_24538.n129 a_35502_24538.n128 1.5005
R47585 a_35502_24538.n59 a_35502_24538.n58 1.5005
R47586 a_35502_24538.n62 a_35502_24538.n61 1.5005
R47587 a_35502_24538.n133 a_35502_24538.n132 1.5005
R47588 a_35502_24538.n138 a_35502_24538.t21 1.4705
R47589 a_35502_24538.n138 a_35502_24538.t13 1.4705
R47590 a_35502_24538.n48 a_35502_24538.t2 1.4705
R47591 a_35502_24538.n48 a_35502_24538.t20 1.4705
R47592 a_35502_24538.n45 a_35502_24538.t22 1.4705
R47593 a_35502_24538.n45 a_35502_24538.t16 1.4705
R47594 a_35502_24538.n53 a_35502_24538.t10 1.4705
R47595 a_35502_24538.n53 a_35502_24538.t19 1.4705
R47596 a_35502_24538.n135 a_35502_24538.t8 1.4705
R47597 a_35502_24538.n135 a_35502_24538.t18 1.4705
R47598 a_35502_24538.n136 a_35502_24538.t14 1.4705
R47599 a_35502_24538.n136 a_35502_24538.t5 1.4705
R47600 a_35502_24538.n83 a_35502_24538.n82 1.39514
R47601 a_35502_24538.n120 a_35502_24538.n117 1.39105
R47602 a_35502_24538.n130 a_35502_24538.n129 1.35453
R47603 a_35502_24538.n47 a_35502_24538.n46 1.27228
R47604 a_35502_24538.n93 a_35502_24538.n92 1.26997
R47605 a_35502_24538.n0 a_35502_24538.n95 1.24392
R47606 a_35502_24538.n113 a_35502_24538.n112 1.24204
R47607 a_35502_24538.n140 a_35502_24538.n137 1.20603
R47608 a_35502_24538.n126 a_35502_24538.n115 1.20414
R47609 a_35502_24538.n99 a_35502_24538.n98 1.14132
R47610 a_35502_24538.n55 a_35502_24538.n52 1.13952
R47611 a_35502_24538.n107 a_35502_24538.n104 1.13598
R47612 a_35502_24538.n37 a_35502_24538.n49 1.20574
R47613 a_35502_24538.n42 a_35502_24538.n34 1.24017
R47614 a_35502_24538.n132 a_35502_24538.n131 0.963743
R47615 a_35502_24538.n49 a_35502_24538.n47 0.937067
R47616 a_35502_24538.n100 a_35502_24538.n1 0.888471
R47617 a_35502_24538.n128 a_35502_24538.n127 0.71825
R47618 a_35502_24538.n94 a_35502_24538.n93 0.663658
R47619 a_35502_24538.n95 a_35502_24538.n94 0.663658
R47620 a_35502_24538.n115 a_35502_24538.n114 0.655156
R47621 a_35502_24538.n114 a_35502_24538.n113 0.655156
R47622 a_35502_24538.n118 a_35502_24538.n117 0.439529
R47623 a_35502_24538.n84 a_35502_24538.n83 0.432797
R47624 a_35502_24538.n123 a_35502_24538.n116 0.379447
R47625 a_35502_24538.n106 a_35502_24538.n103 0.379447
R47626 a_35502_24538.n65 a_35502_24538.n19 0.745981
R47627 a_35502_24538.n9 a_35502_24538.n72 0.745252
R47628 a_35502_24538.n8 a_35502_24538.n73 0.745252
R47629 a_35502_24538.n1 a_35502_24538.n99 0.498861
R47630 a_35502_24538.n67 a_35502_24538.n12 0.756573
R47631 a_35502_24538.n18 a_35502_24538.n64 0.756388
R47632 a_35502_24538.n15 a_35502_24538.n70 0.756711
R47633 a_35502_24538.n75 a_35502_24538.n22 0.756011
R47634 a_35502_24538.n108 a_35502_24538.n107 0.3605
R47635 a_35502_24538.n122 a_35502_24538.n121 0.3605
R47636 a_35502_24538.n98 a_35502_24538.n97 0.335806
R47637 a_35502_24538.n105 a_35502_24538.n104 0.33475
R47638 a_35502_24538.n86 a_35502_24538.n81 0.302474
R47639 a_35502_24538.n88 a_35502_24538.n87 0.287375
R47640 a_35502_24538.n131 a_35502_24538.n62 0.277797
R47641 a_35502_24538.n67 a_35502_24538.n66 0.208888
R47642 a_35502_24538.n75 a_35502_24538.n74 0.20887
R47643 a_35502_24538.n52 a_35502_24538.n44 0.208394
R47644 a_35502_24538.n140 a_35502_24538.n139 0.208357
R47645 a_35502_24538.n62 a_35502_24538.n59 0.168946
R47646 a_35502_24538.n37 a_35502_24538.n44 0.233116
R47647 a_35502_24538.n86 a_35502_24538.n85 0.147342
R47648 a_35502_24538.n90 a_35502_24538.n81 0.147342
R47649 a_35502_24538.n126 a_35502_24538.n125 0.147342
R47650 a_35502_24538.n119 a_35502_24538.n116 0.147342
R47651 a_35502_24538.n110 a_35502_24538.n103 0.147342
R47652 a_35502_24538.n139 a_35502_24538.n42 0.211956
R47653 a_35502_24538.n41 a_35502_24538.n40 0.142388
R47654 a_35502_24538.n56 a_35502_24538.n43 0.14
R47655 a_35502_24538.n66 a_35502_24538.n19 1.12746
R47656 a_35502_24538.n14 a_35502_24538.n12 1.49123
R47657 a_35502_24538.n14 a_35502_24538.n24 0.772202
R47658 a_35502_24538.n18 a_35502_24538.n25 1.21369
R47659 a_35502_24538.n70 a_35502_24538.n27 2.42126
R47660 a_35502_24538.n74 a_35502_24538.n9 1.12837
R47661 a_35502_24538.n4 a_35502_24538.n22 1.49118
R47662 a_35502_24538.n76 a_35502_24538.n4 0.772883
R47663 a_35502_24538.n8 a_35502_24538.n26 1.21186
R47664 a_35502_24538.n5 a_35502_24538.n23 0.772883
R47665 a_35502_24538.n87 a_35502_24538.n82 0.14
R47666 a_35502_24538.n89 a_35502_24538.n88 0.14
R47667 a_35502_24538.n89 a_35502_24538.n80 0.14
R47668 a_35502_24538.n109 a_35502_24538.n108 0.14
R47669 a_35502_24538.n109 a_35502_24538.n101 0.14
R47670 a_35502_24538.n127 a_35502_24538.n102 0.14
R47671 a_35502_24538.n122 a_35502_24538.n102 0.14
R47672 a_35502_24538.n121 a_35502_24538.n120 0.14
R47673 a_35502_24538.n35 a_35502_24538.n39 1.19679
R47674 a_35502_24538.n137 a_35502_24538.n35 0.932624
R47675 a_35502_24538.t4 a_35502_24538.n34 6.53226
R47676 a_35502_24538.n112 a_35502_24538.n111 0.137868
R47677 a_35502_24538.n50 a_35502_24538.n36 0.137318
R47678 a_35502_24538.n134 a_35502_24538.n133 0.131
R47679 a_35502_24538.n97 a_35502_24538.n96 0.128395
R47680 a_35502_24538.n106 a_35502_24538.n105 0.128395
R47681 a_35502_24538.n124 a_35502_24538.n123 0.118921
R47682 a_35502_24538.n92 a_35502_24538.n91 0.114184
R47683 a_35502_24538.n51 a_35502_24538.n50 0.110782
R47684 a_35502_24538.n141 a_35502_24538.n40 0.105711
R47685 a_35502_24538.n56 a_35502_24538.n55 0.0688756
R47686 a_35502_24538.n32 a_35502_24538.n6 0.0402153
R47687 a_35502_24538.n85 a_35502_24538.n84 0.0348421
R47688 a_35502_24538.n20 a_35502_24538.n71 0.0344623
R47689 a_35502_24538.n91 a_35502_24538.n90 0.0336579
R47690 a_35502_24538.n10 a_35502_24538.n63 0.0325285
R47691 a_35502_24538.n30 a_35502_24538.n29 0.0299662
R47692 a_35502_24538.n125 a_35502_24538.n124 0.0289211
R47693 a_35502_24538.n2 a_35502_24538.n77 0.0283648
R47694 a_35502_24538.n68 a_35502_24538.n28 0.0258025
R47695 a_35502_24538.n78 a_35502_24538.n77 0.0226397
R47696 a_35502_24538.n119 a_35502_24538.n118 0.0194474
R47697 a_35502_24538.n69 a_35502_24538.n68 0.0149128
R47698 a_35502_24538.n16 a_35502_24538.n29 0.0107491
R47699 a_35502_24538.n111 a_35502_24538.n110 0.00997368
R47700 a_35502_24538.n133 a_35502_24538.n39 0.0777922
R47701 a_35502_24538.n24 a_35502_24538.n27 2.43637
R47702 a_35502_24538.n0 a_35502_24538.n96 0.6755
R47703 a_35502_24538.n3 a_35502_24538.n2 0.369148
R47704 a_35502_24538.n69 a_35502_24538.n13 0.354735
R47705 a_35502_24538.n7 a_35502_24538.n6 0.347689
R47706 a_35502_24538.n17 a_35502_24538.n16 0.347689
R47707 a_35502_24538.n21 a_35502_24538.n20 0.346915
R47708 a_35502_24538.n11 a_35502_24538.n10 0.32719
R47709 a_41891_4481.n1 a_41891_4481.t4 10.2515
R47710 a_41891_4481.n1 a_41891_4481.t6 10.2515
R47711 a_41891_4481.n1 a_41891_4481.t22 10.2515
R47712 a_41891_4481.n1 a_41891_4481.t16 10.2515
R47713 a_41891_4481.n1 a_41891_4481.t0 10.096
R47714 a_41891_4481.n1 a_41891_4481.t21 10.0935
R47715 a_41891_4481.n1 a_41891_4481.t2 10.0859
R47716 a_41891_4481.n1 a_41891_4481.t15 10.0808
R47717 a_41891_4481.n1 a_41891_4481.t18 9.53981
R47718 a_41891_4481.n1 a_41891_4481.t14 9.53981
R47719 a_41891_4481.n1 a_41891_4481.t20 9.53981
R47720 a_41891_4481.n1 a_41891_4481.t12 9.53981
R47721 a_41891_4481.n1 a_41891_4481.t17 9.53744
R47722 a_41891_4481.n1 a_41891_4481.t13 9.53744
R47723 a_41891_4481.n1 a_41891_4481.t19 9.53744
R47724 a_41891_4481.n1 a_41891_4481.t11 9.53744
R47725 a_41891_4481.n1 a_41891_4481.n0 8.41434
R47726 a_41891_4481.n1 a_41891_4481.t5 8.14082
R47727 a_41891_4481.n0 a_41891_4481.t7 8.13828
R47728 a_41891_4481.t8 a_41891_4481.t10 7.96115
R47729 a_41891_4481.t8 a_41891_4481.t9 7.94694
R47730 a_41891_4481.t8 a_41891_4481.n1 7.50666
R47731 a_41891_4481.n0 a_41891_4481.t1 7.48586
R47732 a_41891_4481.n1 a_41891_4481.t3 7.48333
R47733 a_71281_n8397.n1 a_71281_n8397.n585 13.5116
R47734 a_71281_n8397.n585 a_71281_n8397.t1 10.674
R47735 a_71281_n8397.n710 a_71281_n8397.t89 10.5154
R47736 a_71281_n8397.t89 a_71281_n8397.n705 10.5154
R47737 a_71281_n8397.n724 a_71281_n8397.t163 10.5154
R47738 a_71281_n8397.t163 a_71281_n8397.n719 10.5154
R47739 a_71281_n8397.t83 a_71281_n8397.n802 10.5154
R47740 a_71281_n8397.n806 a_71281_n8397.t83 10.5154
R47741 a_71281_n8397.t156 a_71281_n8397.n789 10.5154
R47742 a_71281_n8397.n793 a_71281_n8397.t156 10.5154
R47743 a_71281_n8397.t120 a_71281_n8397.n588 10.5154
R47744 a_71281_n8397.n592 a_71281_n8397.t120 10.5154
R47745 a_71281_n8397.t195 a_71281_n8397.n601 10.5154
R47746 a_71281_n8397.n605 a_71281_n8397.t195 10.5154
R47747 a_71281_n8397.t182 a_71281_n8397.n615 10.5154
R47748 a_71281_n8397.n619 a_71281_n8397.t182 10.5154
R47749 a_71281_n8397.t251 a_71281_n8397.n629 10.5154
R47750 a_71281_n8397.n633 a_71281_n8397.t251 10.5154
R47751 a_71281_n8397.t241 a_71281_n8397.n646 10.5154
R47752 a_71281_n8397.n650 a_71281_n8397.t241 10.5154
R47753 a_71281_n8397.t308 a_71281_n8397.n660 10.5154
R47754 a_71281_n8397.n664 a_71281_n8397.t308 10.5154
R47755 a_71281_n8397.t287 a_71281_n8397.n677 10.5154
R47756 a_71281_n8397.n681 a_71281_n8397.t287 10.5154
R47757 a_71281_n8397.t100 a_71281_n8397.n691 10.5154
R47758 a_71281_n8397.n695 a_71281_n8397.t100 10.5154
R47759 a_71281_n8397.n126 a_71281_n8397.t318 10.5154
R47760 a_71281_n8397.t318 a_71281_n8397.n121 10.5154
R47761 a_71281_n8397.n140 a_71281_n8397.t131 10.5154
R47762 a_71281_n8397.t131 a_71281_n8397.n135 10.5154
R47763 a_71281_n8397.t200 a_71281_n8397.n162 10.5154
R47764 a_71281_n8397.n166 a_71281_n8397.t200 10.5154
R47765 a_71281_n8397.t264 a_71281_n8397.n149 10.5154
R47766 a_71281_n8397.n153 a_71281_n8397.t264 10.5154
R47767 a_71281_n8397.t81 a_71281_n8397.n4 10.5154
R47768 a_71281_n8397.n8 a_71281_n8397.t81 10.5154
R47769 a_71281_n8397.t154 a_71281_n8397.n17 10.5154
R47770 a_71281_n8397.n21 a_71281_n8397.t154 10.5154
R47771 a_71281_n8397.t151 a_71281_n8397.n31 10.5154
R47772 a_71281_n8397.n35 a_71281_n8397.t151 10.5154
R47773 a_71281_n8397.t222 a_71281_n8397.n45 10.5154
R47774 a_71281_n8397.n49 a_71281_n8397.t222 10.5154
R47775 a_71281_n8397.t214 a_71281_n8397.n62 10.5154
R47776 a_71281_n8397.n66 a_71281_n8397.t214 10.5154
R47777 a_71281_n8397.t281 a_71281_n8397.n76 10.5154
R47778 a_71281_n8397.n80 a_71281_n8397.t281 10.5154
R47779 a_71281_n8397.t261 a_71281_n8397.n93 10.5154
R47780 a_71281_n8397.n97 a_71281_n8397.t261 10.5154
R47781 a_71281_n8397.t326 a_71281_n8397.n107 10.5154
R47782 a_71281_n8397.n111 a_71281_n8397.t326 10.5154
R47783 a_71281_n8397.n285 a_71281_n8397.t143 10.5154
R47784 a_71281_n8397.t143 a_71281_n8397.n280 10.5154
R47785 a_71281_n8397.n271 a_71281_n8397.t215 10.5154
R47786 a_71281_n8397.t215 a_71281_n8397.n266 10.5154
R47787 a_71281_n8397.n257 a_71281_n8397.t198 10.5154
R47788 a_71281_n8397.t198 a_71281_n8397.n252 10.5154
R47789 a_71281_n8397.n243 a_71281_n8397.t204 10.5154
R47790 a_71281_n8397.t204 a_71281_n8397.n238 10.5154
R47791 a_71281_n8397.n226 a_71281_n8397.t197 10.5154
R47792 a_71281_n8397.t197 a_71281_n8397.n221 10.5154
R47793 a_71281_n8397.n212 a_71281_n8397.t262 10.5154
R47794 a_71281_n8397.t262 a_71281_n8397.n207 10.5154
R47795 a_71281_n8397.n195 a_71281_n8397.t253 10.5154
R47796 a_71281_n8397.t253 a_71281_n8397.n190 10.5154
R47797 a_71281_n8397.n181 a_71281_n8397.t319 10.5154
R47798 a_71281_n8397.t319 a_71281_n8397.n176 10.5154
R47799 a_71281_n8397.n417 a_71281_n8397.t97 10.5154
R47800 a_71281_n8397.t97 a_71281_n8397.n412 10.5154
R47801 a_71281_n8397.n431 a_71281_n8397.t170 10.5154
R47802 a_71281_n8397.t170 a_71281_n8397.n426 10.5154
R47803 a_71281_n8397.t101 a_71281_n8397.n453 10.5154
R47804 a_71281_n8397.n457 a_71281_n8397.t101 10.5154
R47805 a_71281_n8397.t173 a_71281_n8397.n440 10.5154
R47806 a_71281_n8397.n444 a_71281_n8397.t173 10.5154
R47807 a_71281_n8397.t126 a_71281_n8397.n295 10.5154
R47808 a_71281_n8397.n299 a_71281_n8397.t126 10.5154
R47809 a_71281_n8397.t201 a_71281_n8397.n308 10.5154
R47810 a_71281_n8397.n312 a_71281_n8397.t201 10.5154
R47811 a_71281_n8397.t192 a_71281_n8397.n322 10.5154
R47812 a_71281_n8397.n326 a_71281_n8397.t192 10.5154
R47813 a_71281_n8397.t260 a_71281_n8397.n336 10.5154
R47814 a_71281_n8397.n340 a_71281_n8397.t260 10.5154
R47815 a_71281_n8397.t248 a_71281_n8397.n353 10.5154
R47816 a_71281_n8397.n357 a_71281_n8397.t248 10.5154
R47817 a_71281_n8397.t316 a_71281_n8397.n367 10.5154
R47818 a_71281_n8397.n371 a_71281_n8397.t316 10.5154
R47819 a_71281_n8397.t293 a_71281_n8397.n384 10.5154
R47820 a_71281_n8397.n388 a_71281_n8397.t293 10.5154
R47821 a_71281_n8397.t110 a_71281_n8397.n398 10.5154
R47822 a_71281_n8397.n402 a_71281_n8397.t110 10.5154
R47823 a_71281_n8397.n576 a_71281_n8397.t304 10.5154
R47824 a_71281_n8397.t304 a_71281_n8397.n571 10.5154
R47825 a_71281_n8397.n562 a_71281_n8397.t123 10.5154
R47826 a_71281_n8397.t123 a_71281_n8397.n557 10.5154
R47827 a_71281_n8397.n548 a_71281_n8397.t95 10.5154
R47828 a_71281_n8397.t95 a_71281_n8397.n543 10.5154
R47829 a_71281_n8397.n534 a_71281_n8397.t108 10.5154
R47830 a_71281_n8397.t108 a_71281_n8397.n529 10.5154
R47831 a_71281_n8397.n517 a_71281_n8397.t94 10.5154
R47832 a_71281_n8397.t94 a_71281_n8397.n512 10.5154
R47833 a_71281_n8397.n503 a_71281_n8397.t168 10.5154
R47834 a_71281_n8397.t168 a_71281_n8397.n498 10.5154
R47835 a_71281_n8397.n486 a_71281_n8397.t162 10.5154
R47836 a_71281_n8397.t162 a_71281_n8397.n481 10.5154
R47837 a_71281_n8397.n472 a_71281_n8397.t232 10.5154
R47838 a_71281_n8397.t232 a_71281_n8397.n467 10.5154
R47839 a_71281_n8397.t290 a_71281_n8397.n733 10.5154
R47840 a_71281_n8397.n737 a_71281_n8397.t290 10.5154
R47841 a_71281_n8397.t104 a_71281_n8397.n747 10.5154
R47842 a_71281_n8397.n751 a_71281_n8397.t104 10.5154
R47843 a_71281_n8397.t79 a_71281_n8397.n761 10.5154
R47844 a_71281_n8397.n765 a_71281_n8397.t79 10.5154
R47845 a_71281_n8397.t87 a_71281_n8397.n775 10.5154
R47846 a_71281_n8397.n779 a_71281_n8397.t87 10.5154
R47847 a_71281_n8397.n866 a_71281_n8397.t78 10.5154
R47848 a_71281_n8397.t78 a_71281_n8397.n861 10.5154
R47849 a_71281_n8397.n852 a_71281_n8397.t153 10.5154
R47850 a_71281_n8397.t153 a_71281_n8397.n847 10.5154
R47851 a_71281_n8397.n835 a_71281_n8397.t149 10.5154
R47852 a_71281_n8397.t149 a_71281_n8397.n830 10.5154
R47853 a_71281_n8397.n821 a_71281_n8397.t220 10.5154
R47854 a_71281_n8397.t220 a_71281_n8397.n816 10.5154
R47855 a_71281_n8397.n589 a_71281_n8397.t206 10.515
R47856 a_71281_n8397.n5 a_71281_n8397.t269 10.515
R47857 a_71281_n8397.n282 a_71281_n8397.t312 10.515
R47858 a_71281_n8397.n296 a_71281_n8397.t226 10.515
R47859 a_71281_n8397.n573 a_71281_n8397.t225 10.515
R47860 a_71281_n8397.n734 a_71281_n8397.t223 10.515
R47861 a_71281_n8397.n706 a_71281_n8397.t176 10.515
R47862 a_71281_n8397.n707 a_71281_n8397.t176 10.515
R47863 a_71281_n8397.n720 a_71281_n8397.t245 10.515
R47864 a_71281_n8397.n721 a_71281_n8397.t245 10.515
R47865 a_71281_n8397.n804 a_71281_n8397.t273 10.515
R47866 a_71281_n8397.n803 a_71281_n8397.t273 10.515
R47867 a_71281_n8397.n791 a_71281_n8397.t337 10.515
R47868 a_71281_n8397.n790 a_71281_n8397.t337 10.515
R47869 a_71281_n8397.n590 a_71281_n8397.t206 10.515
R47870 a_71281_n8397.n603 a_71281_n8397.t270 10.515
R47871 a_71281_n8397.n602 a_71281_n8397.t270 10.515
R47872 a_71281_n8397.n617 a_71281_n8397.t263 10.515
R47873 a_71281_n8397.n616 a_71281_n8397.t263 10.515
R47874 a_71281_n8397.n631 a_71281_n8397.t329 10.515
R47875 a_71281_n8397.n630 a_71281_n8397.t329 10.515
R47876 a_71281_n8397.n648 a_71281_n8397.t322 10.515
R47877 a_71281_n8397.n647 a_71281_n8397.t322 10.515
R47878 a_71281_n8397.n662 a_71281_n8397.t137 10.515
R47879 a_71281_n8397.n661 a_71281_n8397.t137 10.515
R47880 a_71281_n8397.n679 a_71281_n8397.t115 10.515
R47881 a_71281_n8397.n678 a_71281_n8397.t115 10.515
R47882 a_71281_n8397.n693 a_71281_n8397.t185 10.515
R47883 a_71281_n8397.n692 a_71281_n8397.t185 10.515
R47884 a_71281_n8397.n122 a_71281_n8397.t242 10.515
R47885 a_71281_n8397.n123 a_71281_n8397.t242 10.515
R47886 a_71281_n8397.n136 a_71281_n8397.t309 10.515
R47887 a_71281_n8397.n137 a_71281_n8397.t309 10.515
R47888 a_71281_n8397.n164 a_71281_n8397.t111 10.515
R47889 a_71281_n8397.n163 a_71281_n8397.t111 10.515
R47890 a_71281_n8397.n151 a_71281_n8397.t178 10.515
R47891 a_71281_n8397.n150 a_71281_n8397.t178 10.515
R47892 a_71281_n8397.n6 a_71281_n8397.t269 10.515
R47893 a_71281_n8397.n19 a_71281_n8397.t335 10.515
R47894 a_71281_n8397.n18 a_71281_n8397.t335 10.515
R47895 a_71281_n8397.n33 a_71281_n8397.t328 10.515
R47896 a_71281_n8397.n32 a_71281_n8397.t328 10.515
R47897 a_71281_n8397.n47 a_71281_n8397.t141 10.515
R47898 a_71281_n8397.n46 a_71281_n8397.t141 10.515
R47899 a_71281_n8397.n64 a_71281_n8397.t134 10.515
R47900 a_71281_n8397.n63 a_71281_n8397.t134 10.515
R47901 a_71281_n8397.n78 a_71281_n8397.t210 10.515
R47902 a_71281_n8397.n77 a_71281_n8397.t210 10.515
R47903 a_71281_n8397.n95 a_71281_n8397.t184 10.515
R47904 a_71281_n8397.n94 a_71281_n8397.t184 10.515
R47905 a_71281_n8397.n109 a_71281_n8397.t252 10.515
R47906 a_71281_n8397.n108 a_71281_n8397.t252 10.515
R47907 a_71281_n8397.n281 a_71281_n8397.t312 10.515
R47908 a_71281_n8397.n267 a_71281_n8397.t129 10.515
R47909 a_71281_n8397.n268 a_71281_n8397.t129 10.515
R47910 a_71281_n8397.n253 a_71281_n8397.t105 10.515
R47911 a_71281_n8397.n254 a_71281_n8397.t105 10.515
R47912 a_71281_n8397.n239 a_71281_n8397.t116 10.515
R47913 a_71281_n8397.n240 a_71281_n8397.t116 10.515
R47914 a_71281_n8397.n222 a_71281_n8397.t103 10.515
R47915 a_71281_n8397.n223 a_71281_n8397.t103 10.515
R47916 a_71281_n8397.n208 a_71281_n8397.t177 10.515
R47917 a_71281_n8397.n209 a_71281_n8397.t177 10.515
R47918 a_71281_n8397.n191 a_71281_n8397.t164 10.515
R47919 a_71281_n8397.n192 a_71281_n8397.t164 10.515
R47920 a_71281_n8397.n177 a_71281_n8397.t236 10.515
R47921 a_71281_n8397.n178 a_71281_n8397.t236 10.515
R47922 a_71281_n8397.n413 a_71281_n8397.t207 10.515
R47923 a_71281_n8397.n414 a_71281_n8397.t207 10.515
R47924 a_71281_n8397.n427 a_71281_n8397.t274 10.515
R47925 a_71281_n8397.n428 a_71281_n8397.t274 10.515
R47926 a_71281_n8397.n455 a_71281_n8397.t276 10.515
R47927 a_71281_n8397.n454 a_71281_n8397.t276 10.515
R47928 a_71281_n8397.n442 a_71281_n8397.t75 10.515
R47929 a_71281_n8397.n441 a_71281_n8397.t75 10.515
R47930 a_71281_n8397.n297 a_71281_n8397.t226 10.515
R47931 a_71281_n8397.n310 a_71281_n8397.t289 10.515
R47932 a_71281_n8397.n309 a_71281_n8397.t289 10.515
R47933 a_71281_n8397.n324 a_71281_n8397.t283 10.515
R47934 a_71281_n8397.n323 a_71281_n8397.t283 10.515
R47935 a_71281_n8397.n338 a_71281_n8397.t90 10.515
R47936 a_71281_n8397.n337 a_71281_n8397.t90 10.515
R47937 a_71281_n8397.n355 a_71281_n8397.t85 10.515
R47938 a_71281_n8397.n354 a_71281_n8397.t85 10.515
R47939 a_71281_n8397.n369 a_71281_n8397.t158 10.515
R47940 a_71281_n8397.n368 a_71281_n8397.t158 10.515
R47941 a_71281_n8397.n386 a_71281_n8397.t139 10.515
R47942 a_71281_n8397.n385 a_71281_n8397.t139 10.515
R47943 a_71281_n8397.n400 a_71281_n8397.t213 10.515
R47944 a_71281_n8397.n399 a_71281_n8397.t213 10.515
R47945 a_71281_n8397.n572 a_71281_n8397.t225 10.515
R47946 a_71281_n8397.n558 a_71281_n8397.t285 10.515
R47947 a_71281_n8397.n559 a_71281_n8397.t285 10.515
R47948 a_71281_n8397.n544 a_71281_n8397.t272 10.515
R47949 a_71281_n8397.n545 a_71281_n8397.t272 10.515
R47950 a_71281_n8397.n530 a_71281_n8397.t280 10.515
R47951 a_71281_n8397.n531 a_71281_n8397.t280 10.515
R47952 a_71281_n8397.n513 a_71281_n8397.t271 10.515
R47953 a_71281_n8397.n514 a_71281_n8397.t271 10.515
R47954 a_71281_n8397.n499 a_71281_n8397.t336 10.515
R47955 a_71281_n8397.n500 a_71281_n8397.t336 10.515
R47956 a_71281_n8397.n482 a_71281_n8397.t330 10.515
R47957 a_71281_n8397.n483 a_71281_n8397.t330 10.515
R47958 a_71281_n8397.n468 a_71281_n8397.t142 10.515
R47959 a_71281_n8397.n469 a_71281_n8397.t142 10.515
R47960 a_71281_n8397.n735 a_71281_n8397.t223 10.515
R47961 a_71281_n8397.n749 a_71281_n8397.t284 10.515
R47962 a_71281_n8397.n748 a_71281_n8397.t284 10.515
R47963 a_71281_n8397.n763 a_71281_n8397.t267 10.515
R47964 a_71281_n8397.n762 a_71281_n8397.t267 10.515
R47965 a_71281_n8397.n777 a_71281_n8397.t279 10.515
R47966 a_71281_n8397.n776 a_71281_n8397.t279 10.515
R47967 a_71281_n8397.n862 a_71281_n8397.t266 10.515
R47968 a_71281_n8397.n863 a_71281_n8397.t266 10.515
R47969 a_71281_n8397.n848 a_71281_n8397.t334 10.515
R47970 a_71281_n8397.n849 a_71281_n8397.t334 10.515
R47971 a_71281_n8397.n831 a_71281_n8397.t327 10.515
R47972 a_71281_n8397.n832 a_71281_n8397.t327 10.515
R47973 a_71281_n8397.n817 a_71281_n8397.t140 10.515
R47974 a_71281_n8397.n818 a_71281_n8397.t140 10.515
R47975 a_71281_n8397.n710 a_71281_n8397.t296 9.57886
R47976 a_71281_n8397.t296 a_71281_n8397.n705 9.57886
R47977 a_71281_n8397.n707 a_71281_n8397.t228 9.57886
R47978 a_71281_n8397.t228 a_71281_n8397.n706 9.57886
R47979 a_71281_n8397.n724 a_71281_n8397.t112 9.57886
R47980 a_71281_n8397.t112 a_71281_n8397.n719 9.57886
R47981 a_71281_n8397.n721 a_71281_n8397.t297 9.57886
R47982 a_71281_n8397.t297 a_71281_n8397.n720 9.57886
R47983 a_71281_n8397.t186 a_71281_n8397.n802 9.57886
R47984 a_71281_n8397.n806 a_71281_n8397.t186 9.57886
R47985 a_71281_n8397.t174 a_71281_n8397.n803 9.57886
R47986 a_71281_n8397.n804 a_71281_n8397.t174 9.57886
R47987 a_71281_n8397.t254 a_71281_n8397.n789 9.57886
R47988 a_71281_n8397.n793 a_71281_n8397.t254 9.57886
R47989 a_71281_n8397.t243 a_71281_n8397.n790 9.57886
R47990 a_71281_n8397.n791 a_71281_n8397.t243 9.57886
R47991 a_71281_n8397.t321 a_71281_n8397.n588 9.57886
R47992 a_71281_n8397.n592 a_71281_n8397.t321 9.57886
R47993 a_71281_n8397.t256 a_71281_n8397.n589 9.57886
R47994 a_71281_n8397.n590 a_71281_n8397.t256 9.57886
R47995 a_71281_n8397.t136 a_71281_n8397.n601 9.57886
R47996 a_71281_n8397.n605 a_71281_n8397.t136 9.57886
R47997 a_71281_n8397.t323 a_71281_n8397.n602 9.57886
R47998 a_71281_n8397.n603 a_71281_n8397.t323 9.57886
R47999 a_71281_n8397.t128 a_71281_n8397.n615 9.57886
R48000 a_71281_n8397.n619 a_71281_n8397.t128 9.57886
R48001 a_71281_n8397.t313 a_71281_n8397.n616 9.57886
R48002 a_71281_n8397.n617 a_71281_n8397.t313 9.57886
R48003 a_71281_n8397.t203 a_71281_n8397.n629 9.57886
R48004 a_71281_n8397.n633 a_71281_n8397.t203 9.57886
R48005 a_71281_n8397.t130 a_71281_n8397.n630 9.57886
R48006 a_71281_n8397.n631 a_71281_n8397.t130 9.57886
R48007 a_71281_n8397.t34 a_71281_n8397.n646 9.57886
R48008 a_71281_n8397.n650 a_71281_n8397.t34 9.57886
R48009 a_71281_n8397.t60 a_71281_n8397.n647 9.57886
R48010 a_71281_n8397.n648 a_71281_n8397.t60 9.57886
R48011 a_71281_n8397.t14 a_71281_n8397.n660 9.57886
R48012 a_71281_n8397.n664 a_71281_n8397.t14 9.57886
R48013 a_71281_n8397.t32 a_71281_n8397.n661 9.57886
R48014 a_71281_n8397.n662 a_71281_n8397.t32 9.57886
R48015 a_71281_n8397.t235 a_71281_n8397.n677 9.57886
R48016 a_71281_n8397.n681 a_71281_n8397.t235 9.57886
R48017 a_71281_n8397.t165 a_71281_n8397.n678 9.57886
R48018 a_71281_n8397.n679 a_71281_n8397.t165 9.57886
R48019 a_71281_n8397.t302 a_71281_n8397.n691 9.57886
R48020 a_71281_n8397.n695 a_71281_n8397.t302 9.57886
R48021 a_71281_n8397.t237 a_71281_n8397.n692 9.57886
R48022 a_71281_n8397.n693 a_71281_n8397.t237 9.57886
R48023 a_71281_n8397.n126 a_71281_n8397.t118 9.57886
R48024 a_71281_n8397.t118 a_71281_n8397.n121 9.57886
R48025 a_71281_n8397.n123 a_71281_n8397.t217 9.57886
R48026 a_71281_n8397.t217 a_71281_n8397.n122 9.57886
R48027 a_71281_n8397.n140 a_71281_n8397.t191 9.57886
R48028 a_71281_n8397.t191 a_71281_n8397.n135 9.57886
R48029 a_71281_n8397.n137 a_71281_n8397.t282 9.57886
R48030 a_71281_n8397.t282 a_71281_n8397.n136 9.57886
R48031 a_71281_n8397.t187 a_71281_n8397.n162 9.57886
R48032 a_71281_n8397.n166 a_71281_n8397.t187 9.57886
R48033 a_71281_n8397.t298 a_71281_n8397.n163 9.57886
R48034 a_71281_n8397.n164 a_71281_n8397.t298 9.57886
R48035 a_71281_n8397.t255 a_71281_n8397.n149 9.57886
R48036 a_71281_n8397.n153 a_71281_n8397.t255 9.57886
R48037 a_71281_n8397.t113 a_71281_n8397.n150 9.57886
R48038 a_71281_n8397.n151 a_71281_n8397.t113 9.57886
R48039 a_71281_n8397.t144 a_71281_n8397.n4 9.57886
R48040 a_71281_n8397.n8 a_71281_n8397.t144 9.57886
R48041 a_71281_n8397.t234 a_71281_n8397.n5 9.57886
R48042 a_71281_n8397.n6 a_71281_n8397.t234 9.57886
R48043 a_71281_n8397.t216 a_71281_n8397.n17 9.57886
R48044 a_71281_n8397.n21 a_71281_n8397.t216 9.57886
R48045 a_71281_n8397.t300 a_71281_n8397.n18 9.57886
R48046 a_71281_n8397.n19 a_71281_n8397.t300 9.57886
R48047 a_71281_n8397.t212 a_71281_n8397.n31 9.57886
R48048 a_71281_n8397.n35 a_71281_n8397.t212 9.57886
R48049 a_71281_n8397.t292 a_71281_n8397.n32 9.57886
R48050 a_71281_n8397.n33 a_71281_n8397.t292 9.57886
R48051 a_71281_n8397.t278 a_71281_n8397.n45 9.57886
R48052 a_71281_n8397.n49 a_71281_n8397.t278 9.57886
R48053 a_71281_n8397.t109 a_71281_n8397.n46 9.57886
R48054 a_71281_n8397.n47 a_71281_n8397.t109 9.57886
R48055 a_71281_n8397.t10 a_71281_n8397.n62 9.57886
R48056 a_71281_n8397.n66 a_71281_n8397.t10 9.57886
R48057 a_71281_n8397.t66 a_71281_n8397.n63 9.57886
R48058 a_71281_n8397.n64 a_71281_n8397.t66 9.57886
R48059 a_71281_n8397.t2 a_71281_n8397.n76 9.57886
R48060 a_71281_n8397.n80 a_71281_n8397.t2 9.57886
R48061 a_71281_n8397.t46 a_71281_n8397.n77 9.57886
R48062 a_71281_n8397.n78 a_71281_n8397.t46 9.57886
R48063 a_71281_n8397.t310 a_71281_n8397.n93 9.57886
R48064 a_71281_n8397.n97 a_71281_n8397.t310 9.57886
R48065 a_71281_n8397.t152 a_71281_n8397.n94 9.57886
R48066 a_71281_n8397.n95 a_71281_n8397.t152 9.57886
R48067 a_71281_n8397.t125 a_71281_n8397.n107 9.57886
R48068 a_71281_n8397.n111 a_71281_n8397.t125 9.57886
R48069 a_71281_n8397.t224 a_71281_n8397.n108 9.57886
R48070 a_71281_n8397.n109 a_71281_n8397.t224 9.57886
R48071 a_71281_n8397.n285 a_71281_n8397.t133 9.57886
R48072 a_71281_n8397.t133 a_71281_n8397.n280 9.57886
R48073 a_71281_n8397.n282 a_71281_n8397.t249 9.57886
R48074 a_71281_n8397.t249 a_71281_n8397.n281 9.57886
R48075 a_71281_n8397.n271 a_71281_n8397.t209 9.57886
R48076 a_71281_n8397.t209 a_71281_n8397.n266 9.57886
R48077 a_71281_n8397.n268 a_71281_n8397.t317 9.57886
R48078 a_71281_n8397.t317 a_71281_n8397.n267 9.57886
R48079 a_71281_n8397.n257 a_71281_n8397.t183 9.57886
R48080 a_71281_n8397.t183 a_71281_n8397.n252 9.57886
R48081 a_71281_n8397.n254 a_71281_n8397.t294 9.57886
R48082 a_71281_n8397.t294 a_71281_n8397.n253 9.57886
R48083 a_71281_n8397.n243 a_71281_n8397.t196 9.57886
R48084 a_71281_n8397.t196 a_71281_n8397.n238 9.57886
R48085 a_71281_n8397.n240 a_71281_n8397.t301 9.57886
R48086 a_71281_n8397.t301 a_71281_n8397.n239 9.57886
R48087 a_71281_n8397.n226 a_71281_n8397.t38 9.57886
R48088 a_71281_n8397.t38 a_71281_n8397.n221 9.57886
R48089 a_71281_n8397.n223 a_71281_n8397.t6 9.57886
R48090 a_71281_n8397.t6 a_71281_n8397.n222 9.57886
R48091 a_71281_n8397.n212 a_71281_n8397.t16 9.57886
R48092 a_71281_n8397.t16 a_71281_n8397.n207 9.57886
R48093 a_71281_n8397.n209 a_71281_n8397.t64 9.57886
R48094 a_71281_n8397.t64 a_71281_n8397.n208 9.57886
R48095 a_71281_n8397.n195 a_71281_n8397.t240 9.57886
R48096 a_71281_n8397.t240 a_71281_n8397.n190 9.57886
R48097 a_71281_n8397.n192 a_71281_n8397.t96 9.57886
R48098 a_71281_n8397.t96 a_71281_n8397.n191 9.57886
R48099 a_71281_n8397.n181 a_71281_n8397.t307 9.57886
R48100 a_71281_n8397.t307 a_71281_n8397.n176 9.57886
R48101 a_71281_n8397.n178 a_71281_n8397.t169 9.57886
R48102 a_71281_n8397.t169 a_71281_n8397.n177 9.57886
R48103 a_71281_n8397.n417 a_71281_n8397.t331 9.57886
R48104 a_71281_n8397.t331 a_71281_n8397.n412 9.57886
R48105 a_71281_n8397.n414 a_71281_n8397.t161 9.57886
R48106 a_71281_n8397.t161 a_71281_n8397.n413 9.57886
R48107 a_71281_n8397.n431 a_71281_n8397.t145 9.57886
R48108 a_71281_n8397.t145 a_71281_n8397.n426 9.57886
R48109 a_71281_n8397.n428 a_71281_n8397.t231 9.57886
R48110 a_71281_n8397.t231 a_71281_n8397.n427 9.57886
R48111 a_71281_n8397.t84 a_71281_n8397.n453 9.57886
R48112 a_71281_n8397.n457 a_71281_n8397.t84 9.57886
R48113 a_71281_n8397.t117 a_71281_n8397.n454 9.57886
R48114 a_71281_n8397.n455 a_71281_n8397.t117 9.57886
R48115 a_71281_n8397.t157 a_71281_n8397.n440 9.57886
R48116 a_71281_n8397.n444 a_71281_n8397.t157 9.57886
R48117 a_71281_n8397.t188 a_71281_n8397.n441 9.57886
R48118 a_71281_n8397.n442 a_71281_n8397.t188 9.57886
R48119 a_71281_n8397.t91 a_71281_n8397.n295 9.57886
R48120 a_71281_n8397.n299 a_71281_n8397.t91 9.57886
R48121 a_71281_n8397.t190 a_71281_n8397.n296 9.57886
R48122 a_71281_n8397.n297 a_71281_n8397.t190 9.57886
R48123 a_71281_n8397.t166 a_71281_n8397.n308 9.57886
R48124 a_71281_n8397.n312 a_71281_n8397.t166 9.57886
R48125 a_71281_n8397.t258 a_71281_n8397.n309 9.57886
R48126 a_71281_n8397.n310 a_71281_n8397.t258 9.57886
R48127 a_71281_n8397.t160 a_71281_n8397.n322 9.57886
R48128 a_71281_n8397.n326 a_71281_n8397.t160 9.57886
R48129 a_71281_n8397.t247 a_71281_n8397.n323 9.57886
R48130 a_71281_n8397.n324 a_71281_n8397.t247 9.57886
R48131 a_71281_n8397.t230 a_71281_n8397.n336 9.57886
R48132 a_71281_n8397.n340 a_71281_n8397.t230 9.57886
R48133 a_71281_n8397.t315 a_71281_n8397.n337 9.57886
R48134 a_71281_n8397.n338 a_71281_n8397.t315 9.57886
R48135 a_71281_n8397.t24 a_71281_n8397.n353 9.57886
R48136 a_71281_n8397.n357 a_71281_n8397.t24 9.57886
R48137 a_71281_n8397.t4 a_71281_n8397.n354 9.57886
R48138 a_71281_n8397.n355 a_71281_n8397.t4 9.57886
R48139 a_71281_n8397.t8 a_71281_n8397.n367 9.57886
R48140 a_71281_n8397.n371 a_71281_n8397.t8 9.57886
R48141 a_71281_n8397.t58 a_71281_n8397.n368 9.57886
R48142 a_71281_n8397.n369 a_71281_n8397.t58 9.57886
R48143 a_71281_n8397.t275 a_71281_n8397.n384 9.57886
R48144 a_71281_n8397.n388 a_71281_n8397.t275 9.57886
R48145 a_71281_n8397.t93 a_71281_n8397.n385 9.57886
R48146 a_71281_n8397.n386 a_71281_n8397.t93 9.57886
R48147 a_71281_n8397.t74 a_71281_n8397.n398 9.57886
R48148 a_71281_n8397.n402 a_71281_n8397.t74 9.57886
R48149 a_71281_n8397.t167 a_71281_n8397.n399 9.57886
R48150 a_71281_n8397.n400 a_71281_n8397.t167 9.57886
R48151 a_71281_n8397.n576 a_71281_n8397.t291 9.57886
R48152 a_71281_n8397.t291 a_71281_n8397.n571 9.57886
R48153 a_71281_n8397.n573 a_71281_n8397.t320 9.57886
R48154 a_71281_n8397.t320 a_71281_n8397.n572 9.57886
R48155 a_71281_n8397.n562 a_71281_n8397.t106 9.57886
R48156 a_71281_n8397.t106 a_71281_n8397.n557 9.57886
R48157 a_71281_n8397.n559 a_71281_n8397.t135 9.57886
R48158 a_71281_n8397.t135 a_71281_n8397.n558 9.57886
R48159 a_71281_n8397.n548 a_71281_n8397.t80 9.57886
R48160 a_71281_n8397.t80 a_71281_n8397.n543 9.57886
R48161 a_71281_n8397.n545 a_71281_n8397.t114 9.57886
R48162 a_71281_n8397.t114 a_71281_n8397.n544 9.57886
R48163 a_71281_n8397.n534 a_71281_n8397.t88 9.57886
R48164 a_71281_n8397.t88 a_71281_n8397.n529 9.57886
R48165 a_71281_n8397.n531 a_71281_n8397.t122 9.57886
R48166 a_71281_n8397.t122 a_71281_n8397.n530 9.57886
R48167 a_71281_n8397.n517 a_71281_n8397.t70 9.57886
R48168 a_71281_n8397.t70 a_71281_n8397.n512 9.57886
R48169 a_71281_n8397.n514 a_71281_n8397.t62 9.57886
R48170 a_71281_n8397.t62 a_71281_n8397.n513 9.57886
R48171 a_71281_n8397.n503 a_71281_n8397.t50 9.57886
R48172 a_71281_n8397.t50 a_71281_n8397.n498 9.57886
R48173 a_71281_n8397.n500 a_71281_n8397.t36 9.57886
R48174 a_71281_n8397.t36 a_71281_n8397.n499 9.57886
R48175 a_71281_n8397.n486 a_71281_n8397.t150 9.57886
R48176 a_71281_n8397.t150 a_71281_n8397.n481 9.57886
R48177 a_71281_n8397.n483 a_71281_n8397.t175 9.57886
R48178 a_71281_n8397.t175 a_71281_n8397.n482 9.57886
R48179 a_71281_n8397.n472 a_71281_n8397.t221 9.57886
R48180 a_71281_n8397.t221 a_71281_n8397.n467 9.57886
R48181 a_71281_n8397.n469 a_71281_n8397.t244 9.57886
R48182 a_71281_n8397.t244 a_71281_n8397.n468 9.57886
R48183 a_71281_n8397.t132 a_71281_n8397.n733 9.57886
R48184 a_71281_n8397.n737 a_71281_n8397.t132 9.57886
R48185 a_71281_n8397.t124 a_71281_n8397.n734 9.57886
R48186 a_71281_n8397.n735 a_71281_n8397.t124 9.57886
R48187 a_71281_n8397.t208 a_71281_n8397.n747 9.57886
R48188 a_71281_n8397.n751 a_71281_n8397.t208 9.57886
R48189 a_71281_n8397.t199 a_71281_n8397.n748 9.57886
R48190 a_71281_n8397.n749 a_71281_n8397.t199 9.57886
R48191 a_71281_n8397.t181 a_71281_n8397.n761 9.57886
R48192 a_71281_n8397.n765 a_71281_n8397.t181 9.57886
R48193 a_71281_n8397.t171 a_71281_n8397.n762 9.57886
R48194 a_71281_n8397.n763 a_71281_n8397.t171 9.57886
R48195 a_71281_n8397.t194 a_71281_n8397.n775 9.57886
R48196 a_71281_n8397.n779 a_71281_n8397.t194 9.57886
R48197 a_71281_n8397.t179 a_71281_n8397.n776 9.57886
R48198 a_71281_n8397.n777 a_71281_n8397.t179 9.57886
R48199 a_71281_n8397.n866 a_71281_n8397.t40 9.57886
R48200 a_71281_n8397.t40 a_71281_n8397.n861 9.57886
R48201 a_71281_n8397.n863 a_71281_n8397.t44 9.57886
R48202 a_71281_n8397.t44 a_71281_n8397.n862 9.57886
R48203 a_71281_n8397.n852 a_71281_n8397.t18 9.57886
R48204 a_71281_n8397.t18 a_71281_n8397.n847 9.57886
R48205 a_71281_n8397.n849 a_71281_n8397.t22 9.57886
R48206 a_71281_n8397.t22 a_71281_n8397.n848 9.57886
R48207 a_71281_n8397.n835 a_71281_n8397.t239 9.57886
R48208 a_71281_n8397.t239 a_71281_n8397.n830 9.57886
R48209 a_71281_n8397.n832 a_71281_n8397.t233 9.57886
R48210 a_71281_n8397.t233 a_71281_n8397.n831 9.57886
R48211 a_71281_n8397.n821 a_71281_n8397.t306 9.57886
R48212 a_71281_n8397.t306 a_71281_n8397.n816 9.57886
R48213 a_71281_n8397.n818 a_71281_n8397.t299 9.57886
R48214 a_71281_n8397.t299 a_71281_n8397.n817 9.57886
R48215 a_71281_n8397.t238 a_71281_n8397.n712 8.10567
R48216 a_71281_n8397.n713 a_71281_n8397.t238 8.10567
R48217 a_71281_n8397.t305 a_71281_n8397.n726 8.10567
R48218 a_71281_n8397.n727 a_71281_n8397.t305 8.10567
R48219 a_71281_n8397.n810 a_71281_n8397.t82 8.10567
R48220 a_71281_n8397.t82 a_71281_n8397.n809 8.10567
R48221 a_71281_n8397.n796 a_71281_n8397.t155 8.10567
R48222 a_71281_n8397.t155 a_71281_n8397.n795 8.10567
R48223 a_71281_n8397.n595 a_71281_n8397.t265 8.10567
R48224 a_71281_n8397.t265 a_71281_n8397.n594 8.10567
R48225 a_71281_n8397.n609 a_71281_n8397.t333 8.10567
R48226 a_71281_n8397.t333 a_71281_n8397.n608 8.10567
R48227 a_71281_n8397.n623 a_71281_n8397.t325 8.10567
R48228 a_71281_n8397.t325 a_71281_n8397.n622 8.10567
R48229 a_71281_n8397.n637 a_71281_n8397.t138 8.10567
R48230 a_71281_n8397.t138 a_71281_n8397.n636 8.10567
R48231 a_71281_n8397.n654 a_71281_n8397.t56 8.10567
R48232 a_71281_n8397.t56 a_71281_n8397.n653 8.10567
R48233 a_71281_n8397.n668 a_71281_n8397.t28 8.10567
R48234 a_71281_n8397.t28 a_71281_n8397.n667 8.10567
R48235 a_71281_n8397.n685 a_71281_n8397.t180 8.10567
R48236 a_71281_n8397.t180 a_71281_n8397.n684 8.10567
R48237 a_71281_n8397.n699 a_71281_n8397.t250 8.10567
R48238 a_71281_n8397.t250 a_71281_n8397.n698 8.10567
R48239 a_71281_n8397.t286 a_71281_n8397.n128 8.10567
R48240 a_71281_n8397.n129 a_71281_n8397.t286 8.10567
R48241 a_71281_n8397.t98 a_71281_n8397.n142 8.10567
R48242 a_71281_n8397.n143 a_71281_n8397.t98 8.10567
R48243 a_71281_n8397.n170 a_71281_n8397.t205 8.10567
R48244 a_71281_n8397.t205 a_71281_n8397.n169 8.10567
R48245 a_71281_n8397.n156 a_71281_n8397.t268 8.10567
R48246 a_71281_n8397.t268 a_71281_n8397.n155 8.10567
R48247 a_71281_n8397.n11 a_71281_n8397.t311 8.10567
R48248 a_71281_n8397.t311 a_71281_n8397.n10 8.10567
R48249 a_71281_n8397.n25 a_71281_n8397.t127 8.10567
R48250 a_71281_n8397.t127 a_71281_n8397.n24 8.10567
R48251 a_71281_n8397.n39 a_71281_n8397.t119 8.10567
R48252 a_71281_n8397.t119 a_71281_n8397.n38 8.10567
R48253 a_71281_n8397.n53 a_71281_n8397.t193 8.10567
R48254 a_71281_n8397.t193 a_71281_n8397.n52 8.10567
R48255 a_71281_n8397.n70 a_71281_n8397.t42 8.10567
R48256 a_71281_n8397.t42 a_71281_n8397.n69 8.10567
R48257 a_71281_n8397.n84 a_71281_n8397.t20 8.10567
R48258 a_71281_n8397.t20 a_71281_n8397.n83 8.10567
R48259 a_71281_n8397.n101 a_71281_n8397.t227 8.10567
R48260 a_71281_n8397.t227 a_71281_n8397.n100 8.10567
R48261 a_71281_n8397.n115 a_71281_n8397.t295 8.10567
R48262 a_71281_n8397.t295 a_71281_n8397.n114 8.10567
R48263 a_71281_n8397.t148 a_71281_n8397.n287 8.10567
R48264 a_71281_n8397.n288 a_71281_n8397.t148 8.10567
R48265 a_71281_n8397.t219 a_71281_n8397.n273 8.10567
R48266 a_71281_n8397.n274 a_71281_n8397.t219 8.10567
R48267 a_71281_n8397.t202 a_71281_n8397.n259 8.10567
R48268 a_71281_n8397.n260 a_71281_n8397.t202 8.10567
R48269 a_71281_n8397.t211 a_71281_n8397.n245 8.10567
R48270 a_71281_n8397.n246 a_71281_n8397.t211 8.10567
R48271 a_71281_n8397.t30 a_71281_n8397.n228 8.10567
R48272 a_71281_n8397.n229 a_71281_n8397.t30 8.10567
R48273 a_71281_n8397.t12 a_71281_n8397.n214 8.10567
R48274 a_71281_n8397.n215 a_71281_n8397.t12 8.10567
R48275 a_71281_n8397.t259 a_71281_n8397.n197 8.10567
R48276 a_71281_n8397.n198 a_71281_n8397.t259 8.10567
R48277 a_71281_n8397.t324 a_71281_n8397.n183 8.10567
R48278 a_71281_n8397.n184 a_71281_n8397.t324 8.10567
R48279 a_71281_n8397.t246 a_71281_n8397.n419 8.10567
R48280 a_71281_n8397.n420 a_71281_n8397.t246 8.10567
R48281 a_71281_n8397.t314 a_71281_n8397.n433 8.10567
R48282 a_71281_n8397.n434 a_71281_n8397.t314 8.10567
R48283 a_71281_n8397.n461 a_71281_n8397.t99 8.10567
R48284 a_71281_n8397.t99 a_71281_n8397.n460 8.10567
R48285 a_71281_n8397.n447 a_71281_n8397.t172 8.10567
R48286 a_71281_n8397.t172 a_71281_n8397.n446 8.10567
R48287 a_71281_n8397.n302 a_71281_n8397.t277 8.10567
R48288 a_71281_n8397.t277 a_71281_n8397.n301 8.10567
R48289 a_71281_n8397.n316 a_71281_n8397.t76 8.10567
R48290 a_71281_n8397.t76 a_71281_n8397.n315 8.10567
R48291 a_71281_n8397.n330 a_71281_n8397.t332 8.10567
R48292 a_71281_n8397.t332 a_71281_n8397.n329 8.10567
R48293 a_71281_n8397.n344 a_71281_n8397.t146 8.10567
R48294 a_71281_n8397.t146 a_71281_n8397.n343 8.10567
R48295 a_71281_n8397.n361 a_71281_n8397.t54 8.10567
R48296 a_71281_n8397.t54 a_71281_n8397.n360 8.10567
R48297 a_71281_n8397.n375 a_71281_n8397.t26 8.10567
R48298 a_71281_n8397.t26 a_71281_n8397.n374 8.10567
R48299 a_71281_n8397.n392 a_71281_n8397.t189 8.10567
R48300 a_71281_n8397.t189 a_71281_n8397.n391 8.10567
R48301 a_71281_n8397.n406 a_71281_n8397.t257 8.10567
R48302 a_71281_n8397.t257 a_71281_n8397.n405 8.10567
R48303 a_71281_n8397.t303 a_71281_n8397.n578 8.10567
R48304 a_71281_n8397.n579 a_71281_n8397.t303 8.10567
R48305 a_71281_n8397.t121 a_71281_n8397.n564 8.10567
R48306 a_71281_n8397.n565 a_71281_n8397.t121 8.10567
R48307 a_71281_n8397.t92 a_71281_n8397.n550 8.10567
R48308 a_71281_n8397.n551 a_71281_n8397.t92 8.10567
R48309 a_71281_n8397.t107 a_71281_n8397.n536 8.10567
R48310 a_71281_n8397.n537 a_71281_n8397.t107 8.10567
R48311 a_71281_n8397.t68 a_71281_n8397.n519 8.10567
R48312 a_71281_n8397.n520 a_71281_n8397.t68 8.10567
R48313 a_71281_n8397.t48 a_71281_n8397.n505 8.10567
R48314 a_71281_n8397.n506 a_71281_n8397.t48 8.10567
R48315 a_71281_n8397.t159 a_71281_n8397.n488 8.10567
R48316 a_71281_n8397.n489 a_71281_n8397.t159 8.10567
R48317 a_71281_n8397.t229 a_71281_n8397.n474 8.10567
R48318 a_71281_n8397.n475 a_71281_n8397.t229 8.10567
R48319 a_71281_n8397.n741 a_71281_n8397.t288 8.10567
R48320 a_71281_n8397.t288 a_71281_n8397.n740 8.10567
R48321 a_71281_n8397.n755 a_71281_n8397.t102 8.10567
R48322 a_71281_n8397.t102 a_71281_n8397.n754 8.10567
R48323 a_71281_n8397.n769 a_71281_n8397.t77 8.10567
R48324 a_71281_n8397.t77 a_71281_n8397.n768 8.10567
R48325 a_71281_n8397.n783 a_71281_n8397.t86 8.10567
R48326 a_71281_n8397.t86 a_71281_n8397.n782 8.10567
R48327 a_71281_n8397.t72 a_71281_n8397.n868 8.10567
R48328 a_71281_n8397.n869 a_71281_n8397.t72 8.10567
R48329 a_71281_n8397.t52 a_71281_n8397.n854 8.10567
R48330 a_71281_n8397.n855 a_71281_n8397.t52 8.10567
R48331 a_71281_n8397.t147 a_71281_n8397.n837 8.10567
R48332 a_71281_n8397.n838 a_71281_n8397.t147 8.10567
R48333 a_71281_n8397.t218 a_71281_n8397.n823 8.10567
R48334 a_71281_n8397.n824 a_71281_n8397.t218 8.10567
R48335 a_71281_n8397.n585 a_71281_n8397.t0 7.10686
R48336 a_71281_n8397.n673 a_71281_n8397.t15 6.12845
R48337 a_71281_n8397.n843 a_71281_n8397.t19 6.12845
R48338 a_71281_n8397.n89 a_71281_n8397.t3 6.12845
R48339 a_71281_n8397.n203 a_71281_n8397.t17 6.12845
R48340 a_71281_n8397.n380 a_71281_n8397.t9 6.12845
R48341 a_71281_n8397.n494 a_71281_n8397.t51 6.12845
R48342 a_71281_n8397.n874 a_71281_n8397.t45 6.12049
R48343 a_71281_n8397.n642 a_71281_n8397.t61 6.12049
R48344 a_71281_n8397.n58 a_71281_n8397.t67 6.12049
R48345 a_71281_n8397.n234 a_71281_n8397.t7 6.12049
R48346 a_71281_n8397.n349 a_71281_n8397.t5 6.12049
R48347 a_71281_n8397.n525 a_71281_n8397.t63 6.12049
R48348 a_71281_n8397.n712 a_71281_n8397.n708 4.64734
R48349 a_71281_n8397.n713 a_71281_n8397.n704 4.64734
R48350 a_71281_n8397.n726 a_71281_n8397.n722 4.64734
R48351 a_71281_n8397.n727 a_71281_n8397.n718 4.64734
R48352 a_71281_n8397.n810 a_71281_n8397.n801 4.64734
R48353 a_71281_n8397.n809 a_71281_n8397.n805 4.64734
R48354 a_71281_n8397.n796 a_71281_n8397.n788 4.64734
R48355 a_71281_n8397.n795 a_71281_n8397.n792 4.64734
R48356 a_71281_n8397.n595 a_71281_n8397.n587 4.64734
R48357 a_71281_n8397.n594 a_71281_n8397.n591 4.64734
R48358 a_71281_n8397.n609 a_71281_n8397.n600 4.64734
R48359 a_71281_n8397.n608 a_71281_n8397.n604 4.64734
R48360 a_71281_n8397.n623 a_71281_n8397.n614 4.64734
R48361 a_71281_n8397.n622 a_71281_n8397.n618 4.64734
R48362 a_71281_n8397.n637 a_71281_n8397.n628 4.64734
R48363 a_71281_n8397.n636 a_71281_n8397.n632 4.64734
R48364 a_71281_n8397.n654 a_71281_n8397.n645 4.64734
R48365 a_71281_n8397.n653 a_71281_n8397.n649 4.64734
R48366 a_71281_n8397.n668 a_71281_n8397.n659 4.64734
R48367 a_71281_n8397.n667 a_71281_n8397.n663 4.64734
R48368 a_71281_n8397.n685 a_71281_n8397.n676 4.64734
R48369 a_71281_n8397.n684 a_71281_n8397.n680 4.64734
R48370 a_71281_n8397.n699 a_71281_n8397.n690 4.64734
R48371 a_71281_n8397.n698 a_71281_n8397.n694 4.64734
R48372 a_71281_n8397.n128 a_71281_n8397.n124 4.64734
R48373 a_71281_n8397.n129 a_71281_n8397.n120 4.64734
R48374 a_71281_n8397.n142 a_71281_n8397.n138 4.64734
R48375 a_71281_n8397.n143 a_71281_n8397.n134 4.64734
R48376 a_71281_n8397.n170 a_71281_n8397.n161 4.64734
R48377 a_71281_n8397.n169 a_71281_n8397.n165 4.64734
R48378 a_71281_n8397.n156 a_71281_n8397.n148 4.64734
R48379 a_71281_n8397.n155 a_71281_n8397.n152 4.64734
R48380 a_71281_n8397.n11 a_71281_n8397.n3 4.64734
R48381 a_71281_n8397.n10 a_71281_n8397.n7 4.64734
R48382 a_71281_n8397.n25 a_71281_n8397.n16 4.64734
R48383 a_71281_n8397.n24 a_71281_n8397.n20 4.64734
R48384 a_71281_n8397.n39 a_71281_n8397.n30 4.64734
R48385 a_71281_n8397.n38 a_71281_n8397.n34 4.64734
R48386 a_71281_n8397.n53 a_71281_n8397.n44 4.64734
R48387 a_71281_n8397.n52 a_71281_n8397.n48 4.64734
R48388 a_71281_n8397.n70 a_71281_n8397.n61 4.64734
R48389 a_71281_n8397.n69 a_71281_n8397.n65 4.64734
R48390 a_71281_n8397.n84 a_71281_n8397.n75 4.64734
R48391 a_71281_n8397.n83 a_71281_n8397.n79 4.64734
R48392 a_71281_n8397.n101 a_71281_n8397.n92 4.64734
R48393 a_71281_n8397.n100 a_71281_n8397.n96 4.64734
R48394 a_71281_n8397.n115 a_71281_n8397.n106 4.64734
R48395 a_71281_n8397.n114 a_71281_n8397.n110 4.64734
R48396 a_71281_n8397.n287 a_71281_n8397.n283 4.64734
R48397 a_71281_n8397.n288 a_71281_n8397.n279 4.64734
R48398 a_71281_n8397.n273 a_71281_n8397.n269 4.64734
R48399 a_71281_n8397.n274 a_71281_n8397.n265 4.64734
R48400 a_71281_n8397.n259 a_71281_n8397.n255 4.64734
R48401 a_71281_n8397.n260 a_71281_n8397.n251 4.64734
R48402 a_71281_n8397.n245 a_71281_n8397.n241 4.64734
R48403 a_71281_n8397.n246 a_71281_n8397.n237 4.64734
R48404 a_71281_n8397.n228 a_71281_n8397.n224 4.64734
R48405 a_71281_n8397.n229 a_71281_n8397.n220 4.64734
R48406 a_71281_n8397.n214 a_71281_n8397.n210 4.64734
R48407 a_71281_n8397.n215 a_71281_n8397.n206 4.64734
R48408 a_71281_n8397.n197 a_71281_n8397.n193 4.64734
R48409 a_71281_n8397.n198 a_71281_n8397.n189 4.64734
R48410 a_71281_n8397.n183 a_71281_n8397.n179 4.64734
R48411 a_71281_n8397.n184 a_71281_n8397.n175 4.64734
R48412 a_71281_n8397.n419 a_71281_n8397.n415 4.64734
R48413 a_71281_n8397.n420 a_71281_n8397.n411 4.64734
R48414 a_71281_n8397.n433 a_71281_n8397.n429 4.64734
R48415 a_71281_n8397.n434 a_71281_n8397.n425 4.64734
R48416 a_71281_n8397.n461 a_71281_n8397.n452 4.64734
R48417 a_71281_n8397.n460 a_71281_n8397.n456 4.64734
R48418 a_71281_n8397.n447 a_71281_n8397.n439 4.64734
R48419 a_71281_n8397.n446 a_71281_n8397.n443 4.64734
R48420 a_71281_n8397.n302 a_71281_n8397.n294 4.64734
R48421 a_71281_n8397.n301 a_71281_n8397.n298 4.64734
R48422 a_71281_n8397.n316 a_71281_n8397.n307 4.64734
R48423 a_71281_n8397.n315 a_71281_n8397.n311 4.64734
R48424 a_71281_n8397.n330 a_71281_n8397.n321 4.64734
R48425 a_71281_n8397.n329 a_71281_n8397.n325 4.64734
R48426 a_71281_n8397.n344 a_71281_n8397.n335 4.64734
R48427 a_71281_n8397.n343 a_71281_n8397.n339 4.64734
R48428 a_71281_n8397.n361 a_71281_n8397.n352 4.64734
R48429 a_71281_n8397.n360 a_71281_n8397.n356 4.64734
R48430 a_71281_n8397.n375 a_71281_n8397.n366 4.64734
R48431 a_71281_n8397.n374 a_71281_n8397.n370 4.64734
R48432 a_71281_n8397.n392 a_71281_n8397.n383 4.64734
R48433 a_71281_n8397.n391 a_71281_n8397.n387 4.64734
R48434 a_71281_n8397.n406 a_71281_n8397.n397 4.64734
R48435 a_71281_n8397.n405 a_71281_n8397.n401 4.64734
R48436 a_71281_n8397.n578 a_71281_n8397.n574 4.64734
R48437 a_71281_n8397.n579 a_71281_n8397.n570 4.64734
R48438 a_71281_n8397.n564 a_71281_n8397.n560 4.64734
R48439 a_71281_n8397.n565 a_71281_n8397.n556 4.64734
R48440 a_71281_n8397.n550 a_71281_n8397.n546 4.64734
R48441 a_71281_n8397.n551 a_71281_n8397.n542 4.64734
R48442 a_71281_n8397.n536 a_71281_n8397.n532 4.64734
R48443 a_71281_n8397.n537 a_71281_n8397.n528 4.64734
R48444 a_71281_n8397.n519 a_71281_n8397.n515 4.64734
R48445 a_71281_n8397.n520 a_71281_n8397.n511 4.64734
R48446 a_71281_n8397.n505 a_71281_n8397.n501 4.64734
R48447 a_71281_n8397.n506 a_71281_n8397.n497 4.64734
R48448 a_71281_n8397.n488 a_71281_n8397.n484 4.64734
R48449 a_71281_n8397.n489 a_71281_n8397.n480 4.64734
R48450 a_71281_n8397.n474 a_71281_n8397.n470 4.64734
R48451 a_71281_n8397.n475 a_71281_n8397.n466 4.64734
R48452 a_71281_n8397.n741 a_71281_n8397.n732 4.64734
R48453 a_71281_n8397.n740 a_71281_n8397.n736 4.64734
R48454 a_71281_n8397.n755 a_71281_n8397.n746 4.64734
R48455 a_71281_n8397.n754 a_71281_n8397.n750 4.64734
R48456 a_71281_n8397.n769 a_71281_n8397.n760 4.64734
R48457 a_71281_n8397.n768 a_71281_n8397.n764 4.64734
R48458 a_71281_n8397.n783 a_71281_n8397.n774 4.64734
R48459 a_71281_n8397.n782 a_71281_n8397.n778 4.64734
R48460 a_71281_n8397.n868 a_71281_n8397.n864 4.64734
R48461 a_71281_n8397.n869 a_71281_n8397.n860 4.64734
R48462 a_71281_n8397.n854 a_71281_n8397.n850 4.64734
R48463 a_71281_n8397.n855 a_71281_n8397.n846 4.64734
R48464 a_71281_n8397.n837 a_71281_n8397.n833 4.64734
R48465 a_71281_n8397.n838 a_71281_n8397.n829 4.64734
R48466 a_71281_n8397.n823 a_71281_n8397.n819 4.64734
R48467 a_71281_n8397.n824 a_71281_n8397.n815 4.64734
R48468 a_71281_n8397.n642 a_71281_n8397.n641 4.01884
R48469 a_71281_n8397.n58 a_71281_n8397.n57 4.01884
R48470 a_71281_n8397.n234 a_71281_n8397.n233 4.01884
R48471 a_71281_n8397.n349 a_71281_n8397.n348 4.01884
R48472 a_71281_n8397.n525 a_71281_n8397.n524 4.01884
R48473 a_71281_n8397.n875 a_71281_n8397.n874 4.01884
R48474 a_71281_n8397.n673 a_71281_n8397.n672 4.00982
R48475 a_71281_n8397.n843 a_71281_n8397.n842 4.00982
R48476 a_71281_n8397.n89 a_71281_n8397.n88 4.00982
R48477 a_71281_n8397.n203 a_71281_n8397.n202 4.00982
R48478 a_71281_n8397.n380 a_71281_n8397.n379 4.00982
R48479 a_71281_n8397.n494 a_71281_n8397.n493 4.00982
R48480 a_71281_n8397.n584 a_71281_n8397.n292 3.61592
R48481 a_71281_n8397.n0 a_71281_n8397.n584 3.61491
R48482 a_71281_n8397.n714 a_71281_n8397.n713 2.25278
R48483 a_71281_n8397.n712 a_71281_n8397.n711 2.25278
R48484 a_71281_n8397.n728 a_71281_n8397.n727 2.25278
R48485 a_71281_n8397.n726 a_71281_n8397.n725 2.25278
R48486 a_71281_n8397.n809 a_71281_n8397.n808 2.25278
R48487 a_71281_n8397.n811 a_71281_n8397.n810 2.25278
R48488 a_71281_n8397.n795 a_71281_n8397.n794 2.25278
R48489 a_71281_n8397.n797 a_71281_n8397.n796 2.25278
R48490 a_71281_n8397.n594 a_71281_n8397.n593 2.25278
R48491 a_71281_n8397.n596 a_71281_n8397.n595 2.25278
R48492 a_71281_n8397.n608 a_71281_n8397.n607 2.25278
R48493 a_71281_n8397.n610 a_71281_n8397.n609 2.25278
R48494 a_71281_n8397.n622 a_71281_n8397.n621 2.25278
R48495 a_71281_n8397.n624 a_71281_n8397.n623 2.25278
R48496 a_71281_n8397.n636 a_71281_n8397.n635 2.25278
R48497 a_71281_n8397.n638 a_71281_n8397.n637 2.25278
R48498 a_71281_n8397.n653 a_71281_n8397.n652 2.25278
R48499 a_71281_n8397.n655 a_71281_n8397.n654 2.25278
R48500 a_71281_n8397.n667 a_71281_n8397.n666 2.25278
R48501 a_71281_n8397.n669 a_71281_n8397.n668 2.25278
R48502 a_71281_n8397.n684 a_71281_n8397.n683 2.25278
R48503 a_71281_n8397.n686 a_71281_n8397.n685 2.25278
R48504 a_71281_n8397.n698 a_71281_n8397.n697 2.25278
R48505 a_71281_n8397.n700 a_71281_n8397.n699 2.25278
R48506 a_71281_n8397.n130 a_71281_n8397.n129 2.25278
R48507 a_71281_n8397.n128 a_71281_n8397.n127 2.25278
R48508 a_71281_n8397.n144 a_71281_n8397.n143 2.25278
R48509 a_71281_n8397.n142 a_71281_n8397.n141 2.25278
R48510 a_71281_n8397.n169 a_71281_n8397.n168 2.25278
R48511 a_71281_n8397.n171 a_71281_n8397.n170 2.25278
R48512 a_71281_n8397.n155 a_71281_n8397.n154 2.25278
R48513 a_71281_n8397.n157 a_71281_n8397.n156 2.25278
R48514 a_71281_n8397.n10 a_71281_n8397.n9 2.25278
R48515 a_71281_n8397.n12 a_71281_n8397.n11 2.25278
R48516 a_71281_n8397.n24 a_71281_n8397.n23 2.25278
R48517 a_71281_n8397.n26 a_71281_n8397.n25 2.25278
R48518 a_71281_n8397.n38 a_71281_n8397.n37 2.25278
R48519 a_71281_n8397.n40 a_71281_n8397.n39 2.25278
R48520 a_71281_n8397.n52 a_71281_n8397.n51 2.25278
R48521 a_71281_n8397.n54 a_71281_n8397.n53 2.25278
R48522 a_71281_n8397.n69 a_71281_n8397.n68 2.25278
R48523 a_71281_n8397.n71 a_71281_n8397.n70 2.25278
R48524 a_71281_n8397.n83 a_71281_n8397.n82 2.25278
R48525 a_71281_n8397.n85 a_71281_n8397.n84 2.25278
R48526 a_71281_n8397.n100 a_71281_n8397.n99 2.25278
R48527 a_71281_n8397.n102 a_71281_n8397.n101 2.25278
R48528 a_71281_n8397.n114 a_71281_n8397.n113 2.25278
R48529 a_71281_n8397.n116 a_71281_n8397.n115 2.25278
R48530 a_71281_n8397.n289 a_71281_n8397.n288 2.25278
R48531 a_71281_n8397.n287 a_71281_n8397.n286 2.25278
R48532 a_71281_n8397.n275 a_71281_n8397.n274 2.25278
R48533 a_71281_n8397.n273 a_71281_n8397.n272 2.25278
R48534 a_71281_n8397.n261 a_71281_n8397.n260 2.25278
R48535 a_71281_n8397.n259 a_71281_n8397.n258 2.25278
R48536 a_71281_n8397.n247 a_71281_n8397.n246 2.25278
R48537 a_71281_n8397.n245 a_71281_n8397.n244 2.25278
R48538 a_71281_n8397.n230 a_71281_n8397.n229 2.25278
R48539 a_71281_n8397.n228 a_71281_n8397.n227 2.25278
R48540 a_71281_n8397.n216 a_71281_n8397.n215 2.25278
R48541 a_71281_n8397.n214 a_71281_n8397.n213 2.25278
R48542 a_71281_n8397.n199 a_71281_n8397.n198 2.25278
R48543 a_71281_n8397.n197 a_71281_n8397.n196 2.25278
R48544 a_71281_n8397.n185 a_71281_n8397.n184 2.25278
R48545 a_71281_n8397.n183 a_71281_n8397.n182 2.25278
R48546 a_71281_n8397.n421 a_71281_n8397.n420 2.25278
R48547 a_71281_n8397.n419 a_71281_n8397.n418 2.25278
R48548 a_71281_n8397.n435 a_71281_n8397.n434 2.25278
R48549 a_71281_n8397.n433 a_71281_n8397.n432 2.25278
R48550 a_71281_n8397.n460 a_71281_n8397.n459 2.25278
R48551 a_71281_n8397.n462 a_71281_n8397.n461 2.25278
R48552 a_71281_n8397.n446 a_71281_n8397.n445 2.25278
R48553 a_71281_n8397.n448 a_71281_n8397.n447 2.25278
R48554 a_71281_n8397.n301 a_71281_n8397.n300 2.25278
R48555 a_71281_n8397.n303 a_71281_n8397.n302 2.25278
R48556 a_71281_n8397.n315 a_71281_n8397.n314 2.25278
R48557 a_71281_n8397.n317 a_71281_n8397.n316 2.25278
R48558 a_71281_n8397.n329 a_71281_n8397.n328 2.25278
R48559 a_71281_n8397.n331 a_71281_n8397.n330 2.25278
R48560 a_71281_n8397.n343 a_71281_n8397.n342 2.25278
R48561 a_71281_n8397.n345 a_71281_n8397.n344 2.25278
R48562 a_71281_n8397.n360 a_71281_n8397.n359 2.25278
R48563 a_71281_n8397.n362 a_71281_n8397.n361 2.25278
R48564 a_71281_n8397.n374 a_71281_n8397.n373 2.25278
R48565 a_71281_n8397.n376 a_71281_n8397.n375 2.25278
R48566 a_71281_n8397.n391 a_71281_n8397.n390 2.25278
R48567 a_71281_n8397.n393 a_71281_n8397.n392 2.25278
R48568 a_71281_n8397.n405 a_71281_n8397.n404 2.25278
R48569 a_71281_n8397.n407 a_71281_n8397.n406 2.25278
R48570 a_71281_n8397.n580 a_71281_n8397.n579 2.25278
R48571 a_71281_n8397.n578 a_71281_n8397.n577 2.25278
R48572 a_71281_n8397.n566 a_71281_n8397.n565 2.25278
R48573 a_71281_n8397.n564 a_71281_n8397.n563 2.25278
R48574 a_71281_n8397.n552 a_71281_n8397.n551 2.25278
R48575 a_71281_n8397.n550 a_71281_n8397.n549 2.25278
R48576 a_71281_n8397.n538 a_71281_n8397.n537 2.25278
R48577 a_71281_n8397.n536 a_71281_n8397.n535 2.25278
R48578 a_71281_n8397.n521 a_71281_n8397.n520 2.25278
R48579 a_71281_n8397.n519 a_71281_n8397.n518 2.25278
R48580 a_71281_n8397.n507 a_71281_n8397.n506 2.25278
R48581 a_71281_n8397.n505 a_71281_n8397.n504 2.25278
R48582 a_71281_n8397.n490 a_71281_n8397.n489 2.25278
R48583 a_71281_n8397.n488 a_71281_n8397.n487 2.25278
R48584 a_71281_n8397.n476 a_71281_n8397.n475 2.25278
R48585 a_71281_n8397.n474 a_71281_n8397.n473 2.25278
R48586 a_71281_n8397.n740 a_71281_n8397.n739 2.25278
R48587 a_71281_n8397.n742 a_71281_n8397.n741 2.25278
R48588 a_71281_n8397.n754 a_71281_n8397.n753 2.25278
R48589 a_71281_n8397.n756 a_71281_n8397.n755 2.25278
R48590 a_71281_n8397.n768 a_71281_n8397.n767 2.25278
R48591 a_71281_n8397.n770 a_71281_n8397.n769 2.25278
R48592 a_71281_n8397.n782 a_71281_n8397.n781 2.25278
R48593 a_71281_n8397.n784 a_71281_n8397.n783 2.25278
R48594 a_71281_n8397.n870 a_71281_n8397.n869 2.25278
R48595 a_71281_n8397.n868 a_71281_n8397.n867 2.25278
R48596 a_71281_n8397.n856 a_71281_n8397.n855 2.25278
R48597 a_71281_n8397.n854 a_71281_n8397.n853 2.25278
R48598 a_71281_n8397.n839 a_71281_n8397.n838 2.25278
R48599 a_71281_n8397.n837 a_71281_n8397.n836 2.25278
R48600 a_71281_n8397.n825 a_71281_n8397.n824 2.25278
R48601 a_71281_n8397.n823 a_71281_n8397.n822 2.25278
R48602 a_71281_n8397.n1 a_71281_n8397.n0 0.0196917
R48603 a_71281_n8397.n14 a_71281_n8397.n2 1.6802
R48604 a_71281_n8397.n159 a_71281_n8397.n147 1.6802
R48605 a_71281_n8397.n305 a_71281_n8397.n293 1.6802
R48606 a_71281_n8397.n450 a_71281_n8397.n438 1.6802
R48607 a_71281_n8397.n598 a_71281_n8397.n586 1.6802
R48608 a_71281_n8397.n799 a_71281_n8397.n787 1.6802
R48609 a_71281_n8397.n180 a_71281_n8397.n174 1.5005
R48610 a_71281_n8397.n194 a_71281_n8397.n188 1.5005
R48611 a_71281_n8397.n211 a_71281_n8397.n205 1.5005
R48612 a_71281_n8397.n225 a_71281_n8397.n219 1.5005
R48613 a_71281_n8397.n235 a_71281_n8397.n234 1.5005
R48614 a_71281_n8397.n242 a_71281_n8397.n236 1.5005
R48615 a_71281_n8397.n256 a_71281_n8397.n250 1.5005
R48616 a_71281_n8397.n270 a_71281_n8397.n264 1.5005
R48617 a_71281_n8397.n284 a_71281_n8397.n278 1.5005
R48618 a_71281_n8397.n118 a_71281_n8397.n117 1.5005
R48619 a_71281_n8397.n104 a_71281_n8397.n103 1.5005
R48620 a_71281_n8397.n87 a_71281_n8397.n86 1.5005
R48621 a_71281_n8397.n73 a_71281_n8397.n72 1.5005
R48622 a_71281_n8397.n59 a_71281_n8397.n58 1.5005
R48623 a_71281_n8397.n56 a_71281_n8397.n55 1.5005
R48624 a_71281_n8397.n42 a_71281_n8397.n41 1.5005
R48625 a_71281_n8397.n28 a_71281_n8397.n27 1.5005
R48626 a_71281_n8397.n14 a_71281_n8397.n13 1.5005
R48627 a_71281_n8397.n204 a_71281_n8397.n203 1.5005
R48628 a_71281_n8397.n90 a_71281_n8397.n89 1.5005
R48629 a_71281_n8397.n159 a_71281_n8397.n158 1.5005
R48630 a_71281_n8397.n173 a_71281_n8397.n172 1.5005
R48631 a_71281_n8397.n167 a_71281_n8397.n160 1.5005
R48632 a_71281_n8397.n187 a_71281_n8397.n186 1.5005
R48633 a_71281_n8397.n201 a_71281_n8397.n200 1.5005
R48634 a_71281_n8397.n218 a_71281_n8397.n217 1.5005
R48635 a_71281_n8397.n232 a_71281_n8397.n231 1.5005
R48636 a_71281_n8397.n249 a_71281_n8397.n248 1.5005
R48637 a_71281_n8397.n263 a_71281_n8397.n262 1.5005
R48638 a_71281_n8397.n277 a_71281_n8397.n276 1.5005
R48639 a_71281_n8397.n291 a_71281_n8397.n290 1.5005
R48640 a_71281_n8397.n139 a_71281_n8397.n133 1.5005
R48641 a_71281_n8397.n146 a_71281_n8397.n145 1.5005
R48642 a_71281_n8397.n125 a_71281_n8397.n119 1.5005
R48643 a_71281_n8397.n132 a_71281_n8397.n131 1.5005
R48644 a_71281_n8397.n112 a_71281_n8397.n105 1.5005
R48645 a_71281_n8397.n98 a_71281_n8397.n91 1.5005
R48646 a_71281_n8397.n81 a_71281_n8397.n74 1.5005
R48647 a_71281_n8397.n67 a_71281_n8397.n60 1.5005
R48648 a_71281_n8397.n50 a_71281_n8397.n43 1.5005
R48649 a_71281_n8397.n36 a_71281_n8397.n29 1.5005
R48650 a_71281_n8397.n22 a_71281_n8397.n15 1.5005
R48651 a_71281_n8397.n471 a_71281_n8397.n465 1.5005
R48652 a_71281_n8397.n485 a_71281_n8397.n479 1.5005
R48653 a_71281_n8397.n502 a_71281_n8397.n496 1.5005
R48654 a_71281_n8397.n516 a_71281_n8397.n510 1.5005
R48655 a_71281_n8397.n526 a_71281_n8397.n525 1.5005
R48656 a_71281_n8397.n533 a_71281_n8397.n527 1.5005
R48657 a_71281_n8397.n547 a_71281_n8397.n541 1.5005
R48658 a_71281_n8397.n561 a_71281_n8397.n555 1.5005
R48659 a_71281_n8397.n575 a_71281_n8397.n569 1.5005
R48660 a_71281_n8397.n409 a_71281_n8397.n408 1.5005
R48661 a_71281_n8397.n395 a_71281_n8397.n394 1.5005
R48662 a_71281_n8397.n378 a_71281_n8397.n377 1.5005
R48663 a_71281_n8397.n364 a_71281_n8397.n363 1.5005
R48664 a_71281_n8397.n350 a_71281_n8397.n349 1.5005
R48665 a_71281_n8397.n347 a_71281_n8397.n346 1.5005
R48666 a_71281_n8397.n333 a_71281_n8397.n332 1.5005
R48667 a_71281_n8397.n319 a_71281_n8397.n318 1.5005
R48668 a_71281_n8397.n305 a_71281_n8397.n304 1.5005
R48669 a_71281_n8397.n495 a_71281_n8397.n494 1.5005
R48670 a_71281_n8397.n381 a_71281_n8397.n380 1.5005
R48671 a_71281_n8397.n450 a_71281_n8397.n449 1.5005
R48672 a_71281_n8397.n464 a_71281_n8397.n463 1.5005
R48673 a_71281_n8397.n458 a_71281_n8397.n451 1.5005
R48674 a_71281_n8397.n478 a_71281_n8397.n477 1.5005
R48675 a_71281_n8397.n492 a_71281_n8397.n491 1.5005
R48676 a_71281_n8397.n509 a_71281_n8397.n508 1.5005
R48677 a_71281_n8397.n523 a_71281_n8397.n522 1.5005
R48678 a_71281_n8397.n540 a_71281_n8397.n539 1.5005
R48679 a_71281_n8397.n554 a_71281_n8397.n553 1.5005
R48680 a_71281_n8397.n568 a_71281_n8397.n567 1.5005
R48681 a_71281_n8397.n582 a_71281_n8397.n581 1.5005
R48682 a_71281_n8397.n430 a_71281_n8397.n424 1.5005
R48683 a_71281_n8397.n437 a_71281_n8397.n436 1.5005
R48684 a_71281_n8397.n416 a_71281_n8397.n410 1.5005
R48685 a_71281_n8397.n423 a_71281_n8397.n422 1.5005
R48686 a_71281_n8397.n403 a_71281_n8397.n396 1.5005
R48687 a_71281_n8397.n389 a_71281_n8397.n382 1.5005
R48688 a_71281_n8397.n372 a_71281_n8397.n365 1.5005
R48689 a_71281_n8397.n358 a_71281_n8397.n351 1.5005
R48690 a_71281_n8397.n341 a_71281_n8397.n334 1.5005
R48691 a_71281_n8397.n327 a_71281_n8397.n320 1.5005
R48692 a_71281_n8397.n313 a_71281_n8397.n306 1.5005
R48693 a_71281_n8397.n820 a_71281_n8397.n814 1.5005
R48694 a_71281_n8397.n834 a_71281_n8397.n828 1.5005
R48695 a_71281_n8397.n851 a_71281_n8397.n845 1.5005
R48696 a_71281_n8397.n865 a_71281_n8397.n859 1.5005
R48697 a_71281_n8397.n786 a_71281_n8397.n785 1.5005
R48698 a_71281_n8397.n772 a_71281_n8397.n771 1.5005
R48699 a_71281_n8397.n758 a_71281_n8397.n757 1.5005
R48700 a_71281_n8397.n744 a_71281_n8397.n743 1.5005
R48701 a_71281_n8397.n702 a_71281_n8397.n701 1.5005
R48702 a_71281_n8397.n688 a_71281_n8397.n687 1.5005
R48703 a_71281_n8397.n671 a_71281_n8397.n670 1.5005
R48704 a_71281_n8397.n657 a_71281_n8397.n656 1.5005
R48705 a_71281_n8397.n643 a_71281_n8397.n642 1.5005
R48706 a_71281_n8397.n640 a_71281_n8397.n639 1.5005
R48707 a_71281_n8397.n626 a_71281_n8397.n625 1.5005
R48708 a_71281_n8397.n612 a_71281_n8397.n611 1.5005
R48709 a_71281_n8397.n598 a_71281_n8397.n597 1.5005
R48710 a_71281_n8397.n844 a_71281_n8397.n843 1.5005
R48711 a_71281_n8397.n674 a_71281_n8397.n673 1.5005
R48712 a_71281_n8397.n799 a_71281_n8397.n798 1.5005
R48713 a_71281_n8397.n813 a_71281_n8397.n812 1.5005
R48714 a_71281_n8397.n807 a_71281_n8397.n800 1.5005
R48715 a_71281_n8397.n827 a_71281_n8397.n826 1.5005
R48716 a_71281_n8397.n841 a_71281_n8397.n840 1.5005
R48717 a_71281_n8397.n858 a_71281_n8397.n857 1.5005
R48718 a_71281_n8397.n872 a_71281_n8397.n871 1.5005
R48719 a_71281_n8397.n780 a_71281_n8397.n773 1.5005
R48720 a_71281_n8397.n766 a_71281_n8397.n759 1.5005
R48721 a_71281_n8397.n752 a_71281_n8397.n745 1.5005
R48722 a_71281_n8397.n738 a_71281_n8397.n731 1.5005
R48723 a_71281_n8397.n723 a_71281_n8397.n717 1.5005
R48724 a_71281_n8397.n730 a_71281_n8397.n729 1.5005
R48725 a_71281_n8397.n709 a_71281_n8397.n703 1.5005
R48726 a_71281_n8397.n716 a_71281_n8397.n715 1.5005
R48727 a_71281_n8397.n696 a_71281_n8397.n689 1.5005
R48728 a_71281_n8397.n682 a_71281_n8397.n675 1.5005
R48729 a_71281_n8397.n665 a_71281_n8397.n658 1.5005
R48730 a_71281_n8397.n651 a_71281_n8397.n644 1.5005
R48731 a_71281_n8397.n634 a_71281_n8397.n627 1.5005
R48732 a_71281_n8397.n620 a_71281_n8397.n613 1.5005
R48733 a_71281_n8397.n606 a_71281_n8397.n599 1.5005
R48734 a_71281_n8397.n874 a_71281_n8397.n873 1.5005
R48735 a_71281_n8397.n672 a_71281_n8397.t33 1.4705
R48736 a_71281_n8397.n672 a_71281_n8397.t29 1.4705
R48737 a_71281_n8397.n842 a_71281_n8397.t23 1.4705
R48738 a_71281_n8397.n842 a_71281_n8397.t53 1.4705
R48739 a_71281_n8397.n641 a_71281_n8397.t57 1.4705
R48740 a_71281_n8397.n641 a_71281_n8397.t35 1.4705
R48741 a_71281_n8397.n88 a_71281_n8397.t47 1.4705
R48742 a_71281_n8397.n88 a_71281_n8397.t21 1.4705
R48743 a_71281_n8397.n202 a_71281_n8397.t65 1.4705
R48744 a_71281_n8397.n202 a_71281_n8397.t13 1.4705
R48745 a_71281_n8397.n57 a_71281_n8397.t43 1.4705
R48746 a_71281_n8397.n57 a_71281_n8397.t11 1.4705
R48747 a_71281_n8397.n233 a_71281_n8397.t31 1.4705
R48748 a_71281_n8397.n233 a_71281_n8397.t39 1.4705
R48749 a_71281_n8397.n379 a_71281_n8397.t59 1.4705
R48750 a_71281_n8397.n379 a_71281_n8397.t27 1.4705
R48751 a_71281_n8397.n493 a_71281_n8397.t37 1.4705
R48752 a_71281_n8397.n493 a_71281_n8397.t49 1.4705
R48753 a_71281_n8397.n348 a_71281_n8397.t55 1.4705
R48754 a_71281_n8397.n348 a_71281_n8397.t25 1.4705
R48755 a_71281_n8397.n524 a_71281_n8397.t69 1.4705
R48756 a_71281_n8397.n524 a_71281_n8397.t71 1.4705
R48757 a_71281_n8397.t73 a_71281_n8397.n875 1.4705
R48758 a_71281_n8397.n875 a_71281_n8397.t41 1.4705
R48759 a_71281_n8397.n584 a_71281_n8397.n583 0.7505
R48760 a_71281_n8397.n714 a_71281_n8397.n705 0.567403
R48761 a_71281_n8397.n711 a_71281_n8397.n710 0.567403
R48762 a_71281_n8397.n728 a_71281_n8397.n719 0.567403
R48763 a_71281_n8397.n725 a_71281_n8397.n724 0.567403
R48764 a_71281_n8397.n808 a_71281_n8397.n806 0.567403
R48765 a_71281_n8397.n811 a_71281_n8397.n802 0.567403
R48766 a_71281_n8397.n794 a_71281_n8397.n793 0.567403
R48767 a_71281_n8397.n797 a_71281_n8397.n789 0.567403
R48768 a_71281_n8397.n593 a_71281_n8397.n592 0.567403
R48769 a_71281_n8397.n596 a_71281_n8397.n588 0.567403
R48770 a_71281_n8397.n607 a_71281_n8397.n605 0.567403
R48771 a_71281_n8397.n610 a_71281_n8397.n601 0.567403
R48772 a_71281_n8397.n621 a_71281_n8397.n619 0.567403
R48773 a_71281_n8397.n624 a_71281_n8397.n615 0.567403
R48774 a_71281_n8397.n635 a_71281_n8397.n633 0.567403
R48775 a_71281_n8397.n638 a_71281_n8397.n629 0.567403
R48776 a_71281_n8397.n652 a_71281_n8397.n650 0.567403
R48777 a_71281_n8397.n655 a_71281_n8397.n646 0.567403
R48778 a_71281_n8397.n666 a_71281_n8397.n664 0.567403
R48779 a_71281_n8397.n669 a_71281_n8397.n660 0.567403
R48780 a_71281_n8397.n683 a_71281_n8397.n681 0.567403
R48781 a_71281_n8397.n686 a_71281_n8397.n677 0.567403
R48782 a_71281_n8397.n697 a_71281_n8397.n695 0.567403
R48783 a_71281_n8397.n700 a_71281_n8397.n691 0.567403
R48784 a_71281_n8397.n130 a_71281_n8397.n121 0.567403
R48785 a_71281_n8397.n127 a_71281_n8397.n126 0.567403
R48786 a_71281_n8397.n144 a_71281_n8397.n135 0.567403
R48787 a_71281_n8397.n141 a_71281_n8397.n140 0.567403
R48788 a_71281_n8397.n168 a_71281_n8397.n166 0.567403
R48789 a_71281_n8397.n171 a_71281_n8397.n162 0.567403
R48790 a_71281_n8397.n154 a_71281_n8397.n153 0.567403
R48791 a_71281_n8397.n157 a_71281_n8397.n149 0.567403
R48792 a_71281_n8397.n9 a_71281_n8397.n8 0.567403
R48793 a_71281_n8397.n12 a_71281_n8397.n4 0.567403
R48794 a_71281_n8397.n23 a_71281_n8397.n21 0.567403
R48795 a_71281_n8397.n26 a_71281_n8397.n17 0.567403
R48796 a_71281_n8397.n37 a_71281_n8397.n35 0.567403
R48797 a_71281_n8397.n40 a_71281_n8397.n31 0.567403
R48798 a_71281_n8397.n51 a_71281_n8397.n49 0.567403
R48799 a_71281_n8397.n54 a_71281_n8397.n45 0.567403
R48800 a_71281_n8397.n68 a_71281_n8397.n66 0.567403
R48801 a_71281_n8397.n71 a_71281_n8397.n62 0.567403
R48802 a_71281_n8397.n82 a_71281_n8397.n80 0.567403
R48803 a_71281_n8397.n85 a_71281_n8397.n76 0.567403
R48804 a_71281_n8397.n99 a_71281_n8397.n97 0.567403
R48805 a_71281_n8397.n102 a_71281_n8397.n93 0.567403
R48806 a_71281_n8397.n113 a_71281_n8397.n111 0.567403
R48807 a_71281_n8397.n116 a_71281_n8397.n107 0.567403
R48808 a_71281_n8397.n289 a_71281_n8397.n280 0.567403
R48809 a_71281_n8397.n286 a_71281_n8397.n285 0.567403
R48810 a_71281_n8397.n275 a_71281_n8397.n266 0.567403
R48811 a_71281_n8397.n272 a_71281_n8397.n271 0.567403
R48812 a_71281_n8397.n261 a_71281_n8397.n252 0.567403
R48813 a_71281_n8397.n258 a_71281_n8397.n257 0.567403
R48814 a_71281_n8397.n247 a_71281_n8397.n238 0.567403
R48815 a_71281_n8397.n244 a_71281_n8397.n243 0.567403
R48816 a_71281_n8397.n230 a_71281_n8397.n221 0.567403
R48817 a_71281_n8397.n227 a_71281_n8397.n226 0.567403
R48818 a_71281_n8397.n216 a_71281_n8397.n207 0.567403
R48819 a_71281_n8397.n213 a_71281_n8397.n212 0.567403
R48820 a_71281_n8397.n199 a_71281_n8397.n190 0.567403
R48821 a_71281_n8397.n196 a_71281_n8397.n195 0.567403
R48822 a_71281_n8397.n185 a_71281_n8397.n176 0.567403
R48823 a_71281_n8397.n182 a_71281_n8397.n181 0.567403
R48824 a_71281_n8397.n421 a_71281_n8397.n412 0.567403
R48825 a_71281_n8397.n418 a_71281_n8397.n417 0.567403
R48826 a_71281_n8397.n435 a_71281_n8397.n426 0.567403
R48827 a_71281_n8397.n432 a_71281_n8397.n431 0.567403
R48828 a_71281_n8397.n459 a_71281_n8397.n457 0.567403
R48829 a_71281_n8397.n462 a_71281_n8397.n453 0.567403
R48830 a_71281_n8397.n445 a_71281_n8397.n444 0.567403
R48831 a_71281_n8397.n448 a_71281_n8397.n440 0.567403
R48832 a_71281_n8397.n300 a_71281_n8397.n299 0.567403
R48833 a_71281_n8397.n303 a_71281_n8397.n295 0.567403
R48834 a_71281_n8397.n314 a_71281_n8397.n312 0.567403
R48835 a_71281_n8397.n317 a_71281_n8397.n308 0.567403
R48836 a_71281_n8397.n328 a_71281_n8397.n326 0.567403
R48837 a_71281_n8397.n331 a_71281_n8397.n322 0.567403
R48838 a_71281_n8397.n342 a_71281_n8397.n340 0.567403
R48839 a_71281_n8397.n345 a_71281_n8397.n336 0.567403
R48840 a_71281_n8397.n359 a_71281_n8397.n357 0.567403
R48841 a_71281_n8397.n362 a_71281_n8397.n353 0.567403
R48842 a_71281_n8397.n373 a_71281_n8397.n371 0.567403
R48843 a_71281_n8397.n376 a_71281_n8397.n367 0.567403
R48844 a_71281_n8397.n390 a_71281_n8397.n388 0.567403
R48845 a_71281_n8397.n393 a_71281_n8397.n384 0.567403
R48846 a_71281_n8397.n404 a_71281_n8397.n402 0.567403
R48847 a_71281_n8397.n407 a_71281_n8397.n398 0.567403
R48848 a_71281_n8397.n580 a_71281_n8397.n571 0.567403
R48849 a_71281_n8397.n577 a_71281_n8397.n576 0.567403
R48850 a_71281_n8397.n566 a_71281_n8397.n557 0.567403
R48851 a_71281_n8397.n563 a_71281_n8397.n562 0.567403
R48852 a_71281_n8397.n552 a_71281_n8397.n543 0.567403
R48853 a_71281_n8397.n549 a_71281_n8397.n548 0.567403
R48854 a_71281_n8397.n538 a_71281_n8397.n529 0.567403
R48855 a_71281_n8397.n535 a_71281_n8397.n534 0.567403
R48856 a_71281_n8397.n521 a_71281_n8397.n512 0.567403
R48857 a_71281_n8397.n518 a_71281_n8397.n517 0.567403
R48858 a_71281_n8397.n507 a_71281_n8397.n498 0.567403
R48859 a_71281_n8397.n504 a_71281_n8397.n503 0.567403
R48860 a_71281_n8397.n490 a_71281_n8397.n481 0.567403
R48861 a_71281_n8397.n487 a_71281_n8397.n486 0.567403
R48862 a_71281_n8397.n476 a_71281_n8397.n467 0.567403
R48863 a_71281_n8397.n473 a_71281_n8397.n472 0.567403
R48864 a_71281_n8397.n739 a_71281_n8397.n737 0.567403
R48865 a_71281_n8397.n742 a_71281_n8397.n733 0.567403
R48866 a_71281_n8397.n753 a_71281_n8397.n751 0.567403
R48867 a_71281_n8397.n756 a_71281_n8397.n747 0.567403
R48868 a_71281_n8397.n767 a_71281_n8397.n765 0.567403
R48869 a_71281_n8397.n770 a_71281_n8397.n761 0.567403
R48870 a_71281_n8397.n781 a_71281_n8397.n779 0.567403
R48871 a_71281_n8397.n784 a_71281_n8397.n775 0.567403
R48872 a_71281_n8397.n870 a_71281_n8397.n861 0.567403
R48873 a_71281_n8397.n867 a_71281_n8397.n866 0.567403
R48874 a_71281_n8397.n856 a_71281_n8397.n847 0.567403
R48875 a_71281_n8397.n853 a_71281_n8397.n852 0.567403
R48876 a_71281_n8397.n839 a_71281_n8397.n830 0.567403
R48877 a_71281_n8397.n836 a_71281_n8397.n835 0.567403
R48878 a_71281_n8397.n825 a_71281_n8397.n816 0.567403
R48879 a_71281_n8397.n822 a_71281_n8397.n821 0.567403
R48880 a_71281_n8397.n706 a_71281_n8397.n704 0.496742
R48881 a_71281_n8397.n708 a_71281_n8397.n707 0.496742
R48882 a_71281_n8397.n720 a_71281_n8397.n718 0.496742
R48883 a_71281_n8397.n722 a_71281_n8397.n721 0.496742
R48884 a_71281_n8397.n805 a_71281_n8397.n804 0.496742
R48885 a_71281_n8397.n803 a_71281_n8397.n801 0.496742
R48886 a_71281_n8397.n792 a_71281_n8397.n791 0.496742
R48887 a_71281_n8397.n790 a_71281_n8397.n788 0.496742
R48888 a_71281_n8397.n591 a_71281_n8397.n590 0.496742
R48889 a_71281_n8397.n589 a_71281_n8397.n587 0.496742
R48890 a_71281_n8397.n604 a_71281_n8397.n603 0.496742
R48891 a_71281_n8397.n602 a_71281_n8397.n600 0.496742
R48892 a_71281_n8397.n618 a_71281_n8397.n617 0.496742
R48893 a_71281_n8397.n616 a_71281_n8397.n614 0.496742
R48894 a_71281_n8397.n632 a_71281_n8397.n631 0.496742
R48895 a_71281_n8397.n630 a_71281_n8397.n628 0.496742
R48896 a_71281_n8397.n649 a_71281_n8397.n648 0.496742
R48897 a_71281_n8397.n647 a_71281_n8397.n645 0.496742
R48898 a_71281_n8397.n663 a_71281_n8397.n662 0.496742
R48899 a_71281_n8397.n661 a_71281_n8397.n659 0.496742
R48900 a_71281_n8397.n680 a_71281_n8397.n679 0.496742
R48901 a_71281_n8397.n678 a_71281_n8397.n676 0.496742
R48902 a_71281_n8397.n694 a_71281_n8397.n693 0.496742
R48903 a_71281_n8397.n692 a_71281_n8397.n690 0.496742
R48904 a_71281_n8397.n122 a_71281_n8397.n120 0.496742
R48905 a_71281_n8397.n124 a_71281_n8397.n123 0.496742
R48906 a_71281_n8397.n136 a_71281_n8397.n134 0.496742
R48907 a_71281_n8397.n138 a_71281_n8397.n137 0.496742
R48908 a_71281_n8397.n165 a_71281_n8397.n164 0.496742
R48909 a_71281_n8397.n163 a_71281_n8397.n161 0.496742
R48910 a_71281_n8397.n152 a_71281_n8397.n151 0.496742
R48911 a_71281_n8397.n150 a_71281_n8397.n148 0.496742
R48912 a_71281_n8397.n7 a_71281_n8397.n6 0.496742
R48913 a_71281_n8397.n5 a_71281_n8397.n3 0.496742
R48914 a_71281_n8397.n20 a_71281_n8397.n19 0.496742
R48915 a_71281_n8397.n18 a_71281_n8397.n16 0.496742
R48916 a_71281_n8397.n34 a_71281_n8397.n33 0.496742
R48917 a_71281_n8397.n32 a_71281_n8397.n30 0.496742
R48918 a_71281_n8397.n48 a_71281_n8397.n47 0.496742
R48919 a_71281_n8397.n46 a_71281_n8397.n44 0.496742
R48920 a_71281_n8397.n65 a_71281_n8397.n64 0.496742
R48921 a_71281_n8397.n63 a_71281_n8397.n61 0.496742
R48922 a_71281_n8397.n79 a_71281_n8397.n78 0.496742
R48923 a_71281_n8397.n77 a_71281_n8397.n75 0.496742
R48924 a_71281_n8397.n96 a_71281_n8397.n95 0.496742
R48925 a_71281_n8397.n94 a_71281_n8397.n92 0.496742
R48926 a_71281_n8397.n110 a_71281_n8397.n109 0.496742
R48927 a_71281_n8397.n108 a_71281_n8397.n106 0.496742
R48928 a_71281_n8397.n281 a_71281_n8397.n279 0.496742
R48929 a_71281_n8397.n283 a_71281_n8397.n282 0.496742
R48930 a_71281_n8397.n267 a_71281_n8397.n265 0.496742
R48931 a_71281_n8397.n269 a_71281_n8397.n268 0.496742
R48932 a_71281_n8397.n253 a_71281_n8397.n251 0.496742
R48933 a_71281_n8397.n255 a_71281_n8397.n254 0.496742
R48934 a_71281_n8397.n239 a_71281_n8397.n237 0.496742
R48935 a_71281_n8397.n241 a_71281_n8397.n240 0.496742
R48936 a_71281_n8397.n222 a_71281_n8397.n220 0.496742
R48937 a_71281_n8397.n224 a_71281_n8397.n223 0.496742
R48938 a_71281_n8397.n208 a_71281_n8397.n206 0.496742
R48939 a_71281_n8397.n210 a_71281_n8397.n209 0.496742
R48940 a_71281_n8397.n191 a_71281_n8397.n189 0.496742
R48941 a_71281_n8397.n193 a_71281_n8397.n192 0.496742
R48942 a_71281_n8397.n177 a_71281_n8397.n175 0.496742
R48943 a_71281_n8397.n179 a_71281_n8397.n178 0.496742
R48944 a_71281_n8397.n413 a_71281_n8397.n411 0.496742
R48945 a_71281_n8397.n415 a_71281_n8397.n414 0.496742
R48946 a_71281_n8397.n427 a_71281_n8397.n425 0.496742
R48947 a_71281_n8397.n429 a_71281_n8397.n428 0.496742
R48948 a_71281_n8397.n456 a_71281_n8397.n455 0.496742
R48949 a_71281_n8397.n454 a_71281_n8397.n452 0.496742
R48950 a_71281_n8397.n443 a_71281_n8397.n442 0.496742
R48951 a_71281_n8397.n441 a_71281_n8397.n439 0.496742
R48952 a_71281_n8397.n298 a_71281_n8397.n297 0.496742
R48953 a_71281_n8397.n296 a_71281_n8397.n294 0.496742
R48954 a_71281_n8397.n311 a_71281_n8397.n310 0.496742
R48955 a_71281_n8397.n309 a_71281_n8397.n307 0.496742
R48956 a_71281_n8397.n325 a_71281_n8397.n324 0.496742
R48957 a_71281_n8397.n323 a_71281_n8397.n321 0.496742
R48958 a_71281_n8397.n339 a_71281_n8397.n338 0.496742
R48959 a_71281_n8397.n337 a_71281_n8397.n335 0.496742
R48960 a_71281_n8397.n356 a_71281_n8397.n355 0.496742
R48961 a_71281_n8397.n354 a_71281_n8397.n352 0.496742
R48962 a_71281_n8397.n370 a_71281_n8397.n369 0.496742
R48963 a_71281_n8397.n368 a_71281_n8397.n366 0.496742
R48964 a_71281_n8397.n387 a_71281_n8397.n386 0.496742
R48965 a_71281_n8397.n385 a_71281_n8397.n383 0.496742
R48966 a_71281_n8397.n401 a_71281_n8397.n400 0.496742
R48967 a_71281_n8397.n399 a_71281_n8397.n397 0.496742
R48968 a_71281_n8397.n572 a_71281_n8397.n570 0.496742
R48969 a_71281_n8397.n574 a_71281_n8397.n573 0.496742
R48970 a_71281_n8397.n558 a_71281_n8397.n556 0.496742
R48971 a_71281_n8397.n560 a_71281_n8397.n559 0.496742
R48972 a_71281_n8397.n544 a_71281_n8397.n542 0.496742
R48973 a_71281_n8397.n546 a_71281_n8397.n545 0.496742
R48974 a_71281_n8397.n530 a_71281_n8397.n528 0.496742
R48975 a_71281_n8397.n532 a_71281_n8397.n531 0.496742
R48976 a_71281_n8397.n513 a_71281_n8397.n511 0.496742
R48977 a_71281_n8397.n515 a_71281_n8397.n514 0.496742
R48978 a_71281_n8397.n499 a_71281_n8397.n497 0.496742
R48979 a_71281_n8397.n501 a_71281_n8397.n500 0.496742
R48980 a_71281_n8397.n482 a_71281_n8397.n480 0.496742
R48981 a_71281_n8397.n484 a_71281_n8397.n483 0.496742
R48982 a_71281_n8397.n468 a_71281_n8397.n466 0.496742
R48983 a_71281_n8397.n470 a_71281_n8397.n469 0.496742
R48984 a_71281_n8397.n736 a_71281_n8397.n735 0.496742
R48985 a_71281_n8397.n734 a_71281_n8397.n732 0.496742
R48986 a_71281_n8397.n750 a_71281_n8397.n749 0.496742
R48987 a_71281_n8397.n748 a_71281_n8397.n746 0.496742
R48988 a_71281_n8397.n764 a_71281_n8397.n763 0.496742
R48989 a_71281_n8397.n762 a_71281_n8397.n760 0.496742
R48990 a_71281_n8397.n778 a_71281_n8397.n777 0.496742
R48991 a_71281_n8397.n776 a_71281_n8397.n774 0.496742
R48992 a_71281_n8397.n862 a_71281_n8397.n860 0.496742
R48993 a_71281_n8397.n864 a_71281_n8397.n863 0.496742
R48994 a_71281_n8397.n848 a_71281_n8397.n846 0.496742
R48995 a_71281_n8397.n850 a_71281_n8397.n849 0.496742
R48996 a_71281_n8397.n831 a_71281_n8397.n829 0.496742
R48997 a_71281_n8397.n833 a_71281_n8397.n832 0.496742
R48998 a_71281_n8397.n817 a_71281_n8397.n815 0.496742
R48999 a_71281_n8397.n819 a_71281_n8397.n818 0.496742
R49000 a_71281_n8397.n292 a_71281_n8397.n291 0.445939
R49001 a_71281_n8397.n583 a_71281_n8397.n582 0.445939
R49002 a_71281_n8397.n292 a_71281_n8397.n146 0.443507
R49003 a_71281_n8397.n583 a_71281_n8397.n437 0.443507
R49004 a_71281_n8397.n0 a_71281_n8397.n730 0.427392
R49005 a_71281_n8397.n56 a_71281_n8397.n43 0.180804
R49006 a_71281_n8397.n132 a_71281_n8397.n119 0.180804
R49007 a_71281_n8397.n249 a_71281_n8397.n236 0.180804
R49008 a_71281_n8397.n173 a_71281_n8397.n160 0.180804
R49009 a_71281_n8397.n347 a_71281_n8397.n334 0.180804
R49010 a_71281_n8397.n423 a_71281_n8397.n410 0.180804
R49011 a_71281_n8397.n540 a_71281_n8397.n527 0.180804
R49012 a_71281_n8397.n464 a_71281_n8397.n451 0.180804
R49013 a_71281_n8397.n640 a_71281_n8397.n627 0.180804
R49014 a_71281_n8397.n716 a_71281_n8397.n703 0.180804
R49015 a_71281_n8397.n786 a_71281_n8397.n773 0.180804
R49016 a_71281_n8397.n813 a_71281_n8397.n800 0.180804
R49017 a_71281_n8397.n42 a_71281_n8397.n29 0.180196
R49018 a_71281_n8397.n73 a_71281_n8397.n60 0.180196
R49019 a_71281_n8397.n87 a_71281_n8397.n74 0.180196
R49020 a_71281_n8397.n118 a_71281_n8397.n105 0.180196
R49021 a_71281_n8397.n146 a_71281_n8397.n133 0.180196
R49022 a_71281_n8397.n291 a_71281_n8397.n278 0.180196
R49023 a_71281_n8397.n263 a_71281_n8397.n250 0.180196
R49024 a_71281_n8397.n232 a_71281_n8397.n219 0.180196
R49025 a_71281_n8397.n218 a_71281_n8397.n205 0.180196
R49026 a_71281_n8397.n187 a_71281_n8397.n174 0.180196
R49027 a_71281_n8397.n333 a_71281_n8397.n320 0.180196
R49028 a_71281_n8397.n364 a_71281_n8397.n351 0.180196
R49029 a_71281_n8397.n378 a_71281_n8397.n365 0.180196
R49030 a_71281_n8397.n409 a_71281_n8397.n396 0.180196
R49031 a_71281_n8397.n437 a_71281_n8397.n424 0.180196
R49032 a_71281_n8397.n582 a_71281_n8397.n569 0.180196
R49033 a_71281_n8397.n554 a_71281_n8397.n541 0.180196
R49034 a_71281_n8397.n523 a_71281_n8397.n510 0.180196
R49035 a_71281_n8397.n509 a_71281_n8397.n496 0.180196
R49036 a_71281_n8397.n478 a_71281_n8397.n465 0.180196
R49037 a_71281_n8397.n626 a_71281_n8397.n613 0.180196
R49038 a_71281_n8397.n657 a_71281_n8397.n644 0.180196
R49039 a_71281_n8397.n671 a_71281_n8397.n658 0.180196
R49040 a_71281_n8397.n702 a_71281_n8397.n689 0.180196
R49041 a_71281_n8397.n730 a_71281_n8397.n717 0.180196
R49042 a_71281_n8397.n744 a_71281_n8397.n731 0.180196
R49043 a_71281_n8397.n772 a_71281_n8397.n759 0.180196
R49044 a_71281_n8397.n872 a_71281_n8397.n859 0.180196
R49045 a_71281_n8397.n858 a_71281_n8397.n845 0.180196
R49046 a_71281_n8397.n827 a_71281_n8397.n814 0.180196
R49047 a_71281_n8397.n28 a_71281_n8397.n15 0.179892
R49048 a_71281_n8397.n104 a_71281_n8397.n91 0.179892
R49049 a_71281_n8397.n277 a_71281_n8397.n264 0.179892
R49050 a_71281_n8397.n201 a_71281_n8397.n188 0.179892
R49051 a_71281_n8397.n319 a_71281_n8397.n306 0.179892
R49052 a_71281_n8397.n395 a_71281_n8397.n382 0.179892
R49053 a_71281_n8397.n568 a_71281_n8397.n555 0.179892
R49054 a_71281_n8397.n492 a_71281_n8397.n479 0.179892
R49055 a_71281_n8397.n612 a_71281_n8397.n599 0.179892
R49056 a_71281_n8397.n688 a_71281_n8397.n675 0.179892
R49057 a_71281_n8397.n758 a_71281_n8397.n745 0.179892
R49058 a_71281_n8397.n841 a_71281_n8397.n828 0.179892
R49059 a_71281_n8397.n715 a_71281_n8397.n704 0.136625
R49060 a_71281_n8397.n709 a_71281_n8397.n708 0.136625
R49061 a_71281_n8397.n729 a_71281_n8397.n718 0.136625
R49062 a_71281_n8397.n723 a_71281_n8397.n722 0.136625
R49063 a_71281_n8397.n807 a_71281_n8397.n805 0.136625
R49064 a_71281_n8397.n812 a_71281_n8397.n801 0.136625
R49065 a_71281_n8397.n792 a_71281_n8397.n787 0.136625
R49066 a_71281_n8397.n798 a_71281_n8397.n788 0.136625
R49067 a_71281_n8397.n591 a_71281_n8397.n586 0.136625
R49068 a_71281_n8397.n597 a_71281_n8397.n587 0.136625
R49069 a_71281_n8397.n606 a_71281_n8397.n604 0.136625
R49070 a_71281_n8397.n611 a_71281_n8397.n600 0.136625
R49071 a_71281_n8397.n620 a_71281_n8397.n618 0.136625
R49072 a_71281_n8397.n625 a_71281_n8397.n614 0.136625
R49073 a_71281_n8397.n634 a_71281_n8397.n632 0.136625
R49074 a_71281_n8397.n639 a_71281_n8397.n628 0.136625
R49075 a_71281_n8397.n651 a_71281_n8397.n649 0.136625
R49076 a_71281_n8397.n656 a_71281_n8397.n645 0.136625
R49077 a_71281_n8397.n665 a_71281_n8397.n663 0.136625
R49078 a_71281_n8397.n670 a_71281_n8397.n659 0.136625
R49079 a_71281_n8397.n682 a_71281_n8397.n680 0.136625
R49080 a_71281_n8397.n687 a_71281_n8397.n676 0.136625
R49081 a_71281_n8397.n696 a_71281_n8397.n694 0.136625
R49082 a_71281_n8397.n701 a_71281_n8397.n690 0.136625
R49083 a_71281_n8397.n131 a_71281_n8397.n120 0.136625
R49084 a_71281_n8397.n125 a_71281_n8397.n124 0.136625
R49085 a_71281_n8397.n145 a_71281_n8397.n134 0.136625
R49086 a_71281_n8397.n139 a_71281_n8397.n138 0.136625
R49087 a_71281_n8397.n167 a_71281_n8397.n165 0.136625
R49088 a_71281_n8397.n172 a_71281_n8397.n161 0.136625
R49089 a_71281_n8397.n152 a_71281_n8397.n147 0.136625
R49090 a_71281_n8397.n158 a_71281_n8397.n148 0.136625
R49091 a_71281_n8397.n7 a_71281_n8397.n2 0.136625
R49092 a_71281_n8397.n13 a_71281_n8397.n3 0.136625
R49093 a_71281_n8397.n22 a_71281_n8397.n20 0.136625
R49094 a_71281_n8397.n27 a_71281_n8397.n16 0.136625
R49095 a_71281_n8397.n36 a_71281_n8397.n34 0.136625
R49096 a_71281_n8397.n41 a_71281_n8397.n30 0.136625
R49097 a_71281_n8397.n50 a_71281_n8397.n48 0.136625
R49098 a_71281_n8397.n55 a_71281_n8397.n44 0.136625
R49099 a_71281_n8397.n67 a_71281_n8397.n65 0.136625
R49100 a_71281_n8397.n72 a_71281_n8397.n61 0.136625
R49101 a_71281_n8397.n81 a_71281_n8397.n79 0.136625
R49102 a_71281_n8397.n86 a_71281_n8397.n75 0.136625
R49103 a_71281_n8397.n98 a_71281_n8397.n96 0.136625
R49104 a_71281_n8397.n103 a_71281_n8397.n92 0.136625
R49105 a_71281_n8397.n112 a_71281_n8397.n110 0.136625
R49106 a_71281_n8397.n117 a_71281_n8397.n106 0.136625
R49107 a_71281_n8397.n290 a_71281_n8397.n279 0.136625
R49108 a_71281_n8397.n284 a_71281_n8397.n283 0.136625
R49109 a_71281_n8397.n276 a_71281_n8397.n265 0.136625
R49110 a_71281_n8397.n270 a_71281_n8397.n269 0.136625
R49111 a_71281_n8397.n262 a_71281_n8397.n251 0.136625
R49112 a_71281_n8397.n256 a_71281_n8397.n255 0.136625
R49113 a_71281_n8397.n248 a_71281_n8397.n237 0.136625
R49114 a_71281_n8397.n242 a_71281_n8397.n241 0.136625
R49115 a_71281_n8397.n231 a_71281_n8397.n220 0.136625
R49116 a_71281_n8397.n225 a_71281_n8397.n224 0.136625
R49117 a_71281_n8397.n217 a_71281_n8397.n206 0.136625
R49118 a_71281_n8397.n211 a_71281_n8397.n210 0.136625
R49119 a_71281_n8397.n200 a_71281_n8397.n189 0.136625
R49120 a_71281_n8397.n194 a_71281_n8397.n193 0.136625
R49121 a_71281_n8397.n186 a_71281_n8397.n175 0.136625
R49122 a_71281_n8397.n180 a_71281_n8397.n179 0.136625
R49123 a_71281_n8397.n422 a_71281_n8397.n411 0.136625
R49124 a_71281_n8397.n416 a_71281_n8397.n415 0.136625
R49125 a_71281_n8397.n436 a_71281_n8397.n425 0.136625
R49126 a_71281_n8397.n430 a_71281_n8397.n429 0.136625
R49127 a_71281_n8397.n458 a_71281_n8397.n456 0.136625
R49128 a_71281_n8397.n463 a_71281_n8397.n452 0.136625
R49129 a_71281_n8397.n443 a_71281_n8397.n438 0.136625
R49130 a_71281_n8397.n449 a_71281_n8397.n439 0.136625
R49131 a_71281_n8397.n298 a_71281_n8397.n293 0.136625
R49132 a_71281_n8397.n304 a_71281_n8397.n294 0.136625
R49133 a_71281_n8397.n313 a_71281_n8397.n311 0.136625
R49134 a_71281_n8397.n318 a_71281_n8397.n307 0.136625
R49135 a_71281_n8397.n327 a_71281_n8397.n325 0.136625
R49136 a_71281_n8397.n332 a_71281_n8397.n321 0.136625
R49137 a_71281_n8397.n341 a_71281_n8397.n339 0.136625
R49138 a_71281_n8397.n346 a_71281_n8397.n335 0.136625
R49139 a_71281_n8397.n358 a_71281_n8397.n356 0.136625
R49140 a_71281_n8397.n363 a_71281_n8397.n352 0.136625
R49141 a_71281_n8397.n372 a_71281_n8397.n370 0.136625
R49142 a_71281_n8397.n377 a_71281_n8397.n366 0.136625
R49143 a_71281_n8397.n389 a_71281_n8397.n387 0.136625
R49144 a_71281_n8397.n394 a_71281_n8397.n383 0.136625
R49145 a_71281_n8397.n403 a_71281_n8397.n401 0.136625
R49146 a_71281_n8397.n408 a_71281_n8397.n397 0.136625
R49147 a_71281_n8397.n581 a_71281_n8397.n570 0.136625
R49148 a_71281_n8397.n575 a_71281_n8397.n574 0.136625
R49149 a_71281_n8397.n567 a_71281_n8397.n556 0.136625
R49150 a_71281_n8397.n561 a_71281_n8397.n560 0.136625
R49151 a_71281_n8397.n553 a_71281_n8397.n542 0.136625
R49152 a_71281_n8397.n547 a_71281_n8397.n546 0.136625
R49153 a_71281_n8397.n539 a_71281_n8397.n528 0.136625
R49154 a_71281_n8397.n533 a_71281_n8397.n532 0.136625
R49155 a_71281_n8397.n522 a_71281_n8397.n511 0.136625
R49156 a_71281_n8397.n516 a_71281_n8397.n515 0.136625
R49157 a_71281_n8397.n508 a_71281_n8397.n497 0.136625
R49158 a_71281_n8397.n502 a_71281_n8397.n501 0.136625
R49159 a_71281_n8397.n491 a_71281_n8397.n480 0.136625
R49160 a_71281_n8397.n485 a_71281_n8397.n484 0.136625
R49161 a_71281_n8397.n477 a_71281_n8397.n466 0.136625
R49162 a_71281_n8397.n471 a_71281_n8397.n470 0.136625
R49163 a_71281_n8397.n738 a_71281_n8397.n736 0.136625
R49164 a_71281_n8397.n743 a_71281_n8397.n732 0.136625
R49165 a_71281_n8397.n752 a_71281_n8397.n750 0.136625
R49166 a_71281_n8397.n757 a_71281_n8397.n746 0.136625
R49167 a_71281_n8397.n766 a_71281_n8397.n764 0.136625
R49168 a_71281_n8397.n771 a_71281_n8397.n760 0.136625
R49169 a_71281_n8397.n780 a_71281_n8397.n778 0.136625
R49170 a_71281_n8397.n785 a_71281_n8397.n774 0.136625
R49171 a_71281_n8397.n871 a_71281_n8397.n860 0.136625
R49172 a_71281_n8397.n865 a_71281_n8397.n864 0.136625
R49173 a_71281_n8397.n857 a_71281_n8397.n846 0.136625
R49174 a_71281_n8397.n851 a_71281_n8397.n850 0.136625
R49175 a_71281_n8397.n840 a_71281_n8397.n829 0.136625
R49176 a_71281_n8397.n834 a_71281_n8397.n833 0.136625
R49177 a_71281_n8397.n826 a_71281_n8397.n815 0.136625
R49178 a_71281_n8397.n820 a_71281_n8397.n819 0.136625
R49179 a_71281_n8397.n15 a_71281_n8397.n14 0.095973
R49180 a_71281_n8397.n29 a_71281_n8397.n28 0.095973
R49181 a_71281_n8397.n43 a_71281_n8397.n42 0.095973
R49182 a_71281_n8397.n74 a_71281_n8397.n73 0.095973
R49183 a_71281_n8397.n105 a_71281_n8397.n104 0.095973
R49184 a_71281_n8397.n119 a_71281_n8397.n118 0.095973
R49185 a_71281_n8397.n133 a_71281_n8397.n132 0.095973
R49186 a_71281_n8397.n278 a_71281_n8397.n277 0.095973
R49187 a_71281_n8397.n264 a_71281_n8397.n263 0.095973
R49188 a_71281_n8397.n250 a_71281_n8397.n249 0.095973
R49189 a_71281_n8397.n219 a_71281_n8397.n218 0.095973
R49190 a_71281_n8397.n188 a_71281_n8397.n187 0.095973
R49191 a_71281_n8397.n174 a_71281_n8397.n173 0.095973
R49192 a_71281_n8397.n160 a_71281_n8397.n159 0.095973
R49193 a_71281_n8397.n306 a_71281_n8397.n305 0.095973
R49194 a_71281_n8397.n320 a_71281_n8397.n319 0.095973
R49195 a_71281_n8397.n334 a_71281_n8397.n333 0.095973
R49196 a_71281_n8397.n365 a_71281_n8397.n364 0.095973
R49197 a_71281_n8397.n396 a_71281_n8397.n395 0.095973
R49198 a_71281_n8397.n410 a_71281_n8397.n409 0.095973
R49199 a_71281_n8397.n424 a_71281_n8397.n423 0.095973
R49200 a_71281_n8397.n569 a_71281_n8397.n568 0.095973
R49201 a_71281_n8397.n555 a_71281_n8397.n554 0.095973
R49202 a_71281_n8397.n541 a_71281_n8397.n540 0.095973
R49203 a_71281_n8397.n510 a_71281_n8397.n509 0.095973
R49204 a_71281_n8397.n479 a_71281_n8397.n478 0.095973
R49205 a_71281_n8397.n465 a_71281_n8397.n464 0.095973
R49206 a_71281_n8397.n451 a_71281_n8397.n450 0.095973
R49207 a_71281_n8397.n599 a_71281_n8397.n598 0.095973
R49208 a_71281_n8397.n613 a_71281_n8397.n612 0.095973
R49209 a_71281_n8397.n627 a_71281_n8397.n626 0.095973
R49210 a_71281_n8397.n658 a_71281_n8397.n657 0.095973
R49211 a_71281_n8397.n689 a_71281_n8397.n688 0.095973
R49212 a_71281_n8397.n703 a_71281_n8397.n702 0.095973
R49213 a_71281_n8397.n717 a_71281_n8397.n716 0.095973
R49214 a_71281_n8397.n745 a_71281_n8397.n744 0.095973
R49215 a_71281_n8397.n759 a_71281_n8397.n758 0.095973
R49216 a_71281_n8397.n773 a_71281_n8397.n772 0.095973
R49217 a_71281_n8397.n859 a_71281_n8397.n858 0.095973
R49218 a_71281_n8397.n828 a_71281_n8397.n827 0.095973
R49219 a_71281_n8397.n814 a_71281_n8397.n813 0.095973
R49220 a_71281_n8397.n800 a_71281_n8397.n799 0.095973
R49221 a_71281_n8397.n715 a_71281_n8397.n714 0.0719743
R49222 a_71281_n8397.n711 a_71281_n8397.n709 0.0719743
R49223 a_71281_n8397.n729 a_71281_n8397.n728 0.0719743
R49224 a_71281_n8397.n725 a_71281_n8397.n723 0.0719743
R49225 a_71281_n8397.n808 a_71281_n8397.n807 0.0719743
R49226 a_71281_n8397.n812 a_71281_n8397.n811 0.0719743
R49227 a_71281_n8397.n794 a_71281_n8397.n787 0.0719743
R49228 a_71281_n8397.n798 a_71281_n8397.n797 0.0719743
R49229 a_71281_n8397.n593 a_71281_n8397.n586 0.0719743
R49230 a_71281_n8397.n597 a_71281_n8397.n596 0.0719743
R49231 a_71281_n8397.n607 a_71281_n8397.n606 0.0719743
R49232 a_71281_n8397.n611 a_71281_n8397.n610 0.0719743
R49233 a_71281_n8397.n621 a_71281_n8397.n620 0.0719743
R49234 a_71281_n8397.n625 a_71281_n8397.n624 0.0719743
R49235 a_71281_n8397.n635 a_71281_n8397.n634 0.0719743
R49236 a_71281_n8397.n639 a_71281_n8397.n638 0.0719743
R49237 a_71281_n8397.n652 a_71281_n8397.n651 0.0719743
R49238 a_71281_n8397.n656 a_71281_n8397.n655 0.0719743
R49239 a_71281_n8397.n666 a_71281_n8397.n665 0.0719743
R49240 a_71281_n8397.n670 a_71281_n8397.n669 0.0719743
R49241 a_71281_n8397.n683 a_71281_n8397.n682 0.0719743
R49242 a_71281_n8397.n687 a_71281_n8397.n686 0.0719743
R49243 a_71281_n8397.n697 a_71281_n8397.n696 0.0719743
R49244 a_71281_n8397.n701 a_71281_n8397.n700 0.0719743
R49245 a_71281_n8397.n131 a_71281_n8397.n130 0.0719743
R49246 a_71281_n8397.n127 a_71281_n8397.n125 0.0719743
R49247 a_71281_n8397.n145 a_71281_n8397.n144 0.0719743
R49248 a_71281_n8397.n141 a_71281_n8397.n139 0.0719743
R49249 a_71281_n8397.n168 a_71281_n8397.n167 0.0719743
R49250 a_71281_n8397.n172 a_71281_n8397.n171 0.0719743
R49251 a_71281_n8397.n154 a_71281_n8397.n147 0.0719743
R49252 a_71281_n8397.n158 a_71281_n8397.n157 0.0719743
R49253 a_71281_n8397.n9 a_71281_n8397.n2 0.0719743
R49254 a_71281_n8397.n13 a_71281_n8397.n12 0.0719743
R49255 a_71281_n8397.n23 a_71281_n8397.n22 0.0719743
R49256 a_71281_n8397.n27 a_71281_n8397.n26 0.0719743
R49257 a_71281_n8397.n37 a_71281_n8397.n36 0.0719743
R49258 a_71281_n8397.n41 a_71281_n8397.n40 0.0719743
R49259 a_71281_n8397.n51 a_71281_n8397.n50 0.0719743
R49260 a_71281_n8397.n55 a_71281_n8397.n54 0.0719743
R49261 a_71281_n8397.n68 a_71281_n8397.n67 0.0719743
R49262 a_71281_n8397.n72 a_71281_n8397.n71 0.0719743
R49263 a_71281_n8397.n82 a_71281_n8397.n81 0.0719743
R49264 a_71281_n8397.n86 a_71281_n8397.n85 0.0719743
R49265 a_71281_n8397.n99 a_71281_n8397.n98 0.0719743
R49266 a_71281_n8397.n103 a_71281_n8397.n102 0.0719743
R49267 a_71281_n8397.n113 a_71281_n8397.n112 0.0719743
R49268 a_71281_n8397.n117 a_71281_n8397.n116 0.0719743
R49269 a_71281_n8397.n290 a_71281_n8397.n289 0.0719743
R49270 a_71281_n8397.n286 a_71281_n8397.n284 0.0719743
R49271 a_71281_n8397.n276 a_71281_n8397.n275 0.0719743
R49272 a_71281_n8397.n272 a_71281_n8397.n270 0.0719743
R49273 a_71281_n8397.n262 a_71281_n8397.n261 0.0719743
R49274 a_71281_n8397.n258 a_71281_n8397.n256 0.0719743
R49275 a_71281_n8397.n248 a_71281_n8397.n247 0.0719743
R49276 a_71281_n8397.n244 a_71281_n8397.n242 0.0719743
R49277 a_71281_n8397.n231 a_71281_n8397.n230 0.0719743
R49278 a_71281_n8397.n227 a_71281_n8397.n225 0.0719743
R49279 a_71281_n8397.n217 a_71281_n8397.n216 0.0719743
R49280 a_71281_n8397.n213 a_71281_n8397.n211 0.0719743
R49281 a_71281_n8397.n200 a_71281_n8397.n199 0.0719743
R49282 a_71281_n8397.n196 a_71281_n8397.n194 0.0719743
R49283 a_71281_n8397.n186 a_71281_n8397.n185 0.0719743
R49284 a_71281_n8397.n182 a_71281_n8397.n180 0.0719743
R49285 a_71281_n8397.n422 a_71281_n8397.n421 0.0719743
R49286 a_71281_n8397.n418 a_71281_n8397.n416 0.0719743
R49287 a_71281_n8397.n436 a_71281_n8397.n435 0.0719743
R49288 a_71281_n8397.n432 a_71281_n8397.n430 0.0719743
R49289 a_71281_n8397.n459 a_71281_n8397.n458 0.0719743
R49290 a_71281_n8397.n463 a_71281_n8397.n462 0.0719743
R49291 a_71281_n8397.n445 a_71281_n8397.n438 0.0719743
R49292 a_71281_n8397.n449 a_71281_n8397.n448 0.0719743
R49293 a_71281_n8397.n300 a_71281_n8397.n293 0.0719743
R49294 a_71281_n8397.n304 a_71281_n8397.n303 0.0719743
R49295 a_71281_n8397.n314 a_71281_n8397.n313 0.0719743
R49296 a_71281_n8397.n318 a_71281_n8397.n317 0.0719743
R49297 a_71281_n8397.n328 a_71281_n8397.n327 0.0719743
R49298 a_71281_n8397.n332 a_71281_n8397.n331 0.0719743
R49299 a_71281_n8397.n342 a_71281_n8397.n341 0.0719743
R49300 a_71281_n8397.n346 a_71281_n8397.n345 0.0719743
R49301 a_71281_n8397.n359 a_71281_n8397.n358 0.0719743
R49302 a_71281_n8397.n363 a_71281_n8397.n362 0.0719743
R49303 a_71281_n8397.n373 a_71281_n8397.n372 0.0719743
R49304 a_71281_n8397.n377 a_71281_n8397.n376 0.0719743
R49305 a_71281_n8397.n390 a_71281_n8397.n389 0.0719743
R49306 a_71281_n8397.n394 a_71281_n8397.n393 0.0719743
R49307 a_71281_n8397.n404 a_71281_n8397.n403 0.0719743
R49308 a_71281_n8397.n408 a_71281_n8397.n407 0.0719743
R49309 a_71281_n8397.n581 a_71281_n8397.n580 0.0719743
R49310 a_71281_n8397.n577 a_71281_n8397.n575 0.0719743
R49311 a_71281_n8397.n567 a_71281_n8397.n566 0.0719743
R49312 a_71281_n8397.n563 a_71281_n8397.n561 0.0719743
R49313 a_71281_n8397.n553 a_71281_n8397.n552 0.0719743
R49314 a_71281_n8397.n549 a_71281_n8397.n547 0.0719743
R49315 a_71281_n8397.n539 a_71281_n8397.n538 0.0719743
R49316 a_71281_n8397.n535 a_71281_n8397.n533 0.0719743
R49317 a_71281_n8397.n522 a_71281_n8397.n521 0.0719743
R49318 a_71281_n8397.n518 a_71281_n8397.n516 0.0719743
R49319 a_71281_n8397.n508 a_71281_n8397.n507 0.0719743
R49320 a_71281_n8397.n504 a_71281_n8397.n502 0.0719743
R49321 a_71281_n8397.n491 a_71281_n8397.n490 0.0719743
R49322 a_71281_n8397.n487 a_71281_n8397.n485 0.0719743
R49323 a_71281_n8397.n477 a_71281_n8397.n476 0.0719743
R49324 a_71281_n8397.n473 a_71281_n8397.n471 0.0719743
R49325 a_71281_n8397.n739 a_71281_n8397.n738 0.0719743
R49326 a_71281_n8397.n743 a_71281_n8397.n742 0.0719743
R49327 a_71281_n8397.n753 a_71281_n8397.n752 0.0719743
R49328 a_71281_n8397.n757 a_71281_n8397.n756 0.0719743
R49329 a_71281_n8397.n767 a_71281_n8397.n766 0.0719743
R49330 a_71281_n8397.n771 a_71281_n8397.n770 0.0719743
R49331 a_71281_n8397.n781 a_71281_n8397.n780 0.0719743
R49332 a_71281_n8397.n785 a_71281_n8397.n784 0.0719743
R49333 a_71281_n8397.n871 a_71281_n8397.n870 0.0719743
R49334 a_71281_n8397.n867 a_71281_n8397.n865 0.0719743
R49335 a_71281_n8397.n857 a_71281_n8397.n856 0.0719743
R49336 a_71281_n8397.n853 a_71281_n8397.n851 0.0719743
R49337 a_71281_n8397.n840 a_71281_n8397.n839 0.0719743
R49338 a_71281_n8397.n836 a_71281_n8397.n834 0.0719743
R49339 a_71281_n8397.n826 a_71281_n8397.n825 0.0719743
R49340 a_71281_n8397.n822 a_71281_n8397.n820 0.0719743
R49341 a_71281_n8397.n60 a_71281_n8397.n59 0.0485405
R49342 a_71281_n8397.n235 a_71281_n8397.n232 0.0485405
R49343 a_71281_n8397.n351 a_71281_n8397.n350 0.0485405
R49344 a_71281_n8397.n526 a_71281_n8397.n523 0.0485405
R49345 a_71281_n8397.n644 a_71281_n8397.n643 0.0485405
R49346 a_71281_n8397.n873 a_71281_n8397.n872 0.0485405
R49347 a_71281_n8397.n90 a_71281_n8397.n87 0.0482365
R49348 a_71281_n8397.n91 a_71281_n8397.n90 0.0482365
R49349 a_71281_n8397.n205 a_71281_n8397.n204 0.0482365
R49350 a_71281_n8397.n204 a_71281_n8397.n201 0.0482365
R49351 a_71281_n8397.n381 a_71281_n8397.n378 0.0482365
R49352 a_71281_n8397.n382 a_71281_n8397.n381 0.0482365
R49353 a_71281_n8397.n496 a_71281_n8397.n495 0.0482365
R49354 a_71281_n8397.n495 a_71281_n8397.n492 0.0482365
R49355 a_71281_n8397.n674 a_71281_n8397.n671 0.0482365
R49356 a_71281_n8397.n675 a_71281_n8397.n674 0.0482365
R49357 a_71281_n8397.n845 a_71281_n8397.n844 0.0482365
R49358 a_71281_n8397.n844 a_71281_n8397.n841 0.0482365
R49359 a_71281_n8397.n59 a_71281_n8397.n56 0.0479324
R49360 a_71281_n8397.n236 a_71281_n8397.n235 0.0479324
R49361 a_71281_n8397.n350 a_71281_n8397.n347 0.0479324
R49362 a_71281_n8397.n527 a_71281_n8397.n526 0.0479324
R49363 a_71281_n8397.n643 a_71281_n8397.n640 0.0479324
R49364 a_71281_n8397.n873 a_71281_n8397.n786 0.0479324
R49365 a_71281_n8397.n731 a_71281_n8397.n1 0.443549
R49366 a_35922_19591.n237 a_35922_19591.n230 10.6966
R49367 a_35922_19591.n234 a_35922_19591.t104 8.75329
R49368 a_35922_19591.n236 a_35922_19591.t86 8.75329
R49369 a_35922_19591.n233 a_35922_19591.t99 8.75329
R49370 a_35922_19591.n235 a_35922_19591.t51 8.75329
R49371 a_35922_19591.n143 a_35922_19591.t38 8.38704
R49372 a_35922_19591.n132 a_35922_19591.t64 8.38704
R49373 a_35922_19591.n100 a_35922_19591.t150 8.46135
R49374 a_35922_19591.n101 a_35922_19591.t155 8.46135
R49375 a_35922_19591.n0 a_35922_19591.t14 8.39293
R49376 a_35922_19591.n109 a_35922_19591.t168 8.39293
R49377 a_35922_19591.n59 a_35922_19591.t132 8.26625
R49378 a_35922_19591.n61 a_35922_19591.t102 8.26625
R49379 a_35922_19591.n62 a_35922_19591.t71 8.26625
R49380 a_35922_19591.n234 a_35922_19591.t61 8.12045
R49381 a_35922_19591.n236 a_35922_19591.t29 8.12045
R49382 a_35922_19591.n233 a_35922_19591.t58 8.12045
R49383 a_35922_19591.n232 a_35922_19591.t124 8.12045
R49384 a_35922_19591.n235 a_35922_19591.t149 8.12045
R49385 a_35922_19591.n90 a_35922_19591.t80 8.10567
R49386 a_35922_19591.n72 a_35922_19591.t173 8.10567
R49387 a_35922_19591.n72 a_35922_19591.t122 8.10567
R49388 a_35922_19591.n72 a_35922_19591.t84 8.10567
R49389 a_35922_19591.n72 a_35922_19591.t183 8.10567
R49390 a_35922_19591.n31 a_35922_19591.t191 8.10567
R49391 a_35922_19591.n31 a_35922_19591.t13 8.10567
R49392 a_35922_19591.n31 a_35922_19591.t138 8.10567
R49393 a_35922_19591.n31 a_35922_19591.t52 8.10567
R49394 a_35922_19591.n34 a_35922_19591.t15 8.10567
R49395 a_35922_19591.n34 a_35922_19591.t174 8.10567
R49396 a_35922_19591.n34 a_35922_19591.t125 8.10567
R49397 a_35922_19591.n34 a_35922_19591.t26 8.10567
R49398 a_35922_19591.n70 a_35922_19591.t59 8.10567
R49399 a_35922_19591.n70 a_35922_19591.t128 8.10567
R49400 a_35922_19591.n70 a_35922_19591.t76 8.10567
R49401 a_35922_19591.n68 a_35922_19591.t74 8.10567
R49402 a_35922_19591.n68 a_35922_19591.t143 8.10567
R49403 a_35922_19591.n68 a_35922_19591.t131 8.10567
R49404 a_35922_19591.n90 a_35922_19591.t45 8.10567
R49405 a_35922_19591.n90 a_35922_19591.t147 8.10567
R49406 a_35922_19591.n90 a_35922_19591.t44 8.10567
R49407 a_35922_19591.n99 a_35922_19591.t77 8.10567
R49408 a_35922_19591.n86 a_35922_19591.t163 8.10567
R49409 a_35922_19591.n86 a_35922_19591.t116 8.10567
R49410 a_35922_19591.n86 a_35922_19591.t82 8.10567
R49411 a_35922_19591.n86 a_35922_19591.t170 8.10567
R49412 a_35922_19591.n48 a_35922_19591.t178 8.10567
R49413 a_35922_19591.n48 a_35922_19591.t187 8.10567
R49414 a_35922_19591.n48 a_35922_19591.t134 8.10567
R49415 a_35922_19591.n48 a_35922_19591.t37 8.10567
R49416 a_35922_19591.n50 a_35922_19591.t190 8.10567
R49417 a_35922_19591.n50 a_35922_19591.t165 8.10567
R49418 a_35922_19591.n50 a_35922_19591.t117 8.10567
R49419 a_35922_19591.n50 a_35922_19591.t12 8.10567
R49420 a_35922_19591.n82 a_35922_19591.t182 8.10567
R49421 a_35922_19591.n82 a_35922_19591.t87 8.10567
R49422 a_35922_19591.n82 a_35922_19591.t33 8.10567
R49423 a_35922_19591.n80 a_35922_19591.t25 8.10567
R49424 a_35922_19591.n80 a_35922_19591.t98 8.10567
R49425 a_35922_19591.n80 a_35922_19591.t89 8.10567
R49426 a_35922_19591.n99 a_35922_19591.t31 8.10567
R49427 a_35922_19591.n99 a_35922_19591.t144 8.10567
R49428 a_35922_19591.n99 a_35922_19591.t30 8.10567
R49429 a_35922_19591.n91 a_35922_19591.t70 8.10567
R49430 a_35922_19591.n74 a_35922_19591.t152 8.10567
R49431 a_35922_19591.n74 a_35922_19591.t101 8.10567
R49432 a_35922_19591.n74 a_35922_19591.t75 8.10567
R49433 a_35922_19591.n74 a_35922_19591.t158 8.10567
R49434 a_35922_19591.n39 a_35922_19591.t160 8.10567
R49435 a_35922_19591.n39 a_35922_19591.t167 8.10567
R49436 a_35922_19591.n39 a_35922_19591.t119 8.10567
R49437 a_35922_19591.n39 a_35922_19591.t19 8.10567
R49438 a_35922_19591.n43 a_35922_19591.t169 8.10567
R49439 a_35922_19591.n43 a_35922_19591.t154 8.10567
R49440 a_35922_19591.n43 a_35922_19591.t103 8.10567
R49441 a_35922_19591.n43 a_35922_19591.t181 8.10567
R49442 a_35922_19591.n66 a_35922_19591.t34 8.10567
R49443 a_35922_19591.n66 a_35922_19591.t105 8.10567
R49444 a_35922_19591.n66 a_35922_19591.t62 8.10567
R49445 a_35922_19591.n64 a_35922_19591.t57 8.10567
R49446 a_35922_19591.n64 a_35922_19591.t123 8.10567
R49447 a_35922_19591.n64 a_35922_19591.t108 8.10567
R49448 a_35922_19591.n91 a_35922_19591.t9 8.10567
R49449 a_35922_19591.n91 a_35922_19591.t137 8.10567
R49450 a_35922_19591.n91 a_35922_19591.t8 8.10567
R49451 a_35922_19591.n94 a_35922_19591.t81 8.10567
R49452 a_35922_19591.n84 a_35922_19591.t176 8.10567
R49453 a_35922_19591.n84 a_35922_19591.t127 8.10567
R49454 a_35922_19591.n84 a_35922_19591.t85 8.10567
R49455 a_35922_19591.n84 a_35922_19591.t185 8.10567
R49456 a_35922_19591.n54 a_35922_19591.t193 8.10567
R49457 a_35922_19591.n54 a_35922_19591.t17 8.10567
R49458 a_35922_19591.n54 a_35922_19591.t141 8.10567
R49459 a_35922_19591.n54 a_35922_19591.t55 8.10567
R49460 a_35922_19591.n56 a_35922_19591.t21 8.10567
R49461 a_35922_19591.n56 a_35922_19591.t180 8.10567
R49462 a_35922_19591.n56 a_35922_19591.t130 8.10567
R49463 a_35922_19591.n56 a_35922_19591.t28 8.10567
R49464 a_35922_19591.n78 a_35922_19591.t11 8.10567
R49465 a_35922_19591.n78 a_35922_19591.t92 8.10567
R49466 a_35922_19591.n78 a_35922_19591.t50 8.10567
R49467 a_35922_19591.n76 a_35922_19591.t42 8.10567
R49468 a_35922_19591.n76 a_35922_19591.t113 8.10567
R49469 a_35922_19591.n76 a_35922_19591.t93 8.10567
R49470 a_35922_19591.n94 a_35922_19591.t49 8.10567
R49471 a_35922_19591.n94 a_35922_19591.t148 8.10567
R49472 a_35922_19591.n94 a_35922_19591.t47 8.10567
R49473 a_35922_19591.n0 a_35922_19591.t32 8.10567
R49474 a_35922_19591.n0 a_35922_19591.t43 8.10567
R49475 a_35922_19591.n0 a_35922_19591.t146 8.10567
R49476 a_35922_19591.n0 a_35922_19591.t69 8.10567
R49477 a_35922_19591.n0 a_35922_19591.t36 8.10567
R49478 a_35922_19591.n0 a_35922_19591.t109 8.10567
R49479 a_35922_19591.n0 a_35922_19591.t66 8.10567
R49480 a_35922_19591.n0 a_35922_19591.t94 8.10567
R49481 a_35922_19591.n0 a_35922_19591.t24 8.10567
R49482 a_35922_19591.n105 a_35922_19591.t88 8.10567
R49483 a_35922_19591.n103 a_35922_19591.t65 8.10567
R49484 a_35922_19591.n131 a_35922_19591.t157 8.10567
R49485 a_35922_19591.n2 a_35922_19591.t60 8.10567
R49486 a_35922_19591.n228 a_35922_19591.t129 8.10567
R49487 a_35922_19591.n227 a_35922_19591.t111 8.10567
R49488 a_35922_19591.n3 a_35922_19591.t46 8.10567
R49489 a_35922_19591.n3 a_35922_19591.t16 8.10567
R49490 a_35922_19591.n3 a_35922_19591.t140 8.10567
R49491 a_35922_19591.n3 a_35922_19591.t54 8.10567
R49492 a_35922_19591.n12 a_35922_19591.t156 8.10567
R49493 a_35922_19591.n12 a_35922_19591.t162 8.10567
R49494 a_35922_19591.n12 a_35922_19591.t115 8.10567
R49495 a_35922_19591.n12 a_35922_19591.t6 8.10567
R49496 a_35922_19591.n27 a_35922_19591.t23 8.10567
R49497 a_35922_19591.n162 a_35922_19591.t97 8.10567
R49498 a_35922_19591.n161 a_35922_19591.t56 8.10567
R49499 a_35922_19591.n28 a_35922_19591.t95 8.10567
R49500 a_35922_19591.n29 a_35922_19591.t73 8.10567
R49501 a_35922_19591.n29 a_35922_19591.t153 8.10567
R49502 a_35922_19591.n4 a_35922_19591.t67 8.10567
R49503 a_35922_19591.n4 a_35922_19591.t189 8.10567
R49504 a_35922_19591.n4 a_35922_19591.t135 8.10567
R49505 a_35922_19591.n25 a_35922_19591.t53 8.10567
R49506 a_35922_19591.n160 a_35922_19591.t118 8.10567
R49507 a_35922_19591.n159 a_35922_19591.t100 8.10567
R49508 a_35922_19591.n17 a_35922_19591.t164 8.10567
R49509 a_35922_19591.n17 a_35922_19591.t151 8.10567
R49510 a_35922_19591.n16 a_35922_19591.t96 8.10567
R49511 a_35922_19591.n16 a_35922_19591.t171 8.10567
R49512 a_35922_19591.n112 a_35922_19591.t184 8.10567
R49513 a_35922_19591.n111 a_35922_19591.t7 8.10567
R49514 a_35922_19591.n110 a_35922_19591.t136 8.10567
R49515 a_35922_19591.n194 a_35922_19591.t48 8.10567
R49516 a_35922_19591.n177 a_35922_19591.t192 8.10567
R49517 a_35922_19591.n178 a_35922_19591.t90 8.10567
R49518 a_35922_19591.n179 a_35922_19591.t41 8.10567
R49519 a_35922_19591.n108 a_35922_19591.t120 8.10567
R49520 a_35922_19591.n107 a_35922_19591.t83 8.10567
R49521 a_35922_19591.n106 a_35922_19591.t179 8.10567
R49522 a_35922_19591.n126 a_35922_19591.t79 8.10567
R49523 a_35922_19591.n124 a_35922_19591.t39 8.10567
R49524 a_35922_19591.n142 a_35922_19591.t145 8.10567
R49525 a_35922_19591.n153 a_35922_19591.t35 8.10567
R49526 a_35922_19591.n152 a_35922_19591.t106 8.10567
R49527 a_35922_19591.n151 a_35922_19591.t91 8.10567
R49528 a_35922_19591.n120 a_35922_19591.t10 8.10567
R49529 a_35922_19591.n119 a_35922_19591.t172 8.10567
R49530 a_35922_19591.n118 a_35922_19591.t121 8.10567
R49531 a_35922_19591.n115 a_35922_19591.t22 8.10567
R49532 a_35922_19591.n10 a_35922_19591.t166 8.10567
R49533 a_35922_19591.n10 a_35922_19591.t175 8.10567
R49534 a_35922_19591.n10 a_35922_19591.t126 8.10567
R49535 a_35922_19591.n10 a_35922_19591.t27 8.10567
R49536 a_35922_19591.n212 a_35922_19591.t40 8.10567
R49537 a_35922_19591.n213 a_35922_19591.t112 8.10567
R49538 a_35922_19591.n9 a_35922_19591.t68 8.10567
R49539 a_35922_19591.n22 a_35922_19591.t107 8.10567
R49540 a_35922_19591.n23 a_35922_19591.t78 8.10567
R49541 a_35922_19591.n23 a_35922_19591.t161 8.10567
R49542 a_35922_19591.n8 a_35922_19591.t72 8.10567
R49543 a_35922_19591.n8 a_35922_19591.t20 8.10567
R49544 a_35922_19591.n8 a_35922_19591.t142 8.10567
R49545 a_35922_19591.n19 a_35922_19591.t63 8.10567
R49546 a_35922_19591.n210 a_35922_19591.t133 8.10567
R49547 a_35922_19591.n209 a_35922_19591.t114 8.10567
R49548 a_35922_19591.n14 a_35922_19591.t177 8.10567
R49549 a_35922_19591.n14 a_35922_19591.t159 8.10567
R49550 a_35922_19591.n20 a_35922_19591.t110 8.10567
R49551 a_35922_19591.n20 a_35922_19591.t186 8.10567
R49552 a_35922_19591.n231 a_35922_19591.t0 6.69607
R49553 a_35922_19591.n240 a_35922_19591.t2 6.0467
R49554 a_35922_19591.n231 a_35922_19591.t1 5.54843
R49555 a_35922_19591.n238 a_35922_19591.t3 5.44096
R49556 a_35922_19591.n238 a_35922_19591.t4 5.41626
R49557 a_35922_19591.n239 a_35922_19591.n237 4.8989
R49558 a_35922_19591.t5 a_35922_19591.n240 4.79524
R49559 a_35922_19591.n1 a_35922_19591.n3 0.426349
R49560 a_35922_19591.n121 a_35922_19591.n120 2.25163
R49561 a_35922_19591.n18 a_35922_19591.n17 0.607617
R49562 a_35922_19591.n15 a_35922_19591.n14 0.607617
R49563 a_35922_19591.n86 a_35922_19591.n87 0.020246
R49564 a_35922_19591.n85 a_35922_19591.n84 0.020246
R49565 a_35922_19591.n48 a_35922_19591.n47 0.150783
R49566 a_35922_19591.n50 a_35922_19591.n46 0.150803
R49567 a_35922_19591.n99 a_35922_19591.n98 0.0676355
R49568 a_35922_19591.n54 a_35922_19591.n53 0.150803
R49569 a_35922_19591.n58 a_35922_19591.n56 0.150806
R49570 a_35922_19591.n95 a_35922_19591.n94 0.0676255
R49571 a_35922_19591.n34 a_35922_19591.n35 0.153625
R49572 a_35922_19591.n31 a_35922_19591.n32 0.153625
R49573 a_35922_19591.n73 a_35922_19591.n72 0.020088
R49574 a_35922_19591.n51 a_35922_19591.n50 0.246907
R49575 a_35922_19591.n48 a_35922_19591.n49 0.246877
R49576 a_35922_19591.n44 a_35922_19591.n43 0.153625
R49577 a_35922_19591.n40 a_35922_19591.n39 0.153625
R49578 a_35922_19591.n74 a_35922_19591.n75 0.020088
R49579 a_35922_19591.n91 a_35922_19591.n92 0.0201939
R49580 a_35922_19591.n43 a_35922_19591.n42 0.246907
R49581 a_35922_19591.n39 a_35922_19591.n38 0.246907
R49582 a_35922_19591.n56 a_35922_19591.n57 0.246907
R49583 a_35922_19591.n55 a_35922_19591.n54 0.246907
R49584 a_35922_19591.n90 a_35922_19591.n89 0.0201939
R49585 a_35922_19591.n36 a_35922_19591.n34 0.246907
R49586 a_35922_19591.n33 a_35922_19591.n31 0.246907
R49587 a_35922_19591.n4 a_35922_19591.n5 0.260442
R49588 a_35922_19591.n26 a_35922_19591.n16 0.591264
R49589 a_35922_19591.n12 a_35922_19591.n13 0.310971
R49590 a_35922_19591.n30 a_35922_19591.n29 0.591264
R49591 a_35922_19591.n28 a_35922_19591.n100 0.332154
R49592 a_35922_19591.n150 a_35922_19591.n140 4.5005
R49593 a_35922_19591.n126 a_35922_19591.n149 4.5005
R49594 a_35922_19591.n148 a_35922_19591.n125 4.5005
R49595 a_35922_19591.n147 a_35922_19591.n146 4.5005
R49596 a_35922_19591.n124 a_35922_19591.n122 4.5005
R49597 a_35922_19591.n123 a_35922_19591.n145 4.5005
R49598 a_35922_19591.n144 a_35922_19591.n141 4.5005
R49599 a_35922_19591.n206 a_35922_19591.n205 4.5005
R49600 a_35922_19591.n115 a_35922_19591.n113 4.5005
R49601 a_35922_19591.n114 a_35922_19591.n204 4.5005
R49602 a_35922_19591.n203 a_35922_19591.n116 4.5005
R49603 a_35922_19591.n202 a_35922_19591.n118 4.5005
R49604 a_35922_19591.n117 a_35922_19591.n154 4.5005
R49605 a_35922_19591.n201 a_35922_19591.n200 4.5005
R49606 a_35922_19591.n199 a_35922_19591.n119 4.5005
R49607 a_35922_19591.n198 a_35922_19591.n197 4.5005
R49608 a_35922_19591.n196 a_35922_19591.n155 4.5005
R49609 a_35922_19591.n181 a_35922_19591.n180 4.5005
R49610 a_35922_19591.n112 a_35922_19591.n182 4.5005
R49611 a_35922_19591.n183 a_35922_19591.n158 4.5005
R49612 a_35922_19591.n185 a_35922_19591.n184 4.5005
R49613 a_35922_19591.n111 a_35922_19591.n186 4.5005
R49614 a_35922_19591.n187 a_35922_19591.n157 4.5005
R49615 a_35922_19591.n189 a_35922_19591.n188 4.5005
R49616 a_35922_19591.n190 a_35922_19591.n110 4.5005
R49617 a_35922_19591.n192 a_35922_19591.n191 4.5005
R49618 a_35922_19591.n193 a_35922_19591.n156 4.5005
R49619 a_35922_19591.n176 a_35922_19591.n175 4.5005
R49620 a_35922_19591.n174 a_35922_19591.n106 4.5005
R49621 a_35922_19591.n173 a_35922_19591.n172 4.5005
R49622 a_35922_19591.n171 a_35922_19591.n165 4.5005
R49623 a_35922_19591.n107 a_35922_19591.n170 4.5005
R49624 a_35922_19591.n169 a_35922_19591.n168 4.5005
R49625 a_35922_19591.n167 a_35922_19591.n166 4.5005
R49626 a_35922_19591.n8 a_35922_19591.n7 0.260442
R49627 a_35922_19591.n21 a_35922_19591.n20 0.591264
R49628 a_35922_19591.n10 a_35922_19591.n11 0.310971
R49629 a_35922_19591.n23 a_35922_19591.n24 0.591264
R49630 a_35922_19591.n22 a_35922_19591.n101 0.332154
R49631 a_35922_19591.n226 a_35922_19591.n225 4.5005
R49632 a_35922_19591.n138 a_35922_19591.n105 4.5005
R49633 a_35922_19591.n104 a_35922_19591.n129 4.5005
R49634 a_35922_19591.n137 a_35922_19591.n136 4.5005
R49635 a_35922_19591.n135 a_35922_19591.n103 4.5005
R49636 a_35922_19591.n102 a_35922_19591.n130 4.5005
R49637 a_35922_19591.n134 a_35922_19591.n133 4.5005
R49638 a_35922_19591.n222 a_35922_19591.n127 3.97759
R49639 a_35922_19591.n240 a_35922_19591.n239 3.0252
R49640 a_35922_19591.n232 a_35922_19591.n231 2.35922
R49641 a_35922_19591.n237 a_35922_19591.n63 2.34557
R49642 a_35922_19591.n208 a_35922_19591.n139 2.30989
R49643 a_35922_19591.n163 a_35922_19591.n93 2.30989
R49644 a_35922_19591.n195 a_35922_19591.n194 2.25752
R49645 a_35922_19591.n71 a_35922_19591.n70 0.427602
R49646 a_35922_19591.n69 a_35922_19591.n68 0.427602
R49647 a_35922_19591.n67 a_35922_19591.n66 0.427602
R49648 a_35922_19591.n65 a_35922_19591.n64 0.427602
R49649 a_35922_19591.n83 a_35922_19591.n82 0.420727
R49650 a_35922_19591.n81 a_35922_19591.n80 0.420727
R49651 a_35922_19591.n79 a_35922_19591.n78 0.420727
R49652 a_35922_19591.n77 a_35922_19591.n76 0.420727
R49653 a_35922_19591.n207 a_35922_19591.n140 2.16725
R49654 a_35922_19591.n181 a_35922_19591.n164 2.16725
R49655 a_35922_19591.n225 a_35922_19591.n224 2.16725
R49656 a_35922_19591.n42 a_35922_19591.n41 2.96488
R49657 a_35922_19591.n37 a_35922_19591.n75 2.94096
R49658 a_35922_19591.n88 a_35922_19591.n36 2.96488
R49659 a_35922_19591.n73 a_35922_19591.n220 2.94096
R49660 a_35922_19591.n222 a_35922_19591.n221 2.09357
R49661 a_35922_19591.n216 a_35922_19591.n97 2.07182
R49662 a_35922_19591.n217 a_35922_19591.n45 2.07182
R49663 a_35922_19591.n97 a_35922_19591.n46 2.75706
R49664 a_35922_19591.n87 a_35922_19591.n45 2.90773
R49665 a_35922_19591.n58 a_35922_19591.n96 2.75704
R49666 a_35922_19591.n52 a_35922_19591.n85 2.90773
R49667 a_35922_19591.n63 a_35922_19591.n60 1.58959
R49668 a_35922_19591.n96 a_35922_19591.n215 1.5005
R49669 a_35922_19591.n41 a_35922_19591.n216 1.5005
R49670 a_35922_19591.n221 a_35922_19591.n88 1.5005
R49671 a_35922_19591.n220 a_35922_19591.n219 1.5005
R49672 a_35922_19591.n218 a_35922_19591.n52 1.5005
R49673 a_35922_19591.n217 a_35922_19591.n37 1.5005
R49674 a_35922_19591.n214 a_35922_19591.n6 1.5005
R49675 a_35922_19591.n208 a_35922_19591.n207 1.5005
R49676 a_35922_19591.n224 a_35922_19591.n223 1.5005
R49677 a_35922_19591.n211 a_35922_19591.n128 1.5005
R49678 a_35922_19591.n164 a_35922_19591.n163 1.5005
R49679 a_35922_19591.n63 a_35922_19591.n62 1.5005
R49680 a_35922_19591.n63 a_35922_19591.n59 1.5005
R49681 a_35922_19591.n239 a_35922_19591.n238 1.5005
R49682 a_35922_19591.n219 a_35922_19591.n127 1.49172
R49683 a_35922_19591.n216 a_35922_19591.n215 1.47516
R49684 a_35922_19591.n218 a_35922_19591.n217 1.47516
R49685 a_35922_19591.n5 a_35922_19591.t188 9.17619
R49686 a_35922_19591.n7 a_35922_19591.t18 9.17619
R49687 a_35922_19591.n223 a_35922_19591.n222 1.37253
R49688 a_35922_19591.n230 a_35922_19591.n229 1.37253
R49689 a_35922_19591.n29 a_35922_19591.n27 1.24866
R49690 a_35922_19591.n16 a_35922_19591.n25 1.24866
R49691 a_35922_19591.n212 a_35922_19591.n23 1.24866
R49692 a_35922_19591.n20 a_35922_19591.n19 1.24866
R49693 a_35922_19591.n159 a_35922_19591.n4 1.24629
R49694 a_35922_19591.n209 a_35922_19591.n8 1.24629
R49695 a_35922_19591.n214 a_35922_19591.n208 1.23709
R49696 a_35922_19591.n163 a_35922_19591.n128 1.23709
R49697 a_35922_19591.n227 a_35922_19591.n226 1.22261
R49698 a_35922_19591.n180 a_35922_19591.n179 1.22261
R49699 a_35922_19591.n151 a_35922_19591.n150 1.22261
R49700 a_35922_19591.n3 a_35922_19591.n2 1.21313
R49701 a_35922_19591.n177 a_35922_19591.n176 1.21313
R49702 a_35922_19591.n205 a_35922_19591.n153 1.21313
R49703 a_35922_19591.n144 a_35922_19591.n143 1.12904
R49704 a_35922_19591.n133 a_35922_19591.n132 1.12904
R49705 a_35922_19591.n223 a_35922_19591.n214 0.809892
R49706 a_35922_19591.n229 a_35922_19591.n128 0.809892
R49707 a_35922_19591.n26 a_35922_19591.n139 1.14908
R49708 a_35922_19591.n93 a_35922_19591.n30 1.14908
R49709 a_35922_19591.n6 a_35922_19591.n21 1.14908
R49710 a_35922_19591.n24 a_35922_19591.n211 1.14908
R49711 a_35922_19591.n207 a_35922_19591.n206 0.71825
R49712 a_35922_19591.n175 a_35922_19591.n164 0.71825
R49713 a_35922_19591.n224 a_35922_19591.n1 1.69988
R49714 a_35922_19591.n228 a_35922_19591.n227 0.673132
R49715 a_35922_19591.n2 a_35922_19591.n228 0.673132
R49716 a_35922_19591.n162 a_35922_19591.n161 0.673132
R49717 a_35922_19591.n27 a_35922_19591.n162 0.673132
R49718 a_35922_19591.n160 a_35922_19591.n159 0.673132
R49719 a_35922_19591.n25 a_35922_19591.n160 0.673132
R49720 a_35922_19591.n179 a_35922_19591.n178 0.673132
R49721 a_35922_19591.n178 a_35922_19591.n177 0.673132
R49722 a_35922_19591.n152 a_35922_19591.n151 0.673132
R49723 a_35922_19591.n153 a_35922_19591.n152 0.673132
R49724 a_35922_19591.n9 a_35922_19591.n213 0.673132
R49725 a_35922_19591.n213 a_35922_19591.n212 0.673132
R49726 a_35922_19591.n210 a_35922_19591.n209 0.673132
R49727 a_35922_19591.n19 a_35922_19591.n210 0.673132
R49728 a_35922_19591.n230 a_35922_19591.n127 0.602344
R49729 a_35922_19591.n221 a_35922_19591.n215 0.571818
R49730 a_35922_19591.n219 a_35922_19591.n218 0.571818
R49731 a_35922_19591.n59 a_35922_19591.n234 0.487111
R49732 a_35922_19591.n61 a_35922_19591.n236 0.487111
R49733 a_35922_19591.n60 a_35922_19591.n233 0.487111
R49734 a_35922_19591.n62 a_35922_19591.n235 0.487111
R49735 a_35922_19591.n109 a_35922_19591.n108 0.321834
R49736 a_35922_19591.n102 a_35922_19591.n134 0.379447
R49737 a_35922_19591.n104 a_35922_19591.n137 0.379447
R49738 a_35922_19591.n172 a_35922_19591.n171 0.379447
R49739 a_35922_19591.n168 a_35922_19591.n167 0.379447
R49740 a_35922_19591.n193 a_35922_19591.n192 0.379447
R49741 a_35922_19591.n188 a_35922_19591.n187 0.379447
R49742 a_35922_19591.n184 a_35922_19591.n183 0.379447
R49743 a_35922_19591.n114 a_35922_19591.n116 0.379447
R49744 a_35922_19591.n117 a_35922_19591.n201 0.379447
R49745 a_35922_19591.n197 a_35922_19591.n196 0.379447
R49746 a_35922_19591.n123 a_35922_19591.n141 0.379447
R49747 a_35922_19591.n146 a_35922_19591.n125 0.379447
R49748 a_35922_19591.n26 a_35922_19591.n18 1.14166
R49749 a_35922_19591.n93 a_35922_19591.n13 2.75347
R49750 a_35922_19591.n100 a_35922_19591.n30 1.60203
R49751 a_35922_19591.n15 a_35922_19591.n21 1.14166
R49752 a_35922_19591.n211 a_35922_19591.n11 2.75347
R49753 a_35922_19591.n101 a_35922_19591.n24 1.60203
R49754 a_35922_19591.n145 a_35922_19591.n144 0.3605
R49755 a_35922_19591.n148 a_35922_19591.n147 0.3605
R49756 a_35922_19591.n204 a_35922_19591.n203 0.3605
R49757 a_35922_19591.n200 a_35922_19591.n154 0.3605
R49758 a_35922_19591.n198 a_35922_19591.n155 0.3605
R49759 a_35922_19591.n191 a_35922_19591.n156 0.3605
R49760 a_35922_19591.n189 a_35922_19591.n157 0.3605
R49761 a_35922_19591.n185 a_35922_19591.n158 0.3605
R49762 a_35922_19591.n173 a_35922_19591.n165 0.3605
R49763 a_35922_19591.n169 a_35922_19591.n166 0.3605
R49764 a_35922_19591.n133 a_35922_19591.n130 0.3605
R49765 a_35922_19591.n136 a_35922_19591.n129 0.3605
R49766 a_35922_19591.n132 a_35922_19591.n131 0.327481
R49767 a_35922_19591.n143 a_35922_19591.n142 0.327481
R49768 a_35922_19591.n195 a_35922_19591.n156 0.208099
R49769 a_35922_19591.n103 a_35922_19591.n102 0.147342
R49770 a_35922_19591.n105 a_35922_19591.n104 0.147342
R49771 a_35922_19591.n176 a_35922_19591.n106 0.147342
R49772 a_35922_19591.n171 a_35922_19591.n107 0.147342
R49773 a_35922_19591.n192 a_35922_19591.n110 0.147342
R49774 a_35922_19591.n187 a_35922_19591.n111 0.147342
R49775 a_35922_19591.n183 a_35922_19591.n112 0.147342
R49776 a_35922_19591.n205 a_35922_19591.n115 0.147342
R49777 a_35922_19591.n118 a_35922_19591.n116 0.147342
R49778 a_35922_19591.n201 a_35922_19591.n119 0.147342
R49779 a_35922_19591.n124 a_35922_19591.n123 0.147342
R49780 a_35922_19591.n126 a_35922_19591.n125 0.147342
R49781 a_35922_19591.n60 a_35922_19591.n232 0.146729
R49782 a_35922_19591.n134 a_35922_19591.n131 0.142605
R49783 a_35922_19591.n194 a_35922_19591.n193 0.142605
R49784 a_35922_19591.n142 a_35922_19591.n141 0.142605
R49785 a_35922_19591.n69 a_35922_19591.n89 2.03311
R49786 a_35922_19591.n35 a_35922_19591.n69 2.04491
R49787 a_35922_19591.n32 a_35922_19591.n35 4.37762
R49788 a_35922_19591.n71 a_35922_19591.n32 1.87961
R49789 a_35922_19591.n71 a_35922_19591.n73 2.19836
R49790 a_35922_19591.n81 a_35922_19591.n98 2.03667
R49791 a_35922_19591.n51 a_35922_19591.n81 2.2172
R49792 a_35922_19591.n51 a_35922_19591.n49 4.49278
R49793 a_35922_19591.n83 a_35922_19591.n49 1.82125
R49794 a_35922_19591.n83 a_35922_19591.n87 2.19319
R49795 a_35922_19591.n98 a_35922_19591.n97 1.65342
R49796 a_35922_19591.n47 a_35922_19591.n46 4.34534
R49797 a_35922_19591.n47 a_35922_19591.n45 1.50598
R49798 a_35922_19591.n65 a_35922_19591.n92 2.03311
R49799 a_35922_19591.n44 a_35922_19591.n65 2.04491
R49800 a_35922_19591.n40 a_35922_19591.n44 4.37762
R49801 a_35922_19591.n67 a_35922_19591.n40 1.87961
R49802 a_35922_19591.n75 a_35922_19591.n67 2.19836
R49803 a_35922_19591.n41 a_35922_19591.n92 1.65903
R49804 a_35922_19591.n42 a_35922_19591.n38 4.49309
R49805 a_35922_19591.n38 a_35922_19591.n37 1.44546
R49806 a_35922_19591.n77 a_35922_19591.n95 2.03657
R49807 a_35922_19591.n77 a_35922_19591.n57 2.21715
R49808 a_35922_19591.n55 a_35922_19591.n57 4.49317
R49809 a_35922_19591.n79 a_35922_19591.n55 1.82113
R49810 a_35922_19591.n85 a_35922_19591.n79 2.19319
R49811 a_35922_19591.n96 a_35922_19591.n95 1.65366
R49812 a_35922_19591.n53 a_35922_19591.n58 4.34574
R49813 a_35922_19591.n53 a_35922_19591.n52 1.50586
R49814 a_35922_19591.n196 a_35922_19591.n120 0.152079
R49815 a_35922_19591.n150 a_35922_19591.n126 0.147342
R49816 a_35922_19591.n146 a_35922_19591.n124 0.147342
R49817 a_35922_19591.n89 a_35922_19591.n88 1.65903
R49818 a_35922_19591.n36 a_35922_19591.n33 4.49309
R49819 a_35922_19591.n33 a_35922_19591.n220 1.44546
R49820 a_35922_19591.n139 a_35922_19591.n5 2.8103
R49821 a_35922_19591.n13 a_35922_19591.n18 4.38327
R49822 a_35922_19591.n145 a_35922_19591.n122 0.14
R49823 a_35922_19591.n147 a_35922_19591.n122 0.14
R49824 a_35922_19591.n149 a_35922_19591.n148 0.14
R49825 a_35922_19591.n149 a_35922_19591.n140 0.14
R49826 a_35922_19591.n206 a_35922_19591.n113 0.14
R49827 a_35922_19591.n204 a_35922_19591.n113 0.14
R49828 a_35922_19591.n203 a_35922_19591.n202 0.14
R49829 a_35922_19591.n202 a_35922_19591.n154 0.14
R49830 a_35922_19591.n200 a_35922_19591.n199 0.14
R49831 a_35922_19591.n199 a_35922_19591.n198 0.14
R49832 a_35922_19591.n121 a_35922_19591.n155 0.208134
R49833 a_35922_19591.n121 a_35922_19591.n195 3.10882
R49834 a_35922_19591.n167 a_35922_19591.n108 0.152079
R49835 a_35922_19591.n197 a_35922_19591.n119 0.147342
R49836 a_35922_19591.n118 a_35922_19591.n117 0.147342
R49837 a_35922_19591.n115 a_35922_19591.n114 0.147342
R49838 a_35922_19591.n180 a_35922_19591.n112 0.147342
R49839 a_35922_19591.n184 a_35922_19591.n111 0.147342
R49840 a_35922_19591.n188 a_35922_19591.n110 0.147342
R49841 a_35922_19591.n191 a_35922_19591.n190 0.14
R49842 a_35922_19591.n190 a_35922_19591.n189 0.14
R49843 a_35922_19591.n186 a_35922_19591.n157 0.14
R49844 a_35922_19591.n186 a_35922_19591.n185 0.14
R49845 a_35922_19591.n182 a_35922_19591.n158 0.14
R49846 a_35922_19591.n182 a_35922_19591.n181 0.14
R49847 a_35922_19591.n175 a_35922_19591.n174 0.14
R49848 a_35922_19591.n174 a_35922_19591.n173 0.14
R49849 a_35922_19591.n170 a_35922_19591.n165 0.14
R49850 a_35922_19591.n170 a_35922_19591.n169 0.14
R49851 a_35922_19591.n109 a_35922_19591.n166 1.12757
R49852 a_35922_19591.n168 a_35922_19591.n107 0.147342
R49853 a_35922_19591.n172 a_35922_19591.n106 0.147342
R49854 a_35922_19591.n226 a_35922_19591.n105 0.147342
R49855 a_35922_19591.n137 a_35922_19591.n103 0.147342
R49856 a_35922_19591.n7 a_35922_19591.n6 2.8103
R49857 a_35922_19591.n15 a_35922_19591.n11 4.38327
R49858 a_35922_19591.n135 a_35922_19591.n130 0.14
R49859 a_35922_19591.n136 a_35922_19591.n135 0.14
R49860 a_35922_19591.n138 a_35922_19591.n129 0.14
R49861 a_35922_19591.n225 a_35922_19591.n138 0.14
R49862 a_35922_19591.n0 a_35922_19591.n1 5.18575
R49863 a_35922_19591.n161 a_35922_19591.n12 2.13563
R49864 a_35922_19591.n10 a_35922_19591.n9 2.13563
R49865 a_35922_19591.n17 a_35922_19591.n16 2.13445
R49866 a_35922_19591.n20 a_35922_19591.n14 2.13445
R49867 a_35922_19591.n63 a_35922_19591.n61 1.89911
R49868 a_35922_19591.n29 a_35922_19591.n28 1.36353
R49869 a_35922_19591.n23 a_35922_19591.n22 1.36353
R49870 a_35922_19591.n0 a_35922_19591.t139 8.54486
R49871 a_35922_19591.n229 a_35922_19591.n0 3.64386
R49872 a_52635_48695.n83 a_52635_48695.n81 7.22198
R49873 a_52635_48695.n119 a_52635_48695.n118 7.22198
R49874 a_52635_48695.n68 a_52635_48695.t125 6.77653
R49875 a_52635_48695.n54 a_52635_48695.t161 6.77653
R49876 a_52635_48695.n60 a_52635_48695.t142 6.7761
R49877 a_52635_48695.n58 a_52635_48695.t92 6.7761
R49878 a_52635_48695.n23 a_52635_48695.t102 6.77231
R49879 a_52635_48695.n33 a_52635_48695.t130 6.77231
R49880 a_52635_48695.n192 a_52635_48695.n191 6.50088
R49881 a_52635_48695.n162 a_52635_48695.n161 6.50088
R49882 a_52635_48695.n72 a_52635_48695.t135 5.50607
R49883 a_52635_48695.n69 a_52635_48695.t99 5.50607
R49884 a_52635_48695.n99 a_52635_48695.t174 5.50607
R49885 a_52635_48695.n55 a_52635_48695.t144 5.50607
R49886 a_52635_48695.n71 a_52635_48695.t138 5.50475
R49887 a_52635_48695.n75 a_52635_48695.t123 5.50475
R49888 a_52635_48695.n76 a_52635_48695.t131 5.50475
R49889 a_52635_48695.n70 a_52635_48695.t127 5.50475
R49890 a_52635_48695.n98 a_52635_48695.t175 5.50475
R49891 a_52635_48695.n102 a_52635_48695.t157 5.50475
R49892 a_52635_48695.n103 a_52635_48695.t170 5.50475
R49893 a_52635_48695.n56 a_52635_48695.t165 5.50475
R49894 a_52635_48695.n137 a_52635_48695.n135 4.92758
R49895 a_52635_48695.n38 a_52635_48695.n36 4.92758
R49896 a_52635_48695.n6 a_52635_48695.n175 4.92217
R49897 a_52635_48695.n13 a_52635_48695.n142 4.92217
R49898 a_52635_48695.n183 a_52635_48695.n0 3.65107
R49899 a_52635_48695.n182 a_52635_48695.n1 3.65107
R49900 a_52635_48695.n181 a_52635_48695.n2 3.65107
R49901 a_52635_48695.n180 a_52635_48695.n3 3.65107
R49902 a_52635_48695.n178 a_52635_48695.n4 3.65107
R49903 a_52635_48695.n177 a_52635_48695.n5 3.65107
R49904 a_52635_48695.n176 a_52635_48695.n6 3.65107
R49905 a_52635_48695.n7 a_52635_48695.n149 3.65107
R49906 a_52635_48695.n8 a_52635_48695.n148 3.65107
R49907 a_52635_48695.n9 a_52635_48695.n147 3.65107
R49908 a_52635_48695.n10 a_52635_48695.n146 3.65107
R49909 a_52635_48695.n145 a_52635_48695.n11 3.65107
R49910 a_52635_48695.n144 a_52635_48695.n12 3.65107
R49911 a_52635_48695.n143 a_52635_48695.n13 3.65107
R49912 a_52635_48695.n14 a_52635_48695.n125 4.0312
R49913 a_52635_48695.t119 a_52635_48695.n15 5.5012
R49914 a_52635_48695.t116 a_52635_48695.n16 5.5012
R49915 a_52635_48695.n124 a_52635_48695.n17 4.0312
R49916 a_52635_48695.t98 a_52635_48695.n18 5.5012
R49917 a_52635_48695.t111 a_52635_48695.n19 5.5012
R49918 a_52635_48695.n123 a_52635_48695.n20 4.0312
R49919 a_52635_48695.t108 a_52635_48695.n21 5.5012
R49920 a_52635_48695.t88 a_52635_48695.n22 5.5012
R49921 a_52635_48695.n51 a_52635_48695.n23 4.0312
R49922 a_52635_48695.n24 a_52635_48695.n93 4.0312
R49923 a_52635_48695.t147 a_52635_48695.n25 5.5012
R49924 a_52635_48695.t145 a_52635_48695.n26 5.5012
R49925 a_52635_48695.n92 a_52635_48695.n27 4.0312
R49926 a_52635_48695.t126 a_52635_48695.n28 5.5012
R49927 a_52635_48695.t139 a_52635_48695.n29 5.5012
R49928 a_52635_48695.n91 a_52635_48695.n30 4.0312
R49929 a_52635_48695.t136 a_52635_48695.n31 5.5012
R49930 a_52635_48695.t110 a_52635_48695.n32 5.5012
R49931 a_52635_48695.n89 a_52635_48695.n33 4.0312
R49932 a_52635_48695.n82 a_52635_48695.t128 4.24002
R49933 a_52635_48695.n62 a_52635_48695.t95 4.24002
R49934 a_52635_48695.n117 a_52635_48695.t100 4.24002
R49935 a_52635_48695.n108 a_52635_48695.t163 4.24002
R49936 a_52635_48695.n156 a_52635_48695.t71 4.06712
R49937 a_52635_48695.n154 a_52635_48695.t62 4.06712
R49938 a_52635_48695.n186 a_52635_48695.t79 4.06712
R49939 a_52635_48695.n48 a_52635_48695.t66 4.06712
R49940 a_52635_48695.n60 a_52635_48695.n59 4.03475
R49941 a_52635_48695.n74 a_52635_48695.n73 4.03475
R49942 a_52635_48695.n78 a_52635_48695.n77 4.03475
R49943 a_52635_48695.n68 a_52635_48695.n67 4.03475
R49944 a_52635_48695.n58 a_52635_48695.n57 4.03475
R49945 a_52635_48695.n101 a_52635_48695.n100 4.03475
R49946 a_52635_48695.n105 a_52635_48695.n104 4.03475
R49947 a_52635_48695.n54 a_52635_48695.n53 4.03475
R49948 a_52635_48695.n128 a_52635_48695.n43 3.97307
R49949 a_52635_48695.n187 a_52635_48695.n185 3.96014
R49950 a_52635_48695.n157 a_52635_48695.n134 3.96014
R49951 a_52635_48695.n156 a_52635_48695.t74 3.86107
R49952 a_52635_48695.n154 a_52635_48695.t63 3.86107
R49953 a_52635_48695.n186 a_52635_48695.t0 3.86107
R49954 a_52635_48695.n48 a_52635_48695.t75 3.86107
R49955 a_52635_48695.n139 a_52635_48695.n137 3.79678
R49956 a_52635_48695.n171 a_52635_48695.n169 3.79678
R49957 a_52635_48695.n40 a_52635_48695.n38 3.79678
R49958 a_52635_48695.n130 a_52635_48695.n35 3.79678
R49959 a_52635_48695.n82 a_52635_48695.t106 3.68818
R49960 a_52635_48695.n62 a_52635_48695.t166 3.68818
R49961 a_52635_48695.n117 a_52635_48695.t148 3.68818
R49962 a_52635_48695.n108 a_52635_48695.t114 3.68818
R49963 a_52635_48695.n132 a_52635_48695.n131 3.65581
R49964 a_52635_48695.n173 a_52635_48695.n172 3.65581
R49965 a_52635_48695.n171 a_52635_48695.n170 3.65581
R49966 a_52635_48695.n169 a_52635_48695.n168 3.65581
R49967 a_52635_48695.n167 a_52635_48695.n166 3.65581
R49968 a_52635_48695.n141 a_52635_48695.n140 3.65581
R49969 a_52635_48695.n139 a_52635_48695.n138 3.65581
R49970 a_52635_48695.n137 a_52635_48695.n136 3.65581
R49971 a_52635_48695.n130 a_52635_48695.n129 3.65581
R49972 a_52635_48695.n35 a_52635_48695.n34 3.65581
R49973 a_52635_48695.n197 a_52635_48695.n196 3.65581
R49974 a_52635_48695.n42 a_52635_48695.n41 3.65581
R49975 a_52635_48695.n40 a_52635_48695.n39 3.65581
R49976 a_52635_48695.n38 a_52635_48695.n37 3.65581
R49977 a_52635_48695.n167 a_52635_48695.n165 3.64443
R49978 a_52635_48695.n196 a_52635_48695.n195 3.64443
R49979 a_52635_48695.n3 a_52635_48695.n179 3.64223
R49980 a_52635_48695.n150 a_52635_48695.n10 3.64223
R49981 a_52635_48695.n88 a_52635_48695.n87 3.23904
R49982 a_52635_48695.n116 a_52635_48695.n50 3.23904
R49983 a_52635_48695.n86 a_52635_48695.n85 2.77002
R49984 a_52635_48695.n65 a_52635_48695.n64 2.77002
R49985 a_52635_48695.n115 a_52635_48695.n114 2.77002
R49986 a_52635_48695.n111 a_52635_48695.n110 2.77002
R49987 a_52635_48695.n66 a_52635_48695.n62 2.73714
R49988 a_52635_48695.n112 a_52635_48695.n108 2.73714
R49989 a_52635_48695.n49 a_52635_48695.n47 2.73714
R49990 a_52635_48695.n155 a_52635_48695.n153 2.73714
R49991 a_52635_48695.n76 a_52635_48695.n75 2.60203
R49992 a_52635_48695.n103 a_52635_48695.n102 2.60203
R49993 a_52635_48695.n160 a_52635_48695.n158 2.59712
R49994 a_52635_48695.n153 a_52635_48695.n151 2.59712
R49995 a_52635_48695.n190 a_52635_48695.n188 2.59712
R49996 a_52635_48695.n47 a_52635_48695.n45 2.59712
R49997 a_52635_48695.n70 a_52635_48695.n69 2.52436
R49998 a_52635_48695.n72 a_52635_48695.n71 2.52436
R49999 a_52635_48695.n56 a_52635_48695.n55 2.52436
R50000 a_52635_48695.n99 a_52635_48695.n98 2.52436
R50001 a_52635_48695.n192 a_52635_48695.n49 2.46014
R50002 a_52635_48695.n162 a_52635_48695.n155 2.46014
R50003 a_52635_48695.n160 a_52635_48695.n159 2.39107
R50004 a_52635_48695.n153 a_52635_48695.n152 2.39107
R50005 a_52635_48695.n190 a_52635_48695.n189 2.39107
R50006 a_52635_48695.n47 a_52635_48695.n46 2.39107
R50007 a_52635_48695.n86 a_52635_48695.n84 2.21818
R50008 a_52635_48695.n65 a_52635_48695.n63 2.21818
R50009 a_52635_48695.n115 a_52635_48695.n113 2.21818
R50010 a_52635_48695.n111 a_52635_48695.n109 2.21818
R50011 a_52635_48695.n80 a_52635_48695.n79 2.13841
R50012 a_52635_48695.n88 a_52635_48695.n61 2.13841
R50013 a_52635_48695.n163 a_52635_48695.n150 2.0852
R50014 a_52635_48695.n133 a_52635_48695.n128 2.02864
R50015 a_52635_48695.n121 a_52635_48695.n43 1.76168
R50016 a_52635_48695.n81 a_52635_48695.n66 1.73904
R50017 a_52635_48695.n119 a_52635_48695.n112 1.73904
R50018 a_52635_48695.n174 a_52635_48695.n173 1.73609
R50019 a_52635_48695.n133 a_52635_48695.n132 1.73609
R50020 a_52635_48695.n120 a_52635_48695.n119 1.5005
R50021 a_52635_48695.n107 a_52635_48695.n106 1.5005
R50022 a_52635_48695.n90 a_52635_48695.n52 1.5005
R50023 a_52635_48695.n81 a_52635_48695.n80 1.5005
R50024 a_52635_48695.n122 a_52635_48695.n121 1.5005
R50025 a_52635_48695.n127 a_52635_48695.n126 1.5005
R50026 a_52635_48695.n97 a_52635_48695.n96 1.5005
R50027 a_52635_48695.n95 a_52635_48695.n94 1.5005
R50028 a_52635_48695.n163 a_52635_48695.n162 1.5005
R50029 a_52635_48695.n193 a_52635_48695.n192 1.5005
R50030 a_52635_48695.n165 a_52635_48695.n164 1.5005
R50031 a_52635_48695.n179 a_52635_48695.n44 1.5005
R50032 a_52635_48695.n195 a_52635_48695.n194 1.5005
R50033 a_52635_48695.n131 a_52635_48695.t46 1.4705
R50034 a_52635_48695.n131 a_52635_48695.t21 1.4705
R50035 a_52635_48695.n158 a_52635_48695.t57 1.4705
R50036 a_52635_48695.n158 a_52635_48695.t37 1.4705
R50037 a_52635_48695.n159 a_52635_48695.t59 1.4705
R50038 a_52635_48695.n159 a_52635_48695.t40 1.4705
R50039 a_52635_48695.n151 a_52635_48695.t36 1.4705
R50040 a_52635_48695.n151 a_52635_48695.t29 1.4705
R50041 a_52635_48695.n152 a_52635_48695.t38 1.4705
R50042 a_52635_48695.n152 a_52635_48695.t30 1.4705
R50043 a_52635_48695.n183 a_52635_48695.t33 1.4705
R50044 a_52635_48695.n183 a_52635_48695.t10 1.4705
R50045 a_52635_48695.n182 a_52635_48695.t5 1.4705
R50046 a_52635_48695.n182 a_52635_48695.t51 1.4705
R50047 a_52635_48695.n181 a_52635_48695.t86 1.4705
R50048 a_52635_48695.n181 a_52635_48695.t4 1.4705
R50049 a_52635_48695.n180 a_52635_48695.t67 1.4705
R50050 a_52635_48695.n180 a_52635_48695.t27 1.4705
R50051 a_52635_48695.n178 a_52635_48695.t8 1.4705
R50052 a_52635_48695.n178 a_52635_48695.t85 1.4705
R50053 a_52635_48695.n177 a_52635_48695.t80 1.4705
R50054 a_52635_48695.n177 a_52635_48695.t32 1.4705
R50055 a_52635_48695.n176 a_52635_48695.t72 1.4705
R50056 a_52635_48695.n176 a_52635_48695.t52 1.4705
R50057 a_52635_48695.n175 a_52635_48695.t73 1.4705
R50058 a_52635_48695.n175 a_52635_48695.t23 1.4705
R50059 a_52635_48695.n172 a_52635_48695.t41 1.4705
R50060 a_52635_48695.n172 a_52635_48695.t18 1.4705
R50061 a_52635_48695.n170 a_52635_48695.t14 1.4705
R50062 a_52635_48695.n170 a_52635_48695.t53 1.4705
R50063 a_52635_48695.n168 a_52635_48695.t7 1.4705
R50064 a_52635_48695.n168 a_52635_48695.t11 1.4705
R50065 a_52635_48695.n166 a_52635_48695.t77 1.4705
R50066 a_52635_48695.n166 a_52635_48695.t31 1.4705
R50067 a_52635_48695.n140 a_52635_48695.t15 1.4705
R50068 a_52635_48695.n140 a_52635_48695.t6 1.4705
R50069 a_52635_48695.n138 a_52635_48695.t3 1.4705
R50070 a_52635_48695.n138 a_52635_48695.t39 1.4705
R50071 a_52635_48695.n136 a_52635_48695.t81 1.4705
R50072 a_52635_48695.n136 a_52635_48695.t55 1.4705
R50073 a_52635_48695.n135 a_52635_48695.t82 1.4705
R50074 a_52635_48695.n135 a_52635_48695.t24 1.4705
R50075 a_52635_48695.n149 a_52635_48695.t26 1.4705
R50076 a_52635_48695.n149 a_52635_48695.t84 1.4705
R50077 a_52635_48695.n148 a_52635_48695.t78 1.4705
R50078 a_52635_48695.n148 a_52635_48695.t47 1.4705
R50079 a_52635_48695.n147 a_52635_48695.t69 1.4705
R50080 a_52635_48695.n147 a_52635_48695.t76 1.4705
R50081 a_52635_48695.n146 a_52635_48695.t56 1.4705
R50082 a_52635_48695.n146 a_52635_48695.t22 1.4705
R50083 a_52635_48695.n145 a_52635_48695.t83 1.4705
R50084 a_52635_48695.n145 a_52635_48695.t68 1.4705
R50085 a_52635_48695.n144 a_52635_48695.t65 1.4705
R50086 a_52635_48695.n144 a_52635_48695.t25 1.4705
R50087 a_52635_48695.n143 a_52635_48695.t60 1.4705
R50088 a_52635_48695.n143 a_52635_48695.t50 1.4705
R50089 a_52635_48695.n142 a_52635_48695.t61 1.4705
R50090 a_52635_48695.n142 a_52635_48695.t16 1.4705
R50091 a_52635_48695.n125 a_52635_48695.t173 1.4705
R50092 a_52635_48695.n125 a_52635_48695.t153 1.4705
R50093 a_52635_48695.n124 a_52635_48695.t146 1.4705
R50094 a_52635_48695.n124 a_52635_48695.t112 1.4705
R50095 a_52635_48695.n123 a_52635_48695.t152 1.4705
R50096 a_52635_48695.n123 a_52635_48695.t121 1.4705
R50097 a_52635_48695.n51 a_52635_48695.t134 1.4705
R50098 a_52635_48695.n51 a_52635_48695.t101 1.4705
R50099 a_52635_48695.n59 a_52635_48695.t94 1.4705
R50100 a_52635_48695.n59 a_52635_48695.t172 1.4705
R50101 a_52635_48695.n73 a_52635_48695.t162 1.4705
R50102 a_52635_48695.n73 a_52635_48695.t132 1.4705
R50103 a_52635_48695.n77 a_52635_48695.t169 1.4705
R50104 a_52635_48695.n77 a_52635_48695.t141 1.4705
R50105 a_52635_48695.n67 a_52635_48695.t154 1.4705
R50106 a_52635_48695.n67 a_52635_48695.t124 1.4705
R50107 a_52635_48695.n84 a_52635_48695.t167 1.4705
R50108 a_52635_48695.n84 a_52635_48695.t120 1.4705
R50109 a_52635_48695.n85 a_52635_48695.t96 1.4705
R50110 a_52635_48695.n85 a_52635_48695.t143 1.4705
R50111 a_52635_48695.n63 a_52635_48695.t158 1.4705
R50112 a_52635_48695.n63 a_52635_48695.t109 1.4705
R50113 a_52635_48695.n64 a_52635_48695.t93 1.4705
R50114 a_52635_48695.n64 a_52635_48695.t133 1.4705
R50115 a_52635_48695.n93 a_52635_48695.t103 1.4705
R50116 a_52635_48695.n93 a_52635_48695.t91 1.4705
R50117 a_52635_48695.n92 a_52635_48695.t168 1.4705
R50118 a_52635_48695.n92 a_52635_48695.t140 1.4705
R50119 a_52635_48695.n91 a_52635_48695.t89 1.4705
R50120 a_52635_48695.n91 a_52635_48695.t149 1.4705
R50121 a_52635_48695.n89 a_52635_48695.t159 1.4705
R50122 a_52635_48695.n89 a_52635_48695.t129 1.4705
R50123 a_52635_48695.n57 a_52635_48695.t137 1.4705
R50124 a_52635_48695.n57 a_52635_48695.t118 1.4705
R50125 a_52635_48695.n100 a_52635_48695.t107 1.4705
R50126 a_52635_48695.n100 a_52635_48695.t171 1.4705
R50127 a_52635_48695.n104 a_52635_48695.t117 1.4705
R50128 a_52635_48695.n104 a_52635_48695.t90 1.4705
R50129 a_52635_48695.n53 a_52635_48695.t97 1.4705
R50130 a_52635_48695.n53 a_52635_48695.t160 1.4705
R50131 a_52635_48695.n113 a_52635_48695.t115 1.4705
R50132 a_52635_48695.n113 a_52635_48695.t155 1.4705
R50133 a_52635_48695.n114 a_52635_48695.t164 1.4705
R50134 a_52635_48695.n114 a_52635_48695.t113 1.4705
R50135 a_52635_48695.n109 a_52635_48695.t105 1.4705
R50136 a_52635_48695.n109 a_52635_48695.t151 1.4705
R50137 a_52635_48695.n110 a_52635_48695.t156 1.4705
R50138 a_52635_48695.n110 a_52635_48695.t104 1.4705
R50139 a_52635_48695.n188 a_52635_48695.t64 1.4705
R50140 a_52635_48695.n188 a_52635_48695.t44 1.4705
R50141 a_52635_48695.n189 a_52635_48695.t70 1.4705
R50142 a_52635_48695.n189 a_52635_48695.t49 1.4705
R50143 a_52635_48695.n45 a_52635_48695.t43 1.4705
R50144 a_52635_48695.n45 a_52635_48695.t34 1.4705
R50145 a_52635_48695.n46 a_52635_48695.t48 1.4705
R50146 a_52635_48695.n46 a_52635_48695.t42 1.4705
R50147 a_52635_48695.n129 a_52635_48695.t19 1.4705
R50148 a_52635_48695.n129 a_52635_48695.t54 1.4705
R50149 a_52635_48695.n34 a_52635_48695.t13 1.4705
R50150 a_52635_48695.n34 a_52635_48695.t17 1.4705
R50151 a_52635_48695.n41 a_52635_48695.t20 1.4705
R50152 a_52635_48695.n41 a_52635_48695.t12 1.4705
R50153 a_52635_48695.n39 a_52635_48695.t9 1.4705
R50154 a_52635_48695.n39 a_52635_48695.t45 1.4705
R50155 a_52635_48695.n37 a_52635_48695.t1 1.4705
R50156 a_52635_48695.n37 a_52635_48695.t58 1.4705
R50157 a_52635_48695.n36 a_52635_48695.t2 1.4705
R50158 a_52635_48695.n36 a_52635_48695.t28 1.4705
R50159 a_52635_48695.t87 a_52635_48695.n197 1.4705
R50160 a_52635_48695.n197 a_52635_48695.t35 1.4705
R50161 a_52635_48695.n87 a_52635_48695.n86 1.46537
R50162 a_52635_48695.n83 a_52635_48695.n82 1.46537
R50163 a_52635_48695.n66 a_52635_48695.n65 1.46537
R50164 a_52635_48695.n116 a_52635_48695.n115 1.46537
R50165 a_52635_48695.n118 a_52635_48695.n117 1.46537
R50166 a_52635_48695.n112 a_52635_48695.n111 1.46537
R50167 a_52635_48695.n157 a_52635_48695.n156 1.46537
R50168 a_52635_48695.n161 a_52635_48695.n160 1.46537
R50169 a_52635_48695.n155 a_52635_48695.n154 1.46537
R50170 a_52635_48695.n187 a_52635_48695.n186 1.46537
R50171 a_52635_48695.n191 a_52635_48695.n190 1.46537
R50172 a_52635_48695.n49 a_52635_48695.n48 1.46537
R50173 a_52635_48695.n194 a_52635_48695.n43 1.42428
R50174 a_52635_48695.n78 a_52635_48695.n76 1.27228
R50175 a_52635_48695.n75 a_52635_48695.n74 1.27228
R50176 a_52635_48695.n87 a_52635_48695.n83 1.27228
R50177 a_52635_48695.n105 a_52635_48695.n103 1.27228
R50178 a_52635_48695.n102 a_52635_48695.n101 1.27228
R50179 a_52635_48695.n118 a_52635_48695.n116 1.27228
R50180 a_52635_48695.n141 a_52635_48695.n139 1.27228
R50181 a_52635_48695.n169 a_52635_48695.n167 1.27228
R50182 a_52635_48695.n173 a_52635_48695.n171 1.27228
R50183 a_52635_48695.n191 a_52635_48695.n187 1.27228
R50184 a_52635_48695.n161 a_52635_48695.n157 1.27228
R50185 a_52635_48695.n196 a_52635_48695.n35 1.27228
R50186 a_52635_48695.n42 a_52635_48695.n40 1.27228
R50187 a_52635_48695.n132 a_52635_48695.n130 1.27228
R50188 a_52635_48695.n69 a_52635_48695.n68 1.26756
R50189 a_52635_48695.n74 a_52635_48695.n72 1.26756
R50190 a_52635_48695.n55 a_52635_48695.n54 1.26756
R50191 a_52635_48695.n101 a_52635_48695.n99 1.26756
R50192 a_52635_48695.n128 a_52635_48695.n127 1.15732
R50193 a_52635_48695.n184 a_52635_48695.n174 0.822966
R50194 a_52635_48695.n164 a_52635_48695.n44 0.822966
R50195 a_52635_48695.n79 a_52635_48695.n70 0.796291
R50196 a_52635_48695.n71 a_52635_48695.n61 0.796291
R50197 a_52635_48695.n106 a_52635_48695.n56 0.796291
R50198 a_52635_48695.n98 a_52635_48695.n97 0.796291
R50199 a_52635_48695.n80 a_52635_48695.n52 0.780703
R50200 a_52635_48695.n121 a_52635_48695.n120 0.780703
R50201 a_52635_48695.n95 a_52635_48695.n88 0.780703
R50202 a_52635_48695.n127 a_52635_48695.n50 0.780703
R50203 a_52635_48695.n185 a_52635_48695.n133 0.639318
R50204 a_52635_48695.n174 a_52635_48695.n134 0.639318
R50205 a_52635_48695.n194 a_52635_48695.n193 0.639318
R50206 a_52635_48695.n164 a_52635_48695.n163 0.639318
R50207 a_52635_48695.n120 a_52635_48695.n107 0.638405
R50208 a_52635_48695.n96 a_52635_48695.n50 0.638405
R50209 a_52635_48695.n107 a_52635_48695.n52 0.628372
R50210 a_52635_48695.n96 a_52635_48695.n95 0.628372
R50211 a_52635_48695.n185 a_52635_48695.n184 0.585196
R50212 a_52635_48695.n193 a_52635_48695.n44 0.585196
R50213 a_52635_48695.n79 a_52635_48695.n78 0.476484
R50214 a_52635_48695.n61 a_52635_48695.n60 0.476484
R50215 a_52635_48695.n106 a_52635_48695.n105 0.476484
R50216 a_52635_48695.n97 a_52635_48695.n58 0.476484
R50217 a_52635_48695.n30 a_52635_48695.n90 0.478684
R50218 a_52635_48695.n94 a_52635_48695.n24 0.478684
R50219 a_52635_48695.n20 a_52635_48695.n122 0.478684
R50220 a_52635_48695.n126 a_52635_48695.n14 0.478684
R50221 a_52635_48695.n165 a_52635_48695.n141 0.236091
R50222 a_52635_48695.n195 a_52635_48695.n42 0.236091
R50223 a_52635_48695.n5 a_52635_48695.n6 3.79678
R50224 a_52635_48695.n4 a_52635_48695.n5 1.27228
R50225 a_52635_48695.n179 a_52635_48695.n4 0.238291
R50226 a_52635_48695.n2 a_52635_48695.n3 1.27228
R50227 a_52635_48695.n1 a_52635_48695.n2 3.79678
R50228 a_52635_48695.n0 a_52635_48695.n1 1.27228
R50229 a_52635_48695.n184 a_52635_48695.n0 1.73829
R50230 a_52635_48695.n12 a_52635_48695.n13 3.79678
R50231 a_52635_48695.n11 a_52635_48695.n12 1.27228
R50232 a_52635_48695.n150 a_52635_48695.n11 0.238291
R50233 a_52635_48695.n9 a_52635_48695.n10 1.27228
R50234 a_52635_48695.n8 a_52635_48695.n9 3.79678
R50235 a_52635_48695.n7 a_52635_48695.n8 1.27228
R50236 a_52635_48695.n134 a_52635_48695.n7 2.32299
R50237 a_52635_48695.n32 a_52635_48695.n33 1.27228
R50238 a_52635_48695.n31 a_52635_48695.n32 2.51878
R50239 a_52635_48695.n90 a_52635_48695.n31 0.794091
R50240 a_52635_48695.n29 a_52635_48695.n30 1.27228
R50241 a_52635_48695.n28 a_52635_48695.n29 2.60203
R50242 a_52635_48695.n27 a_52635_48695.n28 1.27228
R50243 a_52635_48695.n26 a_52635_48695.n27 1.27228
R50244 a_52635_48695.n25 a_52635_48695.n26 2.51878
R50245 a_52635_48695.n94 a_52635_48695.n25 0.794091
R50246 a_52635_48695.t150 a_52635_48695.n24 6.77266
R50247 a_52635_48695.n22 a_52635_48695.n23 1.27228
R50248 a_52635_48695.n21 a_52635_48695.n22 2.51878
R50249 a_52635_48695.n122 a_52635_48695.n21 0.794091
R50250 a_52635_48695.n19 a_52635_48695.n20 1.27228
R50251 a_52635_48695.n18 a_52635_48695.n19 2.60203
R50252 a_52635_48695.n17 a_52635_48695.n18 1.27228
R50253 a_52635_48695.n16 a_52635_48695.n17 1.27228
R50254 a_52635_48695.n15 a_52635_48695.n16 2.51878
R50255 a_52635_48695.n126 a_52635_48695.n15 0.794091
R50256 a_52635_48695.t122 a_52635_48695.n14 6.77266
R50257 a_50751_n19729.n300 a_50751_n19729.t73 12.6064
R50258 a_50751_n19729.t357 a_50751_n19729.n232 10.1674
R50259 a_50751_n19729.n233 a_50751_n19729.t357 10.1674
R50260 a_50751_n19729.t137 a_50751_n19729.n234 10.1674
R50261 a_50751_n19729.n235 a_50751_n19729.t137 10.1674
R50262 a_50751_n19729.t122 a_50751_n19729.n238 10.1674
R50263 a_50751_n19729.n239 a_50751_n19729.t122 10.1674
R50264 a_50751_n19729.t194 a_50751_n19729.n242 10.1674
R50265 a_50751_n19729.n243 a_50751_n19729.t194 10.1674
R50266 a_50751_n19729.t346 a_50751_n19729.n250 10.1674
R50267 a_50751_n19729.n251 a_50751_n19729.t346 10.1674
R50268 a_50751_n19729.n499 a_50751_n19729.t111 10.1674
R50269 a_50751_n19729.t111 a_50751_n19729.n498 10.1674
R50270 a_50751_n19729.n493 a_50751_n19729.t170 10.1674
R50271 a_50751_n19729.n297 a_50751_n19729.t106 10.1674
R50272 a_50751_n19729.t106 a_50751_n19729.n296 10.1674
R50273 a_50751_n19729.n293 a_50751_n19729.t100 10.1674
R50274 a_50751_n19729.t100 a_50751_n19729.n292 10.1674
R50275 a_50751_n19729.n289 a_50751_n19729.t167 10.1674
R50276 a_50751_n19729.t167 a_50751_n19729.n288 10.1674
R50277 a_50751_n19729.t250 a_50751_n19729.n257 10.1674
R50278 a_50751_n19729.n258 a_50751_n19729.t250 10.1674
R50279 a_50751_n19729.t297 a_50751_n19729.n265 10.1674
R50280 a_50751_n19729.n266 a_50751_n19729.t297 10.1674
R50281 a_50751_n19729.n276 a_50751_n19729.t132 10.1674
R50282 a_50751_n19729.t132 a_50751_n19729.n275 10.1674
R50283 a_50751_n19729.n270 a_50751_n19729.t204 10.1674
R50284 a_50751_n19729.n247 a_50751_n19729.t274 10.1674
R50285 a_50751_n19729.t274 a_50751_n19729.n246 10.1674
R50286 a_50751_n19729.t331 a_50751_n19729.n502 10.1674
R50287 a_50751_n19729.n503 a_50751_n19729.t331 10.1674
R50288 a_50751_n19729.t140 a_50751_n19729.n307 10.1674
R50289 a_50751_n19729.n308 a_50751_n19729.t140 10.1674
R50290 a_50751_n19729.t212 a_50751_n19729.n309 10.1674
R50291 a_50751_n19729.n310 a_50751_n19729.t212 10.1674
R50292 a_50751_n19729.t196 a_50751_n19729.n313 10.1674
R50293 a_50751_n19729.n314 a_50751_n19729.t196 10.1674
R50294 a_50751_n19729.n326 a_50751_n19729.t276 10.1674
R50295 a_50751_n19729.t276 a_50751_n19729.n325 10.1674
R50296 a_50751_n19729.n318 a_50751_n19729.t129 10.1674
R50297 a_50751_n19729.t129 a_50751_n19729.n317 10.1674
R50298 a_50751_n19729.t184 a_50751_n19729.n338 10.1674
R50299 a_50751_n19729.n339 a_50751_n19729.t184 10.1674
R50300 a_50751_n19729.n343 a_50751_n19729.t254 10.1674
R50301 a_50751_n19729.n391 a_50751_n19729.t286 10.1674
R50302 a_50751_n19729.t286 a_50751_n19729.n390 10.1674
R50303 a_50751_n19729.n387 a_50751_n19729.t272 10.1674
R50304 a_50751_n19729.t272 a_50751_n19729.n386 10.1674
R50305 a_50751_n19729.n383 a_50751_n19729.t345 10.1674
R50306 a_50751_n19729.t345 a_50751_n19729.n382 10.1674
R50307 a_50751_n19729.t127 a_50751_n19729.n351 10.1674
R50308 a_50751_n19729.n352 a_50751_n19729.t127 10.1674
R50309 a_50751_n19729.t169 a_50751_n19729.n359 10.1674
R50310 a_50751_n19729.n360 a_50751_n19729.t169 10.1674
R50311 a_50751_n19729.n370 a_50751_n19729.t309 10.1674
R50312 a_50751_n19729.t309 a_50751_n19729.n369 10.1674
R50313 a_50751_n19729.n364 a_50751_n19729.t94 10.1674
R50314 a_50751_n19729.t348 a_50751_n19729.n321 10.1674
R50315 a_50751_n19729.n322 a_50751_n19729.t348 10.1674
R50316 a_50751_n19729.n335 a_50751_n19729.t115 10.1674
R50317 a_50751_n19729.t115 a_50751_n19729.n334 10.1674
R50318 a_50751_n19729.n356 a_50751_n19729.t110 10.1674
R50319 a_50751_n19729.t110 a_50751_n19729.n355 10.1674
R50320 a_50751_n19729.t252 a_50751_n19729.n373 10.1674
R50321 a_50751_n19729.n374 a_50751_n19729.t252 10.1674
R50322 a_50751_n19729.t257 a_50751_n19729.n402 10.1674
R50323 a_50751_n19729.n403 a_50751_n19729.t257 10.1674
R50324 a_50751_n19729.t328 a_50751_n19729.n404 10.1674
R50325 a_50751_n19729.n405 a_50751_n19729.t328 10.1674
R50326 a_50751_n19729.t319 a_50751_n19729.n408 10.1674
R50327 a_50751_n19729.n409 a_50751_n19729.t319 10.1674
R50328 a_50751_n19729.n421 a_50751_n19729.t99 10.1674
R50329 a_50751_n19729.t99 a_50751_n19729.n420 10.1674
R50330 a_50751_n19729.n413 a_50751_n19729.t249 10.1674
R50331 a_50751_n19729.t249 a_50751_n19729.n412 10.1674
R50332 a_50751_n19729.t310 a_50751_n19729.n433 10.1674
R50333 a_50751_n19729.n434 a_50751_n19729.t310 10.1674
R50334 a_50751_n19729.n438 a_50751_n19729.t82 10.1674
R50335 a_50751_n19729.n486 a_50751_n19729.t255 10.1674
R50336 a_50751_n19729.t255 a_50751_n19729.n485 10.1674
R50337 a_50751_n19729.n482 a_50751_n19729.t239 10.1674
R50338 a_50751_n19729.t239 a_50751_n19729.n481 10.1674
R50339 a_50751_n19729.n478 a_50751_n19729.t318 10.1674
R50340 a_50751_n19729.t318 a_50751_n19729.n477 10.1674
R50341 a_50751_n19729.t98 a_50751_n19729.n446 10.1674
R50342 a_50751_n19729.n447 a_50751_n19729.t98 10.1674
R50343 a_50751_n19729.t143 a_50751_n19729.n454 10.1674
R50344 a_50751_n19729.n455 a_50751_n19729.t143 10.1674
R50345 a_50751_n19729.n465 a_50751_n19729.t279 10.1674
R50346 a_50751_n19729.t279 a_50751_n19729.n464 10.1674
R50347 a_50751_n19729.n459 a_50751_n19729.t349 10.1674
R50348 a_50751_n19729.t166 a_50751_n19729.n416 10.1674
R50349 a_50751_n19729.n417 a_50751_n19729.t166 10.1674
R50350 a_50751_n19729.n430 a_50751_n19729.t230 10.1674
R50351 a_50751_n19729.t230 a_50751_n19729.n429 10.1674
R50352 a_50751_n19729.n451 a_50751_n19729.t91 10.1674
R50353 a_50751_n19729.t91 a_50751_n19729.n450 10.1674
R50354 a_50751_n19729.t218 a_50751_n19729.n468 10.1674
R50355 a_50751_n19729.n469 a_50751_n19729.t218 10.1674
R50356 a_50751_n19729.n262 a_50751_n19729.t231 10.1674
R50357 a_50751_n19729.t231 a_50751_n19729.n261 10.1674
R50358 a_50751_n19729.t83 a_50751_n19729.n279 10.1674
R50359 a_50751_n19729.n280 a_50751_n19729.t83 10.1674
R50360 a_50751_n19729.n231 a_50751_n19729.t229 10.1674
R50361 a_50751_n19729.t229 a_50751_n19729.n230 10.1674
R50362 a_50751_n19729.t308 a_50751_n19729.n236 10.1674
R50363 a_50751_n19729.n237 a_50751_n19729.t308 10.1674
R50364 a_50751_n19729.t296 a_50751_n19729.n240 10.1674
R50365 a_50751_n19729.n241 a_50751_n19729.t296 10.1674
R50366 a_50751_n19729.t81 a_50751_n19729.n244 10.1674
R50367 a_50751_n19729.n245 a_50751_n19729.t81 10.1674
R50368 a_50751_n19729.t222 a_50751_n19729.n252 10.1674
R50369 a_50751_n19729.n253 a_50751_n19729.t222 10.1674
R50370 a_50751_n19729.n501 a_50751_n19729.t287 10.1674
R50371 a_50751_n19729.t287 a_50751_n19729.n500 10.1674
R50372 a_50751_n19729.n495 a_50751_n19729.t342 10.1674
R50373 a_50751_n19729.n299 a_50751_n19729.t351 10.1674
R50374 a_50751_n19729.t351 a_50751_n19729.n298 10.1674
R50375 a_50751_n19729.n295 a_50751_n19729.t337 10.1674
R50376 a_50751_n19729.t337 a_50751_n19729.n294 10.1674
R50377 a_50751_n19729.n291 a_50751_n19729.t118 10.1674
R50378 a_50751_n19729.t118 a_50751_n19729.n290 10.1674
R50379 a_50751_n19729.t188 a_50751_n19729.n259 10.1674
R50380 a_50751_n19729.n260 a_50751_n19729.t188 10.1674
R50381 a_50751_n19729.t242 a_50751_n19729.n267 10.1674
R50382 a_50751_n19729.n268 a_50751_n19729.t242 10.1674
R50383 a_50751_n19729.n278 a_50751_n19729.t86 10.1674
R50384 a_50751_n19729.t86 a_50751_n19729.n277 10.1674
R50385 a_50751_n19729.n272 a_50751_n19729.t154 10.1674
R50386 a_50751_n19729.n249 a_50751_n19729.t149 10.1674
R50387 a_50751_n19729.t149 a_50751_n19729.n248 10.1674
R50388 a_50751_n19729.t210 a_50751_n19729.n504 10.1674
R50389 a_50751_n19729.n505 a_50751_n19729.t210 10.1674
R50390 a_50751_n19729.n306 a_50751_n19729.t80 10.1674
R50391 a_50751_n19729.t80 a_50751_n19729.n305 10.1674
R50392 a_50751_n19729.t148 a_50751_n19729.n311 10.1674
R50393 a_50751_n19729.n312 a_50751_n19729.t148 10.1674
R50394 a_50751_n19729.t136 a_50751_n19729.n315 10.1674
R50395 a_50751_n19729.n316 a_50751_n19729.t136 10.1674
R50396 a_50751_n19729.n328 a_50751_n19729.t209 10.1674
R50397 a_50751_n19729.t209 a_50751_n19729.n327 10.1674
R50398 a_50751_n19729.n320 a_50751_n19729.t361 10.1674
R50399 a_50751_n19729.t361 a_50751_n19729.n319 10.1674
R50400 a_50751_n19729.t126 a_50751_n19729.n340 10.1674
R50401 a_50751_n19729.n341 a_50751_n19729.t126 10.1674
R50402 a_50751_n19729.n345 a_50751_n19729.t181 10.1674
R50403 a_50751_n19729.n393 a_50751_n19729.t168 10.1674
R50404 a_50751_n19729.t168 a_50751_n19729.n392 10.1674
R50405 a_50751_n19729.n389 a_50751_n19729.t160 10.1674
R50406 a_50751_n19729.t160 a_50751_n19729.n388 10.1674
R50407 a_50751_n19729.n385 a_50751_n19729.t234 10.1674
R50408 a_50751_n19729.t234 a_50751_n19729.n384 10.1674
R50409 a_50751_n19729.t312 a_50751_n19729.n353 10.1674
R50410 a_50751_n19729.n354 a_50751_n19729.t312 10.1674
R50411 a_50751_n19729.t360 a_50751_n19729.n361 10.1674
R50412 a_50751_n19729.n362 a_50751_n19729.t360 10.1674
R50413 a_50751_n19729.n372 a_50751_n19729.t190 10.1674
R50414 a_50751_n19729.t190 a_50751_n19729.n371 10.1674
R50415 a_50751_n19729.n366 a_50751_n19729.t271 10.1674
R50416 a_50751_n19729.t285 a_50751_n19729.n323 10.1674
R50417 a_50751_n19729.n324 a_50751_n19729.t285 10.1674
R50418 a_50751_n19729.n337 a_50751_n19729.t344 10.1674
R50419 a_50751_n19729.t344 a_50751_n19729.n336 10.1674
R50420 a_50751_n19729.n358 a_50751_n19729.t301 10.1674
R50421 a_50751_n19729.t301 a_50751_n19729.n357 10.1674
R50422 a_50751_n19729.t139 a_50751_n19729.n375 10.1674
R50423 a_50751_n19729.n376 a_50751_n19729.t139 10.1674
R50424 a_50751_n19729.n401 a_50751_n19729.t215 10.1674
R50425 a_50751_n19729.t215 a_50751_n19729.n400 10.1674
R50426 a_50751_n19729.t289 a_50751_n19729.n406 10.1674
R50427 a_50751_n19729.n407 a_50751_n19729.t289 10.1674
R50428 a_50751_n19729.t280 a_50751_n19729.n410 10.1674
R50429 a_50751_n19729.n411 a_50751_n19729.t280 10.1674
R50430 a_50751_n19729.n423 a_50751_n19729.t350 10.1674
R50431 a_50751_n19729.t350 a_50751_n19729.n422 10.1674
R50432 a_50751_n19729.n415 a_50751_n19729.t202 10.1674
R50433 a_50751_n19729.t202 a_50751_n19729.n414 10.1674
R50434 a_50751_n19729.t269 a_50751_n19729.n435 10.1674
R50435 a_50751_n19729.n436 a_50751_n19729.t269 10.1674
R50436 a_50751_n19729.n440 a_50751_n19729.t329 10.1674
R50437 a_50751_n19729.n488 a_50751_n19729.t347 10.1674
R50438 a_50751_n19729.t347 a_50751_n19729.n487 10.1674
R50439 a_50751_n19729.n484 a_50751_n19729.t334 10.1674
R50440 a_50751_n19729.t334 a_50751_n19729.n483 10.1674
R50441 a_50751_n19729.n480 a_50751_n19729.t114 10.1674
R50442 a_50751_n19729.t114 a_50751_n19729.n479 10.1674
R50443 a_50751_n19729.t183 a_50751_n19729.n448 10.1674
R50444 a_50751_n19729.n449 a_50751_n19729.t183 10.1674
R50445 a_50751_n19729.t238 a_50751_n19729.n456 10.1674
R50446 a_50751_n19729.n457 a_50751_n19729.t238 10.1674
R50447 a_50751_n19729.n467 a_50751_n19729.t84 10.1674
R50448 a_50751_n19729.t84 a_50751_n19729.n466 10.1674
R50449 a_50751_n19729.n461 a_50751_n19729.t153 10.1674
R50450 a_50751_n19729.t130 a_50751_n19729.n418 10.1674
R50451 a_50751_n19729.n419 a_50751_n19729.t130 10.1674
R50452 a_50751_n19729.n432 a_50751_n19729.t187 10.1674
R50453 a_50751_n19729.t187 a_50751_n19729.n431 10.1674
R50454 a_50751_n19729.n453 a_50751_n19729.t174 10.1674
R50455 a_50751_n19729.t174 a_50751_n19729.n452 10.1674
R50456 a_50751_n19729.t317 a_50751_n19729.n470 10.1674
R50457 a_50751_n19729.n471 a_50751_n19729.t317 10.1674
R50458 a_50751_n19729.n264 a_50751_n19729.t177 10.1674
R50459 a_50751_n19729.t177 a_50751_n19729.n263 10.1674
R50460 a_50751_n19729.t321 a_50751_n19729.n281 10.1674
R50461 a_50751_n19729.n282 a_50751_n19729.t321 10.1674
R50462 a_50751_n19729.t170 a_50751_n19729.n492 10.1409
R50463 a_50751_n19729.t204 a_50751_n19729.n269 10.1409
R50464 a_50751_n19729.t254 a_50751_n19729.n342 10.1409
R50465 a_50751_n19729.t94 a_50751_n19729.n363 10.1409
R50466 a_50751_n19729.t82 a_50751_n19729.n437 10.1409
R50467 a_50751_n19729.t349 a_50751_n19729.n458 10.1409
R50468 a_50751_n19729.t342 a_50751_n19729.n494 10.1409
R50469 a_50751_n19729.t154 a_50751_n19729.n271 10.1409
R50470 a_50751_n19729.t181 a_50751_n19729.n344 10.1409
R50471 a_50751_n19729.t271 a_50751_n19729.n365 10.1409
R50472 a_50751_n19729.t329 a_50751_n19729.n439 10.1409
R50473 a_50751_n19729.t153 a_50751_n19729.n460 10.1409
R50474 a_50751_n19729.t267 a_50751_n19729.n492 9.54631
R50475 a_50751_n19729.n213 a_50751_n19729.t341 9.54631
R50476 a_50751_n19729.t171 a_50751_n19729.n212 9.54631
R50477 a_50751_n19729.n494 a_50751_n19729.t353 9.54631
R50478 a_50751_n19729.t105 a_50751_n19729.n269 9.54631
R50479 a_50751_n19729.n215 a_50751_n19729.t298 9.54631
R50480 a_50751_n19729.t75 a_50751_n19729.n214 9.54631
R50481 a_50751_n19729.n271 a_50751_n19729.t223 9.54631
R50482 a_50751_n19729.t92 a_50751_n19729.n342 9.54631
R50483 a_50751_n19729.n217 a_50751_n19729.t262 9.54631
R50484 a_50751_n19729.t256 a_50751_n19729.n216 9.54631
R50485 a_50751_n19729.n344 a_50751_n19729.t359 9.54631
R50486 a_50751_n19729.t156 a_50751_n19729.n363 9.54631
R50487 a_50751_n19729.n219 a_50751_n19729.t313 9.54631
R50488 a_50751_n19729.t246 a_50751_n19729.n218 9.54631
R50489 a_50751_n19729.n365 a_50751_n19729.t201 9.54631
R50490 a_50751_n19729.t101 a_50751_n19729.n437 9.54631
R50491 a_50751_n19729.n221 a_50751_n19729.t200 9.54631
R50492 a_50751_n19729.t299 a_50751_n19729.n220 9.54631
R50493 a_50751_n19729.n439 a_50751_n19729.t108 9.54631
R50494 a_50751_n19729.t157 a_50751_n19729.n458 9.54631
R50495 a_50751_n19729.n223 a_50751_n19729.t113 9.54631
R50496 a_50751_n19729.t314 a_50751_n19729.n222 9.54631
R50497 a_50751_n19729.n460 a_50751_n19729.t85 9.54631
R50498 a_50751_n19729.n233 a_50751_n19729.t152 9.54355
R50499 a_50751_n19729.t152 a_50751_n19729.n232 9.54355
R50500 a_50751_n19729.t227 a_50751_n19729.n2 9.54355
R50501 a_50751_n19729.n1 a_50751_n19729.t227 9.54355
R50502 a_50751_n19729.n229 a_50751_n19729.t358 9.54355
R50503 a_50751_n19729.n0 a_50751_n19729.t358 9.54355
R50504 a_50751_n19729.n230 a_50751_n19729.t237 9.54355
R50505 a_50751_n19729.n231 a_50751_n19729.t237 9.54355
R50506 a_50751_n19729.n235 a_50751_n19729.t224 9.54355
R50507 a_50751_n19729.t224 a_50751_n19729.n234 9.54355
R50508 a_50751_n19729.t307 a_50751_n19729.n7 9.54355
R50509 a_50751_n19729.n4 a_50751_n19729.t307 9.54355
R50510 a_50751_n19729.n5 a_50751_n19729.t138 9.54355
R50511 a_50751_n19729.t138 a_50751_n19729.n3 9.54355
R50512 a_50751_n19729.n237 a_50751_n19729.t315 9.54355
R50513 a_50751_n19729.n236 a_50751_n19729.t315 9.54355
R50514 a_50751_n19729.n239 a_50751_n19729.t216 9.54355
R50515 a_50751_n19729.t216 a_50751_n19729.n238 9.54355
R50516 a_50751_n19729.t294 a_50751_n19729.n11 9.54355
R50517 a_50751_n19729.n9 a_50751_n19729.t294 9.54355
R50518 a_50751_n19729.n10 a_50751_n19729.t123 9.54355
R50519 a_50751_n19729.t123 a_50751_n19729.n8 9.54355
R50520 a_50751_n19729.n241 a_50751_n19729.t303 9.54355
R50521 a_50751_n19729.n240 a_50751_n19729.t303 9.54355
R50522 a_50751_n19729.n243 a_50751_n19729.t290 9.54355
R50523 a_50751_n19729.t290 a_50751_n19729.n242 9.54355
R50524 a_50751_n19729.t70 a_50751_n19729.n15 9.54355
R50525 a_50751_n19729.n13 a_50751_n19729.t70 9.54355
R50526 a_50751_n19729.n14 a_50751_n19729.t40 9.54355
R50527 a_50751_n19729.t40 a_50751_n19729.n12 9.54355
R50528 a_50751_n19729.n245 a_50751_n19729.t88 9.54355
R50529 a_50751_n19729.n244 a_50751_n19729.t88 9.54355
R50530 a_50751_n19729.n251 a_50751_n19729.t145 9.54355
R50531 a_50751_n19729.t145 a_50751_n19729.n250 9.54355
R50532 a_50751_n19729.t36 a_50751_n19729.n20 9.54355
R50533 a_50751_n19729.n17 a_50751_n19729.t36 9.54355
R50534 a_50751_n19729.n18 a_50751_n19729.t8 9.54355
R50535 a_50751_n19729.t8 a_50751_n19729.n16 9.54355
R50536 a_50751_n19729.n253 a_50751_n19729.t228 9.54355
R50537 a_50751_n19729.n252 a_50751_n19729.t228 9.54355
R50538 a_50751_n19729.t205 a_50751_n19729.n498 9.54355
R50539 a_50751_n19729.n499 a_50751_n19729.t205 9.54355
R50540 a_50751_n19729.n25 a_50751_n19729.t284 9.54355
R50541 a_50751_n19729.t284 a_50751_n19729.n23 9.54355
R50542 a_50751_n19729.t112 a_50751_n19729.n24 9.54355
R50543 a_50751_n19729.n21 a_50751_n19729.t112 9.54355
R50544 a_50751_n19729.n500 a_50751_n19729.t295 9.54355
R50545 a_50751_n19729.n501 a_50751_n19729.t295 9.54355
R50546 a_50751_n19729.n493 a_50751_n19729.t267 9.54355
R50547 a_50751_n19729.t341 a_50751_n19729.n497 9.54355
R50548 a_50751_n19729.n496 a_50751_n19729.t171 9.54355
R50549 a_50751_n19729.n495 a_50751_n19729.t353 9.54355
R50550 a_50751_n19729.t305 a_50751_n19729.n296 9.54355
R50551 a_50751_n19729.n297 a_50751_n19729.t305 9.54355
R50552 a_50751_n19729.n30 a_50751_n19729.t192 9.54355
R50553 a_50751_n19729.t192 a_50751_n19729.n28 9.54355
R50554 a_50751_n19729.t266 a_50751_n19729.n29 9.54355
R50555 a_50751_n19729.n26 a_50751_n19729.t266 9.54355
R50556 a_50751_n19729.n298 a_50751_n19729.t124 9.54355
R50557 a_50751_n19729.n299 a_50751_n19729.t124 9.54355
R50558 a_50751_n19729.t292 a_50751_n19729.n292 9.54355
R50559 a_50751_n19729.n293 a_50751_n19729.t292 9.54355
R50560 a_50751_n19729.n34 a_50751_n19729.t180 9.54355
R50561 a_50751_n19729.t180 a_50751_n19729.n32 9.54355
R50562 a_50751_n19729.t253 a_50751_n19729.n33 9.54355
R50563 a_50751_n19729.n31 a_50751_n19729.t253 9.54355
R50564 a_50751_n19729.n294 a_50751_n19729.t109 9.54355
R50565 a_50751_n19729.n295 a_50751_n19729.t109 9.54355
R50566 a_50751_n19729.t78 a_50751_n19729.n288 9.54355
R50567 a_50751_n19729.n289 a_50751_n19729.t78 9.54355
R50568 a_50751_n19729.n39 a_50751_n19729.t260 9.54355
R50569 a_50751_n19729.t260 a_50751_n19729.n37 9.54355
R50570 a_50751_n19729.t327 a_50751_n19729.n38 9.54355
R50571 a_50751_n19729.n35 a_50751_n19729.t327 9.54355
R50572 a_50751_n19729.n290 a_50751_n19729.t182 9.54355
R50573 a_50751_n19729.n291 a_50751_n19729.t182 9.54355
R50574 a_50751_n19729.n258 a_50751_n19729.t146 9.54355
R50575 a_50751_n19729.t146 a_50751_n19729.n257 9.54355
R50576 a_50751_n19729.t14 a_50751_n19729.n43 9.54355
R50577 a_50751_n19729.n41 a_50751_n19729.t14 9.54355
R50578 a_50751_n19729.n42 a_50751_n19729.t56 9.54355
R50579 a_50751_n19729.t56 a_50751_n19729.n40 9.54355
R50580 a_50751_n19729.n260 a_50751_n19729.t263 9.54355
R50581 a_50751_n19729.n259 a_50751_n19729.t263 9.54355
R50582 a_50751_n19729.n266 a_50751_n19729.t185 9.54355
R50583 a_50751_n19729.t185 a_50751_n19729.n265 9.54355
R50584 a_50751_n19729.t66 a_50751_n19729.n48 9.54355
R50585 a_50751_n19729.n45 a_50751_n19729.t66 9.54355
R50586 a_50751_n19729.n46 a_50751_n19729.t46 9.54355
R50587 a_50751_n19729.t46 a_50751_n19729.n44 9.54355
R50588 a_50751_n19729.n268 a_50751_n19729.t311 9.54355
R50589 a_50751_n19729.n267 a_50751_n19729.t311 9.54355
R50590 a_50751_n19729.t326 a_50751_n19729.n275 9.54355
R50591 a_50751_n19729.n276 a_50751_n19729.t326 9.54355
R50592 a_50751_n19729.n53 a_50751_n19729.t219 9.54355
R50593 a_50751_n19729.t219 a_50751_n19729.n51 9.54355
R50594 a_50751_n19729.t288 a_50751_n19729.n52 9.54355
R50595 a_50751_n19729.n49 a_50751_n19729.t288 9.54355
R50596 a_50751_n19729.n277 a_50751_n19729.t150 9.54355
R50597 a_50751_n19729.n278 a_50751_n19729.t150 9.54355
R50598 a_50751_n19729.n270 a_50751_n19729.t105 9.54355
R50599 a_50751_n19729.t298 a_50751_n19729.n274 9.54355
R50600 a_50751_n19729.n273 a_50751_n19729.t75 9.54355
R50601 a_50751_n19729.n272 a_50751_n19729.t223 9.54355
R50602 a_50751_n19729.t76 a_50751_n19729.n246 9.54355
R50603 a_50751_n19729.n247 a_50751_n19729.t76 9.54355
R50604 a_50751_n19729.n57 a_50751_n19729.t48 9.54355
R50605 a_50751_n19729.t48 a_50751_n19729.n55 9.54355
R50606 a_50751_n19729.t30 a_50751_n19729.n56 9.54355
R50607 a_50751_n19729.n54 a_50751_n19729.t30 9.54355
R50608 a_50751_n19729.n248 a_50751_n19729.t155 9.54355
R50609 a_50751_n19729.n249 a_50751_n19729.t155 9.54355
R50610 a_50751_n19729.n503 a_50751_n19729.t133 9.54355
R50611 a_50751_n19729.t133 a_50751_n19729.n502 9.54355
R50612 a_50751_n19729.t208 a_50751_n19729.n61 9.54355
R50613 a_50751_n19729.n59 a_50751_n19729.t208 9.54355
R50614 a_50751_n19729.n60 a_50751_n19729.t332 9.54355
R50615 a_50751_n19729.t332 a_50751_n19729.n58 9.54355
R50616 a_50751_n19729.n505 a_50751_n19729.t217 9.54355
R50617 a_50751_n19729.n504 a_50751_n19729.t217 9.54355
R50618 a_50751_n19729.n308 a_50751_n19729.t265 9.54355
R50619 a_50751_n19729.t265 a_50751_n19729.n307 9.54355
R50620 a_50751_n19729.t147 a_50751_n19729.n64 9.54355
R50621 a_50751_n19729.n63 a_50751_n19729.t147 9.54355
R50622 a_50751_n19729.n304 a_50751_n19729.t141 9.54355
R50623 a_50751_n19729.n62 a_50751_n19729.t141 9.54355
R50624 a_50751_n19729.n305 a_50751_n19729.t241 9.54355
R50625 a_50751_n19729.n306 a_50751_n19729.t241 9.54355
R50626 a_50751_n19729.n310 a_50751_n19729.t336 9.54355
R50627 a_50751_n19729.t336 a_50751_n19729.n309 9.54355
R50628 a_50751_n19729.t220 a_50751_n19729.n69 9.54355
R50629 a_50751_n19729.n66 a_50751_n19729.t220 9.54355
R50630 a_50751_n19729.n67 a_50751_n19729.t214 9.54355
R50631 a_50751_n19729.t214 a_50751_n19729.n65 9.54355
R50632 a_50751_n19729.n312 a_50751_n19729.t320 9.54355
R50633 a_50751_n19729.n311 a_50751_n19729.t320 9.54355
R50634 a_50751_n19729.n314 a_50751_n19729.t325 9.54355
R50635 a_50751_n19729.t325 a_50751_n19729.n313 9.54355
R50636 a_50751_n19729.t207 a_50751_n19729.n73 9.54355
R50637 a_50751_n19729.n71 a_50751_n19729.t207 9.54355
R50638 a_50751_n19729.n72 a_50751_n19729.t199 9.54355
R50639 a_50751_n19729.t199 a_50751_n19729.n70 9.54355
R50640 a_50751_n19729.n316 a_50751_n19729.t306 9.54355
R50641 a_50751_n19729.n315 a_50751_n19729.t306 9.54355
R50642 a_50751_n19729.t104 a_50751_n19729.n325 9.54355
R50643 a_50751_n19729.n326 a_50751_n19729.t104 9.54355
R50644 a_50751_n19729.n78 a_50751_n19729.t24 9.54355
R50645 a_50751_n19729.t24 a_50751_n19729.n76 9.54355
R50646 a_50751_n19729.t28 a_50751_n19729.n77 9.54355
R50647 a_50751_n19729.n74 a_50751_n19729.t28 9.54355
R50648 a_50751_n19729.n327 a_50751_n19729.t93 9.54355
R50649 a_50751_n19729.n328 a_50751_n19729.t93 9.54355
R50650 a_50751_n19729.t259 a_50751_n19729.n317 9.54355
R50651 a_50751_n19729.n318 a_50751_n19729.t259 9.54355
R50652 a_50751_n19729.n83 a_50751_n19729.t52 9.54355
R50653 a_50751_n19729.t52 a_50751_n19729.n81 9.54355
R50654 a_50751_n19729.t54 a_50751_n19729.n82 9.54355
R50655 a_50751_n19729.n79 a_50751_n19729.t54 9.54355
R50656 a_50751_n19729.n319 a_50751_n19729.t232 9.54355
R50657 a_50751_n19729.n320 a_50751_n19729.t232 9.54355
R50658 a_50751_n19729.n339 a_50751_n19729.t323 9.54355
R50659 a_50751_n19729.t323 a_50751_n19729.n338 9.54355
R50660 a_50751_n19729.t198 a_50751_n19729.n88 9.54355
R50661 a_50751_n19729.n85 a_50751_n19729.t198 9.54355
R50662 a_50751_n19729.n86 a_50751_n19729.t186 9.54355
R50663 a_50751_n19729.t186 a_50751_n19729.n84 9.54355
R50664 a_50751_n19729.n341 a_50751_n19729.t300 9.54355
R50665 a_50751_n19729.n340 a_50751_n19729.t300 9.54355
R50666 a_50751_n19729.n343 a_50751_n19729.t92 9.54355
R50667 a_50751_n19729.t262 a_50751_n19729.n347 9.54355
R50668 a_50751_n19729.n346 a_50751_n19729.t256 9.54355
R50669 a_50751_n19729.n345 a_50751_n19729.t359 9.54355
R50670 a_50751_n19729.t352 a_50751_n19729.n390 9.54355
R50671 a_50751_n19729.n391 a_50751_n19729.t352 9.54355
R50672 a_50751_n19729.n93 a_50751_n19729.t211 9.54355
R50673 a_50751_n19729.t211 a_50751_n19729.n91 9.54355
R50674 a_50751_n19729.t144 a_50751_n19729.n92 9.54355
R50675 a_50751_n19729.n89 a_50751_n19729.t144 9.54355
R50676 a_50751_n19729.n392 a_50751_n19729.t102 9.54355
R50677 a_50751_n19729.n393 a_50751_n19729.t102 9.54355
R50678 a_50751_n19729.t338 a_50751_n19729.n386 9.54355
R50679 a_50751_n19729.n387 a_50751_n19729.t338 9.54355
R50680 a_50751_n19729.n97 a_50751_n19729.t195 9.54355
R50681 a_50751_n19729.t195 a_50751_n19729.n95 9.54355
R50682 a_50751_n19729.t131 a_50751_n19729.n96 9.54355
R50683 a_50751_n19729.n94 a_50751_n19729.t131 9.54355
R50684 a_50751_n19729.n388 a_50751_n19729.t97 9.54355
R50685 a_50751_n19729.n389 a_50751_n19729.t97 9.54355
R50686 a_50751_n19729.t119 a_50751_n19729.n382 9.54355
R50687 a_50751_n19729.n383 a_50751_n19729.t119 9.54355
R50688 a_50751_n19729.n102 a_50751_n19729.t275 9.54355
R50689 a_50751_n19729.t275 a_50751_n19729.n100 9.54355
R50690 a_50751_n19729.t203 a_50751_n19729.n101 9.54355
R50691 a_50751_n19729.n98 a_50751_n19729.t203 9.54355
R50692 a_50751_n19729.n384 a_50751_n19729.t164 9.54355
R50693 a_50751_n19729.n385 a_50751_n19729.t164 9.54355
R50694 a_50751_n19729.n352 a_50751_n19729.t189 9.54355
R50695 a_50751_n19729.t189 a_50751_n19729.n351 9.54355
R50696 a_50751_n19729.t6 a_50751_n19729.n106 9.54355
R50697 a_50751_n19729.n104 a_50751_n19729.t6 9.54355
R50698 a_50751_n19729.n105 a_50751_n19729.t26 9.54355
R50699 a_50751_n19729.t26 a_50751_n19729.n103 9.54355
R50700 a_50751_n19729.n354 a_50751_n19729.t244 9.54355
R50701 a_50751_n19729.n353 a_50751_n19729.t244 9.54355
R50702 a_50751_n19729.n360 a_50751_n19729.t243 9.54355
R50703 a_50751_n19729.t243 a_50751_n19729.n359 9.54355
R50704 a_50751_n19729.t60 a_50751_n19729.n111 9.54355
R50705 a_50751_n19729.n108 a_50751_n19729.t60 9.54355
R50706 a_50751_n19729.n109 a_50751_n19729.t16 9.54355
R50707 a_50751_n19729.t16 a_50751_n19729.n107 9.54355
R50708 a_50751_n19729.n362 a_50751_n19729.t291 9.54355
R50709 a_50751_n19729.n361 a_50751_n19729.t291 9.54355
R50710 a_50751_n19729.t87 a_50751_n19729.n369 9.54355
R50711 a_50751_n19729.n370 a_50751_n19729.t87 9.54355
R50712 a_50751_n19729.n116 a_50751_n19729.t235 9.54355
R50713 a_50751_n19729.t235 a_50751_n19729.n114 9.54355
R50714 a_50751_n19729.t165 a_50751_n19729.n115 9.54355
R50715 a_50751_n19729.n112 a_50751_n19729.t165 9.54355
R50716 a_50751_n19729.n371 a_50751_n19729.t128 9.54355
R50717 a_50751_n19729.n372 a_50751_n19729.t128 9.54355
R50718 a_50751_n19729.n364 a_50751_n19729.t156 9.54355
R50719 a_50751_n19729.t313 a_50751_n19729.n368 9.54355
R50720 a_50751_n19729.n367 a_50751_n19729.t246 9.54355
R50721 a_50751_n19729.n366 a_50751_n19729.t201 9.54355
R50722 a_50751_n19729.n322 a_50751_n19729.t176 9.54355
R50723 a_50751_n19729.t176 a_50751_n19729.n321 9.54355
R50724 a_50751_n19729.t0 a_50751_n19729.n120 9.54355
R50725 a_50751_n19729.n118 a_50751_n19729.t0 9.54355
R50726 a_50751_n19729.n119 a_50751_n19729.t2 9.54355
R50727 a_50751_n19729.t2 a_50751_n19729.n117 9.54355
R50728 a_50751_n19729.n324 a_50751_n19729.t158 9.54355
R50729 a_50751_n19729.n323 a_50751_n19729.t158 9.54355
R50730 a_50751_n19729.t247 a_50751_n19729.n334 9.54355
R50731 a_50751_n19729.n335 a_50751_n19729.t247 9.54355
R50732 a_50751_n19729.n124 a_50751_n19729.t125 9.54355
R50733 a_50751_n19729.t125 a_50751_n19729.n122 9.54355
R50734 a_50751_n19729.t116 a_50751_n19729.n123 9.54355
R50735 a_50751_n19729.n121 a_50751_n19729.t116 9.54355
R50736 a_50751_n19729.n336 a_50751_n19729.t221 9.54355
R50737 a_50751_n19729.n337 a_50751_n19729.t221 9.54355
R50738 a_50751_n19729.t178 a_50751_n19729.n355 9.54355
R50739 a_50751_n19729.n356 a_50751_n19729.t178 9.54355
R50740 a_50751_n19729.n128 a_50751_n19729.t12 9.54355
R50741 a_50751_n19729.t12 a_50751_n19729.n126 9.54355
R50742 a_50751_n19729.t32 a_50751_n19729.n127 9.54355
R50743 a_50751_n19729.n125 a_50751_n19729.t32 9.54355
R50744 a_50751_n19729.n357 a_50751_n19729.t226 9.54355
R50745 a_50751_n19729.n358 a_50751_n19729.t226 9.54355
R50746 a_50751_n19729.n374 a_50751_n19729.t322 9.54355
R50747 a_50751_n19729.t322 a_50751_n19729.n373 9.54355
R50748 a_50751_n19729.t172 a_50751_n19729.n132 9.54355
R50749 a_50751_n19729.n130 a_50751_n19729.t172 9.54355
R50750 a_50751_n19729.n131 a_50751_n19729.t107 9.54355
R50751 a_50751_n19729.t107 a_50751_n19729.n129 9.54355
R50752 a_50751_n19729.n376 a_50751_n19729.t77 9.54355
R50753 a_50751_n19729.n375 a_50751_n19729.t77 9.54355
R50754 a_50751_n19729.n403 a_50751_n19729.t282 9.54355
R50755 a_50751_n19729.t282 a_50751_n19729.n402 9.54355
R50756 a_50751_n19729.t95 a_50751_n19729.n135 9.54355
R50757 a_50751_n19729.n134 a_50751_n19729.t95 9.54355
R50758 a_50751_n19729.n399 a_50751_n19729.t175 9.54355
R50759 a_50751_n19729.n133 a_50751_n19729.t175 9.54355
R50760 a_50751_n19729.n400 a_50751_n19729.t293 9.54355
R50761 a_50751_n19729.n401 a_50751_n19729.t293 9.54355
R50762 a_50751_n19729.n405 a_50751_n19729.t356 9.54355
R50763 a_50751_n19729.t356 a_50751_n19729.n404 9.54355
R50764 a_50751_n19729.t162 a_50751_n19729.n140 9.54355
R50765 a_50751_n19729.n137 a_50751_n19729.t162 9.54355
R50766 a_50751_n19729.n138 a_50751_n19729.t258 9.54355
R50767 a_50751_n19729.t258 a_50751_n19729.n136 9.54355
R50768 a_50751_n19729.n407 a_50751_n19729.t79 9.54355
R50769 a_50751_n19729.n406 a_50751_n19729.t79 9.54355
R50770 a_50751_n19729.n409 a_50751_n19729.t340 9.54355
R50771 a_50751_n19729.t340 a_50751_n19729.n408 9.54355
R50772 a_50751_n19729.t151 a_50751_n19729.n144 9.54355
R50773 a_50751_n19729.n142 a_50751_n19729.t151 9.54355
R50774 a_50751_n19729.n143 a_50751_n19729.t245 9.54355
R50775 a_50751_n19729.t245 a_50751_n19729.n141 9.54355
R50776 a_50751_n19729.n411 a_50751_n19729.t354 9.54355
R50777 a_50751_n19729.n410 a_50751_n19729.t354 9.54355
R50778 a_50751_n19729.t121 a_50751_n19729.n420 9.54355
R50779 a_50751_n19729.n421 a_50751_n19729.t121 9.54355
R50780 a_50751_n19729.n149 a_50751_n19729.t34 9.54355
R50781 a_50751_n19729.t34 a_50751_n19729.n147 9.54355
R50782 a_50751_n19729.t20 a_50751_n19729.n148 9.54355
R50783 a_50751_n19729.n145 a_50751_n19729.t20 9.54355
R50784 a_50751_n19729.n422 a_50751_n19729.t135 9.54355
R50785 a_50751_n19729.n423 a_50751_n19729.t135 9.54355
R50786 a_50751_n19729.t273 a_50751_n19729.n412 9.54355
R50787 a_50751_n19729.n413 a_50751_n19729.t273 9.54355
R50788 a_50751_n19729.n154 a_50751_n19729.t68 9.54355
R50789 a_50751_n19729.t68 a_50751_n19729.n152 9.54355
R50790 a_50751_n19729.t42 a_50751_n19729.n153 9.54355
R50791 a_50751_n19729.n150 a_50751_n19729.t42 9.54355
R50792 a_50751_n19729.n414 a_50751_n19729.t283 9.54355
R50793 a_50751_n19729.n415 a_50751_n19729.t283 9.54355
R50794 a_50751_n19729.n434 a_50751_n19729.t330 9.54355
R50795 a_50751_n19729.t330 a_50751_n19729.n433 9.54355
R50796 a_50751_n19729.t142 a_50751_n19729.n159 9.54355
R50797 a_50751_n19729.n156 a_50751_n19729.t142 9.54355
R50798 a_50751_n19729.n157 a_50751_n19729.t233 9.54355
R50799 a_50751_n19729.t233 a_50751_n19729.n155 9.54355
R50800 a_50751_n19729.n436 a_50751_n19729.t343 9.54355
R50801 a_50751_n19729.n435 a_50751_n19729.t343 9.54355
R50802 a_50751_n19729.n438 a_50751_n19729.t101 9.54355
R50803 a_50751_n19729.t200 a_50751_n19729.n442 9.54355
R50804 a_50751_n19729.n441 a_50751_n19729.t299 9.54355
R50805 a_50751_n19729.n440 a_50751_n19729.t108 9.54355
R50806 a_50751_n19729.t355 a_50751_n19729.n485 9.54355
R50807 a_50751_n19729.n486 a_50751_n19729.t355 9.54355
R50808 a_50751_n19729.n164 a_50751_n19729.t316 9.54355
R50809 a_50751_n19729.t316 a_50751_n19729.n162 9.54355
R50810 a_50751_n19729.t213 a_50751_n19729.n163 9.54355
R50811 a_50751_n19729.n160 a_50751_n19729.t213 9.54355
R50812 a_50751_n19729.n487 a_50751_n19729.t278 9.54355
R50813 a_50751_n19729.n488 a_50751_n19729.t278 9.54355
R50814 a_50751_n19729.t339 a_50751_n19729.n481 9.54355
R50815 a_50751_n19729.n482 a_50751_n19729.t339 9.54355
R50816 a_50751_n19729.n168 a_50751_n19729.t304 9.54355
R50817 a_50751_n19729.t304 a_50751_n19729.n166 9.54355
R50818 a_50751_n19729.t197 a_50751_n19729.n167 9.54355
R50819 a_50751_n19729.n165 a_50751_n19729.t197 9.54355
R50820 a_50751_n19729.n483 a_50751_n19729.t264 9.54355
R50821 a_50751_n19729.n484 a_50751_n19729.t264 9.54355
R50822 a_50751_n19729.t120 a_50751_n19729.n477 9.54355
R50823 a_50751_n19729.n478 a_50751_n19729.t120 9.54355
R50824 a_50751_n19729.n173 a_50751_n19729.t89 9.54355
R50825 a_50751_n19729.t89 a_50751_n19729.n171 9.54355
R50826 a_50751_n19729.t277 a_50751_n19729.n172 9.54355
R50827 a_50751_n19729.n169 a_50751_n19729.t277 9.54355
R50828 a_50751_n19729.n479 a_50751_n19729.t335 9.54355
R50829 a_50751_n19729.n480 a_50751_n19729.t335 9.54355
R50830 a_50751_n19729.n447 a_50751_n19729.t191 9.54355
R50831 a_50751_n19729.t191 a_50751_n19729.n446 9.54355
R50832 a_50751_n19729.t44 a_50751_n19729.n177 9.54355
R50833 a_50751_n19729.n175 a_50751_n19729.t44 9.54355
R50834 a_50751_n19729.n176 a_50751_n19729.t4 9.54355
R50835 a_50751_n19729.t4 a_50751_n19729.n174 9.54355
R50836 a_50751_n19729.n449 a_50751_n19729.t117 9.54355
R50837 a_50751_n19729.n448 a_50751_n19729.t117 9.54355
R50838 a_50751_n19729.n455 a_50751_n19729.t248 9.54355
R50839 a_50751_n19729.t248 a_50751_n19729.n454 9.54355
R50840 a_50751_n19729.t38 a_50751_n19729.n182 9.54355
R50841 a_50751_n19729.n179 a_50751_n19729.t38 9.54355
R50842 a_50751_n19729.n180 a_50751_n19729.t58 9.54355
R50843 a_50751_n19729.t58 a_50751_n19729.n178 9.54355
R50844 a_50751_n19729.n457 a_50751_n19729.t163 9.54355
R50845 a_50751_n19729.n456 a_50751_n19729.t163 9.54355
R50846 a_50751_n19729.t90 a_50751_n19729.n464 9.54355
R50847 a_50751_n19729.n465 a_50751_n19729.t90 9.54355
R50848 a_50751_n19729.n187 a_50751_n19729.t333 9.54355
R50849 a_50751_n19729.t333 a_50751_n19729.n185 9.54355
R50850 a_50751_n19729.t236 a_50751_n19729.n186 9.54355
R50851 a_50751_n19729.n183 a_50751_n19729.t236 9.54355
R50852 a_50751_n19729.n466 a_50751_n19729.t302 9.54355
R50853 a_50751_n19729.n467 a_50751_n19729.t302 9.54355
R50854 a_50751_n19729.n459 a_50751_n19729.t157 9.54355
R50855 a_50751_n19729.t113 a_50751_n19729.n463 9.54355
R50856 a_50751_n19729.n462 a_50751_n19729.t314 9.54355
R50857 a_50751_n19729.n461 a_50751_n19729.t85 9.54355
R50858 a_50751_n19729.n417 a_50751_n19729.t193 9.54355
R50859 a_50751_n19729.t193 a_50751_n19729.n416 9.54355
R50860 a_50751_n19729.t22 a_50751_n19729.n191 9.54355
R50861 a_50751_n19729.n189 a_50751_n19729.t22 9.54355
R50862 a_50751_n19729.n190 a_50751_n19729.t62 9.54355
R50863 a_50751_n19729.t62 a_50751_n19729.n188 9.54355
R50864 a_50751_n19729.n419 a_50751_n19729.t206 9.54355
R50865 a_50751_n19729.n418 a_50751_n19729.t206 9.54355
R50866 a_50751_n19729.t261 a_50751_n19729.n429 9.54355
R50867 a_50751_n19729.n430 a_50751_n19729.t261 9.54355
R50868 a_50751_n19729.n195 a_50751_n19729.t74 9.54355
R50869 a_50751_n19729.t74 a_50751_n19729.n193 9.54355
R50870 a_50751_n19729.t159 a_50751_n19729.n194 9.54355
R50871 a_50751_n19729.n192 a_50751_n19729.t159 9.54355
R50872 a_50751_n19729.n431 a_50751_n19729.t270 9.54355
R50873 a_50751_n19729.n432 a_50751_n19729.t270 9.54355
R50874 a_50751_n19729.t179 a_50751_n19729.n450 9.54355
R50875 a_50751_n19729.n451 a_50751_n19729.t179 9.54355
R50876 a_50751_n19729.n199 a_50751_n19729.t50 9.54355
R50877 a_50751_n19729.t50 a_50751_n19729.n197 9.54355
R50878 a_50751_n19729.t10 a_50751_n19729.n198 9.54355
R50879 a_50751_n19729.n196 a_50751_n19729.t10 9.54355
R50880 a_50751_n19729.n452 a_50751_n19729.t103 9.54355
R50881 a_50751_n19729.n453 a_50751_n19729.t103 9.54355
R50882 a_50751_n19729.n469 a_50751_n19729.t324 9.54355
R50883 a_50751_n19729.t324 a_50751_n19729.n468 9.54355
R50884 a_50751_n19729.t281 a_50751_n19729.n203 9.54355
R50885 a_50751_n19729.n201 a_50751_n19729.t281 9.54355
R50886 a_50751_n19729.n202 a_50751_n19729.t173 9.54355
R50887 a_50751_n19729.t173 a_50751_n19729.n200 9.54355
R50888 a_50751_n19729.n471 a_50751_n19729.t240 9.54355
R50889 a_50751_n19729.n470 a_50751_n19729.t240 9.54355
R50890 a_50751_n19729.t134 a_50751_n19729.n261 9.54355
R50891 a_50751_n19729.n262 a_50751_n19729.t134 9.54355
R50892 a_50751_n19729.n207 a_50751_n19729.t18 9.54355
R50893 a_50751_n19729.t18 a_50751_n19729.n205 9.54355
R50894 a_50751_n19729.t64 a_50751_n19729.n206 9.54355
R50895 a_50751_n19729.n204 a_50751_n19729.t64 9.54355
R50896 a_50751_n19729.n263 a_50751_n19729.t251 9.54355
R50897 a_50751_n19729.n264 a_50751_n19729.t251 9.54355
R50898 a_50751_n19729.n280 a_50751_n19729.t268 9.54355
R50899 a_50751_n19729.t268 a_50751_n19729.n279 9.54355
R50900 a_50751_n19729.t161 a_50751_n19729.n211 9.54355
R50901 a_50751_n19729.n209 a_50751_n19729.t161 9.54355
R50902 a_50751_n19729.n210 a_50751_n19729.t225 9.54355
R50903 a_50751_n19729.t225 a_50751_n19729.n208 9.54355
R50904 a_50751_n19729.n282 a_50751_n19729.t96 9.54355
R50905 a_50751_n19729.n281 a_50751_n19729.t96 9.54355
R50906 a_50751_n19729.n300 a_50751_n19729.t72 7.11376
R50907 a_50751_n19729.n395 a_50751_n19729.n300 6.02769
R50908 a_50751_n19729.n491 a_50751_n19729.n490 3.90251
R50909 a_50751_n19729.n508 a_50751_n19729.t49 3.3605
R50910 a_50751_n19729.n507 a_50751_n19729.t37 3.3605
R50911 a_50751_n19729.n226 a_50751_n19729.t41 3.3605
R50912 a_50751_n19729.n227 a_50751_n19729.t31 3.3605
R50913 a_50751_n19729.n228 a_50751_n19729.t9 3.3605
R50914 a_50751_n19729.n303 a_50751_n19729.t29 3.3605
R50915 a_50751_n19729.n302 a_50751_n19729.t3 3.3605
R50916 a_50751_n19729.n301 a_50751_n19729.t55 3.3605
R50917 a_50751_n19729.n330 a_50751_n19729.t25 3.3605
R50918 a_50751_n19729.n331 a_50751_n19729.t1 3.3605
R50919 a_50751_n19729.n332 a_50751_n19729.t53 3.3605
R50920 a_50751_n19729.n348 a_50751_n19729.t27 3.3605
R50921 a_50751_n19729.n349 a_50751_n19729.t33 3.3605
R50922 a_50751_n19729.n350 a_50751_n19729.t17 3.3605
R50923 a_50751_n19729.n380 a_50751_n19729.t7 3.3605
R50924 a_50751_n19729.n379 a_50751_n19729.t13 3.3605
R50925 a_50751_n19729.n378 a_50751_n19729.t61 3.3605
R50926 a_50751_n19729.n398 a_50751_n19729.t21 3.3605
R50927 a_50751_n19729.n397 a_50751_n19729.t63 3.3605
R50928 a_50751_n19729.n396 a_50751_n19729.t43 3.3605
R50929 a_50751_n19729.n425 a_50751_n19729.t35 3.3605
R50930 a_50751_n19729.n426 a_50751_n19729.t23 3.3605
R50931 a_50751_n19729.n427 a_50751_n19729.t69 3.3605
R50932 a_50751_n19729.n443 a_50751_n19729.t5 3.3605
R50933 a_50751_n19729.n444 a_50751_n19729.t11 3.3605
R50934 a_50751_n19729.n445 a_50751_n19729.t59 3.3605
R50935 a_50751_n19729.n475 a_50751_n19729.t45 3.3605
R50936 a_50751_n19729.n474 a_50751_n19729.t51 3.3605
R50937 a_50751_n19729.n473 a_50751_n19729.t39 3.3605
R50938 a_50751_n19729.n254 a_50751_n19729.t57 3.3605
R50939 a_50751_n19729.n255 a_50751_n19729.t65 3.3605
R50940 a_50751_n19729.n256 a_50751_n19729.t47 3.3605
R50941 a_50751_n19729.n286 a_50751_n19729.t15 3.3605
R50942 a_50751_n19729.n285 a_50751_n19729.t19 3.3605
R50943 a_50751_n19729.n284 a_50751_n19729.t67 3.3605
R50944 a_50751_n19729.t71 a_50751_n19729.n509 3.3605
R50945 a_50751_n19729.n490 a_50751_n19729.n395 3.14899
R50946 a_50751_n19729.n333 a_50751_n19729.n301 2.59662
R50947 a_50751_n19729.n377 a_50751_n19729.n350 2.59662
R50948 a_50751_n19729.n428 a_50751_n19729.n396 2.59662
R50949 a_50751_n19729.n472 a_50751_n19729.n445 2.59662
R50950 a_50751_n19729.n283 a_50751_n19729.n256 2.59662
R50951 a_50751_n19729.n506 a_50751_n19729.n228 2.59662
R50952 a_50751_n19729.n226 a_50751_n19729.n225 2.59544
R50953 a_50751_n19729.n329 a_50751_n19729.n303 2.59544
R50954 a_50751_n19729.n381 a_50751_n19729.n348 2.59544
R50955 a_50751_n19729.n424 a_50751_n19729.n398 2.59544
R50956 a_50751_n19729.n476 a_50751_n19729.n443 2.59544
R50957 a_50751_n19729.n287 a_50751_n19729.n254 2.59544
R50958 a_50751_n19729.n333 a_50751_n19729.n332 2.58354
R50959 a_50751_n19729.n378 a_50751_n19729.n377 2.58354
R50960 a_50751_n19729.n428 a_50751_n19729.n427 2.58354
R50961 a_50751_n19729.n473 a_50751_n19729.n472 2.58354
R50962 a_50751_n19729.n284 a_50751_n19729.n283 2.58354
R50963 a_50751_n19729.n507 a_50751_n19729.n506 2.58354
R50964 a_50751_n19729.n509 a_50751_n19729.n225 2.58235
R50965 a_50751_n19729.n330 a_50751_n19729.n329 2.58235
R50966 a_50751_n19729.n381 a_50751_n19729.n380 2.58235
R50967 a_50751_n19729.n425 a_50751_n19729.n424 2.58235
R50968 a_50751_n19729.n476 a_50751_n19729.n475 2.58235
R50969 a_50751_n19729.n287 a_50751_n19729.n286 2.58235
R50970 a_50751_n19729.n68 a_50751_n19729.n64 1.6805
R50971 a_50751_n19729.n139 a_50751_n19729.n135 1.6805
R50972 a_50751_n19729.n6 a_50751_n19729.n2 1.6805
R50973 a_50751_n19729.n113 a_50751_n19729.n219 1.59324
R50974 a_50751_n19729.n184 a_50751_n19729.n223 1.59324
R50975 a_50751_n19729.n50 a_50751_n19729.n215 1.59324
R50976 a_50751_n19729.n132 a_50751_n19729.n113 1.5005
R50977 a_50751_n19729.n377 a_50751_n19729.n113 1.5005
R50978 a_50751_n19729.n110 a_50751_n19729.n128 1.5005
R50979 a_50751_n19729.n99 a_50751_n19729.n381 1.5005
R50980 a_50751_n19729.n87 a_50751_n19729.n124 1.5005
R50981 a_50751_n19729.n80 a_50751_n19729.n333 1.5005
R50982 a_50751_n19729.n120 a_50751_n19729.n75 1.5005
R50983 a_50751_n19729.n329 a_50751_n19729.n68 1.5005
R50984 a_50751_n19729.n113 a_50751_n19729.n116 1.5005
R50985 a_50751_n19729.n114 a_50751_n19729.n113 1.5005
R50986 a_50751_n19729.n113 a_50751_n19729.n130 1.5005
R50987 a_50751_n19729.n111 a_50751_n19729.n110 1.5005
R50988 a_50751_n19729.n113 a_50751_n19729.n108 1.5005
R50989 a_50751_n19729.n126 a_50751_n19729.n110 1.5005
R50990 a_50751_n19729.n106 a_50751_n19729.n99 1.5005
R50991 a_50751_n19729.n110 a_50751_n19729.n104 1.5005
R50992 a_50751_n19729.n90 a_50751_n19729.n102 1.5005
R50993 a_50751_n19729.n100 a_50751_n19729.n99 1.5005
R50994 a_50751_n19729.n90 a_50751_n19729.n97 1.5005
R50995 a_50751_n19729.n95 a_50751_n19729.n90 1.5005
R50996 a_50751_n19729.n90 a_50751_n19729.n93 1.5005
R50997 a_50751_n19729.n91 a_50751_n19729.n90 1.5005
R50998 a_50751_n19729.n87 a_50751_n19729.n217 1.5005
R50999 a_50751_n19729.n88 a_50751_n19729.n87 1.5005
R51000 a_50751_n19729.n87 a_50751_n19729.n85 1.5005
R51001 a_50751_n19729.n122 a_50751_n19729.n80 1.5005
R51002 a_50751_n19729.n75 a_50751_n19729.n83 1.5005
R51003 a_50751_n19729.n81 a_50751_n19729.n80 1.5005
R51004 a_50751_n19729.n75 a_50751_n19729.n118 1.5005
R51005 a_50751_n19729.n68 a_50751_n19729.n78 1.5005
R51006 a_50751_n19729.n76 a_50751_n19729.n75 1.5005
R51007 a_50751_n19729.n73 a_50751_n19729.n68 1.5005
R51008 a_50751_n19729.n68 a_50751_n19729.n71 1.5005
R51009 a_50751_n19729.n69 a_50751_n19729.n68 1.5005
R51010 a_50751_n19729.n68 a_50751_n19729.n66 1.5005
R51011 a_50751_n19729.n68 a_50751_n19729.n63 1.5005
R51012 a_50751_n19729.n203 a_50751_n19729.n184 1.5005
R51013 a_50751_n19729.n472 a_50751_n19729.n184 1.5005
R51014 a_50751_n19729.n181 a_50751_n19729.n199 1.5005
R51015 a_50751_n19729.n170 a_50751_n19729.n476 1.5005
R51016 a_50751_n19729.n158 a_50751_n19729.n195 1.5005
R51017 a_50751_n19729.n151 a_50751_n19729.n428 1.5005
R51018 a_50751_n19729.n191 a_50751_n19729.n146 1.5005
R51019 a_50751_n19729.n424 a_50751_n19729.n139 1.5005
R51020 a_50751_n19729.n184 a_50751_n19729.n187 1.5005
R51021 a_50751_n19729.n185 a_50751_n19729.n184 1.5005
R51022 a_50751_n19729.n184 a_50751_n19729.n201 1.5005
R51023 a_50751_n19729.n182 a_50751_n19729.n181 1.5005
R51024 a_50751_n19729.n184 a_50751_n19729.n179 1.5005
R51025 a_50751_n19729.n197 a_50751_n19729.n181 1.5005
R51026 a_50751_n19729.n177 a_50751_n19729.n170 1.5005
R51027 a_50751_n19729.n181 a_50751_n19729.n175 1.5005
R51028 a_50751_n19729.n161 a_50751_n19729.n173 1.5005
R51029 a_50751_n19729.n171 a_50751_n19729.n170 1.5005
R51030 a_50751_n19729.n161 a_50751_n19729.n168 1.5005
R51031 a_50751_n19729.n166 a_50751_n19729.n161 1.5005
R51032 a_50751_n19729.n161 a_50751_n19729.n164 1.5005
R51033 a_50751_n19729.n162 a_50751_n19729.n161 1.5005
R51034 a_50751_n19729.n158 a_50751_n19729.n221 1.5005
R51035 a_50751_n19729.n159 a_50751_n19729.n158 1.5005
R51036 a_50751_n19729.n158 a_50751_n19729.n156 1.5005
R51037 a_50751_n19729.n193 a_50751_n19729.n151 1.5005
R51038 a_50751_n19729.n146 a_50751_n19729.n154 1.5005
R51039 a_50751_n19729.n152 a_50751_n19729.n151 1.5005
R51040 a_50751_n19729.n146 a_50751_n19729.n189 1.5005
R51041 a_50751_n19729.n139 a_50751_n19729.n149 1.5005
R51042 a_50751_n19729.n147 a_50751_n19729.n146 1.5005
R51043 a_50751_n19729.n144 a_50751_n19729.n139 1.5005
R51044 a_50751_n19729.n139 a_50751_n19729.n142 1.5005
R51045 a_50751_n19729.n140 a_50751_n19729.n139 1.5005
R51046 a_50751_n19729.n139 a_50751_n19729.n137 1.5005
R51047 a_50751_n19729.n139 a_50751_n19729.n134 1.5005
R51048 a_50751_n19729.n211 a_50751_n19729.n50 1.5005
R51049 a_50751_n19729.n283 a_50751_n19729.n50 1.5005
R51050 a_50751_n19729.n47 a_50751_n19729.n207 1.5005
R51051 a_50751_n19729.n36 a_50751_n19729.n287 1.5005
R51052 a_50751_n19729.n61 a_50751_n19729.n22 1.5005
R51053 a_50751_n19729.n19 a_50751_n19729.n57 1.5005
R51054 a_50751_n19729.n6 a_50751_n19729.n225 1.5005
R51055 a_50751_n19729.n50 a_50751_n19729.n53 1.5005
R51056 a_50751_n19729.n51 a_50751_n19729.n50 1.5005
R51057 a_50751_n19729.n50 a_50751_n19729.n209 1.5005
R51058 a_50751_n19729.n48 a_50751_n19729.n47 1.5005
R51059 a_50751_n19729.n50 a_50751_n19729.n45 1.5005
R51060 a_50751_n19729.n205 a_50751_n19729.n47 1.5005
R51061 a_50751_n19729.n43 a_50751_n19729.n36 1.5005
R51062 a_50751_n19729.n47 a_50751_n19729.n41 1.5005
R51063 a_50751_n19729.n27 a_50751_n19729.n39 1.5005
R51064 a_50751_n19729.n37 a_50751_n19729.n36 1.5005
R51065 a_50751_n19729.n27 a_50751_n19729.n34 1.5005
R51066 a_50751_n19729.n32 a_50751_n19729.n27 1.5005
R51067 a_50751_n19729.n27 a_50751_n19729.n30 1.5005
R51068 a_50751_n19729.n28 a_50751_n19729.n27 1.5005
R51069 a_50751_n19729.n22 a_50751_n19729.n213 1.5005
R51070 a_50751_n19729.n22 a_50751_n19729.n25 1.5005
R51071 a_50751_n19729.n23 a_50751_n19729.n22 1.5005
R51072 a_50751_n19729.n224 a_50751_n19729.n59 1.5005
R51073 a_50751_n19729.n20 a_50751_n19729.n19 1.5005
R51074 a_50751_n19729.n224 a_50751_n19729.n17 1.5005
R51075 a_50751_n19729.n55 a_50751_n19729.n19 1.5005
R51076 a_50751_n19729.n15 a_50751_n19729.n6 1.5005
R51077 a_50751_n19729.n19 a_50751_n19729.n13 1.5005
R51078 a_50751_n19729.n11 a_50751_n19729.n6 1.5005
R51079 a_50751_n19729.n6 a_50751_n19729.n9 1.5005
R51080 a_50751_n19729.n7 a_50751_n19729.n6 1.5005
R51081 a_50751_n19729.n6 a_50751_n19729.n4 1.5005
R51082 a_50751_n19729.n6 a_50751_n19729.n1 1.5005
R51083 a_50751_n19729.n506 a_50751_n19729.n224 1.5005
R51084 a_50751_n19729.n227 a_50751_n19729.n226 1.06274
R51085 a_50751_n19729.n228 a_50751_n19729.n227 1.06274
R51086 a_50751_n19729.n331 a_50751_n19729.n330 1.06274
R51087 a_50751_n19729.n332 a_50751_n19729.n331 1.06274
R51088 a_50751_n19729.n303 a_50751_n19729.n302 1.06274
R51089 a_50751_n19729.n302 a_50751_n19729.n301 1.06274
R51090 a_50751_n19729.n380 a_50751_n19729.n379 1.06274
R51091 a_50751_n19729.n379 a_50751_n19729.n378 1.06274
R51092 a_50751_n19729.n349 a_50751_n19729.n348 1.06274
R51093 a_50751_n19729.n350 a_50751_n19729.n349 1.06274
R51094 a_50751_n19729.n426 a_50751_n19729.n425 1.06274
R51095 a_50751_n19729.n427 a_50751_n19729.n426 1.06274
R51096 a_50751_n19729.n398 a_50751_n19729.n397 1.06274
R51097 a_50751_n19729.n397 a_50751_n19729.n396 1.06274
R51098 a_50751_n19729.n475 a_50751_n19729.n474 1.06274
R51099 a_50751_n19729.n474 a_50751_n19729.n473 1.06274
R51100 a_50751_n19729.n444 a_50751_n19729.n443 1.06274
R51101 a_50751_n19729.n445 a_50751_n19729.n444 1.06274
R51102 a_50751_n19729.n286 a_50751_n19729.n285 1.06274
R51103 a_50751_n19729.n285 a_50751_n19729.n284 1.06274
R51104 a_50751_n19729.n255 a_50751_n19729.n254 1.06274
R51105 a_50751_n19729.n256 a_50751_n19729.n255 1.06274
R51106 a_50751_n19729.n509 a_50751_n19729.n508 1.06274
R51107 a_50751_n19729.n508 a_50751_n19729.n507 1.06274
R51108 a_50751_n19729.n0 a_50751_n19729.n231 0.97759
R51109 a_50751_n19729.n1 a_50751_n19729.n232 0.97759
R51110 a_50751_n19729.n230 a_50751_n19729.n229 0.97759
R51111 a_50751_n19729.n2 a_50751_n19729.n233 0.97759
R51112 a_50751_n19729.n236 a_50751_n19729.n3 0.97759
R51113 a_50751_n19729.n4 a_50751_n19729.n234 0.97759
R51114 a_50751_n19729.n5 a_50751_n19729.n237 0.97759
R51115 a_50751_n19729.n7 a_50751_n19729.n235 0.97759
R51116 a_50751_n19729.n240 a_50751_n19729.n8 0.97759
R51117 a_50751_n19729.n9 a_50751_n19729.n238 0.97759
R51118 a_50751_n19729.n10 a_50751_n19729.n241 0.97759
R51119 a_50751_n19729.n11 a_50751_n19729.n239 0.97759
R51120 a_50751_n19729.n244 a_50751_n19729.n12 0.97759
R51121 a_50751_n19729.n13 a_50751_n19729.n242 0.97759
R51122 a_50751_n19729.n14 a_50751_n19729.n245 0.97759
R51123 a_50751_n19729.n15 a_50751_n19729.n243 0.97759
R51124 a_50751_n19729.n252 a_50751_n19729.n16 0.97759
R51125 a_50751_n19729.n17 a_50751_n19729.n250 0.97759
R51126 a_50751_n19729.n18 a_50751_n19729.n253 0.97759
R51127 a_50751_n19729.n20 a_50751_n19729.n251 0.97759
R51128 a_50751_n19729.n21 a_50751_n19729.n501 0.97759
R51129 a_50751_n19729.n23 a_50751_n19729.n499 0.97759
R51130 a_50751_n19729.n500 a_50751_n19729.n24 0.97759
R51131 a_50751_n19729.n25 a_50751_n19729.n498 0.97759
R51132 a_50751_n19729.n496 a_50751_n19729.n495 0.97759
R51133 a_50751_n19729.n497 a_50751_n19729.n493 0.97759
R51134 a_50751_n19729.n26 a_50751_n19729.n299 0.97759
R51135 a_50751_n19729.n28 a_50751_n19729.n297 0.97759
R51136 a_50751_n19729.n298 a_50751_n19729.n29 0.97759
R51137 a_50751_n19729.n30 a_50751_n19729.n296 0.97759
R51138 a_50751_n19729.n31 a_50751_n19729.n295 0.97759
R51139 a_50751_n19729.n32 a_50751_n19729.n293 0.97759
R51140 a_50751_n19729.n294 a_50751_n19729.n33 0.97759
R51141 a_50751_n19729.n34 a_50751_n19729.n292 0.97759
R51142 a_50751_n19729.n35 a_50751_n19729.n291 0.97759
R51143 a_50751_n19729.n37 a_50751_n19729.n289 0.97759
R51144 a_50751_n19729.n290 a_50751_n19729.n38 0.97759
R51145 a_50751_n19729.n39 a_50751_n19729.n288 0.97759
R51146 a_50751_n19729.n259 a_50751_n19729.n40 0.97759
R51147 a_50751_n19729.n41 a_50751_n19729.n257 0.97759
R51148 a_50751_n19729.n42 a_50751_n19729.n260 0.97759
R51149 a_50751_n19729.n43 a_50751_n19729.n258 0.97759
R51150 a_50751_n19729.n267 a_50751_n19729.n44 0.97759
R51151 a_50751_n19729.n45 a_50751_n19729.n265 0.97759
R51152 a_50751_n19729.n46 a_50751_n19729.n268 0.97759
R51153 a_50751_n19729.n48 a_50751_n19729.n266 0.97759
R51154 a_50751_n19729.n49 a_50751_n19729.n278 0.97759
R51155 a_50751_n19729.n51 a_50751_n19729.n276 0.97759
R51156 a_50751_n19729.n277 a_50751_n19729.n52 0.97759
R51157 a_50751_n19729.n53 a_50751_n19729.n275 0.97759
R51158 a_50751_n19729.n273 a_50751_n19729.n272 0.97759
R51159 a_50751_n19729.n274 a_50751_n19729.n270 0.97759
R51160 a_50751_n19729.n54 a_50751_n19729.n249 0.97759
R51161 a_50751_n19729.n55 a_50751_n19729.n247 0.97759
R51162 a_50751_n19729.n248 a_50751_n19729.n56 0.97759
R51163 a_50751_n19729.n57 a_50751_n19729.n246 0.97759
R51164 a_50751_n19729.n504 a_50751_n19729.n58 0.97759
R51165 a_50751_n19729.n59 a_50751_n19729.n502 0.97759
R51166 a_50751_n19729.n60 a_50751_n19729.n505 0.97759
R51167 a_50751_n19729.n61 a_50751_n19729.n503 0.97759
R51168 a_50751_n19729.n62 a_50751_n19729.n306 0.97759
R51169 a_50751_n19729.n63 a_50751_n19729.n307 0.97759
R51170 a_50751_n19729.n305 a_50751_n19729.n304 0.97759
R51171 a_50751_n19729.n64 a_50751_n19729.n308 0.97759
R51172 a_50751_n19729.n311 a_50751_n19729.n65 0.97759
R51173 a_50751_n19729.n66 a_50751_n19729.n309 0.97759
R51174 a_50751_n19729.n67 a_50751_n19729.n312 0.97759
R51175 a_50751_n19729.n69 a_50751_n19729.n310 0.97759
R51176 a_50751_n19729.n315 a_50751_n19729.n70 0.97759
R51177 a_50751_n19729.n71 a_50751_n19729.n313 0.97759
R51178 a_50751_n19729.n72 a_50751_n19729.n316 0.97759
R51179 a_50751_n19729.n73 a_50751_n19729.n314 0.97759
R51180 a_50751_n19729.n74 a_50751_n19729.n328 0.97759
R51181 a_50751_n19729.n76 a_50751_n19729.n326 0.97759
R51182 a_50751_n19729.n327 a_50751_n19729.n77 0.97759
R51183 a_50751_n19729.n78 a_50751_n19729.n325 0.97759
R51184 a_50751_n19729.n79 a_50751_n19729.n320 0.97759
R51185 a_50751_n19729.n81 a_50751_n19729.n318 0.97759
R51186 a_50751_n19729.n319 a_50751_n19729.n82 0.97759
R51187 a_50751_n19729.n83 a_50751_n19729.n317 0.97759
R51188 a_50751_n19729.n340 a_50751_n19729.n84 0.97759
R51189 a_50751_n19729.n85 a_50751_n19729.n338 0.97759
R51190 a_50751_n19729.n86 a_50751_n19729.n341 0.97759
R51191 a_50751_n19729.n88 a_50751_n19729.n339 0.97759
R51192 a_50751_n19729.n346 a_50751_n19729.n345 0.97759
R51193 a_50751_n19729.n347 a_50751_n19729.n343 0.97759
R51194 a_50751_n19729.n89 a_50751_n19729.n393 0.97759
R51195 a_50751_n19729.n91 a_50751_n19729.n391 0.97759
R51196 a_50751_n19729.n392 a_50751_n19729.n92 0.97759
R51197 a_50751_n19729.n93 a_50751_n19729.n390 0.97759
R51198 a_50751_n19729.n94 a_50751_n19729.n389 0.97759
R51199 a_50751_n19729.n95 a_50751_n19729.n387 0.97759
R51200 a_50751_n19729.n388 a_50751_n19729.n96 0.97759
R51201 a_50751_n19729.n97 a_50751_n19729.n386 0.97759
R51202 a_50751_n19729.n98 a_50751_n19729.n385 0.97759
R51203 a_50751_n19729.n100 a_50751_n19729.n383 0.97759
R51204 a_50751_n19729.n384 a_50751_n19729.n101 0.97759
R51205 a_50751_n19729.n102 a_50751_n19729.n382 0.97759
R51206 a_50751_n19729.n353 a_50751_n19729.n103 0.97759
R51207 a_50751_n19729.n104 a_50751_n19729.n351 0.97759
R51208 a_50751_n19729.n105 a_50751_n19729.n354 0.97759
R51209 a_50751_n19729.n106 a_50751_n19729.n352 0.97759
R51210 a_50751_n19729.n361 a_50751_n19729.n107 0.97759
R51211 a_50751_n19729.n108 a_50751_n19729.n359 0.97759
R51212 a_50751_n19729.n109 a_50751_n19729.n362 0.97759
R51213 a_50751_n19729.n111 a_50751_n19729.n360 0.97759
R51214 a_50751_n19729.n112 a_50751_n19729.n372 0.97759
R51215 a_50751_n19729.n114 a_50751_n19729.n370 0.97759
R51216 a_50751_n19729.n371 a_50751_n19729.n115 0.97759
R51217 a_50751_n19729.n116 a_50751_n19729.n369 0.97759
R51218 a_50751_n19729.n367 a_50751_n19729.n366 0.97759
R51219 a_50751_n19729.n368 a_50751_n19729.n364 0.97759
R51220 a_50751_n19729.n323 a_50751_n19729.n117 0.97759
R51221 a_50751_n19729.n118 a_50751_n19729.n321 0.97759
R51222 a_50751_n19729.n119 a_50751_n19729.n324 0.97759
R51223 a_50751_n19729.n120 a_50751_n19729.n322 0.97759
R51224 a_50751_n19729.n121 a_50751_n19729.n337 0.97759
R51225 a_50751_n19729.n122 a_50751_n19729.n335 0.97759
R51226 a_50751_n19729.n336 a_50751_n19729.n123 0.97759
R51227 a_50751_n19729.n124 a_50751_n19729.n334 0.97759
R51228 a_50751_n19729.n125 a_50751_n19729.n358 0.97759
R51229 a_50751_n19729.n126 a_50751_n19729.n356 0.97759
R51230 a_50751_n19729.n357 a_50751_n19729.n127 0.97759
R51231 a_50751_n19729.n128 a_50751_n19729.n355 0.97759
R51232 a_50751_n19729.n375 a_50751_n19729.n129 0.97759
R51233 a_50751_n19729.n130 a_50751_n19729.n373 0.97759
R51234 a_50751_n19729.n131 a_50751_n19729.n376 0.97759
R51235 a_50751_n19729.n132 a_50751_n19729.n374 0.97759
R51236 a_50751_n19729.n133 a_50751_n19729.n401 0.97759
R51237 a_50751_n19729.n134 a_50751_n19729.n402 0.97759
R51238 a_50751_n19729.n400 a_50751_n19729.n399 0.97759
R51239 a_50751_n19729.n135 a_50751_n19729.n403 0.97759
R51240 a_50751_n19729.n406 a_50751_n19729.n136 0.97759
R51241 a_50751_n19729.n137 a_50751_n19729.n404 0.97759
R51242 a_50751_n19729.n138 a_50751_n19729.n407 0.97759
R51243 a_50751_n19729.n140 a_50751_n19729.n405 0.97759
R51244 a_50751_n19729.n410 a_50751_n19729.n141 0.97759
R51245 a_50751_n19729.n142 a_50751_n19729.n408 0.97759
R51246 a_50751_n19729.n143 a_50751_n19729.n411 0.97759
R51247 a_50751_n19729.n144 a_50751_n19729.n409 0.97759
R51248 a_50751_n19729.n145 a_50751_n19729.n423 0.97759
R51249 a_50751_n19729.n147 a_50751_n19729.n421 0.97759
R51250 a_50751_n19729.n422 a_50751_n19729.n148 0.97759
R51251 a_50751_n19729.n149 a_50751_n19729.n420 0.97759
R51252 a_50751_n19729.n150 a_50751_n19729.n415 0.97759
R51253 a_50751_n19729.n152 a_50751_n19729.n413 0.97759
R51254 a_50751_n19729.n414 a_50751_n19729.n153 0.97759
R51255 a_50751_n19729.n154 a_50751_n19729.n412 0.97759
R51256 a_50751_n19729.n435 a_50751_n19729.n155 0.97759
R51257 a_50751_n19729.n156 a_50751_n19729.n433 0.97759
R51258 a_50751_n19729.n157 a_50751_n19729.n436 0.97759
R51259 a_50751_n19729.n159 a_50751_n19729.n434 0.97759
R51260 a_50751_n19729.n441 a_50751_n19729.n440 0.97759
R51261 a_50751_n19729.n442 a_50751_n19729.n438 0.97759
R51262 a_50751_n19729.n160 a_50751_n19729.n488 0.97759
R51263 a_50751_n19729.n162 a_50751_n19729.n486 0.97759
R51264 a_50751_n19729.n487 a_50751_n19729.n163 0.97759
R51265 a_50751_n19729.n164 a_50751_n19729.n485 0.97759
R51266 a_50751_n19729.n165 a_50751_n19729.n484 0.97759
R51267 a_50751_n19729.n166 a_50751_n19729.n482 0.97759
R51268 a_50751_n19729.n483 a_50751_n19729.n167 0.97759
R51269 a_50751_n19729.n168 a_50751_n19729.n481 0.97759
R51270 a_50751_n19729.n169 a_50751_n19729.n480 0.97759
R51271 a_50751_n19729.n171 a_50751_n19729.n478 0.97759
R51272 a_50751_n19729.n479 a_50751_n19729.n172 0.97759
R51273 a_50751_n19729.n173 a_50751_n19729.n477 0.97759
R51274 a_50751_n19729.n448 a_50751_n19729.n174 0.97759
R51275 a_50751_n19729.n175 a_50751_n19729.n446 0.97759
R51276 a_50751_n19729.n176 a_50751_n19729.n449 0.97759
R51277 a_50751_n19729.n177 a_50751_n19729.n447 0.97759
R51278 a_50751_n19729.n456 a_50751_n19729.n178 0.97759
R51279 a_50751_n19729.n179 a_50751_n19729.n454 0.97759
R51280 a_50751_n19729.n180 a_50751_n19729.n457 0.97759
R51281 a_50751_n19729.n182 a_50751_n19729.n455 0.97759
R51282 a_50751_n19729.n183 a_50751_n19729.n467 0.97759
R51283 a_50751_n19729.n185 a_50751_n19729.n465 0.97759
R51284 a_50751_n19729.n466 a_50751_n19729.n186 0.97759
R51285 a_50751_n19729.n187 a_50751_n19729.n464 0.97759
R51286 a_50751_n19729.n462 a_50751_n19729.n461 0.97759
R51287 a_50751_n19729.n463 a_50751_n19729.n459 0.97759
R51288 a_50751_n19729.n418 a_50751_n19729.n188 0.97759
R51289 a_50751_n19729.n189 a_50751_n19729.n416 0.97759
R51290 a_50751_n19729.n190 a_50751_n19729.n419 0.97759
R51291 a_50751_n19729.n191 a_50751_n19729.n417 0.97759
R51292 a_50751_n19729.n192 a_50751_n19729.n432 0.97759
R51293 a_50751_n19729.n193 a_50751_n19729.n430 0.97759
R51294 a_50751_n19729.n431 a_50751_n19729.n194 0.97759
R51295 a_50751_n19729.n195 a_50751_n19729.n429 0.97759
R51296 a_50751_n19729.n196 a_50751_n19729.n453 0.97759
R51297 a_50751_n19729.n197 a_50751_n19729.n451 0.97759
R51298 a_50751_n19729.n452 a_50751_n19729.n198 0.97759
R51299 a_50751_n19729.n199 a_50751_n19729.n450 0.97759
R51300 a_50751_n19729.n470 a_50751_n19729.n200 0.97759
R51301 a_50751_n19729.n201 a_50751_n19729.n468 0.97759
R51302 a_50751_n19729.n202 a_50751_n19729.n471 0.97759
R51303 a_50751_n19729.n203 a_50751_n19729.n469 0.97759
R51304 a_50751_n19729.n204 a_50751_n19729.n264 0.97759
R51305 a_50751_n19729.n205 a_50751_n19729.n262 0.97759
R51306 a_50751_n19729.n263 a_50751_n19729.n206 0.97759
R51307 a_50751_n19729.n207 a_50751_n19729.n261 0.97759
R51308 a_50751_n19729.n281 a_50751_n19729.n208 0.97759
R51309 a_50751_n19729.n209 a_50751_n19729.n279 0.97759
R51310 a_50751_n19729.n210 a_50751_n19729.n282 0.97759
R51311 a_50751_n19729.n211 a_50751_n19729.n280 0.97759
R51312 a_50751_n19729.n494 a_50751_n19729.n212 0.931516
R51313 a_50751_n19729.n213 a_50751_n19729.n492 0.931516
R51314 a_50751_n19729.n271 a_50751_n19729.n214 0.931516
R51315 a_50751_n19729.n215 a_50751_n19729.n269 0.931516
R51316 a_50751_n19729.n344 a_50751_n19729.n216 0.931516
R51317 a_50751_n19729.n217 a_50751_n19729.n342 0.931516
R51318 a_50751_n19729.n365 a_50751_n19729.n218 0.931516
R51319 a_50751_n19729.n219 a_50751_n19729.n363 0.931516
R51320 a_50751_n19729.n439 a_50751_n19729.n220 0.931516
R51321 a_50751_n19729.n221 a_50751_n19729.n437 0.931516
R51322 a_50751_n19729.n460 a_50751_n19729.n222 0.931516
R51323 a_50751_n19729.n223 a_50751_n19729.n458 0.931516
R51324 a_50751_n19729.n113 a_50751_n19729.n110 0.82023
R51325 a_50751_n19729.n184 a_50751_n19729.n181 0.82023
R51326 a_50751_n19729.n50 a_50751_n19729.n47 0.82023
R51327 a_50751_n19729.n68 a_50751_n19729.n75 0.818405
R51328 a_50751_n19729.n139 a_50751_n19729.n146 0.818405
R51329 a_50751_n19729.n19 a_50751_n19729.n6 0.818405
R51330 a_50751_n19729.n490 a_50751_n19729.n489 0.7505
R51331 a_50751_n19729.n395 a_50751_n19729.n394 0.7505
R51332 a_50751_n19729.n394 a_50751_n19729.n90 0.717155
R51333 a_50751_n19729.n489 a_50751_n19729.n161 0.717155
R51334 a_50751_n19729.n491 a_50751_n19729.n27 0.717155
R51335 a_50751_n19729.n87 a_50751_n19729.n80 0.639622
R51336 a_50751_n19729.n158 a_50751_n19729.n151 0.639622
R51337 a_50751_n19729.n224 a_50751_n19729.n22 0.639622
R51338 a_50751_n19729.n497 a_50751_n19729.n496 0.62434
R51339 a_50751_n19729.n274 a_50751_n19729.n273 0.62434
R51340 a_50751_n19729.n347 a_50751_n19729.n346 0.62434
R51341 a_50751_n19729.n368 a_50751_n19729.n367 0.62434
R51342 a_50751_n19729.n442 a_50751_n19729.n441 0.62434
R51343 a_50751_n19729.n463 a_50751_n19729.n462 0.62434
R51344 a_50751_n19729.n211 a_50751_n19729.n210 0.62434
R51345 a_50751_n19729.n209 a_50751_n19729.n208 0.62434
R51346 a_50751_n19729.n207 a_50751_n19729.n206 0.62434
R51347 a_50751_n19729.n205 a_50751_n19729.n204 0.62434
R51348 a_50751_n19729.n203 a_50751_n19729.n202 0.62434
R51349 a_50751_n19729.n201 a_50751_n19729.n200 0.62434
R51350 a_50751_n19729.n199 a_50751_n19729.n198 0.62434
R51351 a_50751_n19729.n197 a_50751_n19729.n196 0.62434
R51352 a_50751_n19729.n195 a_50751_n19729.n194 0.62434
R51353 a_50751_n19729.n193 a_50751_n19729.n192 0.62434
R51354 a_50751_n19729.n191 a_50751_n19729.n190 0.62434
R51355 a_50751_n19729.n189 a_50751_n19729.n188 0.62434
R51356 a_50751_n19729.n187 a_50751_n19729.n186 0.62434
R51357 a_50751_n19729.n185 a_50751_n19729.n183 0.62434
R51358 a_50751_n19729.n182 a_50751_n19729.n180 0.62434
R51359 a_50751_n19729.n179 a_50751_n19729.n178 0.62434
R51360 a_50751_n19729.n177 a_50751_n19729.n176 0.62434
R51361 a_50751_n19729.n175 a_50751_n19729.n174 0.62434
R51362 a_50751_n19729.n173 a_50751_n19729.n172 0.62434
R51363 a_50751_n19729.n171 a_50751_n19729.n169 0.62434
R51364 a_50751_n19729.n168 a_50751_n19729.n167 0.62434
R51365 a_50751_n19729.n166 a_50751_n19729.n165 0.62434
R51366 a_50751_n19729.n164 a_50751_n19729.n163 0.62434
R51367 a_50751_n19729.n162 a_50751_n19729.n160 0.62434
R51368 a_50751_n19729.n159 a_50751_n19729.n157 0.62434
R51369 a_50751_n19729.n156 a_50751_n19729.n155 0.62434
R51370 a_50751_n19729.n154 a_50751_n19729.n153 0.62434
R51371 a_50751_n19729.n152 a_50751_n19729.n150 0.62434
R51372 a_50751_n19729.n149 a_50751_n19729.n148 0.62434
R51373 a_50751_n19729.n147 a_50751_n19729.n145 0.62434
R51374 a_50751_n19729.n144 a_50751_n19729.n143 0.62434
R51375 a_50751_n19729.n142 a_50751_n19729.n141 0.62434
R51376 a_50751_n19729.n140 a_50751_n19729.n138 0.62434
R51377 a_50751_n19729.n137 a_50751_n19729.n136 0.62434
R51378 a_50751_n19729.n399 a_50751_n19729.n135 0.62434
R51379 a_50751_n19729.n134 a_50751_n19729.n133 0.62434
R51380 a_50751_n19729.n132 a_50751_n19729.n131 0.62434
R51381 a_50751_n19729.n130 a_50751_n19729.n129 0.62434
R51382 a_50751_n19729.n128 a_50751_n19729.n127 0.62434
R51383 a_50751_n19729.n126 a_50751_n19729.n125 0.62434
R51384 a_50751_n19729.n124 a_50751_n19729.n123 0.62434
R51385 a_50751_n19729.n122 a_50751_n19729.n121 0.62434
R51386 a_50751_n19729.n120 a_50751_n19729.n119 0.62434
R51387 a_50751_n19729.n118 a_50751_n19729.n117 0.62434
R51388 a_50751_n19729.n116 a_50751_n19729.n115 0.62434
R51389 a_50751_n19729.n114 a_50751_n19729.n112 0.62434
R51390 a_50751_n19729.n111 a_50751_n19729.n109 0.62434
R51391 a_50751_n19729.n108 a_50751_n19729.n107 0.62434
R51392 a_50751_n19729.n106 a_50751_n19729.n105 0.62434
R51393 a_50751_n19729.n104 a_50751_n19729.n103 0.62434
R51394 a_50751_n19729.n102 a_50751_n19729.n101 0.62434
R51395 a_50751_n19729.n100 a_50751_n19729.n98 0.62434
R51396 a_50751_n19729.n97 a_50751_n19729.n96 0.62434
R51397 a_50751_n19729.n95 a_50751_n19729.n94 0.62434
R51398 a_50751_n19729.n93 a_50751_n19729.n92 0.62434
R51399 a_50751_n19729.n91 a_50751_n19729.n89 0.62434
R51400 a_50751_n19729.n88 a_50751_n19729.n86 0.62434
R51401 a_50751_n19729.n85 a_50751_n19729.n84 0.62434
R51402 a_50751_n19729.n83 a_50751_n19729.n82 0.62434
R51403 a_50751_n19729.n81 a_50751_n19729.n79 0.62434
R51404 a_50751_n19729.n78 a_50751_n19729.n77 0.62434
R51405 a_50751_n19729.n76 a_50751_n19729.n74 0.62434
R51406 a_50751_n19729.n73 a_50751_n19729.n72 0.62434
R51407 a_50751_n19729.n71 a_50751_n19729.n70 0.62434
R51408 a_50751_n19729.n69 a_50751_n19729.n67 0.62434
R51409 a_50751_n19729.n66 a_50751_n19729.n65 0.62434
R51410 a_50751_n19729.n304 a_50751_n19729.n64 0.62434
R51411 a_50751_n19729.n63 a_50751_n19729.n62 0.62434
R51412 a_50751_n19729.n61 a_50751_n19729.n60 0.62434
R51413 a_50751_n19729.n59 a_50751_n19729.n58 0.62434
R51414 a_50751_n19729.n57 a_50751_n19729.n56 0.62434
R51415 a_50751_n19729.n55 a_50751_n19729.n54 0.62434
R51416 a_50751_n19729.n53 a_50751_n19729.n52 0.62434
R51417 a_50751_n19729.n51 a_50751_n19729.n49 0.62434
R51418 a_50751_n19729.n48 a_50751_n19729.n46 0.62434
R51419 a_50751_n19729.n45 a_50751_n19729.n44 0.62434
R51420 a_50751_n19729.n43 a_50751_n19729.n42 0.62434
R51421 a_50751_n19729.n41 a_50751_n19729.n40 0.62434
R51422 a_50751_n19729.n39 a_50751_n19729.n38 0.62434
R51423 a_50751_n19729.n37 a_50751_n19729.n35 0.62434
R51424 a_50751_n19729.n34 a_50751_n19729.n33 0.62434
R51425 a_50751_n19729.n32 a_50751_n19729.n31 0.62434
R51426 a_50751_n19729.n30 a_50751_n19729.n29 0.62434
R51427 a_50751_n19729.n28 a_50751_n19729.n26 0.62434
R51428 a_50751_n19729.n25 a_50751_n19729.n24 0.62434
R51429 a_50751_n19729.n23 a_50751_n19729.n21 0.62434
R51430 a_50751_n19729.n20 a_50751_n19729.n18 0.62434
R51431 a_50751_n19729.n17 a_50751_n19729.n16 0.62434
R51432 a_50751_n19729.n15 a_50751_n19729.n14 0.62434
R51433 a_50751_n19729.n13 a_50751_n19729.n12 0.62434
R51434 a_50751_n19729.n11 a_50751_n19729.n10 0.62434
R51435 a_50751_n19729.n9 a_50751_n19729.n8 0.62434
R51436 a_50751_n19729.n7 a_50751_n19729.n5 0.62434
R51437 a_50751_n19729.n4 a_50751_n19729.n3 0.62434
R51438 a_50751_n19729.n229 a_50751_n19729.n2 0.62434
R51439 a_50751_n19729.n1 a_50751_n19729.n0 0.62434
R51440 a_50751_n19729.n394 a_50751_n19729.n87 0.617426
R51441 a_50751_n19729.n489 a_50751_n19729.n158 0.617426
R51442 a_50751_n19729.n22 a_50751_n19729.n491 0.617426
R51443 a_50751_n19729.n223 a_50751_n19729.n222 0.595087
R51444 a_50751_n19729.n221 a_50751_n19729.n220 0.595087
R51445 a_50751_n19729.n219 a_50751_n19729.n218 0.595087
R51446 a_50751_n19729.n217 a_50751_n19729.n216 0.595087
R51447 a_50751_n19729.n215 a_50751_n19729.n214 0.595087
R51448 a_50751_n19729.n213 a_50751_n19729.n212 0.595087
R51449 a_50751_n19729.n75 a_50751_n19729.n80 0.545973
R51450 a_50751_n19729.n146 a_50751_n19729.n151 0.545973
R51451 a_50751_n19729.n224 a_50751_n19729.n19 0.545973
R51452 a_50751_n19729.n110 a_50751_n19729.n99 0.545365
R51453 a_50751_n19729.n181 a_50751_n19729.n170 0.545365
R51454 a_50751_n19729.n47 a_50751_n19729.n36 0.545365
R51455 a_50751_n19729.n27 a_50751_n19729.n36 0.452324
R51456 a_50751_n19729.n161 a_50751_n19729.n170 0.452324
R51457 a_50751_n19729.n90 a_50751_n19729.n99 0.452324
R51458 a_65486_n36322.n0 a_65486_n36322.t18 13.7934
R51459 a_65486_n36322.n2 a_65486_n36322.t3 10.7024
R51460 a_65486_n36322.n2 a_65486_n36322.t4 10.1668
R51461 a_65486_n36322.n2 a_65486_n36322.t5 9.64458
R51462 a_65486_n36322.n2 a_65486_n36322.t1 9.27635
R51463 a_65486_n36322.n2 a_65486_n36322.n0 8.75198
R51464 a_65486_n36322.n0 a_65486_n36322.t17 8.14051
R51465 a_65486_n36322.n0 a_65486_n36322.t15 8.14051
R51466 a_65486_n36322.n0 a_65486_n36322.t23 8.14051
R51467 a_65486_n36322.n0 a_65486_n36322.t8 8.14051
R51468 a_65486_n36322.n0 a_65486_n36322.t21 8.06917
R51469 a_65486_n36322.n0 a_65486_n36322.t12 8.06917
R51470 a_65486_n36322.n0 a_65486_n36322.t10 8.06917
R51471 a_65486_n36322.n0 a_65486_n36322.t11 8.06917
R51472 a_65486_n36322.n0 a_65486_n36322.t9 8.06917
R51473 a_65486_n36322.n0 a_65486_n36322.t16 8.06917
R51474 a_65486_n36322.n0 a_65486_n36322.t19 8.06917
R51475 a_65486_n36322.n1 a_65486_n36322.t7 7.94157
R51476 a_65486_n36322.n2 a_65486_n36322.t2 7.72643
R51477 a_65486_n36322.n1 a_65486_n36322.t6 7.22925
R51478 a_65486_n36322.t0 a_65486_n36322.n2 7.17912
R51479 a_65486_n36322.n0 a_65486_n36322.t14 8.33554
R51480 a_65486_n36322.t13 a_65486_n36322.n0 8.33554
R51481 a_65486_n36322.n0 a_65486_n36322.t20 8.33647
R51482 a_65486_n36322.t22 a_65486_n36322.n0 8.33647
R51483 a_65486_n36322.n2 a_65486_n36322.n1 7.46075
R51484 a_71342_n30339.n0 a_71342_n30339.t1 10.3838
R51485 a_71342_n30339.n0 a_71342_n30339.t3 10.3566
R51486 a_71342_n30339.n0 a_71342_n30339.t2 10.0407
R51487 a_71342_n30339.t0 a_71342_n30339.n0 9.57605
R51488 a_106809_n17715.t0 a_106809_n17715.t1 12.8114
R51489 a_33249_48695.n109 a_33249_48695.n106 7.94229
R51490 a_33249_48695.n140 a_33249_48695.n137 7.94229
R51491 a_33249_48695.n394 a_33249_48695.n393 7.22198
R51492 a_33249_48695.n364 a_33249_48695.n363 7.22198
R51493 a_33249_48695.n68 a_33249_48695.t315 6.77653
R51494 a_33249_48695.n47 a_33249_48695.t242 6.77653
R51495 a_33249_48695.n64 a_33249_48695.t176 6.7761
R51496 a_33249_48695.n377 a_33249_48695.t251 6.7761
R51497 a_33249_48695.n9 a_33249_48695.t255 6.77231
R51498 a_33249_48695.n19 a_33249_48695.t203 6.77231
R51499 a_33249_48695.n267 a_33249_48695.t46 6.58663
R51500 a_33249_48695.n223 a_33249_48695.t48 6.58663
R51501 a_33249_48695.n335 a_33249_48695.n334 6.50088
R51502 a_33249_48695.n300 a_33249_48695.n296 6.50088
R51503 a_33249_48695.n268 a_33249_48695.n265 5.95439
R51504 a_33249_48695.n224 a_33249_48695.n221 5.95439
R51505 a_33249_48695.n108 a_33249_48695.t306 5.69423
R51506 a_33249_48695.n90 a_33249_48695.t289 5.69423
R51507 a_33249_48695.n139 a_33249_48695.t199 5.69423
R51508 a_33249_48695.n135 a_33249_48695.t184 5.69423
R51509 a_33249_48695.n61 a_33249_48695.t325 5.50607
R51510 a_33249_48695.n48 a_33249_48695.t264 5.50607
R51511 a_33249_48695.n374 a_33249_48695.t222 5.50607
R51512 a_33249_48695.n69 a_33249_48695.t165 5.50607
R51513 a_33249_48695.n62 a_33249_48695.t213 5.50475
R51514 a_33249_48695.n58 a_33249_48695.t317 5.50475
R51515 a_33249_48695.n57 a_33249_48695.t161 5.50475
R51516 a_33249_48695.n375 a_33249_48695.t287 5.50475
R51517 a_33249_48695.n371 a_33249_48695.t212 5.50475
R51518 a_33249_48695.n370 a_33249_48695.t235 5.50475
R51519 a_33249_48695.n70 a_33249_48695.t227 5.50475
R51520 a_33249_48695.t332 a_33249_48695.n397 5.50475
R51521 a_33249_48695.n108 a_33249_48695.n107 5.49558
R51522 a_33249_48695.n139 a_33249_48695.n138 5.49558
R51523 a_33249_48695.n265 a_33249_48695.t63 5.31528
R51524 a_33249_48695.n221 a_33249_48695.t71 5.31528
R51525 a_33249_48695.n80 a_33249_48695.n78 4.92758
R51526 a_33249_48695.n306 a_33249_48695.n304 4.92758
R51527 a_33249_48695.n38 a_33249_48695.n273 4.92217
R51528 a_33249_48695.n45 a_33249_48695.n286 4.92217
R51529 a_33249_48695.n26 a_33249_48695.n88 4.22068
R51530 a_33249_48695.n27 a_33249_48695.t268 5.69068
R51531 a_33249_48695.n28 a_33249_48695.n87 4.22068
R51532 a_33249_48695.n29 a_33249_48695.n131 4.22068
R51533 a_33249_48695.n30 a_33249_48695.t324 5.69068
R51534 a_33249_48695.n31 a_33249_48695.n130 4.22068
R51535 a_33249_48695.n21 a_33249_48695.n184 3.84173
R51536 a_33249_48695.n24 a_33249_48695.n180 3.84173
R51537 a_33249_48695.n32 a_33249_48695.n280 3.65107
R51538 a_33249_48695.n33 a_33249_48695.n279 3.65107
R51539 a_33249_48695.n34 a_33249_48695.n278 3.65107
R51540 a_33249_48695.n35 a_33249_48695.n277 3.65107
R51541 a_33249_48695.n276 a_33249_48695.n36 3.65107
R51542 a_33249_48695.n275 a_33249_48695.n37 3.65107
R51543 a_33249_48695.n274 a_33249_48695.n38 3.65107
R51544 a_33249_48695.n39 a_33249_48695.n293 3.65107
R51545 a_33249_48695.n40 a_33249_48695.n292 3.65107
R51546 a_33249_48695.n41 a_33249_48695.n291 3.65107
R51547 a_33249_48695.n42 a_33249_48695.n290 3.65107
R51548 a_33249_48695.n289 a_33249_48695.n43 3.65107
R51549 a_33249_48695.n288 a_33249_48695.n44 3.65107
R51550 a_33249_48695.n287 a_33249_48695.n45 3.65107
R51551 a_33249_48695.n0 a_33249_48695.n384 4.0312
R51552 a_33249_48695.t228 a_33249_48695.n1 5.5012
R51553 a_33249_48695.t160 a_33249_48695.n2 5.5012
R51554 a_33249_48695.n383 a_33249_48695.n3 4.0312
R51555 a_33249_48695.t331 a_33249_48695.n4 5.5012
R51556 a_33249_48695.t173 a_33249_48695.n5 5.5012
R51557 a_33249_48695.n382 a_33249_48695.n6 4.0312
R51558 a_33249_48695.t168 a_33249_48695.n7 5.5012
R51559 a_33249_48695.t279 a_33249_48695.n8 5.5012
R51560 a_33249_48695.n380 a_33249_48695.n9 4.0312
R51561 a_33249_48695.n10 a_33249_48695.n75 4.0312
R51562 a_33249_48695.n11 a_33249_48695.t178 5.5012
R51563 a_33249_48695.n12 a_33249_48695.t282 5.5012
R51564 a_33249_48695.n13 a_33249_48695.n74 4.0312
R51565 a_33249_48695.n14 a_33249_48695.t278 5.5012
R51566 a_33249_48695.n15 a_33249_48695.t297 5.5012
R51567 a_33249_48695.n16 a_33249_48695.n73 4.0312
R51568 a_33249_48695.t293 a_33249_48695.n17 5.5012
R51569 a_33249_48695.t229 a_33249_48695.n18 5.5012
R51570 a_33249_48695.n72 a_33249_48695.n19 4.0312
R51571 a_33249_48695.n20 a_33249_48695.t85 5.31173
R51572 a_33249_48695.n22 a_33249_48695.t91 5.31173
R51573 a_33249_48695.n23 a_33249_48695.t80 5.31173
R51574 a_33249_48695.n25 a_33249_48695.t83 5.31173
R51575 a_33249_48695.n264 a_33249_48695.n262 4.50663
R51576 a_33249_48695.n220 a_33249_48695.n179 4.50663
R51577 a_33249_48695.n185 a_33249_48695.n22 4.46113
R51578 a_33249_48695.n392 a_33249_48695.t158 4.24002
R51579 a_33249_48695.n52 a_33249_48695.t318 4.24002
R51580 a_33249_48695.n362 a_33249_48695.t280 4.24002
R51581 a_33249_48695.n353 a_33249_48695.t263 4.24002
R51582 a_33249_48695.n106 a_33249_48695.n105 4.22423
R51583 a_33249_48695.n137 a_33249_48695.n136 4.22423
R51584 a_33249_48695.n301 a_33249_48695.t350 4.06712
R51585 a_33249_48695.n284 a_33249_48695.t130 4.06712
R51586 a_33249_48695.n329 a_33249_48695.t345 4.06712
R51587 a_33249_48695.n327 a_33249_48695.t125 4.06712
R51588 a_33249_48695.n96 a_33249_48695.t205 4.05054
R51589 a_33249_48695.n101 a_33249_48695.t244 4.05054
R51590 a_33249_48695.n103 a_33249_48695.t175 4.05054
R51591 a_33249_48695.n116 a_33249_48695.t170 4.05054
R51592 a_33249_48695.n118 a_33249_48695.t187 4.05054
R51593 a_33249_48695.n124 a_33249_48695.t182 4.05054
R51594 a_33249_48695.n126 a_33249_48695.t296 4.05054
R51595 a_33249_48695.n91 a_33249_48695.t267 4.05054
R51596 a_33249_48695.n164 a_33249_48695.t328 4.05054
R51597 a_33249_48695.n169 a_33249_48695.t192 4.05054
R51598 a_33249_48695.n171 a_33249_48695.t300 4.05054
R51599 a_33249_48695.n158 a_33249_48695.t295 4.05054
R51600 a_33249_48695.n156 a_33249_48695.t312 4.05054
R51601 a_33249_48695.n150 a_33249_48695.t309 4.05054
R51602 a_33249_48695.n148 a_33249_48695.t246 4.05054
R51603 a_33249_48695.n142 a_33249_48695.t221 4.05054
R51604 a_33249_48695.n64 a_33249_48695.n63 4.03475
R51605 a_33249_48695.n60 a_33249_48695.n59 4.03475
R51606 a_33249_48695.n50 a_33249_48695.n49 4.03475
R51607 a_33249_48695.n47 a_33249_48695.n46 4.03475
R51608 a_33249_48695.n377 a_33249_48695.n376 4.03475
R51609 a_33249_48695.n373 a_33249_48695.n372 4.03475
R51610 a_33249_48695.n369 a_33249_48695.n368 4.03475
R51611 a_33249_48695.n68 a_33249_48695.n67 4.03475
R51612 a_33249_48695.n330 a_33249_48695.n77 3.96014
R51613 a_33249_48695.n303 a_33249_48695.n302 3.96014
R51614 a_33249_48695.n96 a_33249_48695.t163 3.87765
R51615 a_33249_48695.n101 a_33249_48695.t197 3.87765
R51616 a_33249_48695.n103 a_33249_48695.t308 3.87765
R51617 a_33249_48695.n116 a_33249_48695.t302 3.87765
R51618 a_33249_48695.n118 a_33249_48695.t321 3.87765
R51619 a_33249_48695.n124 a_33249_48695.t316 3.87765
R51620 a_33249_48695.n126 a_33249_48695.t254 3.87765
R51621 a_33249_48695.n91 a_33249_48695.t225 3.87765
R51622 a_33249_48695.n164 a_33249_48695.t237 3.87765
R51623 a_33249_48695.n169 a_33249_48695.t270 3.87765
R51624 a_33249_48695.n171 a_33249_48695.t204 3.87765
R51625 a_33249_48695.n158 a_33249_48695.t196 3.87765
R51626 a_33249_48695.n156 a_33249_48695.t216 3.87765
R51627 a_33249_48695.n150 a_33249_48695.t210 3.87765
R51628 a_33249_48695.n148 a_33249_48695.t326 3.87765
R51629 a_33249_48695.n142 a_33249_48695.t299 3.87765
R51630 a_33249_48695.n301 a_33249_48695.t349 3.86107
R51631 a_33249_48695.n284 a_33249_48695.t128 3.86107
R51632 a_33249_48695.n329 a_33249_48695.t17 3.86107
R51633 a_33249_48695.n327 a_33249_48695.t11 3.86107
R51634 a_33249_48695.n267 a_33249_48695.n266 3.84528
R51635 a_33249_48695.n264 a_33249_48695.n263 3.84528
R51636 a_33249_48695.n223 a_33249_48695.n222 3.84528
R51637 a_33249_48695.n220 a_33249_48695.n219 3.84528
R51638 a_33249_48695.n256 a_33249_48695.n252 3.79678
R51639 a_33249_48695.n239 a_33249_48695.n235 3.79678
R51640 a_33249_48695.n197 a_33249_48695.n193 3.79678
R51641 a_33249_48695.n212 a_33249_48695.n208 3.79678
R51642 a_33249_48695.n82 a_33249_48695.n80 3.79678
R51643 a_33249_48695.n344 a_33249_48695.n342 3.79678
R51644 a_33249_48695.n308 a_33249_48695.n306 3.79678
R51645 a_33249_48695.n317 a_33249_48695.n315 3.79678
R51646 a_33249_48695.n228 a_33249_48695.n25 3.87644
R51647 a_33249_48695.n248 a_33249_48695.n244 3.73034
R51648 a_33249_48695.n217 a_33249_48695.n201 3.73034
R51649 a_33249_48695.n392 a_33249_48695.t290 3.68818
R51650 a_33249_48695.n52 a_33249_48695.t272 3.68818
R51651 a_33249_48695.n362 a_33249_48695.t185 3.68818
R51652 a_33249_48695.n353 a_33249_48695.t171 3.68818
R51653 a_33249_48695.n346 a_33249_48695.n345 3.65581
R51654 a_33249_48695.n344 a_33249_48695.n343 3.65581
R51655 a_33249_48695.n342 a_33249_48695.n341 3.65581
R51656 a_33249_48695.n340 a_33249_48695.n339 3.65581
R51657 a_33249_48695.n84 a_33249_48695.n83 3.65581
R51658 a_33249_48695.n82 a_33249_48695.n81 3.65581
R51659 a_33249_48695.n80 a_33249_48695.n79 3.65581
R51660 a_33249_48695.n319 a_33249_48695.n318 3.65581
R51661 a_33249_48695.n317 a_33249_48695.n316 3.65581
R51662 a_33249_48695.n315 a_33249_48695.n314 3.65581
R51663 a_33249_48695.n313 a_33249_48695.n312 3.65581
R51664 a_33249_48695.n310 a_33249_48695.n309 3.65581
R51665 a_33249_48695.n308 a_33249_48695.n307 3.65581
R51666 a_33249_48695.n306 a_33249_48695.n305 3.65581
R51667 a_33249_48695.n340 a_33249_48695.n338 3.64443
R51668 a_33249_48695.n313 a_33249_48695.n311 3.64443
R51669 a_33249_48695.n322 a_33249_48695.n35 3.64223
R51670 a_33249_48695.n294 a_33249_48695.n42 3.64223
R51671 a_33249_48695.n129 a_33249_48695.n90 3.25667
R51672 a_33249_48695.n391 a_33249_48695.n387 3.23904
R51673 a_33249_48695.n361 a_33249_48695.n66 3.23904
R51674 a_33249_48695.n133 a_33249_48695.n31 3.15553
R51675 a_33249_48695.n177 a_33249_48695.n28 3.15553
R51676 a_33249_48695.n268 a_33249_48695.n267 3.00663
R51677 a_33249_48695.n224 a_33249_48695.n223 3.00663
R51678 a_33249_48695.n231 a_33249_48695.n229 2.7866
R51679 a_33249_48695.n234 a_33249_48695.n232 2.7866
R51680 a_33249_48695.n238 a_33249_48695.n236 2.7866
R51681 a_33249_48695.n242 a_33249_48695.n240 2.7866
R51682 a_33249_48695.n247 a_33249_48695.n245 2.7866
R51683 a_33249_48695.n251 a_33249_48695.n249 2.7866
R51684 a_33249_48695.n255 a_33249_48695.n253 2.7866
R51685 a_33249_48695.n259 a_33249_48695.n257 2.7866
R51686 a_33249_48695.n204 a_33249_48695.n202 2.7866
R51687 a_33249_48695.n207 a_33249_48695.n205 2.7866
R51688 a_33249_48695.n211 a_33249_48695.n209 2.7866
R51689 a_33249_48695.n215 a_33249_48695.n213 2.7866
R51690 a_33249_48695.n200 a_33249_48695.n198 2.7866
R51691 a_33249_48695.n196 a_33249_48695.n194 2.7866
R51692 a_33249_48695.n192 a_33249_48695.n190 2.7866
R51693 a_33249_48695.n188 a_33249_48695.n186 2.7866
R51694 a_33249_48695.n390 a_33249_48695.n389 2.77002
R51695 a_33249_48695.n55 a_33249_48695.n54 2.77002
R51696 a_33249_48695.n360 a_33249_48695.n359 2.77002
R51697 a_33249_48695.n356 a_33249_48695.n355 2.77002
R51698 a_33249_48695.n56 a_33249_48695.n52 2.73714
R51699 a_33249_48695.n357 a_33249_48695.n353 2.73714
R51700 a_33249_48695.n95 a_33249_48695.n91 2.73714
R51701 a_33249_48695.n146 a_33249_48695.n142 2.73714
R51702 a_33249_48695.n328 a_33249_48695.n326 2.73714
R51703 a_33249_48695.n285 a_33249_48695.n283 2.73714
R51704 a_33249_48695.n235 a_33249_48695.n231 2.73672
R51705 a_33249_48695.n208 a_33249_48695.n204 2.73672
R51706 a_33249_48695.n100 a_33249_48695.n96 2.73672
R51707 a_33249_48695.n168 a_33249_48695.n164 2.73672
R51708 a_33249_48695.n371 a_33249_48695.n370 2.60203
R51709 a_33249_48695.n119 a_33249_48695.n117 2.60203
R51710 a_33249_48695.n159 a_33249_48695.n157 2.60203
R51711 a_33249_48695.n58 a_33249_48695.n57 2.60203
R51712 a_33249_48695.n299 a_33249_48695.n297 2.59712
R51713 a_33249_48695.n283 a_33249_48695.n281 2.59712
R51714 a_33249_48695.n333 a_33249_48695.n331 2.59712
R51715 a_33249_48695.n326 a_33249_48695.n324 2.59712
R51716 a_33249_48695.n99 a_33249_48695.n98 2.58054
R51717 a_33249_48695.n114 a_33249_48695.n113 2.58054
R51718 a_33249_48695.n122 a_33249_48695.n121 2.58054
R51719 a_33249_48695.n94 a_33249_48695.n93 2.58054
R51720 a_33249_48695.n167 a_33249_48695.n166 2.58054
R51721 a_33249_48695.n162 a_33249_48695.n161 2.58054
R51722 a_33249_48695.n154 a_33249_48695.n153 2.58054
R51723 a_33249_48695.n145 a_33249_48695.n144 2.58054
R51724 a_33249_48695.n127 a_33249_48695.n125 2.53418
R51725 a_33249_48695.n104 a_33249_48695.n102 2.53418
R51726 a_33249_48695.n151 a_33249_48695.n149 2.53418
R51727 a_33249_48695.n172 a_33249_48695.n170 2.53418
R51728 a_33249_48695.n397 a_33249_48695.n48 2.52471
R51729 a_33249_48695.n70 a_33249_48695.n69 2.52436
R51730 a_33249_48695.n375 a_33249_48695.n374 2.52436
R51731 a_33249_48695.n62 a_33249_48695.n61 2.52436
R51732 a_33249_48695.n135 a_33249_48695.n134 2.51873
R51733 a_33249_48695.n335 a_33249_48695.n328 2.46014
R51734 a_33249_48695.n296 a_33249_48695.n285 2.46014
R51735 a_33249_48695.n99 a_33249_48695.n97 2.40765
R51736 a_33249_48695.n114 a_33249_48695.n112 2.40765
R51737 a_33249_48695.n122 a_33249_48695.n120 2.40765
R51738 a_33249_48695.n94 a_33249_48695.n92 2.40765
R51739 a_33249_48695.n167 a_33249_48695.n165 2.40765
R51740 a_33249_48695.n162 a_33249_48695.n160 2.40765
R51741 a_33249_48695.n154 a_33249_48695.n152 2.40765
R51742 a_33249_48695.n145 a_33249_48695.n143 2.40765
R51743 a_33249_48695.n299 a_33249_48695.n298 2.39107
R51744 a_33249_48695.n283 a_33249_48695.n282 2.39107
R51745 a_33249_48695.n333 a_33249_48695.n332 2.39107
R51746 a_33249_48695.n326 a_33249_48695.n325 2.39107
R51747 a_33249_48695.n227 a_33249_48695.n23 2.37644
R51748 a_33249_48695.n183 a_33249_48695.n20 2.37644
R51749 a_33249_48695.n110 a_33249_48695.n109 2.23844
R51750 a_33249_48695.n390 a_33249_48695.n388 2.21818
R51751 a_33249_48695.n55 a_33249_48695.n53 2.21818
R51752 a_33249_48695.n360 a_33249_48695.n358 2.21818
R51753 a_33249_48695.n356 a_33249_48695.n354 2.21818
R51754 a_33249_48695.n231 a_33249_48695.n230 2.2016
R51755 a_33249_48695.n234 a_33249_48695.n233 2.2016
R51756 a_33249_48695.n238 a_33249_48695.n237 2.2016
R51757 a_33249_48695.n242 a_33249_48695.n241 2.2016
R51758 a_33249_48695.n247 a_33249_48695.n246 2.2016
R51759 a_33249_48695.n251 a_33249_48695.n250 2.2016
R51760 a_33249_48695.n255 a_33249_48695.n254 2.2016
R51761 a_33249_48695.n259 a_33249_48695.n258 2.2016
R51762 a_33249_48695.n204 a_33249_48695.n203 2.2016
R51763 a_33249_48695.n207 a_33249_48695.n206 2.2016
R51764 a_33249_48695.n211 a_33249_48695.n210 2.2016
R51765 a_33249_48695.n215 a_33249_48695.n214 2.2016
R51766 a_33249_48695.n200 a_33249_48695.n199 2.2016
R51767 a_33249_48695.n196 a_33249_48695.n195 2.2016
R51768 a_33249_48695.n192 a_33249_48695.n191 2.2016
R51769 a_33249_48695.n188 a_33249_48695.n187 2.2016
R51770 a_33249_48695.n396 a_33249_48695.n395 2.13841
R51771 a_33249_48695.n387 a_33249_48695.n65 2.13841
R51772 a_33249_48695.n218 a_33249_48695.n183 2.0852
R51773 a_33249_48695.n295 a_33249_48695.n294 2.0852
R51774 a_33249_48695.n348 a_33249_48695.n347 1.95191
R51775 a_33249_48695.n262 a_33249_48695.n178 1.90397
R51776 a_33249_48695.n348 a_33249_48695.n76 1.80854
R51777 a_33249_48695.n178 a_33249_48695.n71 1.80603
R51778 a_33249_48695.n394 a_33249_48695.n56 1.73904
R51779 a_33249_48695.n364 a_33249_48695.n357 1.73904
R51780 a_33249_48695.n347 a_33249_48695.n346 1.73609
R51781 a_33249_48695.n320 a_33249_48695.n319 1.73609
R51782 a_33249_48695.n261 a_33249_48695.n260 1.65018
R51783 a_33249_48695.n189 a_33249_48695.n185 1.65018
R51784 a_33249_48695.n271 a_33249_48695.n270 1.56167
R51785 a_33249_48695.n132 a_33249_48695.n29 1.65553
R51786 a_33249_48695.n176 a_33249_48695.n26 1.65553
R51787 a_33249_48695.n352 a_33249_48695.n351 1.5005
R51788 a_33249_48695.n365 a_33249_48695.n364 1.5005
R51789 a_33249_48695.n367 a_33249_48695.n366 1.5005
R51790 a_33249_48695.n381 a_33249_48695.n51 1.5005
R51791 a_33249_48695.n395 a_33249_48695.n394 1.5005
R51792 a_33249_48695.n225 a_33249_48695.n224 1.5005
R51793 a_33249_48695.n227 a_33249_48695.n226 1.5005
R51794 a_33249_48695.n269 a_33249_48695.n268 1.5005
R51795 a_33249_48695.n218 a_33249_48695.n217 1.5005
R51796 a_33249_48695.n244 a_33249_48695.n85 1.5005
R51797 a_33249_48695.n147 a_33249_48695.n86 1.5005
R51798 a_33249_48695.n129 a_33249_48695.n128 1.5005
R51799 a_33249_48695.n176 a_33249_48695.n175 1.5005
R51800 a_33249_48695.n174 a_33249_48695.n173 1.5005
R51801 a_33249_48695.n141 a_33249_48695.n140 1.5005
R51802 a_33249_48695.n132 a_33249_48695.n89 1.5005
R51803 a_33249_48695.n111 a_33249_48695.n110 1.5005
R51804 a_33249_48695.n336 a_33249_48695.n335 1.5005
R51805 a_33249_48695.n311 a_33249_48695.n272 1.5005
R51806 a_33249_48695.n323 a_33249_48695.n322 1.5005
R51807 a_33249_48695.n338 a_33249_48695.n337 1.5005
R51808 a_33249_48695.n296 a_33249_48695.n295 1.5005
R51809 a_33249_48695.n350 a_33249_48695.n349 1.5005
R51810 a_33249_48695.n379 a_33249_48695.n378 1.5005
R51811 a_33249_48695.n386 a_33249_48695.n385 1.5005
R51812 a_33249_48695.n63 a_33249_48695.t271 1.4705
R51813 a_33249_48695.n63 a_33249_48695.t211 1.4705
R51814 a_33249_48695.n59 a_33249_48695.t262 1.4705
R51815 a_33249_48695.n59 a_33249_48695.t206 1.4705
R51816 a_33249_48695.n49 a_33249_48695.t256 1.4705
R51817 a_33249_48695.n49 a_33249_48695.t219 1.4705
R51818 a_33249_48695.n46 a_33249_48695.t202 1.4705
R51819 a_33249_48695.n46 a_33249_48695.t322 1.4705
R51820 a_33249_48695.n388 a_33249_48695.t232 1.4705
R51821 a_33249_48695.n388 a_33249_48695.t157 1.4705
R51822 a_33249_48695.n389 a_33249_48695.t273 1.4705
R51823 a_33249_48695.n389 a_33249_48695.t198 1.4705
R51824 a_33249_48695.n53 a_33249_48695.t214 1.4705
R51825 a_33249_48695.n53 a_33249_48695.t294 1.4705
R51826 a_33249_48695.n54 a_33249_48695.t258 1.4705
R51827 a_33249_48695.n54 a_33249_48695.t164 1.4705
R51828 a_33249_48695.n384 a_33249_48695.t284 1.4705
R51829 a_33249_48695.n384 a_33249_48695.t226 1.4705
R51830 a_33249_48695.n383 a_33249_48695.t276 1.4705
R51831 a_33249_48695.n383 a_33249_48695.t218 1.4705
R51832 a_33249_48695.n382 a_33249_48695.t266 1.4705
R51833 a_33249_48695.n382 a_33249_48695.t233 1.4705
R51834 a_33249_48695.n380 a_33249_48695.t215 1.4705
R51835 a_33249_48695.n380 a_33249_48695.t159 1.4705
R51836 a_33249_48695.n376 a_33249_48695.t169 1.4705
R51837 a_33249_48695.n376 a_33249_48695.t286 1.4705
R51838 a_33249_48695.n372 a_33249_48695.t162 1.4705
R51839 a_33249_48695.n372 a_33249_48695.t277 1.4705
R51840 a_33249_48695.n368 a_33249_48695.t329 1.4705
R51841 a_33249_48695.n368 a_33249_48695.t291 1.4705
R51842 a_33249_48695.n67 a_33249_48695.t275 1.4705
R51843 a_33249_48695.n67 a_33249_48695.t217 1.4705
R51844 a_33249_48695.n358 a_33249_48695.t305 1.4705
R51845 a_33249_48695.n358 a_33249_48695.t230 1.4705
R51846 a_33249_48695.n359 a_33249_48695.t223 1.4705
R51847 a_33249_48695.n359 a_33249_48695.t327 1.4705
R51848 a_33249_48695.n354 a_33249_48695.t288 1.4705
R51849 a_33249_48695.n354 a_33249_48695.t190 1.4705
R51850 a_33249_48695.n355 a_33249_48695.t208 1.4705
R51851 a_33249_48695.n355 a_33249_48695.t285 1.4705
R51852 a_33249_48695.n75 a_33249_48695.t239 1.4705
R51853 a_33249_48695.n75 a_33249_48695.t177 1.4705
R51854 a_33249_48695.n74 a_33249_48695.t224 1.4705
R51855 a_33249_48695.n74 a_33249_48695.t167 1.4705
R51856 a_33249_48695.n73 a_33249_48695.t220 1.4705
R51857 a_33249_48695.n73 a_33249_48695.t179 1.4705
R51858 a_33249_48695.n72 a_33249_48695.t166 1.4705
R51859 a_33249_48695.n72 a_33249_48695.t281 1.4705
R51860 a_33249_48695.n182 a_33249_48695.t27 1.4705
R51861 a_33249_48695.n182 a_33249_48695.t62 1.4705
R51862 a_33249_48695.n184 a_33249_48695.t35 1.4705
R51863 a_33249_48695.n184 a_33249_48695.t82 1.4705
R51864 a_33249_48695.n229 a_33249_48695.t31 1.4705
R51865 a_33249_48695.n229 a_33249_48695.t49 1.4705
R51866 a_33249_48695.n230 a_33249_48695.t26 1.4705
R51867 a_33249_48695.n230 a_33249_48695.t47 1.4705
R51868 a_33249_48695.n232 a_33249_48695.t30 1.4705
R51869 a_33249_48695.n232 a_33249_48695.t88 1.4705
R51870 a_33249_48695.n233 a_33249_48695.t25 1.4705
R51871 a_33249_48695.n233 a_33249_48695.t84 1.4705
R51872 a_33249_48695.n236 a_33249_48695.t40 1.4705
R51873 a_33249_48695.n236 a_33249_48695.t65 1.4705
R51874 a_33249_48695.n237 a_33249_48695.t29 1.4705
R51875 a_33249_48695.n237 a_33249_48695.t56 1.4705
R51876 a_33249_48695.n240 a_33249_48695.t69 1.4705
R51877 a_33249_48695.n240 a_33249_48695.t94 1.4705
R51878 a_33249_48695.n241 a_33249_48695.t60 1.4705
R51879 a_33249_48695.n241 a_33249_48695.t87 1.4705
R51880 a_33249_48695.n245 a_33249_48695.t28 1.4705
R51881 a_33249_48695.n245 a_33249_48695.t55 1.4705
R51882 a_33249_48695.n246 a_33249_48695.t23 1.4705
R51883 a_33249_48695.n246 a_33249_48695.t50 1.4705
R51884 a_33249_48695.n249 a_33249_48695.t58 1.4705
R51885 a_33249_48695.n249 a_33249_48695.t98 1.4705
R51886 a_33249_48695.n250 a_33249_48695.t54 1.4705
R51887 a_33249_48695.n250 a_33249_48695.t89 1.4705
R51888 a_33249_48695.n253 a_33249_48695.t67 1.4705
R51889 a_33249_48695.n253 a_33249_48695.t90 1.4705
R51890 a_33249_48695.n254 a_33249_48695.t57 1.4705
R51891 a_33249_48695.n254 a_33249_48695.t86 1.4705
R51892 a_33249_48695.n257 a_33249_48695.t19 1.4705
R51893 a_33249_48695.n257 a_33249_48695.t41 1.4705
R51894 a_33249_48695.n258 a_33249_48695.t102 1.4705
R51895 a_33249_48695.n258 a_33249_48695.t32 1.4705
R51896 a_33249_48695.n202 a_33249_48695.t39 1.4705
R51897 a_33249_48695.n202 a_33249_48695.t53 1.4705
R51898 a_33249_48695.n203 a_33249_48695.t37 1.4705
R51899 a_33249_48695.n203 a_33249_48695.t51 1.4705
R51900 a_33249_48695.n205 a_33249_48695.t38 1.4705
R51901 a_33249_48695.n205 a_33249_48695.t93 1.4705
R51902 a_33249_48695.n206 a_33249_48695.t36 1.4705
R51903 a_33249_48695.n206 a_33249_48695.t92 1.4705
R51904 a_33249_48695.n209 a_33249_48695.t44 1.4705
R51905 a_33249_48695.n209 a_33249_48695.t73 1.4705
R51906 a_33249_48695.n210 a_33249_48695.t42 1.4705
R51907 a_33249_48695.n210 a_33249_48695.t70 1.4705
R51908 a_33249_48695.n213 a_33249_48695.t77 1.4705
R51909 a_33249_48695.n213 a_33249_48695.t100 1.4705
R51910 a_33249_48695.n214 a_33249_48695.t76 1.4705
R51911 a_33249_48695.n214 a_33249_48695.t99 1.4705
R51912 a_33249_48695.n198 a_33249_48695.t34 1.4705
R51913 a_33249_48695.n198 a_33249_48695.t61 1.4705
R51914 a_33249_48695.n199 a_33249_48695.t33 1.4705
R51915 a_33249_48695.n199 a_33249_48695.t59 1.4705
R51916 a_33249_48695.n194 a_33249_48695.t66 1.4705
R51917 a_33249_48695.n194 a_33249_48695.t104 1.4705
R51918 a_33249_48695.n195 a_33249_48695.t64 1.4705
R51919 a_33249_48695.n195 a_33249_48695.t103 1.4705
R51920 a_33249_48695.n190 a_33249_48695.t74 1.4705
R51921 a_33249_48695.n190 a_33249_48695.t97 1.4705
R51922 a_33249_48695.n191 a_33249_48695.t72 1.4705
R51923 a_33249_48695.n191 a_33249_48695.t96 1.4705
R51924 a_33249_48695.n186 a_33249_48695.t22 1.4705
R51925 a_33249_48695.n186 a_33249_48695.t45 1.4705
R51926 a_33249_48695.n187 a_33249_48695.t21 1.4705
R51927 a_33249_48695.n187 a_33249_48695.t43 1.4705
R51928 a_33249_48695.n266 a_33249_48695.t68 1.4705
R51929 a_33249_48695.n266 a_33249_48695.t95 1.4705
R51930 a_33249_48695.n263 a_33249_48695.t78 1.4705
R51931 a_33249_48695.n263 a_33249_48695.t105 1.4705
R51932 a_33249_48695.n181 a_33249_48695.t18 1.4705
R51933 a_33249_48695.n181 a_33249_48695.t52 1.4705
R51934 a_33249_48695.n180 a_33249_48695.t24 1.4705
R51935 a_33249_48695.n180 a_33249_48695.t79 1.4705
R51936 a_33249_48695.n222 a_33249_48695.t75 1.4705
R51937 a_33249_48695.n222 a_33249_48695.t101 1.4705
R51938 a_33249_48695.n219 a_33249_48695.t81 1.4705
R51939 a_33249_48695.n219 a_33249_48695.t20 1.4705
R51940 a_33249_48695.n88 a_33249_48695.t265 1.4705
R51941 a_33249_48695.n88 a_33249_48695.t209 1.4705
R51942 a_33249_48695.n87 a_33249_48695.t253 1.4705
R51943 a_33249_48695.n87 a_33249_48695.t193 1.4705
R51944 a_33249_48695.n107 a_33249_48695.t248 1.4705
R51945 a_33249_48695.n107 a_33249_48695.t172 1.4705
R51946 a_33249_48695.n105 a_33249_48695.t231 1.4705
R51947 a_33249_48695.n105 a_33249_48695.t310 1.4705
R51948 a_33249_48695.n97 a_33249_48695.t257 1.4705
R51949 a_33249_48695.n97 a_33249_48695.t195 1.4705
R51950 a_33249_48695.n98 a_33249_48695.t301 1.4705
R51951 a_33249_48695.n98 a_33249_48695.t243 1.4705
R51952 a_33249_48695.n112 a_33249_48695.t250 1.4705
R51953 a_33249_48695.n112 a_33249_48695.t189 1.4705
R51954 a_33249_48695.n113 a_33249_48695.t292 1.4705
R51955 a_33249_48695.n113 a_33249_48695.t236 1.4705
R51956 a_33249_48695.n120 a_33249_48695.t241 1.4705
R51957 a_33249_48695.n120 a_33249_48695.t201 1.4705
R51958 a_33249_48695.n121 a_33249_48695.t283 1.4705
R51959 a_33249_48695.n121 a_33249_48695.t249 1.4705
R51960 a_33249_48695.n92 a_33249_48695.t186 1.4705
R51961 a_33249_48695.n92 a_33249_48695.t307 1.4705
R51962 a_33249_48695.n93 a_33249_48695.t234 1.4705
R51963 a_33249_48695.n93 a_33249_48695.t174 1.4705
R51964 a_33249_48695.n131 a_33249_48695.t319 1.4705
R51965 a_33249_48695.n131 a_33249_48695.t259 1.4705
R51966 a_33249_48695.n130 a_33249_48695.t303 1.4705
R51967 a_33249_48695.n130 a_33249_48695.t245 1.4705
R51968 a_33249_48695.n138 a_33249_48695.t320 1.4705
R51969 a_33249_48695.n138 a_33249_48695.t247 1.4705
R51970 a_33249_48695.n136 a_33249_48695.t304 1.4705
R51971 a_33249_48695.n136 a_33249_48695.t207 1.4705
R51972 a_33249_48695.n165 a_33249_48695.t330 1.4705
R51973 a_33249_48695.n165 a_33249_48695.t269 1.4705
R51974 a_33249_48695.n166 a_33249_48695.t252 1.4705
R51975 a_33249_48695.n166 a_33249_48695.t191 1.4705
R51976 a_33249_48695.n160 a_33249_48695.t323 1.4705
R51977 a_33249_48695.n160 a_33249_48695.t261 1.4705
R51978 a_33249_48695.n161 a_33249_48695.t240 1.4705
R51979 a_33249_48695.n161 a_33249_48695.t181 1.4705
R51980 a_33249_48695.n152 a_33249_48695.t314 1.4705
R51981 a_33249_48695.n152 a_33249_48695.t274 1.4705
R51982 a_33249_48695.n153 a_33249_48695.t238 1.4705
R51983 a_33249_48695.n153 a_33249_48695.t194 1.4705
R51984 a_33249_48695.n143 a_33249_48695.t260 1.4705
R51985 a_33249_48695.n143 a_33249_48695.t200 1.4705
R51986 a_33249_48695.n144 a_33249_48695.t180 1.4705
R51987 a_33249_48695.n144 a_33249_48695.t298 1.4705
R51988 a_33249_48695.n297 a_33249_48695.t134 1.4705
R51989 a_33249_48695.n297 a_33249_48695.t336 1.4705
R51990 a_33249_48695.n298 a_33249_48695.t133 1.4705
R51991 a_33249_48695.n298 a_33249_48695.t335 1.4705
R51992 a_33249_48695.n281 a_33249_48695.t140 1.4705
R51993 a_33249_48695.n281 a_33249_48695.t0 1.4705
R51994 a_33249_48695.n282 a_33249_48695.t139 1.4705
R51995 a_33249_48695.n282 a_33249_48695.t334 1.4705
R51996 a_33249_48695.n345 a_33249_48695.t111 1.4705
R51997 a_33249_48695.n345 a_33249_48695.t16 1.4705
R51998 a_33249_48695.n343 a_33249_48695.t110 1.4705
R51999 a_33249_48695.n343 a_33249_48695.t137 1.4705
R52000 a_33249_48695.n341 a_33249_48695.t121 1.4705
R52001 a_33249_48695.n341 a_33249_48695.t351 1.4705
R52002 a_33249_48695.n339 a_33249_48695.t4 1.4705
R52003 a_33249_48695.n339 a_33249_48695.t142 1.4705
R52004 a_33249_48695.n83 a_33249_48695.t115 1.4705
R52005 a_33249_48695.n83 a_33249_48695.t344 1.4705
R52006 a_33249_48695.n81 a_33249_48695.t347 1.4705
R52007 a_33249_48695.n81 a_33249_48695.t144 1.4705
R52008 a_33249_48695.n79 a_33249_48695.t3 1.4705
R52009 a_33249_48695.n79 a_33249_48695.t138 1.4705
R52010 a_33249_48695.n78 a_33249_48695.t151 1.4705
R52011 a_33249_48695.n78 a_33249_48695.t112 1.4705
R52012 a_33249_48695.n280 a_33249_48695.t119 1.4705
R52013 a_33249_48695.n280 a_33249_48695.t346 1.4705
R52014 a_33249_48695.n279 a_33249_48695.t118 1.4705
R52015 a_33249_48695.n279 a_33249_48695.t146 1.4705
R52016 a_33249_48695.n278 a_33249_48695.t106 1.4705
R52017 a_33249_48695.n278 a_33249_48695.t12 1.4705
R52018 a_33249_48695.n277 a_33249_48695.t124 1.4705
R52019 a_33249_48695.n277 a_33249_48695.t149 1.4705
R52020 a_33249_48695.n276 a_33249_48695.t113 1.4705
R52021 a_33249_48695.n276 a_33249_48695.t5 1.4705
R52022 a_33249_48695.n275 a_33249_48695.t9 1.4705
R52023 a_33249_48695.n275 a_33249_48695.t152 1.4705
R52024 a_33249_48695.n274 a_33249_48695.t13 1.4705
R52025 a_33249_48695.n274 a_33249_48695.t148 1.4705
R52026 a_33249_48695.n273 a_33249_48695.t337 1.4705
R52027 a_33249_48695.n273 a_33249_48695.t107 1.4705
R52028 a_33249_48695.n318 a_33249_48695.t120 1.4705
R52029 a_33249_48695.n318 a_33249_48695.t342 1.4705
R52030 a_33249_48695.n316 a_33249_48695.t1 1.4705
R52031 a_33249_48695.n316 a_33249_48695.t141 1.4705
R52032 a_33249_48695.n314 a_33249_48695.t114 1.4705
R52033 a_33249_48695.n314 a_33249_48695.t7 1.4705
R52034 a_33249_48695.n312 a_33249_48695.t10 1.4705
R52035 a_33249_48695.n312 a_33249_48695.t145 1.4705
R52036 a_33249_48695.n309 a_33249_48695.t333 1.4705
R52037 a_33249_48695.n309 a_33249_48695.t348 1.4705
R52038 a_33249_48695.n307 a_33249_48695.t2 1.4705
R52039 a_33249_48695.n307 a_33249_48695.t147 1.4705
R52040 a_33249_48695.n305 a_33249_48695.t8 1.4705
R52041 a_33249_48695.n305 a_33249_48695.t143 1.4705
R52042 a_33249_48695.n304 a_33249_48695.t154 1.4705
R52043 a_33249_48695.n304 a_33249_48695.t117 1.4705
R52044 a_33249_48695.n293 a_33249_48695.t15 1.4705
R52045 a_33249_48695.n293 a_33249_48695.t6 1.4705
R52046 a_33249_48695.n292 a_33249_48695.t109 1.4705
R52047 a_33249_48695.n292 a_33249_48695.t153 1.4705
R52048 a_33249_48695.n291 a_33249_48695.t341 1.4705
R52049 a_33249_48695.n291 a_33249_48695.t129 1.4705
R52050 a_33249_48695.n290 a_33249_48695.t135 1.4705
R52051 a_33249_48695.n290 a_33249_48695.t340 1.4705
R52052 a_33249_48695.n289 a_33249_48695.t108 1.4705
R52053 a_33249_48695.n289 a_33249_48695.t123 1.4705
R52054 a_33249_48695.n288 a_33249_48695.t126 1.4705
R52055 a_33249_48695.n288 a_33249_48695.t338 1.4705
R52056 a_33249_48695.n287 a_33249_48695.t132 1.4705
R52057 a_33249_48695.n287 a_33249_48695.t156 1.4705
R52058 a_33249_48695.n286 a_33249_48695.t122 1.4705
R52059 a_33249_48695.n286 a_33249_48695.t343 1.4705
R52060 a_33249_48695.n331 a_33249_48695.t127 1.4705
R52061 a_33249_48695.n331 a_33249_48695.t155 1.4705
R52062 a_33249_48695.n332 a_33249_48695.t14 1.4705
R52063 a_33249_48695.n332 a_33249_48695.t150 1.4705
R52064 a_33249_48695.n324 a_33249_48695.t136 1.4705
R52065 a_33249_48695.n324 a_33249_48695.t116 1.4705
R52066 a_33249_48695.n325 a_33249_48695.t131 1.4705
R52067 a_33249_48695.n325 a_33249_48695.t339 1.4705
R52068 a_33249_48695.n391 a_33249_48695.n390 1.46537
R52069 a_33249_48695.n393 a_33249_48695.n392 1.46537
R52070 a_33249_48695.n56 a_33249_48695.n55 1.46537
R52071 a_33249_48695.n361 a_33249_48695.n360 1.46537
R52072 a_33249_48695.n363 a_33249_48695.n362 1.46537
R52073 a_33249_48695.n357 a_33249_48695.n356 1.46537
R52074 a_33249_48695.n100 a_33249_48695.n99 1.46537
R52075 a_33249_48695.n102 a_33249_48695.n101 1.46537
R52076 a_33249_48695.n115 a_33249_48695.n114 1.46537
R52077 a_33249_48695.n117 a_33249_48695.n116 1.46537
R52078 a_33249_48695.n119 a_33249_48695.n118 1.46537
R52079 a_33249_48695.n123 a_33249_48695.n122 1.46537
R52080 a_33249_48695.n125 a_33249_48695.n124 1.46537
R52081 a_33249_48695.n95 a_33249_48695.n94 1.46537
R52082 a_33249_48695.n168 a_33249_48695.n167 1.46537
R52083 a_33249_48695.n170 a_33249_48695.n169 1.46537
R52084 a_33249_48695.n163 a_33249_48695.n162 1.46537
R52085 a_33249_48695.n159 a_33249_48695.n158 1.46537
R52086 a_33249_48695.n157 a_33249_48695.n156 1.46537
R52087 a_33249_48695.n155 a_33249_48695.n154 1.46537
R52088 a_33249_48695.n151 a_33249_48695.n150 1.46537
R52089 a_33249_48695.n146 a_33249_48695.n145 1.46537
R52090 a_33249_48695.n302 a_33249_48695.n301 1.46537
R52091 a_33249_48695.n300 a_33249_48695.n299 1.46537
R52092 a_33249_48695.n285 a_33249_48695.n284 1.46537
R52093 a_33249_48695.n330 a_33249_48695.n329 1.46537
R52094 a_33249_48695.n334 a_33249_48695.n333 1.46537
R52095 a_33249_48695.n328 a_33249_48695.n327 1.46537
R52096 a_33249_48695.n235 a_33249_48695.n234 1.46537
R52097 a_33249_48695.n239 a_33249_48695.n238 1.46537
R52098 a_33249_48695.n243 a_33249_48695.n242 1.46537
R52099 a_33249_48695.n248 a_33249_48695.n247 1.46537
R52100 a_33249_48695.n252 a_33249_48695.n251 1.46537
R52101 a_33249_48695.n256 a_33249_48695.n255 1.46537
R52102 a_33249_48695.n260 a_33249_48695.n259 1.46537
R52103 a_33249_48695.n208 a_33249_48695.n207 1.46537
R52104 a_33249_48695.n212 a_33249_48695.n211 1.46537
R52105 a_33249_48695.n216 a_33249_48695.n215 1.46537
R52106 a_33249_48695.n201 a_33249_48695.n200 1.46537
R52107 a_33249_48695.n197 a_33249_48695.n196 1.46537
R52108 a_33249_48695.n193 a_33249_48695.n192 1.46537
R52109 a_33249_48695.n189 a_33249_48695.n188 1.46537
R52110 a_33249_48695.n104 a_33249_48695.n103 1.46535
R52111 a_33249_48695.n127 a_33249_48695.n126 1.46535
R52112 a_33249_48695.n172 a_33249_48695.n171 1.46535
R52113 a_33249_48695.n149 a_33249_48695.n148 1.46535
R52114 a_33249_48695.n337 a_33249_48695.n271 1.34705
R52115 a_33249_48695.n270 a_33249_48695.n269 1.2981
R52116 a_33249_48695.n175 a_33249_48695.n76 1.27763
R52117 a_33249_48695.n393 a_33249_48695.n391 1.27228
R52118 a_33249_48695.n370 a_33249_48695.n369 1.27228
R52119 a_33249_48695.n373 a_33249_48695.n371 1.27228
R52120 a_33249_48695.n363 a_33249_48695.n361 1.27228
R52121 a_33249_48695.n106 a_33249_48695.n90 1.27228
R52122 a_33249_48695.n125 a_33249_48695.n123 1.27228
R52123 a_33249_48695.n123 a_33249_48695.n119 1.27228
R52124 a_33249_48695.n117 a_33249_48695.n115 1.27228
R52125 a_33249_48695.n102 a_33249_48695.n100 1.27228
R52126 a_33249_48695.n137 a_33249_48695.n135 1.27228
R52127 a_33249_48695.n155 a_33249_48695.n151 1.27228
R52128 a_33249_48695.n157 a_33249_48695.n155 1.27228
R52129 a_33249_48695.n163 a_33249_48695.n159 1.27228
R52130 a_33249_48695.n170 a_33249_48695.n168 1.27228
R52131 a_33249_48695.n57 a_33249_48695.n50 1.27228
R52132 a_33249_48695.n60 a_33249_48695.n58 1.27228
R52133 a_33249_48695.n260 a_33249_48695.n256 1.27228
R52134 a_33249_48695.n252 a_33249_48695.n248 1.27228
R52135 a_33249_48695.n243 a_33249_48695.n239 1.27228
R52136 a_33249_48695.n193 a_33249_48695.n189 1.27228
R52137 a_33249_48695.n201 a_33249_48695.n197 1.27228
R52138 a_33249_48695.n216 a_33249_48695.n212 1.27228
R52139 a_33249_48695.n265 a_33249_48695.n264 1.27228
R52140 a_33249_48695.n221 a_33249_48695.n220 1.27228
R52141 a_33249_48695.n84 a_33249_48695.n82 1.27228
R52142 a_33249_48695.n342 a_33249_48695.n340 1.27228
R52143 a_33249_48695.n346 a_33249_48695.n344 1.27228
R52144 a_33249_48695.n310 a_33249_48695.n308 1.27228
R52145 a_33249_48695.n315 a_33249_48695.n313 1.27228
R52146 a_33249_48695.n319 a_33249_48695.n317 1.27228
R52147 a_33249_48695.n334 a_33249_48695.n330 1.27228
R52148 a_33249_48695.n302 a_33249_48695.n300 1.27228
R52149 a_33249_48695.n69 a_33249_48695.n68 1.26756
R52150 a_33249_48695.n374 a_33249_48695.n373 1.26756
R52151 a_33249_48695.n48 a_33249_48695.n47 1.26756
R52152 a_33249_48695.n61 a_33249_48695.n60 1.26756
R52153 a_33249_48695.n349 a_33249_48695.n348 1.23567
R52154 a_33249_48695.n352 a_33249_48695.n71 1.23455
R52155 a_33249_48695.n178 a_33249_48695.n177 1.18682
R52156 a_33249_48695.n109 a_33249_48695.n108 1.01873
R52157 a_33249_48695.n140 a_33249_48695.n139 1.01873
R52158 a_33249_48695.n323 a_33249_48695.n272 0.822966
R52159 a_33249_48695.n321 a_33249_48695.n320 0.822966
R52160 a_33249_48695.n367 a_33249_48695.n70 0.796291
R52161 a_33249_48695.n378 a_33249_48695.n375 0.796291
R52162 a_33249_48695.n65 a_33249_48695.n62 0.796291
R52163 a_33249_48695.n397 a_33249_48695.n396 0.795934
R52164 a_33249_48695.n395 a_33249_48695.n51 0.780703
R52165 a_33249_48695.n365 a_33249_48695.n352 0.780703
R52166 a_33249_48695.n387 a_33249_48695.n386 0.780703
R52167 a_33249_48695.n349 a_33249_48695.n66 0.780703
R52168 a_33249_48695.n133 a_33249_48695.n129 0.778574
R52169 a_33249_48695.n177 a_33249_48695.n86 0.778574
R52170 a_33249_48695.n110 a_33249_48695.n89 0.778574
R52171 a_33249_48695.n175 a_33249_48695.n174 0.778574
R52172 a_33249_48695.n134 a_33249_48695.n86 0.738439
R52173 a_33249_48695.n174 a_33249_48695.n141 0.738439
R52174 a_33249_48695.n262 a_33249_48695.n261 0.737223
R52175 a_33249_48695.n185 a_33249_48695.n179 0.737223
R52176 a_33249_48695.n269 a_33249_48695.n85 0.737223
R52177 a_33249_48695.n225 a_33249_48695.n218 0.737223
R52178 a_33249_48695.n228 a_33249_48695.n179 0.725061
R52179 a_33249_48695.n226 a_33249_48695.n225 0.725061
R52180 a_33249_48695.n128 a_33249_48695.n127 0.699581
R52181 a_33249_48695.n111 a_33249_48695.n104 0.699581
R52182 a_33249_48695.n149 a_33249_48695.n147 0.699581
R52183 a_33249_48695.n173 a_33249_48695.n172 0.699581
R52184 a_33249_48695.n337 a_33249_48695.n336 0.639318
R52185 a_33249_48695.n295 a_33249_48695.n272 0.639318
R52186 a_33249_48695.n347 a_33249_48695.n77 0.639318
R52187 a_33249_48695.n320 a_33249_48695.n303 0.639318
R52188 a_33249_48695.n366 a_33249_48695.n365 0.638405
R52189 a_33249_48695.n379 a_33249_48695.n66 0.638405
R52190 a_33249_48695.n366 a_33249_48695.n51 0.628372
R52191 a_33249_48695.n386 a_33249_48695.n379 0.628372
R52192 a_33249_48695.n271 a_33249_48695.n71 0.606869
R52193 a_33249_48695.n270 a_33249_48695.n76 0.60536
R52194 a_33249_48695.n261 a_33249_48695.n228 0.585196
R52195 a_33249_48695.n226 a_33249_48695.n85 0.585196
R52196 a_33249_48695.n336 a_33249_48695.n323 0.585196
R52197 a_33249_48695.n321 a_33249_48695.n77 0.585196
R52198 a_33249_48695.n128 a_33249_48695.n95 0.557791
R52199 a_33249_48695.n115 a_33249_48695.n111 0.557791
R52200 a_33249_48695.n147 a_33249_48695.n146 0.557791
R52201 a_33249_48695.n173 a_33249_48695.n163 0.557791
R52202 a_33249_48695.n134 a_33249_48695.n133 0.530466
R52203 a_33249_48695.n141 a_33249_48695.n89 0.530466
R52204 a_33249_48695.n369 a_33249_48695.n367 0.476484
R52205 a_33249_48695.n378 a_33249_48695.n377 0.476484
R52206 a_33249_48695.n396 a_33249_48695.n50 0.476484
R52207 a_33249_48695.n65 a_33249_48695.n64 0.476484
R52208 a_33249_48695.n6 a_33249_48695.n381 0.478684
R52209 a_33249_48695.n385 a_33249_48695.n0 0.478684
R52210 a_33249_48695.n351 a_33249_48695.n16 0.478684
R52211 a_33249_48695.n350 a_33249_48695.n10 0.478684
R52212 a_33249_48695.n338 a_33249_48695.n84 0.236091
R52213 a_33249_48695.n311 a_33249_48695.n310 0.236091
R52214 a_33249_48695.n244 a_33249_48695.n243 0.150184
R52215 a_33249_48695.n217 a_33249_48695.n216 0.150184
R52216 a_33249_48695.n8 a_33249_48695.n9 1.27228
R52217 a_33249_48695.n7 a_33249_48695.n8 2.51878
R52218 a_33249_48695.n381 a_33249_48695.n7 0.794091
R52219 a_33249_48695.n5 a_33249_48695.n6 1.27228
R52220 a_33249_48695.n4 a_33249_48695.n5 2.60203
R52221 a_33249_48695.n3 a_33249_48695.n4 1.27228
R52222 a_33249_48695.n2 a_33249_48695.n3 1.27228
R52223 a_33249_48695.n1 a_33249_48695.n2 2.51878
R52224 a_33249_48695.n385 a_33249_48695.n1 0.794091
R52225 a_33249_48695.t188 a_33249_48695.n0 6.77266
R52226 a_33249_48695.n18 a_33249_48695.n19 1.27228
R52227 a_33249_48695.n17 a_33249_48695.n18 2.51878
R52228 a_33249_48695.n351 a_33249_48695.n17 0.794091
R52229 a_33249_48695.n15 a_33249_48695.n16 1.27228
R52230 a_33249_48695.n14 a_33249_48695.n15 2.60203
R52231 a_33249_48695.n13 a_33249_48695.n14 1.27228
R52232 a_33249_48695.n12 a_33249_48695.n13 1.27228
R52233 a_33249_48695.n11 a_33249_48695.n12 2.51878
R52234 a_33249_48695.n350 a_33249_48695.n11 0.794091
R52235 a_33249_48695.t313 a_33249_48695.n10 6.77266
R52236 a_33249_48695.n24 a_33249_48695.n25 1.26457
R52237 a_33249_48695.n227 a_33249_48695.n24 6.59229
R52238 a_33249_48695.n181 a_33249_48695.n23 5.10549
R52239 a_33249_48695.n21 a_33249_48695.n22 1.26457
R52240 a_33249_48695.n183 a_33249_48695.n21 6.59229
R52241 a_33249_48695.n182 a_33249_48695.n20 5.10549
R52242 a_33249_48695.n30 a_33249_48695.n31 1.27228
R52243 a_33249_48695.n132 a_33249_48695.n30 7.30549
R52244 a_33249_48695.t183 a_33249_48695.n29 6.96214
R52245 a_33249_48695.n27 a_33249_48695.n28 1.27228
R52246 a_33249_48695.n176 a_33249_48695.n27 7.30549
R52247 a_33249_48695.t311 a_33249_48695.n26 6.96214
R52248 a_33249_48695.n37 a_33249_48695.n38 3.79678
R52249 a_33249_48695.n36 a_33249_48695.n37 1.27228
R52250 a_33249_48695.n322 a_33249_48695.n36 0.238291
R52251 a_33249_48695.n34 a_33249_48695.n35 1.27228
R52252 a_33249_48695.n33 a_33249_48695.n34 3.79678
R52253 a_33249_48695.n32 a_33249_48695.n33 1.27228
R52254 a_33249_48695.n321 a_33249_48695.n32 1.73829
R52255 a_33249_48695.n44 a_33249_48695.n45 3.79678
R52256 a_33249_48695.n43 a_33249_48695.n44 1.27228
R52257 a_33249_48695.n294 a_33249_48695.n43 0.238291
R52258 a_33249_48695.n41 a_33249_48695.n42 1.27228
R52259 a_33249_48695.n40 a_33249_48695.n41 3.79678
R52260 a_33249_48695.n39 a_33249_48695.n40 1.27228
R52261 a_33249_48695.n39 a_33249_48695.n303 2.32299
R52262 OUT.n14 OUT.n13 12.1937
R52263 OUT.n13 OUT.t0 11.5094
R52264 OUT.n13 OUT.t1 9.24966
R52265 OUT.n27 OUT.n20 7.94229
R52266 OUT.n80 OUT.n78 7.94229
R52267 OUT.n117 OUT.n14 7.76579
R52268 OUT.n75 OUT.n68 7.169
R52269 OUT.n142 OUT.n141 7.169
R52270 OUT.n121 OUT.t4 6.96668
R52271 OUT.n8 OUT.t81 6.82564
R52272 OUT.n72 OUT.t92 6.82564
R52273 OUT.n14 OUT.n12 6.28314
R52274 OUT.n137 OUT.t18 5.85326
R52275 OUT.n137 OUT.n136 5.84661
R52276 OUT.n19 OUT.t93 5.69423
R52277 OUT.n28 OUT.t68 5.69423
R52278 OUT.n17 OUT.t85 5.69423
R52279 OUT.n81 OUT.t66 5.69423
R52280 OUT.n19 OUT.n18 5.49558
R52281 OUT.n17 OUT.n16 5.49558
R52282 OUT.n10 OUT.n9 4.61332
R52283 OUT.n144 OUT.n143 4.61332
R52284 OUT.n74 OUT.n73 4.61332
R52285 OUT.n67 OUT.n65 4.61332
R52286 OUT.n63 OUT.n60 4.61332
R52287 OUT.n123 OUT.n122 4.61332
R52288 OUT.n2 OUT.n1 4.61332
R52289 OUT.n9 OUT.n8 4.60571
R52290 OUT.n143 OUT.n142 4.60571
R52291 OUT.n73 OUT.n72 4.60571
R52292 OUT.n68 OUT.n67 4.60571
R52293 OUT.n64 OUT.n63 4.60571
R52294 OUT.n122 OUT.n121 4.60571
R52295 OUT.n145 OUT.n1 4.60571
R52296 OUT.n62 OUT.n59 4.5005
R52297 OUT.n66 OUT.n58 4.5005
R52298 OUT.n71 OUT.n69 4.5005
R52299 OUT.n120 OUT.n118 4.5005
R52300 OUT.n4 OUT.n3 4.5005
R52301 OUT.n7 OUT.n5 4.5005
R52302 OUT.n147 OUT.n146 4.5005
R52303 OUT.n4 OUT.t78 4.22462
R52304 OUT.n66 OUT.t82 4.22462
R52305 OUT.n27 OUT.n26 4.22423
R52306 OUT.n80 OUT.n79 4.22423
R52307 OUT.n130 OUT.t17 4.21195
R52308 OUT.n132 OUT.t2 4.21195
R52309 OUT.n47 OUT.t41 4.05054
R52310 OUT.n52 OUT.t39 4.05054
R52311 OUT.n54 OUT.t38 4.05054
R52312 OUT.n41 OUT.t100 4.05054
R52313 OUT.n39 OUT.t34 4.05054
R52314 OUT.n33 OUT.t27 4.05054
R52315 OUT.n31 OUT.t79 4.05054
R52316 OUT.n21 OUT.t107 4.05054
R52317 OUT.n88 OUT.t32 4.05054
R52318 OUT.n93 OUT.t25 4.05054
R52319 OUT.n95 OUT.t21 4.05054
R52320 OUT.n102 OUT.t84 4.05054
R52321 OUT.n104 OUT.t102 4.05054
R52322 OUT.n110 OUT.t97 4.05054
R52323 OUT.n112 OUT.t74 4.05054
R52324 OUT.n83 OUT.t89 4.05054
R52325 OUT.n130 OUT.t9 4.03668
R52326 OUT.n132 OUT.t11 4.03668
R52327 OUT.n47 OUT.t37 3.87765
R52328 OUT.n52 OUT.t33 3.87765
R52329 OUT.n54 OUT.t29 3.87765
R52330 OUT.n41 OUT.t91 3.87765
R52331 OUT.n39 OUT.t22 3.87765
R52332 OUT.n33 OUT.t104 3.87765
R52333 OUT.n31 OUT.t75 3.87765
R52334 OUT.n21 OUT.t95 3.87765
R52335 OUT.n88 OUT.t30 3.87765
R52336 OUT.n93 OUT.t24 3.87765
R52337 OUT.n95 OUT.t20 3.87765
R52338 OUT.n102 OUT.t83 3.87765
R52339 OUT.n104 OUT.t99 3.87765
R52340 OUT.n110 OUT.t96 3.87765
R52341 OUT.n112 OUT.t73 3.87765
R52342 OUT.n83 OUT.t87 3.87765
R52343 OUT.n135 OUT.n123 3.81532
R52344 OUT.n140 OUT.n139 3.544
R52345 OUT.n29 OUT.n28 3.25667
R52346 OUT.n120 OUT.n119 3.12366
R52347 OUT.n60 OUT.n15 3.01925
R52348 OUT.n116 OUT.n2 3.01925
R52349 OUT.n129 OUT.n128 2.95195
R52350 OUT.n126 OUT.n125 2.95195
R52351 OUT.n129 OUT.n127 2.77668
R52352 OUT.n126 OUT.n124 2.77668
R52353 OUT.n7 OUT.n6 2.75462
R52354 OUT.n71 OUT.n70 2.75462
R52355 OUT.n62 OUT.n61 2.75462
R52356 OUT.n25 OUT.n21 2.73714
R52357 OUT.n87 OUT.n83 2.73714
R52358 OUT.n51 OUT.n47 2.73672
R52359 OUT.n92 OUT.n88 2.73672
R52360 OUT.n131 OUT.n129 2.71872
R52361 OUT.n42 OUT.n40 2.60203
R52362 OUT.n105 OUT.n103 2.60203
R52363 OUT.n50 OUT.n49 2.58054
R52364 OUT.n45 OUT.n44 2.58054
R52365 OUT.n37 OUT.n36 2.58054
R52366 OUT.n24 OUT.n23 2.58054
R52367 OUT.n91 OUT.n90 2.58054
R52368 OUT.n100 OUT.n99 2.58054
R52369 OUT.n108 OUT.n107 2.58054
R52370 OUT.n86 OUT.n85 2.58054
R52371 OUT.n133 OUT.n131 2.56118
R52372 OUT.n138 OUT.n137 2.54573
R52373 OUT.n34 OUT.n32 2.53418
R52374 OUT.n55 OUT.n53 2.53418
R52375 OUT.n113 OUT.n111 2.53418
R52376 OUT.n96 OUT.n94 2.53418
R52377 OUT.n82 OUT.n81 2.51873
R52378 OUT.n50 OUT.n48 2.40765
R52379 OUT.n45 OUT.n43 2.40765
R52380 OUT.n37 OUT.n35 2.40765
R52381 OUT.n24 OUT.n22 2.40765
R52382 OUT.n91 OUT.n89 2.40765
R52383 OUT.n100 OUT.n98 2.40765
R52384 OUT.n108 OUT.n106 2.40765
R52385 OUT.n86 OUT.n84 2.40765
R52386 OUT.n139 OUT.n117 2.25854
R52387 OUT.n57 OUT.n20 2.23844
R52388 OUT OUT.n0 2.05949
R52389 OUT.n134 OUT.n126 2.00466
R52390 OUT.n75 OUT.n74 1.51925
R52391 OUT.n141 OUT.n10 1.51925
R52392 OUT.n115 OUT.n114 1.5005
R52393 OUT.n30 OUT.n29 1.5005
R52394 OUT.n135 OUT.n134 1.5005
R52395 OUT.n97 OUT.n11 1.5005
R52396 OUT.n78 OUT.n77 1.5005
R52397 OUT.n76 OUT.n75 1.5005
R52398 OUT.n57 OUT.n56 1.5005
R52399 OUT.n141 OUT.n140 1.5005
R52400 OUT.n0 OUT.t50 1.4705
R52401 OUT.n0 OUT.t45 1.4705
R52402 OUT.n6 OUT.t76 1.4705
R52403 OUT.n6 OUT.t52 1.4705
R52404 OUT.n18 OUT.t69 1.4705
R52405 OUT.n18 OUT.t26 1.4705
R52406 OUT.n26 OUT.t65 1.4705
R52407 OUT.n26 OUT.t98 1.4705
R52408 OUT.n48 OUT.t72 1.4705
R52409 OUT.n48 OUT.t59 1.4705
R52410 OUT.n49 OUT.t77 1.4705
R52411 OUT.n49 OUT.t64 1.4705
R52412 OUT.n43 OUT.t49 1.4705
R52413 OUT.n43 OUT.t23 1.4705
R52414 OUT.n44 OUT.t57 1.4705
R52415 OUT.n44 OUT.t35 1.4705
R52416 OUT.n35 OUT.t58 1.4705
R52417 OUT.n35 OUT.t36 1.4705
R52418 OUT.n36 OUT.t63 1.4705
R52419 OUT.n36 OUT.t40 1.4705
R52420 OUT.n22 OUT.t44 1.4705
R52421 OUT.n22 OUT.t94 1.4705
R52422 OUT.n23 OUT.t48 1.4705
R52423 OUT.n23 OUT.t106 1.4705
R52424 OUT.n70 OUT.t80 1.4705
R52425 OUT.n70 OUT.t62 1.4705
R52426 OUT.n61 OUT.t61 1.4705
R52427 OUT.n61 OUT.t55 1.4705
R52428 OUT.n16 OUT.t67 1.4705
R52429 OUT.n16 OUT.t105 1.4705
R52430 OUT.n79 OUT.t60 1.4705
R52431 OUT.n79 OUT.t90 1.4705
R52432 OUT.n89 OUT.t70 1.4705
R52433 OUT.n89 OUT.t53 1.4705
R52434 OUT.n90 OUT.t71 1.4705
R52435 OUT.n90 OUT.t56 1.4705
R52436 OUT.n98 OUT.t46 1.4705
R52437 OUT.n98 OUT.t101 1.4705
R52438 OUT.n99 OUT.t47 1.4705
R52439 OUT.n99 OUT.t103 1.4705
R52440 OUT.n106 OUT.t51 1.4705
R52441 OUT.n106 OUT.t28 1.4705
R52442 OUT.n107 OUT.t54 1.4705
R52443 OUT.n107 OUT.t31 1.4705
R52444 OUT.n84 OUT.t42 1.4705
R52445 OUT.n84 OUT.t86 1.4705
R52446 OUT.n85 OUT.t43 1.4705
R52447 OUT.n85 OUT.t88 1.4705
R52448 OUT.n51 OUT.n50 1.46537
R52449 OUT.n53 OUT.n52 1.46537
R52450 OUT.n46 OUT.n45 1.46537
R52451 OUT.n42 OUT.n41 1.46537
R52452 OUT.n40 OUT.n39 1.46537
R52453 OUT.n38 OUT.n37 1.46537
R52454 OUT.n34 OUT.n33 1.46537
R52455 OUT.n25 OUT.n24 1.46537
R52456 OUT.n92 OUT.n91 1.46537
R52457 OUT.n94 OUT.n93 1.46537
R52458 OUT.n101 OUT.n100 1.46537
R52459 OUT.n103 OUT.n102 1.46537
R52460 OUT.n105 OUT.n104 1.46537
R52461 OUT.n109 OUT.n108 1.46537
R52462 OUT.n111 OUT.n110 1.46537
R52463 OUT.n87 OUT.n86 1.46537
R52464 OUT.n131 OUT.n130 1.46537
R52465 OUT.n55 OUT.n54 1.46535
R52466 OUT.n32 OUT.n31 1.46535
R52467 OUT.n96 OUT.n95 1.46535
R52468 OUT.n113 OUT.n112 1.46535
R52469 OUT.n133 OUT.n132 1.46535
R52470 OUT.n28 OUT.n27 1.27228
R52471 OUT.n38 OUT.n34 1.27228
R52472 OUT.n40 OUT.n38 1.27228
R52473 OUT.n46 OUT.n42 1.27228
R52474 OUT.n53 OUT.n51 1.27228
R52475 OUT.n81 OUT.n80 1.27228
R52476 OUT.n111 OUT.n109 1.27228
R52477 OUT.n109 OUT.n105 1.27228
R52478 OUT.n103 OUT.n101 1.27228
R52479 OUT.n94 OUT.n92 1.27228
R52480 OUT.n136 OUT.t5 1.2605
R52481 OUT.n136 OUT.t12 1.2605
R52482 OUT.n127 OUT.t7 1.2605
R52483 OUT.n127 OUT.t13 1.2605
R52484 OUT.n128 OUT.t15 1.2605
R52485 OUT.n128 OUT.t3 1.2605
R52486 OUT.n124 OUT.t19 1.2605
R52487 OUT.n124 OUT.t6 1.2605
R52488 OUT.n125 OUT.t8 1.2605
R52489 OUT.n125 OUT.t14 1.2605
R52490 OUT.n119 OUT.t10 1.2605
R52491 OUT.n119 OUT.t16 1.2605
R52492 OUT.n139 OUT.n138 1.25797
R52493 OUT.n117 OUT.n116 1.22361
R52494 OUT.n20 OUT.n19 1.01873
R52495 OUT.n78 OUT.n17 1.01873
R52496 OUT.n65 OUT.n64 0.9995
R52497 OUT.n145 OUT.n144 0.9995
R52498 OUT.n29 OUT.n15 0.778574
R52499 OUT.n116 OUT.n115 0.778574
R52500 OUT.n76 OUT.n57 0.778574
R52501 OUT.n140 OUT.n11 0.778574
R52502 OUT.n115 OUT.n82 0.738439
R52503 OUT.n138 OUT.n135 0.738439
R52504 OUT.n77 OUT.n11 0.738439
R52505 OUT.n32 OUT.n30 0.699581
R52506 OUT.n56 OUT.n55 0.699581
R52507 OUT.n114 OUT.n113 0.699581
R52508 OUT.n97 OUT.n96 0.699581
R52509 OUT.n134 OUT.n133 0.699581
R52510 OUT OUT.n147 0.695632
R52511 OUT.n30 OUT.n25 0.557791
R52512 OUT.n56 OUT.n46 0.557791
R52513 OUT.n114 OUT.n87 0.557791
R52514 OUT.n101 OUT.n97 0.557791
R52515 OUT.n82 OUT.n15 0.530466
R52516 OUT.n77 OUT.n76 0.530466
R52517 OUT.n60 OUT.n59 0.14
R52518 OUT.n64 OUT.n59 0.14
R52519 OUT.n65 OUT.n58 0.14
R52520 OUT.n68 OUT.n58 0.14
R52521 OUT.n74 OUT.n69 0.14
R52522 OUT.n72 OUT.n69 0.14
R52523 OUT.n123 OUT.n118 0.14
R52524 OUT.n121 OUT.n118 0.14
R52525 OUT.n146 OUT.n2 0.14
R52526 OUT.n146 OUT.n145 0.14
R52527 OUT.n144 OUT.n3 0.14
R52528 OUT.n142 OUT.n3 0.14
R52529 OUT.n10 OUT.n5 0.14
R52530 OUT.n8 OUT.n5 0.14
R52531 OUT.n12 OUT.t109 0.134004
R52532 OUT.n12 OUT.t108 0.03175
R52533 OUT.n9 OUT.n7 0.00168421
R52534 OUT.n143 OUT.n4 0.00168421
R52535 OUT.n73 OUT.n71 0.00168421
R52536 OUT.n67 OUT.n66 0.00168421
R52537 OUT.n63 OUT.n62 0.00168421
R52538 OUT.n122 OUT.n120 0.00168421
R52539 OUT.n147 OUT.n1 0.00168421
R52540 a_30324_n30399.t1 a_30324_n30399.t2 24.9025
R52541 a_30324_n30399.t0 a_30324_n30399.t1 19.5272
R52542 a_31284_n30339.t1 a_31284_n30339.t2 26.4056
R52543 a_31284_n30339.t1 a_31284_n30339.t0 20.6404
R52544 a_100992_n29313.t0 a_100992_n29313.t2 23.2303
R52545 a_100992_n29313.t0 a_100992_n29313.t1 21.6695
R52546 a_38097_n5342.t1 a_38097_n5342.t2 123.341
R52547 a_38097_n5342.t1 a_38097_n5342.t0 20.6404
R52548 a_100992_4421.t2 a_100992_4421.t0 21.6693
R52549 a_100992_4421.t1 a_100992_4421.t0 15.3476
R52550 a_71496_10388.n5 a_71496_10388.n1 10.2377
R52551 a_71496_10388.n4 a_71496_10388.t2 10.2108
R52552 a_71496_10388.n4 a_71496_10388.t0 9.99909
R52553 a_71496_10388.n5 a_71496_10388.t5 9.80443
R52554 a_71496_10388.n5 a_71496_10388.t7 9.55135
R52555 a_71496_10388.n0 a_71496_10388.t19 8.17385
R52556 a_71496_10388.n3 a_71496_10388.t12 8.17299
R52557 a_71496_10388.n3 a_71496_10388.t14 8.17134
R52558 a_71496_10388.n0 a_71496_10388.t10 8.16754
R52559 a_71496_10388.n1 a_71496_10388.t11 8.10567
R52560 a_71496_10388.n1 a_71496_10388.t9 8.10567
R52561 a_71496_10388.n3 a_71496_10388.t22 8.10567
R52562 a_71496_10388.n3 a_71496_10388.t23 8.10567
R52563 a_71496_10388.n1 a_71496_10388.t8 8.10567
R52564 a_71496_10388.n1 a_71496_10388.t17 8.10567
R52565 a_71496_10388.n0 a_71496_10388.t13 8.10567
R52566 a_71496_10388.n0 a_71496_10388.t21 8.10567
R52567 a_71496_10388.n6 a_71496_10388.t3 7.74799
R52568 a_71496_10388.n7 a_71496_10388.t6 7.73052
R52569 a_71496_10388.n6 a_71496_10388.t1 7.46478
R52570 a_71496_10388.t4 a_71496_10388.n7 7.1311
R52571 a_71496_10388.n4 a_71496_10388.n6 2.2505
R52572 a_71496_10388.n7 a_71496_10388.n5 2.2505
R52573 a_71496_10388.n1 a_71496_10388.t15 8.35731
R52574 a_71496_10388.n0 a_71496_10388.t20 8.38107
R52575 a_71496_10388.n1 a_71496_10388.t16 8.37583
R52576 a_71496_10388.n1 a_71496_10388.n0 4.35656
R52577 a_71496_10388.n5 a_71496_10388.n4 2.96863
R52578 a_71496_10388.n2 a_71496_10388.n1 1.0882
R52579 a_71496_10388.n2 a_71496_10388.n3 1.08408
R52580 a_71496_10388.n2 a_71496_10388.t18 8.66753
R52581 a_71342_4481.n0 a_71342_4481.t1 10.6581
R52582 a_71342_4481.n0 a_71342_4481.t3 10.2356
R52583 a_71342_4481.t2 a_71342_4481.n0 9.5019
R52584 a_71342_4481.n0 a_71342_4481.t0 9.34796
R52585 a_30152_10448.t3 a_30152_10448.t11 12.7127
R52586 a_30152_10448.t3 a_30152_10448.t6 10.2828
R52587 a_30152_10448.t3 a_30152_10448.t8 10.2828
R52588 a_30152_10448.t3 a_30152_10448.t19 10.2828
R52589 a_30152_10448.t3 a_30152_10448.t14 10.2828
R52590 a_30152_10448.t3 a_30152_10448.t22 10.1333
R52591 a_30152_10448.t3 a_30152_10448.t23 10.1333
R52592 a_30152_10448.t3 a_30152_10448.t10 10.1333
R52593 a_30152_10448.t3 a_30152_10448.t4 10.1333
R52594 a_30152_10448.t3 a_30152_10448.t0 9.72545
R52595 a_30152_10448.t3 a_30152_10448.t21 9.57156
R52596 a_30152_10448.t3 a_30152_10448.t17 9.57156
R52597 a_30152_10448.t3 a_30152_10448.t18 9.57156
R52598 a_30152_10448.t3 a_30152_10448.t13 9.57156
R52599 a_30152_10448.t3 a_30152_10448.t20 9.57156
R52600 a_30152_10448.t3 a_30152_10448.t15 9.57156
R52601 a_30152_10448.t3 a_30152_10448.t16 9.57156
R52602 a_30152_10448.t3 a_30152_10448.t12 9.57156
R52603 a_30152_10448.t0 a_30152_10448.t2 8.02945
R52604 a_30152_10448.t3 a_30152_10448.t1 8.02708
R52605 a_30152_10448.t3 a_30152_10448.t9 7.90829
R52606 a_30152_10448.t3 a_30152_10448.t7 7.90829
R52607 a_30152_10448.t5 a_30152_10448.t3 7.41776
R52608 a_32913_n8930.t0 a_32913_n8930.t1 103.29
R52609 a_32913_n8930.t1 a_32913_n8930.t2 24.9025
R52610 a_31831_n5342.t1 a_31831_n5342.t2 108.376
R52611 a_31831_n5342.t1 a_31831_n5342.t0 20.6404
R52612 a_51711_n5344.t0 a_51711_n5344.t1 13.2434
R52613 a_33379_34917.n1 a_33379_34917.t2 10.937
R52614 a_33379_34917.n1 a_33379_34917.n0 10.9194
R52615 a_33379_34917.n1 a_33379_34917.t1 9.33982
R52616 a_33379_34917.n6 a_33379_34917.n5 1.21431
R52617 a_33379_34917.n9 a_33379_34917.n1 8.36604
R52618 a_33379_34917.n0 a_33379_34917.t82 8.10567
R52619 a_33379_34917.n3 a_33379_34917.t36 8.10567
R52620 a_33379_34917.n3 a_33379_34917.t22 8.10567
R52621 a_33379_34917.n3 a_33379_34917.t78 8.10567
R52622 a_33379_34917.n3 a_33379_34917.t21 8.10567
R52623 a_33379_34917.n0 a_33379_34917.t55 8.10567
R52624 a_33379_34917.n0 a_33379_34917.t27 8.10567
R52625 a_33379_34917.n0 a_33379_34917.t85 8.10567
R52626 a_33379_34917.n0 a_33379_34917.t61 8.10567
R52627 a_33379_34917.n2 a_33379_34917.t44 8.10567
R52628 a_33379_34917.n2 a_33379_34917.t18 8.10567
R52629 a_33379_34917.n2 a_33379_34917.t89 8.10567
R52630 a_33379_34917.n2 a_33379_34917.t49 8.10567
R52631 a_33379_34917.n3 a_33379_34917.t47 8.10567
R52632 a_33379_34917.n3 a_33379_34917.t12 8.10567
R52633 a_33379_34917.n3 a_33379_34917.t71 8.10567
R52634 a_33379_34917.n2 a_33379_34917.t67 8.10567
R52635 a_33379_34917.n2 a_33379_34917.t20 8.10567
R52636 a_33379_34917.n2 a_33379_34917.t77 8.10567
R52637 a_33379_34917.n0 a_33379_34917.t57 8.10567
R52638 a_33379_34917.n0 a_33379_34917.t28 8.10567
R52639 a_33379_34917.n0 a_33379_34917.t6 8.10567
R52640 a_33379_34917.n4 a_33379_34917.t76 8.10567
R52641 a_33379_34917.n0 a_33379_34917.t34 8.10567
R52642 a_33379_34917.n0 a_33379_34917.t16 8.10567
R52643 a_33379_34917.n0 a_33379_34917.t74 8.10567
R52644 a_33379_34917.n0 a_33379_34917.t15 8.10567
R52645 a_33379_34917.n0 a_33379_34917.t50 8.10567
R52646 a_33379_34917.n0 a_33379_34917.t25 8.10567
R52647 a_33379_34917.n0 a_33379_34917.t80 8.10567
R52648 a_33379_34917.n0 a_33379_34917.t54 8.10567
R52649 a_33379_34917.n6 a_33379_34917.t40 8.10567
R52650 a_33379_34917.n6 a_33379_34917.t13 8.10567
R52651 a_33379_34917.n6 a_33379_34917.t84 8.10567
R52652 a_33379_34917.n6 a_33379_34917.t43 8.10567
R52653 a_33379_34917.n0 a_33379_34917.t31 8.10567
R52654 a_33379_34917.n0 a_33379_34917.t81 8.10567
R52655 a_33379_34917.n0 a_33379_34917.t53 8.10567
R52656 a_33379_34917.n4 a_33379_34917.t48 8.10567
R52657 a_33379_34917.n4 a_33379_34917.t91 8.10567
R52658 a_33379_34917.n4 a_33379_34917.t63 8.10567
R52659 a_33379_34917.n4 a_33379_34917.t52 8.10567
R52660 a_33379_34917.n4 a_33379_34917.t26 8.10567
R52661 a_33379_34917.n4 a_33379_34917.t4 8.10567
R52662 a_33379_34917.n0 a_33379_34917.t72 8.10567
R52663 a_33379_34917.n7 a_33379_34917.t32 8.10567
R52664 a_33379_34917.n7 a_33379_34917.t11 8.10567
R52665 a_33379_34917.n7 a_33379_34917.t70 8.10567
R52666 a_33379_34917.n7 a_33379_34917.t10 8.10567
R52667 a_33379_34917.n0 a_33379_34917.t41 8.10567
R52668 a_33379_34917.n0 a_33379_34917.t14 8.10567
R52669 a_33379_34917.n0 a_33379_34917.t73 8.10567
R52670 a_33379_34917.n0 a_33379_34917.t45 8.10567
R52671 a_33379_34917.n0 a_33379_34917.t35 8.10567
R52672 a_33379_34917.n0 a_33379_34917.t8 8.10567
R52673 a_33379_34917.n0 a_33379_34917.t75 8.10567
R52674 a_33379_34917.n0 a_33379_34917.t39 8.10567
R52675 a_33379_34917.n0 a_33379_34917.t37 8.10567
R52676 a_33379_34917.n0 a_33379_34917.t3 8.10567
R52677 a_33379_34917.n0 a_33379_34917.t65 8.10567
R52678 a_33379_34917.n0 a_33379_34917.t64 8.10567
R52679 a_33379_34917.n0 a_33379_34917.t9 8.10567
R52680 a_33379_34917.n0 a_33379_34917.t69 8.10567
R52681 a_33379_34917.n0 a_33379_34917.t42 8.10567
R52682 a_33379_34917.n0 a_33379_34917.t17 8.10567
R52683 a_33379_34917.n0 a_33379_34917.t88 8.10567
R52684 a_33379_34917.n0 a_33379_34917.t83 8.10567
R52685 a_33379_34917.n8 a_33379_34917.t38 8.10567
R52686 a_33379_34917.n8 a_33379_34917.t24 8.10567
R52687 a_33379_34917.n8 a_33379_34917.t79 8.10567
R52688 a_33379_34917.n8 a_33379_34917.t23 8.10567
R52689 a_33379_34917.n0 a_33379_34917.t58 8.10567
R52690 a_33379_34917.n0 a_33379_34917.t29 8.10567
R52691 a_33379_34917.n0 a_33379_34917.t86 8.10567
R52692 a_33379_34917.n0 a_33379_34917.t62 8.10567
R52693 a_33379_34917.n0 a_33379_34917.t46 8.10567
R52694 a_33379_34917.n0 a_33379_34917.t19 8.10567
R52695 a_33379_34917.n0 a_33379_34917.t90 8.10567
R52696 a_33379_34917.n0 a_33379_34917.t51 8.10567
R52697 a_33379_34917.n0 a_33379_34917.t33 8.10567
R52698 a_33379_34917.n0 a_33379_34917.t87 8.10567
R52699 a_33379_34917.n0 a_33379_34917.t60 8.10567
R52700 a_33379_34917.n0 a_33379_34917.t56 8.10567
R52701 a_33379_34917.n0 a_33379_34917.t5 8.10567
R52702 a_33379_34917.n0 a_33379_34917.t66 8.10567
R52703 a_33379_34917.n0 a_33379_34917.t59 8.10567
R52704 a_33379_34917.n0 a_33379_34917.t30 8.10567
R52705 a_33379_34917.n0 a_33379_34917.t7 8.10567
R52706 a_33379_34917.t0 a_33379_34917.n9 6.76216
R52707 a_33379_34917.n9 a_33379_34917.t68 6.15224
R52708 a_33379_34917.n0 a_33379_34917.n2 6.81859
R52709 a_33379_34917.n3 a_33379_34917.n0 6.66138
R52710 a_33379_34917.n5 a_33379_34917.n4 0.358927
R52711 a_33379_34917.n0 a_33379_34917.n5 1.88254
R52712 a_33379_34917.n0 a_33379_34917.n8 5.10926
R52713 a_33379_34917.n7 a_33379_34917.n0 5.07392
R52714 a_45445_n19595.t0 a_45445_n19595.t1 49.4223
R52715 a_45445_n19595.t1 a_45445_n19595.t2 24.9025
R52716 a_71281_n10073.n21 a_71281_n10073.t173 10.5154
R52717 a_71281_n10073.t173 a_71281_n10073.n16 10.5154
R52718 a_71281_n10073.n35 a_71281_n10073.t168 10.5154
R52719 a_71281_n10073.t168 a_71281_n10073.n30 10.5154
R52720 a_71281_n10073.n49 a_71281_n10073.t239 10.5154
R52721 a_71281_n10073.t239 a_71281_n10073.n44 10.5154
R52722 a_71281_n10073.t225 a_71281_n10073.n861 10.5154
R52723 a_71281_n10073.n865 a_71281_n10073.t225 10.5154
R52724 a_71281_n10073.t310 a_71281_n10073.n847 10.5154
R52725 a_71281_n10073.n851 a_71281_n10073.t310 10.5154
R52726 a_71281_n10073.t279 a_71281_n10073.n830 10.5154
R52727 a_71281_n10073.n834 a_71281_n10073.t279 10.5154
R52728 a_71281_n10073.t85 a_71281_n10073.n816 10.5154
R52729 a_71281_n10073.n820 a_71281_n10073.t85 10.5154
R52730 a_71281_n10073.t81 a_71281_n10073.n802 10.5154
R52731 a_71281_n10073.n806 a_71281_n10073.t81 10.5154
R52732 a_71281_n10073.t146 a_71281_n10073.n788 10.5154
R52733 a_71281_n10073.n792 a_71281_n10073.t146 10.5154
R52734 a_71281_n10073.t330 a_71281_n10073.n175 10.5154
R52735 a_71281_n10073.n179 a_71281_n10073.t330 10.5154
R52736 a_71281_n10073.t294 a_71281_n10073.n161 10.5154
R52737 a_71281_n10073.n165 a_71281_n10073.t294 10.5154
R52738 a_71281_n10073.t309 a_71281_n10073.n147 10.5154
R52739 a_71281_n10073.n151 a_71281_n10073.t309 10.5154
R52740 a_71281_n10073.t293 a_71281_n10073.n130 10.5154
R52741 a_71281_n10073.n134 a_71281_n10073.t293 10.5154
R52742 a_71281_n10073.t101 a_71281_n10073.n116 10.5154
R52743 a_71281_n10073.n120 a_71281_n10073.t101 10.5154
R52744 a_71281_n10073.t94 a_71281_n10073.n99 10.5154
R52745 a_71281_n10073.n103 a_71281_n10073.t94 10.5154
R52746 a_71281_n10073.t161 a_71281_n10073.n85 10.5154
R52747 a_71281_n10073.n89 a_71281_n10073.t161 10.5154
R52748 a_71281_n10073.t300 a_71281_n10073.n71 10.5154
R52749 a_71281_n10073.n75 a_71281_n10073.t300 10.5154
R52750 a_71281_n10073.t106 a_71281_n10073.n58 10.5154
R52751 a_71281_n10073.n62 a_71281_n10073.t106 10.5154
R52752 a_71281_n10073.t108 a_71281_n10073.n3 10.5154
R52753 a_71281_n10073.n7 a_71281_n10073.t108 10.5154
R52754 a_71281_n10073.n221 a_71281_n10073.t177 10.5154
R52755 a_71281_n10073.t177 a_71281_n10073.n216 10.5154
R52756 a_71281_n10073.n235 a_71281_n10073.t172 10.5154
R52757 a_71281_n10073.t172 a_71281_n10073.n230 10.5154
R52758 a_71281_n10073.n249 a_71281_n10073.t247 10.5154
R52759 a_71281_n10073.t247 a_71281_n10073.n244 10.5154
R52760 a_71281_n10073.n266 a_71281_n10073.t231 10.5154
R52761 a_71281_n10073.t231 a_71281_n10073.n261 10.5154
R52762 a_71281_n10073.n280 a_71281_n10073.t316 10.5154
R52763 a_71281_n10073.t316 a_71281_n10073.n275 10.5154
R52764 a_71281_n10073.n297 a_71281_n10073.t284 10.5154
R52765 a_71281_n10073.t284 a_71281_n10073.n292 10.5154
R52766 a_71281_n10073.n311 a_71281_n10073.t89 10.5154
R52767 a_71281_n10073.t89 a_71281_n10073.n306 10.5154
R52768 a_71281_n10073.n325 a_71281_n10073.t83 10.5154
R52769 a_71281_n10073.t83 a_71281_n10073.n320 10.5154
R52770 a_71281_n10073.n339 a_71281_n10073.t149 10.5154
R52771 a_71281_n10073.t149 a_71281_n10073.n334 10.5154
R52772 a_71281_n10073.t243 a_71281_n10073.n465 10.5154
R52773 a_71281_n10073.n469 a_71281_n10073.t243 10.5154
R52774 a_71281_n10073.t207 a_71281_n10073.n451 10.5154
R52775 a_71281_n10073.n455 a_71281_n10073.t207 10.5154
R52776 a_71281_n10073.t219 a_71281_n10073.n437 10.5154
R52777 a_71281_n10073.n441 a_71281_n10073.t219 10.5154
R52778 a_71281_n10073.t206 a_71281_n10073.n420 10.5154
R52779 a_71281_n10073.n424 a_71281_n10073.t206 10.5154
R52780 a_71281_n10073.t286 a_71281_n10073.n406 10.5154
R52781 a_71281_n10073.n410 a_71281_n10073.t286 10.5154
R52782 a_71281_n10073.t280 a_71281_n10073.n389 10.5154
R52783 a_71281_n10073.n393 a_71281_n10073.t280 10.5154
R52784 a_71281_n10073.t87 a_71281_n10073.n375 10.5154
R52785 a_71281_n10073.n379 a_71281_n10073.t87 10.5154
R52786 a_71281_n10073.t212 a_71281_n10073.n361 10.5154
R52787 a_71281_n10073.n365 a_71281_n10073.t212 10.5154
R52788 a_71281_n10073.t291 a_71281_n10073.n348 10.5154
R52789 a_71281_n10073.n352 a_71281_n10073.t291 10.5154
R52790 a_71281_n10073.t112 a_71281_n10073.n203 10.5154
R52791 a_71281_n10073.n207 a_71281_n10073.t112 10.5154
R52792 a_71281_n10073.n484 a_71281_n10073.t170 10.5154
R52793 a_71281_n10073.t170 a_71281_n10073.n479 10.5154
R52794 a_71281_n10073.n512 a_71281_n10073.t109 10.5154
R52795 a_71281_n10073.t109 a_71281_n10073.n507 10.5154
R52796 a_71281_n10073.n526 a_71281_n10073.t100 10.5154
R52797 a_71281_n10073.t100 a_71281_n10073.n521 10.5154
R52798 a_71281_n10073.n540 a_71281_n10073.t169 10.5154
R52799 a_71281_n10073.t169 a_71281_n10073.n535 10.5154
R52800 a_71281_n10073.n557 a_71281_n10073.t154 10.5154
R52801 a_71281_n10073.t154 a_71281_n10073.n552 10.5154
R52802 a_71281_n10073.n571 a_71281_n10073.t227 10.5154
R52803 a_71281_n10073.t227 a_71281_n10073.n566 10.5154
R52804 a_71281_n10073.n588 a_71281_n10073.t198 10.5154
R52805 a_71281_n10073.t198 a_71281_n10073.n583 10.5154
R52806 a_71281_n10073.n602 a_71281_n10073.t281 10.5154
R52807 a_71281_n10073.t281 a_71281_n10073.n597 10.5154
R52808 a_71281_n10073.n616 a_71281_n10073.t272 10.5154
R52809 a_71281_n10073.t272 a_71281_n10073.n611 10.5154
R52810 a_71281_n10073.n630 a_71281_n10073.t82 10.5154
R52811 a_71281_n10073.t82 a_71281_n10073.n625 10.5154
R52812 a_71281_n10073.t263 a_71281_n10073.n756 10.5154
R52813 a_71281_n10073.n760 a_71281_n10073.t263 10.5154
R52814 a_71281_n10073.t232 a_71281_n10073.n742 10.5154
R52815 a_71281_n10073.n746 a_71281_n10073.t232 10.5154
R52816 a_71281_n10073.t246 a_71281_n10073.n728 10.5154
R52817 a_71281_n10073.n732 a_71281_n10073.t246 10.5154
R52818 a_71281_n10073.t230 a_71281_n10073.n711 10.5154
R52819 a_71281_n10073.n715 a_71281_n10073.t230 10.5154
R52820 a_71281_n10073.t315 a_71281_n10073.n697 10.5154
R52821 a_71281_n10073.n701 a_71281_n10073.t315 10.5154
R52822 a_71281_n10073.t302 a_71281_n10073.n680 10.5154
R52823 a_71281_n10073.n684 a_71281_n10073.t302 10.5154
R52824 a_71281_n10073.t107 a_71281_n10073.n666 10.5154
R52825 a_71281_n10073.n670 a_71281_n10073.t107 10.5154
R52826 a_71281_n10073.t237 a_71281_n10073.n652 10.5154
R52827 a_71281_n10073.n656 a_71281_n10073.t237 10.5154
R52828 a_71281_n10073.t319 a_71281_n10073.n639 10.5154
R52829 a_71281_n10073.n643 a_71281_n10073.t319 10.5154
R52830 a_71281_n10073.t304 a_71281_n10073.n494 10.5154
R52831 a_71281_n10073.n498 a_71281_n10073.t304 10.5154
R52832 a_71281_n10073.n775 a_71281_n10073.t184 10.5154
R52833 a_71281_n10073.t184 a_71281_n10073.n770 10.5154
R52834 a_71281_n10073.n194 a_71281_n10073.t251 10.5154
R52835 a_71281_n10073.t251 a_71281_n10073.n189 10.5154
R52836 a_71281_n10073.n789 a_71281_n10073.t214 10.515
R52837 a_71281_n10073.n59 a_71281_n10073.t126 10.515
R52838 a_71281_n10073.n336 a_71281_n10073.t218 10.515
R52839 a_71281_n10073.n349 a_71281_n10073.t325 10.515
R52840 a_71281_n10073.n627 a_71281_n10073.t181 10.515
R52841 a_71281_n10073.n640 a_71281_n10073.t202 10.515
R52842 a_71281_n10073.n17 a_71281_n10073.t254 10.515
R52843 a_71281_n10073.n18 a_71281_n10073.t254 10.515
R52844 a_71281_n10073.n31 a_71281_n10073.t241 10.515
R52845 a_71281_n10073.n32 a_71281_n10073.t241 10.515
R52846 a_71281_n10073.n45 a_71281_n10073.t321 10.515
R52847 a_71281_n10073.n46 a_71281_n10073.t321 10.515
R52848 a_71281_n10073.n863 a_71281_n10073.t312 10.515
R52849 a_71281_n10073.n862 a_71281_n10073.t312 10.515
R52850 a_71281_n10073.n849 a_71281_n10073.t114 10.515
R52851 a_71281_n10073.n848 a_71281_n10073.t114 10.515
R52852 a_71281_n10073.n832 a_71281_n10073.t86 10.515
R52853 a_71281_n10073.n831 a_71281_n10073.t86 10.515
R52854 a_71281_n10073.n818 a_71281_n10073.t152 10.515
R52855 a_71281_n10073.n817 a_71281_n10073.t152 10.515
R52856 a_71281_n10073.n804 a_71281_n10073.t148 10.515
R52857 a_71281_n10073.n803 a_71281_n10073.t148 10.515
R52858 a_71281_n10073.n790 a_71281_n10073.t214 10.515
R52859 a_71281_n10073.n177 a_71281_n10073.t76 10.515
R52860 a_71281_n10073.n176 a_71281_n10073.t76 10.515
R52861 a_71281_n10073.n163 a_71281_n10073.t329 10.515
R52862 a_71281_n10073.n162 a_71281_n10073.t329 10.515
R52863 a_71281_n10073.n149 a_71281_n10073.t336 10.515
R52864 a_71281_n10073.n148 a_71281_n10073.t336 10.515
R52865 a_71281_n10073.n132 a_71281_n10073.t328 10.515
R52866 a_71281_n10073.n131 a_71281_n10073.t328 10.515
R52867 a_71281_n10073.n118 a_71281_n10073.t124 10.515
R52868 a_71281_n10073.n117 a_71281_n10073.t124 10.515
R52869 a_71281_n10073.n101 a_71281_n10073.t119 10.515
R52870 a_71281_n10073.n100 a_71281_n10073.t119 10.515
R52871 a_71281_n10073.n87 a_71281_n10073.t183 10.515
R52872 a_71281_n10073.n86 a_71281_n10073.t183 10.515
R52873 a_71281_n10073.n73 a_71281_n10073.t333 10.515
R52874 a_71281_n10073.n72 a_71281_n10073.t333 10.515
R52875 a_71281_n10073.n60 a_71281_n10073.t126 10.515
R52876 a_71281_n10073.n5 a_71281_n10073.t174 10.515
R52877 a_71281_n10073.n4 a_71281_n10073.t174 10.515
R52878 a_71281_n10073.n217 a_71281_n10073.t259 10.515
R52879 a_71281_n10073.n218 a_71281_n10073.t259 10.515
R52880 a_71281_n10073.n231 a_71281_n10073.t250 10.515
R52881 a_71281_n10073.n232 a_71281_n10073.t250 10.515
R52882 a_71281_n10073.n245 a_71281_n10073.t327 10.515
R52883 a_71281_n10073.n246 a_71281_n10073.t327 10.515
R52884 a_71281_n10073.n262 a_71281_n10073.t317 10.515
R52885 a_71281_n10073.n263 a_71281_n10073.t317 10.515
R52886 a_71281_n10073.n276 a_71281_n10073.t118 10.515
R52887 a_71281_n10073.n277 a_71281_n10073.t118 10.515
R52888 a_71281_n10073.n293 a_71281_n10073.t93 10.515
R52889 a_71281_n10073.n294 a_71281_n10073.t93 10.515
R52890 a_71281_n10073.n307 a_71281_n10073.t159 10.515
R52891 a_71281_n10073.n308 a_71281_n10073.t159 10.515
R52892 a_71281_n10073.n321 a_71281_n10073.t150 10.515
R52893 a_71281_n10073.n322 a_71281_n10073.t150 10.515
R52894 a_71281_n10073.n335 a_71281_n10073.t218 10.515
R52895 a_71281_n10073.n467 a_71281_n10073.t264 10.515
R52896 a_71281_n10073.n466 a_71281_n10073.t264 10.515
R52897 a_71281_n10073.n453 a_71281_n10073.t242 10.515
R52898 a_71281_n10073.n452 a_71281_n10073.t242 10.515
R52899 a_71281_n10073.n439 a_71281_n10073.t253 10.515
R52900 a_71281_n10073.n438 a_71281_n10073.t253 10.515
R52901 a_71281_n10073.n422 a_71281_n10073.t240 10.515
R52902 a_71281_n10073.n421 a_71281_n10073.t240 10.515
R52903 a_71281_n10073.n408 a_71281_n10073.t320 10.515
R52904 a_71281_n10073.n407 a_71281_n10073.t320 10.515
R52905 a_71281_n10073.n391 a_71281_n10073.t311 10.515
R52906 a_71281_n10073.n390 a_71281_n10073.t311 10.515
R52907 a_71281_n10073.n377 a_71281_n10073.t113 10.515
R52908 a_71281_n10073.n376 a_71281_n10073.t113 10.515
R52909 a_71281_n10073.n363 a_71281_n10073.t249 10.515
R52910 a_71281_n10073.n362 a_71281_n10073.t249 10.515
R52911 a_71281_n10073.n350 a_71281_n10073.t325 10.515
R52912 a_71281_n10073.n205 a_71281_n10073.t178 10.515
R52913 a_71281_n10073.n204 a_71281_n10073.t178 10.515
R52914 a_71281_n10073.n480 a_71281_n10073.t186 10.515
R52915 a_71281_n10073.n481 a_71281_n10073.t186 10.515
R52916 a_71281_n10073.n508 a_71281_n10073.t195 10.515
R52917 a_71281_n10073.n509 a_71281_n10073.t195 10.515
R52918 a_71281_n10073.n522 a_71281_n10073.t189 10.515
R52919 a_71281_n10073.n523 a_71281_n10073.t189 10.515
R52920 a_71281_n10073.n536 a_71281_n10073.t270 10.515
R52921 a_71281_n10073.n537 a_71281_n10073.t270 10.515
R52922 a_71281_n10073.n553 a_71281_n10073.t267 10.515
R52923 a_71281_n10073.n554 a_71281_n10073.t267 10.515
R52924 a_71281_n10073.n567 a_71281_n10073.t74 10.515
R52925 a_71281_n10073.n568 a_71281_n10073.t74 10.515
R52926 a_71281_n10073.n584 a_71281_n10073.t323 10.515
R52927 a_71281_n10073.n585 a_71281_n10073.t323 10.515
R52928 a_71281_n10073.n598 a_71281_n10073.t122 10.515
R52929 a_71281_n10073.n599 a_71281_n10073.t122 10.515
R52930 a_71281_n10073.n612 a_71281_n10073.t117 10.515
R52931 a_71281_n10073.n613 a_71281_n10073.t117 10.515
R52932 a_71281_n10073.n626 a_71281_n10073.t181 10.515
R52933 a_71281_n10073.n758 a_71281_n10073.t157 10.515
R52934 a_71281_n10073.n757 a_71281_n10073.t157 10.515
R52935 a_71281_n10073.n744 a_71281_n10073.t135 10.515
R52936 a_71281_n10073.n743 a_71281_n10073.t135 10.515
R52937 a_71281_n10073.n730 a_71281_n10073.t145 10.515
R52938 a_71281_n10073.n729 a_71281_n10073.t145 10.515
R52939 a_71281_n10073.n713 a_71281_n10073.t132 10.515
R52940 a_71281_n10073.n712 a_71281_n10073.t132 10.515
R52941 a_71281_n10073.n699 a_71281_n10073.t200 10.515
R52942 a_71281_n10073.n698 a_71281_n10073.t200 10.515
R52943 a_71281_n10073.n682 a_71281_n10073.t192 10.515
R52944 a_71281_n10073.n681 a_71281_n10073.t192 10.515
R52945 a_71281_n10073.n668 a_71281_n10073.t274 10.515
R52946 a_71281_n10073.n667 a_71281_n10073.t274 10.515
R52947 a_71281_n10073.n654 a_71281_n10073.t138 10.515
R52948 a_71281_n10073.n653 a_71281_n10073.t138 10.515
R52949 a_71281_n10073.n641 a_71281_n10073.t202 10.515
R52950 a_71281_n10073.n496 a_71281_n10073.t130 10.515
R52951 a_71281_n10073.n495 a_71281_n10073.t130 10.515
R52952 a_71281_n10073.n771 a_71281_n10073.t92 10.515
R52953 a_71281_n10073.n772 a_71281_n10073.t92 10.515
R52954 a_71281_n10073.n190 a_71281_n10073.t268 10.515
R52955 a_71281_n10073.n191 a_71281_n10073.t268 10.515
R52956 a_71281_n10073.n21 a_71281_n10073.t121 9.57886
R52957 a_71281_n10073.t121 a_71281_n10073.n16 9.57886
R52958 a_71281_n10073.n18 a_71281_n10073.t313 9.57886
R52959 a_71281_n10073.t313 a_71281_n10073.n17 9.57886
R52960 a_71281_n10073.n35 a_71281_n10073.t116 9.57886
R52961 a_71281_n10073.t116 a_71281_n10073.n30 9.57886
R52962 a_71281_n10073.n32 a_71281_n10073.t299 9.57886
R52963 a_71281_n10073.t299 a_71281_n10073.n31 9.57886
R52964 a_71281_n10073.n49 a_71281_n10073.t180 9.57886
R52965 a_71281_n10073.t180 a_71281_n10073.n44 9.57886
R52966 a_71281_n10073.n46 a_71281_n10073.t105 9.57886
R52967 a_71281_n10073.t105 a_71281_n10073.n45 9.57886
R52968 a_71281_n10073.t44 a_71281_n10073.n861 9.57886
R52969 a_71281_n10073.n865 a_71281_n10073.t44 9.57886
R52970 a_71281_n10073.t72 a_71281_n10073.n862 9.57886
R52971 a_71281_n10073.n863 a_71281_n10073.t72 9.57886
R52972 a_71281_n10073.t16 a_71281_n10073.n847 9.57886
R52973 a_71281_n10073.n851 a_71281_n10073.t16 9.57886
R52974 a_71281_n10073.t48 a_71281_n10073.n848 9.57886
R52975 a_71281_n10073.n849 a_71281_n10073.t48 9.57886
R52976 a_71281_n10073.t215 a_71281_n10073.n830 9.57886
R52977 a_71281_n10073.n834 a_71281_n10073.t215 9.57886
R52978 a_71281_n10073.t139 a_71281_n10073.n831 9.57886
R52979 a_71281_n10073.n832 a_71281_n10073.t139 9.57886
R52980 a_71281_n10073.t297 a_71281_n10073.n816 9.57886
R52981 a_71281_n10073.n820 a_71281_n10073.t297 9.57886
R52982 a_71281_n10073.t203 a_71281_n10073.n817 9.57886
R52983 a_71281_n10073.n818 a_71281_n10073.t203 9.57886
R52984 a_71281_n10073.t285 a_71281_n10073.n802 9.57886
R52985 a_71281_n10073.n806 a_71281_n10073.t285 9.57886
R52986 a_71281_n10073.t196 a_71281_n10073.n803 9.57886
R52987 a_71281_n10073.n804 a_71281_n10073.t196 9.57886
R52988 a_71281_n10073.t98 a_71281_n10073.n788 9.57886
R52989 a_71281_n10073.n792 a_71281_n10073.t98 9.57886
R52990 a_71281_n10073.t277 a_71281_n10073.n789 9.57886
R52991 a_71281_n10073.n790 a_71281_n10073.t277 9.57886
R52992 a_71281_n10073.t142 a_71281_n10073.n175 9.57886
R52993 a_71281_n10073.n179 a_71281_n10073.t142 9.57886
R52994 a_71281_n10073.t238 a_71281_n10073.n176 9.57886
R52995 a_71281_n10073.n177 a_71281_n10073.t238 9.57886
R52996 a_71281_n10073.t127 a_71281_n10073.n161 9.57886
R52997 a_71281_n10073.n165 a_71281_n10073.t127 9.57886
R52998 a_71281_n10073.t204 a_71281_n10073.n162 9.57886
R52999 a_71281_n10073.n163 a_71281_n10073.t204 9.57886
R53000 a_71281_n10073.t129 a_71281_n10073.n147 9.57886
R53001 a_71281_n10073.n151 a_71281_n10073.t129 9.57886
R53002 a_71281_n10073.t216 a_71281_n10073.n148 9.57886
R53003 a_71281_n10073.n149 a_71281_n10073.t216 9.57886
R53004 a_71281_n10073.t60 a_71281_n10073.n130 9.57886
R53005 a_71281_n10073.n134 a_71281_n10073.t60 9.57886
R53006 a_71281_n10073.t30 a_71281_n10073.n131 9.57886
R53007 a_71281_n10073.n132 a_71281_n10073.t30 9.57886
R53008 a_71281_n10073.t38 a_71281_n10073.n116 9.57886
R53009 a_71281_n10073.n120 a_71281_n10073.t38 9.57886
R53010 a_71281_n10073.t14 a_71281_n10073.n117 9.57886
R53011 a_71281_n10073.n118 a_71281_n10073.t14 9.57886
R53012 a_71281_n10073.t187 a_71281_n10073.n99 9.57886
R53013 a_71281_n10073.n103 a_71281_n10073.t187 9.57886
R53014 a_71281_n10073.t278 a_71281_n10073.n100 9.57886
R53015 a_71281_n10073.n101 a_71281_n10073.t278 9.57886
R53016 a_71281_n10073.t265 a_71281_n10073.n85 9.57886
R53017 a_71281_n10073.n89 a_71281_n10073.t265 9.57886
R53018 a_71281_n10073.t84 a_71281_n10073.n86 9.57886
R53019 a_71281_n10073.n87 a_71281_n10073.t84 9.57886
R53020 a_71281_n10073.t128 a_71281_n10073.n71 9.57886
R53021 a_71281_n10073.n75 a_71281_n10073.t128 9.57886
R53022 a_71281_n10073.t210 a_71281_n10073.n72 9.57886
R53023 a_71281_n10073.n73 a_71281_n10073.t210 9.57886
R53024 a_71281_n10073.t190 a_71281_n10073.n58 9.57886
R53025 a_71281_n10073.n62 a_71281_n10073.t190 9.57886
R53026 a_71281_n10073.t288 a_71281_n10073.n59 9.57886
R53027 a_71281_n10073.n60 a_71281_n10073.t288 9.57886
R53028 a_71281_n10073.t322 a_71281_n10073.n3 9.57886
R53029 a_71281_n10073.n7 a_71281_n10073.t322 9.57886
R53030 a_71281_n10073.t228 a_71281_n10073.n4 9.57886
R53031 a_71281_n10073.n5 a_71281_n10073.t228 9.57886
R53032 a_71281_n10073.n221 a_71281_n10073.t185 9.57886
R53033 a_71281_n10073.t185 a_71281_n10073.n216 9.57886
R53034 a_71281_n10073.n218 a_71281_n10073.t318 9.57886
R53035 a_71281_n10073.t318 a_71281_n10073.n217 9.57886
R53036 a_71281_n10073.n235 a_71281_n10073.t179 9.57886
R53037 a_71281_n10073.t179 a_71281_n10073.n230 9.57886
R53038 a_71281_n10073.n232 a_71281_n10073.t305 9.57886
R53039 a_71281_n10073.t305 a_71281_n10073.n231 9.57886
R53040 a_71281_n10073.n249 a_71281_n10073.t260 9.57886
R53041 a_71281_n10073.t260 a_71281_n10073.n244 9.57886
R53042 a_71281_n10073.n246 a_71281_n10073.t110 9.57886
R53043 a_71281_n10073.t110 a_71281_n10073.n245 9.57886
R53044 a_71281_n10073.n266 a_71281_n10073.t18 9.57886
R53045 a_71281_n10073.t18 a_71281_n10073.n261 9.57886
R53046 a_71281_n10073.n263 a_71281_n10073.t68 9.57886
R53047 a_71281_n10073.t68 a_71281_n10073.n262 9.57886
R53048 a_71281_n10073.n280 a_71281_n10073.t2 9.57886
R53049 a_71281_n10073.t2 a_71281_n10073.n275 9.57886
R53050 a_71281_n10073.n277 a_71281_n10073.t46 9.57886
R53051 a_71281_n10073.t46 a_71281_n10073.n276 9.57886
R53052 a_71281_n10073.n297 a_71281_n10073.t295 9.57886
R53053 a_71281_n10073.t295 a_71281_n10073.n292 9.57886
R53054 a_71281_n10073.n294 a_71281_n10073.t143 9.57886
R53055 a_71281_n10073.t143 a_71281_n10073.n293 9.57886
R53056 a_71281_n10073.n311 a_71281_n10073.t102 9.57886
R53057 a_71281_n10073.t102 a_71281_n10073.n306 9.57886
R53058 a_71281_n10073.n308 a_71281_n10073.t209 9.57886
R53059 a_71281_n10073.t209 a_71281_n10073.n307 9.57886
R53060 a_71281_n10073.n325 a_71281_n10073.t95 9.57886
R53061 a_71281_n10073.t95 a_71281_n10073.n320 9.57886
R53062 a_71281_n10073.n322 a_71281_n10073.t199 9.57886
R53063 a_71281_n10073.t199 a_71281_n10073.n321 9.57886
R53064 a_71281_n10073.n339 a_71281_n10073.t162 9.57886
R53065 a_71281_n10073.t162 a_71281_n10073.n334 9.57886
R53066 a_71281_n10073.n336 a_71281_n10073.t283 9.57886
R53067 a_71281_n10073.t283 a_71281_n10073.n335 9.57886
R53068 a_71281_n10073.t256 a_71281_n10073.n465 9.57886
R53069 a_71281_n10073.n469 a_71281_n10073.t256 9.57886
R53070 a_71281_n10073.t156 a_71281_n10073.n466 9.57886
R53071 a_71281_n10073.n467 a_71281_n10073.t156 9.57886
R53072 a_71281_n10073.t222 a_71281_n10073.n451 9.57886
R53073 a_71281_n10073.n455 a_71281_n10073.t222 9.57886
R53074 a_71281_n10073.t133 a_71281_n10073.n452 9.57886
R53075 a_71281_n10073.n453 a_71281_n10073.t133 9.57886
R53076 a_71281_n10073.t234 a_71281_n10073.n437 9.57886
R53077 a_71281_n10073.n441 a_71281_n10073.t234 9.57886
R53078 a_71281_n10073.t144 a_71281_n10073.n438 9.57886
R53079 a_71281_n10073.n439 a_71281_n10073.t144 9.57886
R53080 a_71281_n10073.t26 a_71281_n10073.n420 9.57886
R53081 a_71281_n10073.n424 a_71281_n10073.t26 9.57886
R53082 a_71281_n10073.t56 a_71281_n10073.n421 9.57886
R53083 a_71281_n10073.n422 a_71281_n10073.t56 9.57886
R53084 a_71281_n10073.t6 a_71281_n10073.n406 9.57886
R53085 a_71281_n10073.n410 a_71281_n10073.t6 9.57886
R53086 a_71281_n10073.t34 a_71281_n10073.n407 9.57886
R53087 a_71281_n10073.n408 a_71281_n10073.t34 9.57886
R53088 a_71281_n10073.t287 a_71281_n10073.n389 9.57886
R53089 a_71281_n10073.n393 a_71281_n10073.t287 9.57886
R53090 a_71281_n10073.t191 a_71281_n10073.n390 9.57886
R53091 a_71281_n10073.n391 a_71281_n10073.t191 9.57886
R53092 a_71281_n10073.t99 a_71281_n10073.n375 9.57886
R53093 a_71281_n10073.n379 a_71281_n10073.t99 9.57886
R53094 a_71281_n10073.t273 a_71281_n10073.n376 9.57886
R53095 a_71281_n10073.n377 a_71281_n10073.t273 9.57886
R53096 a_71281_n10073.t224 a_71281_n10073.n361 9.57886
R53097 a_71281_n10073.n365 a_71281_n10073.t224 9.57886
R53098 a_71281_n10073.t137 a_71281_n10073.n362 9.57886
R53099 a_71281_n10073.n363 a_71281_n10073.t137 9.57886
R53100 a_71281_n10073.t308 a_71281_n10073.n348 9.57886
R53101 a_71281_n10073.n352 a_71281_n10073.t308 9.57886
R53102 a_71281_n10073.t201 a_71281_n10073.n349 9.57886
R53103 a_71281_n10073.n350 a_71281_n10073.t201 9.57886
R53104 a_71281_n10073.t120 a_71281_n10073.n203 9.57886
R53105 a_71281_n10073.n207 a_71281_n10073.t120 9.57886
R53106 a_71281_n10073.t235 a_71281_n10073.n204 9.57886
R53107 a_71281_n10073.n205 a_71281_n10073.t235 9.57886
R53108 a_71281_n10073.n484 a_71281_n10073.t175 9.57886
R53109 a_71281_n10073.t175 a_71281_n10073.n479 9.57886
R53110 a_71281_n10073.n481 a_71281_n10073.t91 9.57886
R53111 a_71281_n10073.t91 a_71281_n10073.n480 9.57886
R53112 a_71281_n10073.n512 a_71281_n10073.t80 9.57886
R53113 a_71281_n10073.t80 a_71281_n10073.n507 9.57886
R53114 a_71281_n10073.n509 a_71281_n10073.t233 9.57886
R53115 a_71281_n10073.t233 a_71281_n10073.n508 9.57886
R53116 a_71281_n10073.n526 a_71281_n10073.t75 9.57886
R53117 a_71281_n10073.t75 a_71281_n10073.n521 9.57886
R53118 a_71281_n10073.n523 a_71281_n10073.t220 9.57886
R53119 a_71281_n10073.t220 a_71281_n10073.n522 9.57886
R53120 a_71281_n10073.n540 a_71281_n10073.t134 9.57886
R53121 a_71281_n10073.t134 a_71281_n10073.n535 9.57886
R53122 a_71281_n10073.n537 a_71281_n10073.t303 9.57886
R53123 a_71281_n10073.t303 a_71281_n10073.n536 9.57886
R53124 a_71281_n10073.n557 a_71281_n10073.t58 9.57886
R53125 a_71281_n10073.t58 a_71281_n10073.n552 9.57886
R53126 a_71281_n10073.n554 a_71281_n10073.t12 9.57886
R53127 a_71281_n10073.t12 a_71281_n10073.n553 9.57886
R53128 a_71281_n10073.n571 a_71281_n10073.t36 9.57886
R53129 a_71281_n10073.t36 a_71281_n10073.n566 9.57886
R53130 a_71281_n10073.n568 a_71281_n10073.t70 9.57886
R53131 a_71281_n10073.t70 a_71281_n10073.n567 9.57886
R53132 a_71281_n10073.n588 a_71281_n10073.t182 9.57886
R53133 a_71281_n10073.t182 a_71281_n10073.n583 9.57886
R53134 a_71281_n10073.n585 a_71281_n10073.t77 9.57886
R53135 a_71281_n10073.t77 a_71281_n10073.n584 9.57886
R53136 a_71281_n10073.n602 a_71281_n10073.t262 9.57886
R53137 a_71281_n10073.t262 a_71281_n10073.n597 9.57886
R53138 a_71281_n10073.n599 a_71281_n10073.t141 9.57886
R53139 a_71281_n10073.t141 a_71281_n10073.n598 9.57886
R53140 a_71281_n10073.n616 a_71281_n10073.t255 9.57886
R53141 a_71281_n10073.t255 a_71281_n10073.n611 9.57886
R53142 a_71281_n10073.n613 a_71281_n10073.t131 9.57886
R53143 a_71281_n10073.t131 a_71281_n10073.n612 9.57886
R53144 a_71281_n10073.n630 a_71281_n10073.t334 9.57886
R53145 a_71281_n10073.t334 a_71281_n10073.n625 9.57886
R53146 a_71281_n10073.n627 a_71281_n10073.t197 9.57886
R53147 a_71281_n10073.t197 a_71281_n10073.n626 9.57886
R53148 a_71281_n10073.t244 a_71281_n10073.n756 9.57886
R53149 a_71281_n10073.n760 a_71281_n10073.t244 9.57886
R53150 a_71281_n10073.t176 a_71281_n10073.n757 9.57886
R53151 a_71281_n10073.n758 a_71281_n10073.t176 9.57886
R53152 a_71281_n10073.t208 a_71281_n10073.n742 9.57886
R53153 a_71281_n10073.n746 a_71281_n10073.t208 9.57886
R53154 a_71281_n10073.t151 a_71281_n10073.n743 9.57886
R53155 a_71281_n10073.n744 a_71281_n10073.t151 9.57886
R53156 a_71281_n10073.t221 a_71281_n10073.n728 9.57886
R53157 a_71281_n10073.n732 a_71281_n10073.t221 9.57886
R53158 a_71281_n10073.t165 a_71281_n10073.n729 9.57886
R53159 a_71281_n10073.n730 a_71281_n10073.t165 9.57886
R53160 a_71281_n10073.t28 a_71281_n10073.n711 9.57886
R53161 a_71281_n10073.n715 a_71281_n10073.t28 9.57886
R53162 a_71281_n10073.t50 a_71281_n10073.n712 9.57886
R53163 a_71281_n10073.n713 a_71281_n10073.t50 9.57886
R53164 a_71281_n10073.t10 a_71281_n10073.n697 9.57886
R53165 a_71281_n10073.n701 a_71281_n10073.t10 9.57886
R53166 a_71281_n10073.t22 a_71281_n10073.n698 9.57886
R53167 a_71281_n10073.n699 a_71281_n10073.t22 9.57886
R53168 a_71281_n10073.t282 a_71281_n10073.n680 9.57886
R53169 a_71281_n10073.n684 a_71281_n10073.t282 9.57886
R53170 a_71281_n10073.t211 a_71281_n10073.n681 9.57886
R53171 a_71281_n10073.n682 a_71281_n10073.t211 9.57886
R53172 a_71281_n10073.t88 a_71281_n10073.n666 9.57886
R53173 a_71281_n10073.n670 a_71281_n10073.t88 9.57886
R53174 a_71281_n10073.t289 a_71281_n10073.n667 9.57886
R53175 a_71281_n10073.n668 a_71281_n10073.t289 9.57886
R53176 a_71281_n10073.t213 a_71281_n10073.n652 9.57886
R53177 a_71281_n10073.n656 a_71281_n10073.t213 9.57886
R53178 a_71281_n10073.t153 a_71281_n10073.n653 9.57886
R53179 a_71281_n10073.n654 a_71281_n10073.t153 9.57886
R53180 a_71281_n10073.t292 a_71281_n10073.n639 9.57886
R53181 a_71281_n10073.n643 a_71281_n10073.t292 9.57886
R53182 a_71281_n10073.t226 a_71281_n10073.n640 9.57886
R53183 a_71281_n10073.n641 a_71281_n10073.t226 9.57886
R53184 a_71281_n10073.t271 a_71281_n10073.n494 9.57886
R53185 a_71281_n10073.n498 a_71281_n10073.t271 9.57886
R53186 a_71281_n10073.t160 a_71281_n10073.n495 9.57886
R53187 a_71281_n10073.n496 a_71281_n10073.t160 9.57886
R53188 a_71281_n10073.n775 a_71281_n10073.t171 9.57886
R53189 a_71281_n10073.t171 a_71281_n10073.n770 9.57886
R53190 a_71281_n10073.n772 a_71281_n10073.t111 9.57886
R53191 a_71281_n10073.t111 a_71281_n10073.n771 9.57886
R53192 a_71281_n10073.n194 a_71281_n10073.t79 9.57886
R53193 a_71281_n10073.t79 a_71281_n10073.n189 9.57886
R53194 a_71281_n10073.n191 a_71281_n10073.t167 9.57886
R53195 a_71281_n10073.t167 a_71281_n10073.n190 9.57886
R53196 a_71281_n10073.t337 a_71281_n10073.n23 8.10567
R53197 a_71281_n10073.n24 a_71281_n10073.t337 8.10567
R53198 a_71281_n10073.t332 a_71281_n10073.n37 8.10567
R53199 a_71281_n10073.n38 a_71281_n10073.t332 8.10567
R53200 a_71281_n10073.t125 a_71281_n10073.n51 8.10567
R53201 a_71281_n10073.n52 a_71281_n10073.t125 8.10567
R53202 a_71281_n10073.n869 a_71281_n10073.t62 8.10567
R53203 a_71281_n10073.t62 a_71281_n10073.n868 8.10567
R53204 a_71281_n10073.n855 a_71281_n10073.t40 8.10567
R53205 a_71281_n10073.t40 a_71281_n10073.n854 8.10567
R53206 a_71281_n10073.n838 a_71281_n10073.t166 8.10567
R53207 a_71281_n10073.t166 a_71281_n10073.n837 8.10567
R53208 a_71281_n10073.n824 a_71281_n10073.t236 8.10567
R53209 a_71281_n10073.t236 a_71281_n10073.n823 8.10567
R53210 a_71281_n10073.n810 a_71281_n10073.t223 8.10567
R53211 a_71281_n10073.t223 a_71281_n10073.n809 8.10567
R53212 a_71281_n10073.n796 a_71281_n10073.t307 8.10567
R53213 a_71281_n10073.t307 a_71281_n10073.n795 8.10567
R53214 a_71281_n10073.n183 a_71281_n10073.t324 8.10567
R53215 a_71281_n10073.t324 a_71281_n10073.n182 8.10567
R53216 a_71281_n10073.n169 a_71281_n10073.t290 8.10567
R53217 a_71281_n10073.t290 a_71281_n10073.n168 8.10567
R53218 a_71281_n10073.n155 a_71281_n10073.t306 8.10567
R53219 a_71281_n10073.t306 a_71281_n10073.n154 8.10567
R53220 a_71281_n10073.n138 a_71281_n10073.t8 8.10567
R53221 a_71281_n10073.t8 a_71281_n10073.n137 8.10567
R53222 a_71281_n10073.n124 a_71281_n10073.t66 8.10567
R53223 a_71281_n10073.t66 a_71281_n10073.n123 8.10567
R53224 a_71281_n10073.n107 a_71281_n10073.t90 8.10567
R53225 a_71281_n10073.t90 a_71281_n10073.n106 8.10567
R53226 a_71281_n10073.n93 a_71281_n10073.t155 8.10567
R53227 a_71281_n10073.t155 a_71281_n10073.n92 8.10567
R53228 a_71281_n10073.n79 a_71281_n10073.t298 8.10567
R53229 a_71281_n10073.t298 a_71281_n10073.n78 8.10567
R53230 a_71281_n10073.n65 a_71281_n10073.t104 8.10567
R53231 a_71281_n10073.t104 a_71281_n10073.n64 8.10567
R53232 a_71281_n10073.n10 a_71281_n10073.t261 8.10567
R53233 a_71281_n10073.t261 a_71281_n10073.n9 8.10567
R53234 a_71281_n10073.t103 a_71281_n10073.n223 8.10567
R53235 a_71281_n10073.n224 a_71281_n10073.t103 8.10567
R53236 a_71281_n10073.t96 a_71281_n10073.n237 8.10567
R53237 a_71281_n10073.n238 a_71281_n10073.t96 8.10567
R53238 a_71281_n10073.t163 a_71281_n10073.n251 8.10567
R53239 a_71281_n10073.n252 a_71281_n10073.t163 8.10567
R53240 a_71281_n10073.t52 a_71281_n10073.n268 8.10567
R53241 a_71281_n10073.n269 a_71281_n10073.t52 8.10567
R53242 a_71281_n10073.t24 a_71281_n10073.n282 8.10567
R53243 a_71281_n10073.n283 a_71281_n10073.t24 8.10567
R53244 a_71281_n10073.t194 a_71281_n10073.n299 8.10567
R53245 a_71281_n10073.n300 a_71281_n10073.t194 8.10567
R53246 a_71281_n10073.t276 a_71281_n10073.n313 8.10567
R53247 a_71281_n10073.n314 a_71281_n10073.t276 8.10567
R53248 a_71281_n10073.t269 a_71281_n10073.n327 8.10567
R53249 a_71281_n10073.n328 a_71281_n10073.t269 8.10567
R53250 a_71281_n10073.t78 a_71281_n10073.n341 8.10567
R53251 a_71281_n10073.n342 a_71281_n10073.t78 8.10567
R53252 a_71281_n10073.n473 a_71281_n10073.t266 8.10567
R53253 a_71281_n10073.t266 a_71281_n10073.n472 8.10567
R53254 a_71281_n10073.n459 a_71281_n10073.t245 8.10567
R53255 a_71281_n10073.t245 a_71281_n10073.n458 8.10567
R53256 a_71281_n10073.n445 a_71281_n10073.t257 8.10567
R53257 a_71281_n10073.t257 a_71281_n10073.n444 8.10567
R53258 a_71281_n10073.n428 a_71281_n10073.t20 8.10567
R53259 a_71281_n10073.t20 a_71281_n10073.n427 8.10567
R53260 a_71281_n10073.n414 a_71281_n10073.t4 8.10567
R53261 a_71281_n10073.t4 a_71281_n10073.n413 8.10567
R53262 a_71281_n10073.n397 a_71281_n10073.t314 8.10567
R53263 a_71281_n10073.t314 a_71281_n10073.n396 8.10567
R53264 a_71281_n10073.n383 a_71281_n10073.t115 8.10567
R53265 a_71281_n10073.t115 a_71281_n10073.n382 8.10567
R53266 a_71281_n10073.n369 a_71281_n10073.t252 8.10567
R53267 a_71281_n10073.t252 a_71281_n10073.n368 8.10567
R53268 a_71281_n10073.n355 a_71281_n10073.t331 8.10567
R53269 a_71281_n10073.t331 a_71281_n10073.n354 8.10567
R53270 a_71281_n10073.n210 a_71281_n10073.t296 8.10567
R53271 a_71281_n10073.t296 a_71281_n10073.n209 8.10567
R53272 a_71281_n10073.t188 a_71281_n10073.n486 8.10567
R53273 a_71281_n10073.n487 a_71281_n10073.t188 8.10567
R53274 a_71281_n10073.t335 a_71281_n10073.n514 8.10567
R53275 a_71281_n10073.n515 a_71281_n10073.t335 8.10567
R53276 a_71281_n10073.t326 a_71281_n10073.n528 8.10567
R53277 a_71281_n10073.n529 a_71281_n10073.t326 8.10567
R53278 a_71281_n10073.t123 a_71281_n10073.n542 8.10567
R53279 a_71281_n10073.n543 a_71281_n10073.t123 8.10567
R53280 a_71281_n10073.t64 a_71281_n10073.n559 8.10567
R53281 a_71281_n10073.n560 a_71281_n10073.t64 8.10567
R53282 a_71281_n10073.t42 a_71281_n10073.n573 8.10567
R53283 a_71281_n10073.n574 a_71281_n10073.t42 8.10567
R53284 a_71281_n10073.t158 a_71281_n10073.n590 8.10567
R53285 a_71281_n10073.n591 a_71281_n10073.t158 8.10567
R53286 a_71281_n10073.t229 a_71281_n10073.n604 8.10567
R53287 a_71281_n10073.n605 a_71281_n10073.t229 8.10567
R53288 a_71281_n10073.t217 a_71281_n10073.n618 8.10567
R53289 a_71281_n10073.n619 a_71281_n10073.t217 8.10567
R53290 a_71281_n10073.t301 a_71281_n10073.n632 8.10567
R53291 a_71281_n10073.n633 a_71281_n10073.t301 8.10567
R53292 a_71281_n10073.n764 a_71281_n10073.t164 8.10567
R53293 a_71281_n10073.t164 a_71281_n10073.n763 8.10567
R53294 a_71281_n10073.n750 a_71281_n10073.t136 8.10567
R53295 a_71281_n10073.t136 a_71281_n10073.n749 8.10567
R53296 a_71281_n10073.n736 a_71281_n10073.t147 8.10567
R53297 a_71281_n10073.t147 a_71281_n10073.n735 8.10567
R53298 a_71281_n10073.n719 a_71281_n10073.t54 8.10567
R53299 a_71281_n10073.t54 a_71281_n10073.n718 8.10567
R53300 a_71281_n10073.n705 a_71281_n10073.t32 8.10567
R53301 a_71281_n10073.t32 a_71281_n10073.n704 8.10567
R53302 a_71281_n10073.n688 a_71281_n10073.t193 8.10567
R53303 a_71281_n10073.t193 a_71281_n10073.n687 8.10567
R53304 a_71281_n10073.n674 a_71281_n10073.t275 8.10567
R53305 a_71281_n10073.t275 a_71281_n10073.n673 8.10567
R53306 a_71281_n10073.n660 a_71281_n10073.t140 8.10567
R53307 a_71281_n10073.t140 a_71281_n10073.n659 8.10567
R53308 a_71281_n10073.n646 a_71281_n10073.t205 8.10567
R53309 a_71281_n10073.t205 a_71281_n10073.n645 8.10567
R53310 a_71281_n10073.n501 a_71281_n10073.t258 8.10567
R53311 a_71281_n10073.t258 a_71281_n10073.n500 8.10567
R53312 a_71281_n10073.t97 a_71281_n10073.n777 8.10567
R53313 a_71281_n10073.n778 a_71281_n10073.t97 8.10567
R53314 a_71281_n10073.t248 a_71281_n10073.n196 8.10567
R53315 a_71281_n10073.n197 a_71281_n10073.t248 8.10567
R53316 a_71281_n10073.n143 a_71281_n10073.t61 6.12845
R53317 a_71281_n10073.n257 a_71281_n10073.t19 6.12845
R53318 a_71281_n10073.n433 a_71281_n10073.t27 6.12845
R53319 a_71281_n10073.n548 a_71281_n10073.t59 6.12845
R53320 a_71281_n10073.n724 a_71281_n10073.t29 6.12845
R53321 a_71281_n10073.n874 a_71281_n10073.t45 6.12845
R53322 a_71281_n10073.n843 a_71281_n10073.t49 6.12049
R53323 a_71281_n10073.n288 a_71281_n10073.t47 6.12049
R53324 a_71281_n10073.n402 a_71281_n10073.t35 6.12049
R53325 a_71281_n10073.n579 a_71281_n10073.t71 6.12049
R53326 a_71281_n10073.n693 a_71281_n10073.t23 6.12049
R53327 a_71281_n10073.n112 a_71281_n10073.t15 6.12049
R53328 a_71281_n10073.n23 a_71281_n10073.n19 4.64734
R53329 a_71281_n10073.n24 a_71281_n10073.n15 4.64734
R53330 a_71281_n10073.n37 a_71281_n10073.n33 4.64734
R53331 a_71281_n10073.n38 a_71281_n10073.n29 4.64734
R53332 a_71281_n10073.n51 a_71281_n10073.n47 4.64734
R53333 a_71281_n10073.n52 a_71281_n10073.n43 4.64734
R53334 a_71281_n10073.n869 a_71281_n10073.n860 4.64734
R53335 a_71281_n10073.n868 a_71281_n10073.n864 4.64734
R53336 a_71281_n10073.n855 a_71281_n10073.n846 4.64734
R53337 a_71281_n10073.n854 a_71281_n10073.n850 4.64734
R53338 a_71281_n10073.n838 a_71281_n10073.n829 4.64734
R53339 a_71281_n10073.n837 a_71281_n10073.n833 4.64734
R53340 a_71281_n10073.n824 a_71281_n10073.n815 4.64734
R53341 a_71281_n10073.n823 a_71281_n10073.n819 4.64734
R53342 a_71281_n10073.n810 a_71281_n10073.n801 4.64734
R53343 a_71281_n10073.n809 a_71281_n10073.n805 4.64734
R53344 a_71281_n10073.n796 a_71281_n10073.n787 4.64734
R53345 a_71281_n10073.n795 a_71281_n10073.n791 4.64734
R53346 a_71281_n10073.n183 a_71281_n10073.n174 4.64734
R53347 a_71281_n10073.n182 a_71281_n10073.n178 4.64734
R53348 a_71281_n10073.n169 a_71281_n10073.n160 4.64734
R53349 a_71281_n10073.n168 a_71281_n10073.n164 4.64734
R53350 a_71281_n10073.n155 a_71281_n10073.n146 4.64734
R53351 a_71281_n10073.n154 a_71281_n10073.n150 4.64734
R53352 a_71281_n10073.n138 a_71281_n10073.n129 4.64734
R53353 a_71281_n10073.n137 a_71281_n10073.n133 4.64734
R53354 a_71281_n10073.n124 a_71281_n10073.n115 4.64734
R53355 a_71281_n10073.n123 a_71281_n10073.n119 4.64734
R53356 a_71281_n10073.n107 a_71281_n10073.n98 4.64734
R53357 a_71281_n10073.n106 a_71281_n10073.n102 4.64734
R53358 a_71281_n10073.n93 a_71281_n10073.n84 4.64734
R53359 a_71281_n10073.n92 a_71281_n10073.n88 4.64734
R53360 a_71281_n10073.n79 a_71281_n10073.n70 4.64734
R53361 a_71281_n10073.n78 a_71281_n10073.n74 4.64734
R53362 a_71281_n10073.n65 a_71281_n10073.n57 4.64734
R53363 a_71281_n10073.n64 a_71281_n10073.n61 4.64734
R53364 a_71281_n10073.n10 a_71281_n10073.n2 4.64734
R53365 a_71281_n10073.n9 a_71281_n10073.n6 4.64734
R53366 a_71281_n10073.n223 a_71281_n10073.n219 4.64734
R53367 a_71281_n10073.n224 a_71281_n10073.n215 4.64734
R53368 a_71281_n10073.n237 a_71281_n10073.n233 4.64734
R53369 a_71281_n10073.n238 a_71281_n10073.n229 4.64734
R53370 a_71281_n10073.n251 a_71281_n10073.n247 4.64734
R53371 a_71281_n10073.n252 a_71281_n10073.n243 4.64734
R53372 a_71281_n10073.n268 a_71281_n10073.n264 4.64734
R53373 a_71281_n10073.n269 a_71281_n10073.n260 4.64734
R53374 a_71281_n10073.n282 a_71281_n10073.n278 4.64734
R53375 a_71281_n10073.n283 a_71281_n10073.n274 4.64734
R53376 a_71281_n10073.n299 a_71281_n10073.n295 4.64734
R53377 a_71281_n10073.n300 a_71281_n10073.n291 4.64734
R53378 a_71281_n10073.n313 a_71281_n10073.n309 4.64734
R53379 a_71281_n10073.n314 a_71281_n10073.n305 4.64734
R53380 a_71281_n10073.n327 a_71281_n10073.n323 4.64734
R53381 a_71281_n10073.n328 a_71281_n10073.n319 4.64734
R53382 a_71281_n10073.n341 a_71281_n10073.n337 4.64734
R53383 a_71281_n10073.n342 a_71281_n10073.n333 4.64734
R53384 a_71281_n10073.n473 a_71281_n10073.n464 4.64734
R53385 a_71281_n10073.n472 a_71281_n10073.n468 4.64734
R53386 a_71281_n10073.n459 a_71281_n10073.n450 4.64734
R53387 a_71281_n10073.n458 a_71281_n10073.n454 4.64734
R53388 a_71281_n10073.n445 a_71281_n10073.n436 4.64734
R53389 a_71281_n10073.n444 a_71281_n10073.n440 4.64734
R53390 a_71281_n10073.n428 a_71281_n10073.n419 4.64734
R53391 a_71281_n10073.n427 a_71281_n10073.n423 4.64734
R53392 a_71281_n10073.n414 a_71281_n10073.n405 4.64734
R53393 a_71281_n10073.n413 a_71281_n10073.n409 4.64734
R53394 a_71281_n10073.n397 a_71281_n10073.n388 4.64734
R53395 a_71281_n10073.n396 a_71281_n10073.n392 4.64734
R53396 a_71281_n10073.n383 a_71281_n10073.n374 4.64734
R53397 a_71281_n10073.n382 a_71281_n10073.n378 4.64734
R53398 a_71281_n10073.n369 a_71281_n10073.n360 4.64734
R53399 a_71281_n10073.n368 a_71281_n10073.n364 4.64734
R53400 a_71281_n10073.n355 a_71281_n10073.n347 4.64734
R53401 a_71281_n10073.n354 a_71281_n10073.n351 4.64734
R53402 a_71281_n10073.n210 a_71281_n10073.n202 4.64734
R53403 a_71281_n10073.n209 a_71281_n10073.n206 4.64734
R53404 a_71281_n10073.n486 a_71281_n10073.n482 4.64734
R53405 a_71281_n10073.n487 a_71281_n10073.n478 4.64734
R53406 a_71281_n10073.n514 a_71281_n10073.n510 4.64734
R53407 a_71281_n10073.n515 a_71281_n10073.n506 4.64734
R53408 a_71281_n10073.n528 a_71281_n10073.n524 4.64734
R53409 a_71281_n10073.n529 a_71281_n10073.n520 4.64734
R53410 a_71281_n10073.n542 a_71281_n10073.n538 4.64734
R53411 a_71281_n10073.n543 a_71281_n10073.n534 4.64734
R53412 a_71281_n10073.n559 a_71281_n10073.n555 4.64734
R53413 a_71281_n10073.n560 a_71281_n10073.n551 4.64734
R53414 a_71281_n10073.n573 a_71281_n10073.n569 4.64734
R53415 a_71281_n10073.n574 a_71281_n10073.n565 4.64734
R53416 a_71281_n10073.n590 a_71281_n10073.n586 4.64734
R53417 a_71281_n10073.n591 a_71281_n10073.n582 4.64734
R53418 a_71281_n10073.n604 a_71281_n10073.n600 4.64734
R53419 a_71281_n10073.n605 a_71281_n10073.n596 4.64734
R53420 a_71281_n10073.n618 a_71281_n10073.n614 4.64734
R53421 a_71281_n10073.n619 a_71281_n10073.n610 4.64734
R53422 a_71281_n10073.n632 a_71281_n10073.n628 4.64734
R53423 a_71281_n10073.n633 a_71281_n10073.n624 4.64734
R53424 a_71281_n10073.n764 a_71281_n10073.n755 4.64734
R53425 a_71281_n10073.n763 a_71281_n10073.n759 4.64734
R53426 a_71281_n10073.n750 a_71281_n10073.n741 4.64734
R53427 a_71281_n10073.n749 a_71281_n10073.n745 4.64734
R53428 a_71281_n10073.n736 a_71281_n10073.n727 4.64734
R53429 a_71281_n10073.n735 a_71281_n10073.n731 4.64734
R53430 a_71281_n10073.n719 a_71281_n10073.n710 4.64734
R53431 a_71281_n10073.n718 a_71281_n10073.n714 4.64734
R53432 a_71281_n10073.n705 a_71281_n10073.n696 4.64734
R53433 a_71281_n10073.n704 a_71281_n10073.n700 4.64734
R53434 a_71281_n10073.n688 a_71281_n10073.n679 4.64734
R53435 a_71281_n10073.n687 a_71281_n10073.n683 4.64734
R53436 a_71281_n10073.n674 a_71281_n10073.n665 4.64734
R53437 a_71281_n10073.n673 a_71281_n10073.n669 4.64734
R53438 a_71281_n10073.n660 a_71281_n10073.n651 4.64734
R53439 a_71281_n10073.n659 a_71281_n10073.n655 4.64734
R53440 a_71281_n10073.n646 a_71281_n10073.n638 4.64734
R53441 a_71281_n10073.n645 a_71281_n10073.n642 4.64734
R53442 a_71281_n10073.n501 a_71281_n10073.n493 4.64734
R53443 a_71281_n10073.n500 a_71281_n10073.n497 4.64734
R53444 a_71281_n10073.n777 a_71281_n10073.n773 4.64734
R53445 a_71281_n10073.n778 a_71281_n10073.n769 4.64734
R53446 a_71281_n10073.n196 a_71281_n10073.n192 4.64734
R53447 a_71281_n10073.n197 a_71281_n10073.n188 4.64734
R53448 a_71281_n10073.n784 a_71281_n10073.n0 18.9036
R53449 a_71281_n10073.n843 a_71281_n10073.n842 4.01884
R53450 a_71281_n10073.n288 a_71281_n10073.n287 4.01884
R53451 a_71281_n10073.n402 a_71281_n10073.n401 4.01884
R53452 a_71281_n10073.n579 a_71281_n10073.n578 4.01884
R53453 a_71281_n10073.n693 a_71281_n10073.n692 4.01884
R53454 a_71281_n10073.n112 a_71281_n10073.n111 4.01884
R53455 a_71281_n10073.n143 a_71281_n10073.n142 4.00982
R53456 a_71281_n10073.n257 a_71281_n10073.n256 4.00982
R53457 a_71281_n10073.n433 a_71281_n10073.n432 4.00982
R53458 a_71281_n10073.n548 a_71281_n10073.n547 4.00982
R53459 a_71281_n10073.n724 a_71281_n10073.n723 4.00982
R53460 a_71281_n10073.n875 a_71281_n10073.n874 4.00982
R53461 a_71281_n10073.n0 a_71281_n10073.t0 3.7215
R53462 a_71281_n10073.n783 a_71281_n10073.n491 3.61592
R53463 a_71281_n10073.n784 a_71281_n10073.n783 2.86491
R53464 a_71281_n10073.n25 a_71281_n10073.n24 2.25278
R53465 a_71281_n10073.n23 a_71281_n10073.n22 2.25278
R53466 a_71281_n10073.n39 a_71281_n10073.n38 2.25278
R53467 a_71281_n10073.n37 a_71281_n10073.n36 2.25278
R53468 a_71281_n10073.n53 a_71281_n10073.n52 2.25278
R53469 a_71281_n10073.n51 a_71281_n10073.n50 2.25278
R53470 a_71281_n10073.n868 a_71281_n10073.n867 2.25278
R53471 a_71281_n10073.n870 a_71281_n10073.n869 2.25278
R53472 a_71281_n10073.n854 a_71281_n10073.n853 2.25278
R53473 a_71281_n10073.n856 a_71281_n10073.n855 2.25278
R53474 a_71281_n10073.n837 a_71281_n10073.n836 2.25278
R53475 a_71281_n10073.n839 a_71281_n10073.n838 2.25278
R53476 a_71281_n10073.n823 a_71281_n10073.n822 2.25278
R53477 a_71281_n10073.n825 a_71281_n10073.n824 2.25278
R53478 a_71281_n10073.n809 a_71281_n10073.n808 2.25278
R53479 a_71281_n10073.n811 a_71281_n10073.n810 2.25278
R53480 a_71281_n10073.n795 a_71281_n10073.n794 2.25278
R53481 a_71281_n10073.n797 a_71281_n10073.n796 2.25278
R53482 a_71281_n10073.n182 a_71281_n10073.n181 2.25278
R53483 a_71281_n10073.n184 a_71281_n10073.n183 2.25278
R53484 a_71281_n10073.n168 a_71281_n10073.n167 2.25278
R53485 a_71281_n10073.n170 a_71281_n10073.n169 2.25278
R53486 a_71281_n10073.n154 a_71281_n10073.n153 2.25278
R53487 a_71281_n10073.n156 a_71281_n10073.n155 2.25278
R53488 a_71281_n10073.n137 a_71281_n10073.n136 2.25278
R53489 a_71281_n10073.n139 a_71281_n10073.n138 2.25278
R53490 a_71281_n10073.n123 a_71281_n10073.n122 2.25278
R53491 a_71281_n10073.n125 a_71281_n10073.n124 2.25278
R53492 a_71281_n10073.n106 a_71281_n10073.n105 2.25278
R53493 a_71281_n10073.n108 a_71281_n10073.n107 2.25278
R53494 a_71281_n10073.n92 a_71281_n10073.n91 2.25278
R53495 a_71281_n10073.n94 a_71281_n10073.n93 2.25278
R53496 a_71281_n10073.n78 a_71281_n10073.n77 2.25278
R53497 a_71281_n10073.n80 a_71281_n10073.n79 2.25278
R53498 a_71281_n10073.n64 a_71281_n10073.n63 2.25278
R53499 a_71281_n10073.n66 a_71281_n10073.n65 2.25278
R53500 a_71281_n10073.n9 a_71281_n10073.n8 2.25278
R53501 a_71281_n10073.n11 a_71281_n10073.n10 2.25278
R53502 a_71281_n10073.n225 a_71281_n10073.n224 2.25278
R53503 a_71281_n10073.n223 a_71281_n10073.n222 2.25278
R53504 a_71281_n10073.n239 a_71281_n10073.n238 2.25278
R53505 a_71281_n10073.n237 a_71281_n10073.n236 2.25278
R53506 a_71281_n10073.n253 a_71281_n10073.n252 2.25278
R53507 a_71281_n10073.n251 a_71281_n10073.n250 2.25278
R53508 a_71281_n10073.n270 a_71281_n10073.n269 2.25278
R53509 a_71281_n10073.n268 a_71281_n10073.n267 2.25278
R53510 a_71281_n10073.n284 a_71281_n10073.n283 2.25278
R53511 a_71281_n10073.n282 a_71281_n10073.n281 2.25278
R53512 a_71281_n10073.n301 a_71281_n10073.n300 2.25278
R53513 a_71281_n10073.n299 a_71281_n10073.n298 2.25278
R53514 a_71281_n10073.n315 a_71281_n10073.n314 2.25278
R53515 a_71281_n10073.n313 a_71281_n10073.n312 2.25278
R53516 a_71281_n10073.n329 a_71281_n10073.n328 2.25278
R53517 a_71281_n10073.n327 a_71281_n10073.n326 2.25278
R53518 a_71281_n10073.n343 a_71281_n10073.n342 2.25278
R53519 a_71281_n10073.n341 a_71281_n10073.n340 2.25278
R53520 a_71281_n10073.n472 a_71281_n10073.n471 2.25278
R53521 a_71281_n10073.n474 a_71281_n10073.n473 2.25278
R53522 a_71281_n10073.n458 a_71281_n10073.n457 2.25278
R53523 a_71281_n10073.n460 a_71281_n10073.n459 2.25278
R53524 a_71281_n10073.n444 a_71281_n10073.n443 2.25278
R53525 a_71281_n10073.n446 a_71281_n10073.n445 2.25278
R53526 a_71281_n10073.n427 a_71281_n10073.n426 2.25278
R53527 a_71281_n10073.n429 a_71281_n10073.n428 2.25278
R53528 a_71281_n10073.n413 a_71281_n10073.n412 2.25278
R53529 a_71281_n10073.n415 a_71281_n10073.n414 2.25278
R53530 a_71281_n10073.n396 a_71281_n10073.n395 2.25278
R53531 a_71281_n10073.n398 a_71281_n10073.n397 2.25278
R53532 a_71281_n10073.n382 a_71281_n10073.n381 2.25278
R53533 a_71281_n10073.n384 a_71281_n10073.n383 2.25278
R53534 a_71281_n10073.n368 a_71281_n10073.n367 2.25278
R53535 a_71281_n10073.n370 a_71281_n10073.n369 2.25278
R53536 a_71281_n10073.n354 a_71281_n10073.n353 2.25278
R53537 a_71281_n10073.n356 a_71281_n10073.n355 2.25278
R53538 a_71281_n10073.n209 a_71281_n10073.n208 2.25278
R53539 a_71281_n10073.n211 a_71281_n10073.n210 2.25278
R53540 a_71281_n10073.n488 a_71281_n10073.n487 2.25278
R53541 a_71281_n10073.n486 a_71281_n10073.n485 2.25278
R53542 a_71281_n10073.n516 a_71281_n10073.n515 2.25278
R53543 a_71281_n10073.n514 a_71281_n10073.n513 2.25278
R53544 a_71281_n10073.n530 a_71281_n10073.n529 2.25278
R53545 a_71281_n10073.n528 a_71281_n10073.n527 2.25278
R53546 a_71281_n10073.n544 a_71281_n10073.n543 2.25278
R53547 a_71281_n10073.n542 a_71281_n10073.n541 2.25278
R53548 a_71281_n10073.n561 a_71281_n10073.n560 2.25278
R53549 a_71281_n10073.n559 a_71281_n10073.n558 2.25278
R53550 a_71281_n10073.n575 a_71281_n10073.n574 2.25278
R53551 a_71281_n10073.n573 a_71281_n10073.n572 2.25278
R53552 a_71281_n10073.n592 a_71281_n10073.n591 2.25278
R53553 a_71281_n10073.n590 a_71281_n10073.n589 2.25278
R53554 a_71281_n10073.n606 a_71281_n10073.n605 2.25278
R53555 a_71281_n10073.n604 a_71281_n10073.n603 2.25278
R53556 a_71281_n10073.n620 a_71281_n10073.n619 2.25278
R53557 a_71281_n10073.n618 a_71281_n10073.n617 2.25278
R53558 a_71281_n10073.n634 a_71281_n10073.n633 2.25278
R53559 a_71281_n10073.n632 a_71281_n10073.n631 2.25278
R53560 a_71281_n10073.n763 a_71281_n10073.n762 2.25278
R53561 a_71281_n10073.n765 a_71281_n10073.n764 2.25278
R53562 a_71281_n10073.n749 a_71281_n10073.n748 2.25278
R53563 a_71281_n10073.n751 a_71281_n10073.n750 2.25278
R53564 a_71281_n10073.n735 a_71281_n10073.n734 2.25278
R53565 a_71281_n10073.n737 a_71281_n10073.n736 2.25278
R53566 a_71281_n10073.n718 a_71281_n10073.n717 2.25278
R53567 a_71281_n10073.n720 a_71281_n10073.n719 2.25278
R53568 a_71281_n10073.n704 a_71281_n10073.n703 2.25278
R53569 a_71281_n10073.n706 a_71281_n10073.n705 2.25278
R53570 a_71281_n10073.n687 a_71281_n10073.n686 2.25278
R53571 a_71281_n10073.n689 a_71281_n10073.n688 2.25278
R53572 a_71281_n10073.n673 a_71281_n10073.n672 2.25278
R53573 a_71281_n10073.n675 a_71281_n10073.n674 2.25278
R53574 a_71281_n10073.n659 a_71281_n10073.n658 2.25278
R53575 a_71281_n10073.n661 a_71281_n10073.n660 2.25278
R53576 a_71281_n10073.n645 a_71281_n10073.n644 2.25278
R53577 a_71281_n10073.n647 a_71281_n10073.n646 2.25278
R53578 a_71281_n10073.n500 a_71281_n10073.n499 2.25278
R53579 a_71281_n10073.n502 a_71281_n10073.n501 2.25278
R53580 a_71281_n10073.n779 a_71281_n10073.n778 2.25278
R53581 a_71281_n10073.n777 a_71281_n10073.n776 2.25278
R53582 a_71281_n10073.n198 a_71281_n10073.n197 2.25278
R53583 a_71281_n10073.n196 a_71281_n10073.n195 2.25278
R53584 a_71281_n10073.n213 a_71281_n10073.n201 1.6802
R53585 a_71281_n10073.n358 a_71281_n10073.n346 1.6802
R53586 a_71281_n10073.n504 a_71281_n10073.n492 1.6802
R53587 a_71281_n10073.n649 a_71281_n10073.n637 1.6802
R53588 a_71281_n10073.n13 a_71281_n10073.n1 1.6802
R53589 a_71281_n10073.n68 a_71281_n10073.n56 1.6802
R53590 a_71281_n10073.n403 a_71281_n10073.n402 1.5005
R53591 a_71281_n10073.n483 a_71281_n10073.n477 1.5005
R53592 a_71281_n10073.n289 a_71281_n10073.n288 1.5005
R53593 a_71281_n10073.n213 a_71281_n10073.n212 1.5005
R53594 a_71281_n10073.n434 a_71281_n10073.n433 1.5005
R53595 a_71281_n10073.n258 a_71281_n10073.n257 1.5005
R53596 a_71281_n10073.n358 a_71281_n10073.n357 1.5005
R53597 a_71281_n10073.n372 a_71281_n10073.n371 1.5005
R53598 a_71281_n10073.n366 a_71281_n10073.n359 1.5005
R53599 a_71281_n10073.n386 a_71281_n10073.n385 1.5005
R53600 a_71281_n10073.n380 a_71281_n10073.n373 1.5005
R53601 a_71281_n10073.n400 a_71281_n10073.n399 1.5005
R53602 a_71281_n10073.n394 a_71281_n10073.n387 1.5005
R53603 a_71281_n10073.n417 a_71281_n10073.n416 1.5005
R53604 a_71281_n10073.n411 a_71281_n10073.n404 1.5005
R53605 a_71281_n10073.n431 a_71281_n10073.n430 1.5005
R53606 a_71281_n10073.n425 a_71281_n10073.n418 1.5005
R53607 a_71281_n10073.n448 a_71281_n10073.n447 1.5005
R53608 a_71281_n10073.n442 a_71281_n10073.n435 1.5005
R53609 a_71281_n10073.n462 a_71281_n10073.n461 1.5005
R53610 a_71281_n10073.n456 a_71281_n10073.n449 1.5005
R53611 a_71281_n10073.n476 a_71281_n10073.n475 1.5005
R53612 a_71281_n10073.n470 a_71281_n10073.n463 1.5005
R53613 a_71281_n10073.n490 a_71281_n10073.n489 1.5005
R53614 a_71281_n10073.n338 a_71281_n10073.n332 1.5005
R53615 a_71281_n10073.n345 a_71281_n10073.n344 1.5005
R53616 a_71281_n10073.n324 a_71281_n10073.n318 1.5005
R53617 a_71281_n10073.n331 a_71281_n10073.n330 1.5005
R53618 a_71281_n10073.n310 a_71281_n10073.n304 1.5005
R53619 a_71281_n10073.n317 a_71281_n10073.n316 1.5005
R53620 a_71281_n10073.n296 a_71281_n10073.n290 1.5005
R53621 a_71281_n10073.n303 a_71281_n10073.n302 1.5005
R53622 a_71281_n10073.n279 a_71281_n10073.n273 1.5005
R53623 a_71281_n10073.n286 a_71281_n10073.n285 1.5005
R53624 a_71281_n10073.n265 a_71281_n10073.n259 1.5005
R53625 a_71281_n10073.n272 a_71281_n10073.n271 1.5005
R53626 a_71281_n10073.n248 a_71281_n10073.n242 1.5005
R53627 a_71281_n10073.n255 a_71281_n10073.n254 1.5005
R53628 a_71281_n10073.n234 a_71281_n10073.n228 1.5005
R53629 a_71281_n10073.n241 a_71281_n10073.n240 1.5005
R53630 a_71281_n10073.n220 a_71281_n10073.n214 1.5005
R53631 a_71281_n10073.n227 a_71281_n10073.n226 1.5005
R53632 a_71281_n10073.n694 a_71281_n10073.n693 1.5005
R53633 a_71281_n10073.n774 a_71281_n10073.n768 1.5005
R53634 a_71281_n10073.n580 a_71281_n10073.n579 1.5005
R53635 a_71281_n10073.n504 a_71281_n10073.n503 1.5005
R53636 a_71281_n10073.n725 a_71281_n10073.n724 1.5005
R53637 a_71281_n10073.n549 a_71281_n10073.n548 1.5005
R53638 a_71281_n10073.n649 a_71281_n10073.n648 1.5005
R53639 a_71281_n10073.n663 a_71281_n10073.n662 1.5005
R53640 a_71281_n10073.n657 a_71281_n10073.n650 1.5005
R53641 a_71281_n10073.n677 a_71281_n10073.n676 1.5005
R53642 a_71281_n10073.n671 a_71281_n10073.n664 1.5005
R53643 a_71281_n10073.n691 a_71281_n10073.n690 1.5005
R53644 a_71281_n10073.n685 a_71281_n10073.n678 1.5005
R53645 a_71281_n10073.n708 a_71281_n10073.n707 1.5005
R53646 a_71281_n10073.n702 a_71281_n10073.n695 1.5005
R53647 a_71281_n10073.n722 a_71281_n10073.n721 1.5005
R53648 a_71281_n10073.n716 a_71281_n10073.n709 1.5005
R53649 a_71281_n10073.n739 a_71281_n10073.n738 1.5005
R53650 a_71281_n10073.n733 a_71281_n10073.n726 1.5005
R53651 a_71281_n10073.n753 a_71281_n10073.n752 1.5005
R53652 a_71281_n10073.n747 a_71281_n10073.n740 1.5005
R53653 a_71281_n10073.n767 a_71281_n10073.n766 1.5005
R53654 a_71281_n10073.n761 a_71281_n10073.n754 1.5005
R53655 a_71281_n10073.n781 a_71281_n10073.n780 1.5005
R53656 a_71281_n10073.n629 a_71281_n10073.n623 1.5005
R53657 a_71281_n10073.n636 a_71281_n10073.n635 1.5005
R53658 a_71281_n10073.n615 a_71281_n10073.n609 1.5005
R53659 a_71281_n10073.n622 a_71281_n10073.n621 1.5005
R53660 a_71281_n10073.n601 a_71281_n10073.n595 1.5005
R53661 a_71281_n10073.n608 a_71281_n10073.n607 1.5005
R53662 a_71281_n10073.n587 a_71281_n10073.n581 1.5005
R53663 a_71281_n10073.n594 a_71281_n10073.n593 1.5005
R53664 a_71281_n10073.n570 a_71281_n10073.n564 1.5005
R53665 a_71281_n10073.n577 a_71281_n10073.n576 1.5005
R53666 a_71281_n10073.n556 a_71281_n10073.n550 1.5005
R53667 a_71281_n10073.n563 a_71281_n10073.n562 1.5005
R53668 a_71281_n10073.n539 a_71281_n10073.n533 1.5005
R53669 a_71281_n10073.n546 a_71281_n10073.n545 1.5005
R53670 a_71281_n10073.n525 a_71281_n10073.n519 1.5005
R53671 a_71281_n10073.n532 a_71281_n10073.n531 1.5005
R53672 a_71281_n10073.n511 a_71281_n10073.n505 1.5005
R53673 a_71281_n10073.n518 a_71281_n10073.n517 1.5005
R53674 a_71281_n10073.n113 a_71281_n10073.n112 1.5005
R53675 a_71281_n10073.n193 a_71281_n10073.n187 1.5005
R53676 a_71281_n10073.n844 a_71281_n10073.n843 1.5005
R53677 a_71281_n10073.n13 a_71281_n10073.n12 1.5005
R53678 a_71281_n10073.n144 a_71281_n10073.n143 1.5005
R53679 a_71281_n10073.n68 a_71281_n10073.n67 1.5005
R53680 a_71281_n10073.n82 a_71281_n10073.n81 1.5005
R53681 a_71281_n10073.n76 a_71281_n10073.n69 1.5005
R53682 a_71281_n10073.n96 a_71281_n10073.n95 1.5005
R53683 a_71281_n10073.n90 a_71281_n10073.n83 1.5005
R53684 a_71281_n10073.n110 a_71281_n10073.n109 1.5005
R53685 a_71281_n10073.n104 a_71281_n10073.n97 1.5005
R53686 a_71281_n10073.n127 a_71281_n10073.n126 1.5005
R53687 a_71281_n10073.n121 a_71281_n10073.n114 1.5005
R53688 a_71281_n10073.n141 a_71281_n10073.n140 1.5005
R53689 a_71281_n10073.n135 a_71281_n10073.n128 1.5005
R53690 a_71281_n10073.n158 a_71281_n10073.n157 1.5005
R53691 a_71281_n10073.n152 a_71281_n10073.n145 1.5005
R53692 a_71281_n10073.n172 a_71281_n10073.n171 1.5005
R53693 a_71281_n10073.n166 a_71281_n10073.n159 1.5005
R53694 a_71281_n10073.n186 a_71281_n10073.n185 1.5005
R53695 a_71281_n10073.n180 a_71281_n10073.n173 1.5005
R53696 a_71281_n10073.n200 a_71281_n10073.n199 1.5005
R53697 a_71281_n10073.n799 a_71281_n10073.n798 1.5005
R53698 a_71281_n10073.n793 a_71281_n10073.n786 1.5005
R53699 a_71281_n10073.n813 a_71281_n10073.n812 1.5005
R53700 a_71281_n10073.n807 a_71281_n10073.n800 1.5005
R53701 a_71281_n10073.n827 a_71281_n10073.n826 1.5005
R53702 a_71281_n10073.n821 a_71281_n10073.n814 1.5005
R53703 a_71281_n10073.n841 a_71281_n10073.n840 1.5005
R53704 a_71281_n10073.n835 a_71281_n10073.n828 1.5005
R53705 a_71281_n10073.n858 a_71281_n10073.n857 1.5005
R53706 a_71281_n10073.n852 a_71281_n10073.n845 1.5005
R53707 a_71281_n10073.n872 a_71281_n10073.n871 1.5005
R53708 a_71281_n10073.n866 a_71281_n10073.n859 1.5005
R53709 a_71281_n10073.n48 a_71281_n10073.n42 1.5005
R53710 a_71281_n10073.n55 a_71281_n10073.n54 1.5005
R53711 a_71281_n10073.n34 a_71281_n10073.n28 1.5005
R53712 a_71281_n10073.n41 a_71281_n10073.n40 1.5005
R53713 a_71281_n10073.n20 a_71281_n10073.n14 1.5005
R53714 a_71281_n10073.n27 a_71281_n10073.n26 1.5005
R53715 a_71281_n10073.n874 a_71281_n10073.n873 1.5005
R53716 a_71281_n10073.n142 a_71281_n10073.t31 1.4705
R53717 a_71281_n10073.n142 a_71281_n10073.t9 1.4705
R53718 a_71281_n10073.n842 a_71281_n10073.t41 1.4705
R53719 a_71281_n10073.n842 a_71281_n10073.t17 1.4705
R53720 a_71281_n10073.n256 a_71281_n10073.t69 1.4705
R53721 a_71281_n10073.n256 a_71281_n10073.t53 1.4705
R53722 a_71281_n10073.n432 a_71281_n10073.t57 1.4705
R53723 a_71281_n10073.n432 a_71281_n10073.t21 1.4705
R53724 a_71281_n10073.n287 a_71281_n10073.t25 1.4705
R53725 a_71281_n10073.n287 a_71281_n10073.t3 1.4705
R53726 a_71281_n10073.n401 a_71281_n10073.t5 1.4705
R53727 a_71281_n10073.n401 a_71281_n10073.t7 1.4705
R53728 a_71281_n10073.n547 a_71281_n10073.t13 1.4705
R53729 a_71281_n10073.n547 a_71281_n10073.t65 1.4705
R53730 a_71281_n10073.n723 a_71281_n10073.t51 1.4705
R53731 a_71281_n10073.n723 a_71281_n10073.t55 1.4705
R53732 a_71281_n10073.n578 a_71281_n10073.t43 1.4705
R53733 a_71281_n10073.n578 a_71281_n10073.t37 1.4705
R53734 a_71281_n10073.n692 a_71281_n10073.t33 1.4705
R53735 a_71281_n10073.n692 a_71281_n10073.t11 1.4705
R53736 a_71281_n10073.n111 a_71281_n10073.t67 1.4705
R53737 a_71281_n10073.n111 a_71281_n10073.t39 1.4705
R53738 a_71281_n10073.t73 a_71281_n10073.n875 1.4705
R53739 a_71281_n10073.n875 a_71281_n10073.t63 1.4705
R53740 a_71281_n10073.n783 a_71281_n10073.n782 0.7505
R53741 a_71281_n10073.n785 a_71281_n10073.n784 0.7505
R53742 a_71281_n10073.n25 a_71281_n10073.n16 0.567403
R53743 a_71281_n10073.n22 a_71281_n10073.n21 0.567403
R53744 a_71281_n10073.n39 a_71281_n10073.n30 0.567403
R53745 a_71281_n10073.n36 a_71281_n10073.n35 0.567403
R53746 a_71281_n10073.n53 a_71281_n10073.n44 0.567403
R53747 a_71281_n10073.n50 a_71281_n10073.n49 0.567403
R53748 a_71281_n10073.n867 a_71281_n10073.n865 0.567403
R53749 a_71281_n10073.n870 a_71281_n10073.n861 0.567403
R53750 a_71281_n10073.n853 a_71281_n10073.n851 0.567403
R53751 a_71281_n10073.n856 a_71281_n10073.n847 0.567403
R53752 a_71281_n10073.n836 a_71281_n10073.n834 0.567403
R53753 a_71281_n10073.n839 a_71281_n10073.n830 0.567403
R53754 a_71281_n10073.n822 a_71281_n10073.n820 0.567403
R53755 a_71281_n10073.n825 a_71281_n10073.n816 0.567403
R53756 a_71281_n10073.n808 a_71281_n10073.n806 0.567403
R53757 a_71281_n10073.n811 a_71281_n10073.n802 0.567403
R53758 a_71281_n10073.n794 a_71281_n10073.n792 0.567403
R53759 a_71281_n10073.n797 a_71281_n10073.n788 0.567403
R53760 a_71281_n10073.n181 a_71281_n10073.n179 0.567403
R53761 a_71281_n10073.n184 a_71281_n10073.n175 0.567403
R53762 a_71281_n10073.n167 a_71281_n10073.n165 0.567403
R53763 a_71281_n10073.n170 a_71281_n10073.n161 0.567403
R53764 a_71281_n10073.n153 a_71281_n10073.n151 0.567403
R53765 a_71281_n10073.n156 a_71281_n10073.n147 0.567403
R53766 a_71281_n10073.n136 a_71281_n10073.n134 0.567403
R53767 a_71281_n10073.n139 a_71281_n10073.n130 0.567403
R53768 a_71281_n10073.n122 a_71281_n10073.n120 0.567403
R53769 a_71281_n10073.n125 a_71281_n10073.n116 0.567403
R53770 a_71281_n10073.n105 a_71281_n10073.n103 0.567403
R53771 a_71281_n10073.n108 a_71281_n10073.n99 0.567403
R53772 a_71281_n10073.n91 a_71281_n10073.n89 0.567403
R53773 a_71281_n10073.n94 a_71281_n10073.n85 0.567403
R53774 a_71281_n10073.n77 a_71281_n10073.n75 0.567403
R53775 a_71281_n10073.n80 a_71281_n10073.n71 0.567403
R53776 a_71281_n10073.n63 a_71281_n10073.n62 0.567403
R53777 a_71281_n10073.n66 a_71281_n10073.n58 0.567403
R53778 a_71281_n10073.n8 a_71281_n10073.n7 0.567403
R53779 a_71281_n10073.n11 a_71281_n10073.n3 0.567403
R53780 a_71281_n10073.n225 a_71281_n10073.n216 0.567403
R53781 a_71281_n10073.n222 a_71281_n10073.n221 0.567403
R53782 a_71281_n10073.n239 a_71281_n10073.n230 0.567403
R53783 a_71281_n10073.n236 a_71281_n10073.n235 0.567403
R53784 a_71281_n10073.n253 a_71281_n10073.n244 0.567403
R53785 a_71281_n10073.n250 a_71281_n10073.n249 0.567403
R53786 a_71281_n10073.n270 a_71281_n10073.n261 0.567403
R53787 a_71281_n10073.n267 a_71281_n10073.n266 0.567403
R53788 a_71281_n10073.n284 a_71281_n10073.n275 0.567403
R53789 a_71281_n10073.n281 a_71281_n10073.n280 0.567403
R53790 a_71281_n10073.n301 a_71281_n10073.n292 0.567403
R53791 a_71281_n10073.n298 a_71281_n10073.n297 0.567403
R53792 a_71281_n10073.n315 a_71281_n10073.n306 0.567403
R53793 a_71281_n10073.n312 a_71281_n10073.n311 0.567403
R53794 a_71281_n10073.n329 a_71281_n10073.n320 0.567403
R53795 a_71281_n10073.n326 a_71281_n10073.n325 0.567403
R53796 a_71281_n10073.n343 a_71281_n10073.n334 0.567403
R53797 a_71281_n10073.n340 a_71281_n10073.n339 0.567403
R53798 a_71281_n10073.n471 a_71281_n10073.n469 0.567403
R53799 a_71281_n10073.n474 a_71281_n10073.n465 0.567403
R53800 a_71281_n10073.n457 a_71281_n10073.n455 0.567403
R53801 a_71281_n10073.n460 a_71281_n10073.n451 0.567403
R53802 a_71281_n10073.n443 a_71281_n10073.n441 0.567403
R53803 a_71281_n10073.n446 a_71281_n10073.n437 0.567403
R53804 a_71281_n10073.n426 a_71281_n10073.n424 0.567403
R53805 a_71281_n10073.n429 a_71281_n10073.n420 0.567403
R53806 a_71281_n10073.n412 a_71281_n10073.n410 0.567403
R53807 a_71281_n10073.n415 a_71281_n10073.n406 0.567403
R53808 a_71281_n10073.n395 a_71281_n10073.n393 0.567403
R53809 a_71281_n10073.n398 a_71281_n10073.n389 0.567403
R53810 a_71281_n10073.n381 a_71281_n10073.n379 0.567403
R53811 a_71281_n10073.n384 a_71281_n10073.n375 0.567403
R53812 a_71281_n10073.n367 a_71281_n10073.n365 0.567403
R53813 a_71281_n10073.n370 a_71281_n10073.n361 0.567403
R53814 a_71281_n10073.n353 a_71281_n10073.n352 0.567403
R53815 a_71281_n10073.n356 a_71281_n10073.n348 0.567403
R53816 a_71281_n10073.n208 a_71281_n10073.n207 0.567403
R53817 a_71281_n10073.n211 a_71281_n10073.n203 0.567403
R53818 a_71281_n10073.n488 a_71281_n10073.n479 0.567403
R53819 a_71281_n10073.n485 a_71281_n10073.n484 0.567403
R53820 a_71281_n10073.n516 a_71281_n10073.n507 0.567403
R53821 a_71281_n10073.n513 a_71281_n10073.n512 0.567403
R53822 a_71281_n10073.n530 a_71281_n10073.n521 0.567403
R53823 a_71281_n10073.n527 a_71281_n10073.n526 0.567403
R53824 a_71281_n10073.n544 a_71281_n10073.n535 0.567403
R53825 a_71281_n10073.n541 a_71281_n10073.n540 0.567403
R53826 a_71281_n10073.n561 a_71281_n10073.n552 0.567403
R53827 a_71281_n10073.n558 a_71281_n10073.n557 0.567403
R53828 a_71281_n10073.n575 a_71281_n10073.n566 0.567403
R53829 a_71281_n10073.n572 a_71281_n10073.n571 0.567403
R53830 a_71281_n10073.n592 a_71281_n10073.n583 0.567403
R53831 a_71281_n10073.n589 a_71281_n10073.n588 0.567403
R53832 a_71281_n10073.n606 a_71281_n10073.n597 0.567403
R53833 a_71281_n10073.n603 a_71281_n10073.n602 0.567403
R53834 a_71281_n10073.n620 a_71281_n10073.n611 0.567403
R53835 a_71281_n10073.n617 a_71281_n10073.n616 0.567403
R53836 a_71281_n10073.n634 a_71281_n10073.n625 0.567403
R53837 a_71281_n10073.n631 a_71281_n10073.n630 0.567403
R53838 a_71281_n10073.n762 a_71281_n10073.n760 0.567403
R53839 a_71281_n10073.n765 a_71281_n10073.n756 0.567403
R53840 a_71281_n10073.n748 a_71281_n10073.n746 0.567403
R53841 a_71281_n10073.n751 a_71281_n10073.n742 0.567403
R53842 a_71281_n10073.n734 a_71281_n10073.n732 0.567403
R53843 a_71281_n10073.n737 a_71281_n10073.n728 0.567403
R53844 a_71281_n10073.n717 a_71281_n10073.n715 0.567403
R53845 a_71281_n10073.n720 a_71281_n10073.n711 0.567403
R53846 a_71281_n10073.n703 a_71281_n10073.n701 0.567403
R53847 a_71281_n10073.n706 a_71281_n10073.n697 0.567403
R53848 a_71281_n10073.n686 a_71281_n10073.n684 0.567403
R53849 a_71281_n10073.n689 a_71281_n10073.n680 0.567403
R53850 a_71281_n10073.n672 a_71281_n10073.n670 0.567403
R53851 a_71281_n10073.n675 a_71281_n10073.n666 0.567403
R53852 a_71281_n10073.n658 a_71281_n10073.n656 0.567403
R53853 a_71281_n10073.n661 a_71281_n10073.n652 0.567403
R53854 a_71281_n10073.n644 a_71281_n10073.n643 0.567403
R53855 a_71281_n10073.n647 a_71281_n10073.n639 0.567403
R53856 a_71281_n10073.n499 a_71281_n10073.n498 0.567403
R53857 a_71281_n10073.n502 a_71281_n10073.n494 0.567403
R53858 a_71281_n10073.n779 a_71281_n10073.n770 0.567403
R53859 a_71281_n10073.n776 a_71281_n10073.n775 0.567403
R53860 a_71281_n10073.n198 a_71281_n10073.n189 0.567403
R53861 a_71281_n10073.n195 a_71281_n10073.n194 0.567403
R53862 a_71281_n10073.n17 a_71281_n10073.n15 0.496742
R53863 a_71281_n10073.n19 a_71281_n10073.n18 0.496742
R53864 a_71281_n10073.n31 a_71281_n10073.n29 0.496742
R53865 a_71281_n10073.n33 a_71281_n10073.n32 0.496742
R53866 a_71281_n10073.n45 a_71281_n10073.n43 0.496742
R53867 a_71281_n10073.n47 a_71281_n10073.n46 0.496742
R53868 a_71281_n10073.n864 a_71281_n10073.n863 0.496742
R53869 a_71281_n10073.n862 a_71281_n10073.n860 0.496742
R53870 a_71281_n10073.n850 a_71281_n10073.n849 0.496742
R53871 a_71281_n10073.n848 a_71281_n10073.n846 0.496742
R53872 a_71281_n10073.n833 a_71281_n10073.n832 0.496742
R53873 a_71281_n10073.n831 a_71281_n10073.n829 0.496742
R53874 a_71281_n10073.n819 a_71281_n10073.n818 0.496742
R53875 a_71281_n10073.n817 a_71281_n10073.n815 0.496742
R53876 a_71281_n10073.n805 a_71281_n10073.n804 0.496742
R53877 a_71281_n10073.n803 a_71281_n10073.n801 0.496742
R53878 a_71281_n10073.n791 a_71281_n10073.n790 0.496742
R53879 a_71281_n10073.n789 a_71281_n10073.n787 0.496742
R53880 a_71281_n10073.n178 a_71281_n10073.n177 0.496742
R53881 a_71281_n10073.n176 a_71281_n10073.n174 0.496742
R53882 a_71281_n10073.n164 a_71281_n10073.n163 0.496742
R53883 a_71281_n10073.n162 a_71281_n10073.n160 0.496742
R53884 a_71281_n10073.n150 a_71281_n10073.n149 0.496742
R53885 a_71281_n10073.n148 a_71281_n10073.n146 0.496742
R53886 a_71281_n10073.n133 a_71281_n10073.n132 0.496742
R53887 a_71281_n10073.n131 a_71281_n10073.n129 0.496742
R53888 a_71281_n10073.n119 a_71281_n10073.n118 0.496742
R53889 a_71281_n10073.n117 a_71281_n10073.n115 0.496742
R53890 a_71281_n10073.n102 a_71281_n10073.n101 0.496742
R53891 a_71281_n10073.n100 a_71281_n10073.n98 0.496742
R53892 a_71281_n10073.n88 a_71281_n10073.n87 0.496742
R53893 a_71281_n10073.n86 a_71281_n10073.n84 0.496742
R53894 a_71281_n10073.n74 a_71281_n10073.n73 0.496742
R53895 a_71281_n10073.n72 a_71281_n10073.n70 0.496742
R53896 a_71281_n10073.n61 a_71281_n10073.n60 0.496742
R53897 a_71281_n10073.n59 a_71281_n10073.n57 0.496742
R53898 a_71281_n10073.n6 a_71281_n10073.n5 0.496742
R53899 a_71281_n10073.n4 a_71281_n10073.n2 0.496742
R53900 a_71281_n10073.n217 a_71281_n10073.n215 0.496742
R53901 a_71281_n10073.n219 a_71281_n10073.n218 0.496742
R53902 a_71281_n10073.n231 a_71281_n10073.n229 0.496742
R53903 a_71281_n10073.n233 a_71281_n10073.n232 0.496742
R53904 a_71281_n10073.n245 a_71281_n10073.n243 0.496742
R53905 a_71281_n10073.n247 a_71281_n10073.n246 0.496742
R53906 a_71281_n10073.n262 a_71281_n10073.n260 0.496742
R53907 a_71281_n10073.n264 a_71281_n10073.n263 0.496742
R53908 a_71281_n10073.n276 a_71281_n10073.n274 0.496742
R53909 a_71281_n10073.n278 a_71281_n10073.n277 0.496742
R53910 a_71281_n10073.n293 a_71281_n10073.n291 0.496742
R53911 a_71281_n10073.n295 a_71281_n10073.n294 0.496742
R53912 a_71281_n10073.n307 a_71281_n10073.n305 0.496742
R53913 a_71281_n10073.n309 a_71281_n10073.n308 0.496742
R53914 a_71281_n10073.n321 a_71281_n10073.n319 0.496742
R53915 a_71281_n10073.n323 a_71281_n10073.n322 0.496742
R53916 a_71281_n10073.n335 a_71281_n10073.n333 0.496742
R53917 a_71281_n10073.n337 a_71281_n10073.n336 0.496742
R53918 a_71281_n10073.n468 a_71281_n10073.n467 0.496742
R53919 a_71281_n10073.n466 a_71281_n10073.n464 0.496742
R53920 a_71281_n10073.n454 a_71281_n10073.n453 0.496742
R53921 a_71281_n10073.n452 a_71281_n10073.n450 0.496742
R53922 a_71281_n10073.n440 a_71281_n10073.n439 0.496742
R53923 a_71281_n10073.n438 a_71281_n10073.n436 0.496742
R53924 a_71281_n10073.n423 a_71281_n10073.n422 0.496742
R53925 a_71281_n10073.n421 a_71281_n10073.n419 0.496742
R53926 a_71281_n10073.n409 a_71281_n10073.n408 0.496742
R53927 a_71281_n10073.n407 a_71281_n10073.n405 0.496742
R53928 a_71281_n10073.n392 a_71281_n10073.n391 0.496742
R53929 a_71281_n10073.n390 a_71281_n10073.n388 0.496742
R53930 a_71281_n10073.n378 a_71281_n10073.n377 0.496742
R53931 a_71281_n10073.n376 a_71281_n10073.n374 0.496742
R53932 a_71281_n10073.n364 a_71281_n10073.n363 0.496742
R53933 a_71281_n10073.n362 a_71281_n10073.n360 0.496742
R53934 a_71281_n10073.n351 a_71281_n10073.n350 0.496742
R53935 a_71281_n10073.n349 a_71281_n10073.n347 0.496742
R53936 a_71281_n10073.n206 a_71281_n10073.n205 0.496742
R53937 a_71281_n10073.n204 a_71281_n10073.n202 0.496742
R53938 a_71281_n10073.n480 a_71281_n10073.n478 0.496742
R53939 a_71281_n10073.n482 a_71281_n10073.n481 0.496742
R53940 a_71281_n10073.n508 a_71281_n10073.n506 0.496742
R53941 a_71281_n10073.n510 a_71281_n10073.n509 0.496742
R53942 a_71281_n10073.n522 a_71281_n10073.n520 0.496742
R53943 a_71281_n10073.n524 a_71281_n10073.n523 0.496742
R53944 a_71281_n10073.n536 a_71281_n10073.n534 0.496742
R53945 a_71281_n10073.n538 a_71281_n10073.n537 0.496742
R53946 a_71281_n10073.n553 a_71281_n10073.n551 0.496742
R53947 a_71281_n10073.n555 a_71281_n10073.n554 0.496742
R53948 a_71281_n10073.n567 a_71281_n10073.n565 0.496742
R53949 a_71281_n10073.n569 a_71281_n10073.n568 0.496742
R53950 a_71281_n10073.n584 a_71281_n10073.n582 0.496742
R53951 a_71281_n10073.n586 a_71281_n10073.n585 0.496742
R53952 a_71281_n10073.n598 a_71281_n10073.n596 0.496742
R53953 a_71281_n10073.n600 a_71281_n10073.n599 0.496742
R53954 a_71281_n10073.n612 a_71281_n10073.n610 0.496742
R53955 a_71281_n10073.n614 a_71281_n10073.n613 0.496742
R53956 a_71281_n10073.n626 a_71281_n10073.n624 0.496742
R53957 a_71281_n10073.n628 a_71281_n10073.n627 0.496742
R53958 a_71281_n10073.n759 a_71281_n10073.n758 0.496742
R53959 a_71281_n10073.n757 a_71281_n10073.n755 0.496742
R53960 a_71281_n10073.n745 a_71281_n10073.n744 0.496742
R53961 a_71281_n10073.n743 a_71281_n10073.n741 0.496742
R53962 a_71281_n10073.n731 a_71281_n10073.n730 0.496742
R53963 a_71281_n10073.n729 a_71281_n10073.n727 0.496742
R53964 a_71281_n10073.n714 a_71281_n10073.n713 0.496742
R53965 a_71281_n10073.n712 a_71281_n10073.n710 0.496742
R53966 a_71281_n10073.n700 a_71281_n10073.n699 0.496742
R53967 a_71281_n10073.n698 a_71281_n10073.n696 0.496742
R53968 a_71281_n10073.n683 a_71281_n10073.n682 0.496742
R53969 a_71281_n10073.n681 a_71281_n10073.n679 0.496742
R53970 a_71281_n10073.n669 a_71281_n10073.n668 0.496742
R53971 a_71281_n10073.n667 a_71281_n10073.n665 0.496742
R53972 a_71281_n10073.n655 a_71281_n10073.n654 0.496742
R53973 a_71281_n10073.n653 a_71281_n10073.n651 0.496742
R53974 a_71281_n10073.n642 a_71281_n10073.n641 0.496742
R53975 a_71281_n10073.n640 a_71281_n10073.n638 0.496742
R53976 a_71281_n10073.n497 a_71281_n10073.n496 0.496742
R53977 a_71281_n10073.n495 a_71281_n10073.n493 0.496742
R53978 a_71281_n10073.n771 a_71281_n10073.n769 0.496742
R53979 a_71281_n10073.n773 a_71281_n10073.n772 0.496742
R53980 a_71281_n10073.n190 a_71281_n10073.n188 0.496742
R53981 a_71281_n10073.n192 a_71281_n10073.n191 0.496742
R53982 a_71281_n10073.n491 a_71281_n10073.n345 0.445939
R53983 a_71281_n10073.n782 a_71281_n10073.n636 0.445939
R53984 a_71281_n10073.n786 a_71281_n10073.n785 0.445939
R53985 a_71281_n10073.n491 a_71281_n10073.n490 0.443507
R53986 a_71281_n10073.n782 a_71281_n10073.n781 0.443507
R53987 a_71281_n10073.n785 a_71281_n10073.n200 0.443507
R53988 a_71281_n10073.n227 a_71281_n10073.n214 0.180804
R53989 a_71281_n10073.n303 a_71281_n10073.n290 0.180804
R53990 a_71281_n10073.n476 a_71281_n10073.n463 0.180804
R53991 a_71281_n10073.n400 a_71281_n10073.n387 0.180804
R53992 a_71281_n10073.n518 a_71281_n10073.n505 0.180804
R53993 a_71281_n10073.n594 a_71281_n10073.n581 0.180804
R53994 a_71281_n10073.n767 a_71281_n10073.n754 0.180804
R53995 a_71281_n10073.n691 a_71281_n10073.n678 0.180804
R53996 a_71281_n10073.n27 a_71281_n10073.n14 0.180804
R53997 a_71281_n10073.n841 a_71281_n10073.n828 0.180804
R53998 a_71281_n10073.n186 a_71281_n10073.n173 0.180804
R53999 a_71281_n10073.n110 a_71281_n10073.n97 0.180804
R54000 a_71281_n10073.n241 a_71281_n10073.n228 0.180196
R54001 a_71281_n10073.n272 a_71281_n10073.n259 0.180196
R54002 a_71281_n10073.n286 a_71281_n10073.n273 0.180196
R54003 a_71281_n10073.n317 a_71281_n10073.n304 0.180196
R54004 a_71281_n10073.n345 a_71281_n10073.n332 0.180196
R54005 a_71281_n10073.n490 a_71281_n10073.n477 0.180196
R54006 a_71281_n10073.n462 a_71281_n10073.n449 0.180196
R54007 a_71281_n10073.n431 a_71281_n10073.n418 0.180196
R54008 a_71281_n10073.n417 a_71281_n10073.n404 0.180196
R54009 a_71281_n10073.n386 a_71281_n10073.n373 0.180196
R54010 a_71281_n10073.n532 a_71281_n10073.n519 0.180196
R54011 a_71281_n10073.n563 a_71281_n10073.n550 0.180196
R54012 a_71281_n10073.n577 a_71281_n10073.n564 0.180196
R54013 a_71281_n10073.n608 a_71281_n10073.n595 0.180196
R54014 a_71281_n10073.n636 a_71281_n10073.n623 0.180196
R54015 a_71281_n10073.n781 a_71281_n10073.n768 0.180196
R54016 a_71281_n10073.n753 a_71281_n10073.n740 0.180196
R54017 a_71281_n10073.n722 a_71281_n10073.n709 0.180196
R54018 a_71281_n10073.n708 a_71281_n10073.n695 0.180196
R54019 a_71281_n10073.n677 a_71281_n10073.n664 0.180196
R54020 a_71281_n10073.n41 a_71281_n10073.n28 0.180196
R54021 a_71281_n10073.n872 a_71281_n10073.n859 0.180196
R54022 a_71281_n10073.n858 a_71281_n10073.n845 0.180196
R54023 a_71281_n10073.n827 a_71281_n10073.n814 0.180196
R54024 a_71281_n10073.n799 a_71281_n10073.n786 0.180196
R54025 a_71281_n10073.n200 a_71281_n10073.n187 0.180196
R54026 a_71281_n10073.n172 a_71281_n10073.n159 0.180196
R54027 a_71281_n10073.n141 a_71281_n10073.n128 0.180196
R54028 a_71281_n10073.n127 a_71281_n10073.n114 0.180196
R54029 a_71281_n10073.n96 a_71281_n10073.n83 0.180196
R54030 a_71281_n10073.n255 a_71281_n10073.n242 0.179892
R54031 a_71281_n10073.n331 a_71281_n10073.n318 0.179892
R54032 a_71281_n10073.n448 a_71281_n10073.n435 0.179892
R54033 a_71281_n10073.n372 a_71281_n10073.n359 0.179892
R54034 a_71281_n10073.n546 a_71281_n10073.n533 0.179892
R54035 a_71281_n10073.n622 a_71281_n10073.n609 0.179892
R54036 a_71281_n10073.n739 a_71281_n10073.n726 0.179892
R54037 a_71281_n10073.n663 a_71281_n10073.n650 0.179892
R54038 a_71281_n10073.n55 a_71281_n10073.n42 0.179892
R54039 a_71281_n10073.n813 a_71281_n10073.n800 0.179892
R54040 a_71281_n10073.n158 a_71281_n10073.n145 0.179892
R54041 a_71281_n10073.n82 a_71281_n10073.n69 0.179892
R54042 a_71281_n10073.n26 a_71281_n10073.n15 0.136625
R54043 a_71281_n10073.n20 a_71281_n10073.n19 0.136625
R54044 a_71281_n10073.n40 a_71281_n10073.n29 0.136625
R54045 a_71281_n10073.n34 a_71281_n10073.n33 0.136625
R54046 a_71281_n10073.n54 a_71281_n10073.n43 0.136625
R54047 a_71281_n10073.n48 a_71281_n10073.n47 0.136625
R54048 a_71281_n10073.n866 a_71281_n10073.n864 0.136625
R54049 a_71281_n10073.n871 a_71281_n10073.n860 0.136625
R54050 a_71281_n10073.n852 a_71281_n10073.n850 0.136625
R54051 a_71281_n10073.n857 a_71281_n10073.n846 0.136625
R54052 a_71281_n10073.n835 a_71281_n10073.n833 0.136625
R54053 a_71281_n10073.n840 a_71281_n10073.n829 0.136625
R54054 a_71281_n10073.n821 a_71281_n10073.n819 0.136625
R54055 a_71281_n10073.n826 a_71281_n10073.n815 0.136625
R54056 a_71281_n10073.n807 a_71281_n10073.n805 0.136625
R54057 a_71281_n10073.n812 a_71281_n10073.n801 0.136625
R54058 a_71281_n10073.n793 a_71281_n10073.n791 0.136625
R54059 a_71281_n10073.n798 a_71281_n10073.n787 0.136625
R54060 a_71281_n10073.n180 a_71281_n10073.n178 0.136625
R54061 a_71281_n10073.n185 a_71281_n10073.n174 0.136625
R54062 a_71281_n10073.n166 a_71281_n10073.n164 0.136625
R54063 a_71281_n10073.n171 a_71281_n10073.n160 0.136625
R54064 a_71281_n10073.n152 a_71281_n10073.n150 0.136625
R54065 a_71281_n10073.n157 a_71281_n10073.n146 0.136625
R54066 a_71281_n10073.n135 a_71281_n10073.n133 0.136625
R54067 a_71281_n10073.n140 a_71281_n10073.n129 0.136625
R54068 a_71281_n10073.n121 a_71281_n10073.n119 0.136625
R54069 a_71281_n10073.n126 a_71281_n10073.n115 0.136625
R54070 a_71281_n10073.n104 a_71281_n10073.n102 0.136625
R54071 a_71281_n10073.n109 a_71281_n10073.n98 0.136625
R54072 a_71281_n10073.n90 a_71281_n10073.n88 0.136625
R54073 a_71281_n10073.n95 a_71281_n10073.n84 0.136625
R54074 a_71281_n10073.n76 a_71281_n10073.n74 0.136625
R54075 a_71281_n10073.n81 a_71281_n10073.n70 0.136625
R54076 a_71281_n10073.n61 a_71281_n10073.n56 0.136625
R54077 a_71281_n10073.n67 a_71281_n10073.n57 0.136625
R54078 a_71281_n10073.n6 a_71281_n10073.n1 0.136625
R54079 a_71281_n10073.n12 a_71281_n10073.n2 0.136625
R54080 a_71281_n10073.n226 a_71281_n10073.n215 0.136625
R54081 a_71281_n10073.n220 a_71281_n10073.n219 0.136625
R54082 a_71281_n10073.n240 a_71281_n10073.n229 0.136625
R54083 a_71281_n10073.n234 a_71281_n10073.n233 0.136625
R54084 a_71281_n10073.n254 a_71281_n10073.n243 0.136625
R54085 a_71281_n10073.n248 a_71281_n10073.n247 0.136625
R54086 a_71281_n10073.n271 a_71281_n10073.n260 0.136625
R54087 a_71281_n10073.n265 a_71281_n10073.n264 0.136625
R54088 a_71281_n10073.n285 a_71281_n10073.n274 0.136625
R54089 a_71281_n10073.n279 a_71281_n10073.n278 0.136625
R54090 a_71281_n10073.n302 a_71281_n10073.n291 0.136625
R54091 a_71281_n10073.n296 a_71281_n10073.n295 0.136625
R54092 a_71281_n10073.n316 a_71281_n10073.n305 0.136625
R54093 a_71281_n10073.n310 a_71281_n10073.n309 0.136625
R54094 a_71281_n10073.n330 a_71281_n10073.n319 0.136625
R54095 a_71281_n10073.n324 a_71281_n10073.n323 0.136625
R54096 a_71281_n10073.n344 a_71281_n10073.n333 0.136625
R54097 a_71281_n10073.n338 a_71281_n10073.n337 0.136625
R54098 a_71281_n10073.n470 a_71281_n10073.n468 0.136625
R54099 a_71281_n10073.n475 a_71281_n10073.n464 0.136625
R54100 a_71281_n10073.n456 a_71281_n10073.n454 0.136625
R54101 a_71281_n10073.n461 a_71281_n10073.n450 0.136625
R54102 a_71281_n10073.n442 a_71281_n10073.n440 0.136625
R54103 a_71281_n10073.n447 a_71281_n10073.n436 0.136625
R54104 a_71281_n10073.n425 a_71281_n10073.n423 0.136625
R54105 a_71281_n10073.n430 a_71281_n10073.n419 0.136625
R54106 a_71281_n10073.n411 a_71281_n10073.n409 0.136625
R54107 a_71281_n10073.n416 a_71281_n10073.n405 0.136625
R54108 a_71281_n10073.n394 a_71281_n10073.n392 0.136625
R54109 a_71281_n10073.n399 a_71281_n10073.n388 0.136625
R54110 a_71281_n10073.n380 a_71281_n10073.n378 0.136625
R54111 a_71281_n10073.n385 a_71281_n10073.n374 0.136625
R54112 a_71281_n10073.n366 a_71281_n10073.n364 0.136625
R54113 a_71281_n10073.n371 a_71281_n10073.n360 0.136625
R54114 a_71281_n10073.n351 a_71281_n10073.n346 0.136625
R54115 a_71281_n10073.n357 a_71281_n10073.n347 0.136625
R54116 a_71281_n10073.n206 a_71281_n10073.n201 0.136625
R54117 a_71281_n10073.n212 a_71281_n10073.n202 0.136625
R54118 a_71281_n10073.n489 a_71281_n10073.n478 0.136625
R54119 a_71281_n10073.n483 a_71281_n10073.n482 0.136625
R54120 a_71281_n10073.n517 a_71281_n10073.n506 0.136625
R54121 a_71281_n10073.n511 a_71281_n10073.n510 0.136625
R54122 a_71281_n10073.n531 a_71281_n10073.n520 0.136625
R54123 a_71281_n10073.n525 a_71281_n10073.n524 0.136625
R54124 a_71281_n10073.n545 a_71281_n10073.n534 0.136625
R54125 a_71281_n10073.n539 a_71281_n10073.n538 0.136625
R54126 a_71281_n10073.n562 a_71281_n10073.n551 0.136625
R54127 a_71281_n10073.n556 a_71281_n10073.n555 0.136625
R54128 a_71281_n10073.n576 a_71281_n10073.n565 0.136625
R54129 a_71281_n10073.n570 a_71281_n10073.n569 0.136625
R54130 a_71281_n10073.n593 a_71281_n10073.n582 0.136625
R54131 a_71281_n10073.n587 a_71281_n10073.n586 0.136625
R54132 a_71281_n10073.n607 a_71281_n10073.n596 0.136625
R54133 a_71281_n10073.n601 a_71281_n10073.n600 0.136625
R54134 a_71281_n10073.n621 a_71281_n10073.n610 0.136625
R54135 a_71281_n10073.n615 a_71281_n10073.n614 0.136625
R54136 a_71281_n10073.n635 a_71281_n10073.n624 0.136625
R54137 a_71281_n10073.n629 a_71281_n10073.n628 0.136625
R54138 a_71281_n10073.n761 a_71281_n10073.n759 0.136625
R54139 a_71281_n10073.n766 a_71281_n10073.n755 0.136625
R54140 a_71281_n10073.n747 a_71281_n10073.n745 0.136625
R54141 a_71281_n10073.n752 a_71281_n10073.n741 0.136625
R54142 a_71281_n10073.n733 a_71281_n10073.n731 0.136625
R54143 a_71281_n10073.n738 a_71281_n10073.n727 0.136625
R54144 a_71281_n10073.n716 a_71281_n10073.n714 0.136625
R54145 a_71281_n10073.n721 a_71281_n10073.n710 0.136625
R54146 a_71281_n10073.n702 a_71281_n10073.n700 0.136625
R54147 a_71281_n10073.n707 a_71281_n10073.n696 0.136625
R54148 a_71281_n10073.n685 a_71281_n10073.n683 0.136625
R54149 a_71281_n10073.n690 a_71281_n10073.n679 0.136625
R54150 a_71281_n10073.n671 a_71281_n10073.n669 0.136625
R54151 a_71281_n10073.n676 a_71281_n10073.n665 0.136625
R54152 a_71281_n10073.n657 a_71281_n10073.n655 0.136625
R54153 a_71281_n10073.n662 a_71281_n10073.n651 0.136625
R54154 a_71281_n10073.n642 a_71281_n10073.n637 0.136625
R54155 a_71281_n10073.n648 a_71281_n10073.n638 0.136625
R54156 a_71281_n10073.n497 a_71281_n10073.n492 0.136625
R54157 a_71281_n10073.n503 a_71281_n10073.n493 0.136625
R54158 a_71281_n10073.n780 a_71281_n10073.n769 0.136625
R54159 a_71281_n10073.n774 a_71281_n10073.n773 0.136625
R54160 a_71281_n10073.n199 a_71281_n10073.n188 0.136625
R54161 a_71281_n10073.n193 a_71281_n10073.n192 0.136625
R54162 a_71281_n10073.n214 a_71281_n10073.n213 0.095973
R54163 a_71281_n10073.n228 a_71281_n10073.n227 0.095973
R54164 a_71281_n10073.n242 a_71281_n10073.n241 0.095973
R54165 a_71281_n10073.n273 a_71281_n10073.n272 0.095973
R54166 a_71281_n10073.n304 a_71281_n10073.n303 0.095973
R54167 a_71281_n10073.n318 a_71281_n10073.n317 0.095973
R54168 a_71281_n10073.n332 a_71281_n10073.n331 0.095973
R54169 a_71281_n10073.n477 a_71281_n10073.n476 0.095973
R54170 a_71281_n10073.n463 a_71281_n10073.n462 0.095973
R54171 a_71281_n10073.n449 a_71281_n10073.n448 0.095973
R54172 a_71281_n10073.n418 a_71281_n10073.n417 0.095973
R54173 a_71281_n10073.n387 a_71281_n10073.n386 0.095973
R54174 a_71281_n10073.n373 a_71281_n10073.n372 0.095973
R54175 a_71281_n10073.n359 a_71281_n10073.n358 0.095973
R54176 a_71281_n10073.n505 a_71281_n10073.n504 0.095973
R54177 a_71281_n10073.n519 a_71281_n10073.n518 0.095973
R54178 a_71281_n10073.n533 a_71281_n10073.n532 0.095973
R54179 a_71281_n10073.n564 a_71281_n10073.n563 0.095973
R54180 a_71281_n10073.n595 a_71281_n10073.n594 0.095973
R54181 a_71281_n10073.n609 a_71281_n10073.n608 0.095973
R54182 a_71281_n10073.n623 a_71281_n10073.n622 0.095973
R54183 a_71281_n10073.n768 a_71281_n10073.n767 0.095973
R54184 a_71281_n10073.n754 a_71281_n10073.n753 0.095973
R54185 a_71281_n10073.n740 a_71281_n10073.n739 0.095973
R54186 a_71281_n10073.n709 a_71281_n10073.n708 0.095973
R54187 a_71281_n10073.n678 a_71281_n10073.n677 0.095973
R54188 a_71281_n10073.n664 a_71281_n10073.n663 0.095973
R54189 a_71281_n10073.n650 a_71281_n10073.n649 0.095973
R54190 a_71281_n10073.n14 a_71281_n10073.n13 0.095973
R54191 a_71281_n10073.n28 a_71281_n10073.n27 0.095973
R54192 a_71281_n10073.n42 a_71281_n10073.n41 0.095973
R54193 a_71281_n10073.n859 a_71281_n10073.n858 0.095973
R54194 a_71281_n10073.n828 a_71281_n10073.n827 0.095973
R54195 a_71281_n10073.n814 a_71281_n10073.n813 0.095973
R54196 a_71281_n10073.n800 a_71281_n10073.n799 0.095973
R54197 a_71281_n10073.n187 a_71281_n10073.n186 0.095973
R54198 a_71281_n10073.n173 a_71281_n10073.n172 0.095973
R54199 a_71281_n10073.n159 a_71281_n10073.n158 0.095973
R54200 a_71281_n10073.n128 a_71281_n10073.n127 0.095973
R54201 a_71281_n10073.n97 a_71281_n10073.n96 0.095973
R54202 a_71281_n10073.n83 a_71281_n10073.n82 0.095973
R54203 a_71281_n10073.n69 a_71281_n10073.n68 0.095973
R54204 a_71281_n10073.n26 a_71281_n10073.n25 0.0719743
R54205 a_71281_n10073.n22 a_71281_n10073.n20 0.0719743
R54206 a_71281_n10073.n40 a_71281_n10073.n39 0.0719743
R54207 a_71281_n10073.n36 a_71281_n10073.n34 0.0719743
R54208 a_71281_n10073.n54 a_71281_n10073.n53 0.0719743
R54209 a_71281_n10073.n50 a_71281_n10073.n48 0.0719743
R54210 a_71281_n10073.n867 a_71281_n10073.n866 0.0719743
R54211 a_71281_n10073.n871 a_71281_n10073.n870 0.0719743
R54212 a_71281_n10073.n853 a_71281_n10073.n852 0.0719743
R54213 a_71281_n10073.n857 a_71281_n10073.n856 0.0719743
R54214 a_71281_n10073.n836 a_71281_n10073.n835 0.0719743
R54215 a_71281_n10073.n840 a_71281_n10073.n839 0.0719743
R54216 a_71281_n10073.n822 a_71281_n10073.n821 0.0719743
R54217 a_71281_n10073.n826 a_71281_n10073.n825 0.0719743
R54218 a_71281_n10073.n808 a_71281_n10073.n807 0.0719743
R54219 a_71281_n10073.n812 a_71281_n10073.n811 0.0719743
R54220 a_71281_n10073.n794 a_71281_n10073.n793 0.0719743
R54221 a_71281_n10073.n798 a_71281_n10073.n797 0.0719743
R54222 a_71281_n10073.n181 a_71281_n10073.n180 0.0719743
R54223 a_71281_n10073.n185 a_71281_n10073.n184 0.0719743
R54224 a_71281_n10073.n167 a_71281_n10073.n166 0.0719743
R54225 a_71281_n10073.n171 a_71281_n10073.n170 0.0719743
R54226 a_71281_n10073.n153 a_71281_n10073.n152 0.0719743
R54227 a_71281_n10073.n157 a_71281_n10073.n156 0.0719743
R54228 a_71281_n10073.n136 a_71281_n10073.n135 0.0719743
R54229 a_71281_n10073.n140 a_71281_n10073.n139 0.0719743
R54230 a_71281_n10073.n122 a_71281_n10073.n121 0.0719743
R54231 a_71281_n10073.n126 a_71281_n10073.n125 0.0719743
R54232 a_71281_n10073.n105 a_71281_n10073.n104 0.0719743
R54233 a_71281_n10073.n109 a_71281_n10073.n108 0.0719743
R54234 a_71281_n10073.n91 a_71281_n10073.n90 0.0719743
R54235 a_71281_n10073.n95 a_71281_n10073.n94 0.0719743
R54236 a_71281_n10073.n77 a_71281_n10073.n76 0.0719743
R54237 a_71281_n10073.n81 a_71281_n10073.n80 0.0719743
R54238 a_71281_n10073.n63 a_71281_n10073.n56 0.0719743
R54239 a_71281_n10073.n67 a_71281_n10073.n66 0.0719743
R54240 a_71281_n10073.n8 a_71281_n10073.n1 0.0719743
R54241 a_71281_n10073.n12 a_71281_n10073.n11 0.0719743
R54242 a_71281_n10073.n226 a_71281_n10073.n225 0.0719743
R54243 a_71281_n10073.n222 a_71281_n10073.n220 0.0719743
R54244 a_71281_n10073.n240 a_71281_n10073.n239 0.0719743
R54245 a_71281_n10073.n236 a_71281_n10073.n234 0.0719743
R54246 a_71281_n10073.n254 a_71281_n10073.n253 0.0719743
R54247 a_71281_n10073.n250 a_71281_n10073.n248 0.0719743
R54248 a_71281_n10073.n271 a_71281_n10073.n270 0.0719743
R54249 a_71281_n10073.n267 a_71281_n10073.n265 0.0719743
R54250 a_71281_n10073.n285 a_71281_n10073.n284 0.0719743
R54251 a_71281_n10073.n281 a_71281_n10073.n279 0.0719743
R54252 a_71281_n10073.n302 a_71281_n10073.n301 0.0719743
R54253 a_71281_n10073.n298 a_71281_n10073.n296 0.0719743
R54254 a_71281_n10073.n316 a_71281_n10073.n315 0.0719743
R54255 a_71281_n10073.n312 a_71281_n10073.n310 0.0719743
R54256 a_71281_n10073.n330 a_71281_n10073.n329 0.0719743
R54257 a_71281_n10073.n326 a_71281_n10073.n324 0.0719743
R54258 a_71281_n10073.n344 a_71281_n10073.n343 0.0719743
R54259 a_71281_n10073.n340 a_71281_n10073.n338 0.0719743
R54260 a_71281_n10073.n471 a_71281_n10073.n470 0.0719743
R54261 a_71281_n10073.n475 a_71281_n10073.n474 0.0719743
R54262 a_71281_n10073.n457 a_71281_n10073.n456 0.0719743
R54263 a_71281_n10073.n461 a_71281_n10073.n460 0.0719743
R54264 a_71281_n10073.n443 a_71281_n10073.n442 0.0719743
R54265 a_71281_n10073.n447 a_71281_n10073.n446 0.0719743
R54266 a_71281_n10073.n426 a_71281_n10073.n425 0.0719743
R54267 a_71281_n10073.n430 a_71281_n10073.n429 0.0719743
R54268 a_71281_n10073.n412 a_71281_n10073.n411 0.0719743
R54269 a_71281_n10073.n416 a_71281_n10073.n415 0.0719743
R54270 a_71281_n10073.n395 a_71281_n10073.n394 0.0719743
R54271 a_71281_n10073.n399 a_71281_n10073.n398 0.0719743
R54272 a_71281_n10073.n381 a_71281_n10073.n380 0.0719743
R54273 a_71281_n10073.n385 a_71281_n10073.n384 0.0719743
R54274 a_71281_n10073.n367 a_71281_n10073.n366 0.0719743
R54275 a_71281_n10073.n371 a_71281_n10073.n370 0.0719743
R54276 a_71281_n10073.n353 a_71281_n10073.n346 0.0719743
R54277 a_71281_n10073.n357 a_71281_n10073.n356 0.0719743
R54278 a_71281_n10073.n208 a_71281_n10073.n201 0.0719743
R54279 a_71281_n10073.n212 a_71281_n10073.n211 0.0719743
R54280 a_71281_n10073.n489 a_71281_n10073.n488 0.0719743
R54281 a_71281_n10073.n485 a_71281_n10073.n483 0.0719743
R54282 a_71281_n10073.n517 a_71281_n10073.n516 0.0719743
R54283 a_71281_n10073.n513 a_71281_n10073.n511 0.0719743
R54284 a_71281_n10073.n531 a_71281_n10073.n530 0.0719743
R54285 a_71281_n10073.n527 a_71281_n10073.n525 0.0719743
R54286 a_71281_n10073.n545 a_71281_n10073.n544 0.0719743
R54287 a_71281_n10073.n541 a_71281_n10073.n539 0.0719743
R54288 a_71281_n10073.n562 a_71281_n10073.n561 0.0719743
R54289 a_71281_n10073.n558 a_71281_n10073.n556 0.0719743
R54290 a_71281_n10073.n576 a_71281_n10073.n575 0.0719743
R54291 a_71281_n10073.n572 a_71281_n10073.n570 0.0719743
R54292 a_71281_n10073.n593 a_71281_n10073.n592 0.0719743
R54293 a_71281_n10073.n589 a_71281_n10073.n587 0.0719743
R54294 a_71281_n10073.n607 a_71281_n10073.n606 0.0719743
R54295 a_71281_n10073.n603 a_71281_n10073.n601 0.0719743
R54296 a_71281_n10073.n621 a_71281_n10073.n620 0.0719743
R54297 a_71281_n10073.n617 a_71281_n10073.n615 0.0719743
R54298 a_71281_n10073.n635 a_71281_n10073.n634 0.0719743
R54299 a_71281_n10073.n631 a_71281_n10073.n629 0.0719743
R54300 a_71281_n10073.n762 a_71281_n10073.n761 0.0719743
R54301 a_71281_n10073.n766 a_71281_n10073.n765 0.0719743
R54302 a_71281_n10073.n748 a_71281_n10073.n747 0.0719743
R54303 a_71281_n10073.n752 a_71281_n10073.n751 0.0719743
R54304 a_71281_n10073.n734 a_71281_n10073.n733 0.0719743
R54305 a_71281_n10073.n738 a_71281_n10073.n737 0.0719743
R54306 a_71281_n10073.n717 a_71281_n10073.n716 0.0719743
R54307 a_71281_n10073.n721 a_71281_n10073.n720 0.0719743
R54308 a_71281_n10073.n703 a_71281_n10073.n702 0.0719743
R54309 a_71281_n10073.n707 a_71281_n10073.n706 0.0719743
R54310 a_71281_n10073.n686 a_71281_n10073.n685 0.0719743
R54311 a_71281_n10073.n690 a_71281_n10073.n689 0.0719743
R54312 a_71281_n10073.n672 a_71281_n10073.n671 0.0719743
R54313 a_71281_n10073.n676 a_71281_n10073.n675 0.0719743
R54314 a_71281_n10073.n658 a_71281_n10073.n657 0.0719743
R54315 a_71281_n10073.n662 a_71281_n10073.n661 0.0719743
R54316 a_71281_n10073.n644 a_71281_n10073.n637 0.0719743
R54317 a_71281_n10073.n648 a_71281_n10073.n647 0.0719743
R54318 a_71281_n10073.n499 a_71281_n10073.n492 0.0719743
R54319 a_71281_n10073.n503 a_71281_n10073.n502 0.0719743
R54320 a_71281_n10073.n780 a_71281_n10073.n779 0.0719743
R54321 a_71281_n10073.n776 a_71281_n10073.n774 0.0719743
R54322 a_71281_n10073.n199 a_71281_n10073.n198 0.0719743
R54323 a_71281_n10073.n195 a_71281_n10073.n193 0.0719743
R54324 a_71281_n10073.n289 a_71281_n10073.n286 0.0485405
R54325 a_71281_n10073.n404 a_71281_n10073.n403 0.0485405
R54326 a_71281_n10073.n580 a_71281_n10073.n577 0.0485405
R54327 a_71281_n10073.n695 a_71281_n10073.n694 0.0485405
R54328 a_71281_n10073.n845 a_71281_n10073.n844 0.0485405
R54329 a_71281_n10073.n114 a_71281_n10073.n113 0.0485405
R54330 a_71281_n10073.n258 a_71281_n10073.n255 0.0482365
R54331 a_71281_n10073.n259 a_71281_n10073.n258 0.0482365
R54332 a_71281_n10073.n435 a_71281_n10073.n434 0.0482365
R54333 a_71281_n10073.n434 a_71281_n10073.n431 0.0482365
R54334 a_71281_n10073.n549 a_71281_n10073.n546 0.0482365
R54335 a_71281_n10073.n550 a_71281_n10073.n549 0.0482365
R54336 a_71281_n10073.n726 a_71281_n10073.n725 0.0482365
R54337 a_71281_n10073.n725 a_71281_n10073.n722 0.0482365
R54338 a_71281_n10073.n873 a_71281_n10073.n55 0.0482365
R54339 a_71281_n10073.n873 a_71281_n10073.n872 0.0482365
R54340 a_71281_n10073.n145 a_71281_n10073.n144 0.0482365
R54341 a_71281_n10073.n144 a_71281_n10073.n141 0.0482365
R54342 a_71281_n10073.n290 a_71281_n10073.n289 0.0479324
R54343 a_71281_n10073.n403 a_71281_n10073.n400 0.0479324
R54344 a_71281_n10073.n581 a_71281_n10073.n580 0.0479324
R54345 a_71281_n10073.n694 a_71281_n10073.n691 0.0479324
R54346 a_71281_n10073.n844 a_71281_n10073.n841 0.0479324
R54347 a_71281_n10073.n113 a_71281_n10073.n110 0.0479324
R54348 a_71281_n10073.t1 a_71281_n10073.n0 3.76597
R54349 a_60677_10448.t2 a_60677_10448.t4 60.937
R54350 a_60677_10448.t0 a_60677_10448.t2 12.9273
R54351 a_60677_10448.t2 a_60677_10448.t5 10.1307
R54352 a_60677_10448.t2 a_60677_10448.t1 8.54643
R54353 a_60677_10448.t2 a_60677_10448.t3 7.50895
R54354 a_33379_34007.t2 a_33379_34007.n351 10.937
R54355 a_33379_34007.t27 a_33379_34007.n350 9.74618
R54356 a_33379_34007.n351 a_33379_34007.t3 9.33982
R54357 a_33379_34007.n180 a_33379_34007.t8 8.38704
R54358 a_33379_34007.n305 a_33379_34007.t20 8.38704
R54359 a_33379_34007.n139 a_33379_34007.t33 8.37857
R54360 a_33379_34007.n286 a_33379_34007.t36 8.37857
R54361 a_33379_34007.n55 a_33379_34007.t40 8.39293
R54362 a_33379_34007.n83 a_33379_34007.t50 8.39293
R54363 a_33379_34007.n37 a_33379_34007.t45 8.10567
R54364 a_33379_34007.n133 a_33379_34007.t19 8.10567
R54365 a_33379_34007.n6 a_33379_34007.t78 8.10567
R54366 a_33379_34007.n25 a_33379_34007.t48 8.10567
R54367 a_33379_34007.n148 a_33379_34007.t39 8.10567
R54368 a_33379_34007.n149 a_33379_34007.t91 8.10567
R54369 a_33379_34007.n150 a_33379_34007.t63 8.10567
R54370 a_33379_34007.n138 a_33379_34007.t13 8.10567
R54371 a_33379_34007.n3 a_33379_34007.t73 8.10567
R54372 a_33379_34007.n23 a_33379_34007.t12 8.10567
R54373 a_33379_34007.n42 a_33379_34007.t74 8.10567
R54374 a_33379_34007.n120 a_33379_34007.t47 8.10567
R54375 a_33379_34007.n12 a_33379_34007.t21 8.10567
R54376 a_33379_34007.n128 a_33379_34007.t61 8.10567
R54377 a_33379_34007.n127 a_33379_34007.t11 8.10567
R54378 a_33379_34007.n126 a_33379_34007.t72 8.10567
R54379 a_33379_34007.n38 a_33379_34007.t38 8.10567
R54380 a_33379_34007.n130 a_33379_34007.t10 8.10567
R54381 a_33379_34007.n9 a_33379_34007.t80 8.10567
R54382 a_33379_34007.n29 a_33379_34007.t41 8.10567
R54383 a_33379_34007.n60 a_33379_34007.t56 8.10567
R54384 a_33379_34007.n58 a_33379_34007.t28 8.10567
R54385 a_33379_34007.n56 a_33379_34007.t85 8.10567
R54386 a_33379_34007.n222 a_33379_34007.t60 8.10567
R54387 a_33379_34007.n207 a_33379_34007.t34 8.10567
R54388 a_33379_34007.n208 a_33379_34007.t86 8.10567
R54389 a_33379_34007.n209 a_33379_34007.t58 8.10567
R54390 a_33379_34007.n54 a_33379_34007.t26 8.10567
R54391 a_33379_34007.n53 a_33379_34007.t82 8.10567
R54392 a_33379_34007.n51 a_33379_34007.t25 8.10567
R54393 a_33379_34007.n75 a_33379_34007.t84 8.10567
R54394 a_33379_34007.n72 a_33379_34007.t57 8.10567
R54395 a_33379_34007.n179 a_33379_34007.t29 8.10567
R54396 a_33379_34007.n189 a_33379_34007.t55 8.10567
R54397 a_33379_34007.n188 a_33379_34007.t4 8.10567
R54398 a_33379_34007.n187 a_33379_34007.t67 8.10567
R54399 a_33379_34007.n68 a_33379_34007.t49 8.10567
R54400 a_33379_34007.n67 a_33379_34007.t22 8.10567
R54401 a_33379_34007.n66 a_33379_34007.t88 8.10567
R54402 a_33379_34007.n63 a_33379_34007.t53 8.10567
R54403 a_33379_34007.n45 a_33379_34007.t51 8.10567
R54404 a_33379_34007.n275 a_33379_34007.t23 8.10567
R54405 a_33379_34007.n18 a_33379_34007.t81 8.10567
R54406 a_33379_34007.n33 a_33379_34007.t54 8.10567
R54407 a_33379_34007.n283 a_33379_34007.t44 8.10567
R54408 a_33379_34007.n282 a_33379_34007.t7 8.10567
R54409 a_33379_34007.n281 a_33379_34007.t70 8.10567
R54410 a_33379_34007.n285 a_33379_34007.t18 8.10567
R54411 a_33379_34007.n15 a_33379_34007.t77 8.10567
R54412 a_33379_34007.n32 a_33379_34007.t17 8.10567
R54413 a_33379_34007.n50 a_33379_34007.t79 8.10567
R54414 a_33379_34007.n243 a_33379_34007.t52 8.10567
R54415 a_33379_34007.n20 a_33379_34007.t24 8.10567
R54416 a_33379_34007.n254 a_33379_34007.t66 8.10567
R54417 a_33379_34007.n253 a_33379_34007.t16 8.10567
R54418 a_33379_34007.n252 a_33379_34007.t76 8.10567
R54419 a_33379_34007.n47 a_33379_34007.t42 8.10567
R54420 a_33379_34007.n264 a_33379_34007.t14 8.10567
R54421 a_33379_34007.n19 a_33379_34007.t83 8.10567
R54422 a_33379_34007.n36 a_33379_34007.t46 8.10567
R54423 a_33379_34007.n92 a_33379_34007.t65 8.10567
R54424 a_33379_34007.n89 a_33379_34007.t35 8.10567
R54425 a_33379_34007.n86 a_33379_34007.t5 8.10567
R54426 a_33379_34007.n298 a_33379_34007.t71 8.10567
R54427 a_33379_34007.n339 a_33379_34007.t43 8.10567
R54428 a_33379_34007.n338 a_33379_34007.t6 8.10567
R54429 a_33379_34007.n337 a_33379_34007.t69 8.10567
R54430 a_33379_34007.n82 a_33379_34007.t32 8.10567
R54431 a_33379_34007.n81 a_33379_34007.t89 8.10567
R54432 a_33379_34007.n78 a_33379_34007.t31 8.10567
R54433 a_33379_34007.n106 a_33379_34007.t92 8.10567
R54434 a_33379_34007.n104 a_33379_34007.t68 8.10567
R54435 a_33379_34007.n304 a_33379_34007.t37 8.10567
R54436 a_33379_34007.n317 a_33379_34007.t64 8.10567
R54437 a_33379_34007.n316 a_33379_34007.t15 8.10567
R54438 a_33379_34007.n315 a_33379_34007.t75 8.10567
R54439 a_33379_34007.n101 a_33379_34007.t59 8.10567
R54440 a_33379_34007.n99 a_33379_34007.t30 8.10567
R54441 a_33379_34007.n96 a_33379_34007.t9 8.10567
R54442 a_33379_34007.n94 a_33379_34007.t62 8.10567
R54443 a_33379_34007.n350 a_33379_34007.n349 6.72496
R54444 a_33379_34007.n69 a_33379_34007.n68 2.25163
R54445 a_33379_34007.n102 a_33379_34007.n101 2.25163
R54446 a_33379_34007.n39 a_33379_34007.n38 2.24588
R54447 a_33379_34007.n48 a_33379_34007.n47 2.24588
R54448 a_33379_34007.n26 a_33379_34007.n25 2.2453
R54449 a_33379_34007.n34 a_33379_34007.n33 2.2453
R54450 a_33379_34007.n117 a_33379_34007.n11 4.5005
R54451 a_33379_34007.n119 a_33379_34007.n118 4.5005
R54452 a_33379_34007.n121 a_33379_34007.n116 4.5005
R54453 a_33379_34007.n123 a_33379_34007.n122 4.5005
R54454 a_33379_34007.n124 a_33379_34007.n41 4.5005
R54455 a_33379_34007.n42 a_33379_34007.n40 4.5005
R54456 a_33379_34007.n125 a_33379_34007.n115 4.5005
R54457 a_33379_34007.n175 a_33379_34007.n174 4.5005
R54458 a_33379_34007.n29 a_33379_34007.n27 4.5005
R54459 a_33379_34007.n28 a_33379_34007.n173 4.5005
R54460 a_33379_34007.n172 a_33379_34007.n8 4.5005
R54461 a_33379_34007.n171 a_33379_34007.n9 4.5005
R54462 a_33379_34007.n7 a_33379_34007.n129 4.5005
R54463 a_33379_34007.n170 a_33379_34007.n169 4.5005
R54464 a_33379_34007.n168 a_33379_34007.n167 4.5005
R54465 a_33379_34007.n166 a_33379_34007.n131 4.5005
R54466 a_33379_34007.n165 a_33379_34007.n164 4.5005
R54467 a_33379_34007.n24 a_33379_34007.n163 4.5005
R54468 a_33379_34007.n162 a_33379_34007.n5 4.5005
R54469 a_33379_34007.n161 a_33379_34007.n6 4.5005
R54470 a_33379_34007.n4 a_33379_34007.n132 4.5005
R54471 a_33379_34007.n160 a_33379_34007.n159 4.5005
R54472 a_33379_34007.n158 a_33379_34007.n157 4.5005
R54473 a_33379_34007.n156 a_33379_34007.n134 4.5005
R54474 a_33379_34007.n155 a_33379_34007.n154 4.5005
R54475 a_33379_34007.n153 a_33379_34007.n37 4.5005
R54476 a_33379_34007.n152 a_33379_34007.n151 4.5005
R54477 a_33379_34007.n147 a_33379_34007.n146 4.5005
R54478 a_33379_34007.n145 a_33379_34007.n23 4.5005
R54479 a_33379_34007.n22 a_33379_34007.n136 4.5005
R54480 a_33379_34007.n144 a_33379_34007.n143 4.5005
R54481 a_33379_34007.n142 a_33379_34007.n3 4.5005
R54482 a_33379_34007.n2 a_33379_34007.n137 4.5005
R54483 a_33379_34007.n141 a_33379_34007.n140 4.5005
R54484 a_33379_34007.n186 a_33379_34007.n177 4.5005
R54485 a_33379_34007.n75 a_33379_34007.n73 4.5005
R54486 a_33379_34007.n185 a_33379_34007.n74 4.5005
R54487 a_33379_34007.n184 a_33379_34007.n183 4.5005
R54488 a_33379_34007.n72 a_33379_34007.n70 4.5005
R54489 a_33379_34007.n71 a_33379_34007.n182 4.5005
R54490 a_33379_34007.n181 a_33379_34007.n178 4.5005
R54491 a_33379_34007.n234 a_33379_34007.n233 4.5005
R54492 a_33379_34007.n63 a_33379_34007.n61 4.5005
R54493 a_33379_34007.n62 a_33379_34007.n232 4.5005
R54494 a_33379_34007.n231 a_33379_34007.n64 4.5005
R54495 a_33379_34007.n230 a_33379_34007.n66 4.5005
R54496 a_33379_34007.n65 a_33379_34007.n190 4.5005
R54497 a_33379_34007.n229 a_33379_34007.n228 4.5005
R54498 a_33379_34007.n227 a_33379_34007.n67 4.5005
R54499 a_33379_34007.n226 a_33379_34007.n225 4.5005
R54500 a_33379_34007.n224 a_33379_34007.n191 4.5005
R54501 a_33379_34007.n211 a_33379_34007.n210 4.5005
R54502 a_33379_34007.n60 a_33379_34007.n59 4.5005
R54503 a_33379_34007.n212 a_33379_34007.n194 4.5005
R54504 a_33379_34007.n214 a_33379_34007.n213 4.5005
R54505 a_33379_34007.n58 a_33379_34007.n57 4.5005
R54506 a_33379_34007.n215 a_33379_34007.n193 4.5005
R54507 a_33379_34007.n217 a_33379_34007.n216 4.5005
R54508 a_33379_34007.n218 a_33379_34007.n56 4.5005
R54509 a_33379_34007.n220 a_33379_34007.n219 4.5005
R54510 a_33379_34007.n221 a_33379_34007.n192 4.5005
R54511 a_33379_34007.n206 a_33379_34007.n205 4.5005
R54512 a_33379_34007.n204 a_33379_34007.n51 4.5005
R54513 a_33379_34007.n203 a_33379_34007.n202 4.5005
R54514 a_33379_34007.n201 a_33379_34007.n196 4.5005
R54515 a_33379_34007.n53 a_33379_34007.n52 4.5005
R54516 a_33379_34007.n200 a_33379_34007.n199 4.5005
R54517 a_33379_34007.n198 a_33379_34007.n197 4.5005
R54518 a_33379_34007.n242 a_33379_34007.n241 4.5005
R54519 a_33379_34007.n245 a_33379_34007.n244 4.5005
R54520 a_33379_34007.n246 a_33379_34007.n240 4.5005
R54521 a_33379_34007.n248 a_33379_34007.n247 4.5005
R54522 a_33379_34007.n49 a_33379_34007.n239 4.5005
R54523 a_33379_34007.n249 a_33379_34007.n50 4.5005
R54524 a_33379_34007.n251 a_33379_34007.n250 4.5005
R54525 a_33379_34007.n256 a_33379_34007.n255 4.5005
R54526 a_33379_34007.n36 a_33379_34007.n35 4.5005
R54527 a_33379_34007.n257 a_33379_34007.n114 4.5005
R54528 a_33379_34007.n259 a_33379_34007.n258 4.5005
R54529 a_33379_34007.n260 a_33379_34007.n19 4.5005
R54530 a_33379_34007.n262 a_33379_34007.n261 4.5005
R54531 a_33379_34007.n263 a_33379_34007.n113 4.5005
R54532 a_33379_34007.n266 a_33379_34007.n265 4.5005
R54533 a_33379_34007.n267 a_33379_34007.n112 4.5005
R54534 a_33379_34007.n46 a_33379_34007.n268 4.5005
R54535 a_33379_34007.n270 a_33379_34007.n269 4.5005
R54536 a_33379_34007.n17 a_33379_34007.n111 4.5005
R54537 a_33379_34007.n271 a_33379_34007.n18 4.5005
R54538 a_33379_34007.n272 a_33379_34007.n16 4.5005
R54539 a_33379_34007.n274 a_33379_34007.n273 4.5005
R54540 a_33379_34007.n276 a_33379_34007.n110 4.5005
R54541 a_33379_34007.n278 a_33379_34007.n277 4.5005
R54542 a_33379_34007.n279 a_33379_34007.n44 4.5005
R54543 a_33379_34007.n45 a_33379_34007.n43 4.5005
R54544 a_33379_34007.n280 a_33379_34007.n109 4.5005
R54545 a_33379_34007.n293 a_33379_34007.n292 4.5005
R54546 a_33379_34007.n32 a_33379_34007.n30 4.5005
R54547 a_33379_34007.n31 a_33379_34007.n291 4.5005
R54548 a_33379_34007.n290 a_33379_34007.n14 4.5005
R54549 a_33379_34007.n289 a_33379_34007.n15 4.5005
R54550 a_33379_34007.n13 a_33379_34007.n284 4.5005
R54551 a_33379_34007.n288 a_33379_34007.n287 4.5005
R54552 a_33379_34007.n314 a_33379_34007.n313 4.5005
R54553 a_33379_34007.n311 a_33379_34007.n106 4.5005
R54554 a_33379_34007.n105 a_33379_34007.n302 4.5005
R54555 a_33379_34007.n310 a_33379_34007.n309 4.5005
R54556 a_33379_34007.n308 a_33379_34007.n104 4.5005
R54557 a_33379_34007.n103 a_33379_34007.n303 4.5005
R54558 a_33379_34007.n307 a_33379_34007.n306 4.5005
R54559 a_33379_34007.n93 a_33379_34007.n301 4.5005
R54560 a_33379_34007.n318 a_33379_34007.n94 4.5005
R54561 a_33379_34007.n320 a_33379_34007.n319 4.5005
R54562 a_33379_34007.n95 a_33379_34007.n300 4.5005
R54563 a_33379_34007.n321 a_33379_34007.n96 4.5005
R54564 a_33379_34007.n323 a_33379_34007.n322 4.5005
R54565 a_33379_34007.n97 a_33379_34007.n299 4.5005
R54566 a_33379_34007.n324 a_33379_34007.n99 4.5005
R54567 a_33379_34007.n325 a_33379_34007.n98 4.5005
R54568 a_33379_34007.n100 a_33379_34007.n326 4.5005
R54569 a_33379_34007.n336 a_33379_34007.n296 4.5005
R54570 a_33379_34007.n92 a_33379_34007.n90 4.5005
R54571 a_33379_34007.n335 a_33379_34007.n91 4.5005
R54572 a_33379_34007.n334 a_33379_34007.n333 4.5005
R54573 a_33379_34007.n89 a_33379_34007.n87 4.5005
R54574 a_33379_34007.n88 a_33379_34007.n332 4.5005
R54575 a_33379_34007.n331 a_33379_34007.n85 4.5005
R54576 a_33379_34007.n330 a_33379_34007.n86 4.5005
R54577 a_33379_34007.n84 a_33379_34007.n297 4.5005
R54578 a_33379_34007.n329 a_33379_34007.n328 4.5005
R54579 a_33379_34007.n347 a_33379_34007.n346 4.5005
R54580 a_33379_34007.n78 a_33379_34007.n76 4.5005
R54581 a_33379_34007.n77 a_33379_34007.n345 4.5005
R54582 a_33379_34007.n344 a_33379_34007.n79 4.5005
R54583 a_33379_34007.n343 a_33379_34007.n81 4.5005
R54584 a_33379_34007.n80 a_33379_34007.n340 4.5005
R54585 a_33379_34007.n342 a_33379_34007.n341 4.5005
R54586 a_33379_34007.n1 a_33379_34007.n0 0.49013
R54587 a_33379_34007.t27 a_33379_34007.n1 7.88634
R54588 a_33379_34007.n135 a_33379_34007.n108 2.30989
R54589 a_33379_34007.n236 a_33379_34007.n176 2.30989
R54590 a_33379_34007.n223 a_33379_34007.n222 2.25752
R54591 a_33379_34007.n327 a_33379_34007.n298 2.25752
R54592 a_33379_34007.n176 a_33379_34007.n115 2.18975
R54593 a_33379_34007.n152 a_33379_34007.n135 2.18975
R54594 a_33379_34007.n250 a_33379_34007.n238 2.18975
R54595 a_33379_34007.n294 a_33379_34007.n109 2.18975
R54596 a_33379_34007.n235 a_33379_34007.n177 2.16725
R54597 a_33379_34007.n211 a_33379_34007.n195 2.16725
R54598 a_33379_34007.n313 a_33379_34007.n312 2.16725
R54599 a_33379_34007.n348 a_33379_34007.n296 2.16725
R54600 a_33379_34007.n349 a_33379_34007.n348 1.5005
R54601 a_33379_34007.n295 a_33379_34007.n294 1.5005
R54602 a_33379_34007.n195 a_33379_34007.n108 1.5005
R54603 a_33379_34007.n312 a_33379_34007.n107 1.5005
R54604 a_33379_34007.n238 a_33379_34007.n237 1.5005
R54605 a_33379_34007.n236 a_33379_34007.n235 1.5005
R54606 a_33379_34007.n10 a_33379_34007.t87 8.40801
R54607 a_33379_34007.n21 a_33379_34007.t90 8.40801
R54608 a_33379_34007.n148 a_33379_34007.n147 1.24866
R54609 a_33379_34007.n174 a_33379_34007.n128 1.24866
R54610 a_33379_34007.n292 a_33379_34007.n283 1.24866
R54611 a_33379_34007.n255 a_33379_34007.n254 1.24866
R54612 a_33379_34007.n151 a_33379_34007.n150 1.24629
R54613 a_33379_34007.n126 a_33379_34007.n125 1.24629
R54614 a_33379_34007.n281 a_33379_34007.n280 1.24629
R54615 a_33379_34007.n252 a_33379_34007.n251 1.24629
R54616 a_33379_34007.n295 a_33379_34007.n108 1.23709
R54617 a_33379_34007.n237 a_33379_34007.n236 1.23709
R54618 a_33379_34007.n210 a_33379_34007.n209 1.22261
R54619 a_33379_34007.n187 a_33379_34007.n186 1.22261
R54620 a_33379_34007.n337 a_33379_34007.n336 1.22261
R54621 a_33379_34007.n315 a_33379_34007.n314 1.22261
R54622 a_33379_34007.n207 a_33379_34007.n206 1.21313
R54623 a_33379_34007.n233 a_33379_34007.n189 1.21313
R54624 a_33379_34007.n346 a_33379_34007.n339 1.21313
R54625 a_33379_34007.n93 a_33379_34007.n317 1.21313
R54626 a_33379_34007.n181 a_33379_34007.n180 1.12904
R54627 a_33379_34007.n306 a_33379_34007.n305 1.12904
R54628 a_33379_34007.n140 a_33379_34007.n139 1.11862
R54629 a_33379_34007.n287 a_33379_34007.n286 1.11862
R54630 a_33379_34007.n349 a_33379_34007.n295 0.809892
R54631 a_33379_34007.n237 a_33379_34007.n107 0.809892
R54632 a_33379_34007.t0 a_33379_34007.n1 0.311051
R54633 a_33379_34007.n176 a_33379_34007.n175 0.752
R54634 a_33379_34007.n146 a_33379_34007.n135 0.752
R54635 a_33379_34007.n256 a_33379_34007.n238 0.752
R54636 a_33379_34007.n294 a_33379_34007.n293 0.752
R54637 a_33379_34007.n235 a_33379_34007.n234 0.71825
R54638 a_33379_34007.n205 a_33379_34007.n195 0.71825
R54639 a_33379_34007.n312 a_33379_34007.n301 0.71825
R54640 a_33379_34007.n348 a_33379_34007.n347 0.71825
R54641 a_33379_34007.n150 a_33379_34007.n149 0.673132
R54642 a_33379_34007.n149 a_33379_34007.n148 0.673132
R54643 a_33379_34007.n127 a_33379_34007.n126 0.673132
R54644 a_33379_34007.n128 a_33379_34007.n127 0.673132
R54645 a_33379_34007.n209 a_33379_34007.n208 0.673132
R54646 a_33379_34007.n208 a_33379_34007.n207 0.673132
R54647 a_33379_34007.n188 a_33379_34007.n187 0.673132
R54648 a_33379_34007.n189 a_33379_34007.n188 0.673132
R54649 a_33379_34007.n282 a_33379_34007.n281 0.673132
R54650 a_33379_34007.n283 a_33379_34007.n282 0.673132
R54651 a_33379_34007.n253 a_33379_34007.n252 0.673132
R54652 a_33379_34007.n254 a_33379_34007.n253 0.673132
R54653 a_33379_34007.n338 a_33379_34007.n337 0.673132
R54654 a_33379_34007.n339 a_33379_34007.n338 0.673132
R54655 a_33379_34007.n316 a_33379_34007.n315 0.673132
R54656 a_33379_34007.n317 a_33379_34007.n316 0.673132
R54657 a_33379_34007.n350 a_33379_34007.n107 0.647527
R54658 a_33379_34007.n55 a_33379_34007.n54 0.321834
R54659 a_33379_34007.n83 a_33379_34007.n82 0.321834
R54660 a_33379_34007.n12 a_33379_34007.n10 0.307602
R54661 a_33379_34007.n21 a_33379_34007.n20 0.307602
R54662 a_33379_34007.n2 a_33379_34007.n141 0.394842
R54663 a_33379_34007.n4 a_33379_34007.n160 0.394842
R54664 a_33379_34007.n7 a_33379_34007.n170 0.394842
R54665 a_33379_34007.n119 a_33379_34007.n11 0.394842
R54666 a_33379_34007.n13 a_33379_34007.n288 0.394842
R54667 a_33379_34007.n274 a_33379_34007.n16 0.394842
R54668 a_33379_34007.n263 a_33379_34007.n262 0.394842
R54669 a_33379_34007.n244 a_33379_34007.n242 0.394842
R54670 a_33379_34007.n22 a_33379_34007.n144 0.381816
R54671 a_33379_34007.n24 a_33379_34007.n5 0.381816
R54672 a_33379_34007.n28 a_33379_34007.n8 0.381816
R54673 a_33379_34007.n31 a_33379_34007.n14 0.381816
R54674 a_33379_34007.n17 a_33379_34007.n270 0.381816
R54675 a_33379_34007.n258 a_33379_34007.n257 0.381816
R54676 a_33379_34007.n202 a_33379_34007.n201 0.379447
R54677 a_33379_34007.n199 a_33379_34007.n198 0.379447
R54678 a_33379_34007.n221 a_33379_34007.n220 0.379447
R54679 a_33379_34007.n216 a_33379_34007.n215 0.379447
R54680 a_33379_34007.n213 a_33379_34007.n212 0.379447
R54681 a_33379_34007.n62 a_33379_34007.n64 0.379447
R54682 a_33379_34007.n65 a_33379_34007.n229 0.379447
R54683 a_33379_34007.n225 a_33379_34007.n224 0.379447
R54684 a_33379_34007.n71 a_33379_34007.n178 0.379447
R54685 a_33379_34007.n183 a_33379_34007.n74 0.379447
R54686 a_33379_34007.n77 a_33379_34007.n79 0.379447
R54687 a_33379_34007.n80 a_33379_34007.n342 0.379447
R54688 a_33379_34007.n84 a_33379_34007.n329 0.379447
R54689 a_33379_34007.n88 a_33379_34007.n85 0.379447
R54690 a_33379_34007.n333 a_33379_34007.n91 0.379447
R54691 a_33379_34007.n95 a_33379_34007.n320 0.379447
R54692 a_33379_34007.n97 a_33379_34007.n323 0.379447
R54693 a_33379_34007.n100 a_33379_34007.n98 0.379447
R54694 a_33379_34007.n103 a_33379_34007.n307 0.379447
R54695 a_33379_34007.n105 a_33379_34007.n310 0.379447
R54696 a_33379_34007.n118 a_33379_34007.n117 0.375125
R54697 a_33379_34007.n169 a_33379_34007.n129 0.375125
R54698 a_33379_34007.n159 a_33379_34007.n132 0.375125
R54699 a_33379_34007.n140 a_33379_34007.n137 0.375125
R54700 a_33379_34007.n245 a_33379_34007.n241 0.375125
R54701 a_33379_34007.n261 a_33379_34007.n113 0.375125
R54702 a_33379_34007.n273 a_33379_34007.n272 0.375125
R54703 a_33379_34007.n287 a_33379_34007.n284 0.375125
R54704 a_33379_34007.n173 a_33379_34007.n172 0.36275
R54705 a_33379_34007.n163 a_33379_34007.n162 0.36275
R54706 a_33379_34007.n143 a_33379_34007.n136 0.36275
R54707 a_33379_34007.n259 a_33379_34007.n114 0.36275
R54708 a_33379_34007.n269 a_33379_34007.n111 0.36275
R54709 a_33379_34007.n291 a_33379_34007.n290 0.36275
R54710 a_33379_34007.n182 a_33379_34007.n181 0.3605
R54711 a_33379_34007.n185 a_33379_34007.n184 0.3605
R54712 a_33379_34007.n232 a_33379_34007.n231 0.3605
R54713 a_33379_34007.n228 a_33379_34007.n190 0.3605
R54714 a_33379_34007.n226 a_33379_34007.n191 0.3605
R54715 a_33379_34007.n219 a_33379_34007.n192 0.3605
R54716 a_33379_34007.n217 a_33379_34007.n193 0.3605
R54717 a_33379_34007.n214 a_33379_34007.n194 0.3605
R54718 a_33379_34007.n203 a_33379_34007.n196 0.3605
R54719 a_33379_34007.n200 a_33379_34007.n197 0.3605
R54720 a_33379_34007.n306 a_33379_34007.n303 0.3605
R54721 a_33379_34007.n309 a_33379_34007.n302 0.3605
R54722 a_33379_34007.n319 a_33379_34007.n300 0.3605
R54723 a_33379_34007.n322 a_33379_34007.n299 0.3605
R54724 a_33379_34007.n326 a_33379_34007.n325 0.3605
R54725 a_33379_34007.n328 a_33379_34007.n297 0.3605
R54726 a_33379_34007.n332 a_33379_34007.n331 0.3605
R54727 a_33379_34007.n335 a_33379_34007.n334 0.3605
R54728 a_33379_34007.n345 a_33379_34007.n344 0.3605
R54729 a_33379_34007.n341 a_33379_34007.n340 0.3605
R54730 a_33379_34007.n139 a_33379_34007.n138 0.348488
R54731 a_33379_34007.n286 a_33379_34007.n285 0.348488
R54732 a_33379_34007.n180 a_33379_34007.n179 0.327481
R54733 a_33379_34007.n305 a_33379_34007.n304 0.327481
R54734 a_33379_34007.n156 a_33379_34007.n155 0.302474
R54735 a_33379_34007.n166 a_33379_34007.n165 0.302474
R54736 a_33379_34007.n122 a_33379_34007.n41 0.302474
R54737 a_33379_34007.n277 a_33379_34007.n44 0.302474
R54738 a_33379_34007.n46 a_33379_34007.n112 0.302474
R54739 a_33379_34007.n49 a_33379_34007.n248 0.302474
R54740 a_33379_34007.n124 a_33379_34007.n123 0.287375
R54741 a_33379_34007.n164 a_33379_34007.n131 0.287375
R54742 a_33379_34007.n154 a_33379_34007.n134 0.287375
R54743 a_33379_34007.n247 a_33379_34007.n239 0.287375
R54744 a_33379_34007.n268 a_33379_34007.n267 0.287375
R54745 a_33379_34007.n279 a_33379_34007.n278 0.287375
R54746 a_33379_34007.n223 a_33379_34007.n192 0.208099
R54747 a_33379_34007.n328 a_33379_34007.n327 0.208099
R54748 a_33379_34007.n101 a_33379_34007.n100 0.152079
R54749 a_33379_34007.n314 a_33379_34007.n106 0.147342
R54750 a_33379_34007.n310 a_33379_34007.n104 0.147342
R54751 a_33379_34007.n23 a_33379_34007.n22 0.147342
R54752 a_33379_34007.n3 a_33379_34007.n2 0.147342
R54753 a_33379_34007.n6 a_33379_34007.n4 0.147342
R54754 a_33379_34007.n157 a_33379_34007.n156 0.147342
R54755 a_33379_34007.n155 a_33379_34007.n37 0.147342
R54756 a_33379_34007.n29 a_33379_34007.n28 0.147342
R54757 a_33379_34007.n9 a_33379_34007.n7 0.147342
R54758 a_33379_34007.n167 a_33379_34007.n166 0.147342
R54759 a_33379_34007.n122 a_33379_34007.n121 0.147342
R54760 a_33379_34007.n42 a_33379_34007.n41 0.147342
R54761 a_33379_34007.n206 a_33379_34007.n51 0.147342
R54762 a_33379_34007.n201 a_33379_34007.n53 0.147342
R54763 a_33379_34007.n220 a_33379_34007.n56 0.147342
R54764 a_33379_34007.n215 a_33379_34007.n58 0.147342
R54765 a_33379_34007.n212 a_33379_34007.n60 0.147342
R54766 a_33379_34007.n233 a_33379_34007.n63 0.147342
R54767 a_33379_34007.n66 a_33379_34007.n64 0.147342
R54768 a_33379_34007.n229 a_33379_34007.n67 0.147342
R54769 a_33379_34007.n72 a_33379_34007.n71 0.147342
R54770 a_33379_34007.n75 a_33379_34007.n74 0.147342
R54771 a_33379_34007.n32 a_33379_34007.n31 0.147342
R54772 a_33379_34007.n15 a_33379_34007.n13 0.147342
R54773 a_33379_34007.n18 a_33379_34007.n16 0.147342
R54774 a_33379_34007.n277 a_33379_34007.n276 0.147342
R54775 a_33379_34007.n45 a_33379_34007.n44 0.147342
R54776 a_33379_34007.n257 a_33379_34007.n36 0.147342
R54777 a_33379_34007.n262 a_33379_34007.n19 0.147342
R54778 a_33379_34007.n265 a_33379_34007.n112 0.147342
R54779 a_33379_34007.n248 a_33379_34007.n240 0.147342
R54780 a_33379_34007.n50 a_33379_34007.n49 0.147342
R54781 a_33379_34007.n346 a_33379_34007.n78 0.147342
R54782 a_33379_34007.n81 a_33379_34007.n79 0.147342
R54783 a_33379_34007.n86 a_33379_34007.n84 0.147342
R54784 a_33379_34007.n89 a_33379_34007.n88 0.147342
R54785 a_33379_34007.n92 a_33379_34007.n91 0.147342
R54786 a_33379_34007.n94 a_33379_34007.n93 0.147342
R54787 a_33379_34007.n96 a_33379_34007.n95 0.147342
R54788 a_33379_34007.n99 a_33379_34007.n97 0.147342
R54789 a_33379_34007.n104 a_33379_34007.n103 0.147342
R54790 a_33379_34007.n106 a_33379_34007.n105 0.147342
R54791 a_33379_34007.n222 a_33379_34007.n221 0.142605
R54792 a_33379_34007.n179 a_33379_34007.n178 0.142605
R54793 a_33379_34007.n329 a_33379_34007.n298 0.142605
R54794 a_33379_34007.n307 a_33379_34007.n304 0.142605
R54795 a_33379_34007.n117 a_33379_34007.n10 1.12843
R54796 a_33379_34007.n118 a_33379_34007.n116 0.14
R54797 a_33379_34007.n123 a_33379_34007.n116 0.14
R54798 a_33379_34007.n40 a_33379_34007.n124 0.14
R54799 a_33379_34007.n40 a_33379_34007.n115 0.14
R54800 a_33379_34007.n175 a_33379_34007.n27 0.14
R54801 a_33379_34007.n173 a_33379_34007.n27 0.14
R54802 a_33379_34007.n172 a_33379_34007.n171 0.14
R54803 a_33379_34007.n171 a_33379_34007.n129 0.14
R54804 a_33379_34007.n169 a_33379_34007.n168 0.14
R54805 a_33379_34007.n168 a_33379_34007.n131 0.14
R54806 a_33379_34007.n164 a_33379_34007.n39 0.208307
R54807 a_33379_34007.n39 a_33379_34007.n26 3.16466
R54808 a_33379_34007.n163 a_33379_34007.n26 0.208324
R54809 a_33379_34007.n162 a_33379_34007.n161 0.14
R54810 a_33379_34007.n161 a_33379_34007.n132 0.14
R54811 a_33379_34007.n159 a_33379_34007.n158 0.14
R54812 a_33379_34007.n158 a_33379_34007.n134 0.14
R54813 a_33379_34007.n154 a_33379_34007.n153 0.14
R54814 a_33379_34007.n153 a_33379_34007.n152 0.14
R54815 a_33379_34007.n146 a_33379_34007.n145 0.14
R54816 a_33379_34007.n145 a_33379_34007.n136 0.14
R54817 a_33379_34007.n143 a_33379_34007.n142 0.14
R54818 a_33379_34007.n142 a_33379_34007.n137 0.14
R54819 a_33379_34007.n182 a_33379_34007.n70 0.14
R54820 a_33379_34007.n184 a_33379_34007.n70 0.14
R54821 a_33379_34007.n73 a_33379_34007.n185 0.14
R54822 a_33379_34007.n73 a_33379_34007.n177 0.14
R54823 a_33379_34007.n234 a_33379_34007.n61 0.14
R54824 a_33379_34007.n232 a_33379_34007.n61 0.14
R54825 a_33379_34007.n231 a_33379_34007.n230 0.14
R54826 a_33379_34007.n230 a_33379_34007.n190 0.14
R54827 a_33379_34007.n228 a_33379_34007.n227 0.14
R54828 a_33379_34007.n227 a_33379_34007.n226 0.14
R54829 a_33379_34007.n69 a_33379_34007.n191 0.208134
R54830 a_33379_34007.n69 a_33379_34007.n223 3.10882
R54831 a_33379_34007.n219 a_33379_34007.n218 0.14
R54832 a_33379_34007.n218 a_33379_34007.n217 0.14
R54833 a_33379_34007.n57 a_33379_34007.n193 0.14
R54834 a_33379_34007.n57 a_33379_34007.n214 0.14
R54835 a_33379_34007.n59 a_33379_34007.n194 0.14
R54836 a_33379_34007.n59 a_33379_34007.n211 0.14
R54837 a_33379_34007.n205 a_33379_34007.n204 0.14
R54838 a_33379_34007.n204 a_33379_34007.n203 0.14
R54839 a_33379_34007.n52 a_33379_34007.n196 0.14
R54840 a_33379_34007.n52 a_33379_34007.n200 0.14
R54841 a_33379_34007.n55 a_33379_34007.n197 1.12757
R54842 a_33379_34007.n21 a_33379_34007.n241 1.12843
R54843 a_33379_34007.n246 a_33379_34007.n245 0.14
R54844 a_33379_34007.n247 a_33379_34007.n246 0.14
R54845 a_33379_34007.n249 a_33379_34007.n239 0.14
R54846 a_33379_34007.n250 a_33379_34007.n249 0.14
R54847 a_33379_34007.n35 a_33379_34007.n256 0.14
R54848 a_33379_34007.n35 a_33379_34007.n114 0.14
R54849 a_33379_34007.n260 a_33379_34007.n259 0.14
R54850 a_33379_34007.n261 a_33379_34007.n260 0.14
R54851 a_33379_34007.n266 a_33379_34007.n113 0.14
R54852 a_33379_34007.n267 a_33379_34007.n266 0.14
R54853 a_33379_34007.n268 a_33379_34007.n48 0.208307
R54854 a_33379_34007.n34 a_33379_34007.n48 3.16466
R54855 a_33379_34007.n269 a_33379_34007.n34 0.208324
R54856 a_33379_34007.n271 a_33379_34007.n111 0.14
R54857 a_33379_34007.n272 a_33379_34007.n271 0.14
R54858 a_33379_34007.n273 a_33379_34007.n110 0.14
R54859 a_33379_34007.n278 a_33379_34007.n110 0.14
R54860 a_33379_34007.n43 a_33379_34007.n279 0.14
R54861 a_33379_34007.n43 a_33379_34007.n109 0.14
R54862 a_33379_34007.n293 a_33379_34007.n30 0.14
R54863 a_33379_34007.n291 a_33379_34007.n30 0.14
R54864 a_33379_34007.n290 a_33379_34007.n289 0.14
R54865 a_33379_34007.n289 a_33379_34007.n284 0.14
R54866 a_33379_34007.n308 a_33379_34007.n303 0.14
R54867 a_33379_34007.n309 a_33379_34007.n308 0.14
R54868 a_33379_34007.n311 a_33379_34007.n302 0.14
R54869 a_33379_34007.n313 a_33379_34007.n311 0.14
R54870 a_33379_34007.n318 a_33379_34007.n301 0.14
R54871 a_33379_34007.n319 a_33379_34007.n318 0.14
R54872 a_33379_34007.n321 a_33379_34007.n300 0.14
R54873 a_33379_34007.n322 a_33379_34007.n321 0.14
R54874 a_33379_34007.n324 a_33379_34007.n299 0.14
R54875 a_33379_34007.n325 a_33379_34007.n324 0.14
R54876 a_33379_34007.n326 a_33379_34007.n102 0.208134
R54877 a_33379_34007.n327 a_33379_34007.n102 3.10882
R54878 a_33379_34007.n342 a_33379_34007.n82 0.152079
R54879 a_33379_34007.n99 a_33379_34007.n98 0.147342
R54880 a_33379_34007.n323 a_33379_34007.n96 0.147342
R54881 a_33379_34007.n320 a_33379_34007.n94 0.147342
R54882 a_33379_34007.n336 a_33379_34007.n92 0.147342
R54883 a_33379_34007.n333 a_33379_34007.n89 0.147342
R54884 a_33379_34007.n86 a_33379_34007.n85 0.147342
R54885 a_33379_34007.n330 a_33379_34007.n297 0.14
R54886 a_33379_34007.n331 a_33379_34007.n330 0.14
R54887 a_33379_34007.n332 a_33379_34007.n87 0.14
R54888 a_33379_34007.n334 a_33379_34007.n87 0.14
R54889 a_33379_34007.n90 a_33379_34007.n335 0.14
R54890 a_33379_34007.n90 a_33379_34007.n296 0.14
R54891 a_33379_34007.n347 a_33379_34007.n76 0.14
R54892 a_33379_34007.n345 a_33379_34007.n76 0.14
R54893 a_33379_34007.n344 a_33379_34007.n343 0.14
R54894 a_33379_34007.n343 a_33379_34007.n340 0.14
R54895 a_33379_34007.n341 a_33379_34007.n83 1.12757
R54896 a_33379_34007.n242 a_33379_34007.n20 0.1805
R54897 a_33379_34007.n12 a_33379_34007.n11 0.1805
R54898 a_33379_34007.n270 a_33379_34007.n33 0.178132
R54899 a_33379_34007.n25 a_33379_34007.n24 0.178132
R54900 a_33379_34007.n47 a_33379_34007.n46 0.175763
R54901 a_33379_34007.n165 a_33379_34007.n38 0.175763
R54902 a_33379_34007.n224 a_33379_34007.n68 0.152079
R54903 a_33379_34007.n198 a_33379_34007.n54 0.152079
R54904 a_33379_34007.n81 a_33379_34007.n80 0.147342
R54905 a_33379_34007.n78 a_33379_34007.n77 0.147342
R54906 a_33379_34007.n186 a_33379_34007.n75 0.147342
R54907 a_33379_34007.n183 a_33379_34007.n72 0.147342
R54908 a_33379_34007.n225 a_33379_34007.n67 0.147342
R54909 a_33379_34007.n66 a_33379_34007.n65 0.147342
R54910 a_33379_34007.n63 a_33379_34007.n62 0.147342
R54911 a_33379_34007.n210 a_33379_34007.n60 0.147342
R54912 a_33379_34007.n213 a_33379_34007.n58 0.147342
R54913 a_33379_34007.n216 a_33379_34007.n56 0.147342
R54914 a_33379_34007.n199 a_33379_34007.n53 0.147342
R54915 a_33379_34007.n202 a_33379_34007.n51 0.147342
R54916 a_33379_34007.n251 a_33379_34007.n50 0.147342
R54917 a_33379_34007.n280 a_33379_34007.n45 0.147342
R54918 a_33379_34007.n125 a_33379_34007.n42 0.147342
R54919 a_33379_34007.n151 a_33379_34007.n37 0.147342
R54920 a_33379_34007.n255 a_33379_34007.n36 0.147342
R54921 a_33379_34007.n292 a_33379_34007.n32 0.147342
R54922 a_33379_34007.n174 a_33379_34007.n29 0.147342
R54923 a_33379_34007.n147 a_33379_34007.n23 0.147342
R54924 a_33379_34007.n258 a_33379_34007.n19 0.147342
R54925 a_33379_34007.n18 a_33379_34007.n17 0.147342
R54926 a_33379_34007.n15 a_33379_34007.n14 0.147342
R54927 a_33379_34007.n9 a_33379_34007.n8 0.147342
R54928 a_33379_34007.n6 a_33379_34007.n5 0.147342
R54929 a_33379_34007.n144 a_33379_34007.n3 0.147342
R54930 a_33379_34007.n141 a_33379_34007.n138 0.0987895
R54931 a_33379_34007.n160 a_33379_34007.n133 0.0987895
R54932 a_33379_34007.n170 a_33379_34007.n130 0.0987895
R54933 a_33379_34007.n120 a_33379_34007.n119 0.0987895
R54934 a_33379_34007.n288 a_33379_34007.n285 0.0987895
R54935 a_33379_34007.n275 a_33379_34007.n274 0.0987895
R54936 a_33379_34007.n264 a_33379_34007.n263 0.0987895
R54937 a_33379_34007.n244 a_33379_34007.n243 0.0987895
R54938 a_33379_34007.n157 a_33379_34007.n133 0.0490526
R54939 a_33379_34007.n167 a_33379_34007.n130 0.0490526
R54940 a_33379_34007.n121 a_33379_34007.n120 0.0490526
R54941 a_33379_34007.n276 a_33379_34007.n275 0.0490526
R54942 a_33379_34007.n265 a_33379_34007.n264 0.0490526
R54943 a_33379_34007.n243 a_33379_34007.n240 0.0490526
R54944 a_33379_34007.n0 a_33379_34007.t1 0.295568
R54945 a_33379_34007.n0 a_33379_34007.n351 16.9974
R54946 a_33249_34067.n114 a_33249_34067.n113 8.18538
R54947 a_33249_34067.n125 a_33249_34067.n123 7.22198
R54948 a_33249_34067.n153 a_33249_34067.n28 7.22198
R54949 a_33249_34067.n30 a_33249_34067.t23 6.77653
R54950 a_33249_34067.n132 a_33249_34067.t20 6.77653
R54951 a_33249_34067.n48 a_33249_34067.t77 6.7761
R54952 a_33249_34067.n145 a_33249_34067.t74 6.7761
R54953 a_33249_34067.n25 a_33249_34067.t133 6.86989
R54954 a_33249_34067.n9 a_33249_34067.t101 6.77231
R54955 a_33249_34067.n19 a_33249_34067.t89 6.77231
R54956 a_33249_34067.n109 a_33249_34067.t7 6.53862
R54957 a_33249_34067.n114 a_33249_34067.n55 5.95467
R54958 a_33249_34067.n79 a_33249_34067.n77 5.89898
R54959 a_33249_34067.n93 a_33249_34067.t126 5.66511
R54960 a_33249_34067.n86 a_33249_34067.t111 5.66511
R54961 a_33249_34067.n94 a_33249_34067.t131 5.66379
R54962 a_33249_34067.n87 a_33249_34067.t116 5.66379
R54963 a_33249_34067.n86 a_33249_34067.n85 5.65285
R54964 a_33249_34067.n73 a_33249_34067.t130 5.61877
R54965 a_33249_34067.n74 a_33249_34067.t109 5.61877
R54966 a_33249_34067.n70 a_33249_34067.t114 5.61877
R54967 a_33249_34067.n45 a_33249_34067.t65 5.50607
R54968 a_33249_34067.n31 a_33249_34067.t36 5.50607
R54969 a_33249_34067.n142 a_33249_34067.t59 5.50607
R54970 a_33249_34067.n133 a_33249_34067.t31 5.50607
R54971 a_33249_34067.n46 a_33249_34067.t97 5.50475
R54972 a_33249_34067.n42 a_33249_34067.t62 5.50475
R54973 a_33249_34067.n41 a_33249_34067.t72 5.50475
R54974 a_33249_34067.n32 a_33249_34067.t69 5.50475
R54975 a_33249_34067.n143 a_33249_34067.t92 5.50475
R54976 a_33249_34067.n139 a_33249_34067.t56 5.50475
R54977 a_33249_34067.n138 a_33249_34067.t68 5.50475
R54978 a_33249_34067.n134 a_33249_34067.t64 5.50475
R54979 a_33249_34067.n112 a_33249_34067.t1 5.28484
R54980 a_33249_34067.n22 a_33249_34067.n99 5.29079
R54981 a_33249_34067.n96 a_33249_34067.n95 4.88835
R54982 a_33249_34067.n63 a_33249_34067.n62 4.88517
R54983 a_33249_34067.n100 a_33249_34067.n21 4.02009
R54984 a_33249_34067.t11 a_33249_34067.n20 5.28011
R54985 a_33249_34067.t10 a_33249_34067.n22 5.28011
R54986 a_33249_34067.n0 a_33249_34067.n38 4.0312
R54987 a_33249_34067.n1 a_33249_34067.t84 5.5012
R54988 a_33249_34067.n2 a_33249_34067.t54 5.5012
R54989 a_33249_34067.n3 a_33249_34067.n37 4.0312
R54990 a_33249_34067.n4 a_33249_34067.t50 5.5012
R54991 a_33249_34067.n5 a_33249_34067.t61 5.5012
R54992 a_33249_34067.n6 a_33249_34067.n36 4.0312
R54993 a_33249_34067.t57 a_33249_34067.n7 5.5012
R54994 a_33249_34067.t26 a_33249_34067.n8 5.5012
R54995 a_33249_34067.n35 a_33249_34067.n9 4.0312
R54996 a_33249_34067.n10 a_33249_34067.n118 4.0312
R54997 a_33249_34067.n11 a_33249_34067.t79 5.5012
R54998 a_33249_34067.n12 a_33249_34067.t45 5.5012
R54999 a_33249_34067.n13 a_33249_34067.n117 4.0312
R55000 a_33249_34067.n14 a_33249_34067.t39 5.5012
R55001 a_33249_34067.n15 a_33249_34067.t51 5.5012
R55002 a_33249_34067.n16 a_33249_34067.n116 4.0312
R55003 a_33249_34067.t48 a_33249_34067.n17 5.5012
R55004 a_33249_34067.t18 a_33249_34067.n18 5.5012
R55005 a_33249_34067.n115 a_33249_34067.n19 4.0312
R55006 a_33249_34067.n23 a_33249_34067.n72 4.40099
R55007 a_33249_34067.n24 a_33249_34067.n71 4.40099
R55008 a_33249_34067.n69 a_33249_34067.n25 4.40099
R55009 a_33249_34067.n92 a_33249_34067.n91 4.40379
R55010 a_33249_34067.n90 a_33249_34067.n89 4.40379
R55011 a_33249_34067.n78 a_33249_34067.t136 4.40142
R55012 a_33249_34067.n64 a_33249_34067.t125 4.40142
R55013 a_33249_34067.n27 a_33249_34067.t52 4.24002
R55014 a_33249_34067.n26 a_33249_34067.t43 4.24002
R55015 a_33249_34067.n124 a_33249_34067.t41 4.24002
R55016 a_33249_34067.n56 a_33249_34067.t35 4.24002
R55017 a_33249_34067.n105 a_33249_34067.t3 4.22616
R55018 a_33249_34067.n48 a_33249_34067.n47 4.03475
R55019 a_33249_34067.n44 a_33249_34067.n43 4.03475
R55020 a_33249_34067.n40 a_33249_34067.n39 4.03475
R55021 a_33249_34067.n30 a_33249_34067.n29 4.03475
R55022 a_33249_34067.n145 a_33249_34067.n144 4.03475
R55023 a_33249_34067.n141 a_33249_34067.n140 4.03475
R55024 a_33249_34067.n137 a_33249_34067.n136 4.03475
R55025 a_33249_34067.n132 a_33249_34067.n131 4.03475
R55026 a_33249_34067.n111 a_33249_34067.n110 4.02484
R55027 a_33249_34067.n109 a_33249_34067.n108 4.02484
R55028 a_33249_34067.n105 a_33249_34067.t9 4.02247
R55029 a_33249_34067.n107 a_33249_34067.n106 3.96014
R55030 a_33249_34067.n98 a_33249_34067.n61 3.94195
R55031 a_33249_34067.n78 a_33249_34067.t141 3.84721
R55032 a_33249_34067.n64 a_33249_34067.t129 3.84721
R55033 a_33249_34067.n92 a_33249_34067.n90 3.81703
R55034 a_33249_34067.n111 a_33249_34067.n109 3.80578
R55035 a_33249_34067.n27 a_33249_34067.t47 3.68818
R55036 a_33249_34067.n26 a_33249_34067.t38 3.68818
R55037 a_33249_34067.n124 a_33249_34067.t40 3.68818
R55038 a_33249_34067.n56 a_33249_34067.t34 3.68818
R55039 a_33249_34067.n130 a_33249_34067.n129 3.23904
R55040 a_33249_34067.n54 a_33249_34067.n53 3.23904
R55041 a_33249_34067.n84 a_33249_34067.n83 3.23004
R55042 a_33249_34067.n82 a_33249_34067.n81 3.14142
R55043 a_33249_34067.n67 a_33249_34067.n66 3.14142
R55044 a_33249_34067.n104 a_33249_34067.n102 2.96616
R55045 a_33249_34067.n52 a_33249_34067.n51 2.77002
R55046 a_33249_34067.n128 a_33249_34067.n127 2.77002
R55047 a_33249_34067.n59 a_33249_34067.n58 2.77002
R55048 a_33249_34067.n157 a_33249_34067.n156 2.77002
R55049 a_33249_34067.n104 a_33249_34067.n103 2.76247
R55050 a_33249_34067.n154 a_33249_34067.n26 2.7375
R55051 a_33249_34067.n60 a_33249_34067.n56 2.73714
R55052 a_33249_34067.n106 a_33249_34067.n104 2.71914
R55053 a_33249_34067.n68 a_33249_34067.n64 2.71914
R55054 a_33249_34067.n98 a_33249_34067.n97 2.64424
R55055 a_33249_34067.n42 a_33249_34067.n41 2.60203
R55056 a_33249_34067.n139 a_33249_34067.n138 2.60203
R55057 a_33249_34067.n82 a_33249_34067.n80 2.58721
R55058 a_33249_34067.n67 a_33249_34067.n65 2.58721
R55059 a_33249_34067.n87 a_33249_34067.n86 2.55136
R55060 a_33249_34067.n94 a_33249_34067.n93 2.55136
R55061 a_33249_34067.n32 a_33249_34067.n31 2.52436
R55062 a_33249_34067.n46 a_33249_34067.n45 2.52436
R55063 a_33249_34067.n134 a_33249_34067.n133 2.52436
R55064 a_33249_34067.n143 a_33249_34067.n142 2.52436
R55065 a_33249_34067.n76 a_33249_34067.n75 2.2807
R55066 a_33249_34067.n84 a_33249_34067.n63 2.2807
R55067 a_33249_34067.n52 a_33249_34067.n50 2.21818
R55068 a_33249_34067.n128 a_33249_34067.n126 2.21818
R55069 a_33249_34067.n59 a_33249_34067.n57 2.21818
R55070 a_33249_34067.n156 a_33249_34067.n155 2.21818
R55071 a_33249_34067.n152 a_33249_34067.n33 2.13841
R55072 a_33249_34067.n54 a_33249_34067.n49 2.13841
R55073 a_33249_34067.n123 a_33249_34067.n60 1.73904
R55074 a_33249_34067.n154 a_33249_34067.n153 1.73868
R55075 a_33249_34067.n113 a_33249_34067.n112 1.73609
R55076 a_33249_34067.n77 a_33249_34067.n68 1.73004
R55077 a_33249_34067.n121 a_33249_34067.n120 1.5005
R55078 a_33249_34067.n123 a_33249_34067.n122 1.5005
R55079 a_33249_34067.n135 a_33249_34067.n34 1.5005
R55080 a_33249_34067.n151 a_33249_34067.n150 1.5005
R55081 a_33249_34067.n77 a_33249_34067.n76 1.5005
R55082 a_33249_34067.n88 a_33249_34067.n61 1.5005
R55083 a_33249_34067.n97 a_33249_34067.n96 1.5005
R55084 a_33249_34067.n119 a_33249_34067.n55 1.5005
R55085 a_33249_34067.n147 a_33249_34067.n146 1.5005
R55086 a_33249_34067.n149 a_33249_34067.n148 1.5005
R55087 a_33249_34067.n153 a_33249_34067.n152 1.5005
R55088 a_33249_34067.n155 a_33249_34067.t98 1.4705
R55089 a_33249_34067.n155 a_33249_34067.t49 1.4705
R55090 a_33249_34067.n50 a_33249_34067.t19 1.4705
R55091 a_33249_34067.n50 a_33249_34067.t71 1.4705
R55092 a_33249_34067.n51 a_33249_34067.t24 1.4705
R55093 a_33249_34067.n51 a_33249_34067.t76 1.4705
R55094 a_33249_34067.n47 a_33249_34067.t37 1.4705
R55095 a_33249_34067.n47 a_33249_34067.t96 1.4705
R55096 a_33249_34067.n43 a_33249_34067.t32 1.4705
R55097 a_33249_34067.n43 a_33249_34067.t90 1.4705
R55098 a_33249_34067.n39 a_33249_34067.t30 1.4705
R55099 a_33249_34067.n39 a_33249_34067.t99 1.4705
R55100 a_33249_34067.n29 a_33249_34067.t88 1.4705
R55101 a_33249_34067.n29 a_33249_34067.t63 1.4705
R55102 a_33249_34067.n38 a_33249_34067.t28 1.4705
R55103 a_33249_34067.n38 a_33249_34067.t83 1.4705
R55104 a_33249_34067.n37 a_33249_34067.t25 1.4705
R55105 a_33249_34067.n37 a_33249_34067.t82 1.4705
R55106 a_33249_34067.n36 a_33249_34067.t22 1.4705
R55107 a_33249_34067.n36 a_33249_34067.t87 1.4705
R55108 a_33249_34067.n35 a_33249_34067.t81 1.4705
R55109 a_33249_34067.n35 a_33249_34067.t53 1.4705
R55110 a_33249_34067.n144 a_33249_34067.t33 1.4705
R55111 a_33249_34067.n144 a_33249_34067.t91 1.4705
R55112 a_33249_34067.n140 a_33249_34067.t29 1.4705
R55113 a_33249_34067.n140 a_33249_34067.t86 1.4705
R55114 a_33249_34067.n136 a_33249_34067.t27 1.4705
R55115 a_33249_34067.n136 a_33249_34067.t95 1.4705
R55116 a_33249_34067.n131 a_33249_34067.t85 1.4705
R55117 a_33249_34067.n131 a_33249_34067.t58 1.4705
R55118 a_33249_34067.n126 a_33249_34067.t102 1.4705
R55119 a_33249_34067.n126 a_33249_34067.t66 1.4705
R55120 a_33249_34067.n127 a_33249_34067.t103 1.4705
R55121 a_33249_34067.n127 a_33249_34067.t67 1.4705
R55122 a_33249_34067.n57 a_33249_34067.t93 1.4705
R55123 a_33249_34067.n57 a_33249_34067.t44 1.4705
R55124 a_33249_34067.n58 a_33249_34067.t94 1.4705
R55125 a_33249_34067.n58 a_33249_34067.t46 1.4705
R55126 a_33249_34067.n118 a_33249_34067.t21 1.4705
R55127 a_33249_34067.n118 a_33249_34067.t78 1.4705
R55128 a_33249_34067.n117 a_33249_34067.t104 1.4705
R55129 a_33249_34067.n117 a_33249_34067.t75 1.4705
R55130 a_33249_34067.n116 a_33249_34067.t100 1.4705
R55131 a_33249_34067.n116 a_33249_34067.t80 1.4705
R55132 a_33249_34067.n115 a_33249_34067.t73 1.4705
R55133 a_33249_34067.n115 a_33249_34067.t42 1.4705
R55134 a_33249_34067.t105 a_33249_34067.n157 1.4705
R55135 a_33249_34067.n157 a_33249_34067.t55 1.4705
R55136 a_33249_34067.n53 a_33249_34067.n52 1.46537
R55137 a_33249_34067.n28 a_33249_34067.n27 1.46537
R55138 a_33249_34067.n129 a_33249_34067.n128 1.46537
R55139 a_33249_34067.n125 a_33249_34067.n124 1.46537
R55140 a_33249_34067.n60 a_33249_34067.n59 1.46537
R55141 a_33249_34067.n83 a_33249_34067.n82 1.46537
R55142 a_33249_34067.n79 a_33249_34067.n78 1.46537
R55143 a_33249_34067.n68 a_33249_34067.n67 1.46537
R55144 a_33249_34067.n156 a_33249_34067.n154 1.46537
R55145 a_33249_34067.n106 a_33249_34067.n105 1.46537
R55146 a_33249_34067.n121 a_33249_34067.n114 1.37875
R55147 a_33249_34067.n41 a_33249_34067.n40 1.27228
R55148 a_33249_34067.n44 a_33249_34067.n42 1.27228
R55149 a_33249_34067.n138 a_33249_34067.n137 1.27228
R55150 a_33249_34067.n141 a_33249_34067.n139 1.27228
R55151 a_33249_34067.n129 a_33249_34067.n125 1.27228
R55152 a_33249_34067.n53 a_33249_34067.n28 1.27228
R55153 a_33249_34067.n31 a_33249_34067.n30 1.26756
R55154 a_33249_34067.n45 a_33249_34067.n44 1.26756
R55155 a_33249_34067.n133 a_33249_34067.n132 1.26756
R55156 a_33249_34067.n142 a_33249_34067.n141 1.26756
R55157 a_33249_34067.n101 a_33249_34067.n98 1.26344
R55158 a_33249_34067.n110 a_33249_34067.t15 1.2605
R55159 a_33249_34067.n110 a_33249_34067.t14 1.2605
R55160 a_33249_34067.n108 a_33249_34067.t12 1.2605
R55161 a_33249_34067.n108 a_33249_34067.t0 1.2605
R55162 a_33249_34067.n100 a_33249_34067.t6 1.2605
R55163 a_33249_34067.n100 a_33249_34067.t5 1.2605
R55164 a_33249_34067.n99 a_33249_34067.t17 1.2605
R55165 a_33249_34067.n99 a_33249_34067.t4 1.2605
R55166 a_33249_34067.n102 a_33249_34067.t8 1.2605
R55167 a_33249_34067.n102 a_33249_34067.t13 1.2605
R55168 a_33249_34067.n103 a_33249_34067.t16 1.2605
R55169 a_33249_34067.n103 a_33249_34067.t2 1.2605
R55170 a_33249_34067.n62 a_33249_34067.t106 1.2605
R55171 a_33249_34067.n62 a_33249_34067.t120 1.2605
R55172 a_33249_34067.n72 a_33249_34067.t118 1.2605
R55173 a_33249_34067.n72 a_33249_34067.t122 1.2605
R55174 a_33249_34067.n71 a_33249_34067.t123 1.2605
R55175 a_33249_34067.n71 a_33249_34067.t135 1.2605
R55176 a_33249_34067.n69 a_33249_34067.t110 1.2605
R55177 a_33249_34067.n69 a_33249_34067.t108 1.2605
R55178 a_33249_34067.n95 a_33249_34067.t107 1.2605
R55179 a_33249_34067.n95 a_33249_34067.t124 1.2605
R55180 a_33249_34067.n91 a_33249_34067.t112 1.2605
R55181 a_33249_34067.n91 a_33249_34067.t119 1.2605
R55182 a_33249_34067.n89 a_33249_34067.t127 1.2605
R55183 a_33249_34067.n89 a_33249_34067.t138 1.2605
R55184 a_33249_34067.n85 a_33249_34067.t137 1.2605
R55185 a_33249_34067.n85 a_33249_34067.t113 1.2605
R55186 a_33249_34067.n80 a_33249_34067.t139 1.2605
R55187 a_33249_34067.n80 a_33249_34067.t117 1.2605
R55188 a_33249_34067.n81 a_33249_34067.t132 1.2605
R55189 a_33249_34067.n81 a_33249_34067.t115 1.2605
R55190 a_33249_34067.n65 a_33249_34067.t128 1.2605
R55191 a_33249_34067.n65 a_33249_34067.t140 1.2605
R55192 a_33249_34067.n66 a_33249_34067.t121 1.2605
R55193 a_33249_34067.n66 a_33249_34067.t134 1.2605
R55194 a_33249_34067.n83 a_33249_34067.n79 1.25428
R55195 a_33249_34067.n112 a_33249_34067.n111 1.25428
R55196 a_33249_34067.n93 a_33249_34067.n92 1.24956
R55197 a_33249_34067.n74 a_33249_34067.n23 1.25162
R55198 a_33249_34067.n33 a_33249_34067.n32 0.796291
R55199 a_33249_34067.n49 a_33249_34067.n46 0.796291
R55200 a_33249_34067.n135 a_33249_34067.n134 0.796291
R55201 a_33249_34067.n146 a_33249_34067.n143 0.796291
R55202 a_33249_34067.n152 a_33249_34067.n151 0.780703
R55203 a_33249_34067.n122 a_33249_34067.n121 0.780703
R55204 a_33249_34067.n148 a_33249_34067.n54 0.780703
R55205 a_33249_34067.n130 a_33249_34067.n55 0.780703
R55206 a_33249_34067.n88 a_33249_34067.n87 0.769291
R55207 a_33249_34067.n96 a_33249_34067.n94 0.769291
R55208 a_33249_34067.n75 a_33249_34067.n70 0.767125
R55209 a_33249_34067.n73 a_33249_34067.n63 0.767125
R55210 a_33249_34067.n113 a_33249_34067.n107 0.639318
R55211 a_33249_34067.n122 a_33249_34067.n34 0.638405
R55212 a_33249_34067.n76 a_33249_34067.n61 0.638405
R55213 a_33249_34067.n97 a_33249_34067.n84 0.638405
R55214 a_33249_34067.n147 a_33249_34067.n130 0.638405
R55215 a_33249_34067.n151 a_33249_34067.n34 0.628372
R55216 a_33249_34067.n148 a_33249_34067.n147 0.628372
R55217 a_33249_34067.n107 a_33249_34067.n101 0.585196
R55218 a_33249_34067.n90 a_33249_34067.n88 0.485484
R55219 a_33249_34067.n40 a_33249_34067.n33 0.476484
R55220 a_33249_34067.n49 a_33249_34067.n48 0.476484
R55221 a_33249_34067.n137 a_33249_34067.n135 0.476484
R55222 a_33249_34067.n146 a_33249_34067.n145 0.476484
R55223 a_33249_34067.n75 a_33249_34067.n24 0.484998
R55224 a_33249_34067.n150 a_33249_34067.n6 0.478684
R55225 a_33249_34067.n149 a_33249_34067.n0 0.478684
R55226 a_33249_34067.n120 a_33249_34067.n16 0.478684
R55227 a_33249_34067.n119 a_33249_34067.n10 0.478684
R55228 a_33249_34067.n8 a_33249_34067.n9 1.27228
R55229 a_33249_34067.n7 a_33249_34067.n8 2.51878
R55230 a_33249_34067.n150 a_33249_34067.n7 0.794091
R55231 a_33249_34067.n5 a_33249_34067.n6 1.27228
R55232 a_33249_34067.n4 a_33249_34067.n5 2.60203
R55233 a_33249_34067.n3 a_33249_34067.n4 1.27228
R55234 a_33249_34067.n2 a_33249_34067.n3 1.27228
R55235 a_33249_34067.n1 a_33249_34067.n2 2.51878
R55236 a_33249_34067.n149 a_33249_34067.n1 0.794091
R55237 a_33249_34067.t70 a_33249_34067.n0 6.77266
R55238 a_33249_34067.n18 a_33249_34067.n19 1.27228
R55239 a_33249_34067.n17 a_33249_34067.n18 2.51878
R55240 a_33249_34067.n120 a_33249_34067.n17 0.794091
R55241 a_33249_34067.n15 a_33249_34067.n16 1.27228
R55242 a_33249_34067.n14 a_33249_34067.n15 2.60203
R55243 a_33249_34067.n13 a_33249_34067.n14 1.27228
R55244 a_33249_34067.n12 a_33249_34067.n13 1.27228
R55245 a_33249_34067.n11 a_33249_34067.n12 2.51878
R55246 a_33249_34067.n119 a_33249_34067.n11 0.794091
R55247 a_33249_34067.t60 a_33249_34067.n10 6.77266
R55248 a_33249_34067.n21 a_33249_34067.n22 3.15817
R55249 a_33249_34067.n20 a_33249_34067.n21 1.27188
R55250 a_33249_34067.n101 a_33249_34067.n20 1.73829
R55251 a_33249_34067.n70 a_33249_34067.n25 3.17898
R55252 a_33249_34067.n74 a_33249_34067.n24 3.19023
R55253 a_33249_34067.n73 a_33249_34067.n23 3.17898
R55254 a_65486_n35156.t8 a_65486_n35156.t5 12.7136
R55255 a_65486_n35156.t8 a_65486_n35156.t14 10.2828
R55256 a_65486_n35156.t8 a_65486_n35156.t0 10.2828
R55257 a_65486_n35156.t8 a_65486_n35156.t13 10.2828
R55258 a_65486_n35156.t8 a_65486_n35156.t2 10.2828
R55259 a_65486_n35156.t8 a_65486_n35156.t6 10.1333
R55260 a_65486_n35156.t8 a_65486_n35156.t21 10.1333
R55261 a_65486_n35156.t8 a_65486_n35156.t4 10.1333
R55262 a_65486_n35156.t8 a_65486_n35156.t22 10.1333
R55263 a_65486_n35156.t8 a_65486_n35156.t11 9.72545
R55264 a_65486_n35156.t8 a_65486_n35156.t20 9.57156
R55265 a_65486_n35156.t8 a_65486_n35156.t17 9.57156
R55266 a_65486_n35156.t8 a_65486_n35156.t19 9.57156
R55267 a_65486_n35156.t8 a_65486_n35156.t18 9.57156
R55268 a_65486_n35156.t8 a_65486_n35156.t16 9.57156
R55269 a_65486_n35156.t8 a_65486_n35156.t23 9.57156
R55270 a_65486_n35156.t8 a_65486_n35156.t15 9.57156
R55271 a_65486_n35156.t8 a_65486_n35156.t12 9.57156
R55272 a_65486_n35156.t11 a_65486_n35156.t10 8.02827
R55273 a_65486_n35156.t8 a_65486_n35156.t9 8.0259
R55274 a_65486_n35156.t8 a_65486_n35156.t3 7.90799
R55275 a_65486_n35156.t1 a_65486_n35156.t8 7.90799
R55276 a_65486_n35156.t8 a_65486_n35156.t7 7.41865
R55277 a_100820_n36322.n0 a_100820_n36322.t16 13.7934
R55278 a_100820_n36322.n2 a_100820_n36322.t1 10.7024
R55279 a_100820_n36322.n2 a_100820_n36322.t7 10.1668
R55280 a_100820_n36322.n2 a_100820_n36322.t5 9.64458
R55281 a_100820_n36322.n2 a_100820_n36322.t3 9.27635
R55282 a_100820_n36322.n2 a_100820_n36322.n0 8.75198
R55283 a_100820_n36322.n0 a_100820_n36322.t20 8.14051
R55284 a_100820_n36322.n0 a_100820_n36322.t18 8.14051
R55285 a_100820_n36322.n0 a_100820_n36322.t10 8.14051
R55286 a_100820_n36322.n0 a_100820_n36322.t11 8.14051
R55287 a_100820_n36322.n0 a_100820_n36322.t17 8.06917
R55288 a_100820_n36322.n0 a_100820_n36322.t15 8.06917
R55289 a_100820_n36322.n0 a_100820_n36322.t14 8.06917
R55290 a_100820_n36322.n0 a_100820_n36322.t9 8.06917
R55291 a_100820_n36322.n0 a_100820_n36322.t23 8.06917
R55292 a_100820_n36322.n0 a_100820_n36322.t19 8.06917
R55293 a_100820_n36322.n0 a_100820_n36322.t22 8.06917
R55294 a_100820_n36322.n1 a_100820_n36322.t4 7.94157
R55295 a_100820_n36322.t0 a_100820_n36322.n2 7.72643
R55296 a_100820_n36322.n1 a_100820_n36322.t6 7.22925
R55297 a_100820_n36322.n2 a_100820_n36322.t2 7.17912
R55298 a_100820_n36322.n0 a_100820_n36322.t8 8.33554
R55299 a_100820_n36322.t21 a_100820_n36322.n0 8.33554
R55300 a_100820_n36322.n0 a_100820_n36322.t12 8.33647
R55301 a_100820_n36322.t13 a_100820_n36322.n0 8.33647
R55302 a_100820_n36322.n2 a_100820_n36322.n1 7.46075
R55303 a_106676_n30339.t2 a_106676_n30339.n0 10.3838
R55304 a_106676_n30339.n0 a_106676_n30339.t0 10.3566
R55305 a_106676_n30339.n0 a_106676_n30339.t1 10.0407
R55306 a_106676_n30339.n0 a_106676_n30339.t3 9.57605
R55307 a_83153_11614.n2 a_83153_11614.t15 12.8637
R55308 a_83153_11614.n1 a_83153_11614.t6 10.7018
R55309 a_83153_11614.n1 a_83153_11614.t2 10.1659
R55310 a_83153_11614.n1 a_83153_11614.t0 9.64387
R55311 a_83153_11614.t4 a_83153_11614.n1 9.27665
R55312 a_83153_11614.n1 a_83153_11614.n2 8.75198
R55313 a_83153_11614.n2 a_83153_11614.t14 8.14051
R55314 a_83153_11614.n2 a_83153_11614.t10 8.14051
R55315 a_83153_11614.n2 a_83153_11614.t22 8.14051
R55316 a_83153_11614.n2 a_83153_11614.t16 8.14051
R55317 a_83153_11614.n2 a_83153_11614.t23 8.06917
R55318 a_83153_11614.n2 a_83153_11614.t20 8.06917
R55319 a_83153_11614.n2 a_83153_11614.t9 8.06917
R55320 a_83153_11614.n2 a_83153_11614.t12 8.06917
R55321 a_83153_11614.n2 a_83153_11614.t19 8.06917
R55322 a_83153_11614.n2 a_83153_11614.t11 8.06917
R55323 a_83153_11614.n2 a_83153_11614.t21 8.06917
R55324 a_83153_11614.n0 a_83153_11614.t3 7.94068
R55325 a_83153_11614.n1 a_83153_11614.t7 7.72524
R55326 a_83153_11614.n0 a_83153_11614.t1 7.22855
R55327 a_83153_11614.n1 a_83153_11614.t5 7.17942
R55328 a_83153_11614.t13 a_83153_11614.n2 8.33649
R55329 a_83153_11614.n2 a_83153_11614.t17 8.33649
R55330 a_83153_11614.t18 a_83153_11614.n2 8.33556
R55331 a_83153_11614.n2 a_83153_11614.t8 8.33556
R55332 a_83153_11614.n1 a_83153_11614.n0 7.46075
R55333 a_86903_n14095.t0 a_86903_n14095.t2 61.4377
R55334 a_86903_n14095.t0 a_86903_n14095.n0 13.0169
R55335 a_86903_n14095.n1 a_86903_n14095.n0 10.9309
R55336 a_86903_n14095.t0 a_86903_n14095.t1 8.5021
R55337 a_86903_n14095.n1 a_86903_n14095.t6 8.44198
R55338 a_86903_n14095.n1 a_86903_n14095.t8 8.44198
R55339 a_86903_n14095.n0 a_86903_n14095.t3 8.44198
R55340 a_86903_n14095.n0 a_86903_n14095.t7 8.44198
R55341 a_86903_n14095.n1 a_86903_n14095.t9 8.10567
R55342 a_86903_n14095.n0 a_86903_n14095.t10 9.26955
R55343 a_86903_n14095.n1 a_86903_n14095.t4 8.65823
R55344 a_86903_n14095.n0 a_86903_n14095.t5 8.77493
R55345 a_89715_n17715.t1 a_89715_n17715.t5 64.7464
R55346 a_89715_n17715.t1 a_89715_n17715.t4 12.9273
R55347 a_89715_n17715.t0 a_89715_n17715.t1 10.1307
R55348 a_89715_n17715.t1 a_89715_n17715.t3 8.54643
R55349 a_89715_n17715.t1 a_89715_n17715.t2 7.50895
R55350 a_112559_4481.n1 a_112559_4481.t7 10.2515
R55351 a_112559_4481.n1 a_112559_4481.t5 10.2515
R55352 a_112559_4481.n1 a_112559_4481.t12 10.2515
R55353 a_112559_4481.n1 a_112559_4481.t17 10.2515
R55354 a_112559_4481.n1 a_112559_4481.t3 10.096
R55355 a_112559_4481.n1 a_112559_4481.t22 10.0935
R55356 a_112559_4481.n1 a_112559_4481.t9 10.0859
R55357 a_112559_4481.n1 a_112559_4481.t15 10.0808
R55358 a_112559_4481.n1 a_112559_4481.t19 9.53981
R55359 a_112559_4481.n1 a_112559_4481.t16 9.53981
R55360 a_112559_4481.n1 a_112559_4481.t11 9.53981
R55361 a_112559_4481.n1 a_112559_4481.t13 9.53981
R55362 a_112559_4481.n1 a_112559_4481.t21 9.53744
R55363 a_112559_4481.n1 a_112559_4481.t20 9.53744
R55364 a_112559_4481.n1 a_112559_4481.t14 9.53744
R55365 a_112559_4481.n1 a_112559_4481.t18 9.53744
R55366 a_112559_4481.n1 a_112559_4481.n0 8.41434
R55367 a_112559_4481.n1 a_112559_4481.t8 8.14082
R55368 a_112559_4481.n0 a_112559_4481.t6 8.13828
R55369 a_112559_4481.t1 a_112559_4481.t2 7.96115
R55370 a_112559_4481.t0 a_112559_4481.t1 7.94694
R55371 a_112559_4481.t1 a_112559_4481.n1 7.50666
R55372 a_112559_4481.n0 a_112559_4481.t4 7.48586
R55373 a_112559_4481.n1 a_112559_4481.t10 7.48333
R55374 a_30152_n36322.n0 a_30152_n36322.t14 13.7934
R55375 a_30152_n36322.n2 a_30152_n36322.t5 10.7024
R55376 a_30152_n36322.n2 a_30152_n36322.t3 10.1668
R55377 a_30152_n36322.n2 a_30152_n36322.t4 9.64458
R55378 a_30152_n36322.n2 a_30152_n36322.t6 9.27635
R55379 a_30152_n36322.n2 a_30152_n36322.n0 8.75198
R55380 a_30152_n36322.n0 a_30152_n36322.t13 8.14051
R55381 a_30152_n36322.n0 a_30152_n36322.t11 8.14051
R55382 a_30152_n36322.n0 a_30152_n36322.t18 8.14051
R55383 a_30152_n36322.n0 a_30152_n36322.t21 8.14051
R55384 a_30152_n36322.n0 a_30152_n36322.t15 8.06917
R55385 a_30152_n36322.n0 a_30152_n36322.t20 8.06917
R55386 a_30152_n36322.n0 a_30152_n36322.t17 8.06917
R55387 a_30152_n36322.n0 a_30152_n36322.t23 8.06917
R55388 a_30152_n36322.n0 a_30152_n36322.t22 8.06917
R55389 a_30152_n36322.n0 a_30152_n36322.t8 8.06917
R55390 a_30152_n36322.n0 a_30152_n36322.t9 8.06917
R55391 a_30152_n36322.n1 a_30152_n36322.t2 7.94157
R55392 a_30152_n36322.n2 a_30152_n36322.t7 7.72643
R55393 a_30152_n36322.n1 a_30152_n36322.t1 7.22925
R55394 a_30152_n36322.t0 a_30152_n36322.n2 7.17912
R55395 a_30152_n36322.n0 a_30152_n36322.t12 8.33554
R55396 a_30152_n36322.t10 a_30152_n36322.n0 8.33554
R55397 a_30152_n36322.n0 a_30152_n36322.t16 8.33647
R55398 a_30152_n36322.t19 a_30152_n36322.n0 8.33647
R55399 a_30152_n36322.n2 a_30152_n36322.n1 7.46075
R55400 a_47819_n35156.n0 a_47819_n35156.t12 10.2828
R55401 a_47819_n35156.t8 a_47819_n35156.t4 10.2828
R55402 a_47819_n35156.n0 a_47819_n35156.t11 10.2828
R55403 a_47819_n35156.n0 a_47819_n35156.t0 10.2828
R55404 a_47819_n35156.n0 a_47819_n35156.t6 10.1333
R55405 a_47819_n35156.t8 a_47819_n35156.t19 10.1333
R55406 a_47819_n35156.n0 a_47819_n35156.t2 10.1333
R55407 a_47819_n35156.n0 a_47819_n35156.t21 10.1333
R55408 a_47819_n35156.n0 a_47819_n35156.t18 9.57156
R55409 a_47819_n35156.t8 a_47819_n35156.t15 9.57156
R55410 a_47819_n35156.n0 a_47819_n35156.t17 9.57156
R55411 a_47819_n35156.n0 a_47819_n35156.t16 9.57156
R55412 a_47819_n35156.n0 a_47819_n35156.t14 9.57156
R55413 a_47819_n35156.t8 a_47819_n35156.t20 9.57156
R55414 a_47819_n35156.n0 a_47819_n35156.t13 9.57156
R55415 a_47819_n35156.n0 a_47819_n35156.t22 9.57156
R55416 a_47819_n35156.t8 a_47819_n35156.n1 8.94763
R55417 a_47819_n35156.t8 a_47819_n35156.t9 8.02827
R55418 a_47819_n35156.t8 a_47819_n35156.t10 8.0259
R55419 a_47819_n35156.n1 a_47819_n35156.t5 7.90799
R55420 a_47819_n35156.t1 a_47819_n35156.t8 7.90799
R55421 a_47819_n35156.n1 a_47819_n35156.t7 7.41865
R55422 a_47819_n35156.t8 a_47819_n35156.t3 7.41865
R55423 a_47819_n35156.t8 a_47819_n35156.n0 7.31642
R55424 a_51711_n12421.t0 a_51711_n12421.t1 78.206
R55425 a_51711_n12421.t0 a_51711_n12421.t2 24.9014
R55426 a_100820_n35156.n0 a_100820_n35156.t20 10.2828
R55427 a_100820_n35156.t1 a_100820_n35156.t7 10.2828
R55428 a_100820_n35156.n0 a_100820_n35156.t19 10.2828
R55429 a_100820_n35156.n0 a_100820_n35156.t3 10.2828
R55430 a_100820_n35156.n0 a_100820_n35156.t9 10.1333
R55431 a_100820_n35156.t1 a_100820_n35156.t11 10.1333
R55432 a_100820_n35156.n0 a_100820_n35156.t5 10.1333
R55433 a_100820_n35156.n0 a_100820_n35156.t12 10.1333
R55434 a_100820_n35156.n0 a_100820_n35156.t16 9.57156
R55435 a_100820_n35156.t1 a_100820_n35156.t13 9.57156
R55436 a_100820_n35156.n0 a_100820_n35156.t15 9.57156
R55437 a_100820_n35156.n0 a_100820_n35156.t14 9.57156
R55438 a_100820_n35156.n0 a_100820_n35156.t22 9.57156
R55439 a_100820_n35156.t1 a_100820_n35156.t17 9.57156
R55440 a_100820_n35156.n0 a_100820_n35156.t21 9.57156
R55441 a_100820_n35156.n0 a_100820_n35156.t18 9.57156
R55442 a_100820_n35156.t1 a_100820_n35156.n1 8.94763
R55443 a_100820_n35156.t1 a_100820_n35156.t0 8.02827
R55444 a_100820_n35156.t1 a_100820_n35156.t2 8.0259
R55445 a_100820_n35156.n1 a_100820_n35156.t8 7.90799
R55446 a_100820_n35156.t4 a_100820_n35156.t1 7.90799
R55447 a_100820_n35156.n1 a_100820_n35156.t10 7.41865
R55448 a_100820_n35156.t1 a_100820_n35156.t6 7.41865
R55449 a_100820_n35156.t1 a_100820_n35156.n0 7.31642
R55450 a_77225_4481.n1 a_77225_4481.t6 10.2515
R55451 a_77225_4481.n1 a_77225_4481.t0 10.2515
R55452 a_77225_4481.n1 a_77225_4481.t13 10.2515
R55453 a_77225_4481.n1 a_77225_4481.t16 10.2515
R55454 a_77225_4481.n1 a_77225_4481.t2 10.096
R55455 a_77225_4481.n1 a_77225_4481.t19 10.0935
R55456 a_77225_4481.n1 a_77225_4481.t4 10.0859
R55457 a_77225_4481.n1 a_77225_4481.t11 10.0808
R55458 a_77225_4481.n1 a_77225_4481.t21 9.53981
R55459 a_77225_4481.n1 a_77225_4481.t20 9.53981
R55460 a_77225_4481.n1 a_77225_4481.t17 9.53981
R55461 a_77225_4481.n1 a_77225_4481.t18 9.53981
R55462 a_77225_4481.n1 a_77225_4481.t15 9.53744
R55463 a_77225_4481.n1 a_77225_4481.t14 9.53744
R55464 a_77225_4481.n1 a_77225_4481.t22 9.53744
R55465 a_77225_4481.n1 a_77225_4481.t12 9.53744
R55466 a_77225_4481.n1 a_77225_4481.n0 8.41434
R55467 a_77225_4481.n1 a_77225_4481.t7 8.14082
R55468 a_77225_4481.n0 a_77225_4481.t1 8.13828
R55469 a_77225_4481.t8 a_77225_4481.t10 7.96115
R55470 a_77225_4481.t8 a_77225_4481.t9 7.94694
R55471 a_77225_4481.t8 a_77225_4481.n1 7.50666
R55472 a_77225_4481.n0 a_77225_4481.t3 7.48586
R55473 a_77225_4481.n1 a_77225_4481.t5 7.48333
R55474 a_106830_10388.n6 a_106830_10388.n1 10.2377
R55475 a_106830_10388.n5 a_106830_10388.t7 10.2108
R55476 a_106830_10388.n5 a_106830_10388.t4 9.99909
R55477 a_106830_10388.t0 a_106830_10388.n6 9.80443
R55478 a_106830_10388.n6 a_106830_10388.t2 9.55135
R55479 a_106830_10388.n0 a_106830_10388.t18 8.17385
R55480 a_106830_10388.n3 a_106830_10388.t15 8.17299
R55481 a_106830_10388.n3 a_106830_10388.t17 8.17134
R55482 a_106830_10388.n0 a_106830_10388.t14 8.16754
R55483 a_106830_10388.n1 a_106830_10388.t11 8.10567
R55484 a_106830_10388.n1 a_106830_10388.t10 8.10567
R55485 a_106830_10388.n3 a_106830_10388.t23 8.10567
R55486 a_106830_10388.n3 a_106830_10388.t8 8.10567
R55487 a_106830_10388.n1 a_106830_10388.t9 8.10567
R55488 a_106830_10388.n1 a_106830_10388.t16 8.10567
R55489 a_106830_10388.n0 a_106830_10388.t13 8.10567
R55490 a_106830_10388.n0 a_106830_10388.t21 8.10567
R55491 a_106830_10388.n7 a_106830_10388.t5 7.74799
R55492 a_106830_10388.n4 a_106830_10388.t1 7.73052
R55493 a_106830_10388.n7 a_106830_10388.t6 7.46478
R55494 a_106830_10388.n4 a_106830_10388.t3 7.1311
R55495 a_106830_10388.n5 a_106830_10388.n7 2.2505
R55496 a_106830_10388.n6 a_106830_10388.n4 2.2505
R55497 a_106830_10388.n1 a_106830_10388.t19 8.35731
R55498 a_106830_10388.n0 a_106830_10388.t12 8.38107
R55499 a_106830_10388.n1 a_106830_10388.t20 8.37583
R55500 a_106830_10388.n1 a_106830_10388.n0 4.35656
R55501 a_106830_10388.n6 a_106830_10388.n5 2.96863
R55502 a_106830_10388.n2 a_106830_10388.n1 1.0882
R55503 a_106830_10388.n2 a_106830_10388.n3 1.08408
R55504 a_106830_10388.n2 a_106830_10388.t22 8.66753
R55505 a_106676_4481.n0 a_106676_4481.t1 10.6581
R55506 a_106676_4481.n0 a_106676_4481.t3 10.2356
R55507 a_106676_4481.t2 a_106676_4481.n0 9.5019
R55508 a_106676_4481.n0 a_106676_4481.t0 9.34796
R55509 a_36032_n35156.t0 a_36032_n35156.n3 96.9245
R55510 a_36032_n35156.n1 a_36032_n35156.n0 10.9327
R55511 a_36032_n35156.n0 a_36032_n35156.t8 8.44198
R55512 a_36032_n35156.n0 a_36032_n35156.t10 8.44198
R55513 a_36032_n35156.n1 a_36032_n35156.t7 8.44198
R55514 a_36032_n35156.n1 a_36032_n35156.t9 8.44198
R55515 a_36032_n35156.n0 a_36032_n35156.t5 9.26917
R55516 a_36032_n35156.n1 a_36032_n35156.t6 8.10567
R55517 a_36032_n35156.n3 a_36032_n35156.t1 6.51122
R55518 a_36032_n35156.n3 a_36032_n35156.n0 6.50622
R55519 a_36032_n35156.t1 a_36032_n35156.t2 6.36267
R55520 a_36032_n35156.t1 a_36032_n35156.n2 4.84877
R55521 a_36032_n35156.n2 a_36032_n35156.t4 3.65383
R55522 a_36032_n35156.n1 a_36032_n35156.t12 8.65827
R55523 a_36032_n35156.n2 a_36032_n35156.t3 3.57094
R55524 a_36032_n35156.n0 a_36032_n35156.t11 8.77499
R55525 a_30152_n35156.t8 a_30152_n35156.t5 12.7136
R55526 a_30152_n35156.t8 a_30152_n35156.t18 10.2828
R55527 a_30152_n35156.t8 a_30152_n35156.t0 10.2828
R55528 a_30152_n35156.t8 a_30152_n35156.t17 10.2828
R55529 a_30152_n35156.t8 a_30152_n35156.t6 10.2828
R55530 a_30152_n35156.t8 a_30152_n35156.t2 10.1333
R55531 a_30152_n35156.t8 a_30152_n35156.t19 10.1333
R55532 a_30152_n35156.t8 a_30152_n35156.t4 10.1333
R55533 a_30152_n35156.t8 a_30152_n35156.t20 10.1333
R55534 a_30152_n35156.t8 a_30152_n35156.t11 9.72545
R55535 a_30152_n35156.t8 a_30152_n35156.t16 9.57156
R55536 a_30152_n35156.t8 a_30152_n35156.t22 9.57156
R55537 a_30152_n35156.t8 a_30152_n35156.t15 9.57156
R55538 a_30152_n35156.t8 a_30152_n35156.t12 9.57156
R55539 a_30152_n35156.t8 a_30152_n35156.t14 9.57156
R55540 a_30152_n35156.t8 a_30152_n35156.t21 9.57156
R55541 a_30152_n35156.t8 a_30152_n35156.t13 9.57156
R55542 a_30152_n35156.t8 a_30152_n35156.t23 9.57156
R55543 a_30152_n35156.t11 a_30152_n35156.t9 8.02827
R55544 a_30152_n35156.t8 a_30152_n35156.t10 8.0259
R55545 a_30152_n35156.t8 a_30152_n35156.t7 7.90799
R55546 a_30152_n35156.t1 a_30152_n35156.t8 7.90799
R55547 a_30152_n35156.t8 a_30152_n35156.t3 7.41865
R55548 a_89163_10388.n6 a_89163_10388.n1 10.2377
R55549 a_89163_10388.n5 a_89163_10388.t3 10.2108
R55550 a_89163_10388.n5 a_89163_10388.t2 9.99909
R55551 a_89163_10388.n6 a_89163_10388.t6 9.80443
R55552 a_89163_10388.t4 a_89163_10388.n6 9.55135
R55553 a_89163_10388.n0 a_89163_10388.t17 8.17385
R55554 a_89163_10388.n3 a_89163_10388.t9 8.17299
R55555 a_89163_10388.n3 a_89163_10388.t11 8.17134
R55556 a_89163_10388.n0 a_89163_10388.t8 8.16754
R55557 a_89163_10388.n1 a_89163_10388.t16 8.10567
R55558 a_89163_10388.n1 a_89163_10388.t14 8.10567
R55559 a_89163_10388.n3 a_89163_10388.t20 8.10567
R55560 a_89163_10388.n3 a_89163_10388.t21 8.10567
R55561 a_89163_10388.n1 a_89163_10388.t13 8.10567
R55562 a_89163_10388.n1 a_89163_10388.t18 8.10567
R55563 a_89163_10388.n0 a_89163_10388.t12 8.10567
R55564 a_89163_10388.n0 a_89163_10388.t19 8.10567
R55565 a_89163_10388.n7 a_89163_10388.t0 7.74799
R55566 a_89163_10388.n4 a_89163_10388.t7 7.73052
R55567 a_89163_10388.n7 a_89163_10388.t1 7.46478
R55568 a_89163_10388.n4 a_89163_10388.t5 7.1311
R55569 a_89163_10388.n5 a_89163_10388.n7 2.2505
R55570 a_89163_10388.n6 a_89163_10388.n4 2.2505
R55571 a_89163_10388.n1 a_89163_10388.t22 8.35731
R55572 a_89163_10388.n0 a_89163_10388.t15 8.38107
R55573 a_89163_10388.n1 a_89163_10388.t23 8.37583
R55574 a_89163_10388.n1 a_89163_10388.n0 4.35656
R55575 a_89163_10388.n6 a_89163_10388.n5 2.96863
R55576 a_89163_10388.n2 a_89163_10388.n1 1.0882
R55577 a_89163_10388.n2 a_89163_10388.n3 1.08408
R55578 a_89163_10388.n2 a_89163_10388.t10 8.66753
R55579 a_89033_13546.n1 a_89033_13546.n0 26.5215
R55580 a_89033_13546.t0 a_89033_13546.n1 11.5094
R55581 a_89033_13546.n0 a_89033_13546.t3 10.937
R55582 a_89033_13546.n0 a_89033_13546.t2 9.33982
R55583 a_89033_13546.n1 a_89033_13546.t1 9.24966
R55584 a_65486_10448.n0 a_65486_10448.t2 10.2828
R55585 a_65486_10448.t10 a_65486_10448.t6 10.2828
R55586 a_65486_10448.n0 a_65486_10448.t19 10.2828
R55587 a_65486_10448.n0 a_65486_10448.t16 10.2828
R55588 a_65486_10448.n0 a_65486_10448.t17 10.1333
R55589 a_65486_10448.t10 a_65486_10448.t18 10.1333
R55590 a_65486_10448.n0 a_65486_10448.t0 10.1333
R55591 a_65486_10448.n0 a_65486_10448.t4 10.1333
R55592 a_65486_10448.n0 a_65486_10448.t13 9.57156
R55593 a_65486_10448.n0 a_65486_10448.t11 9.57156
R55594 a_65486_10448.t10 a_65486_10448.t12 9.57156
R55595 a_65486_10448.n0 a_65486_10448.t15 9.57156
R55596 a_65486_10448.n0 a_65486_10448.t22 9.57156
R55597 a_65486_10448.n0 a_65486_10448.t20 9.57156
R55598 a_65486_10448.t10 a_65486_10448.t21 9.57156
R55599 a_65486_10448.n0 a_65486_10448.t14 9.57156
R55600 a_65486_10448.t10 a_65486_10448.n1 8.94763
R55601 a_65486_10448.t10 a_65486_10448.t9 8.02945
R55602 a_65486_10448.t10 a_65486_10448.t8 8.02708
R55603 a_65486_10448.t10 a_65486_10448.t3 7.90829
R55604 a_65486_10448.n1 a_65486_10448.t7 7.90829
R55605 a_65486_10448.n1 a_65486_10448.t5 7.41776
R55606 a_65486_10448.t1 a_65486_10448.t10 7.41776
R55607 a_65486_10448.t10 a_65486_10448.n0 7.31642
R55608 a_36032_11614.t0 a_36032_11614.t2 74.3465
R55609 a_36032_11614.t0 a_36032_11614.n0 13.0169
R55610 a_36032_11614.n1 a_36032_11614.n0 10.9309
R55611 a_36032_11614.t0 a_36032_11614.t1 8.5021
R55612 a_36032_11614.n1 a_36032_11614.t9 8.44198
R55613 a_36032_11614.n1 a_36032_11614.t5 8.44198
R55614 a_36032_11614.n0 a_36032_11614.t6 8.44198
R55615 a_36032_11614.n0 a_36032_11614.t10 8.44198
R55616 a_36032_11614.n1 a_36032_11614.t3 8.10567
R55617 a_36032_11614.n0 a_36032_11614.t4 9.26955
R55618 a_36032_11614.n1 a_36032_11614.t7 8.65823
R55619 a_36032_11614.n0 a_36032_11614.t8 8.77493
R55620 a_43010_10448.t0 a_43010_10448.t4 76.8811
R55621 a_43010_10448.t0 a_43010_10448.t1 8.54643
R55622 a_43010_10448.t0 a_43010_10448.t2 8.17727
R55623 a_43010_10448.t0 a_43010_10448.t3 7.03425
R55624 a_81205_n14095.t0 a_81205_n14095.t2 45.7073
R55625 a_81205_n14095.t0 a_81205_n14095.n0 13.0169
R55626 a_81205_n14095.n1 a_81205_n14095.n0 10.9309
R55627 a_81205_n14095.t0 a_81205_n14095.t1 8.5021
R55628 a_81205_n14095.n1 a_81205_n14095.t3 8.44198
R55629 a_81205_n14095.n1 a_81205_n14095.t7 8.44198
R55630 a_81205_n14095.n0 a_81205_n14095.t8 8.44198
R55631 a_81205_n14095.n0 a_81205_n14095.t4 8.44198
R55632 a_81205_n14095.n1 a_81205_n14095.t5 8.10567
R55633 a_81205_n14095.n0 a_81205_n14095.t6 9.26955
R55634 a_81205_n14095.n1 a_81205_n14095.t9 8.65823
R55635 a_81205_n14095.n0 a_81205_n14095.t10 8.77493
R55636 a_89163_n36382.n5 a_89163_n36382.n1 10.2377
R55637 a_89163_n36382.n4 a_89163_n36382.t6 10.2105
R55638 a_89163_n36382.n4 a_89163_n36382.t5 9.99998
R55639 a_89163_n36382.n5 a_89163_n36382.t1 9.80532
R55640 a_89163_n36382.n5 a_89163_n36382.t3 9.55206
R55641 a_89163_n36382.n0 a_89163_n36382.t12 8.17385
R55642 a_89163_n36382.n3 a_89163_n36382.t10 8.17299
R55643 a_89163_n36382.n3 a_89163_n36382.t13 8.17134
R55644 a_89163_n36382.n0 a_89163_n36382.t11 8.16754
R55645 a_89163_n36382.n1 a_89163_n36382.t14 8.10567
R55646 a_89163_n36382.n1 a_89163_n36382.t19 8.10567
R55647 a_89163_n36382.n3 a_89163_n36382.t9 8.10567
R55648 a_89163_n36382.n3 a_89163_n36382.t22 8.10567
R55649 a_89163_n36382.n1 a_89163_n36382.t16 8.10567
R55650 a_89163_n36382.n1 a_89163_n36382.t18 8.10567
R55651 a_89163_n36382.n0 a_89163_n36382.t8 8.10567
R55652 a_89163_n36382.n0 a_89163_n36382.t23 8.10567
R55653 a_89163_n36382.n6 a_89163_n36382.t4 7.74888
R55654 a_89163_n36382.t0 a_89163_n36382.n7 7.73041
R55655 a_89163_n36382.n6 a_89163_n36382.t7 7.46359
R55656 a_89163_n36382.n7 a_89163_n36382.t2 7.13181
R55657 a_89163_n36382.n4 a_89163_n36382.n6 2.2505
R55658 a_89163_n36382.n7 a_89163_n36382.n5 2.2505
R55659 a_89163_n36382.t17 a_89163_n36382.n1 8.35729
R55660 a_89163_n36382.n1 a_89163_n36382.t15 8.37586
R55661 a_89163_n36382.n0 a_89163_n36382.t20 8.38104
R55662 a_89163_n36382.n1 a_89163_n36382.n0 4.35658
R55663 a_89163_n36382.n5 a_89163_n36382.n4 2.96863
R55664 a_89163_n36382.n2 a_89163_n36382.n1 1.08819
R55665 a_89163_n36382.n2 a_89163_n36382.n3 1.08408
R55666 a_89163_n36382.n2 a_89163_n36382.t21 8.6675
R55667 a_106809_n5150.t0 a_106809_n5150.t2 42.6538
R55668 a_106809_n5150.t2 a_106809_n5150.t3 9.77323
R55669 a_106809_n5150.t2 a_106809_n5150.t1 8.17727
R55670 a_41891_n29181.n0 a_41891_n29181.t14 10.2515
R55671 a_41891_n29181.n1 a_41891_n29181.t9 10.2515
R55672 a_41891_n29181.n0 a_41891_n29181.t18 10.2515
R55673 a_41891_n29181.n0 a_41891_n29181.t7 10.2515
R55674 a_41891_n29181.n0 a_41891_n29181.t3 10.096
R55675 a_41891_n29181.n1 a_41891_n29181.t19 10.0935
R55676 a_41891_n29181.n0 a_41891_n29181.t5 10.0859
R55677 a_41891_n29181.n0 a_41891_n29181.t12 10.0808
R55678 a_41891_n29181.n0 a_41891_n29181.t11 9.53981
R55679 a_41891_n29181.n1 a_41891_n29181.t22 9.53981
R55680 a_41891_n29181.n0 a_41891_n29181.t16 9.53981
R55681 a_41891_n29181.n0 a_41891_n29181.t17 9.53981
R55682 a_41891_n29181.n0 a_41891_n29181.t21 9.53744
R55683 a_41891_n29181.n1 a_41891_n29181.t20 9.53744
R55684 a_41891_n29181.n0 a_41891_n29181.t13 9.53744
R55685 a_41891_n29181.n0 a_41891_n29181.t15 9.53744
R55686 a_41891_n29181.n1 a_41891_n29181.n0 9.16839
R55687 a_41891_n29181.n1 a_41891_n29181.t8 8.14051
R55688 a_41891_n29181.n1 a_41891_n29181.t10 8.13798
R55689 a_41891_n29181.t0 a_41891_n29181.t1 7.95997
R55690 a_41891_n29181.t0 a_41891_n29181.t2 7.94576
R55691 a_41891_n29181.t0 a_41891_n29181.n1 7.50666
R55692 a_41891_n29181.n1 a_41891_n29181.t4 7.48675
R55693 a_41891_n29181.n1 a_41891_n29181.t6 7.48422
R55694 a_89009_n27257.n0 a_89009_n27257.t3 10.6581
R55695 a_89009_n27257.n0 a_89009_n27257.t1 10.2358
R55696 a_89009_n27257.t0 a_89009_n27257.n0 9.50202
R55697 a_89009_n27257.n0 a_89009_n27257.t2 9.34796
R55698 a_71496_n36382.n5 a_71496_n36382.n1 10.2377
R55699 a_71496_n36382.n4 a_71496_n36382.t1 10.2105
R55700 a_71496_n36382.n4 a_71496_n36382.t2 9.99998
R55701 a_71496_n36382.n5 a_71496_n36382.t5 9.80532
R55702 a_71496_n36382.n5 a_71496_n36382.t7 9.55206
R55703 a_71496_n36382.n0 a_71496_n36382.t10 8.17385
R55704 a_71496_n36382.n3 a_71496_n36382.t18 8.17299
R55705 a_71496_n36382.n3 a_71496_n36382.t11 8.17134
R55706 a_71496_n36382.n0 a_71496_n36382.t23 8.16754
R55707 a_71496_n36382.n1 a_71496_n36382.t16 8.10567
R55708 a_71496_n36382.n1 a_71496_n36382.t20 8.10567
R55709 a_71496_n36382.n3 a_71496_n36382.t15 8.10567
R55710 a_71496_n36382.n3 a_71496_n36382.t22 8.10567
R55711 a_71496_n36382.n1 a_71496_n36382.t17 8.10567
R55712 a_71496_n36382.n1 a_71496_n36382.t19 8.10567
R55713 a_71496_n36382.n0 a_71496_n36382.t14 8.10567
R55714 a_71496_n36382.n0 a_71496_n36382.t9 8.10567
R55715 a_71496_n36382.n6 a_71496_n36382.t0 7.74888
R55716 a_71496_n36382.t4 a_71496_n36382.n7 7.73041
R55717 a_71496_n36382.n6 a_71496_n36382.t3 7.46359
R55718 a_71496_n36382.n7 a_71496_n36382.t6 7.13181
R55719 a_71496_n36382.n4 a_71496_n36382.n6 2.2505
R55720 a_71496_n36382.n7 a_71496_n36382.n5 2.2505
R55721 a_71496_n36382.t8 a_71496_n36382.n1 8.35729
R55722 a_71496_n36382.n1 a_71496_n36382.t21 8.37586
R55723 a_71496_n36382.n0 a_71496_n36382.t12 8.38104
R55724 a_71496_n36382.n1 a_71496_n36382.n0 4.35658
R55725 a_71496_n36382.n5 a_71496_n36382.n4 2.96863
R55726 a_71496_n36382.n2 a_71496_n36382.n1 1.08819
R55727 a_71496_n36382.n2 a_71496_n36382.n3 1.08408
R55728 a_71496_n36382.n2 a_71496_n36382.t13 8.6675
R55729 a_53699_n36322.n1 a_53699_n36322.n0 26.5254
R55730 a_53699_n36322.n0 a_53699_n36322.t2 11.5094
R55731 a_53699_n36322.n1 a_53699_n36322.t1 10.937
R55732 a_53699_n36322.t0 a_53699_n36322.n1 9.33982
R55733 a_53699_n36322.n0 a_53699_n36322.t3 9.24966
R55734 a_44363_n16007.t0 a_44363_n16007.t2 56.3087
R55735 a_44363_n16007.t2 a_44363_n16007.t1 18.4133
R55736 a_71366_n35156.t0 a_71366_n35156.n3 69.4088
R55737 a_71366_n35156.n1 a_71366_n35156.n0 10.9327
R55738 a_71366_n35156.n0 a_71366_n35156.t9 8.44198
R55739 a_71366_n35156.n0 a_71366_n35156.t11 8.44198
R55740 a_71366_n35156.n1 a_71366_n35156.t8 8.44198
R55741 a_71366_n35156.n1 a_71366_n35156.t10 8.44198
R55742 a_71366_n35156.n0 a_71366_n35156.t12 9.26917
R55743 a_71366_n35156.n1 a_71366_n35156.t5 8.10567
R55744 a_71366_n35156.n3 a_71366_n35156.t4 6.51122
R55745 a_71366_n35156.n3 a_71366_n35156.n0 6.50622
R55746 a_71366_n35156.t4 a_71366_n35156.t2 6.36267
R55747 a_71366_n35156.t4 a_71366_n35156.n2 4.84877
R55748 a_71366_n35156.n2 a_71366_n35156.t3 3.65383
R55749 a_71366_n35156.n1 a_71366_n35156.t7 8.65827
R55750 a_71366_n35156.n2 a_71366_n35156.t1 3.57094
R55751 a_71366_n35156.n0 a_71366_n35156.t6 8.77499
R55752 a_78344_n36322.t0 a_78344_n36322.t2 67.5623
R55753 a_78344_n36322.t2 a_78344_n36322.t1 9.77323
R55754 a_78344_n36322.t2 a_78344_n36322.t3 8.17727
R55755 a_39179_n19595.t0 a_39179_n19595.t1 34.4821
R55756 a_39179_n19595.t0 a_39179_n19595.t2 24.9025
R55757 a_59558_4481.n1 a_59558_4481.t5 10.2515
R55758 a_59558_4481.n1 a_59558_4481.t7 10.2515
R55759 a_59558_4481.n1 a_59558_4481.t14 10.2515
R55760 a_59558_4481.n1 a_59558_4481.t19 10.2515
R55761 a_59558_4481.n1 a_59558_4481.t9 10.096
R55762 a_59558_4481.n1 a_59558_4481.t13 10.0935
R55763 a_59558_4481.n1 a_59558_4481.t3 10.0859
R55764 a_59558_4481.n1 a_59558_4481.t18 10.0808
R55765 a_59558_4481.n1 a_59558_4481.t21 9.53981
R55766 a_59558_4481.n1 a_59558_4481.t17 9.53981
R55767 a_59558_4481.n1 a_59558_4481.t12 9.53981
R55768 a_59558_4481.n1 a_59558_4481.t15 9.53981
R55769 a_59558_4481.n1 a_59558_4481.t11 9.53744
R55770 a_59558_4481.n1 a_59558_4481.t22 9.53744
R55771 a_59558_4481.n1 a_59558_4481.t16 9.53744
R55772 a_59558_4481.n1 a_59558_4481.t20 9.53744
R55773 a_59558_4481.n1 a_59558_4481.n0 8.41434
R55774 a_59558_4481.n1 a_59558_4481.t6 8.14082
R55775 a_59558_4481.n0 a_59558_4481.t8 8.13828
R55776 a_59558_4481.t0 a_59558_4481.t2 7.96115
R55777 a_59558_4481.t2 a_59558_4481.t1 7.94694
R55778 a_59558_4481.t2 a_59558_4481.n1 7.50666
R55779 a_59558_4481.n0 a_59558_4481.t10 7.48586
R55780 a_59558_4481.n1 a_59558_4481.t4 7.48333
R55781 a_53699_n35156.t0 a_53699_n35156.n3 80.9771
R55782 a_53699_n35156.n1 a_53699_n35156.n0 10.9327
R55783 a_53699_n35156.n0 a_53699_n35156.t12 8.44198
R55784 a_53699_n35156.n0 a_53699_n35156.t8 8.44198
R55785 a_53699_n35156.n1 a_53699_n35156.t11 8.44198
R55786 a_53699_n35156.n1 a_53699_n35156.t7 8.44198
R55787 a_53699_n35156.n0 a_53699_n35156.t5 9.26917
R55788 a_53699_n35156.n1 a_53699_n35156.t6 8.10567
R55789 a_53699_n35156.n3 a_53699_n35156.t3 6.51122
R55790 a_53699_n35156.n3 a_53699_n35156.n0 6.50622
R55791 a_53699_n35156.t3 a_53699_n35156.t4 6.36267
R55792 a_53699_n35156.t3 a_53699_n35156.n2 4.84877
R55793 a_53699_n35156.n2 a_53699_n35156.t1 3.65383
R55794 a_53699_n35156.n1 a_53699_n35156.t10 8.65827
R55795 a_53699_n35156.n2 a_53699_n35156.t2 3.57094
R55796 a_53699_n35156.n0 a_53699_n35156.t9 8.77499
R55797 a_83325_n29313.t0 a_83325_n29313.t1 23.2303
R55798 a_83325_n29313.t0 a_83325_n29313.t2 21.6695
R55799 a_94892_n29181.n0 a_94892_n29181.t18 10.2515
R55800 a_94892_n29181.n1 a_94892_n29181.t0 10.2515
R55801 a_94892_n29181.n0 a_94892_n29181.t22 10.2515
R55802 a_94892_n29181.n0 a_94892_n29181.t2 10.2515
R55803 a_94892_n29181.n0 a_94892_n29181.t4 10.096
R55804 a_94892_n29181.n1 a_94892_n29181.t11 10.0935
R55805 a_94892_n29181.n0 a_94892_n29181.t6 10.0859
R55806 a_94892_n29181.n0 a_94892_n29181.t16 10.0808
R55807 a_94892_n29181.n0 a_94892_n29181.t15 9.53981
R55808 a_94892_n29181.n1 a_94892_n29181.t14 9.53981
R55809 a_94892_n29181.n0 a_94892_n29181.t20 9.53981
R55810 a_94892_n29181.n0 a_94892_n29181.t21 9.53981
R55811 a_94892_n29181.n0 a_94892_n29181.t13 9.53744
R55812 a_94892_n29181.n1 a_94892_n29181.t12 9.53744
R55813 a_94892_n29181.n0 a_94892_n29181.t17 9.53744
R55814 a_94892_n29181.n0 a_94892_n29181.t19 9.53744
R55815 a_94892_n29181.n1 a_94892_n29181.n0 9.16839
R55816 a_94892_n29181.n1 a_94892_n29181.t3 8.14051
R55817 a_94892_n29181.n1 a_94892_n29181.t1 8.13798
R55818 a_94892_n29181.t9 a_94892_n29181.t10 7.95997
R55819 a_94892_n29181.t8 a_94892_n29181.t9 7.94576
R55820 a_94892_n29181.t9 a_94892_n29181.n1 7.50666
R55821 a_94892_n29181.n1 a_94892_n29181.t5 7.48675
R55822 a_94892_n29181.n1 a_94892_n29181.t7 7.48422
R55823 I1U I1U.t1 3.63879
R55824 I1U.n0 I1U.t5 2.56243
R55825 I1U.n0 I1U.t4 2.32184
R55826 I1U.n1 I1U.t2 2.32184
R55827 I1U.n2 I1U.t3 2.32184
R55828 I1U.n3 I1U.t6 2.32184
R55829 I1U.n4 I1U.t0 1.34815
R55830 I1U.n4 I1U.n3 1.20346
R55831 I1U I1U.n4 1.12236
R55832 I1U.n1 I1U.n0 0.242306
R55833 I1U.n3 I1U.n2 0.241697
R55834 I1U.n2 I1U.n1 0.241089
R55835 a_77225_n29181.n0 a_77225_n29181.t15 10.2515
R55836 a_77225_n29181.n1 a_77225_n29181.t6 10.2515
R55837 a_77225_n29181.n0 a_77225_n29181.t19 10.2515
R55838 a_77225_n29181.n0 a_77225_n29181.t4 10.2515
R55839 a_77225_n29181.n0 a_77225_n29181.t2 10.096
R55840 a_77225_n29181.n1 a_77225_n29181.t13 10.0935
R55841 a_77225_n29181.n0 a_77225_n29181.t0 10.0859
R55842 a_77225_n29181.n0 a_77225_n29181.t18 10.0808
R55843 a_77225_n29181.n0 a_77225_n29181.t16 9.53981
R55844 a_77225_n29181.n1 a_77225_n29181.t14 9.53981
R55845 a_77225_n29181.n0 a_77225_n29181.t21 9.53981
R55846 a_77225_n29181.n0 a_77225_n29181.t22 9.53981
R55847 a_77225_n29181.n0 a_77225_n29181.t20 9.53744
R55848 a_77225_n29181.n1 a_77225_n29181.t17 9.53744
R55849 a_77225_n29181.n0 a_77225_n29181.t11 9.53744
R55850 a_77225_n29181.n0 a_77225_n29181.t12 9.53744
R55851 a_77225_n29181.n1 a_77225_n29181.n0 9.16839
R55852 a_77225_n29181.n1 a_77225_n29181.t5 8.14051
R55853 a_77225_n29181.n1 a_77225_n29181.t7 8.13798
R55854 a_77225_n29181.t8 a_77225_n29181.t9 7.95997
R55855 a_77225_n29181.t9 a_77225_n29181.t10 7.94576
R55856 a_77225_n29181.t9 a_77225_n29181.n1 7.50666
R55857 a_77225_n29181.n1 a_77225_n29181.t3 7.48675
R55858 a_77225_n29181.n1 a_77225_n29181.t1 7.48422
R55859 a_64243_n1756.t1 a_64243_n1756.t2 24.9014
R55860 a_64243_n1756.t0 a_64243_n1756.t1 23.8039
R55861 a_63161_n5344.t0 a_63161_n5344.t1 30.6913
R55862 a_63161_n5344.t1 a_63161_n5344.t2 15.0742
R55863 a_30152_11614.n2 a_30152_11614.t22 12.8637
R55864 a_30152_11614.t4 a_30152_11614.n1 10.7018
R55865 a_30152_11614.n1 a_30152_11614.t1 10.1659
R55866 a_30152_11614.n1 a_30152_11614.t0 9.64387
R55867 a_30152_11614.n1 a_30152_11614.t7 9.27665
R55868 a_30152_11614.n1 a_30152_11614.n2 8.75198
R55869 a_30152_11614.n2 a_30152_11614.t19 8.14051
R55870 a_30152_11614.n2 a_30152_11614.t15 8.14051
R55871 a_30152_11614.n2 a_30152_11614.t12 8.14051
R55872 a_30152_11614.n2 a_30152_11614.t23 8.14051
R55873 a_30152_11614.n2 a_30152_11614.t16 8.06917
R55874 a_30152_11614.n2 a_30152_11614.t13 8.06917
R55875 a_30152_11614.n2 a_30152_11614.t14 8.06917
R55876 a_30152_11614.n2 a_30152_11614.t18 8.06917
R55877 a_30152_11614.n2 a_30152_11614.t10 8.06917
R55878 a_30152_11614.n2 a_30152_11614.t20 8.06917
R55879 a_30152_11614.n2 a_30152_11614.t11 8.06917
R55880 a_30152_11614.n0 a_30152_11614.t2 7.94068
R55881 a_30152_11614.n1 a_30152_11614.t6 7.72524
R55882 a_30152_11614.n0 a_30152_11614.t3 7.22855
R55883 a_30152_11614.n1 a_30152_11614.t5 7.17942
R55884 a_30152_11614.t21 a_30152_11614.n2 8.33649
R55885 a_30152_11614.n2 a_30152_11614.t8 8.33649
R55886 a_30152_11614.t9 a_30152_11614.n2 8.33556
R55887 a_30152_11614.n2 a_30152_11614.t17 8.33556
R55888 a_30152_11614.n1 a_30152_11614.n0 7.46075
R55889 a_36008_4481.n0 a_36008_4481.t1 10.6581
R55890 a_36008_4481.t2 a_36008_4481.n0 10.2346
R55891 a_36008_4481.n0 a_36008_4481.t3 9.5029
R55892 a_36008_4481.n0 a_36008_4481.t0 9.34796
R55893 a_96011_n36322.t0 a_96011_n36322.t1 39.0132
R55894 a_96011_n36322.t1 a_96011_n36322.t3 9.77323
R55895 a_96011_n36322.t1 a_96011_n36322.t2 8.17727
R55896 a_89033_n35156.t0 a_89033_n35156.n3 36.8446
R55897 a_89033_n35156.n1 a_89033_n35156.n0 10.9327
R55898 a_89033_n35156.n0 a_89033_n35156.t6 8.44198
R55899 a_89033_n35156.n0 a_89033_n35156.t8 8.44198
R55900 a_89033_n35156.n1 a_89033_n35156.t5 8.44198
R55901 a_89033_n35156.n1 a_89033_n35156.t7 8.44198
R55902 a_89033_n35156.n0 a_89033_n35156.t11 9.26917
R55903 a_89033_n35156.n1 a_89033_n35156.t12 8.10567
R55904 a_89033_n35156.n3 a_89033_n35156.t4 6.51122
R55905 a_89033_n35156.n3 a_89033_n35156.n0 6.50622
R55906 a_89033_n35156.t4 a_89033_n35156.t3 6.36267
R55907 a_89033_n35156.t4 a_89033_n35156.n2 4.84877
R55908 a_89033_n35156.n2 a_89033_n35156.t2 3.65383
R55909 a_89033_n35156.n1 a_89033_n35156.t10 8.65827
R55910 a_89033_n35156.n2 a_89033_n35156.t1 3.57094
R55911 a_89033_n35156.n0 a_89033_n35156.t9 8.77499
R55912 a_83153_n35156.t10 a_83153_n35156.t3 12.7136
R55913 a_83153_n35156.t10 a_83153_n35156.t21 10.2828
R55914 a_83153_n35156.t10 a_83153_n35156.t0 10.2828
R55915 a_83153_n35156.t10 a_83153_n35156.t20 10.2828
R55916 a_83153_n35156.t10 a_83153_n35156.t6 10.2828
R55917 a_83153_n35156.t10 a_83153_n35156.t4 10.1333
R55918 a_83153_n35156.t10 a_83153_n35156.t22 10.1333
R55919 a_83153_n35156.t10 a_83153_n35156.t2 10.1333
R55920 a_83153_n35156.t10 a_83153_n35156.t23 10.1333
R55921 a_83153_n35156.t10 a_83153_n35156.t11 9.72545
R55922 a_83153_n35156.t10 a_83153_n35156.t19 9.57156
R55923 a_83153_n35156.t10 a_83153_n35156.t13 9.57156
R55924 a_83153_n35156.t10 a_83153_n35156.t18 9.57156
R55925 a_83153_n35156.t10 a_83153_n35156.t15 9.57156
R55926 a_83153_n35156.t10 a_83153_n35156.t17 9.57156
R55927 a_83153_n35156.t10 a_83153_n35156.t12 9.57156
R55928 a_83153_n35156.t10 a_83153_n35156.t16 9.57156
R55929 a_83153_n35156.t10 a_83153_n35156.t14 9.57156
R55930 a_83153_n35156.t11 a_83153_n35156.t8 8.02827
R55931 a_83153_n35156.t10 a_83153_n35156.t9 8.0259
R55932 a_83153_n35156.t10 a_83153_n35156.t7 7.90799
R55933 a_83153_n35156.t1 a_83153_n35156.t10 7.90799
R55934 a_83153_n35156.t10 a_83153_n35156.t5 7.41865
R55935 a_56895_n16009.t0 a_56895_n16009.t1 97.9575
R55936 a_30324_n29313.t0 a_30324_n29313.t2 23.2303
R55937 a_30324_n29313.t0 a_30324_n29313.t1 21.6695
R55938 a_112559_n29181.n0 a_112559_n29181.t14 10.2515
R55939 a_112559_n29181.n1 a_112559_n29181.t9 10.2515
R55940 a_112559_n29181.n0 a_112559_n29181.t20 10.2515
R55941 a_112559_n29181.n0 a_112559_n29181.t3 10.2515
R55942 a_112559_n29181.n0 a_112559_n29181.t7 10.096
R55943 a_112559_n29181.n1 a_112559_n29181.t16 10.0935
R55944 a_112559_n29181.n0 a_112559_n29181.t5 10.0859
R55945 a_112559_n29181.n0 a_112559_n29181.t21 10.0808
R55946 a_112559_n29181.n0 a_112559_n29181.t13 9.53981
R55947 a_112559_n29181.n1 a_112559_n29181.t11 9.53981
R55948 a_112559_n29181.n0 a_112559_n29181.t17 9.53981
R55949 a_112559_n29181.n0 a_112559_n29181.t19 9.53981
R55950 a_112559_n29181.n0 a_112559_n29181.t12 9.53744
R55951 a_112559_n29181.n1 a_112559_n29181.t22 9.53744
R55952 a_112559_n29181.n0 a_112559_n29181.t15 9.53744
R55953 a_112559_n29181.n0 a_112559_n29181.t18 9.53744
R55954 a_112559_n29181.n1 a_112559_n29181.n0 9.16839
R55955 a_112559_n29181.n1 a_112559_n29181.t4 8.14051
R55956 a_112559_n29181.n1 a_112559_n29181.t10 8.13798
R55957 a_112559_n29181.t0 a_112559_n29181.t1 7.95997
R55958 a_112559_n29181.t1 a_112559_n29181.t2 7.94576
R55959 a_112559_n29181.t1 a_112559_n29181.n1 7.50666
R55960 a_112559_n29181.n1 a_112559_n29181.t8 7.48675
R55961 a_112559_n29181.n1 a_112559_n29181.t6 7.48422
R55962 a_47819_10448.n0 a_47819_10448.t3 10.2828
R55963 a_47819_10448.t1 a_47819_10448.t5 10.2828
R55964 a_47819_10448.n0 a_47819_10448.t19 10.2828
R55965 a_47819_10448.n0 a_47819_10448.t15 10.2828
R55966 a_47819_10448.n0 a_47819_10448.t12 10.1333
R55967 a_47819_10448.t1 a_47819_10448.t13 10.1333
R55968 a_47819_10448.n0 a_47819_10448.t9 10.1333
R55969 a_47819_10448.n0 a_47819_10448.t7 10.1333
R55970 a_47819_10448.n0 a_47819_10448.t18 9.57156
R55971 a_47819_10448.n0 a_47819_10448.t16 9.57156
R55972 a_47819_10448.t1 a_47819_10448.t17 9.57156
R55973 a_47819_10448.n0 a_47819_10448.t11 9.57156
R55974 a_47819_10448.n0 a_47819_10448.t22 9.57156
R55975 a_47819_10448.n0 a_47819_10448.t20 9.57156
R55976 a_47819_10448.t1 a_47819_10448.t21 9.57156
R55977 a_47819_10448.n0 a_47819_10448.t14 9.57156
R55978 a_47819_10448.t1 a_47819_10448.n1 8.94763
R55979 a_47819_10448.t1 a_47819_10448.t2 8.02945
R55980 a_47819_10448.t1 a_47819_10448.t0 8.02708
R55981 a_47819_10448.n1 a_47819_10448.t6 7.90829
R55982 a_47819_10448.t4 a_47819_10448.t1 7.90829
R55983 a_47819_10448.n1 a_47819_10448.t8 7.41776
R55984 a_47819_10448.t1 a_47819_10448.t10 7.41776
R55985 a_47819_10448.t1 a_47819_10448.n0 7.31642
R55986 a_47819_n36322.n0 a_47819_n36322.t13 13.7934
R55987 a_47819_n36322.t0 a_47819_n36322.n2 10.7024
R55988 a_47819_n36322.n2 a_47819_n36322.t7 10.1668
R55989 a_47819_n36322.n2 a_47819_n36322.t5 9.64458
R55990 a_47819_n36322.n2 a_47819_n36322.t2 9.27635
R55991 a_47819_n36322.n2 a_47819_n36322.n0 8.75198
R55992 a_47819_n36322.n0 a_47819_n36322.t17 8.14051
R55993 a_47819_n36322.n0 a_47819_n36322.t15 8.14051
R55994 a_47819_n36322.n0 a_47819_n36322.t23 8.14051
R55995 a_47819_n36322.n0 a_47819_n36322.t8 8.14051
R55996 a_47819_n36322.n0 a_47819_n36322.t14 8.06917
R55997 a_47819_n36322.n0 a_47819_n36322.t12 8.06917
R55998 a_47819_n36322.n0 a_47819_n36322.t11 8.06917
R55999 a_47819_n36322.n0 a_47819_n36322.t22 8.06917
R56000 a_47819_n36322.n0 a_47819_n36322.t20 8.06917
R56001 a_47819_n36322.n0 a_47819_n36322.t16 8.06917
R56002 a_47819_n36322.n0 a_47819_n36322.t19 8.06917
R56003 a_47819_n36322.n1 a_47819_n36322.t6 7.94157
R56004 a_47819_n36322.n2 a_47819_n36322.t1 7.72643
R56005 a_47819_n36322.n1 a_47819_n36322.t4 7.22925
R56006 a_47819_n36322.n2 a_47819_n36322.t3 7.17912
R56007 a_47819_n36322.n0 a_47819_n36322.t21 8.33554
R56008 a_47819_n36322.t18 a_47819_n36322.n0 8.33554
R56009 a_47819_n36322.n0 a_47819_n36322.t9 8.33647
R56010 a_47819_n36322.t10 a_47819_n36322.n0 8.33647
R56011 a_47819_n36322.n2 a_47819_n36322.n1 7.46075
R56012 a_83325_4421.t2 a_83325_4421.t0 21.6693
R56013 a_83325_4421.t1 a_83325_4421.t0 15.3476
R56014 a_84017_n17715.t2 a_84017_n17715.t4 49.024
R56015 a_84017_n17715.t2 a_84017_n17715.t1 13.8923
R56016 a_84017_n17715.t2 a_84017_n17715.t3 10.1307
R56017 a_84017_n17715.t0 a_84017_n17715.t2 8.54643
R56018 a_83153_n36322.n0 a_83153_n36322.t16 13.7934
R56019 a_83153_n36322.n2 a_83153_n36322.t5 10.7024
R56020 a_83153_n36322.n2 a_83153_n36322.t2 10.1668
R56021 a_83153_n36322.n2 a_83153_n36322.t3 9.64458
R56022 a_83153_n36322.n2 a_83153_n36322.t6 9.27635
R56023 a_83153_n36322.n2 a_83153_n36322.n0 8.75198
R56024 a_83153_n36322.n0 a_83153_n36322.t22 8.14051
R56025 a_83153_n36322.n0 a_83153_n36322.t20 8.14051
R56026 a_83153_n36322.n0 a_83153_n36322.t10 8.14051
R56027 a_83153_n36322.n0 a_83153_n36322.t13 8.14051
R56028 a_83153_n36322.n0 a_83153_n36322.t17 8.06917
R56029 a_83153_n36322.n0 a_83153_n36322.t11 8.06917
R56030 a_83153_n36322.n0 a_83153_n36322.t9 8.06917
R56031 a_83153_n36322.n0 a_83153_n36322.t8 8.06917
R56032 a_83153_n36322.n0 a_83153_n36322.t23 8.06917
R56033 a_83153_n36322.n0 a_83153_n36322.t15 8.06917
R56034 a_83153_n36322.n0 a_83153_n36322.t18 8.06917
R56035 a_83153_n36322.n1 a_83153_n36322.t0 7.94157
R56036 a_83153_n36322.t4 a_83153_n36322.n2 7.72643
R56037 a_83153_n36322.n1 a_83153_n36322.t1 7.22925
R56038 a_83153_n36322.n2 a_83153_n36322.t7 7.17912
R56039 a_83153_n36322.n0 a_83153_n36322.t14 8.33554
R56040 a_83153_n36322.t12 a_83153_n36322.n0 8.33554
R56041 a_83153_n36322.n0 a_83153_n36322.t19 8.33647
R56042 a_83153_n36322.t21 a_83153_n36322.n0 8.33647
R56043 a_83153_n36322.n2 a_83153_n36322.n1 7.46075
R56044 a_83153_10448.t1 a_83153_10448.t7 12.7127
R56045 a_83153_10448.t1 a_83153_10448.t8 10.2828
R56046 a_83153_10448.t1 a_83153_10448.t10 10.2828
R56047 a_83153_10448.t1 a_83153_10448.t17 10.2828
R56048 a_83153_10448.t1 a_83153_10448.t12 10.2828
R56049 a_83153_10448.t1 a_83153_10448.t20 10.1333
R56050 a_83153_10448.t1 a_83153_10448.t21 10.1333
R56051 a_83153_10448.t1 a_83153_10448.t6 10.1333
R56052 a_83153_10448.t1 a_83153_10448.t4 10.1333
R56053 a_83153_10448.t1 a_83153_10448.t2 9.72545
R56054 a_83153_10448.t1 a_83153_10448.t19 9.57156
R56055 a_83153_10448.t1 a_83153_10448.t15 9.57156
R56056 a_83153_10448.t1 a_83153_10448.t16 9.57156
R56057 a_83153_10448.t1 a_83153_10448.t23 9.57156
R56058 a_83153_10448.t1 a_83153_10448.t18 9.57156
R56059 a_83153_10448.t1 a_83153_10448.t13 9.57156
R56060 a_83153_10448.t1 a_83153_10448.t14 9.57156
R56061 a_83153_10448.t1 a_83153_10448.t22 9.57156
R56062 a_83153_10448.t2 a_83153_10448.t3 8.02945
R56063 a_83153_10448.t1 a_83153_10448.t0 8.02708
R56064 a_83153_10448.t1 a_83153_10448.t11 7.90829
R56065 a_83153_10448.t1 a_83153_10448.t9 7.90829
R56066 a_83153_10448.t5 a_83153_10448.t1 7.41776
R56067 a_47819_11614.n2 a_47819_11614.t12 12.8637
R56068 a_47819_11614.t0 a_47819_11614.n1 10.7018
R56069 a_47819_11614.n1 a_47819_11614.t4 10.1659
R56070 a_47819_11614.n1 a_47819_11614.t6 9.64387
R56071 a_47819_11614.n1 a_47819_11614.t3 9.27665
R56072 a_47819_11614.n1 a_47819_11614.n2 8.75198
R56073 a_47819_11614.n2 a_47819_11614.t23 8.14051
R56074 a_47819_11614.n2 a_47819_11614.t19 8.14051
R56075 a_47819_11614.n2 a_47819_11614.t17 8.14051
R56076 a_47819_11614.n2 a_47819_11614.t10 8.14051
R56077 a_47819_11614.n2 a_47819_11614.t14 8.06917
R56078 a_47819_11614.n2 a_47819_11614.t11 8.06917
R56079 a_47819_11614.n2 a_47819_11614.t20 8.06917
R56080 a_47819_11614.n2 a_47819_11614.t8 8.06917
R56081 a_47819_11614.n2 a_47819_11614.t22 8.06917
R56082 a_47819_11614.n2 a_47819_11614.t16 8.06917
R56083 a_47819_11614.n2 a_47819_11614.t18 8.06917
R56084 a_47819_11614.n0 a_47819_11614.t7 7.94068
R56085 a_47819_11614.n1 a_47819_11614.t1 7.72524
R56086 a_47819_11614.n0 a_47819_11614.t5 7.22855
R56087 a_47819_11614.n1 a_47819_11614.t2 7.17942
R56088 a_47819_11614.t9 a_47819_11614.n2 8.33649
R56089 a_47819_11614.n2 a_47819_11614.t13 8.33649
R56090 a_47819_11614.t15 a_47819_11614.n2 8.33556
R56091 a_47819_11614.n2 a_47819_11614.t21 8.33556
R56092 a_47819_11614.n1 a_47819_11614.n0 7.46075
R56093 a_47991_4421.t2 a_47991_4421.t0 21.6693
R56094 a_47991_4421.t1 a_47991_4421.t0 15.3476
R56095 a_57977_n5344.t0 a_57977_n5344.t1 13.2434
R56096 a_103997_n8770.t0 a_103997_n8770.n3 39.3605
R56097 a_103997_n8770.n1 a_103997_n8770.n0 10.9327
R56098 a_103997_n8770.n0 a_103997_n8770.t12 8.44198
R56099 a_103997_n8770.n0 a_103997_n8770.t8 8.44198
R56100 a_103997_n8770.n1 a_103997_n8770.t11 8.44198
R56101 a_103997_n8770.n1 a_103997_n8770.t7 8.44198
R56102 a_103997_n8770.n0 a_103997_n8770.t5 9.26917
R56103 a_103997_n8770.n1 a_103997_n8770.t6 8.10567
R56104 a_103997_n8770.n3 a_103997_n8770.t1 6.51122
R56105 a_103997_n8770.n3 a_103997_n8770.n0 6.50622
R56106 a_103997_n8770.t1 a_103997_n8770.t2 6.36267
R56107 a_103997_n8770.t1 a_103997_n8770.n2 4.84877
R56108 a_103997_n8770.n2 a_103997_n8770.t4 3.65383
R56109 a_103997_n8770.n1 a_103997_n8770.t10 8.65827
R56110 a_103997_n8770.n2 a_103997_n8770.t3 3.57094
R56111 a_103997_n8770.n0 a_103997_n8770.t9 8.77499
R56112 a_47991_5507.t0 a_47991_5507.t2 24.9014
R56113 a_47991_5507.t0 a_47991_5507.t1 15.5881
R56114 a_48951_4481.t0 a_48951_4481.t1 26.1287
R56115 a_48951_4481.t1 a_48951_4481.t2 15.0742
R56116 a_47991_n29313.t0 a_47991_n29313.t1 23.2303
R56117 a_47991_n29313.t0 a_47991_n29313.t2 21.6695
R56118 a_59558_n29181.n0 a_59558_n29181.t11 10.2515
R56119 a_59558_n29181.n1 a_59558_n29181.t2 10.2515
R56120 a_59558_n29181.n0 a_59558_n29181.t17 10.2515
R56121 a_59558_n29181.n0 a_59558_n29181.t0 10.2515
R56122 a_59558_n29181.n0 a_59558_n29181.t4 10.096
R56123 a_59558_n29181.n1 a_59558_n29181.t18 10.0935
R56124 a_59558_n29181.n0 a_59558_n29181.t6 10.0859
R56125 a_59558_n29181.n0 a_59558_n29181.t12 10.0808
R56126 a_59558_n29181.n0 a_59558_n29181.t22 9.53981
R56127 a_59558_n29181.n1 a_59558_n29181.t20 9.53981
R56128 a_59558_n29181.n0 a_59558_n29181.t14 9.53981
R56129 a_59558_n29181.n0 a_59558_n29181.t16 9.53981
R56130 a_59558_n29181.n0 a_59558_n29181.t21 9.53744
R56131 a_59558_n29181.n1 a_59558_n29181.t19 9.53744
R56132 a_59558_n29181.n0 a_59558_n29181.t13 9.53744
R56133 a_59558_n29181.n0 a_59558_n29181.t15 9.53744
R56134 a_59558_n29181.n1 a_59558_n29181.n0 9.16839
R56135 a_59558_n29181.n1 a_59558_n29181.t1 8.14051
R56136 a_59558_n29181.n1 a_59558_n29181.t3 8.13798
R56137 a_59558_n29181.t8 a_59558_n29181.t10 7.95997
R56138 a_59558_n29181.t8 a_59558_n29181.t9 7.94576
R56139 a_59558_n29181.t8 a_59558_n29181.n1 7.50666
R56140 a_59558_n29181.n1 a_59558_n29181.t5 7.48675
R56141 a_59558_n29181.n1 a_59558_n29181.t7 7.48422
R56142 a_53675_n30339.n0 a_53675_n30339.t3 10.3838
R56143 a_53675_n30339.n0 a_53675_n30339.t1 10.3566
R56144 a_53675_n30339.n0 a_53675_n30339.t0 10.0407
R56145 a_53675_n30339.t2 a_53675_n30339.n0 9.57605
R56146 a_60677_n36322.t0 a_60677_n36322.t1 83.5159
R56147 a_60677_n36322.t1 a_60677_n36322.t3 9.77323
R56148 a_60677_n36322.t1 a_60677_n36322.t2 8.17727
R56149 a_65486_11614.n2 a_65486_11614.t23 12.8637
R56150 a_65486_11614.n1 a_65486_11614.t1 10.7018
R56151 a_65486_11614.n1 a_65486_11614.t6 10.1659
R56152 a_65486_11614.n1 a_65486_11614.t4 9.64387
R56153 a_65486_11614.t0 a_65486_11614.n1 9.27665
R56154 a_65486_11614.n1 a_65486_11614.n2 8.75198
R56155 a_65486_11614.n2 a_65486_11614.t18 8.14051
R56156 a_65486_11614.n2 a_65486_11614.t14 8.14051
R56157 a_65486_11614.n2 a_65486_11614.t10 8.14051
R56158 a_65486_11614.n2 a_65486_11614.t22 8.14051
R56159 a_65486_11614.n2 a_65486_11614.t15 8.06917
R56160 a_65486_11614.n2 a_65486_11614.t11 8.06917
R56161 a_65486_11614.n2 a_65486_11614.t16 8.06917
R56162 a_65486_11614.n2 a_65486_11614.t20 8.06917
R56163 a_65486_11614.n2 a_65486_11614.t8 8.06917
R56164 a_65486_11614.n2 a_65486_11614.t19 8.06917
R56165 a_65486_11614.n2 a_65486_11614.t12 8.06917
R56166 a_65486_11614.n0 a_65486_11614.t7 7.94068
R56167 a_65486_11614.n1 a_65486_11614.t2 7.72524
R56168 a_65486_11614.n0 a_65486_11614.t5 7.22855
R56169 a_65486_11614.n1 a_65486_11614.t3 7.17942
R56170 a_65486_11614.t13 a_65486_11614.n2 8.33649
R56171 a_65486_11614.n2 a_65486_11614.t17 8.33649
R56172 a_65486_11614.t21 a_65486_11614.n2 8.33556
R56173 a_65486_11614.n2 a_65486_11614.t9 8.33556
R56174 a_65486_11614.n1 a_65486_11614.n0 7.46075
R56175 a_53829_10388.n5 a_53829_10388.n1 10.2377
R56176 a_53829_10388.n4 a_53829_10388.t3 10.2108
R56177 a_53829_10388.n4 a_53829_10388.t1 9.99909
R56178 a_53829_10388.n5 a_53829_10388.t7 9.80443
R56179 a_53829_10388.n5 a_53829_10388.t5 9.55135
R56180 a_53829_10388.n0 a_53829_10388.t16 8.17385
R56181 a_53829_10388.n3 a_53829_10388.t9 8.17299
R56182 a_53829_10388.n3 a_53829_10388.t10 8.17134
R56183 a_53829_10388.n0 a_53829_10388.t8 8.16754
R56184 a_53829_10388.n1 a_53829_10388.t20 8.10567
R56185 a_53829_10388.n1 a_53829_10388.t19 8.10567
R56186 a_53829_10388.n3 a_53829_10388.t15 8.10567
R56187 a_53829_10388.n3 a_53829_10388.t17 8.10567
R56188 a_53829_10388.n1 a_53829_10388.t18 8.10567
R56189 a_53829_10388.n1 a_53829_10388.t23 8.10567
R56190 a_53829_10388.n0 a_53829_10388.t22 8.10567
R56191 a_53829_10388.n0 a_53829_10388.t13 8.10567
R56192 a_53829_10388.n6 a_53829_10388.t2 7.74799
R56193 a_53829_10388.t4 a_53829_10388.n7 7.73052
R56194 a_53829_10388.n6 a_53829_10388.t0 7.46478
R56195 a_53829_10388.n7 a_53829_10388.t6 7.1311
R56196 a_53829_10388.n4 a_53829_10388.n6 2.2505
R56197 a_53829_10388.n7 a_53829_10388.n5 2.2505
R56198 a_53829_10388.n1 a_53829_10388.t11 8.35731
R56199 a_53829_10388.n0 a_53829_10388.t21 8.38107
R56200 a_53829_10388.n1 a_53829_10388.t12 8.37583
R56201 a_53829_10388.n1 a_53829_10388.n0 4.35656
R56202 a_53829_10388.n5 a_53829_10388.n4 2.96863
R56203 a_53829_10388.n2 a_53829_10388.n1 1.0882
R56204 a_53829_10388.n2 a_53829_10388.n3 1.08408
R56205 a_53829_10388.n2 a_53829_10388.t14 8.66753
R56206 a_53699_13546.n1 a_53699_13546.n0 26.5254
R56207 a_53699_13546.n1 a_53699_13546.t1 11.5094
R56208 a_53699_13546.n0 a_53699_13546.t3 10.937
R56209 a_53699_13546.n0 a_53699_13546.t2 9.33982
R56210 a_53699_13546.t0 a_53699_13546.n1 9.24966
R56211 a_53699_11614.t0 a_53699_11614.t2 58.3955
R56212 a_53699_11614.t0 a_53699_11614.n0 13.0169
R56213 a_53699_11614.n1 a_53699_11614.n0 10.9309
R56214 a_53699_11614.t0 a_53699_11614.t1 8.5021
R56215 a_53699_11614.n1 a_53699_11614.t9 8.44198
R56216 a_53699_11614.n1 a_53699_11614.t3 8.44198
R56217 a_53699_11614.n0 a_53699_11614.t6 8.44198
R56218 a_53699_11614.n0 a_53699_11614.t10 8.44198
R56219 a_53699_11614.n1 a_53699_11614.t4 8.10567
R56220 a_53699_11614.n0 a_53699_11614.t5 9.26955
R56221 a_53699_11614.n1 a_53699_11614.t7 8.65823
R56222 a_53699_11614.n0 a_53699_11614.t8 8.77493
R56223 a_65658_4421.t1 a_65658_4421.t0 21.6693
R56224 a_65658_4421.t2 a_65658_4421.t0 15.3476
R56225 I1N.n8 I1N.t1 10.2879
R56226 I1N.n32 I1N.n31 6.37738
R56227 I1N.t0 I1N.n9 4.39661
R56228 I1N.n7 I1N.t12 4.39661
R56229 I1N.t17 I1N.n1 4.39661
R56230 I1N.t6 I1N.n25 4.39661
R56231 I1N.n10 I1N.t0 4.39661
R56232 I1N.n26 I1N.t6 4.39661
R56233 I1N.n13 I1N.t7 4.39651
R56234 I1N.n12 I1N.t7 4.39651
R56235 I1N.n21 I1N.t4 4.39651
R56236 I1N.n19 I1N.t10 4.39651
R56237 I1N.n29 I1N.t2 4.39651
R56238 I1N.n28 I1N.t2 4.39651
R56239 I1N.n32 I1N.t3 3.9368
R56240 I1N.n13 I1N.t9 2.96638
R56241 I1N.t9 I1N.n12 2.96638
R56242 I1N.t14 I1N.n9 2.96638
R56243 I1N.n10 I1N.t14 2.96638
R56244 I1N.t8 I1N.n1 2.96638
R56245 I1N.n7 I1N.t5 2.96638
R56246 I1N.n21 I1N.t11 2.96638
R56247 I1N.n29 I1N.t16 2.96638
R56248 I1N.t16 I1N.n28 2.96638
R56249 I1N.t13 I1N.n25 2.96638
R56250 I1N.n26 I1N.t13 2.96638
R56251 I1N.t15 I1N.n19 2.96638
R56252 I1N.n6 I1N.t8 2.52844
R56253 I1N.n18 I1N.t4 2.52844
R56254 I1N.t10 I1N.n18 2.52844
R56255 I1N.t5 I1N.n6 2.52844
R56256 I1N.n3 I1N.t12 2.52844
R56257 I1N.n20 I1N.t15 2.52844
R56258 I1N.t11 I1N.n20 2.52844
R56259 I1N.n3 I1N.t17 2.52844
R56260 I1N.n31 I1N.n30 1.5005
R56261 I1N.n27 I1N.n24 1.5005
R56262 I1N.n23 I1N.n22 1.5005
R56263 I1N.n4 I1N.n0 1.5005
R56264 I1N.n17 I1N.n16 1.5005
R56265 I1N.n15 I1N.n14 1.5005
R56266 I1N.n11 I1N.n8 1.5005
R56267 I1N.n5 I1N.n4 1.19221
R56268 I1N.n4 I1N.n2 1.16411
R56269 I1N.n11 I1N.n10 0.88285
R56270 I1N.n14 I1N.n9 0.88285
R56271 I1N.n17 I1N.n7 0.88285
R56272 I1N.n22 I1N.n1 0.88285
R56273 I1N.n27 I1N.n26 0.88285
R56274 I1N.n30 I1N.n25 0.88285
R56275 I1N.n12 I1N.n11 0.858643
R56276 I1N.n14 I1N.n13 0.858643
R56277 I1N.n19 I1N.n17 0.858643
R56278 I1N.n22 I1N.n21 0.858643
R56279 I1N.n28 I1N.n27 0.858643
R56280 I1N.n30 I1N.n29 0.858643
R56281 I1N.n18 I1N.n2 0.367144
R56282 I1N.n5 I1N.n3 0.365787
R56283 I1N.n16 I1N.n0 0.210297
R56284 I1N.n23 I1N.n0 0.207257
R56285 I1N.n31 I1N.n24 0.1805
R56286 I1N.n15 I1N.n8 0.179588
R56287 I1N.n16 I1N.n15 0.0935405
R56288 I1N.n24 I1N.n23 0.0935405
R56289 I1N.n6 I1N.n5 0.0804816
R56290 I1N.n20 I1N.n2 0.0795377
R56291 I1N I1N.n32 0.0159334
R56292 a_89715_n16810.t0 a_89715_n16810.t1 12.8122
R56293 a_71366_13546.n1 a_71366_13546.n0 26.5281
R56294 a_71366_13546.n0 a_71366_13546.t3 11.5094
R56295 a_71366_13546.t0 a_71366_13546.n1 10.937
R56296 a_71366_13546.n1 a_71366_13546.t1 9.33982
R56297 a_71366_13546.n0 a_71366_13546.t2 9.24966
R56298 a_36162_n36382.n6 a_36162_n36382.n1 10.2377
R56299 a_36162_n36382.n5 a_36162_n36382.t7 10.2105
R56300 a_36162_n36382.n5 a_36162_n36382.t5 9.99998
R56301 a_36162_n36382.t0 a_36162_n36382.n6 9.80432
R56302 a_36162_n36382.n6 a_36162_n36382.t3 9.55206
R56303 a_36162_n36382.n0 a_36162_n36382.t22 8.17385
R56304 a_36162_n36382.n3 a_36162_n36382.t20 8.17299
R56305 a_36162_n36382.n3 a_36162_n36382.t23 8.17134
R56306 a_36162_n36382.n0 a_36162_n36382.t21 8.16754
R56307 a_36162_n36382.n1 a_36162_n36382.t9 8.10567
R56308 a_36162_n36382.n1 a_36162_n36382.t17 8.10567
R56309 a_36162_n36382.n3 a_36162_n36382.t15 8.10567
R56310 a_36162_n36382.n3 a_36162_n36382.t8 8.10567
R56311 a_36162_n36382.n1 a_36162_n36382.t12 8.10567
R56312 a_36162_n36382.n1 a_36162_n36382.t16 8.10567
R56313 a_36162_n36382.n0 a_36162_n36382.t14 8.10567
R56314 a_36162_n36382.n0 a_36162_n36382.t10 8.10567
R56315 a_36162_n36382.n7 a_36162_n36382.t4 7.74888
R56316 a_36162_n36382.n4 a_36162_n36382.t2 7.73141
R56317 a_36162_n36382.n7 a_36162_n36382.t6 7.46359
R56318 a_36162_n36382.n4 a_36162_n36382.t1 7.13181
R56319 a_36162_n36382.n6 a_36162_n36382.n4 2.2505
R56320 a_36162_n36382.n5 a_36162_n36382.n7 2.2505
R56321 a_36162_n36382.t13 a_36162_n36382.n1 8.35729
R56322 a_36162_n36382.n1 a_36162_n36382.t11 8.37586
R56323 a_36162_n36382.n0 a_36162_n36382.t18 8.38104
R56324 a_36162_n36382.n1 a_36162_n36382.n0 4.35658
R56325 a_36162_n36382.n6 a_36162_n36382.n5 2.96863
R56326 a_36162_n36382.n2 a_36162_n36382.n1 1.08819
R56327 a_36162_n36382.n2 a_36162_n36382.n3 1.08408
R56328 a_36162_n36382.n2 a_36162_n36382.t19 8.6675
R56329 a_71342_7563.t2 a_71342_7563.n0 10.3829
R56330 a_71342_7563.n0 a_71342_7563.t0 10.3566
R56331 a_71342_7563.n0 a_71342_7563.t1 10.0407
R56332 a_71342_7563.n0 a_71342_7563.t3 9.57605
R56333 a_71366_11614.n1 a_71366_11614.t2 42.1702
R56334 a_71366_11614.t1 a_71366_11614.n1 11.3595
R56335 a_71366_11614.n2 a_71366_11614.n0 10.9309
R56336 a_71366_11614.n2 a_71366_11614.t7 8.44198
R56337 a_71366_11614.n2 a_71366_11614.t3 8.44198
R56338 a_71366_11614.n0 a_71366_11614.t4 8.44198
R56339 a_71366_11614.n0 a_71366_11614.t10 8.44198
R56340 a_71366_11614.n2 a_71366_11614.t5 8.10567
R56341 a_71366_11614.n0 a_71366_11614.t6 9.26955
R56342 a_71366_11614.n1 a_71366_11614.n0 6.50622
R56343 a_71366_11614.n2 a_71366_11614.t8 8.65823
R56344 a_71366_11614.t0 a_71366_11614.t1 3.57094
R56345 a_71366_11614.n0 a_71366_11614.t9 8.77493
R56346 a_78344_10448.t0 a_78344_10448.t4 44.9824
R56347 a_78344_10448.t0 a_78344_10448.t2 13.8923
R56348 a_78344_10448.t0 a_78344_10448.t3 10.1307
R56349 a_78344_10448.t0 a_78344_10448.t1 8.54643
R56350 a_38097_n16007.t0 a_38097_n16007.t2 41.3378
R56351 a_38097_n16007.t2 a_38097_n16007.t1 18.4133
R56352 a_53675_4481.n0 a_53675_4481.t0 10.6581
R56353 a_53675_4481.n0 a_53675_4481.t3 10.2356
R56354 a_53675_4481.t2 a_53675_4481.n0 9.5019
R56355 a_53675_4481.n0 a_53675_4481.t1 9.34796
R56356 a_36162_10388.n5 a_36162_10388.n1 10.2377
R56357 a_36162_10388.n4 a_36162_10388.t2 10.2108
R56358 a_36162_10388.n4 a_36162_10388.t3 9.99909
R56359 a_36162_10388.n5 a_36162_10388.t5 9.80443
R56360 a_36162_10388.n5 a_36162_10388.t7 9.55135
R56361 a_36162_10388.n0 a_36162_10388.t20 8.17385
R56362 a_36162_10388.n3 a_36162_10388.t16 8.17299
R56363 a_36162_10388.n3 a_36162_10388.t17 8.17134
R56364 a_36162_10388.n0 a_36162_10388.t15 8.16754
R56365 a_36162_10388.n1 a_36162_10388.t14 8.10567
R56366 a_36162_10388.n1 a_36162_10388.t11 8.10567
R56367 a_36162_10388.n3 a_36162_10388.t9 8.10567
R56368 a_36162_10388.n3 a_36162_10388.t13 8.10567
R56369 a_36162_10388.n1 a_36162_10388.t10 8.10567
R56370 a_36162_10388.n1 a_36162_10388.t19 8.10567
R56371 a_36162_10388.n0 a_36162_10388.t18 8.10567
R56372 a_36162_10388.n0 a_36162_10388.t8 8.10567
R56373 a_36162_10388.n6 a_36162_10388.t1 7.74799
R56374 a_36162_10388.n7 a_36162_10388.t6 7.73052
R56375 a_36162_10388.n6 a_36162_10388.t0 7.46478
R56376 a_36162_10388.t4 a_36162_10388.n7 7.1311
R56377 a_36162_10388.n4 a_36162_10388.n6 2.2505
R56378 a_36162_10388.n7 a_36162_10388.n5 2.2505
R56379 a_36162_10388.n1 a_36162_10388.t21 8.35731
R56380 a_36162_10388.n0 a_36162_10388.t12 8.38107
R56381 a_36162_10388.n1 a_36162_10388.t22 8.37583
R56382 a_36162_10388.n1 a_36162_10388.n0 4.35656
R56383 a_36162_10388.n5 a_36162_10388.n4 2.96863
R56384 a_36162_10388.n2 a_36162_10388.n1 1.0882
R56385 a_36162_10388.n2 a_36162_10388.n3 1.08408
R56386 a_36162_10388.n2 a_36162_10388.t23 8.66753
R56387 a_32913_n5342.t0 a_32913_n5342.t1 13.2434
R56388 a_65658_n29313.t0 a_65658_n29313.t1 23.2303
R56389 a_65658_n29313.t0 a_65658_n29313.t2 21.6695
R56390 a_39179_n16007.t0 a_39179_n16007.t1 13.2434
R56391 a_71366_n36322.n1 a_71366_n36322.n0 26.5281
R56392 a_71366_n36322.n0 a_71366_n36322.t2 11.5094
R56393 a_71366_n36322.n1 a_71366_n36322.t1 10.937
R56394 a_71366_n36322.t0 a_71366_n36322.n1 9.33982
R56395 a_71366_n36322.n0 a_71366_n36322.t3 9.24966
R56396 a_30324_5507.t0 a_30324_5507.t1 30.2725
R56397 a_30324_5507.t1 a_30324_5507.t2 24.9014
R56398 a_71342_n27257.n0 a_71342_n27257.t0 10.6581
R56399 a_71342_n27257.n0 a_71342_n27257.t3 10.2358
R56400 a_71342_n27257.t2 a_71342_n27257.n0 9.50202
R56401 a_71342_n27257.n0 a_71342_n27257.t1 9.34796
R56402 a_50629_n16009.t1 a_50629_n16009.t2 82.9933
R56403 a_50629_n16009.t0 a_50629_n16009.t1 17.244
R56404 a_39179_n8930.t0 a_39179_n8930.t1 118.243
R56405 a_39179_n8930.t1 a_39179_n8930.t2 24.9025
R56406 a_106676_7563.t2 a_106676_7563.n0 10.3829
R56407 a_106676_7563.n0 a_106676_7563.t0 10.3566
R56408 a_106676_7563.n0 a_106676_7563.t1 10.0407
R56409 a_106676_7563.n0 a_106676_7563.t3 9.57605
R56410 a_106830_n36382.n5 a_106830_n36382.n1 10.2377
R56411 a_106830_n36382.n4 a_106830_n36382.t2 10.2105
R56412 a_106830_n36382.n4 a_106830_n36382.t1 9.99998
R56413 a_106830_n36382.n5 a_106830_n36382.t5 9.80532
R56414 a_106830_n36382.n5 a_106830_n36382.t7 9.55206
R56415 a_106830_n36382.n0 a_106830_n36382.t20 8.17385
R56416 a_106830_n36382.n3 a_106830_n36382.t16 8.17299
R56417 a_106830_n36382.n3 a_106830_n36382.t21 8.17134
R56418 a_106830_n36382.n0 a_106830_n36382.t17 8.16754
R56419 a_106830_n36382.n1 a_106830_n36382.t18 8.10567
R56420 a_106830_n36382.n1 a_106830_n36382.t23 8.10567
R56421 a_106830_n36382.n3 a_106830_n36382.t15 8.10567
R56422 a_106830_n36382.n3 a_106830_n36382.t10 8.10567
R56423 a_106830_n36382.n1 a_106830_n36382.t19 8.10567
R56424 a_106830_n36382.n1 a_106830_n36382.t22 8.10567
R56425 a_106830_n36382.n0 a_106830_n36382.t14 8.10567
R56426 a_106830_n36382.n0 a_106830_n36382.t13 8.10567
R56427 a_106830_n36382.n6 a_106830_n36382.t3 7.74888
R56428 a_106830_n36382.n7 a_106830_n36382.t6 7.73141
R56429 a_106830_n36382.n6 a_106830_n36382.t0 7.46359
R56430 a_106830_n36382.t4 a_106830_n36382.n7 7.13081
R56431 a_106830_n36382.n4 a_106830_n36382.n6 2.2505
R56432 a_106830_n36382.n7 a_106830_n36382.n5 2.2505
R56433 a_106830_n36382.t9 a_106830_n36382.n1 8.35729
R56434 a_106830_n36382.n1 a_106830_n36382.t8 8.37586
R56435 a_106830_n36382.n0 a_106830_n36382.t11 8.38104
R56436 a_106830_n36382.n1 a_106830_n36382.n0 4.35658
R56437 a_106830_n36382.n5 a_106830_n36382.n4 2.96863
R56438 a_106830_n36382.n2 a_106830_n36382.n1 1.08819
R56439 a_106830_n36382.n2 a_106830_n36382.n3 1.08408
R56440 a_106830_n36382.n2 a_106830_n36382.t12 8.6675
R56441 a_36008_7563.t0 a_36008_7563.n0 10.3829
R56442 a_36008_7563.n0 a_36008_7563.t3 10.3566
R56443 a_36008_7563.n0 a_36008_7563.t2 10.0407
R56444 a_36008_7563.n0 a_36008_7563.t1 9.57605
R56445 a_89009_7563.n0 a_89009_7563.t3 10.3829
R56446 a_89009_7563.n0 a_89009_7563.t1 10.3566
R56447 a_89009_7563.n0 a_89009_7563.t0 10.0407
R56448 a_89009_7563.t2 a_89009_7563.n0 9.57605
R56449 a_36032_13546.n1 a_36032_13546.n0 26.5241
R56450 a_36032_13546.n1 a_36032_13546.t1 11.5094
R56451 a_36032_13546.n0 a_36032_13546.t3 10.937
R56452 a_36032_13546.n0 a_36032_13546.t2 9.33982
R56453 a_36032_13546.t0 a_36032_13546.n1 9.24966
R56454 a_101111_n6055.t0 a_101111_n6055.t1 12.8122
R56455 IN_POS.n32 IN_POS.n31 17.0316
R56456 IN_POS.n15 IN_POS.n1 3.06497
R56457 IN_POS.n27 IN_POS.n0 2.80204
R56458 IN_POS.n23 IN_POS.n22 2.55189
R56459 IN_POS.n29 IN_POS.n28 2.44888
R56460 IN_POS.n13 IN_POS.n12 2.44888
R56461 IN_POS.n11 IN_POS.n10 2.44888
R56462 IN_POS.n17 IN_POS.n16 2.44888
R56463 IN_POS.n20 IN_POS.n19 2.44888
R56464 IN_POS.n25 IN_POS.n24 2.44888
R56465 IN_POS IN_POS.n32 2.30113
R56466 IN_POS IN_POS.n32 2.27938
R56467 IN_POS.n31 IN_POS.n0 1.75374
R56468 IN_POS.t0 IN_POS.n8 1.1935
R56469 IN_POS.t0 IN_POS.n18 1.19272
R56470 IN_POS.n23 IN_POS.n9 1.18175
R56471 IN_POS.n27 IN_POS.t0 1.0998
R56472 IN_POS.t0 IN_POS.n15 1.08916
R56473 IN_POS.n28 IN_POS.n27 0.958371
R56474 IN_POS.n17 IN_POS.n15 0.907386
R56475 IN_POS.t0 IN_POS.n9 0.752643
R56476 IN_POS.n13 IN_POS.n8 0.706267
R56477 IN_POS.n20 IN_POS.n18 0.672835
R56478 IN_POS.n16 IN_POS.n1 0.66672
R56479 IN_POS.t0 IN_POS.n14 0.629953
R56480 IN_POS.n30 IN_POS.n29 0.622487
R56481 IN_POS.t0 IN_POS.n21 0.604576
R56482 IN_POS.n25 IN_POS.n21 0.585642
R56483 IN_POS.n14 IN_POS.n11 0.583689
R56484 IN_POS.n21 IN_POS.n20 0.559641
R56485 IN_POS.n26 IN_POS.n25 0.549445
R56486 IN_POS.n28 IN_POS.n8 0.540673
R56487 IN_POS.n14 IN_POS.n13 0.529423
R56488 IN_POS.n18 IN_POS.n17 0.519089
R56489 IN_POS.n12 IN_POS.n7 0.514976
R56490 IN_POS.n19 IN_POS.n4 0.499862
R56491 IN_POS.t1 IN_POS.n30 0.47657
R56492 IN_POS.n30 IN_POS.n0 0.424689
R56493 IN_POS.n29 IN_POS.n7 0.383261
R56494 IN_POS.n16 IN_POS.n4 0.36773
R56495 IN_POS.n10 IN_POS.n6 0.365351
R56496 IN_POS.n24 IN_POS.n3 0.362981
R56497 IN_POS.n19 IN_POS.n3 0.348693
R56498 IN_POS.n12 IN_POS.n6 0.337682
R56499 IN_POS.t1 IN_POS.n1 0.323064
R56500 IN_POS.t1 IN_POS.n4 0.304037
R56501 IN_POS.t1 IN_POS.n7 0.300094
R56502 IN_POS.n10 IN_POS.n5 0.256772
R56503 IN_POS.n24 IN_POS.n2 0.246737
R56504 IN_POS.t1 IN_POS.n6 0.136362
R56505 IN_POS.t1 IN_POS.n3 0.128975
R56506 IN_POS.n11 IN_POS.n9 0.104562
R56507 IN_POS.n22 IN_POS.n2 0.0290825
R56508 IN_POS.n22 IN_POS.n5 0.0207691
R56509 IN_POS.n26 IN_POS.n23 0.00666077
R56510 IN_POS.t1 IN_POS.n2 0.00482948
R56511 IN_POS.t0 IN_POS.n26 0.00449532
R56512 IN_POS.t1 IN_POS.n5 0.00410811
R56513 IN_POS.n31 IN_POS.t1 0.00330619
R56514 a_94892_4481.n1 a_94892_4481.t4 10.2515
R56515 a_94892_4481.n1 a_94892_4481.t0 10.2515
R56516 a_94892_4481.n1 a_94892_4481.t14 10.2515
R56517 a_94892_4481.n1 a_94892_4481.t20 10.2515
R56518 a_94892_4481.n1 a_94892_4481.t2 10.096
R56519 a_94892_4481.n1 a_94892_4481.t13 10.0935
R56520 a_94892_4481.n1 a_94892_4481.t6 10.0859
R56521 a_94892_4481.n1 a_94892_4481.t19 10.0808
R56522 a_94892_4481.n1 a_94892_4481.t22 9.53981
R56523 a_94892_4481.n1 a_94892_4481.t18 9.53981
R56524 a_94892_4481.n1 a_94892_4481.t12 9.53981
R56525 a_94892_4481.n1 a_94892_4481.t16 9.53981
R56526 a_94892_4481.n1 a_94892_4481.t21 9.53744
R56527 a_94892_4481.n1 a_94892_4481.t17 9.53744
R56528 a_94892_4481.n1 a_94892_4481.t11 9.53744
R56529 a_94892_4481.n1 a_94892_4481.t15 9.53744
R56530 a_94892_4481.n1 a_94892_4481.n0 8.41434
R56531 a_94892_4481.n1 a_94892_4481.t5 8.14082
R56532 a_94892_4481.n0 a_94892_4481.t1 8.13828
R56533 a_94892_4481.t8 a_94892_4481.t9 7.96115
R56534 a_94892_4481.t8 a_94892_4481.t10 7.94694
R56535 a_94892_4481.t8 a_94892_4481.n1 7.50666
R56536 a_94892_4481.n0 a_94892_4481.t3 7.48586
R56537 a_94892_4481.n1 a_94892_4481.t7 7.48333
R56538 a_89033_n36322.n1 a_89033_n36322.n0 26.5215
R56539 a_89033_n36322.n0 a_89033_n36322.t3 11.5094
R56540 a_89033_n36322.n1 a_89033_n36322.t1 10.937
R56541 a_89033_n36322.t0 a_89033_n36322.n1 9.33982
R56542 a_89033_n36322.n0 a_89033_n36322.t2 9.24966
R56543 a_53675_n27257.n0 a_53675_n27257.t1 10.6581
R56544 a_53675_n27257.t2 a_53675_n27257.n0 10.2348
R56545 a_53675_n27257.n0 a_53675_n27257.t3 9.50202
R56546 a_53675_n27257.n0 a_53675_n27257.t0 9.34796
R56547 a_51711_n16009.t0 a_51711_n16009.t1 13.2434
R56548 a_89715_n5150.t0 a_89715_n5150.t1 12.8122
R56549 a_64243_n5344.t0 a_64243_n5344.t1 13.2434
R56550 a_89009_4481.n0 a_89009_4481.t0 10.6581
R56551 a_89009_4481.t2 a_89009_4481.n0 10.2346
R56552 a_89009_4481.n0 a_89009_4481.t3 9.5029
R56553 a_89009_4481.n0 a_89009_4481.t1 9.34796
R56554 a_39179_n5342.t0 a_39179_n5342.t1 13.2434
R56555 a_106809_n6055.t0 a_106809_n6055.t1 12.8114
R56556 VCM.n1 VCM.t1 11.5094
R56557 VCM.n2 VCM.n1 10.2743
R56558 VCM.n1 VCM.t0 9.24966
R56559 VCM VCM.n2 4.98085
R56560 VCM.n2 VCM.n0 4.18387
R56561 VCM.n0 VCM.t2 0.111029
R56562 VCM.n0 VCM.t3 0.03175
R56563 a_36008_n30339.t0 a_36008_n30339.n0 10.3838
R56564 a_36008_n30339.n0 a_36008_n30339.t3 10.3566
R56565 a_36008_n30339.n0 a_36008_n30339.t2 10.0407
R56566 a_36008_n30339.n0 a_36008_n30339.t1 9.57605
R56567 a_89009_n30339.t2 a_89009_n30339.n0 10.3838
R56568 a_89009_n30339.n0 a_89009_n30339.t0 10.3566
R56569 a_89009_n30339.n0 a_89009_n30339.t1 10.0407
R56570 a_89009_n30339.n0 a_89009_n30339.t3 9.57605
R56571 a_112507_n17715.t0 a_112507_n17715.t1 12.8114
R56572 a_53675_7563.t2 a_53675_7563.n0 10.3829
R56573 a_53675_7563.n0 a_53675_7563.t1 10.3566
R56574 a_53675_7563.n0 a_53675_7563.t0 10.0407
R56575 a_53675_7563.n0 a_53675_7563.t3 9.57605
R56576 a_45445_n5342.t0 a_45445_n5342.t1 13.2434
R56577 a_43010_n36322.t2 a_43010_n36322.t3 99.46
R56578 a_43010_n36322.t2 a_43010_n36322.t1 9.77323
R56579 a_43010_n36322.t0 a_43010_n36322.t2 8.17727
R56580 a_64243_n16009.t0 a_64243_n16009.t1 13.2434
R56581 a_57977_n16009.t0 a_57977_n16009.t1 13.2434
R56582 a_36008_n27257.n0 a_36008_n27257.t2 10.6581
R56583 a_36008_n27257.t0 a_36008_n27257.n0 10.2348
R56584 a_36008_n27257.n0 a_36008_n27257.t1 9.50202
R56585 a_36008_n27257.n0 a_36008_n27257.t3 9.34796
R56586 a_71266_n4019.t1 a_71266_n4019.t0 9.72448
R56587 a_84017_n5150.t0 a_84017_n5150.t1 12.8114
R56588 a_106676_n27257.n0 a_106676_n27257.t0 10.6581
R56589 a_106676_n27257.n0 a_106676_n27257.t3 10.2358
R56590 a_106676_n27257.t2 a_106676_n27257.n0 9.50202
R56591 a_106676_n27257.n0 a_106676_n27257.t1 9.34796
R56592 a_95413_n5150.t0 a_95413_n5150.t1 12.8114
R56593 a_112507_n6055.t0 a_112507_n6055.t1 12.8114
R56594 a_95413_n16810.t0 a_95413_n16810.t1 12.8114
R56595 a_32913_n16007.t0 a_32913_n16007.t1 13.2434
R56596 a_45445_n16007.t0 a_45445_n16007.t1 13.2434
R56597 IBPOUT IBPOUT.t0 3.31278
R56598 a_84017_n16810.t0 a_84017_n16810.t1 12.8114
R56599 IN_NEG.n30 IN_NEG.t0 24.6019
R56600 IN_NEG.n8 IN_NEG.n0 3.09085
R56601 IN_NEG.n29 IN_NEG.n7 3.06463
R56602 IN_NEG.n19 IN_NEG.n18 2.55189
R56603 IN_NEG.n13 IN_NEG.n12 2.44888
R56604 IN_NEG.n10 IN_NEG.n9 2.44888
R56605 IN_NEG.n22 IN_NEG.n21 2.44888
R56606 IN_NEG.n25 IN_NEG.n24 2.44888
R56607 IN_NEG.n28 IN_NEG.n27 2.44888
R56608 IN_NEG.n16 IN_NEG.n15 2.44888
R56609 IN_NEG IN_NEG.n30 2.29437
R56610 IN_NEG IN_NEG.n30 2.28612
R56611 IN_NEG.t0 IN_NEG.n1 1.1935
R56612 IN_NEG.t0 IN_NEG.n6 1.19272
R56613 IN_NEG.t0 IN_NEG.n0 1.0998
R56614 IN_NEG.t0 IN_NEG.n29 1.08916
R56615 IN_NEG.n9 IN_NEG.n0 0.958371
R56616 IN_NEG.n29 IN_NEG.n28 0.907386
R56617 IN_NEG.n12 IN_NEG.n1 0.706267
R56618 IN_NEG.n10 IN_NEG.n8 0.694516
R56619 IN_NEG.n24 IN_NEG.n6 0.672835
R56620 IN_NEG.n27 IN_NEG.n7 0.66725
R56621 IN_NEG.t0 IN_NEG.n2 0.629953
R56622 IN_NEG.t0 IN_NEG.n5 0.604576
R56623 IN_NEG.n21 IN_NEG.n5 0.585642
R56624 IN_NEG.n15 IN_NEG.n2 0.583689
R56625 IN_NEG.n15 IN_NEG.n3 0.563066
R56626 IN_NEG.n24 IN_NEG.n5 0.559641
R56627 IN_NEG.n9 IN_NEG.n1 0.540673
R56628 IN_NEG.n12 IN_NEG.n2 0.529423
R56629 IN_NEG.n28 IN_NEG.n6 0.519089
R56630 IN_NEG.n13 IN_NEG.n11 0.514976
R56631 IN_NEG.n21 IN_NEG.n4 0.513594
R56632 IN_NEG.n26 IN_NEG.n25 0.500509
R56633 IN_NEG.n11 IN_NEG.n10 0.383261
R56634 IN_NEG.n27 IN_NEG.n26 0.367123
R56635 IN_NEG.n16 IN_NEG.n14 0.365351
R56636 IN_NEG.n23 IN_NEG.n22 0.3637
R56637 IN_NEG.n25 IN_NEG.n23 0.347986
R56638 IN_NEG.n14 IN_NEG.n13 0.337682
R56639 IN_NEG.n8 IN_NEG.t1 0.323963
R56640 IN_NEG.t1 IN_NEG.n7 0.323141
R56641 IN_NEG.n26 IN_NEG.t1 0.304079
R56642 IN_NEG.n11 IN_NEG.t1 0.300094
R56643 IN_NEG.n22 IN_NEG.n20 0.247682
R56644 IN_NEG.n17 IN_NEG.n16 0.229987
R56645 IN_NEG.n19 IN_NEG.n17 0.222212
R56646 IN_NEG.n14 IN_NEG.t1 0.136362
R56647 IN_NEG.n23 IN_NEG.t1 0.129075
R56648 IN_NEG.n18 IN_NEG.n4 0.100573
R56649 IN_NEG.t0 IN_NEG.n4 0.0624826
R56650 IN_NEG.n17 IN_NEG.t1 0.0337966
R56651 IN_NEG.n20 IN_NEG.n19 0.0147343
R56652 IN_NEG.n18 IN_NEG.n3 0.00689777
R56653 IN_NEG.t0 IN_NEG.n3 0.00476406
R56654 IN_NEG.n20 IN_NEG.t1 0.00295152
R56655 IBNOUT IBNOUT.t0 3.42291
R56656 a_101111_n17715.t0 a_101111_n17715.t1 12.8114
C0 a_66016_n35156# a_66016_n36322# 0.004007f
C1 a_34347_n2651# a_35221_n2651# 5.43e-19
C2 a_59411_n2653# a_59763_n3550# 0.053799f
C3 a_57417_n2653# a_57977_n3550# 0.0284f
C4 a_32088_12380# VDD 0.061113f
C5 a_44363_n13316# a_45445_n12419# 5.37e-19
C6 a_75585_n8397# a_75585_n9297# 0.005955f
C7 a_81205_n16810# VDD 1.20767f
C8 a_93969_n19525# a_94537_n19525# 0.027101f
C9 a_92601_n21335# a_93131_n21335# 0.044257f
C10 a_101350_11614# a_101350_10448# 0.004007f
C11 a_34347_n7136# a_35221_n7136# 0.004425f
C12 a_56895_n7138# a_56895_n8932# 0.005987f
C13 a_55635_12380# VDD 0.009062f
C14 a_47753_n15110# a_47753_n16007# 0.005987f
C15 a_45445_n16904# a_44885_n16904# 0.035468f
C16 a_83709_n3340# a_83709_n4245# 0.024773f
C17 a_36562_n34390# VDD 0.009062f
C18 a_31831_n8930# I1U 1.08e-34
C19 a_30377_19942# a_30377_18342# 0.007227f
C20 a_102756_n33224# a_102756_n34390# 0.004007f
C21 a_40613_n2651# a_40053_n2651# 0.0284f
C22 a_64243_n3550# a_64595_n3550# 0.210644f
C23 a_67111_n2653# a_66029_n3550# 5.37e-19
C24 a_79182_11614# VDD 0.011958f
C25 a_66551_n1756# a_66551_n2653# 0.005987f
C26 a_83141_n9675# a_83709_n9675# 0.027101f
C27 a_95943_n15000# VDD 0.39614f
C28 a_30682_10448# I1U 0.005416f
C29 a_111631_n3340# a_111631_n4245# 0.005903f
C30 a_71896_n33224# VDD 0.021515f
C31 a_42413_6405# a_42413_5639# 0.00778f
C32 a_38619_n6239# a_38619_n7136# 0.005987f
C33 a_40613_n7136# a_40053_n7136# 0.037577f
C34 a_38097_n7136# a_39179_n8033# 5.37e-19
C35 a_41487_n6239# a_42047_n7136# 0.0284f
C36 a_67111_n7138# a_66551_n7138# 0.0284f
C37 a_108636_n36322# VCM 0.004624f
C38 a_65677_n7138# a_65677_n8932# 0.01664f
C39 a_51711_n16906# a_51151_n16906# 0.034628f
C40 a_84547_n6960# VDD 1.15365f
C41 a_87433_n6055# a_86903_n9675# 0.03483f
C42 a_98829_n15905# VDD 0.137705f
C43 a_110225_n9675# a_111063_n9675# 0.027101f
C44 a_105933_n15000# a_105933_n15905# 0.005903f
C45 a_102756_n35156# VDD 0.061113f
C46 a_46879_n2651# a_45445_n3548# 1.57e-19
C47 a_72603_n10973# OUT 2.78e-19
C48 a_32913_n12419# a_33787_n12419# 0.001405f
C49 a_94537_n1530# a_95105_n1530# 0.027101f
C50 a_93131_n1530# a_93131_n2435# 0.024773f
C51 a_92601_n5150# a_93969_n2435# 0.002134f
C52 a_87433_n6960# VDD 0.137705f
C53 a_106501_n15905# VDD 0.112244f
C54 a_105933_n20430# a_106501_n20430# 0.027101f
C55 a_47753_n6239# a_48313_n7136# 0.0284f
C56 a_44885_n6239# a_44885_n7136# 0.005987f
C57 a_44363_n7136# a_45445_n8033# 5.37e-19
C58 a_46879_n7136# a_46319_n7136# 0.037577f
C59 a_34699_n16904# a_35781_n17801# 0.002917f
C60 a_60285_n16009# a_59411_n17803# 0.034652f
C61 a_59763_n16906# a_60285_n16906# 0.034714f
C62 a_93131_n6960# a_93131_n7865# 0.024773f
C63 a_93969_n7865# VDD 0.016281f
C64 a_92601_n7865# a_93969_n7865# 2.31e-19
C65 a_87433_n13190# a_88271_n13190# 0.027101f
C66 a_65117_n13318# IBNOUT -8.11e-35
C67 a_111631_n15905# a_113037_n18620# 0.002302f
C68 a_67422_13546# a_67422_12380# 0.004007f
C69 a_53145_n2653# a_51711_n3550# 1.57e-19
C70 a_107198_5639# VDD 0.042519f
C71 a_38619_n12419# a_39179_n12419# 0.0284f
C72 a_100803_n2435# a_101641_n3340# 0.028522f
C73 a_86903_n19525# a_88271_n18620# 2.31e-19
C74 a_111063_n21335# a_111631_n21335# 0.027101f
C75 a_49755_n35156# a_49755_n36322# 0.004007f
C76 a_53145_n7138# a_53497_n8035# 0.16936f
C77 a_64243_n16906# a_64243_n18700# 0.008933f
C78 a_98299_n9675# a_99667_n9675# 7.4e-19
C79 a_105933_n8770# VDD 0.016652f
C80 a_92601_n16810# a_93969_n15000# 0.002134f
C81 a_93131_n14095# a_93969_n14095# 0.027101f
C82 a_73302_n35156# I1N 0.002533f
C83 a_95105_n13190# a_95105_n14095# 0.024773f
C84 a_32353_n17801# I1U 0.002649f
C85 a_34347_n2651# a_34699_n3548# 0.053799f
C86 a_32353_n2651# a_32913_n3548# 0.0284f
C87 a_30682_12380# VDD 0.076387f
C88 a_59411_n2653# a_58851_n2653# 0.0284f
C89 a_44363_n13316# a_44885_n12419# 0.0284f
C90 a_103997_n5150# a_103997_n9675# 0.032645f
C91 a_104527_n3340# a_105365_n3340# 0.027101f
C92 a_107339_n3340# a_106501_n3340# 0.028522f
C93 a_112199_n9675# VDD 0.209912f
C94 a_95105_n18620# a_95105_n19525# 0.024773f
C95 a_83683_n34390# a_83683_n35156# 0.00778f
C96 a_34347_n7136# a_34699_n8033# 0.062551f
C97 a_31831_n7136# a_33265_n8033# 1.57e-19
C98 a_57417_n7138# a_57977_n8035# 0.0284f
C99 a_54229_12380# VDD 0.009062f
C100 a_47231_n16904# a_47753_n16007# 0.005903f
C101 a_45445_n16904# a_44363_n17801# 0.001037f
C102 a_81735_n4245# a_82573_n4245# 0.027101f
C103 a_89407_n13190# VDD 0.150485f
C104 a_105933_n7865# a_105933_n8770# 0.005903f
C105 a_101641_n15000# a_100803_n15000# 0.028522f
C106 a_98829_n15000# a_99667_n15000# 0.027101f
C107 a_98299_n16810# a_98299_n21335# 0.032645f
C108 a_30377_19942# a_31699_19142# 0.009898f
C109 a_66058_n28415# a_66058_n29181# 0.00778f
C110 a_113110_11614# a_113110_10448# 0.004007f
C111 a_40613_n2651# a_39531_n3548# 5.37e-19
C112 a_40053_n1754# a_40053_n2651# 0.005987f
C113 a_38097_n2651# a_38097_n4445# 0.005987f
C114 a_77776_n33224# VCM 0.002508f
C115 a_39179_n1754# a_40965_n3548# 0.006457f
C116 a_77776_11614# VDD 0.017204f
C117 a_65677_n2653# a_66551_n2653# 5.43e-19
C118 a_95105_n14095# VDD 0.180629f
C119 a_67422_n36322# VDD 0.05845f
C120 a_32088_11614# I1U 0.003282f
C121 IBPOUT VCM 0.360724f
C122 a_100235_n19525# a_100235_n20430# 0.005903f
C123 a_38097_n7136# a_38619_n7136# 0.0284f
C124 a_40613_n7136# a_39531_n8033# 0.00117f
C125 a_107230_n36322# VCM 0.02891f
C126 a_66551_n6241# a_66551_n7138# 0.005987f
C127 a_67111_n7138# a_66029_n8035# 5.37e-19
C128 a_102756_10448# VDD 0.05812f
C129 a_64243_n8035# a_64595_n8035# 0.210644f
C130 a_53497_n16906# a_53145_n17803# 0.070243f
C131 a_54019_n15112# a_54019_n16009# 0.005987f
C132 a_51711_n16906# a_50629_n17803# 0.002568f
C133 a_83709_n4245# VDD 0.138244f
C134 a_111631_n8770# a_111631_n9675# 0.005903f
C135 a_100803_n15000# VDD 0.121044f
C136 a_101350_n35156# VDD 0.076387f
C137 a_47753_n1754# a_48313_n2651# 0.0284f
C138 a_56895_n13318# a_57417_n12421# 0.0284f
C139 a_86903_n7865# VDD 0.399575f
C140 a_92601_n5150# a_93131_n2435# 0.012586f
C141 a_105933_n15905# VDD 0.023105f
C142 a_83709_n15905# a_84547_n18620# 0.032618f
C143 a_87433_n3340# IN_POS 0.00603f
C144 a_104527_n20430# a_104527_n21335# 0.024773f
C145 a_46879_n7136# a_45797_n8033# 0.00117f
C146 a_44363_n7136# a_44885_n7136# 0.0284f
C147 a_34699_n16904# a_35221_n16904# 0.035574f
C148 a_93969_n6960# a_94537_n6960# 0.027101f
C149 a_92601_n9675# a_93969_n7865# 0.002134f
C150 a_93131_n7865# VDD 0.121044f
C151 a_95943_n6960# a_95943_n8770# 0.011861f
C152 a_92601_n7865# a_93131_n7865# 0.028522f
C153 a_110225_n17715# VDD 0.41764f
C154 a_86903_n16810# a_88271_n13190# 7.4e-19
C155 a_64595_n14215# IBNOUT 0.002725f
C156 a_110225_n15905# a_110225_n17715# 0.006141f
C157 a_111631_n15905# a_112199_n15905# 0.027101f
C158 a_89531_6405# a_89531_5639# 0.00778f
C159 a_54019_n1756# a_54579_n2653# 0.0284f
C160 a_108602_6405# VDD 0.034176f
C161 a_38097_n13316# a_39179_n12419# 5.37e-19
C162 a_101641_n8770# VDD 0.392932f
C163 a_100235_n2435# a_101641_n3340# 2.31e-19
C164 a_98299_n5150# a_99667_n4245# 0.002134f
C165 a_98829_n2435# a_98829_n3340# 0.024773f
C166 w_27790_n38888# VCM 0.210753f
C167 a_86903_n19525# a_87433_n18620# 0.028522f
C168 a_86903_n21335# a_88271_n18620# 0.002134f
C169 a_112199_n20430# a_112199_n21335# 0.024773f
C170 a_53145_n7138# a_52585_n7138# 0.0284f
C171 a_50629_n7138# a_52063_n8035# 1.57e-19
C172 a_41487_n15110# a_41487_n16007# 0.005987f
C173 a_39179_n16904# a_38619_n16904# 0.035468f
C174 a_63683_n16009# a_63683_n16906# 0.005987f
C175 a_66029_n16906# a_67111_n17803# 0.001641f
C176 a_98299_n9675# a_98829_n9675# 0.032766f
C177 a_99667_n7865# a_100235_n7865# 0.027101f
C178 a_105365_n8770# VDD 0.016652f
C179 a_92601_n16810# a_93131_n15000# 0.012586f
C180 a_67422_n34390# a_67422_n35156# 0.00778f
C181 a_34347_n2651# a_33787_n2651# 0.0284f
C182 a_56895_n2653# a_56895_n4447# 0.005987f
C183 a_59411_n2653# a_58329_n3550# 5.37e-19
C184 a_58851_n1756# a_58851_n2653# 0.005987f
C185 a_32088_13546# VDD 0.05845f
C186 a_72603_n8397# a_72603_n9297# 0.005955f
C187 a_107339_n3340# a_105933_n3340# 2.31e-19
C188 a_111631_n9675# VDD 0.031519f
C189 a_106501_n2435# a_106501_n3340# 0.024773f
C190 a_103997_n4245# a_105365_n3340# 2.31e-19
C191 a_93131_n19525# a_93969_n19525# 0.027101f
C192 a_102756_12380# a_102756_11614# 0.00778f
C193 a_34347_n7136# a_33787_n7136# 0.037577f
C194 a_31831_n7136# a_32913_n8033# 5.37e-19
C195 a_32353_n6239# a_32353_n7136# 0.005987f
C196 a_35221_n6239# a_35781_n7136# 0.0284f
C197 a_59411_n7138# a_60285_n7138# 0.006769f
C198 a_94537_n21335# IBPOUT 0.00243f
C199 a_47231_n16904# a_46879_n17801# 0.534125f
C200 a_46879_n14213# a_48313_n17801# 0.009477f
C201 a_83141_n3340# a_83141_n4245# 0.005903f
C202 a_88839_n13190# VDD 0.02546f
C203 a_37968_n33224# VDD 0.021515f
C204 a_84547_n20430# IN_POS 0.004986f
C205 a_101641_n15000# a_100235_n15000# 2.31e-19
C206 a_100803_n14095# a_100803_n15000# 0.024773f
C207 a_98299_n15905# a_99667_n15000# 2.31e-19
C208 a_101350_n33224# a_101350_n34390# 0.004007f
C209 a_40613_n2651# a_39179_n3548# 1.57e-19
C210 a_63683_n2653# a_64243_n3550# 0.0284f
C211 a_79182_12380# VDD 0.009062f
C212 a_65677_n2653# a_66029_n3550# 0.053799f
C213 a_82573_n9675# a_83141_n9675# 0.027101f
C214 a_111063_n3340# a_111063_n4245# 0.005903f
C215 a_113037_n3340# a_113037_n6960# 0.011861f
C216 a_94537_n14095# VDD 0.022711f
C217 a_30682_11614# I1U 0.005416f
C218 a_66016_n36322# VDD 0.073724f
C219 a_87433_n21335# IN_POS 0.00603f
C220 a_79151_n29181# a_79151_n30339# 0.004047f
C221 a_43817_7563# a_43817_6405# 0.004047f
C222 a_40613_n7136# a_39179_n8033# 5.12e-19
C223 a_108636_n35156# VCM 0.003165f
C224 a_101350_10448# VDD 0.073394f
C225 a_63161_n7138# a_63161_n8932# 0.005987f
C226 a_53497_n16906# a_54019_n16009# 0.005903f
C227 a_83141_n4245# VDD 0.01295f
C228 a_90245_n6960# a_90245_n6055# 0.088786f
C229 a_100235_n15000# VDD 0.016281f
C230 a_102756_n34390# VDD 0.046892f
C231 a_105365_n15000# a_105365_n15905# 0.005903f
C232 a_107339_n15000# a_107339_n18620# 0.011861f
C233 a_45445_n1754# a_45445_n3548# 0.006457f
C234 a_46879_n2651# a_48313_n2651# 0.014106f
C235 a_32353_n12419# a_32913_n12419# 0.0284f
C236 a_72603_n10073# OUT 2.78e-19
C237 a_93969_n1530# a_94537_n1530# 0.027101f
C238 a_86903_n9675# VDD 1.03237f
C239 a_105365_n15905# VDD 0.012916f
C240 a_83141_n15905# a_84547_n18620# 7.35e-19
C241 a_86903_n4245# IN_POS 0.001743f
C242 a_105365_n20430# a_105933_n20430# 0.027101f
C243 a_46879_n7136# a_45445_n8033# 5.12e-19
C244 a_57977_n16906# a_57417_n16906# 0.034628f
C245 a_92601_n9675# a_93131_n7865# 0.012586f
C246 a_95105_n6960# VDD 0.112244f
C247 a_113037_n18620# VDD 1.1868f
C248 a_86903_n16810# a_87433_n13190# 0.032766f
C249 a_64243_n14215# IBNOUT 0.041483f
C250 a_66016_13546# a_66016_12380# 0.004007f
C251 a_53145_n2653# a_54579_n2653# 0.014106f
C252 a_38097_n13316# a_38619_n12419# 0.0284f
C253 a_107198_6405# VDD 0.029136f
C254 a_100235_n2435# a_100803_n2435# 0.027101f
C255 a_98299_n5150# a_98829_n4245# 0.012586f
C256 a_100803_n7865# VDD 0.121044f
C257 a_86903_n21335# a_87433_n18620# 0.012586f
C258 a_90245_n18620# a_89407_n18620# 0.042385f
C259 a_110225_n21335# a_111063_n21335# 0.027101f
C260 a_48349_n35156# a_48349_n36322# 0.004007f
C261 a_54019_n6241# a_54579_n7138# 0.0284f
C262 a_51151_n6241# a_51151_n7138# 0.005987f
C263 a_50629_n7138# a_51711_n8035# 5.37e-19
C264 a_53145_n7138# a_52063_n8035# 0.011365f
C265 a_39179_n16904# a_38097_n17801# 0.001037f
C266 a_40965_n16904# a_41487_n16007# 0.005903f
C267 a_66029_n16906# a_66551_n16906# 0.034714f
C268 a_66551_n16009# a_65677_n17803# 0.034652f
C269 a_100803_n6960# a_100803_n7865# 0.024773f
C270 a_104527_n8770# VDD 0.121415f
C271 a_73302_n34390# I1N 0.003565f
C272 a_92601_n16810# a_92601_n15905# 0.086339f
C273 a_94537_n13190# a_94537_n14095# 0.005903f
C274 a_33787_n1754# a_33787_n2651# 0.005987f
C275 a_31831_n2651# a_31831_n4445# 0.005987f
C276 a_34347_n2651# a_33265_n3548# 5.37e-19
C277 a_32913_n1754# a_34699_n3548# 0.006457f
C278 a_59411_n2653# a_57977_n3550# 1.57e-19
C279 a_30682_13546# VDD 0.073724f
C280 a_103997_n4245# a_104527_n3340# 0.028522f
C281 a_111063_n9675# VDD 0.029377f
C282 a_92601_n21335# a_93969_n20430# 0.002134f
C283 a_94537_n18620# a_94537_n19525# 0.005903f
C284 a_85089_n33224# a_85089_n34390# 0.004007f
C285 a_34347_n7136# a_33265_n8033# 0.00117f
C286 a_31831_n7136# a_32353_n7136# 0.0284f
C287 a_59411_n7138# a_59763_n8035# 0.16936f
C288 a_55635_13546# VDD 0.021314f
C289 a_93969_n21335# IBPOUT 0.003499f
C290 a_45445_n16904# a_46879_n17801# 4.66e-19
C291 a_88271_n13190# VDD 0.02546f
C292 a_105365_n7865# a_105365_n8770# 0.005903f
C293 a_36562_n33224# VDD 0.021515f
C294 a_98299_n15905# a_98829_n15000# 0.028522f
C295 a_114516_12380# a_114516_11614# 0.00778f
C296 a_41487_n1754# a_42047_n2651# 0.0284f
C297 a_65677_n2653# a_65117_n2653# 0.0284f
C298 a_77776_12380# VDD 0.017204f
C299 a_83709_n8770# a_83709_n9675# 0.024773f
C300 a_111631_n3340# a_112199_n3340# 0.027101f
C301 a_93969_n14095# VDD 0.016652f
C302 a_32088_12380# I1U 0.003282f
C303 a_67422_n35156# VDD 0.061113f
C304 a_99667_n19525# a_99667_n20430# 0.005903f
C305 a_63683_n7138# a_64243_n8035# 0.0284f
C306 a_102756_11614# VDD 0.046892f
C307 a_82573_n4245# VDD 0.023101f
C308 a_111063_n8770# a_111063_n9675# 0.005903f
C309 a_99667_n15000# VDD 0.016281f
C310 a_101350_n34390# VDD 0.062166f
C311 a_105933_n15000# a_106501_n15000# 0.027101f
C312 a_46879_n2651# a_47753_n1754# 5.43e-19
C313 a_44363_n2651# a_45797_n3548# 1.57e-19
C314 a_31831_n13316# a_32913_n12419# 5.37e-19
C315 a_90245_n6055# VDD 0.472471f
C316 a_83141_n15905# a_83709_n15905# 0.027101f
C317 a_73268_n27257# I1N -8.11e-35
C318 a_104527_n15905# VDD 0.137705f
C319 a_81735_n15905# a_81735_n17715# 0.006141f
C320 a_47231_n6239# a_47231_n8033# 0.009483f
C321 a_32913_n16904# a_32353_n16904# 0.035468f
C322 a_35221_n15110# a_35221_n16007# 0.005987f
C323 a_59763_n16906# a_59411_n17803# 0.070243f
C324 a_60285_n15112# a_60285_n16009# 0.005987f
C325 a_57977_n16906# a_56895_n17803# 0.002568f
C326 a_94537_n6960# VDD 0.023105f
C327 a_93131_n6960# a_93969_n6960# 0.027101f
C328 a_112199_n15905# VDD 0.112244f
C329 a_63683_n13318# IBNOUT 0.004735f
C330 a_111063_n15905# a_111631_n15905# 0.027101f
C331 a_32088_n35156# a_32088_n36322# 0.004007f
C332 a_53145_n2653# a_54019_n1756# 5.43e-19
C333 a_50629_n2653# a_52063_n3550# 1.57e-19
C334 a_108602_7563# VDD 0.00658f
C335 a_63161_n13318# a_63683_n12421# 0.0284f
C336 a_100235_n7865# VDD 0.016281f
C337 a_90245_n18620# a_88839_n18620# 0.002302f
C338 a_86903_n21335# a_86903_n19525# 0.086469f
C339 a_111631_n20430# a_111631_n21335# 0.005903f
C340 a_77776_13546# a_77776_12380# 0.004007f
C341 a_53145_n7138# a_51711_n8035# 9.78e-20
C342 a_50629_n7138# a_51151_n7138# 0.0284f
C343 a_40965_n16904# a_40613_n17801# 0.534125f
C344 a_40613_n14213# a_42047_n17801# 0.009477f
C345 a_98829_n7865# a_99667_n7865# 0.027101f
C346 a_32353_n16904# I1U 0.002649f
C347 a_66016_n34390# a_66016_n35156# 0.00778f
C348 a_34347_n2651# a_32913_n3548# 1.57e-19
C349 a_60285_n1756# a_60845_n2653# 0.0284f
C350 a_110225_n9675# VDD 0.188021f
C351 a_103997_n5150# a_104527_n6055# 0.03483f
C352 a_105933_n2435# a_105933_n3340# 0.005903f
C353 a_92601_n21335# a_93131_n20430# 0.012586f
C354 a_85129_n30339# IN_POS 6.24e-19
C355 a_101350_12380# a_101350_11614# 0.00778f
C356 a_34347_n7136# a_32913_n8033# 5.12e-19
C357 a_56895_n7138# a_58329_n8035# 1.57e-19
C358 a_59411_n7138# a_58851_n7138# 0.0284f
C359 a_93131_n21335# IBPOUT 0.018739f
C360 a_82573_n3340# a_82573_n4245# 0.005903f
C361 a_84547_n3340# a_84547_n6960# 0.012104f
C362 a_106501_n7865# a_107339_n8770# 0.028522f
C363 a_87433_n13190# VDD 0.150485f
C364 a_100235_n14095# a_100235_n15000# 0.005903f
C365 a_32088_n36322# VDD 0.05845f
C366 a_98299_n16810# a_98829_n17715# 0.03483f
C367 a_39179_n1754# a_39179_n3548# 0.006457f
C368 a_40613_n2651# a_42047_n2651# 0.014106f
C369 a_65117_n1756# a_65117_n2653# 0.005987f
C370 a_65677_n2653# a_64595_n3550# 5.37e-19
C371 a_63161_n2653# a_63161_n4447# 0.005987f
C372 a_81735_n9675# a_82573_n9675# 0.027101f
C373 a_110225_n3340# a_110225_n4245# 0.024773f
C374 a_93131_n14095# VDD 0.121415f
C375 a_109695_n4245# a_111063_n4245# 2.31e-19
C376 a_30682_12380# I1U 0.005416f
C377 a_66016_n35156# VDD 0.076387f
C378 a_100803_n19525# a_101641_n20430# 0.028522f
C379 a_77747_n29181# a_77747_n30339# 0.004047f
C380 a_42413_7563# a_42413_6405# 0.004047f
C381 a_108636_n34390# VCM 0.009172f
C382 a_41487_n5342# a_41487_n6239# 0.005987f
C383 a_38097_n7136# a_38619_n6239# 0.0284f
C384 a_40613_n7136# a_42047_n7136# 0.003256f
C385 a_40965_n6239# a_40965_n8033# 0.009483f
C386 a_65677_n7138# a_66551_n7138# 0.006769f
C387 a_101350_11614# VDD 0.062166f
C388 a_53497_n16906# a_54019_n15112# 0.035574f
C389 a_54579_n15112# a_53145_n17803# 0.009477f
C390 a_51711_n16906# a_51151_n16009# 0.00587f
C391 a_81735_n4245# VDD 0.113729f
C392 a_98829_n15000# VDD 0.121044f
C393 a_111631_n8770# a_112199_n8770# 0.027101f
C394 a_102756_n33224# VDD 0.05812f
C395 a_103997_n15905# a_105365_n15905# 2.31e-19
C396 a_104527_n15000# a_104527_n15905# 0.024773f
C397 a_72603_n9297# OUT 2.78e-19
C398 a_45445_n1754# a_48313_n2651# 5.37e-19
C399 a_44885_n1754# a_44885_n2651# 0.005987f
C400 a_44363_n2651# a_45445_n3548# 5.37e-19
C401 a_31831_n13316# a_32353_n12419# 0.0284f
C402 a_93131_n1530# a_93969_n1530# 0.027101f
C403 a_87433_n6055# VDD 0.41764f
C404 a_106501_n15000# VDD 0.121044f
C405 a_104527_n20430# a_105365_n20430# 0.027101f
C406 a_107339_n20430# a_106501_n20430# 0.028522f
C407 a_73268_6405# a_73268_5639# 0.00778f
C408 VCM IN_POS 0.3453f
C409 a_47753_n5342# a_47753_n6239# 0.005987f
C410 a_46879_n7136# a_48313_n7136# 0.003256f
C411 a_44363_n7136# a_44885_n6239# 0.0284f
C412 a_73268_5639# VDD 0.042519f
C413 a_32913_n16904# a_31831_n17801# 0.001037f
C414 a_34699_n16904# a_35221_n16007# 0.005903f
C415 a_59763_n16906# a_60285_n16009# 0.005903f
C416 a_92601_n7865# a_93969_n6960# 2.31e-19
C417 a_93969_n6960# VDD 0.012916f
C418 a_111631_n15905# VDD 0.023105f
C419 a_112199_n15000# a_112199_n15905# 0.024773f
C420 a_50629_n2653# a_51711_n3550# 5.37e-19
C421 a_51151_n1756# a_51151_n2653# 0.005987f
C422 a_99667_n2435# a_100235_n2435# 0.027101f
C423 a_99667_n7865# VDD 0.016281f
C424 a_37934_n30339# VDD 0.00658f
C425 a_87433_n17715# a_87433_n18620# 0.006141f
C426 a_49755_n34390# a_49755_n35156# 0.00778f
C427 a_53497_n6241# a_53497_n8035# 0.0089f
C428 a_39179_n16904# a_40613_n17801# 4.66e-19
C429 a_64243_n16906# a_63683_n16906# 0.034628f
C430 a_100235_n6960# a_100235_n7865# 0.005903f
C431 a_98299_n9675# a_99667_n8770# 0.002134f
C432 a_107339_n8770# VDD 0.392932f
C433 a_93969_n13190# a_93969_n14095# 0.005903f
C434 a_31831_n17801# I1U -2.34e-34
C435 a_35221_n1754# a_35781_n2651# 0.0284f
C436 a_59411_n2653# a_60845_n2653# 0.014106f
C437 a_112199_n8770# VDD 0.180629f
C438 a_93969_n18620# a_93969_n19525# 0.005903f
C439 a_83683_n33224# a_83683_n34390# 0.004007f
C440 w_27790_n38888# IN_NEG 0.395442f
C441 a_56895_n7138# a_57977_n8035# 5.37e-19
C442 a_60285_n6241# a_60845_n7138# 0.0284f
C443 a_59411_n7138# a_58329_n8035# 0.011365f
C444 a_57417_n6241# a_57417_n7138# 0.005987f
C445 a_45445_n16904# a_44885_n16007# 0.00587f
C446 a_83141_n3340# a_83709_n3340# 0.027101f
C447 a_105933_n7865# a_107339_n8770# 2.31e-19
C448 a_86903_n16810# VDD 1.27745f
C449 a_104527_n7865# a_104527_n8770# 0.024773f
C450 a_30682_n36322# VDD 0.073724f
C451 a_113110_12380# a_113110_11614# 0.00778f
C452 a_38097_n2651# a_39531_n3548# 1.57e-19
C453 a_40613_n2651# a_41487_n1754# 5.43e-19
C454 a_79182_13546# VDD 0.024605f
C455 a_65677_n2653# a_64243_n3550# 1.57e-19
C456 a_83141_n8770# a_83141_n9675# 0.005903f
C457 a_111063_n3340# a_111631_n3340# 0.027101f
C458 a_109695_n4245# a_110225_n4245# 0.028522f
C459 a_100235_n19525# a_101641_n20430# 2.31e-19
C460 a_67422_n34390# VDD 0.046892f
C461 a_98829_n19525# a_98829_n20430# 0.024773f
C462 a_32088_13546# I1U 0.003282f
C463 a_40613_n7136# a_41487_n6239# 4.96e-19
C464 a_65677_n7138# a_66029_n8035# 0.16936f
C465 a_102756_12380# VDD 0.061113f
C466 a_51151_n15112# a_51151_n16009# 0.005987f
C467 a_83709_n3340# VDD 0.121044f
C468 a_89407_n4245# a_90245_n6960# 0.032618f
C469 a_98299_n15905# VDD 0.399575f
C470 a_110225_n8770# a_110225_n9675# 0.024773f
C471 a_105365_n15000# a_105933_n15000# 0.027101f
C472 a_103997_n15905# a_104527_n15905# 0.028522f
C473 a_101350_n33224# VDD 0.073394f
C474 a_44363_n2651# a_44885_n2651# 0.0284f
C475 a_45445_n1754# a_47753_n1754# 0.0284f
C476 a_46319_n1754# a_46879_n2651# 0.0284f
C477 a_90245_n6960# VDD 1.18674f
C478 a_92601_n5150# a_93969_n1530# 7.4e-19
C479 a_82573_n15905# a_83141_n15905# 0.027101f
C480 a_105933_n15000# VDD 0.016281f
C481 a_107339_n20430# a_105933_n20430# 2.31e-19
C482 a_106501_n19525# a_106501_n20430# 0.024773f
C483 a_46879_n7136# a_47753_n6239# 4.96e-19
C484 a_34699_n16904# a_34347_n17801# 0.534125f
C485 a_34347_n14213# a_35781_n17801# 0.009477f
C486 a_71864_5639# VDD 0.042519f
C487 a_93131_n6960# VDD 0.137705f
C488 a_92601_n7865# a_93131_n6960# 0.028522f
C489 a_92601_n9675# a_93969_n6960# 0.002134f
C490 a_111063_n15905# VDD 0.012916f
C491 a_110225_n15905# a_111063_n15905# 0.027101f
C492 a_30682_n35156# a_30682_n36322# 0.004007f
C493 a_50629_n2653# a_51151_n2653# 0.0284f
C494 a_52585_n1756# a_53145_n2653# 0.0284f
C495 a_100803_n1530# a_100803_n2435# 0.024773f
C496 a_98829_n7865# VDD 0.121044f
C497 a_98299_n5150# a_99667_n3340# 0.002134f
C498 a_111063_n20430# a_111063_n21335# 0.005903f
C499 a_53145_n7138# a_54579_n7138# 0.08885f
C500 a_66029_n16906# a_65677_n17803# 0.070243f
C501 a_64243_n16906# a_63161_n17803# 0.002568f
C502 a_66551_n15112# a_66551_n16009# 0.005987f
C503 a_106501_n7865# VDD 0.121044f
C504 a_98299_n9675# a_98829_n8770# 0.012586f
C505 a_73302_n33224# I1N 0.00386f
C506 a_67422_n33224# a_67422_n34390# 0.004007f
C507 a_34347_n2651# a_35781_n2651# 0.014106f
C508 a_32913_n1754# a_32913_n3548# 0.006457f
C509 a_56895_n2653# a_58329_n3550# 1.57e-19
C510 a_59411_n2653# a_60285_n1756# 5.43e-19
C511 a_105365_n2435# a_105365_n3340# 0.005903f
C512 a_111631_n8770# VDD 0.022711f
C513 a_90935_n30339# VDD 0.00658f
C514 a_94537_n18620# a_95105_n18620# 0.027101f
C515 a_85129_n29181# IN_POS 6.24e-19
C516 a_102756_13546# a_102756_12380# 0.004007f
C517 a_34347_n7136# a_35781_n7136# 0.003256f
C518 a_31831_n7136# a_32353_n6239# 0.0284f
C519 a_34699_n6239# a_34699_n8033# 0.009483f
C520 a_35221_n5342# a_35221_n6239# 0.005987f
C521 a_59411_n7138# a_57977_n8035# 9.78e-20
C522 a_54229_13546# VDD 0.021314f
C523 a_56895_n7138# a_57417_n7138# 0.0284f
C524 a_47231_n16904# a_47753_n15110# 0.034714f
C525 a_46879_n14213# a_47753_n16007# 0.034652f
C526 a_44885_n15110# a_44885_n16007# 0.005987f
C527 a_94537_n20430# IBPOUT 0.00243f
C528 a_81735_n3340# a_81735_n4245# 0.024773f
C529 a_81205_n4245# a_82573_n4245# 2.31e-19
C530 a_83709_n21335# VDD 0.177586f
C531 a_105933_n7865# a_106501_n7865# 0.027101f
C532 a_32088_n35156# VDD 0.061113f
C533 a_99667_n14095# a_99667_n15000# 0.005903f
C534 a_32353_n7136# I1U 0.002649f
C535 a_66058_n27257# a_66058_n28415# 0.004047f
C536 a_38097_n2651# a_39179_n3548# 5.37e-19
C537 a_38619_n1754# a_38619_n2651# 0.005987f
C538 a_39179_n1754# a_42047_n2651# 5.37e-19
C539 a_66551_n1756# a_67111_n2653# 0.0284f
C540 a_48313_n19595# a_47753_n19595# 0.0284f
C541 a_30682_13546# I1U 0.005416f
C542 a_95105_n13190# VDD 0.209912f
C543 a_100235_n19525# a_100803_n19525# 0.027101f
C544 a_66016_n34390# VDD 0.062166f
C545 a_87433_n20430# IN_POS 0.00603f
C546 a_41100_19698# a_41100_19075# 0.007809f
C547 a_79151_n28415# a_79151_n29181# 0.00778f
C548 a_108636_n33224# VCM 0.02829f
C549 a_65677_n7138# a_65117_n7138# 0.0284f
C550 a_101350_12380# VDD 0.076387f
C551 a_63161_n7138# a_64595_n8035# 1.57e-19
C552 a_53145_n14215# a_53145_n17803# 0.00969f
C553 a_51711_n16906# a_53497_n16906# 0.012473f
C554 a_83141_n3340# VDD 0.016281f
C555 a_88839_n4245# a_90245_n6960# 7.35e-19
C556 a_111063_n8770# a_111631_n8770# 0.027101f
C557 a_101641_n15000# VDD 0.399226f
C558 a_96849_n36322# VDD 0.024605f
C559 a_45445_n1754# a_46879_n2651# 0.054819f
C560 a_51711_n19597# a_54019_n19597# 0.0284f
C561 a_89407_n4245# VDD 0.138244f
C562 a_92601_n5150# a_93131_n1530# 0.032766f
C563 a_105365_n15000# VDD 0.016281f
C564 a_83709_n15000# a_83709_n15905# 0.024773f
C565 a_71864_6405# a_71864_5639# 0.00778f
C566 a_32913_n16904# a_34347_n17801# 4.66e-19
C567 a_73268_6405# VDD 0.034176f
C568 a_59763_n16906# a_60285_n15112# 0.035574f
C569 a_60845_n15112# a_59411_n17803# 0.009477f
C570 a_57977_n16906# a_57417_n16009# 0.00587f
C571 a_92601_n7865# VDD 0.399575f
C572 a_95943_n6960# a_95105_n6960# 0.042385f
C573 a_92601_n9675# a_93131_n6960# 0.012586f
C574 a_110225_n15905# VDD 0.137705f
C575 a_65677_n13318# IBNOUT 0.006509f
C576 a_83141_n21335# a_83709_n21335# 0.027101f
C577 a_111631_n15000# a_111631_n15905# 0.005903f
C578 a_100803_n6960# VDD 0.138244f
C579 a_98299_n5150# a_98829_n3340# 0.012586f
C580 a_98829_n2435# a_99667_n2435# 0.027101f
C581 a_87433_n17715# a_86903_n21335# 0.03483f
C582 a_37934_n29181# VDD 0.034176f
C583 a_111631_n20430# a_112199_n20430# 0.027101f
C584 a_48349_n34390# a_48349_n35156# 0.00778f
C585 a_53145_n7138# a_54019_n6241# 0.005903f
C586 a_50629_n7138# a_51151_n6241# 0.0284f
C587 a_39179_n16904# a_38619_n16007# 0.00587f
C588 a_66029_n16906# a_66551_n16009# 0.005903f
C589 a_105933_n7865# VDD 0.016281f
C590 a_99667_n6960# a_99667_n7865# 0.005903f
C591 a_94537_n13190# a_95105_n13190# 0.027101f
C592 a_92601_n16810# a_93969_n14095# 0.002134f
C593 a_93131_n13190# a_93131_n14095# 0.024773f
C594 a_31831_n2651# a_33265_n3548# 1.57e-19
C595 a_34347_n2651# a_35221_n1754# 5.43e-19
C596 a_57417_n1756# a_57417_n2653# 0.005987f
C597 a_56895_n2653# a_57977_n3550# 5.37e-19
C598 a_106501_n2435# a_107339_n3340# 0.028522f
C599 a_111063_n8770# VDD 0.016883f
C600 a_93131_n18620# a_93131_n19525# 0.024773f
C601 a_92601_n19525# a_93969_n19525# 2.31e-19
C602 a_34347_n7136# a_35221_n6239# 4.96e-19
C603 a_59763_n6241# a_59763_n8035# 0.0089f
C604 a_93969_n20430# IBPOUT 0.003499f
C605 a_46879_n14213# a_46879_n17801# 0.00969f
C606 a_82573_n3340# a_83141_n3340# 0.027101f
C607 a_81205_n4245# a_81735_n4245# 0.028522f
C608 a_83141_n21335# VDD 0.02546f
C609 a_103997_n9675# a_105365_n9675# 7.4e-19
C610 a_30682_n35156# VDD 0.076387f
C611 a_100803_n14095# a_101641_n15000# 0.028522f
C612 a_38097_n2651# a_38619_n2651# 0.0284f
C613 a_39179_n1754# a_41487_n1754# 0.0284f
C614 a_40053_n1754# a_40613_n2651# 0.0284f
C615 a_77776_13546# VDD 0.029536f
C616 a_65677_n2653# a_67111_n2653# 0.014106f
C617 a_47753_n18698# a_47753_n19595# 0.005987f
C618 a_82573_n8770# a_82573_n9675# 0.005903f
C619 a_113037_n3340# a_112199_n3340# 0.028522f
C620 a_94537_n13190# VDD 0.031519f
C621 a_110225_n3340# a_111063_n3340# 0.027101f
C622 a_98299_n21335# a_99667_n21335# 7.4e-19
C623 a_67422_n33224# VDD 0.05812f
C624 a_40578_19075# a_41100_19075# 0.017917f
C625 a_102756_13546# VDD 0.05845f
C626 a_63683_n6241# a_63683_n7138# 0.005987f
C627 a_65677_n7138# a_64595_n8035# 0.011365f
C628 a_63161_n7138# a_64243_n8035# 5.37e-19
C629 a_66551_n6241# a_67111_n7138# 0.0284f
C630 a_54579_n15112# a_54019_n15112# 0.0284f
C631 a_53145_n14215# a_54019_n16009# 0.030444f
C632 a_82573_n3340# VDD 0.016281f
C633 a_87433_n4245# a_87433_n6055# 0.006141f
C634 a_88839_n4245# a_89407_n4245# 0.027101f
C635 a_100803_n14095# VDD 0.121415f
C636 a_113037_n8770# a_112199_n8770# 0.028522f
C637 a_104527_n15000# a_105365_n15000# 0.027101f
C638 a_95443_n36322# VDD 0.029536f
C639 a_103997_n16810# a_103997_n21335# 0.032645f
C640 a_107339_n15000# a_106501_n15000# 0.028522f
C641 a_45445_n1754# a_46319_n1754# 0.001405f
C642 a_32088_n36322# I1U 0.003282f
C643 a_72603_n8397# OUT 2.78e-19
C644 a_51711_n19597# a_52585_n19597# 0.001405f
C645 a_88839_n4245# VDD 0.01295f
C646 a_87433_n2435# IN_POS 0.00603f
C647 a_81735_n15905# a_82573_n15905# 0.027101f
C648 a_104527_n15000# VDD 0.121044f
C649 a_105933_n19525# a_105933_n20430# 0.005903f
C650 a_45445_n6239# a_45445_n8033# 0.009307f
C651 a_71864_6405# VDD 0.029136f
C652 a_57417_n15112# a_57417_n16009# 0.005987f
C653 a_92601_n9675# VDD 1.40063f
C654 a_92601_n9675# a_92601_n7865# 0.086469f
C655 a_95943_n6960# a_94537_n6960# 0.002302f
C656 a_65117_n12421# IBNOUT -2.71e-34
C657 a_112199_n15000# VDD 0.121044f
C658 a_32088_n34390# a_32088_n35156# 0.00778f
C659 a_100235_n6960# VDD 0.01295f
C660 a_100235_n1530# a_100235_n2435# 0.005903f
C661 a_98299_n5150# a_98299_n4245# 0.086469f
C662 a_36530_n29181# VDD 0.029136f
C663 a_110225_n20430# a_110225_n21335# 0.024773f
C664 a_54019_n5344# a_54019_n6241# 0.005987f
C665 a_40965_n16904# a_41487_n15110# 0.034714f
C666 a_38619_n15110# a_38619_n16007# 0.005987f
C667 a_40613_n14213# a_41487_n16007# 0.034652f
C668 a_105365_n7865# VDD 0.016281f
C669 IN_POS IN_NEG 3.17862f
C670 a_100235_n6960# a_100803_n6960# 0.027101f
C671 a_92601_n16810# a_93131_n14095# 0.012586f
C672 a_66016_n33224# a_66016_n34390# 0.004007f
C673 a_31831_n2651# a_32913_n3548# 5.37e-19
C674 a_32913_n1754# a_35781_n2651# 5.37e-19
C675 a_32353_n1754# a_32353_n2651# 0.005987f
C676 a_56895_n2653# a_57417_n2653# 0.0284f
C677 a_58851_n1756# a_59411_n2653# 0.0284f
C678 a_42047_n19595# a_41487_n19595# 0.0284f
C679 a_110225_n8770# VDD 0.152953f
C680 a_103997_n5150# a_105365_n4245# 0.002134f
C681 a_105933_n2435# a_107339_n3340# 2.31e-19
C682 a_104527_n2435# a_104527_n3340# 0.024773f
C683 a_95943_n18620# a_95943_n20430# 0.011861f
C684 a_92601_n19525# a_93131_n19525# 0.028522f
C685 a_93969_n18620# a_94537_n18620# 0.027101f
C686 a_92601_n21335# a_93969_n19525# 0.002134f
C687 a_90935_n29181# VDD 0.034176f
C688 a_85129_n28415# IN_POS 6.24e-19
C689 a_101350_13546# a_101350_12380# 0.004007f
C690 a_59411_n7138# a_60845_n7138# 0.08885f
C691 a_93131_n20430# IBPOUT 0.01873f
C692 a_45445_n16904# a_47231_n16904# 0.012473f
C693 a_82573_n21335# VDD 0.02546f
C694 a_105365_n7865# a_105933_n7865# 0.027101f
C695 a_103997_n9675# a_104527_n9675# 0.032766f
C696 a_98829_n14095# a_98829_n15000# 0.024773f
C697 a_98299_n16810# a_99667_n15905# 0.002134f
C698 a_100235_n14095# a_101641_n15000# 2.31e-19
C699 a_32088_n34390# VDD 0.046892f
C700 a_39179_n1754# a_40613_n2651# 0.054819f
C701 a_65677_n2653# a_66551_n1756# 5.43e-19
C702 a_63161_n2653# a_64595_n3550# 1.57e-19
C703 a_46879_n19595# a_47753_n19595# 5.43e-19
C704 a_83141_n8770# a_83709_n8770# 0.027101f
C705 a_109695_n4245# a_111063_n3340# 2.31e-19
C706 a_113037_n3340# a_111631_n3340# 2.31e-19
C707 a_109695_n5150# a_109695_n9675# 0.032645f
C708 a_112199_n2435# a_112199_n3340# 0.024773f
C709 a_93969_n13190# VDD 0.02546f
C710 a_98299_n21335# a_98829_n21335# 0.032766f
C711 a_66016_n33224# VDD 0.073394f
C712 a_99667_n19525# a_100235_n19525# 0.027101f
C713 a_40578_19075# a_41100_19698# 0.017917f
C714 a_77747_n28415# a_77747_n29181# 0.00778f
C715 a_39179_n6239# a_39179_n8033# 0.009307f
C716 a_38619_n5342# a_38619_n6239# 0.005987f
C717 a_40613_n7136# a_41487_n5342# 0.030444f
C718 a_101350_13546# VDD 0.073724f
C719 a_102756_n36322# VCM 0.002253f
C720 a_65677_n7138# a_64243_n8035# 9.78e-20
C721 a_63161_n7138# a_63683_n7138# 0.0284f
C722 a_54019_n14215# a_54019_n15112# 0.005987f
C723 a_54579_n15112# a_53497_n16906# 0.002917f
C724 a_51151_n15112# a_51711_n16906# 0.035468f
C725 a_81735_n3340# VDD 0.121044f
C726 a_113037_n8770# a_111631_n8770# 2.31e-19
C727 a_112199_n7865# a_112199_n8770# 0.024773f
C728 a_110225_n8770# a_111063_n8770# 0.027101f
C729 a_100235_n14095# VDD 0.016652f
C730 a_96849_n35156# VDD 0.009062f
C731 a_106501_n14095# a_106501_n15000# 0.024773f
C732 a_107339_n15000# a_105933_n15000# 2.31e-19
C733 a_103997_n15905# a_105365_n15000# 2.31e-19
C734 a_30682_n36322# I1U 0.005416f
C735 a_54579_n19597# a_54019_n19597# 0.0284f
C736 a_88271_n4245# VDD 0.023101f
C737 a_83141_n15000# a_83141_n15905# 0.005903f
C738 a_103997_n15905# VDD 0.399575f
C739 a_46879_n7136# a_47753_n5342# 0.030444f
C740 a_44885_n5342# a_44885_n6239# 0.005987f
C741 a_47231_n6239# a_48313_n7136# 0.002917f
C742 a_73268_7563# VDD 0.00658f
C743 a_32913_n16904# a_32353_n16007# 0.00587f
C744 a_57977_n16906# a_59763_n16906# 0.012473f
C745 a_59411_n14215# a_59411_n17803# 0.00969f
C746 a_95943_n6055# VDD 0.472471f
C747 a_93131_n6055# a_93131_n6960# 0.006141f
C748 a_82573_n21335# a_83141_n21335# 0.027101f
C749 a_111631_n15000# VDD 0.016281f
C750 a_111063_n15000# a_111063_n15905# 0.005903f
C751 a_113037_n15000# a_113037_n18620# 0.011861f
C752 a_57977_n19597# a_60285_n19597# 0.0284f
C753 a_99667_n6960# VDD 0.023101f
C754 a_90245_n18620# a_90245_n17715# 0.088786f
C755 a_37934_n28415# VDD 0.042519f
C756 a_111063_n20430# a_111631_n20430# 0.027101f
C757 a_49755_n33224# a_49755_n34390# 0.004007f
C758 a_101392_5639# a_101392_4481# 0.004047f
C759 a_51711_n6241# a_51711_n8035# 0.008933f
C760 a_40613_n14213# a_40613_n17801# 0.00969f
C761 a_66029_n16906# a_66551_n15112# 0.035574f
C762 a_64243_n16906# a_63683_n16009# 0.00587f
C763 a_67111_n15112# a_65677_n17803# 0.009477f
C764 a_104527_n7865# VDD 0.121044f
C765 a_98829_n6960# a_98829_n7865# 0.024773f
C766 a_98299_n7865# a_99667_n7865# 2.31e-19
C767 a_93969_n13190# a_94537_n13190# 0.027101f
C768 a_37934_n28415# a_37934_n29181# 0.00778f
C769 a_32353_n16007# I1U 0.002649f
C770 a_33787_n1754# a_34347_n2651# 0.0284f
C771 a_32913_n1754# a_35221_n1754# 0.0284f
C772 a_31831_n2651# a_32353_n2651# 0.0284f
C773 a_41487_n18698# a_41487_n19595# 0.005987f
C774 a_113037_n8770# VDD 0.39614f
C775 a_103997_n5150# a_104527_n4245# 0.012586f
C776 a_105933_n2435# a_106501_n2435# 0.027101f
C777 a_92601_n21335# a_93131_n19525# 0.012586f
C778 a_89531_n29181# VDD 0.029136f
C779 a_49755_10448# VDD 0.05812f
C780 a_59411_n7138# a_60285_n6241# 0.005903f
C781 a_56895_n7138# a_57417_n6241# 0.0284f
C782 a_48313_n15110# a_47753_n15110# 0.0284f
C783 a_84547_n3340# a_83709_n3340# 0.028522f
C784 a_81735_n3340# a_82573_n3340# 0.027101f
C785 a_81735_n21335# VDD 0.150485f
C786 a_106501_n6960# a_106501_n7865# 0.024773f
C787 a_98299_n16810# a_98829_n15905# 0.012586f
C788 a_30682_n34390# VDD 0.062166f
C789 a_100235_n14095# a_100803_n14095# 0.027101f
C790 a_32353_n6239# I1U 0.002649f
C791 a_39179_n1754# a_40053_n1754# 0.001405f
C792 a_73302_10448# VDD 0.021515f
C793 a_63683_n1756# a_63683_n2653# 0.005987f
C794 a_63161_n2653# a_64243_n3550# 5.37e-19
C795 a_46879_n19595# a_46319_n19595# 0.0284f
C796 a_81735_n8770# a_81735_n9675# 0.024773f
C797 a_93131_n13190# VDD 0.150485f
C798 a_109695_n4245# a_110225_n3340# 0.028522f
C799 a_61515_n36322# VDD 0.024605f
C800 a_100803_n18620# a_100803_n19525# 0.024773f
C801 a_41660_19698# a_41100_19698# 0.017917f
C802 a_113110_n35156# a_113110_n36322# 0.004007f
C803 a_40965_n6239# a_42047_n7136# 0.002917f
C804 a_101350_n36322# VCM 0.002253f
C805 a_66029_n6241# a_66029_n8035# 0.0089f
C806 a_53145_n14215# a_54019_n15112# 4.96e-19
C807 a_88271_n4245# a_88839_n4245# 0.027101f
C808 a_81205_n4245# VDD 0.393432f
C809 a_99667_n14095# VDD 0.016652f
C810 a_103997_n15905# a_104527_n15000# 0.028522f
C811 a_95443_n35156# VDD 0.017204f
C812 a_55601_6405# a_55601_5639# 0.00778f
C813 a_44885_n1754# a_45445_n1754# 0.0284f
C814 a_37934_5639# VDD 0.042519f
C815 a_32088_n35156# I1U 0.003282f
C816 a_75602_n4019# a_75602_n4978# 0.005385f
C817 a_51151_n19597# a_51711_n19597# 0.0284f
C818 a_54019_n18700# a_54019_n19597# 0.005987f
C819 a_87433_n4245# VDD 0.113729f
C820 a_107339_n15000# VDD 0.399226f
C821 a_105365_n19525# a_105365_n20430# 0.005903f
C822 a_47231_n6239# a_47753_n6239# 0.035574f
C823 a_34699_n16904# a_35221_n15110# 0.034714f
C824 a_34347_n14213# a_35221_n16007# 0.034652f
C825 a_32353_n15110# a_32353_n16007# 0.005987f
C826 a_60845_n15112# a_60285_n15112# 0.0284f
C827 a_59411_n14215# a_60285_n16009# 0.030444f
C828 a_93131_n6055# VDD 0.41764f
C829 a_83709_n20430# a_83709_n21335# 0.024773f
C830 a_63683_n12421# IBNOUT 0.041834f
C831 a_111063_n15000# VDD 0.016281f
C832 a_111631_n15000# a_112199_n15000# 0.027101f
C833 a_30682_n34390# a_30682_n35156# 0.00778f
C834 a_72596_n4978# OUT 3.16e-19
C835 a_35781_n19595# a_35221_n19595# 0.0284f
C836 a_57977_n19597# a_58851_n19597# 0.001405f
C837 a_98829_n6960# VDD 0.113729f
C838 a_99667_n1530# a_99667_n2435# 0.005903f
C839 a_36530_n28415# VDD 0.042519f
C840 a_53497_n6241# a_54579_n7138# 0.001641f
C841 a_51151_n5344# a_51151_n6241# 0.005987f
C842 a_39179_n16904# a_40965_n16904# 0.012473f
C843 a_63683_n15112# a_63683_n16009# 0.005987f
C844 a_106501_n6960# VDD 0.138244f
C845 a_98299_n7865# a_98829_n7865# 0.028522f
C846 a_99667_n6960# a_100235_n6960# 0.027101f
C847 VDD I1U 1.71173f
C848 a_32913_n1754# a_34347_n2651# 0.054819f
C849 a_40613_n19595# a_41487_n19595# 5.43e-19
C850 a_112199_n7865# VDD 0.180258f
C851 a_93131_n18620# a_93969_n18620# 0.027101f
C852 a_90935_n28415# VDD 0.042519f
C853 a_34347_n7136# a_35221_n5342# 0.030444f
C854 a_32353_n5342# a_32353_n6239# 0.005987f
C855 a_32913_n6239# a_32913_n8033# 0.009307f
C856 a_60285_n5344# a_60285_n6241# 0.005987f
C857 a_48349_10448# VDD 0.073394f
C858 a_47753_n14213# a_47753_n15110# 0.005987f
C859 a_48313_n15110# a_47231_n16904# 0.001641f
C860 a_44885_n15110# a_45445_n16904# 0.034628f
C861 a_81205_n4245# a_82573_n3340# 2.31e-19
C862 a_84547_n3340# a_83141_n3340# 2.31e-19
C863 a_83709_n2435# a_83709_n3340# 0.024773f
C864 a_83709_n20430# VDD 0.121415f
C865 a_104527_n7865# a_105365_n7865# 0.027101f
C866 a_32088_n33224# VDD 0.05812f
C867 a_31831_n7136# I1U -9.82e-34
C868 a_95443_n35156# a_95443_n36322# 0.004007f
C869 a_71896_10448# VDD 0.021515f
C870 a_65117_n1756# a_65677_n2653# 0.0284f
C871 a_63161_n2653# a_63683_n2653# 0.0284f
C872 a_46319_n18698# a_46319_n19595# 0.005987f
C873 a_82573_n8770# a_83141_n8770# 0.027101f
C874 a_92601_n16810# VDD 1.28143f
C875 a_109695_n5150# a_110225_n6055# 0.03483f
C876 a_111631_n2435# a_111631_n3340# 0.005903f
C877 a_98829_n19525# a_99667_n19525# 0.027101f
C878 a_60109_n36322# VDD 0.029536f
C879 a_41660_19698# a_40578_19075# 2.78e-19
C880 a_41100_20251# a_41100_19698# 0.009337f
C881 a_40965_n6239# a_41487_n6239# 0.035574f
C882 a_65677_n7138# a_67111_n7138# 0.08885f
C883 a_53145_n14215# a_53497_n16906# 0.534125f
C884 a_84547_n3340# VDD 0.392932f
C885 a_89407_n3340# a_89407_n4245# 0.024773f
C886 a_98829_n14095# VDD 0.149203f
C887 a_111631_n7865# a_111631_n8770# 0.005903f
C888 a_96849_n34390# VDD 0.011958f
C889 a_103997_n16810# a_104527_n17715# 0.03483f
C890 a_105933_n14095# a_105933_n15000# 0.005903f
C891 a_44363_n2651# a_45445_n1754# 5.37e-19
C892 a_36530_5639# VDD 0.042519f
C893 a_30682_n35156# I1U 0.005416f
C894 a_54579_n19597# a_51711_n19597# 5.37e-19
C895 a_53145_n19597# a_54019_n19597# 5.43e-19
C896 a_89407_n3340# VDD 0.121044f
C897 a_88839_n9675# a_89407_n9675# 0.027101f
C898 a_106501_n14095# VDD 0.121415f
C899 a_84547_n15000# a_84547_n18620# 0.012104f
C900 a_82573_n15000# a_82573_n15905# 0.005903f
C901 a_106501_n19525# a_107339_n20430# 0.028522f
C902 a_34347_n14213# a_34347_n17801# 0.00969f
C903 a_60285_n14215# a_60285_n15112# 0.005987f
C904 a_57417_n15112# a_57977_n16906# 0.035468f
C905 a_60845_n15112# a_59763_n16906# 0.002917f
C906 a_93131_n6055# a_92601_n9675# 0.03483f
C907 a_95943_n6960# VDD 1.18674f
C908 a_110225_n15000# VDD 0.121044f
C909 a_81735_n21335# a_82573_n21335# 0.027101f
C910 a_63161_n13318# IBNOUT 0.002932f
C911 a_110225_n15000# a_110225_n15905# 0.024773f
C912 a_109695_n15905# a_111063_n15905# 2.31e-19
C913 a_35221_n18698# a_35221_n19595# 0.005987f
C914 a_60845_n19597# a_60285_n19597# 0.0284f
C915 a_100235_n1530# a_100803_n1530# 0.027101f
C916 a_98299_n7865# VDD 0.393432f
C917 a_110225_n20430# a_111063_n20430# 0.027101f
C918 a_113037_n20430# a_112199_n20430# 0.028522f
C919 a_48349_n33224# a_48349_n34390# 0.004007f
C920 a_102796_6405# a_102796_5639# 0.00778f
C921 a_53497_n6241# a_54019_n6241# 0.034714f
C922 a_54019_n5344# a_53145_n7138# 0.034652f
C923 a_42047_n15110# a_41487_n15110# 0.0284f
C924 a_65677_n14215# a_65677_n17803# 0.00969f
C925 a_64243_n16906# a_66029_n16906# 0.012473f
C926 a_98299_n9675# a_99667_n7865# 0.002134f
C927 a_105933_n6960# VDD 0.01295f
C928 a_93131_n13190# a_93969_n13190# 0.027101f
C929 a_36530_n28415# a_36530_n29181# 0.00778f
C930 a_32913_n1754# a_33787_n1754# 0.001405f
C931 a_45706_22884# VDD 0.04859f
C932 a_40613_n19595# a_40053_n19595# 0.0284f
C933 a_64243_n19597# a_66551_n19597# 0.0284f
C934 a_105365_n2435# a_105933_n2435# 0.027101f
C935 a_111631_n7865# VDD 0.02234f
C936 a_89531_n28415# VDD 0.042519f
C937 a_92601_n19525# a_93969_n18620# 2.31e-19
C938 a_85129_n27257# IN_POS 6.24e-19
C939 a_34699_n6239# a_35781_n7136# 0.002917f
C940 a_49755_11614# VDD 0.046892f
C941 a_57977_n6241# a_57977_n8035# 0.008933f
C942 a_94537_n19525# IBPOUT 0.00243f
C943 a_46879_n14213# a_47753_n15110# 0.005903f
C944 a_81205_n5150# a_81205_n9675# 0.032645f
C945 a_81205_n4245# a_81735_n3340# 0.028522f
C946 a_83141_n20430# VDD 0.016652f
C947 a_105933_n6960# a_105933_n7865# 0.005903f
C948 a_103997_n9675# a_105365_n8770# 0.002134f
C949 a_99667_n14095# a_100235_n14095# 0.027101f
C950 a_30682_n33224# VDD 0.073394f
C951 a_113110_13546# a_113110_12380# 0.004007f
C952 a_38619_n1754# a_39179_n1754# 0.0284f
C953 a_73302_11614# VDD 0.009062f
C954 a_47753_n18698# a_48313_n19595# 0.0284f
C955 a_84547_n8770# a_83709_n8770# 0.028522f
C956 a_89407_n21335# VDD 0.177586f
C957 a_98299_n21335# a_99667_n20430# 0.002134f
C958 a_87433_n19525# IN_POS 0.00603f
C959 a_100235_n18620# a_100235_n19525# 0.005903f
C960 a_61515_n35156# VDD 0.009062f
C961 a_79151_n27257# a_79151_n28415# 0.004047f
C962 a_114516_n34390# a_114516_n35156# 0.00778f
C963 a_65677_n7138# a_66551_n6241# 0.005903f
C964 a_96849_10448# VDD 0.021515f
C965 a_63161_n7138# a_63683_n6241# 0.0284f
C966 a_53145_n14215# a_51711_n16906# 4.66e-19
C967 a_87433_n4245# a_88271_n4245# 0.027101f
C968 a_83709_n2435# VDD 0.121415f
C969 a_100803_n13190# VDD 0.177586f
C970 a_95443_n34390# VDD 0.017204f
C971 a_90935_n28415# a_90935_n29181# 0.00778f
C972 a_85089_n36322# IN_POS 0.003316f
C973 a_54197_6405# a_54197_5639# 0.00778f
C974 a_44363_n2651# a_44885_n1754# 0.0284f
C975 a_32088_n34390# I1U 0.003282f
C976 a_37934_6405# VDD 0.034176f
C977 a_72596_n4019# a_72596_n4978# 0.005385f
C978 a_53145_n19597# a_52585_n19597# 0.0284f
C979 a_88839_n3340# VDD 0.016281f
C980 a_105933_n14095# VDD 0.016652f
C981 a_83141_n15000# a_83709_n15000# 0.027101f
C982 a_104527_n19525# a_104527_n20430# 0.024773f
C983 a_105933_n19525# a_107339_n20430# 2.31e-19
C984 a_45445_n6239# a_44885_n6239# 0.035468f
C985 a_47753_n4445# a_47753_n5342# 0.005987f
C986 a_32913_n16904# a_34699_n16904# 0.012473f
C987 a_59411_n14215# a_60285_n15112# 4.96e-19
C988 a_95105_n4245# VDD 0.138244f
C989 a_109695_n15905# VDD 0.399575f
C990 a_83141_n20430# a_83141_n21335# 0.005903f
C991 a_111063_n15000# a_111631_n15000# 0.027101f
C992 a_109695_n15905# a_110225_n15905# 0.028522f
C993 a_32088_n33224# a_32088_n34390# 0.004007f
C994 a_72596_n4019# OUT 3.16e-19
C995 a_50629_n2653# a_51151_n1756# 0.0284f
C996 a_34347_n19595# a_35221_n19595# 5.43e-19
C997 a_57417_n19597# a_57977_n19597# 0.0284f
C998 a_60285_n18700# a_60285_n19597# 0.005987f
C999 a_98829_n1530# a_98829_n2435# 0.024773f
C1000 a_98299_n5150# a_99667_n2435# 0.002134f
C1001 a_89407_n15905# a_90245_n18620# 0.032618f
C1002 a_113037_n20430# a_111631_n20430# 2.31e-19
C1003 a_112199_n19525# a_112199_n20430# 0.024773f
C1004 a_41487_n14213# a_41487_n15110# 0.005987f
C1005 a_42047_n15110# a_40965_n16904# 0.001641f
C1006 a_38619_n15110# a_39179_n16904# 0.034628f
C1007 a_65677_n14215# a_66551_n16009# 0.030444f
C1008 a_67111_n15112# a_66551_n15112# 0.0284f
C1009 a_98299_n9675# a_98829_n7865# 0.012586f
C1010 a_101641_n6960# a_101641_n8770# 0.012104f
C1011 a_98829_n6960# a_99667_n6960# 0.027101f
C1012 a_105365_n6960# VDD 0.023101f
C1013 a_92601_n16810# a_93969_n13190# 7.4e-19
C1014 a_45138_22884# VDD 0.040003f
C1015 a_40053_n18698# a_40053_n19595# 0.005987f
C1016 a_64243_n19597# a_65117_n19597# 0.001405f
C1017 a_111063_n7865# VDD 0.016281f
C1018 a_106501_n1530# a_106501_n2435# 0.024773f
C1019 a_103997_n5150# a_105365_n3340# 0.002134f
C1020 a_92601_n21335# a_93969_n18620# 0.002134f
C1021 a_92601_n19525# a_93131_n18620# 0.028522f
C1022 a_48391_n29181# a_48391_n30339# 0.004047f
C1023 a_34699_n6239# a_35221_n6239# 0.035574f
C1024 a_48349_11614# VDD 0.062166f
C1025 a_57417_n5344# a_57417_n6241# 0.005987f
C1026 a_59763_n6241# a_60845_n7138# 0.001641f
C1027 a_93969_n19525# IBPOUT 0.003499f
C1028 a_46879_n14213# a_47231_n16904# 0.070243f
C1029 a_83141_n2435# a_83141_n3340# 0.005903f
C1030 a_103997_n9675# a_104527_n8770# 0.012586f
C1031 a_82573_n20430# VDD 0.016652f
C1032 a_114485_n30339# VDD 0.002225f
C1033 a_98299_n16810# a_99667_n15000# 0.002134f
C1034 a_100803_n13190# a_100803_n14095# 0.024773f
C1035 a_96849_n34390# a_96849_n35156# 0.00778f
C1036 a_38097_n2651# a_39179_n1754# 5.37e-19
C1037 a_71896_11614# VDD 0.009062f
C1038 a_46879_n19595# a_48313_n19595# 0.014106f
C1039 a_81735_n8770# a_82573_n8770# 0.027101f
C1040 a_83709_n7865# a_83709_n8770# 0.024773f
C1041 a_84547_n8770# a_83141_n8770# 2.31e-19
C1042 a_111063_n2435# a_111063_n3340# 0.005903f
C1043 a_88839_n21335# VDD 0.02546f
C1044 a_60109_n35156# VDD 0.017204f
C1045 a_98299_n21335# a_98829_n20430# 0.012586f
C1046 a_41100_20251# a_41660_19698# 0.017917f
C1047 a_41487_n4445# a_41487_n5342# 0.005987f
C1048 a_39179_n6239# a_38619_n6239# 0.035468f
C1049 a_66551_n5344# a_66551_n6241# 0.005987f
C1050 a_95443_10448# VDD 0.029536f
C1051 a_54019_n14215# a_54579_n15112# 0.0284f
C1052 a_88839_n3340# a_88839_n4245# 0.005903f
C1053 a_83141_n2435# VDD 0.016652f
C1054 a_100235_n13190# VDD 0.02546f
C1055 a_112199_n7865# a_113037_n8770# 0.028522f
C1056 a_111063_n7865# a_111063_n8770# 0.005903f
C1057 a_96849_n33224# VDD 0.021515f
C1058 a_105365_n14095# a_105365_n15000# 0.005903f
C1059 a_37968_12380# a_37968_11614# 0.00778f
C1060 a_30682_n34390# I1U 0.005416f
C1061 a_36530_6405# VDD 0.029136f
C1062 a_52585_n18700# a_52585_n19597# 0.005987f
C1063 a_53145_n19597# a_51711_n19597# 0.054819f
C1064 a_88271_n3340# VDD 0.016281f
C1065 a_88271_n9675# a_88839_n9675# 0.027101f
C1066 a_105365_n14095# VDD 0.016652f
C1067 a_81735_n15000# a_81735_n15905# 0.024773f
C1068 a_87433_n1530# IN_POS 0.004984f
C1069 a_81205_n15905# a_82573_n15905# 2.31e-19
C1070 a_105933_n19525# a_106501_n19525# 0.027101f
C1071 a_47231_n6239# a_47753_n5342# 0.005903f
C1072 a_45445_n6239# a_44363_n7136# 0.001037f
C1073 a_35781_n15110# a_35221_n15110# 0.0284f
C1074 a_59411_n14215# a_59763_n16906# 0.534125f
C1075 a_94537_n4245# VDD 0.01295f
C1076 a_95943_n6960# a_95943_n6055# 0.088786f
C1077 a_113037_n15000# VDD 0.399226f
C1078 a_34347_n19595# a_33787_n19595# 0.0284f
C1079 a_60845_n19597# a_57977_n19597# 5.37e-19
C1080 a_59411_n19597# a_60285_n19597# 5.43e-19
C1081 a_98299_n5150# a_98829_n2435# 0.012586f
C1082 a_98299_n9675# VDD 1.27279f
C1083 a_99667_n1530# a_100235_n1530# 0.027101f
C1084 a_88839_n15905# a_90245_n18620# 7.35e-19
C1085 a_101392_6405# a_101392_5639# 0.00778f
C1086 a_51711_n6241# a_51151_n6241# 0.034628f
C1087 a_40613_n14213# a_41487_n15110# 0.005903f
C1088 a_63683_n15112# a_64243_n16906# 0.035468f
C1089 a_67111_n15112# a_66029_n16906# 0.002917f
C1090 a_66551_n14215# a_66551_n15112# 0.005987f
C1091 a_104527_n6960# VDD 0.113729f
C1092 a_98299_n7865# a_99667_n6960# 2.31e-19
C1093 a_92601_n16810# a_93131_n13190# 0.032766f
C1094 a_32353_n1754# a_32913_n1754# 0.0284f
C1095 a_45706_23609# VDD 0.016884f
C1096 a_41487_n18698# a_42047_n19595# 0.0284f
C1097 a_67111_n19597# a_66551_n19597# 0.0284f
C1098 a_104527_n2435# a_105365_n2435# 0.027101f
C1099 a_110225_n7865# VDD 0.121907f
C1100 a_103997_n5150# a_104527_n3340# 0.012586f
C1101 a_92601_n21335# a_93131_n18620# 0.012586f
C1102 a_95943_n18620# a_95105_n18620# 0.042385f
C1103 a_77776_n35156# a_77776_n36322# 0.004007f
C1104 a_59763_n6241# a_60285_n6241# 0.034714f
C1105 a_49755_12380# VDD 0.061113f
C1106 a_60285_n5344# a_59411_n7138# 0.034652f
C1107 a_93131_n19525# IBPOUT 0.01873f
C1108 a_81205_n5150# a_81735_n6055# 0.035071f
C1109 a_81735_n20430# VDD 0.149203f
C1110 a_105365_n6960# a_105365_n7865# 0.005903f
C1111 a_84547_n17715# IN_POS 0.001247f
C1112 a_98829_n14095# a_99667_n14095# 0.027101f
C1113 a_98299_n16810# a_98829_n15000# 0.012586f
C1114 a_38097_n2651# a_38619_n1754# 0.0284f
C1115 a_73302_12380# VDD 0.009062f
C1116 a_46879_n19595# a_47753_n18698# 5.43e-19
C1117 a_44885_n18698# a_44885_n19595# 0.005987f
C1118 VDD I1N 1.34057f
C1119 a_112199_n2435# a_113037_n3340# 0.028522f
C1120 a_88271_n21335# VDD 0.02546f
C1121 a_61515_n34390# VDD 0.011958f
C1122 a_99667_n18620# a_99667_n19525# 0.005903f
C1123 a_77747_n27257# a_77747_n28415# 0.004047f
C1124 a_113110_n34390# a_113110_n35156# 0.00778f
C1125 a_40965_n6239# a_41487_n5342# 0.005903f
C1126 a_39179_n6239# a_38097_n7136# 0.001037f
C1127 a_96849_11614# VDD 0.011958f
C1128 a_64243_n6241# a_64243_n8035# 0.008933f
C1129 a_53145_n14215# a_54579_n15112# 0.003256f
C1130 a_82573_n2435# VDD 0.016652f
C1131 a_99667_n13190# VDD 0.02546f
C1132 a_111631_n7865# a_113037_n8770# 2.31e-19
C1133 a_95443_n33224# VDD 0.029536f
C1134 a_106501_n14095# a_107339_n15000# 0.028522f
C1135 a_85089_n35156# IN_POS 0.003316f
C1136 a_89531_n28415# a_89531_n29181# 0.00778f
C1137 a_32088_n33224# I1U 0.003282f
C1138 a_37934_7563# VDD 0.00658f
C1139 a_75602_n3060# a_75602_n4019# 0.005385f
C1140 a_54019_n18700# a_54579_n19597# 0.0284f
C1141 a_89407_n8770# a_89407_n9675# 0.024773f
C1142 a_87433_n3340# VDD 0.121044f
C1143 a_81205_n15905# a_81735_n15905# 0.028522f
C1144 a_104527_n14095# VDD 0.149203f
C1145 a_82573_n15000# a_83141_n15000# 0.027101f
C1146 a_86903_n5150# IN_POS 0.092815f
C1147 a_103997_n21335# a_105365_n21335# 7.4e-19
C1148 a_49755_11614# a_49755_10448# 0.004007f
C1149 a_46879_n3548# a_48313_n7136# 0.009477f
C1150 a_47231_n6239# a_46879_n7136# 0.534125f
C1151 a_35781_n15110# a_34699_n16904# 0.001641f
C1152 a_32353_n15110# a_32913_n16904# 0.034628f
C1153 a_35221_n14213# a_35221_n15110# 0.005987f
C1154 a_59411_n14215# a_57977_n16906# 4.66e-19
C1155 a_93969_n4245# VDD 0.023101f
C1156 a_82573_n20430# a_82573_n21335# 0.005903f
C1157 a_112199_n14095# VDD 0.121415f
C1158 a_113037_n15000# a_112199_n15000# 0.028522f
C1159 a_110225_n15000# a_111063_n15000# 0.027101f
C1160 a_109695_n16810# a_109695_n21335# 0.032645f
C1161 a_30682_n33224# a_30682_n34390# 0.004007f
C1162 a_83725_5639# a_83725_4481# 0.004047f
C1163 a_72596_n3060# OUT 3.16e-19
C1164 a_33787_n18698# a_33787_n19595# 0.005987f
C1165 a_59411_n19597# a_58851_n19597# 0.0284f
C1166 a_101641_n6055# VDD 0.472471f
C1167 a_88839_n15905# a_89407_n15905# 0.027101f
C1168 a_65117_n19597# IBNOUT -8.11e-35
C1169 a_87433_n15905# a_87433_n17715# 0.006141f
C1170 a_111631_n19525# a_111631_n20430# 0.005903f
C1171 a_54019_n4447# a_54019_n5344# 0.005987f
C1172 a_53497_n6241# a_53145_n7138# 0.070243f
C1173 a_51711_n6241# a_50629_n7138# 0.002568f
C1174 a_40613_n14213# a_40965_n16904# 0.070243f
C1175 a_65677_n14215# a_66551_n15112# 4.96e-19
C1176 a_98299_n7865# a_98829_n6960# 0.028522f
C1177 a_103997_n7865# VDD 0.393432f
C1178 a_32353_n15110# I1U 0.002649f
C1179 a_31831_n2651# a_32913_n1754# 5.37e-19
C1180 a_45138_23609# VDD 0.018612f
C1181 a_56895_n2653# a_57417_n1756# 0.0284f
C1182 a_40613_n19595# a_42047_n19595# 0.014106f
C1183 a_66551_n18700# a_66551_n19597# 0.005987f
C1184 a_63683_n19597# a_64243_n19597# 0.0284f
C1185 a_112199_n6960# VDD 0.201f
C1186 a_103997_n5150# a_103997_n4245# 0.086469f
C1187 a_105933_n1530# a_105933_n2435# 0.005903f
C1188 a_95943_n18620# a_94537_n18620# 0.002302f
C1189 a_92601_n21335# a_92601_n19525# 0.086469f
C1190 a_49795_n28415# a_49795_n29181# 0.00778f
C1191 a_35221_n4445# a_35221_n5342# 0.005987f
C1192 a_32913_n6239# a_32353_n6239# 0.035468f
C1193 a_48349_12380# VDD 0.076387f
C1194 a_47753_n14213# a_48313_n15110# 0.0284f
C1195 a_82573_n2435# a_82573_n3340# 0.005903f
C1196 a_105933_n6960# a_106501_n6960# 0.027101f
C1197 a_84547_n20430# VDD 0.399226f
C1198 a_114485_n29181# VDD 0.002225f
C1199 a_98299_n16810# a_98299_n15905# 0.086469f
C1200 a_100235_n13190# a_100235_n14095# 0.005903f
C1201 a_32353_n5342# I1U 0.002649f
C1202 a_95443_n34390# a_95443_n35156# 0.00778f
C1203 a_71896_12380# VDD 0.009062f
C1204 a_44363_n19595# a_44885_n19595# 0.0284f
C1205 a_83141_n7865# a_83141_n8770# 0.005903f
C1206 a_87433_n21335# VDD 0.150485f
C1207 a_110225_n2435# a_110225_n3340# 0.024773f
C1208 a_111631_n2435# a_113037_n3340# 2.31e-19
C1209 a_109695_n5150# a_111063_n4245# 0.002134f
C1210 a_60109_n34390# VDD 0.017204f
C1211 a_100235_n18620# a_100803_n18620# 0.027101f
C1212 a_37934_6405# a_37934_5639# 0.00778f
C1213 a_40965_n6239# a_40613_n7136# 0.534125f
C1214 a_40613_n3548# a_42047_n7136# 0.009477f
C1215 a_95443_11614# VDD 0.017204f
C1216 a_63683_n5344# a_63683_n6241# 0.005987f
C1217 a_66029_n6241# a_67111_n7138# 0.001641f
C1218 a_50629_n15112# a_51711_n16906# 0.001037f
C1219 a_51151_n14215# a_51151_n15112# 0.005987f
C1220 a_53145_n14215# a_54019_n14215# 0.004425f
C1221 a_90245_n3340# a_90245_n6960# 0.012104f
C1222 a_81735_n2435# VDD 0.121415f
C1223 a_88271_n3340# a_88271_n4245# 0.005903f
C1224 a_111631_n7865# a_112199_n7865# 0.027101f
C1225 a_98829_n13190# VDD 0.150485f
C1226 a_110225_n7865# a_110225_n8770# 0.024773f
C1227 a_90969_n36322# VDD 0.021314f
C1228 a_103997_n16810# a_105365_n15905# 0.002134f
C1229 a_104527_n14095# a_104527_n15000# 0.024773f
C1230 a_105933_n14095# a_107339_n15000# 2.31e-19
C1231 a_36562_12380# a_36562_11614# 0.00778f
C1232 a_30682_n33224# I1U 0.005416f
C1233 a_53145_n19597# a_54579_n19597# 0.014106f
C1234 a_87433_n9675# a_88271_n9675# 0.027101f
C1235 a_86903_n4245# VDD 0.393432f
C1236 a_106501_n13190# VDD 0.177586f
C1237 a_105365_n19525# a_105933_n19525# 0.027101f
C1238 a_103997_n21335# a_104527_n21335# 0.032766f
C1239 a_101392_n29181# a_101392_n30339# 0.004047f
C1240 a_108636_10448# OUT 0.02829f
C1241 a_45445_n6239# a_46879_n7136# 4.66e-19
C1242 a_34347_n14213# a_35221_n15110# 0.005903f
C1243 a_60285_n14215# a_60845_n15112# 0.0284f
C1244 a_93131_n4245# VDD 0.113729f
C1245 a_83141_n20430# a_83709_n20430# 0.027101f
C1246 a_111631_n14095# VDD 0.016652f
C1247 a_109695_n15905# a_111063_n15000# 2.31e-19
C1248 a_112199_n14095# a_112199_n15000# 0.024773f
C1249 a_113037_n15000# a_111631_n15000# 2.31e-19
C1250 a_60109_11614# a_60109_10448# 0.004007f
C1251 a_35221_n18698# a_35781_n19595# 0.0284f
C1252 a_59411_n19597# a_57977_n19597# 0.054819f
C1253 a_58851_n18700# a_58851_n19597# 0.005987f
C1254 a_98829_n1530# a_99667_n1530# 0.027101f
C1255 a_64243_n19597# IBNOUT 0.051f
C1256 a_53497_n6241# a_54019_n5344# 0.005903f
C1257 a_65677_n14215# a_66029_n16906# 0.534125f
C1258 a_98299_n9675# a_99667_n6960# 0.002134f
C1259 a_31831_n2651# a_32353_n1754# 0.0284f
C1260 a_44608_22884# VDD 0.378896f
C1261 a_40613_n19595# a_41487_n18698# 5.43e-19
C1262 a_38619_n18698# a_38619_n19595# 0.005987f
C1263 a_65677_n19597# a_66551_n19597# 5.43e-19
C1264 a_67111_n19597# a_64243_n19597# 5.37e-19
C1265 a_111631_n6960# VDD 0.01901f
C1266 a_93131_n17715# a_93131_n18620# 0.006141f
C1267 a_79182_n34390# a_79182_n35156# 0.00778f
C1268 a_34699_n6239# a_35221_n5342# 0.005903f
C1269 a_32913_n6239# a_31831_n7136# 0.001037f
C1270 a_57977_n6241# a_57417_n6241# 0.034628f
C1271 a_49755_13546# VDD 0.05845f
C1272 a_94537_n18620# IBPOUT 0.00243f
C1273 a_46879_n14213# a_48313_n15110# 0.08885f
C1274 a_83709_n2435# a_84547_n3340# 0.028522f
C1275 a_103997_n7865# a_105365_n7865# 2.31e-19
C1276 a_104527_n6960# a_104527_n7865# 0.024773f
C1277 a_83709_n19525# VDD 0.121044f
C1278 a_84547_n18620# IN_POS 0.036003f
C1279 a_46319_n18698# a_46879_n19595# 0.0284f
C1280 a_89407_n20430# VDD 0.121415f
C1281 a_111631_n2435# a_112199_n2435# 0.027101f
C1282 a_109695_n5150# a_110225_n4245# 0.012586f
C1283 a_61515_n33224# VDD 0.021515f
C1284 a_87433_n18620# IN_POS 0.00603f
C1285 a_98299_n19525# a_99667_n19525# 2.31e-19
C1286 a_98829_n18620# a_98829_n19525# 0.024773f
C1287 a_39179_n6239# a_40613_n7136# 4.66e-19
C1288 a_96849_12380# VDD 0.009062f
C1289 a_66029_n6241# a_66551_n6241# 0.034714f
C1290 a_66551_n5344# a_65677_n7138# 0.034652f
C1291 a_53497_n14215# a_53497_n16906# 0.009483f
C1292 a_50629_n15112# a_51151_n15112# 0.0284f
C1293 a_88839_n3340# a_89407_n3340# 0.027101f
C1294 a_98299_n16810# VDD 1.03823f
C1295 a_89563_n36322# VDD 0.021314f
C1296 a_103997_n16810# a_104527_n15905# 0.012586f
C1297 a_105933_n14095# a_106501_n14095# 0.027101f
C1298 a_85089_n34390# IN_POS 0.003316f
C1299 a_72596_n3060# a_72596_n4019# 0.005385f
C1300 a_50629_n19597# a_51711_n19597# 5.37e-19
C1301 a_51151_n18700# a_51151_n19597# 0.005987f
C1302 a_53145_n19597# a_54019_n18700# 5.43e-19
C1303 a_90245_n3340# VDD 0.392932f
C1304 a_88839_n8770# a_88839_n9675# 0.005903f
C1305 a_84547_n15000# a_83709_n15000# 0.028522f
C1306 a_81735_n15000# a_82573_n15000# 0.027101f
C1307 a_105933_n13190# VDD 0.02546f
C1308 a_106501_n18620# a_106501_n19525# 0.024773f
C1309 a_48349_11614# a_48349_10448# 0.004007f
C1310 a_34347_n14213# a_34699_n16904# 0.070243f
C1311 a_59411_n14215# a_60845_n15112# 0.003256f
C1312 a_95105_n3340# VDD 0.121044f
C1313 a_95105_n4245# a_95943_n6960# 0.032618f
C1314 a_81735_n20430# a_81735_n21335# 0.024773f
C1315 a_111063_n14095# VDD 0.016652f
C1316 a_109695_n15905# a_110225_n15000# 0.028522f
C1317 a_85129_6405# a_85129_5639# 0.00778f
C1318 a_34347_n19595# a_35781_n19595# 0.014106f
C1319 a_60285_n18700# a_60845_n19597# 0.0284f
C1320 a_98829_n6055# VDD 0.41764f
C1321 a_98299_n5150# a_99667_n1530# 0.002563f
C1322 a_88271_n15905# a_88839_n15905# 0.027101f
C1323 a_63683_n19597# IBNOUT 0.004735f
C1324 a_111063_n19525# a_111063_n20430# 0.005903f
C1325 a_41487_n14213# a_42047_n15110# 0.0284f
C1326 a_65677_n14215# a_64243_n16906# 4.66e-19
C1327 a_98299_n9675# a_98829_n6960# 0.012586f
C1328 a_103997_n9675# VDD 1.27279f
C1329 a_60109_n35156# a_60109_n36322# 0.004007f
C1330 a_46274_23609# VDD 0.328969f
C1331 a_38097_n19595# a_38619_n19595# 0.0284f
C1332 a_65677_n19597# a_65117_n19597# 0.0284f
C1333 a_111063_n6960# VDD 0.023101f
C1334 a_105365_n1530# a_105365_n2435# 0.005903f
C1335 a_48391_n28415# a_48391_n29181# 0.00778f
C1336 a_34699_n6239# a_34347_n7136# 0.534125f
C1337 a_34347_n3548# a_35781_n7136# 0.009477f
C1338 a_57977_n6241# a_56895_n7138# 0.002568f
C1339 a_59763_n6241# a_59411_n7138# 0.070243f
C1340 a_60285_n4447# a_60285_n5344# 0.005987f
C1341 a_48349_13546# VDD 0.073724f
C1342 a_46879_n14213# a_47753_n14213# 0.006769f
C1343 a_44363_n15110# a_45445_n16904# 0.002568f
C1344 a_44885_n14213# a_44885_n15110# 0.005987f
C1345 a_93969_n18620# IBPOUT 0.003499f
C1346 a_71864_n30339# OUT 0.003757f
C1347 a_81735_n2435# a_81735_n3340# 0.024773f
C1348 a_83141_n2435# a_84547_n3340# 2.31e-19
C1349 a_83141_n19525# VDD 0.016281f
C1350 a_105365_n6960# a_105933_n6960# 0.027101f
C1351 a_103997_n7865# a_104527_n7865# 0.028522f
C1352 a_99667_n13190# a_99667_n14095# 0.005903f
C1353 a_114485_n28415# VDD 0.002225f
C1354 a_73302_13546# VDD 0.021314f
C1355 a_63161_n2653# a_63683_n1756# 0.0284f
C1356 a_82573_n7865# a_82573_n8770# 0.005903f
C1357 a_83709_n7865# a_84547_n8770# 0.028522f
C1358 a_88839_n20430# VDD 0.016652f
C1359 a_60109_n33224# VDD 0.029536f
C1360 a_98299_n19525# a_98829_n19525# 0.028522f
C1361 a_86903_n19525# IN_POS 0.001743f
C1362 a_99667_n18620# a_100235_n18620# 0.027101f
C1363 a_45138_22884# a_45706_22884# 0.017228f
C1364 a_36530_6405# a_36530_5639# 0.00778f
C1365 a_96849_n36322# VCM 0.001273f
C1366 a_95443_12380# VDD 0.017204f
C1367 a_52585_n14215# a_53145_n14215# 0.037577f
C1368 a_83709_n1530# VDD 0.150485f
C1369 a_87433_n3340# a_87433_n4245# 0.024773f
C1370 a_86903_n4245# a_88271_n4245# 2.31e-19
C1371 a_95105_n21335# VDD 0.177586f
C1372 a_109695_n9675# a_111063_n9675# 7.4e-19
C1373 a_111063_n7865# a_111631_n7865# 0.027101f
C1374 a_90969_n35156# VDD 0.009062f
C1375 a_50629_n19597# a_51151_n19597# 0.0284f
C1376 a_89407_n2435# VDD 0.121415f
C1377 a_105365_n13190# VDD 0.02546f
C1378 a_84547_n15000# a_83141_n15000# 2.31e-19
C1379 a_81205_n15905# a_82573_n15000# 2.31e-19
C1380 a_83709_n14095# a_83709_n15000# 0.024773f
C1381 a_104527_n19525# a_105365_n19525# 0.027101f
C1382 VDD VCM 6.7918f
C1383 a_102796_n28415# a_102796_n29181# 0.00778f
C1384 a_108636_11614# OUT 0.009172f
C1385 a_47231_n6239# a_47753_n4445# 0.034714f
C1386 a_45445_n6239# a_44885_n5342# 0.00587f
C1387 a_59411_n14215# a_60285_n14215# 0.004425f
C1388 a_57417_n14215# a_57417_n15112# 0.005987f
C1389 a_56895_n15112# a_57977_n16906# 0.001037f
C1390 a_94537_n4245# a_95943_n6960# 7.35e-19
C1391 a_94537_n3340# VDD 0.016281f
C1392 a_110225_n14095# VDD 0.149203f
C1393 a_82573_n20430# a_83141_n20430# 0.027101f
C1394 a_111631_n14095# a_111631_n15000# 0.005903f
C1395 a_109695_n16810# a_110225_n17715# 0.03483f
C1396 a_61515_12380# a_61515_11614# 0.00778f
C1397 a_34347_n19595# a_35221_n18698# 5.43e-19
C1398 a_32353_n18698# a_32353_n19595# 0.005987f
C1399 a_59411_n19597# a_60845_n19597# 0.014106f
C1400 a_101641_n6960# VDD 1.18674f
C1401 a_98299_n5150# a_98829_n1530# 0.044257f
C1402 a_89407_n15000# a_89407_n15905# 0.024773f
C1403 a_112199_n19525# a_113037_n20430# 0.028522f
C1404 a_51711_n6241# a_51151_n5344# 0.00587f
C1405 a_54579_n4447# a_53145_n7138# 0.009477f
C1406 a_53497_n6241# a_54019_n4447# 0.035574f
C1407 a_40613_n14213# a_42047_n15110# 0.08885f
C1408 a_66551_n14215# a_67111_n15112# 0.0284f
C1409 a_107339_n6055# VDD 0.472471f
C1410 a_98299_n9675# a_98299_n7865# 0.086339f
C1411 a_101641_n6960# a_100803_n6960# 0.032618f
C1412 a_88839_n21335# a_89407_n21335# 0.027101f
C1413 a_45706_24195# VDD 0.016884f
C1414 a_40053_n18698# a_40613_n19595# 0.0284f
C1415 a_65117_n18700# a_65117_n19597# 0.005987f
C1416 a_65677_n19597# a_64243_n19597# 0.054819f
C1417 a_105933_n1530# a_106501_n1530# 0.027101f
C1418 a_110225_n6960# VDD 0.113729f
C1419 a_93131_n17715# a_92601_n21335# 0.03483f
C1420 w_27790_n38888# OUT 0.022266f
C1421 a_77776_n34390# a_77776_n35156# 0.00778f
C1422 a_32913_n6239# a_34347_n7136# 4.66e-19
C1423 a_59763_n6241# a_60285_n5344# 0.005903f
C1424 a_44363_n15110# a_44885_n15110# 0.0284f
C1425 a_93131_n18620# IBPOUT 0.01873f
C1426 a_47231_n14213# a_47231_n16904# 0.0089f
C1427 a_83141_n2435# a_83709_n2435# 0.027101f
C1428 a_81205_n5150# a_82573_n4245# 0.002134f
C1429 a_82573_n19525# VDD 0.016281f
C1430 a_103997_n9675# a_105365_n7865# 0.002134f
C1431 a_100235_n13190# a_100803_n13190# 0.027101f
C1432 a_61484_n29181# a_61484_n30339# 0.004047f
C1433 a_47753_n17801# a_47753_n18698# 0.005987f
C1434 a_47231_n18698# a_48313_n19595# 5.37e-19
C1435 a_83141_n7865# a_84547_n8770# 2.31e-19
C1436 a_111063_n2435# a_111631_n2435# 0.027101f
C1437 a_88271_n20430# VDD 0.016652f
C1438 a_55635_n36322# VDD 0.021314f
C1439 a_98299_n21335# a_99667_n19525# 0.002134f
C1440 a_86903_n21335# IN_POS 0.157025f
C1441 a_45706_23609# a_45706_22884# 0.006281f
C1442 a_113110_n33224# a_113110_n34390# 0.004007f
C1443 a_95443_n36322# VCM 0.001246f
C1444 a_39179_n6239# a_38619_n5342# 0.00587f
C1445 a_64243_n6241# a_63683_n6241# 0.034628f
C1446 a_83141_n1530# VDD 0.02546f
C1447 a_86903_n4245# a_87433_n4245# 0.028522f
C1448 a_88271_n3340# a_88839_n3340# 0.027101f
C1449 a_109695_n9675# a_110225_n9675# 0.032766f
C1450 a_112199_n6960# a_112199_n7865# 0.024773f
C1451 a_94537_n21335# VDD 0.02546f
C1452 a_105365_n14095# a_105933_n14095# 0.027101f
C1453 a_89563_n35156# VDD 0.009062f
C1454 a_85089_n33224# IN_POS 0.003316f
C1455 a_52585_n18700# a_53145_n19597# 0.0284f
C1456 a_53497_n18700# a_51711_n19597# 0.006457f
C1457 a_88839_n2435# VDD 0.016652f
C1458 a_88271_n8770# a_88271_n9675# 0.005903f
C1459 a_81205_n16810# a_81205_n21335# 0.032645f
C1460 a_104527_n13190# VDD 0.150485f
C1461 a_81205_n15905# a_81735_n15000# 0.028522f
C1462 a_103997_n21335# a_105365_n20430# 0.002134f
C1463 a_105933_n18620# a_105933_n19525# 0.005903f
C1464 a_49755_12380# a_49755_11614# 0.00778f
C1465 a_44885_n4445# a_44885_n5342# 0.005987f
C1466 a_46879_n3548# a_47753_n5342# 0.034652f
C1467 a_35221_n14213# a_35781_n15110# 0.0284f
C1468 a_56895_n15112# a_57417_n15112# 0.0284f
C1469 a_59763_n14215# a_59763_n16906# 0.009483f
C1470 a_93969_n3340# VDD 0.016281f
C1471 a_93131_n4245# a_93131_n6055# 0.006141f
C1472 a_94537_n4245# a_95105_n4245# 0.027101f
C1473 a_84547_n20430# a_83709_n20430# 0.028522f
C1474 a_112199_n13190# VDD 0.177586f
C1475 a_83725_6405# a_83725_5639# 0.00778f
C1476 a_31831_n19595# a_32353_n19595# 0.0284f
C1477 a_56895_n19597# a_57977_n19597# 5.37e-19
C1478 a_57417_n18700# a_57417_n19597# 0.005987f
C1479 a_59411_n19597# a_60285_n18700# 5.43e-19
C1480 a_100803_n4245# VDD 0.112244f
C1481 a_87433_n15905# a_88271_n15905# 0.027101f
C1482 a_110225_n19525# a_110225_n20430# 0.024773f
C1483 a_111631_n19525# a_113037_n20430# 2.31e-19
C1484 a_73302_12380# a_73302_11614# 0.00778f
C1485 a_101392_7563# a_101392_6405# 0.004047f
C1486 a_51151_n4447# a_51151_n5344# 0.005987f
C1487 a_40613_n14213# a_41487_n14213# 0.006769f
C1488 a_38619_n14213# a_38619_n15110# 0.005987f
C1489 a_38097_n15110# a_39179_n16904# 0.002568f
C1490 a_65677_n14215# a_67111_n15112# 0.003256f
C1491 a_101641_n6960# a_100235_n6960# 7.35e-19
C1492 a_61515_n34390# a_61515_n35156# 0.00778f
C1493 a_45138_24195# VDD 0.017047f
C1494 a_66551_n18700# a_67111_n19597# 0.0284f
C1495 a_109695_n7865# VDD 0.401168f
C1496 a_103997_n5150# a_105365_n2435# 0.002134f
C1497 a_104527_n1530# a_104527_n2435# 0.024773f
C1498 a_32128_n30339# I1U 5.57e-19
C1499 a_92601_n19525# IBPOUT 0.007901f
C1500 a_46319_n14213# a_46879_n14213# 0.0284f
C1501 a_71864_n29181# OUT 0.001942f
C1502 a_81205_n5150# a_81735_n4245# 0.012586f
C1503 a_104527_n6960# a_105365_n6960# 0.027101f
C1504 a_81735_n19525# VDD 0.121044f
C1505 a_107339_n6960# a_107339_n8770# 0.012104f
C1506 a_103997_n9675# a_104527_n7865# 0.012586f
C1507 a_98829_n13190# a_98829_n14095# 0.024773f
C1508 a_98299_n16810# a_99667_n14095# 0.002134f
C1509 a_95443_n33224# a_95443_n34390# 0.004007f
C1510 a_47231_n18698# a_47753_n18698# 0.0284f
C1511 a_81735_n7865# a_81735_n8770# 0.024773f
C1512 a_83141_n7865# a_83709_n7865# 0.027101f
C1513 a_87433_n20430# VDD 0.149203f
C1514 a_112199_n1530# a_112199_n2435# 0.024773f
C1515 a_109695_n5150# a_111063_n3340# 0.002134f
C1516 a_101641_n18620# a_101641_n20430# 0.012104f
C1517 a_98829_n18620# a_99667_n18620# 0.027101f
C1518 a_98299_n21335# a_98829_n19525# 0.012586f
C1519 a_54229_n36322# VDD 0.021314f
C1520 a_38619_n4445# a_38619_n5342# 0.005987f
C1521 a_40613_n3548# a_41487_n5342# 0.034652f
C1522 a_40965_n6239# a_41487_n4445# 0.034714f
C1523 a_66029_n6241# a_65677_n7138# 0.070243f
C1524 a_64243_n6241# a_63161_n7138# 0.002568f
C1525 a_66551_n4447# a_66551_n5344# 0.005987f
C1526 a_96849_13546# VDD 0.024605f
C1527 a_53497_n14215# a_54579_n15112# 5.37e-19
C1528 a_54019_n13318# a_54019_n14215# 0.005987f
C1529 a_82573_n1530# VDD 0.02546f
C1530 a_93969_n21335# VDD 0.02546f
C1531 a_110225_n7865# a_111063_n7865# 0.027101f
C1532 a_103997_n16810# a_105365_n15000# 0.002134f
C1533 a_106501_n13190# a_106501_n14095# 0.024773f
C1534 a_90969_n34390# VDD 0.009062f
C1535 a_42047_n8930# a_41487_n8930# 0.0284f
C1536 a_88271_n2435# VDD 0.016652f
C1537 a_71896_n36322# OUT 0.001027f
C1538 a_88839_n8770# a_89407_n8770# 0.027101f
C1539 a_103997_n16810# VDD 1.04258f
C1540 a_83141_n14095# a_83141_n15000# 0.005903f
C1541 a_103997_n21335# a_104527_n20430# 0.012586f
C1542 a_101392_n28415# a_101392_n29181# 0.00778f
C1543 a_66058_5639# a_66058_4481# 0.004047f
C1544 a_108636_12380# OUT 0.003165f
C1545 a_45445_n6239# a_47231_n6239# 0.012473f
C1546 a_46879_n3548# a_46879_n7136# 0.00969f
C1547 a_34347_n14213# a_35781_n15110# 0.08885f
C1548 a_58851_n14215# a_59411_n14215# 0.037577f
C1549 a_93131_n3340# VDD 0.121044f
C1550 a_81735_n20430# a_82573_n20430# 0.027101f
C1551 a_83709_n19525# a_83709_n20430# 0.024773f
C1552 a_84547_n20430# a_83141_n20430# 2.31e-19
C1553 a_111631_n13190# VDD 0.02546f
C1554 a_111063_n14095# a_111063_n15000# 0.005903f
C1555 a_60109_12380# a_60109_11614# 0.00778f
C1556 a_33787_n18698# a_34347_n19595# 0.0284f
C1557 a_56895_n19597# a_57417_n19597# 0.0284f
C1558 a_100235_n4245# VDD 0.023105f
C1559 a_88839_n15000# a_88839_n15905# 0.005903f
C1560 a_65677_n19597# IBNOUT 0.006327f
C1561 a_32128_4481# I1U 5.57e-19
C1562 a_111631_n19525# a_112199_n19525# 0.027101f
C1563 a_42442_n35156# a_42442_n36322# 0.004007f
C1564 a_51711_n6241# a_53497_n6241# 0.012473f
C1565 a_53145_n3550# a_53145_n7138# 0.00969f
C1566 a_40965_n14213# a_40965_n16904# 0.0089f
C1567 a_38097_n15110# a_38619_n15110# 0.0284f
C1568 a_63161_n15112# a_64243_n16906# 0.001037f
C1569 a_63683_n14215# a_63683_n15112# 0.005987f
C1570 a_65677_n14215# a_66551_n14215# 0.004425f
C1571 a_104527_n6055# VDD 0.41764f
C1572 a_98829_n6055# a_98829_n6960# 0.006141f
C1573 a_88271_n21335# a_88839_n21335# 0.027101f
C1574 a_32353_n14213# I1U 0.002649f
C1575 a_85089_11614# a_85089_10448# 0.004007f
C1576 a_46274_24920# VDD 0.165281f
C1577 a_51711_n8932# a_54019_n8932# 0.0284f
C1578 a_41487_n17801# a_41487_n18698# 0.005987f
C1579 a_40965_n18698# a_42047_n19595# 5.37e-19
C1580 a_65677_n19597# a_67111_n19597# 0.014106f
C1581 a_103997_n5150# a_104527_n2435# 0.012586f
C1582 a_105365_n1530# a_105933_n1530# 0.027101f
C1583 a_95943_n18620# a_95943_n17715# 0.088786f
C1584 a_32913_n6239# a_32353_n5342# 0.00587f
C1585 a_43848_10448# VDD 0.023325f
C1586 a_30724_n30339# I1U 0.004931f
C1587 a_60845_n4447# a_59411_n7138# 0.009477f
C1588 a_57977_n6241# a_57417_n5344# 0.00587f
C1589 a_59763_n6241# a_60285_n4447# 0.035574f
C1590 a_92601_n21335# IBPOUT 0.2259f
C1591 a_82573_n2435# a_83141_n2435# 0.027101f
C1592 a_83709_n18620# VDD 0.112244f
C1593 a_103997_n7865# a_105365_n6960# 2.31e-19
C1594 a_98299_n16810# a_98829_n14095# 0.012586f
C1595 a_114485_n27257# VDD 0.002225f
C1596 a_99667_n13190# a_100235_n13190# 0.027101f
C1597 a_32353_n4445# I1U 0.002649f
C1598 a_60080_n29181# a_60080_n30339# 0.004047f
C1599 a_71896_13546# VDD 0.021314f
C1600 a_44363_n19595# a_44885_n18698# 0.0284f
C1601 a_47231_n18698# a_46879_n19595# 0.053799f
C1602 a_81205_n9675# a_82573_n9675# 0.002563f
C1603 a_90245_n20430# VDD 0.399226f
C1604 a_110225_n2435# a_111063_n2435# 0.027101f
C1605 a_109695_n5150# a_110225_n3340# 0.012586f
C1606 a_98299_n19525# a_99667_n18620# 2.31e-19
C1607 a_55635_n35156# VDD 0.009062f
C1608 a_87433_n17715# IN_POS 0.005369f
C1609 a_44608_22884# a_45706_22884# 1.81e-19
C1610 a_45138_23609# a_45138_22884# 0.006281f
C1611 a_40613_n3548# a_40613_n7136# 0.00969f
C1612 a_66029_n6241# a_66551_n5344# 0.005903f
C1613 a_51711_n14215# a_51711_n16906# 0.009307f
C1614 a_53497_n14215# a_54019_n14215# 0.0284f
C1615 a_81735_n1530# VDD 0.150485f
C1616 a_90245_n3340# a_89407_n3340# 0.028522f
C1617 a_87433_n3340# a_88271_n3340# 0.027101f
C1618 a_93131_n21335# VDD 0.150485f
C1619 a_111631_n6960# a_111631_n7865# 0.005903f
C1620 a_89563_n34390# VDD 0.009062f
C1621 a_104527_n14095# a_105365_n14095# 0.027101f
C1622 a_103997_n16810# a_104527_n15000# 0.012586f
C1623 a_41487_n8033# a_41487_n8930# 0.005987f
C1624 a_53497_n18700# a_54579_n19597# 5.37e-19
C1625 a_54019_n17803# a_54019_n18700# 0.005987f
C1626 a_87433_n2435# VDD 0.121415f
C1627 a_87433_n8770# a_87433_n9675# 0.024773f
C1628 a_81205_n16810# a_81735_n17715# 0.035071f
C1629 a_100803_n21335# VDD 0.150485f
C1630 a_105365_n18620# a_105365_n19525# 0.005903f
C1631 a_48349_12380# a_48349_11614# 0.00778f
C1632 a_48313_n4445# a_47753_n4445# 0.0284f
C1633 a_32353_n14213# a_32353_n15110# 0.005987f
C1634 a_31831_n15110# a_32913_n16904# 0.002568f
C1635 a_34347_n14213# a_35221_n14213# 0.006769f
C1636 a_92601_n4245# VDD 0.393432f
C1637 a_93969_n4245# a_94537_n4245# 0.027101f
C1638 a_111063_n13190# VDD 0.02546f
C1639 a_112199_n14095# a_113037_n15000# 0.028522f
C1640 a_114485_n29181# a_114485_n30339# 0.004047f
C1641 a_48313_n8930# a_47753_n8930# 0.0284f
C1642 a_58851_n18700# a_59411_n19597# 0.0284f
C1643 a_59763_n18700# a_57977_n19597# 0.006457f
C1644 a_85129_4481# IN_POS 6.24e-19
C1645 a_99667_n4245# VDD 0.012916f
C1646 a_30724_4481# I1U 0.004931f
C1647 a_109695_n21335# a_111063_n21335# 7.4e-19
C1648 a_71896_12380# a_71896_11614# 0.00778f
C1649 a_53145_n3550# a_54019_n5344# 0.030444f
C1650 a_54579_n4447# a_54019_n4447# 0.0284f
C1651 a_40053_n14213# a_40613_n14213# 0.0284f
C1652 a_66029_n14215# a_66029_n16906# 0.009483f
C1653 a_63161_n15112# a_63683_n15112# 0.0284f
C1654 VDD IN_NEG 2.89387f
C1655 OUT IN_POS 0.390657f
C1656 a_107339_n6960# VDD 1.18674f
C1657 a_89407_n20430# a_89407_n21335# 0.024773f
C1658 a_31831_n15110# I1U 0.008518f
C1659 a_60109_n34390# a_60109_n35156# 0.00778f
C1660 a_45706_24920# VDD 0.030148f
C1661 a_51711_n8932# a_52585_n8932# 0.001405f
C1662 a_40965_n18698# a_41487_n18698# 0.0284f
C1663 a_65677_n19597# a_66551_n18700# 5.43e-19
C1664 a_63161_n19597# a_64243_n19597# 5.37e-19
C1665 a_63683_n18700# a_63683_n19597# 0.005987f
C1666 a_109695_n9675# VDD 1.60209f
C1667 a_95443_11614# a_95443_10448# 0.004007f
C1668 a_34347_n3548# a_35221_n5342# 0.034652f
C1669 a_34699_n6239# a_35221_n4445# 0.034714f
C1670 a_32353_n4445# a_32353_n5342# 0.005987f
C1671 a_42442_10448# VDD 0.029536f
C1672 a_32128_n29181# I1U 5.57e-19
C1673 a_57417_n4447# a_57417_n5344# 0.005987f
C1674 a_47231_n14213# a_48313_n15110# 5.37e-19
C1675 a_47753_n13316# a_47753_n14213# 0.005987f
C1676 a_71864_n28415# OUT 0.001942f
C1677 a_83141_n18620# VDD 0.023105f
C1678 a_103997_n7865# a_104527_n6960# 0.028522f
C1679 a_35781_n8930# a_35221_n8930# 0.0284f
C1680 a_47231_n18698# a_46319_n18698# 5.43e-19
C1681 a_81205_n9675# a_81735_n9675# 0.044257f
C1682 a_82573_n7865# a_83141_n7865# 0.027101f
C1683 a_89407_n19525# VDD 0.121044f
C1684 a_111631_n1530# a_111631_n2435# 0.005903f
C1685 a_109695_n5150# a_109695_n4245# 0.086469f
C1686 a_54229_n35156# VDD 0.009062f
C1687 a_98299_n19525# a_98829_n18620# 0.028522f
C1688 a_45138_23609# a_45706_23609# 0.017228f
C1689 a_44608_22884# a_45138_22884# 0.017843f
C1690 a_39179_n6239# a_40965_n6239# 0.012473f
C1691 a_95443_13546# VDD 0.029536f
C1692 w_27790_n38888# IBNOUT 0.022266f
C1693 a_50629_n15112# a_51151_n14215# 0.0284f
C1694 a_53497_n14215# a_53145_n14215# 0.062551f
C1695 a_81205_n5150# VDD 0.916148f
C1696 a_89407_n2435# a_89407_n3340# 0.024773f
C1697 a_86903_n4245# a_88271_n3340# 2.31e-19
C1698 a_90245_n3340# a_88839_n3340# 2.31e-19
C1699 a_95105_n20430# VDD 0.121415f
C1700 a_109695_n9675# a_111063_n8770# 0.002134f
C1701 a_105933_n13190# a_105933_n14095# 0.005903f
C1702 a_103997_n16810# a_103997_n15905# 0.086469f
C1703 a_40613_n8930# a_41487_n8930# 5.43e-19
C1704 a_53497_n18700# a_54019_n18700# 0.0284f
C1705 a_51711_n18700# a_51711_n19597# 0.006457f
C1706 a_71896_n35156# OUT 0.001027f
C1707 a_88271_n8770# a_88839_n8770# 0.027101f
C1708 a_100235_n21335# VDD 0.02546f
C1709 a_82573_n14095# a_82573_n15000# 0.005903f
C1710 a_105933_n18620# a_106501_n18620# 0.027101f
C1711 a_67462_6405# a_67462_5639# 0.00778f
C1712 a_47753_n3548# a_47753_n4445# 0.005987f
C1713 a_48313_n4445# a_47231_n6239# 0.001641f
C1714 a_44885_n4445# a_45445_n6239# 0.034628f
C1715 a_34699_n14213# a_34699_n16904# 0.0089f
C1716 a_31831_n15110# a_32353_n15110# 0.0284f
C1717 a_59763_n14215# a_60845_n15112# 5.37e-19
C1718 a_60285_n13318# a_60285_n14215# 0.005987f
C1719 a_95943_n3340# VDD 0.392932f
C1720 a_95105_n3340# a_95105_n4245# 0.024773f
C1721 a_83141_n19525# a_83141_n20430# 0.005903f
C1722 a_110225_n13190# VDD 0.150485f
C1723 a_111631_n14095# a_113037_n15000# 2.31e-19
C1724 a_110225_n14095# a_110225_n15000# 0.024773f
C1725 a_109695_n16810# a_111063_n15905# 0.002134f
C1726 a_47753_n8033# a_47753_n8930# 0.005987f
C1727 a_34699_n18698# a_35781_n19595# 5.37e-19
C1728 a_35221_n17801# a_35221_n18698# 0.005987f
C1729 a_98829_n4245# VDD 0.137705f
C1730 a_94537_n9675# a_95105_n9675# 0.027101f
C1731 a_88271_n15000# a_88271_n15905# 0.005903f
C1732 a_32128_5639# I1U 5.57e-19
C1733 a_90245_n15000# a_90245_n18620# 0.012104f
C1734 a_63683_n18700# IBNOUT 0.004735f
C1735 a_109695_n21335# a_110225_n21335# 0.032766f
C1736 a_111063_n19525# a_111631_n19525# 0.027101f
C1737 a_43848_n34390# a_43848_n35156# 0.00778f
C1738 a_54579_n4447# a_53497_n6241# 0.002917f
C1739 a_54019_n3550# a_54019_n4447# 0.005987f
C1740 a_51151_n4447# a_51711_n6241# 0.035468f
C1741 a_65117_n14215# a_65677_n14215# 0.037577f
C1742 a_106501_n4245# VDD 0.112244f
C1743 a_87433_n21335# a_88271_n21335# 0.027101f
C1744 a_55601_n30339# VDD 0.00658f
C1745 a_83683_11614# a_83683_10448# 0.004007f
C1746 a_45138_24920# VDD 0.030305f
C1747 a_54579_n8932# a_54019_n8932# 0.0284f
C1748 a_38097_n19595# a_38619_n18698# 0.0284f
C1749 a_40965_n18698# a_40613_n19595# 0.053799f
C1750 a_63161_n19597# a_63683_n19597# 0.0284f
C1751 a_113037_n6055# VDD 0.509696f
C1752 a_64243_n8932# IBNOUT 0.001252f
C1753 a_104527_n1530# a_105365_n1530# 0.027101f
C1754 a_48391_n27257# a_48391_n28415# 0.004047f
C1755 a_77776_n33224# a_77776_n34390# 0.004007f
C1756 a_34347_n3548# a_34347_n7136# 0.00969f
C1757 a_30724_n29181# I1U 0.004931f
C1758 a_43848_11614# VDD 0.013768f
C1759 a_59411_n3550# a_59411_n7138# 0.00969f
C1760 a_57977_n6241# a_59763_n6241# 0.012473f
C1761 a_93131_n17715# IBPOUT 0.026429f
C1762 a_47753_n13316# a_46879_n14213# 8.45e-19
C1763 a_47231_n14213# a_47753_n14213# 0.0284f
C1764 a_45445_n14213# a_45445_n16904# 0.008933f
C1765 a_83709_n1530# a_83709_n2435# 0.024773f
C1766 a_81735_n2435# a_82573_n2435# 0.027101f
C1767 a_81205_n5150# a_82573_n3340# 0.002134f
C1768 a_82573_n18620# VDD 0.012916f
C1769 a_103997_n9675# a_105365_n6960# 0.002134f
C1770 a_98829_n13190# a_99667_n13190# 0.027101f
C1771 a_61484_n28415# a_61484_n29181# 0.00778f
C1772 a_35221_n8033# a_35221_n8930# 0.005987f
C1773 a_57977_n8932# a_60285_n8932# 0.0284f
C1774 a_45797_n18698# a_46879_n19595# 5.37e-19
C1775 a_46319_n17801# a_46319_n18698# 0.005987f
C1776 a_83709_n6960# a_83709_n7865# 0.024773f
C1777 a_88839_n19525# VDD 0.016281f
C1778 a_98299_n21335# a_99667_n18620# 0.002134f
C1779 a_55635_n34390# VDD 0.009062f
C1780 a_44608_22884# a_45706_23609# 1.81e-19
C1781 a_42047_n4445# a_41487_n4445# 0.0284f
C1782 a_67111_n4447# a_65677_n7138# 0.009477f
C1783 a_64243_n6241# a_63683_n5344# 0.00587f
C1784 a_66029_n6241# a_66551_n4447# 0.035574f
C1785 a_53497_n14215# a_52585_n14215# 5.43e-19
C1786 a_86903_n4245# a_87433_n3340# 0.028522f
C1787 a_86903_n5150# a_86903_n9675# 0.032645f
C1788 a_94537_n20430# VDD 0.016652f
C1789 a_109695_n9675# a_110225_n8770# 0.012586f
C1790 a_111063_n6960# a_111063_n7865# 0.005903f
C1791 a_90969_n33224# VDD 0.021515f
C1792 a_40613_n8930# a_40053_n8930# 0.0284f
C1793 a_50629_n19597# a_51151_n18700# 0.0284f
C1794 a_53497_n18700# a_53145_n19597# 0.053799f
C1795 a_90245_n8770# a_89407_n8770# 0.028522f
C1796 a_89407_n1530# VDD 0.150485f
C1797 a_99667_n21335# VDD 0.02546f
C1798 a_83709_n14095# a_84547_n15000# 0.028522f
C1799 a_103997_n19525# a_105365_n19525# 2.31e-19
C1800 a_104527_n18620# a_104527_n19525# 0.024773f
C1801 a_108636_13546# OUT 0.003165f
C1802 a_49755_13546# a_49755_12380# 0.004007f
C1803 a_46879_n3548# a_47753_n4445# 0.005903f
C1804 a_33787_n14213# a_34347_n14213# 0.0284f
C1805 a_59763_n14215# a_60285_n14215# 0.0284f
C1806 a_57977_n14215# a_57977_n16906# 0.009307f
C1807 a_95105_n2435# VDD 0.121415f
C1808 a_93131_n4245# a_93969_n4245# 0.027101f
C1809 a_109695_n16810# VDD 1.40063f
C1810 a_109695_n16810# a_110225_n15905# 0.012586f
C1811 a_111631_n14095# a_112199_n14095# 0.027101f
C1812 a_113081_n29181# a_113081_n30339# 0.004047f
C1813 a_46879_n8930# a_47753_n8930# 5.43e-19
C1814 a_34699_n18698# a_35221_n18698# 0.0284f
C1815 a_60285_n17803# a_60285_n18700# 0.005987f
C1816 a_59763_n18700# a_60845_n19597# 5.37e-19
C1817 a_85129_5639# IN_POS 6.24e-19
C1818 a_100803_n3340# VDD 0.121044f
C1819 a_30724_5639# I1U 0.004931f
C1820 a_63161_n19597# IBNOUT 0.008659f
C1821 a_88839_n15000# a_89407_n15000# 0.027101f
C1822 a_112199_n18620# a_112199_n19525# 0.024773f
C1823 a_53145_n3550# a_54019_n4447# 4.96e-19
C1824 a_40965_n14213# a_42047_n15110# 5.37e-19
C1825 a_41487_n13316# a_41487_n14213# 0.005987f
C1826 a_105933_n4245# VDD 0.023105f
C1827 a_98829_n6055# a_98299_n9675# 0.035071f
C1828 a_88839_n20430# a_88839_n21335# 0.005903f
C1829 a_114485_5639# a_114485_4481# 0.004047f
C1830 a_54019_n8035# a_54019_n8932# 0.005987f
C1831 a_51151_n8932# a_51711_n8932# 0.0284f
C1832 a_44608_24195# VDD 0.378914f
C1833 a_40965_n18698# a_40053_n18698# 5.43e-19
C1834 a_66029_n18700# a_64243_n19597# 0.006457f
C1835 a_65117_n18700# a_65677_n19597# 0.0284f
C1836 a_110225_n6055# VDD 0.41764f
C1837 a_103997_n5150# a_105365_n1530# 0.002563f
C1838 a_95105_n15905# a_95943_n18620# 0.032618f
C1839 a_96849_12380# a_96849_11614# 0.00778f
C1840 a_32913_n6239# a_34699_n6239# 0.012473f
C1841 a_60845_n4447# a_60285_n4447# 0.0284f
C1842 a_42442_11614# VDD 0.017204f
C1843 a_59411_n3550# a_60285_n5344# 0.030444f
C1844 a_32128_n28415# I1U 5.57e-19
C1845 a_44363_n15110# a_44885_n14213# 0.0284f
C1846 a_47231_n14213# a_46879_n14213# 0.16936f
C1847 a_81205_n5150# a_81735_n3340# 0.012586f
C1848 a_81735_n18620# VDD 0.137705f
C1849 a_103997_n9675# a_104527_n6960# 0.012586f
C1850 a_98299_n16810# a_99667_n13190# 0.002563f
C1851 a_108602_n30339# VDD 0.00658f
C1852 a_34347_n8930# a_35221_n8930# 5.43e-19
C1853 a_67422_10448# VDD 0.05812f
C1854 a_57977_n8932# a_58851_n8932# 0.001405f
C1855 a_45445_n18698# a_46879_n19595# 1.57e-19
C1856 a_45797_n18698# a_46319_n18698# 0.0284f
C1857 a_48313_n17801# a_48313_n19595# 0.005987f
C1858 a_81735_n7865# a_82573_n7865# 0.027101f
C1859 a_88271_n19525# VDD 0.016281f
C1860 a_111063_n1530# a_111063_n2435# 0.005903f
C1861 a_54229_n34390# VDD 0.009062f
C1862 a_98299_n21335# a_98829_n18620# 0.012586f
C1863 a_46274_23609# a_45706_23609# 0.018349f
C1864 a_44608_22884# a_45138_23609# 0.017843f
C1865 a_38619_n4445# a_39179_n6239# 0.034628f
C1866 a_41487_n3548# a_41487_n4445# 0.005987f
C1867 a_42047_n4445# a_40965_n6239# 0.001641f
C1868 a_90969_10448# VDD 0.021515f
C1869 a_63683_n4447# a_63683_n5344# 0.005987f
C1870 a_52585_n13318# a_52585_n14215# 0.005987f
C1871 a_52063_n14215# a_53145_n14215# 0.00117f
C1872 a_88839_n2435# a_88839_n3340# 0.005903f
C1873 a_93969_n20430# VDD 0.016652f
C1874 a_111631_n6960# a_112199_n6960# 0.027101f
C1875 a_105365_n13190# a_105365_n14095# 0.005903f
C1876 a_89563_n33224# VDD 0.021515f
C1877 a_40053_n8033# a_40053_n8930# 0.005987f
C1878 a_53497_n18700# a_52585_n18700# 5.43e-19
C1879 a_88839_n1530# VDD 0.02546f
C1880 a_71896_n34390# OUT 0.001027f
C1881 a_87433_n8770# a_88271_n8770# 0.027101f
C1882 a_89407_n7865# a_89407_n8770# 0.024773f
C1883 a_90245_n8770# a_88839_n8770# 2.31e-19
C1884 a_98829_n21335# VDD 0.150485f
C1885 a_84547_n8770# IN_POS 0.004986f
C1886 a_81735_n14095# a_81735_n15000# 0.024773f
C1887 a_83141_n14095# a_84547_n15000# 2.31e-19
C1888 a_103997_n19525# a_104527_n19525# 0.028522f
C1889 a_105365_n18620# a_105933_n18620# 0.027101f
C1890 a_66058_6405# a_66058_5639# 0.00778f
C1891 a_46879_n3548# a_47231_n6239# 0.070243f
C1892 a_56895_n15112# a_57417_n14215# 0.0284f
C1893 a_59763_n14215# a_59411_n14215# 0.062551f
C1894 a_94537_n3340# a_94537_n4245# 0.005903f
C1895 a_94537_n2435# VDD 0.016652f
C1896 a_106501_n21335# VDD 0.150485f
C1897 a_83709_n19525# a_84547_n20430# 0.028522f
C1898 a_82573_n19525# a_82573_n20430# 0.005903f
C1899 a_87433_n9675# IN_POS 0.00603f
C1900 a_83725_7563# a_83725_6405# 0.004047f
C1901 a_46879_n8930# a_46319_n8930# 0.0284f
C1902 a_31831_n19595# a_32353_n18698# 0.0284f
C1903 a_34699_n18698# a_34347_n19595# 0.053799f
C1904 a_59763_n18700# a_60285_n18700# 0.0284f
C1905 a_57977_n18700# a_57977_n19597# 0.006457f
C1906 a_100235_n3340# VDD 0.016281f
C1907 a_93969_n9675# a_94537_n9675# 0.027101f
C1908 a_32128_6405# I1U 5.57e-19
C1909 a_86903_n15905# a_88271_n15905# 2.31e-19
C1910 a_87433_n15000# a_87433_n15905# 0.024773f
C1911 a_110225_n19525# a_111063_n19525# 0.027101f
C1912 a_42442_n34390# a_42442_n35156# 0.00778f
C1913 a_53145_n3550# a_53497_n6241# 0.534125f
C1914 a_40965_n14213# a_41487_n14213# 0.0284f
C1915 a_41487_n13316# a_40613_n14213# 8.45e-19
C1916 a_39179_n14213# a_39179_n16904# 0.008933f
C1917 a_66029_n14215# a_67111_n15112# 5.37e-19
C1918 a_66551_n13318# a_66551_n14215# 0.005987f
C1919 a_105365_n4245# VDD 0.012916f
C1920 a_55601_n29181# VDD 0.034176f
C1921 a_85089_12380# a_85089_11614# 0.00778f
C1922 a_54579_n8932# a_51711_n8932# 5.37e-19
C1923 a_53145_n8932# a_54019_n8932# 5.43e-19
C1924 a_39531_n18698# a_40613_n19595# 5.37e-19
C1925 a_40053_n17801# a_40053_n18698# 0.005987f
C1926 a_113037_n6960# VDD 1.28333f
C1927 a_103997_n5150# a_104527_n1530# 0.044257f
C1928 a_94537_n15905# a_95943_n18620# 7.35e-19
C1929 a_30724_n28415# I1U 0.004931f
C1930 a_35781_n4445# a_35221_n4445# 0.0284f
C1931 a_57417_n4447# a_57977_n6241# 0.035468f
C1932 a_60285_n3550# a_60285_n4447# 0.005987f
C1933 a_60845_n4447# a_59763_n6241# 0.002917f
C1934 a_43848_12380# VDD 0.010872f
C1935 a_71864_n27257# OUT 0.001942f
C1936 a_81205_n5150# a_81205_n4245# 0.086339f
C1937 a_83141_n1530# a_83141_n2435# 0.005903f
C1938 a_81205_n19525# VDD 0.399575f
C1939 a_103997_n9675# a_103997_n7865# 0.086339f
C1940 a_107339_n6960# a_106501_n6960# 0.032618f
C1941 a_98299_n16810# a_98829_n13190# 0.044257f
C1942 a_60080_n28415# a_60080_n29181# 0.00778f
C1943 a_34347_n8930# a_33787_n8930# 0.0284f
C1944 a_60845_n8932# a_60285_n8932# 0.0284f
C1945 a_66016_10448# VDD 0.073394f
C1946 a_47231_n18698# a_47753_n17801# 0.0284f
C1947 a_81205_n9675# a_82573_n8770# 0.002134f
C1948 a_83141_n6960# a_83141_n7865# 0.005903f
C1949 a_87433_n19525# VDD 0.121044f
C1950 a_111631_n1530# a_112199_n1530# 0.027101f
C1951 a_101641_n18620# a_100803_n18620# 0.032618f
C1952 a_98299_n21335# a_98299_n19525# 0.086339f
C1953 a_46274_23609# a_45138_23609# 1.92e-19
C1954 a_45706_24195# a_45706_23609# 0.008552f
C1955 a_40613_n3548# a_41487_n4445# 0.005903f
C1956 a_89563_10448# VDD 0.021515f
C1957 a_64243_n6241# a_66029_n6241# 0.012473f
C1958 a_65677_n3550# a_65677_n7138# 0.00969f
C1959 a_85089_10448# IN_POS 0.003316f
C1960 a_51711_n14215# a_53145_n14215# 5.12e-19
C1961 a_54579_n13318# a_54579_n15112# 0.005987f
C1962 a_52063_n14215# a_52585_n14215# 0.0284f
C1963 a_86903_n5150# a_87433_n6055# 0.035071f
C1964 a_93131_n20430# VDD 0.149203f
C1965 a_109695_n7865# a_111063_n7865# 2.31e-19
C1966 a_110225_n6960# a_110225_n7865# 0.024773f
C1967 a_85089_n36322# VDD 0.05845f
C1968 a_105933_n13190# a_106501_n13190# 0.027101f
C1969 a_48391_5639# a_48391_4481# 0.004047f
C1970 a_41487_n8033# a_42047_n8930# 0.0284f
C1971 a_64243_n8932# a_66551_n8932# 0.0284f
C1972 a_52585_n17803# a_52585_n18700# 0.005987f
C1973 a_52063_n18700# a_53145_n19597# 5.37e-19
C1974 a_88271_n1530# VDD 0.02546f
C1975 a_100803_n20430# VDD 0.121415f
C1976 a_81205_n16810# a_82573_n15905# 0.002134f
C1977 a_83141_n14095# a_83709_n14095# 0.027101f
C1978 a_103997_n21335# a_105365_n19525# 0.002134f
C1979 a_101392_n27257# a_101392_n28415# 0.004047f
C1980 a_48349_13546# a_48349_12380# 0.004007f
C1981 a_34699_n14213# a_35781_n15110# 5.37e-19
C1982 a_35221_n13316# a_35221_n14213# 0.005987f
C1983 a_59763_n14215# a_58851_n14215# 5.43e-19
C1984 a_93969_n2435# VDD 0.016652f
C1985 a_105933_n21335# VDD 0.02546f
C1986 a_83141_n19525# a_84547_n20430# 2.31e-19
C1987 a_111063_n14095# a_111631_n14095# 0.027101f
C1988 w_27790_n38888# IBPOUT 0.022266f
C1989 a_114485_n28415# a_114485_n29181# 0.00778f
C1990 a_46319_n8033# a_46319_n8930# 0.005987f
C1991 a_47753_n8033# a_48313_n8930# 0.0284f
C1992 a_34699_n18698# a_33787_n18698# 5.43e-19
C1993 a_59763_n18700# a_59411_n19597# 0.053799f
C1994 a_56895_n19597# a_57417_n18700# 0.0284f
C1995 a_85129_6405# IN_POS 6.24e-19
C1996 a_95105_n8770# a_95105_n9675# 0.024773f
C1997 a_99667_n3340# VDD 0.016281f
C1998 a_30724_6405# I1U 0.004931f
C1999 a_88271_n15000# a_88839_n15000# 0.027101f
C2000 a_66029_n18700# IBNOUT 0.001124f
C2001 a_86903_n15905# a_87433_n15905# 0.028522f
C2002 a_111631_n18620# a_111631_n19525# 0.005903f
C2003 a_109695_n21335# a_111063_n20430# 0.002134f
C2004 a_53145_n3550# a_51711_n6241# 4.66e-19
C2005 a_38097_n15110# a_38619_n14213# 0.0284f
C2006 a_40965_n14213# a_40613_n14213# 0.16936f
C2007 a_66029_n14215# a_66551_n14215# 0.0284f
C2008 a_64243_n14215# a_64243_n16906# 0.009307f
C2009 a_101641_n6960# a_101641_n6055# 0.088786f
C2010 a_104527_n4245# VDD 0.137705f
C2011 a_54197_n29181# VDD 0.029136f
C2012 a_88271_n20430# a_88271_n21335# 0.005903f
C2013 a_60109_n33224# a_60109_n34390# 0.004007f
C2014 a_113081_5639# a_113081_4481# 0.004047f
C2015 a_53145_n8932# a_52585_n8932# 0.0284f
C2016 a_42047_n17801# a_42047_n19595# 0.005987f
C2017 a_39179_n18698# a_40613_n19595# 1.57e-19
C2018 a_39531_n18698# a_40053_n18698# 0.0284f
C2019 a_66029_n18700# a_67111_n19597# 5.37e-19
C2020 a_66551_n17803# a_66551_n18700# 0.005987f
C2021 a_112199_n4245# VDD 0.128099f
C2022 a_93131_n15905# a_93131_n17715# 0.006141f
C2023 a_94537_n15905# a_95105_n15905# 0.027101f
C2024 a_95443_12380# a_95443_11614# 0.00778f
C2025 a_35221_n3548# a_35221_n4445# 0.005987f
C2026 a_35781_n4445# a_34699_n6239# 0.001641f
C2027 a_32353_n4445# a_32913_n6239# 0.034628f
C2028 a_59411_n3550# a_60285_n4447# 4.96e-19
C2029 a_42442_12380# VDD 0.017204f
C2030 a_94537_n15905# IBPOUT 0.00243f
C2031 a_46319_n13316# a_46319_n14213# 0.005987f
C2032 a_45797_n14213# a_46879_n14213# 0.011365f
C2033 a_81205_n21335# VDD 1.33016f
C2034 a_107339_n6960# a_105933_n6960# 7.35e-19
C2035 a_108602_n29181# VDD 0.034176f
C2036 a_32353_n3548# I1U 0.002649f
C2037 a_33787_n8033# a_33787_n8930# 0.005987f
C2038 a_60285_n8035# a_60285_n8932# 0.005987f
C2039 a_67422_11614# VDD 0.046892f
C2040 a_57417_n8932# a_57977_n8932# 0.0284f
C2041 a_45445_n18698# a_44885_n18698# 0.0284f
C2042 a_45797_n18698# a_44363_n19595# 1.57e-19
C2043 a_81205_n9675# a_81735_n8770# 0.012586f
C2044 a_89407_n18620# VDD 0.112244f
C2045 a_110225_n1530# a_110225_n2435# 0.024773f
C2046 a_109695_n5150# a_111063_n2435# 0.002134f
C2047 a_55635_n33224# VDD 0.021515f
C2048 a_87433_n15905# IN_POS 0.00603f
C2049 a_101641_n18620# a_100235_n18620# 7.35e-19
C2050 a_46274_23609# a_44608_22884# 3.84e-20
C2051 a_40613_n3548# a_40965_n6239# 0.070243f
C2052 a_90969_11614# VDD 0.009062f
C2053 a_90969_n36322# VCM 0.001459f
C2054 a_67111_n4447# a_66551_n4447# 0.0284f
C2055 a_65677_n3550# a_66551_n5344# 0.030444f
C2056 a_53497_n14215# a_54019_n13318# 0.0284f
C2057 a_88271_n2435# a_88271_n3340# 0.005903f
C2058 a_111063_n6960# a_111631_n6960# 0.027101f
C2059 a_95943_n20430# VDD 0.399226f
C2060 a_109695_n7865# a_110225_n7865# 0.028522f
C2061 a_103997_n16810# a_105365_n14095# 0.002134f
C2062 a_83683_n36322# VDD 0.073724f
C2063 a_104527_n13190# a_104527_n14095# 0.024773f
C2064 a_40613_n8930# a_42047_n8930# 0.014106f
C2065 a_64243_n8932# a_65117_n8932# 0.001405f
C2066 a_54579_n17803# a_54579_n19597# 0.005987f
C2067 a_51711_n18700# a_53145_n19597# 1.57e-19
C2068 a_52063_n18700# a_52585_n18700# 0.0284f
C2069 a_87433_n1530# VDD 0.150485f
C2070 a_88839_n7865# a_88839_n8770# 0.005903f
C2071 a_100235_n20430# VDD 0.016652f
C2072 a_81205_n16810# a_81735_n15905# 0.012586f
C2073 a_104527_n18620# a_105365_n18620# 0.027101f
C2074 a_107339_n18620# a_107339_n20430# 0.012104f
C2075 a_103997_n21335# a_104527_n19525# 0.012586f
C2076 a_107230_13546# OUT 0.02829f
C2077 a_47753_n3548# a_48313_n4445# 0.0284f
C2078 a_32913_n14213# a_32913_n16904# 0.008933f
C2079 a_34699_n14213# a_35221_n14213# 0.0284f
C2080 a_35221_n13316# a_34347_n14213# 8.45e-19
C2081 a_58851_n13318# a_58851_n14215# 0.005987f
C2082 a_58329_n14215# a_59411_n14215# 0.00117f
C2083 a_93969_n3340# a_93969_n4245# 0.005903f
C2084 a_95943_n3340# a_95943_n6960# 0.012104f
C2085 a_93131_n2435# VDD 0.121415f
C2086 a_105365_n21335# VDD 0.02546f
C2087 a_83141_n19525# a_83709_n19525# 0.027101f
C2088 a_81735_n19525# a_81735_n20430# 0.024773f
C2089 a_109695_n16810# a_111063_n15000# 0.002134f
C2090 a_112199_n13190# a_112199_n14095# 0.024773f
C2091 a_60109_13546# a_60109_12380# 0.004007f
C2092 a_46879_n8930# a_48313_n8930# 0.014106f
C2093 a_33265_n18698# a_34347_n19595# 5.37e-19
C2094 a_33787_n17801# a_33787_n18698# 0.005987f
C2095 a_59763_n18700# a_58851_n18700# 5.43e-19
C2096 a_93131_n9675# a_93969_n9675# 0.027101f
C2097 a_98829_n3340# VDD 0.121044f
C2098 a_65117_n17803# IBNOUT -7.22e-35
C2099 a_32128_7563# I1U 5.57e-19
C2100 a_109695_n21335# a_110225_n20430# 0.012586f
C2101 a_54019_n3550# a_54579_n4447# 0.0284f
C2102 a_66029_n14215# a_65677_n14215# 0.062551f
C2103 a_63161_n15112# a_63683_n14215# 0.0284f
C2104 a_106501_n3340# VDD 0.121044f
C2105 a_55601_n28415# VDD 0.042519f
C2106 a_88839_n20430# a_89407_n20430# 0.027101f
C2107 a_83683_12380# a_83683_11614# 0.00778f
C2108 a_52585_n8035# a_52585_n8932# 0.005987f
C2109 a_53145_n8932# a_51711_n8932# 0.054819f
C2110 a_40965_n18698# a_41487_n17801# 0.0284f
C2111 a_64243_n18700# a_64243_n19597# 0.006457f
C2112 a_66029_n18700# a_66551_n18700# 0.0284f
C2113 a_111631_n4245# VDD 0.023105f
C2114 a_32128_n27257# I1U 5.57e-19
C2115 a_34347_n3548# a_35221_n4445# 0.005903f
C2116 a_59411_n3550# a_59763_n6241# 0.534125f
C2117 a_93969_n15905# IBPOUT 0.003499f
C2118 a_45445_n14213# a_46879_n14213# 9.78e-20
C2119 a_45797_n14213# a_46319_n14213# 0.0284f
C2120 a_48313_n13316# a_48313_n15110# 0.005987f
C2121 a_82573_n1530# a_82573_n2435# 0.005903f
C2122 a_104527_n6055# a_104527_n6960# 0.006141f
C2123 a_84547_n17715# VDD 0.472471f
C2124 a_107198_n29181# VDD 0.029136f
C2125 a_31831_n4445# I1U 0.008518f
C2126 a_84547_n15000# IN_POS 0.004986f
C2127 a_108636_12380# a_108636_11614# 0.00778f
C2128 a_35221_n8033# a_35781_n8930# 0.0284f
C2129 a_66016_11614# VDD 0.062166f
C2130 a_60845_n8932# a_57977_n8932# 5.37e-19
C2131 a_59411_n8932# a_60285_n8932# 5.43e-19
C2132 a_45445_n18698# a_44363_n19595# 5.37e-19
C2133 a_46319_n17801# a_47231_n18698# 5.43e-19
C2134 a_44885_n17801# a_44885_n18698# 0.005987f
C2135 a_82573_n6960# a_82573_n7865# 0.005903f
C2136 a_111063_n1530# a_111631_n1530# 0.027101f
C2137 a_88839_n18620# VDD 0.023105f
C2138 a_109695_n5150# a_110225_n2435# 0.012586f
C2139 a_54229_n33224# VDD 0.021515f
C2140 a_98829_n17715# a_98829_n18620# 0.006141f
C2141 a_45138_24195# a_45138_23609# 0.008552f
C2142 a_89563_n36322# VCM 6.2e-19
C2143 a_89563_11614# VDD 0.009062f
C2144 a_66551_n3550# a_66551_n4447# 0.005987f
C2145 a_63683_n4447# a_64243_n6241# 0.035468f
C2146 a_67111_n4447# a_66029_n6241# 0.002917f
C2147 a_51711_n14215# a_51151_n14215# 0.0284f
C2148 a_85089_11614# IN_POS 0.003316f
C2149 a_52063_n14215# a_50629_n15112# 1.57e-19
C2150 a_89407_n2435# a_90245_n3340# 0.028522f
C2151 a_113037_n6960# a_113037_n8770# 0.012104f
C2152 a_109695_n9675# a_111063_n7865# 0.002134f
C2153 a_95105_n19525# VDD 0.121371f
C2154 a_85089_n35156# VDD 0.061113f
C2155 a_103997_n16810# a_104527_n14095# 0.012586f
C2156 a_105365_n13190# a_105933_n13190# 0.027101f
C2157 a_49795_6405# a_49795_5639# 0.00778f
C2158 a_40613_n8930# a_41487_n8033# 5.43e-19
C2159 a_38619_n8033# a_38619_n8930# 0.005987f
C2160 a_67111_n8932# a_66551_n8932# 0.0284f
C2161 a_114516_10448# VDD 0.02294f
C2162 a_71896_n33224# OUT 0.003436f
C2163 a_53497_n18700# a_54019_n17803# 0.0284f
C2164 a_86903_n5150# VDD 0.916148f
C2165 a_99667_n20430# VDD 0.016652f
C2166 a_82573_n14095# a_83141_n14095# 0.027101f
C2167 a_103997_n19525# a_105365_n18620# 2.31e-19
C2168 a_46879_n3548# a_48313_n4445# 0.08885f
C2169 a_34699_n14213# a_34347_n14213# 0.16936f
C2170 a_31831_n15110# a_32353_n14213# 0.0284f
C2171 a_58329_n14215# a_58851_n14215# 0.0284f
C2172 a_60845_n13318# a_60845_n15112# 0.005987f
C2173 a_57977_n14215# a_59411_n14215# 5.12e-19
C2174 a_94537_n3340# a_95105_n3340# 0.027101f
C2175 a_81205_n21335# a_82573_n21335# 0.002563f
C2176 a_104527_n21335# VDD 0.150485f
C2177 a_110225_n14095# a_111063_n14095# 0.027101f
C2178 a_109695_n16810# a_110225_n15000# 0.012586f
C2179 a_113081_n28415# a_113081_n29181# 0.00778f
C2180 a_44885_n8033# a_44885_n8930# 0.005987f
C2181 a_46879_n8930# a_47753_n8033# 5.43e-19
C2182 a_35781_n17801# a_35781_n19595# 0.005987f
C2183 a_33265_n18698# a_33787_n18698# 0.0284f
C2184 a_32913_n18698# a_34347_n19595# 1.57e-19
C2185 a_90935_5639# VDD 0.042519f
C2186 a_58851_n17803# a_58851_n18700# 0.005987f
C2187 a_85129_7563# IN_POS 6.24e-19
C2188 a_58329_n18700# a_59411_n19597# 5.37e-19
C2189 a_98299_n4245# VDD 0.399575f
C2190 a_94537_n8770# a_94537_n9675# 0.005903f
C2191 a_112199_n21335# VDD 0.150485f
C2192 a_90245_n15000# a_89407_n15000# 0.028522f
C2193 a_64595_n18700# IBNOUT 0.011856f
C2194 a_87433_n15000# a_88271_n15000# 0.027101f
C2195 a_111063_n18620# a_111063_n19525# 0.005903f
C2196 a_53145_n3550# a_54579_n4447# 0.003256f
C2197 a_39531_n14213# a_40613_n14213# 0.011365f
C2198 a_40053_n13316# a_40053_n14213# 0.005987f
C2199 a_66029_n14215# a_65117_n14215# 5.43e-19
C2200 a_105933_n3340# VDD 0.016281f
C2201 a_54197_n28415# VDD 0.042519f
C2202 a_87433_n20430# a_87433_n21335# 0.024773f
C2203 a_32353_n13316# I1U 0.002649f
C2204 a_114485_6405# a_114485_5639# 0.00778f
C2205 a_54019_n8035# a_54579_n8932# 0.0284f
C2206 a_39531_n18698# a_38097_n19595# 1.57e-19
C2207 a_39179_n18698# a_38619_n18698# 0.0284f
C2208 a_63161_n19597# a_63683_n18700# 0.0284f
C2209 a_66029_n18700# a_65677_n19597# 0.053799f
C2210 a_111063_n4245# VDD 0.012916f
C2211 a_93969_n15905# a_94537_n15905# 0.027101f
C2212 a_30724_n27257# I1U 0.004931f
C2213 a_34347_n3548# a_34699_n6239# 0.070243f
C2214 a_59411_n3550# a_57977_n6241# 4.66e-19
C2215 a_43848_13546# VDD 0.026416f
C2216 a_93131_n15905# IBPOUT 0.01873f
C2217 a_47231_n14213# a_47753_n13316# 0.0284f
C2218 a_81735_n17715# VDD 0.41764f
C2219 a_108602_n28415# VDD 0.042519f
C2220 a_61484_n27257# a_61484_n28415# 0.004047f
C2221 a_34347_n8930# a_35781_n8930# 0.014106f
C2222 a_67422_12380# VDD 0.061113f
C2223 a_59411_n8932# a_58851_n8932# 0.0284f
C2224 a_45797_n18698# a_47231_n18698# 0.014106f
C2225 a_83141_n6960# a_83709_n6960# 0.027101f
C2226 a_88271_n18620# VDD 0.012916f
C2227 a_49755_n36322# VDD 0.05845f
C2228 a_73268_n28415# a_73268_n29181# 0.00778f
C2229 a_45706_24195# a_46274_23609# 0.018349f
C2230 a_41487_n3548# a_42047_n4445# 0.0284f
C2231 a_65677_n3550# a_66551_n4447# 4.96e-19
C2232 a_90969_12380# VDD 0.009062f
C2233 a_51151_n13318# a_51151_n14215# 0.005987f
C2234 a_51711_n14215# a_50629_n15112# 5.37e-19
C2235 a_52585_n13318# a_53497_n14215# 5.43e-19
C2236 a_88839_n2435# a_90245_n3340# 2.31e-19
C2237 a_87433_n2435# a_87433_n3340# 0.024773f
C2238 a_94537_n19525# VDD 0.016281f
C2239 a_110225_n6960# a_111063_n6960# 0.027101f
C2240 a_109695_n9675# a_110225_n7865# 0.012586f
C2241 a_83683_n35156# VDD 0.076387f
C2242 a_38097_n8930# a_38619_n8930# 0.0284f
C2243 a_113110_10448# VDD 0.029536f
C2244 a_66551_n8035# a_66551_n8932# 0.005987f
C2245 a_63683_n8932# a_64243_n8932# 0.0284f
C2246 a_51711_n18700# a_51151_n18700# 0.0284f
C2247 a_52063_n18700# a_50629_n19597# 1.57e-19
C2248 a_89407_n7865# a_90245_n8770# 0.028522f
C2249 a_88271_n7865# a_88271_n8770# 0.005903f
C2250 a_83709_n9675# VDD 0.177586f
C2251 a_98829_n20430# VDD 0.121415f
C2252 a_103997_n19525# a_104527_n18620# 0.028522f
C2253 a_44363_n4445# a_45445_n6239# 0.002568f
C2254 a_44885_n3548# a_44885_n4445# 0.005987f
C2255 a_46879_n3548# a_47753_n3548# 0.006769f
C2256 a_59763_n14215# a_60285_n13318# 0.0284f
C2257 a_95105_n1530# VDD 0.150485f
C2258 a_92601_n4245# a_93969_n4245# 2.31e-19
C2259 a_93131_n3340# a_93131_n4245# 0.024773f
C2260 a_106501_n20430# VDD 0.121415f
C2261 a_82573_n19525# a_83141_n19525# 0.027101f
C2262 a_81205_n21335# a_81735_n21335# 0.044257f
C2263 a_87433_n8770# IN_POS 0.00603f
C2264 a_111631_n13190# a_111631_n14095# 0.005903f
C2265 a_109695_n16810# a_109695_n15905# 0.086469f
C2266 a_44363_n8930# a_44885_n8930# 0.0284f
C2267 a_89531_5639# VDD 0.042519f
C2268 a_34699_n18698# a_35221_n17801# 0.0284f
C2269 a_60845_n17803# a_60845_n19597# 0.005987f
C2270 a_57977_n18700# a_59411_n19597# 1.57e-19
C2271 a_58329_n18700# a_58851_n18700# 0.0284f
C2272 a_101641_n3340# VDD 0.399226f
C2273 a_111631_n21335# VDD 0.02546f
C2274 a_86903_n15905# a_88271_n15000# 2.31e-19
C2275 a_90245_n15000# a_88839_n15000# 2.31e-19
C2276 a_89407_n14095# a_89407_n15000# 0.024773f
C2277 a_64243_n18700# IBNOUT 0.029699f
C2278 a_30724_7563# I1U 0.004931f
C2279 a_111631_n18620# a_112199_n18620# 0.027101f
C2280 a_42442_n33224# a_42442_n34390# 0.004007f
C2281 a_96818_5639# a_96818_4481# 0.004047f
C2282 a_53145_n3550# a_54019_n3550# 0.004425f
C2283 a_51151_n3550# a_51151_n4447# 0.005987f
C2284 a_50629_n4447# a_51711_n6241# 0.001037f
C2285 a_39531_n14213# a_40053_n14213# 0.0284f
C2286 a_42047_n13316# a_42047_n15110# 0.005987f
C2287 a_39179_n14213# a_40613_n14213# 9.78e-20
C2288 a_64595_n14215# a_65677_n14215# 0.00117f
C2289 a_65117_n13318# a_65117_n14215# 0.005987f
C2290 a_105365_n3340# VDD 0.016281f
C2291 a_88271_n20430# a_88839_n20430# 0.027101f
C2292 a_30724_n29181# a_30724_n30339# 0.004047f
C2293 a_85089_13546# a_85089_12380# 0.004007f
C2294 a_53145_n8932# a_54579_n8932# 0.014106f
C2295 a_40053_n17801# a_40965_n18698# 5.43e-19
C2296 a_38619_n17801# a_38619_n18698# 0.005987f
C2297 a_39179_n18698# a_38097_n19595# 5.37e-19
C2298 w_27790_n38888# IN_POS 0.024701f
C2299 a_66029_n18700# a_65117_n18700# 5.43e-19
C2300 a_110225_n4245# VDD 0.137705f
C2301 a_100235_n9675# a_100803_n9675# 0.027101f
C2302 a_95105_n15000# a_95105_n15905# 0.024773f
C2303 a_60285_n3550# a_60845_n4447# 0.0284f
C2304 a_48313_n13316# a_46879_n14213# 0.018216f
C2305 a_45797_n14213# a_44363_n15110# 1.57e-19
C2306 a_45445_n14213# a_44885_n14213# 0.0284f
C2307 a_83141_n1530# a_83709_n1530# 0.027101f
C2308 a_81205_n5150# a_82573_n2435# 0.002134f
C2309 a_81735_n1530# a_81735_n2435# 0.024773f
C2310 a_84547_n18620# VDD 1.18674f
C2311 a_107198_n28415# VDD 0.042519f
C2312 a_94537_n21335# a_95105_n21335# 0.027101f
C2313 a_107230_12380# a_107230_11614# 0.00778f
C2314 a_32353_n8033# a_32353_n8930# 0.005987f
C2315 a_34347_n8930# a_35221_n8033# 5.43e-19
C2316 a_59411_n8932# a_57977_n8932# 0.054819f
C2317 a_58851_n8035# a_58851_n8932# 0.005987f
C2318 a_66016_12380# VDD 0.076387f
C2319 a_45797_n18698# a_46319_n17801# 0.0284f
C2320 a_81735_n6960# a_81735_n7865# 0.024773f
C2321 a_81205_n7865# a_82573_n7865# 2.31e-19
C2322 a_110225_n1530# a_111063_n1530# 0.027101f
C2323 a_87433_n18620# VDD 0.137705f
C2324 a_48349_n36322# VDD 0.073724f
C2325 a_45138_24195# a_46274_23609# 1.92e-19
C2326 a_108636_n34390# a_108636_n35156# 0.00778f
C2327 a_40613_n3548# a_42047_n4445# 0.08885f
C2328 a_89563_12380# VDD 0.009062f
C2329 a_65677_n3550# a_66029_n6241# 0.534125f
C2330 a_53145_n13318# a_53145_n14215# 0.011408f
C2331 a_52063_n14215# a_53497_n14215# 0.014106f
C2332 a_85089_12380# IN_POS 0.003316f
C2333 a_86903_n5150# a_88271_n4245# 0.002134f
C2334 a_88839_n2435# a_89407_n2435# 0.027101f
C2335 a_109695_n7865# a_111063_n6960# 2.31e-19
C2336 a_93969_n19525# VDD 0.016281f
C2337 a_85089_n34390# VDD 0.046892f
C2338 a_104527_n13190# a_105365_n13190# 0.027101f
C2339 a_48391_6405# a_48391_5639# 0.00778f
C2340 a_40053_n8033# a_40613_n8930# 0.0284f
C2341 a_65677_n8932# a_66551_n8932# 5.43e-19
C2342 a_67111_n8932# a_64243_n8932# 5.37e-19
C2343 a_114516_11614# VDD 0.013383f
C2344 a_51151_n17803# a_51151_n18700# 0.005987f
C2345 a_51711_n18700# a_50629_n19597# 5.37e-19
C2346 a_88839_n7865# a_90245_n8770# 2.31e-19
C2347 a_83141_n9675# VDD 0.02546f
C2348 a_83709_n13190# a_83709_n14095# 0.024773f
C2349 a_81735_n14095# a_82573_n14095# 0.027101f
C2350 a_81205_n16810# a_82573_n15000# 0.002134f
C2351 a_103997_n21335# a_105365_n18620# 0.002134f
C2352 a_66058_7563# a_66058_6405# 0.004047f
C2353 a_44363_n4445# a_44885_n4445# 0.0284f
C2354 a_47231_n3548# a_47231_n6239# 0.0089f
C2355 a_33265_n14213# a_34347_n14213# 0.011365f
C2356 a_33787_n13316# a_33787_n14213# 0.005987f
C2357 a_57977_n14215# a_57417_n14215# 0.0284f
C2358 a_58329_n14215# a_56895_n15112# 1.57e-19
C2359 a_93969_n3340# a_94537_n3340# 0.027101f
C2360 a_94537_n1530# VDD 0.02546f
C2361 a_92601_n4245# a_93131_n4245# 0.028522f
C2362 a_83709_n18620# a_83709_n19525# 0.024773f
C2363 a_105933_n20430# VDD 0.016652f
C2364 a_46319_n8033# a_46879_n8930# 0.0284f
C2365 a_90935_6405# VDD 0.034176f
C2366 a_33265_n18698# a_31831_n19595# 1.57e-19
C2367 a_32913_n18698# a_32353_n18698# 0.0284f
C2368 a_59763_n18700# a_60285_n17803# 0.0284f
C2369 a_100803_n2435# VDD 0.121415f
C2370 a_93969_n8770# a_93969_n9675# 0.005903f
C2371 a_86903_n16810# a_86903_n21335# 0.032645f
C2372 a_63683_n17803# IBNOUT 0.004735f
C2373 a_86903_n15905# a_87433_n15000# 0.028522f
C2374 a_111063_n21335# VDD 0.02546f
C2375 a_110225_n18620# a_110225_n19525# 0.024773f
C2376 a_109695_n19525# a_111063_n19525# 2.31e-19
C2377 a_53497_n3550# a_53497_n6241# 0.009483f
C2378 a_50629_n4447# a_51151_n4447# 0.0284f
C2379 a_40965_n14213# a_41487_n13316# 0.0284f
C2380 a_64243_n14215# a_65677_n14215# 5.12e-19
C2381 a_64595_n14215# a_65117_n14215# 0.0284f
C2382 a_67111_n13318# a_67111_n15112# 0.005987f
C2383 a_104527_n3340# VDD 0.121044f
C2384 a_100803_n4245# a_101641_n6960# 0.042385f
C2385 a_90245_n20430# a_89407_n20430# 0.028522f
C2386 a_113081_6405# a_113081_5639# 0.00778f
C2387 a_53145_n8932# a_54019_n8035# 5.43e-19
C2388 a_50629_n8932# a_51711_n8932# 5.37e-19
C2389 a_51151_n8035# a_51151_n8932# 0.005987f
C2390 a_39531_n18698# a_40965_n18698# 0.014106f
C2391 a_75585_n10973# I1N 0.134577f
C2392 a_65117_n17803# a_65117_n18700# 0.005987f
C2393 a_64595_n18700# a_65677_n19597# 5.37e-19
C2394 a_112199_n3340# VDD 0.121371f
C2395 a_93131_n15905# a_93969_n15905# 0.027101f
C2396 a_35221_n3548# a_35781_n4445# 0.0284f
C2397 a_59411_n3550# a_60845_n4447# 0.003256f
C2398 a_42442_13546# VDD 0.029536f
C2399 a_45445_n14213# a_44363_n15110# 5.37e-19
C2400 a_46319_n13316# a_47231_n14213# 5.43e-19
C2401 a_44885_n13316# a_44885_n14213# 0.005987f
C2402 a_94537_n15000# IBPOUT 0.00243f
C2403 a_81205_n5150# a_81735_n2435# 0.012586f
C2404 a_104527_n6055# a_103997_n9675# 0.035071f
C2405 a_83709_n15905# VDD 0.138244f
C2406 a_60080_n27257# a_60080_n28415# 0.004047f
C2407 a_90969_n34390# a_90969_n35156# 0.00778f
C2408 a_31831_n8930# a_32353_n8930# 0.0284f
C2409 a_67422_13546# VDD 0.05845f
C2410 a_60285_n8035# a_60845_n8932# 0.0284f
C2411 a_48313_n17801# a_47753_n17801# 0.0284f
C2412 a_84547_n6960# a_84547_n8770# 0.011861f
C2413 a_81205_n7865# a_81735_n7865# 0.028522f
C2414 a_82573_n6960# a_83141_n6960# 0.027101f
C2415 a_81205_n9675# a_82573_n7865# 0.002134f
C2416 a_109695_n5150# a_111063_n1530# 0.002563f
C2417 a_86903_n19525# VDD 0.399575f
C2418 a_98829_n17715# a_98299_n21335# 0.035071f
C2419 a_31699_17542# I1U 0.269982f
C2420 a_49755_n35156# VDD 0.061113f
C2421 a_87433_n15000# IN_POS 0.00603f
C2422 a_71864_n28415# a_71864_n29181# 0.00778f
C2423 a_45138_24195# a_45706_24195# 0.017228f
C2424 a_46274_24920# a_46274_23609# 0.007268f
C2425 a_30724_5639# a_30724_4481# 0.004047f
C2426 a_40613_n3548# a_41487_n3548# 0.006769f
C2427 a_38619_n3548# a_38619_n4445# 0.005987f
C2428 a_38097_n4445# a_39179_n6239# 0.002568f
C2429 a_65677_n3550# a_64243_n6241# 4.66e-19
C2430 a_52063_n14215# a_52585_n13318# 0.0284f
C2431 a_86903_n5150# a_87433_n4245# 0.012586f
C2432 a_93131_n19525# VDD 0.121044f
C2433 a_109695_n7865# a_110225_n6960# 0.028522f
C2434 a_83683_n34390# VDD 0.062166f
C2435 a_103997_n16810# a_105365_n13190# 0.002563f
C2436 a_113110_11614# VDD 0.017204f
C2437 a_65677_n8932# a_65117_n8932# 0.0284f
C2438 a_53145_n17803# a_54579_n19597# 0.018216f
C2439 a_52063_n18700# a_53497_n18700# 0.005986f
C2440 a_82573_n9675# VDD 0.02546f
C2441 a_88839_n7865# a_89407_n7865# 0.027101f
C2442 a_87433_n7865# a_87433_n8770# 0.024773f
C2443 a_81205_n16810# a_81735_n15000# 0.012586f
C2444 a_101641_n20430# VDD 0.392932f
C2445 a_103997_n21335# a_104527_n18620# 0.012586f
C2446 a_46319_n3548# a_46879_n3548# 0.0284f
C2447 a_32913_n14213# a_34347_n14213# 9.78e-20
C2448 a_33265_n14213# a_33787_n14213# 0.0284f
C2449 a_35781_n13316# a_35781_n15110# 0.005987f
C2450 a_57977_n14215# a_56895_n15112# 5.37e-19
C2451 a_58851_n13318# a_59763_n14215# 5.43e-19
C2452 a_57417_n13318# a_57417_n14215# 0.005987f
C2453 a_93969_n1530# VDD 0.02546f
C2454 a_81735_n19525# a_82573_n19525# 0.027101f
C2455 a_105365_n20430# VDD 0.016652f
C2456 a_111063_n13190# a_111063_n14095# 0.005903f
C2457 a_114485_n27257# a_114485_n28415# 0.004047f
C2458 a_33787_n17801# a_34699_n18698# 5.43e-19
C2459 a_32353_n17801# a_32353_n18698# 0.005987f
C2460 a_89531_6405# VDD 0.029136f
C2461 a_32913_n18698# a_31831_n19595# 5.37e-19
C2462 a_58329_n18700# a_56895_n19597# 1.57e-19
C2463 a_57977_n18700# a_57417_n18700# 0.0284f
C2464 a_94537_n8770# a_95105_n8770# 0.027101f
C2465 a_100235_n2435# VDD 0.016652f
C2466 a_88839_n14095# a_88839_n15000# 0.005903f
C2467 a_110225_n21335# VDD 0.150485f
C2468 a_109695_n19525# a_110225_n19525# 0.028522f
C2469 a_111063_n18620# a_111631_n18620# 0.027101f
C2470 a_71864_4481# OUT 0.001942f
C2471 a_95414_5639# a_95414_4481# 0.004047f
C2472 a_52585_n3550# a_53145_n3550# 0.037577f
C2473 a_39179_n14213# a_38619_n14213# 0.0284f
C2474 a_39531_n14213# a_38097_n15110# 1.57e-19
C2475 a_42047_n13316# a_40613_n14213# 0.018216f
C2476 a_66029_n14215# a_66551_n13318# 0.0284f
C2477 a_103997_n4245# VDD 0.399575f
C2478 a_100235_n4245# a_101641_n6960# 0.002302f
C2479 a_87433_n20430# a_88271_n20430# 0.027101f
C2480 a_89407_n19525# a_89407_n20430# 0.024773f
C2481 a_90245_n20430# a_88839_n20430# 2.31e-19
C2482 a_32128_n28415# a_32128_n29181# 0.00778f
C2483 a_83683_13546# a_83683_12380# 0.004007f
C2484 a_50629_n8932# a_51151_n8932# 0.0284f
C2485 a_39531_n18698# a_40053_n17801# 0.0284f
C2486 a_72603_n10973# I1N 0.14436f
C2487 a_64243_n18700# a_65677_n19597# 1.57e-19
C2488 a_67111_n17803# a_67111_n19597# 0.005987f
C2489 a_64595_n18700# a_65117_n18700# 0.0284f
C2490 a_111631_n3340# VDD 0.016281f
C2491 a_99667_n9675# a_100235_n9675# 0.027101f
C2492 a_94537_n15000# a_94537_n15905# 0.005903f
C2493 a_34347_n3548# a_35781_n4445# 0.08885f
C2494 a_56895_n4447# a_57977_n6241# 0.001037f
C2495 a_59411_n3550# a_60285_n3550# 0.004425f
C2496 a_57417_n3550# a_57417_n4447# 0.005987f
C2497 a_93969_n15000# IBPOUT 0.003499f
C2498 a_45797_n14213# a_47231_n14213# 0.005986f
C2499 a_46879_n13316# a_46879_n14213# 0.01664f
C2500 a_82573_n1530# a_83141_n1530# 0.027101f
C2501 a_83141_n15905# VDD 0.01295f
C2502 a_93969_n21335# a_94537_n21335# 0.027101f
C2503 a_33787_n8033# a_34347_n8930# 0.0284f
C2504 a_59411_n8932# a_60845_n8932# 0.014106f
C2505 a_66016_13546# VDD 0.073724f
C2506 a_45445_n18698# a_45797_n18698# 0.210644f
C2507 a_46879_n17801# a_46879_n19595# 0.011408f
C2508 a_47753_n16904# a_47753_n17801# 0.005987f
C2509 a_48313_n17801# a_47231_n18698# 5.37e-19
C2510 a_81205_n9675# a_81735_n7865# 0.012586f
C2511 a_86903_n21335# VDD 1.40049f
C2512 a_109695_n5150# a_110225_n1530# 0.044257f
C2513 a_30377_18342# I1U 0.258844f
C2514 a_48349_n35156# VDD 0.076387f
C2515 a_86903_n15905# IN_POS 0.001743f
C2516 a_107230_n34390# a_107230_n35156# 0.00778f
C2517 a_40965_n3548# a_40965_n6239# 0.0089f
C2518 a_38097_n4445# a_38619_n4445# 0.0284f
C2519 a_90969_13546# VDD 0.021314f
C2520 a_66551_n3550# a_67111_n4447# 0.0284f
C2521 a_54579_n13318# a_54019_n13318# 0.0284f
C2522 a_85089_13546# IN_POS 0.003316f
C2523 a_88271_n2435# a_88839_n2435# 0.027101f
C2524 a_109695_n9675# a_111063_n6960# 0.002134f
C2525 a_95105_n18620# VDD 0.128099f
C2526 a_103997_n16810# a_104527_n13190# 0.044257f
C2527 a_85089_n33224# VDD 0.05812f
C2528 a_83725_n29181# a_83725_n30339# 0.004047f
C2529 a_66058_n30339# IBNOUT 6.21e-20
C2530 a_41487_n7136# a_41487_n8033# 0.005987f
C2531 a_40965_n8033# a_42047_n8930# 5.37e-19
C2532 a_65677_n8932# a_64243_n8932# 0.054819f
C2533 a_65117_n8035# a_65117_n8932# 0.005987f
C2534 a_114516_12380# VDD 0.010487f
C2535 a_53145_n17803# a_54019_n18700# 8.45e-19
C2536 a_52063_n18700# a_52585_n17803# 0.0284f
C2537 a_81735_n9675# VDD 0.150485f
C2538 a_86903_n9675# a_88271_n9675# 0.002563f
C2539 a_83141_n13190# a_83141_n14095# 0.005903f
C2540 a_81205_n16810# a_81205_n15905# 0.086339f
C2541 a_100803_n19525# VDD 0.121044f
C2542 a_103997_n21335# a_103997_n19525# 0.086339f
C2543 a_107339_n18620# a_106501_n18620# 0.032618f
C2544 a_114516_n36322# VDD 0.02603f
C2545 a_34699_n14213# a_35221_n13316# 0.0284f
C2546 a_58329_n14215# a_59763_n14215# 0.014106f
C2547 a_59411_n13318# a_59411_n14215# 0.011408f
C2548 a_93131_n1530# VDD 0.150485f
C2549 a_93131_n3340# a_93969_n3340# 0.027101f
C2550 a_95943_n3340# a_95105_n3340# 0.028522f
C2551 a_104527_n20430# VDD 0.121415f
C2552 a_81205_n21335# a_82573_n20430# 0.002134f
C2553 a_83141_n18620# a_83141_n19525# 0.005903f
C2554 a_111631_n13190# a_112199_n13190# 0.027101f
C2555 a_47753_n7136# a_47753_n8033# 0.005987f
C2556 a_47231_n8033# a_48313_n8930# 5.37e-19
C2557 a_33265_n18698# a_34699_n18698# 0.014106f
C2558 a_90935_7563# VDD 0.00658f
C2559 a_57977_n18700# a_56895_n19597# 5.37e-19
C2560 a_57417_n17803# a_57417_n18700# 0.005987f
C2561 a_99667_n2435# VDD 0.016652f
C2562 a_93131_n8770# a_93131_n9675# 0.024773f
C2563 a_86903_n16810# a_87433_n17715# 0.035071f
C2564 a_112199_n20430# VDD 0.121415f
C2565 a_109695_n21335# a_111063_n19525# 0.002134f
C2566 a_39179_n14213# a_38097_n15110# 5.37e-19
C2567 a_40053_n13316# a_40965_n14213# 5.43e-19
C2568 a_38619_n13316# a_38619_n14213# 0.005987f
C2569 a_64595_n14215# a_63161_n15112# 1.57e-19
C2570 a_64243_n14215# a_63683_n14215# 0.0284f
C2571 a_100235_n4245# a_100803_n4245# 0.027101f
C2572 a_107339_n3340# VDD 0.399226f
C2573 a_98829_n4245# a_98829_n6055# 0.006141f
C2574 a_114485_7563# a_114485_6405# 0.004047f
C2575 a_53497_n8035# a_51711_n8932# 0.006457f
C2576 a_52585_n8035# a_53145_n8932# 0.0284f
C2577 a_42047_n17801# a_41487_n17801# 0.0284f
C2578 a_66029_n18700# a_66551_n17803# 0.0284f
C2579 a_75585_n10073# I1N 0.159921f
C2580 a_111063_n3340# VDD 0.016281f
C2581 a_100803_n8770# a_100803_n9675# 0.024773f
C2582 a_95443_13546# a_95443_12380# 0.004007f
C2583 a_31831_n4445# a_32913_n6239# 0.002568f
C2584 a_32353_n3548# a_32353_n4445# 0.005987f
C2585 a_34347_n3548# a_35221_n3548# 0.006769f
C2586 a_37968_10448# VDD 0.021515f
C2587 a_59763_n3550# a_59763_n6241# 0.009483f
C2588 a_56895_n4447# a_57417_n4447# 0.0284f
C2589 a_45797_n14213# a_46319_n13316# 0.0284f
C2590 a_93131_n15000# IBPOUT 0.019592f
C2591 a_107339_n6960# a_107339_n6055# 0.088786f
C2592 a_82573_n15905# VDD 0.023101f
C2593 a_95105_n20430# a_95105_n21335# 0.024773f
C2594 a_89563_n34390# a_89563_n35156# 0.00778f
C2595 a_59411_n8932# a_60285_n8035# 5.43e-19
C2596 a_56895_n8932# a_57977_n8932# 5.37e-19
C2597 a_57417_n8035# a_57417_n8932# 0.005987f
C2598 a_44363_n17801# a_44363_n19595# 0.005987f
C2599 a_81735_n6960# a_82573_n6960# 0.027101f
C2600 a_90245_n17715# VDD 0.472471f
C2601 a_31699_19142# I1U 0.260073f
C2602 a_101641_n18620# a_101641_n17715# 0.088786f
C2603 a_49755_n34390# VDD 0.046892f
C2604 a_44608_24195# a_44608_22884# 0.012404f
C2605 a_45706_24920# a_45706_24195# 0.006281f
C2606 a_32128_6405# a_32128_5639# 0.00778f
C2607 a_40053_n3548# a_40613_n3548# 0.0284f
C2608 a_65677_n3550# a_67111_n4447# 0.003256f
C2609 a_51711_n14215# a_52063_n14215# 0.210644f
C2610 a_54019_n12421# a_54019_n13318# 0.005987f
C2611 a_54579_n13318# a_53497_n14215# 5.37e-19
C2612 a_94537_n18620# VDD 0.023105f
C2613 a_113037_n6960# a_112199_n6960# 0.032618f
C2614 a_109695_n9675# a_110225_n6960# 0.012586f
C2615 a_83683_n33224# VDD 0.073394f
C2616 a_40965_n8033# a_41487_n8033# 0.0284f
C2617 a_66551_n8035# a_67111_n8932# 0.0284f
C2618 a_113110_12380# VDD 0.017204f
C2619 a_54579_n17803# a_54019_n17803# 0.0284f
C2620 a_53145_n17803# a_53145_n19597# 0.01664f
C2621 a_83709_n8770# VDD 0.121415f
C2622 a_88271_n7865# a_88839_n7865# 0.027101f
C2623 a_86903_n9675# a_87433_n9675# 0.044257f
C2624 a_100235_n19525# VDD 0.016281f
C2625 a_113110_n36322# VDD 0.029536f
C2626 a_107339_n18620# a_105933_n18620# 7.35e-19
C2627 a_47753_n2651# a_47753_n3548# 0.005987f
C2628 a_47231_n3548# a_48313_n4445# 5.37e-19
C2629 a_33265_n14213# a_31831_n15110# 1.57e-19
C2630 a_35781_n13316# a_34347_n14213# 0.018216f
C2631 a_32913_n14213# a_32353_n14213# 0.0284f
C2632 a_55601_5639# VDD 0.042519f
C2633 a_58329_n14215# a_58851_n13318# 0.0284f
C2634 a_75602_n4978# VDD 0.03531f
C2635 a_92601_n5150# VDD 1.28138f
C2636 a_92601_n4245# a_93969_n3340# 2.31e-19
C2637 a_95943_n3340# a_94537_n3340# 2.31e-19
C2638 a_95105_n2435# a_95105_n3340# 0.024773f
C2639 a_81205_n21335# a_81735_n20430# 0.012586f
C2640 a_110225_n13190# a_110225_n14095# 0.024773f
C2641 a_109695_n16810# a_111063_n14095# 0.002134f
C2642 a_113081_n27257# a_113081_n28415# 0.004047f
C2643 a_47231_n8033# a_47753_n8033# 0.0284f
C2644 a_33265_n18698# a_33787_n17801# 0.0284f
C2645 a_59411_n17803# a_60845_n19597# 0.018216f
C2646 a_58329_n18700# a_59763_n18700# 0.005986f
C2647 a_98829_n2435# VDD 0.149203f
C2648 a_93969_n8770# a_94537_n8770# 0.027101f
C2649 a_88271_n14095# a_88271_n15000# 0.005903f
C2650 a_63683_n16906# IBNOUT 0.004735f
C2651 a_111631_n20430# VDD 0.016652f
C2652 a_110225_n18620# a_111063_n18620# 0.027101f
C2653 a_113037_n18620# a_113037_n20430# 0.012104f
C2654 a_109695_n21335# a_110225_n19525# 0.012586f
C2655 a_66016_n36322# IBNOUT 5.91e-19
C2656 a_71864_5639# OUT 0.001942f
C2657 a_96818_6405# a_96818_5639# 0.00778f
C2658 a_54019_n2653# a_54019_n3550# 0.005987f
C2659 a_53497_n3550# a_54579_n4447# 5.37e-19
C2660 a_40613_n13316# a_40613_n14213# 0.01664f
C2661 a_39531_n14213# a_40965_n14213# 0.005986f
C2662 a_63683_n13318# a_63683_n14215# 0.005987f
C2663 a_65117_n13318# a_66029_n14215# 5.43e-19
C2664 a_64243_n14215# a_63161_n15112# 5.37e-19
C2665 a_106501_n2435# VDD 0.121415f
C2666 a_88839_n19525# a_88839_n20430# 0.005903f
C2667 a_30724_n28415# a_30724_n29181# 0.00778f
C2668 a_32913_n12419# I1U 2.01e-19
C2669 a_42047_n17801# a_40965_n18698# 5.37e-19
C2670 a_39179_n18698# a_39531_n18698# 0.210644f
C2671 a_41487_n16904# a_41487_n17801# 0.005987f
C2672 a_40613_n17801# a_40613_n19595# 0.011408f
C2673 a_64243_n18700# a_63683_n18700# 0.0284f
C2674 a_72603_n10073# I1N 0.158537f
C2675 a_64595_n18700# a_63161_n19597# 1.57e-19
C2676 a_110225_n3340# VDD 0.121044f
C2677 a_98829_n9675# a_99667_n9675# 0.027101f
C2678 a_93969_n15000# a_93969_n15905# 0.005903f
C2679 a_95943_n15000# a_95943_n18620# 0.012104f
C2680 a_73302_n34390# a_73302_n35156# 0.00778f
C2681 a_31831_n4445# a_32353_n4445# 0.0284f
C2682 a_34699_n3548# a_34699_n6239# 0.0089f
C2683 a_36562_10448# VDD 0.021515f
C2684 a_58851_n3550# a_59411_n3550# 0.037577f
C2685 a_92601_n15905# IBPOUT 0.015637f
C2686 a_48313_n13316# a_47753_n13316# 0.0284f
C2687 a_81735_n1530# a_82573_n1530# 0.027101f
C2688 a_81735_n15905# VDD 0.113729f
C2689 a_93131_n21335# a_93969_n21335# 0.027101f
C2690 a_32353_n2651# I1U 0.002649f
C2691 a_35221_n7136# a_35221_n8033# 0.005987f
C2692 a_34699_n8033# a_35781_n8930# 5.37e-19
C2693 a_56895_n8932# a_57417_n8932# 0.0284f
C2694 a_44885_n17801# a_45445_n18698# 0.0284f
C2695 a_81205_n7865# a_82573_n6960# 2.31e-19
C2696 a_30377_19942# I1U 0.258645f
C2697 a_87433_n17715# VDD 0.41764f
C2698 a_48349_n34390# VDD 0.062166f
C2699 a_44608_24195# a_46274_23609# 3.84e-20
C2700 a_63683_n3550# a_63683_n4447# 0.005987f
C2701 a_65677_n3550# a_66551_n3550# 0.004425f
C2702 a_63161_n4447# a_64243_n6241# 0.001037f
C2703 a_53145_n13318# a_54019_n13318# 5.43e-19
C2704 a_86903_n5150# a_88271_n3340# 0.002134f
C2705 a_89407_n1530# a_89407_n2435# 0.024773f
C2706 a_87433_n2435# a_88271_n2435# 0.027101f
C2707 a_109695_n9675# a_109695_n7865# 0.086339f
C2708 a_113037_n6960# a_111631_n6960# 7.35e-19
C2709 a_93969_n18620# VDD 0.012916f
C2710 a_79182_n36322# VDD 0.024605f
C2711 a_85129_n28415# a_85129_n29181# 0.00778f
C2712 a_66058_n29181# IBNOUT 6.21e-20
C2713 a_40965_n8033# a_40613_n8930# 0.053799f
C2714 a_38097_n8930# a_38619_n8033# 0.0284f
C2715 a_65677_n8932# a_67111_n8932# 0.014106f
C2716 a_54019_n16906# a_54019_n17803# 0.005987f
C2717 a_51711_n18700# a_52063_n18700# 0.210644f
C2718 a_54579_n17803# a_53497_n18700# 5.37e-19
C2719 a_83141_n8770# VDD 0.016652f
C2720 a_89407_n6960# a_89407_n7865# 0.024773f
C2721 a_82573_n13190# a_82573_n14095# 0.005903f
C2722 a_99667_n19525# VDD 0.016281f
C2723 a_104527_n17715# a_104527_n18620# 0.006141f
C2724 a_114516_n35156# VDD 0.010487f
C2725 a_45445_n3548# a_45445_n6239# 0.008933f
C2726 a_47231_n3548# a_47753_n3548# 0.0284f
C2727 a_47753_n2651# a_46879_n3548# 8.45e-19
C2728 a_32353_n13316# a_32353_n14213# 0.005987f
C2729 a_33787_n13316# a_34699_n14213# 5.43e-19
C2730 a_54197_5639# VDD 0.042519f
C2731 a_32913_n14213# a_31831_n15110# 5.37e-19
C2732 a_60845_n13318# a_60285_n13318# 0.0284f
C2733 a_72596_n4978# VDD 0.03531f
C2734 a_89407_n9675# VDD 0.177586f
C2735 a_92601_n5150# a_92601_n9675# 0.032645f
C2736 a_92601_n4245# a_93131_n3340# 0.028522f
C2737 a_107339_n20430# VDD 0.392932f
C2738 a_82573_n18620# a_82573_n19525# 0.005903f
C2739 a_87433_n7865# IN_POS 0.00603f
C2740 a_109695_n16810# a_110225_n14095# 0.012586f
C2741 a_111063_n13190# a_111631_n13190# 0.027101f
C2742 a_79151_5639# a_79151_4481# 0.004047f
C2743 a_44363_n8930# a_44885_n8033# 0.0284f
C2744 a_47231_n8033# a_46879_n8930# 0.053799f
C2745 a_35781_n17801# a_35221_n17801# 0.0284f
C2746 a_58329_n18700# a_58851_n17803# 0.0284f
C2747 a_59411_n17803# a_60285_n18700# 8.45e-19
C2748 a_100803_n1530# VDD 0.177586f
C2749 a_95943_n8770# a_95105_n8770# 0.028522f
C2750 a_89407_n14095# a_90245_n15000# 0.028522f
C2751 a_63161_n17803# IBNOUT 0.008675f
C2752 a_111063_n20430# VDD 0.016652f
C2753 a_109695_n19525# a_111063_n18620# 2.31e-19
C2754 VDD OUT 47.331f
C2755 a_53497_n3550# a_54019_n3550# 0.0284f
C2756 a_51711_n3550# a_51711_n6241# 0.009307f
C2757 a_39531_n14213# a_40053_n13316# 0.0284f
C2758 a_65677_n13318# a_65677_n14215# 0.011408f
C2759 a_64595_n14215# a_66029_n14215# 0.014106f
C2760 a_105933_n2435# VDD 0.016652f
C2761 a_99667_n4245# a_100235_n4245# 0.027101f
C2762 a_32353_n12419# I1U 0.002649f
C2763 a_113081_7563# a_113081_6405# 0.004047f
C2764 a_54019_n7138# a_54019_n8035# 0.005987f
C2765 a_53497_n8035# a_54579_n8932# 5.37e-19
C2766 a_38097_n17801# a_38097_n19595# 0.005987f
C2767 a_64243_n18700# a_63161_n19597# 5.37e-19
C2768 a_75585_n9297# I1N 0.159888f
C2769 a_63683_n17803# a_63683_n18700# 0.005987f
C2770 a_109695_n4245# VDD 0.399575f
C2771 a_100235_n8770# a_100235_n9675# 0.005903f
C2772 a_94537_n15000# a_95105_n15000# 0.027101f
C2773 a_43817_n29181# a_43817_n30339# 0.004047f
C2774 a_33787_n3548# a_34347_n3548# 0.0284f
C2775 a_37968_11614# VDD 0.009062f
C2776 a_47753_n12419# a_47753_n13316# 0.005987f
C2777 a_45445_n14213# a_45797_n14213# 0.210644f
C2778 a_48313_n13316# a_47231_n14213# 5.37e-19
C2779 a_81205_n5150# a_82573_n1530# 7.4e-19
C2780 a_83709_n15000# VDD 0.121044f
C2781 a_94537_n20430# a_94537_n21335# 0.005903f
C2782 a_34699_n8033# a_35221_n8033# 0.0284f
C2783 a_61515_10448# VDD 0.021515f
C2784 a_59763_n8035# a_57977_n8932# 0.006457f
C2785 a_58851_n8035# a_59411_n8932# 0.0284f
C2786 a_81205_n9675# a_82573_n6960# 0.002134f
C2787 a_81205_n7865# a_81735_n6960# 0.028522f
C2788 a_90245_n18620# VDD 1.18674f
C2789 a_49755_n33224# VDD 0.05812f
C2790 a_45138_24920# a_45138_24195# 0.006281f
C2791 a_45706_24920# a_46274_24920# 0.017228f
C2792 a_44608_24195# a_45706_24195# 1.81e-19
C2793 a_30724_6405# a_30724_5639# 0.00778f
C2794 a_40965_n3548# a_42047_n4445# 5.37e-19
C2795 a_41487_n2651# a_41487_n3548# 0.005987f
C2796 a_89563_13546# VDD 0.021314f
C2797 a_66029_n3550# a_66029_n6241# 0.009483f
C2798 a_63161_n4447# a_63683_n4447# 0.0284f
C2799 a_51151_n13318# a_51711_n14215# 0.0284f
C2800 a_53145_n13318# a_53497_n14215# 0.053799f
C2801 a_86903_n5150# a_87433_n3340# 0.012586f
C2802 a_93131_n18620# VDD 0.137705f
C2803 a_110225_n6055# a_110225_n6960# 0.006141f
C2804 a_77776_n36322# VDD 0.029536f
C2805 a_48391_7563# a_48391_6405# 0.004047f
C2806 a_40965_n8033# a_40053_n8033# 5.43e-19
C2807 a_114516_13546# VDD 0.02603f
C2808 a_63161_n8932# a_64243_n8932# 5.37e-19
C2809 a_63683_n8035# a_63683_n8932# 0.005987f
C2810 a_65677_n8932# a_66551_n8035# 5.43e-19
C2811 a_50629_n17803# a_50629_n19597# 0.005987f
C2812 a_87433_n7865# a_88271_n7865# 0.027101f
C2813 a_82573_n8770# VDD 0.016652f
C2814 a_98829_n19525# VDD 0.121044f
C2815 a_113110_n35156# VDD 0.017204f
C2816 a_47231_n3548# a_46879_n3548# 0.16936f
C2817 a_44363_n4445# a_44885_n3548# 0.0284f
C2818 a_55601_6405# VDD 0.034176f
C2819 a_33265_n14213# a_34699_n14213# 0.005986f
C2820 a_34347_n13316# a_34347_n14213# 0.01664f
C2821 a_60285_n12421# a_60285_n13318# 0.005987f
C2822 a_60845_n13318# a_59763_n14215# 5.37e-19
C2823 a_57977_n14215# a_58329_n14215# 0.210644f
C2824 a_75602_n4019# VDD 0.027393f
C2825 a_94537_n2435# a_94537_n3340# 0.005903f
C2826 a_88839_n9675# VDD 0.02546f
C2827 a_106501_n19525# VDD 0.121044f
C2828 a_83141_n18620# a_83709_n18620# 0.027101f
C2829 a_47231_n8033# a_46319_n8033# 5.43e-19
C2830 a_32913_n18698# a_33265_n18698# 0.210644f
C2831 a_34347_n17801# a_34347_n19595# 0.011408f
C2832 a_35781_n17801# a_34699_n18698# 5.37e-19
C2833 a_35221_n16904# a_35221_n17801# 0.005987f
C2834 a_60845_n17803# a_60285_n17803# 0.0284f
C2835 a_59411_n17803# a_59411_n19597# 0.01664f
C2836 a_100235_n1530# VDD 0.02546f
C2837 a_95105_n7865# a_95105_n8770# 0.024773f
C2838 a_95943_n8770# a_94537_n8770# 2.31e-19
C2839 a_93131_n8770# a_93969_n8770# 0.027101f
C2840 a_65677_n17803# IBNOUT 0.004325f
C2841 a_87433_n14095# a_87433_n15000# 0.024773f
C2842 a_88839_n14095# a_90245_n15000# 2.31e-19
C2843 a_110225_n20430# VDD 0.121415f
C2844 a_109695_n19525# a_110225_n18620# 0.028522f
C2845 a_66016_n35156# IBNOUT 5.91e-19
C2846 a_71864_6405# OUT 0.001942f
C2847 a_95414_6405# a_95414_5639# 0.00778f
C2848 a_50629_n4447# a_51151_n3550# 0.0284f
C2849 a_53497_n3550# a_53145_n3550# 0.062551f
C2850 a_42047_n13316# a_41487_n13316# 0.0284f
C2851 a_64595_n14215# a_65117_n13318# 0.0284f
C2852 a_105365_n2435# VDD 0.016652f
C2853 a_100803_n3340# a_100803_n4245# 0.024773f
C2854 a_88271_n19525# a_88271_n20430# 0.005903f
C2855 a_89407_n19525# a_90245_n20430# 0.028522f
C2856 a_31831_n13316# I1U 0.008518f
C2857 a_51711_n8035# a_51711_n8932# 0.006457f
C2858 a_53497_n8035# a_54019_n8035# 0.0284f
C2859 a_38619_n17801# a_39179_n18698# 0.0284f
C2860 a_65677_n17803# a_67111_n19597# 0.018216f
C2861 a_64595_n18700# a_66029_n18700# 0.005986f
C2862 a_72603_n9297# I1N 0.158318f
C2863 a_113037_n3340# VDD 0.399226f
C2864 a_92601_n15905# a_93969_n15905# 2.31e-19
C2865 a_93131_n15000# a_93131_n15905# 0.024773f
C2866 a_71896_n34390# a_71896_n35156# 0.00778f
C2867 a_36562_11614# VDD 0.009062f
C2868 a_60285_n2653# a_60285_n3550# 0.005987f
C2869 a_59763_n3550# a_60845_n4447# 5.37e-19
C2870 a_46879_n13316# a_47753_n13316# 5.43e-19
C2871 a_81205_n5150# a_81735_n1530# 0.032766f
C2872 a_83141_n15000# VDD 0.016281f
C2873 a_34699_n8033# a_34347_n8930# 0.053799f
C2874 a_31831_n8930# a_32353_n8033# 0.0284f
C2875 a_60109_10448# VDD 0.029536f
C2876 a_46879_n17801# a_47753_n17801# 0.004425f
C2877 a_84547_n6960# a_83709_n6960# 0.042385f
C2878 a_81205_n9675# a_81735_n6960# 0.012586f
C2879 a_89407_n15905# VDD 0.138244f
C2880 a_105933_n9675# a_106501_n9675# 0.027101f
C2881 a_48349_n33224# VDD 0.073394f
C2882 a_44608_24195# a_45138_24195# 0.017843f
C2883 a_41487_n2651# a_40613_n3548# 8.45e-19
C2884 a_39179_n3548# a_39179_n6239# 0.008933f
C2885 a_40965_n3548# a_41487_n3548# 0.0284f
C2886 a_85089_n36322# VCM 0.002253f
C2887 a_65117_n3550# a_65677_n3550# 0.037577f
C2888 a_53145_n13318# a_52585_n13318# 0.0284f
C2889 a_86903_n5150# a_86903_n4245# 0.086339f
C2890 a_88839_n1530# a_88839_n2435# 0.005903f
C2891 a_92601_n19525# VDD 0.399575f
C2892 a_79182_n35156# VDD 0.009062f
C2893 a_100235_n21335# a_100803_n21335# 0.027101f
C2894 a_83725_n28415# a_83725_n29181# 0.00778f
C2895 a_66058_n28415# IBNOUT 6.21e-20
C2896 a_39531_n8033# a_40613_n8930# 5.37e-19
C2897 a_40053_n7136# a_40053_n8033# 0.005987f
C2898 a_63161_n8932# a_63683_n8932# 0.0284f
C2899 a_51151_n17803# a_51711_n18700# 0.0284f
C2900 a_86903_n9675# a_88271_n8770# 0.002134f
C2901 a_81735_n8770# VDD 0.149203f
C2902 a_88839_n6960# a_88839_n7865# 0.005903f
C2903 a_100803_n18620# VDD 0.138244f
C2904 a_83141_n13190# a_83709_n13190# 0.027101f
C2905 a_84547_n6055# IN_POS 0.001247f
C2906 a_81735_n13190# a_81735_n14095# 0.024773f
C2907 a_81205_n16810# a_82573_n14095# 0.002134f
C2908 a_114516_n34390# VDD 0.013383f
C2909 a_54197_6405# VDD 0.029136f
C2910 a_33265_n14213# a_33787_n13316# 0.0284f
C2911 a_59411_n13318# a_60285_n13318# 5.43e-19
C2912 a_72596_n4019# VDD 0.027393f
C2913 a_88271_n9675# VDD 0.02546f
C2914 a_92601_n5150# a_93131_n6055# 0.035071f
C2915 a_105933_n19525# VDD 0.016281f
C2916 a_81205_n19525# a_82573_n19525# 2.31e-19
C2917 a_81735_n18620# a_81735_n19525# 0.024773f
C2918 a_110225_n13190# a_111063_n13190# 0.027101f
C2919 a_77747_5639# a_77747_4481# 0.004047f
C2920 a_45797_n8033# a_46879_n8930# 5.37e-19
C2921 a_46319_n7136# a_46319_n8033# 0.005987f
C2922 a_31831_n17801# a_31831_n19595# 0.005987f
C2923 a_60285_n16906# a_60285_n17803# 0.005987f
C2924 a_57977_n18700# a_58329_n18700# 0.210644f
C2925 a_60845_n17803# a_59763_n18700# 5.37e-19
C2926 a_99667_n1530# VDD 0.02546f
C2927 a_88839_n14095# a_89407_n14095# 0.027101f
C2928 a_86903_n16810# a_88271_n15905# 0.002134f
C2929 a_109695_n21335# a_111063_n18620# 0.002134f
C2930 a_53497_n3550# a_52585_n3550# 5.43e-19
C2931 a_42047_n13316# a_40965_n14213# 5.37e-19
C2932 a_39179_n14213# a_39531_n14213# 0.210644f
C2933 a_41487_n12419# a_41487_n13316# 0.005987f
C2934 a_67111_n13318# a_66551_n13318# 0.0284f
C2935 a_98829_n4245# a_99667_n4245# 0.027101f
C2936 a_104527_n2435# VDD 0.149203f
C2937 a_88839_n19525# a_90245_n20430# 2.31e-19
C2938 a_55635_n34390# a_55635_n35156# 0.00778f
C2939 a_50629_n8932# a_51151_n8035# 0.0284f
C2940 a_53497_n8035# a_53145_n8932# 0.053799f
C2941 a_64595_n18700# a_65117_n17803# 0.0284f
C2942 a_65677_n17803# a_66551_n18700# 8.45e-19
C2943 a_112199_n2435# VDD 0.121415f
C2944 a_99667_n8770# a_99667_n9675# 0.005903f
C2945 a_92601_n15905# a_93131_n15905# 0.028522f
C2946 a_93969_n15000# a_94537_n15000# 0.027101f
C2947 a_42413_n29181# a_42413_n30339# 0.004047f
C2948 a_35221_n2651# a_35221_n3548# 0.005987f
C2949 a_34699_n3548# a_35781_n4445# 5.37e-19
C2950 a_57977_n3550# a_57977_n6241# 0.009307f
C2951 a_59763_n3550# a_60285_n3550# 0.0284f
C2952 a_37968_12380# VDD 0.009062f
C2953 a_94537_n14095# IBPOUT 0.00243f
C2954 a_44885_n13316# a_45445_n14213# 0.0284f
C2955 a_46879_n13316# a_47231_n14213# 0.053799f
C2956 a_82573_n15000# VDD 0.016281f
C2957 a_106501_n4245# a_107339_n6960# 0.042385f
C2958 a_93969_n20430# a_93969_n21335# 0.005903f
C2959 a_34699_n8033# a_33787_n8033# 5.43e-19
C2960 a_60285_n7138# a_60285_n8035# 0.005987f
C2961 a_59763_n8035# a_60845_n8932# 5.37e-19
C2962 a_61515_11614# VDD 0.011958f
C2963 a_46879_n17801# a_47231_n18698# 0.062551f
C2964 a_44363_n17801# a_45797_n18698# 1.57e-19
C2965 a_84547_n6960# a_83141_n6960# 0.002302f
C2966 a_81205_n9675# a_81205_n7865# 0.086469f
C2967 a_88839_n15905# VDD 0.01295f
C2968 a_87433_n14095# IN_POS 0.00603f
C2969 a_43848_n36322# VDD 0.024605f
C2970 a_100803_n15905# a_101641_n18620# 0.042385f
C2971 a_45138_24920# a_45706_24920# 0.017228f
C2972 a_44608_24195# a_46274_24920# 9.58e-21
C2973 a_38097_n4445# a_38619_n3548# 0.0284f
C2974 a_40965_n3548# a_40613_n3548# 0.16936f
C2975 a_83683_n36322# VCM 0.002253f
C2976 a_50629_n13318# a_50629_n15112# 0.005987f
C2977 a_52585_n12421# a_52585_n13318# 0.005987f
C2978 a_53145_n13318# a_52063_n14215# 5.37e-19
C2979 a_92601_n21335# VDD 1.40049f
C2980 a_77776_n35156# VDD 0.017204f
C2981 a_32088_11614# a_32088_10448# 0.004007f
C2982 a_39531_n8033# a_40053_n8033# 0.0284f
C2983 a_39179_n8033# a_40613_n8930# 1.57e-19
C2984 a_42047_n7136# a_42047_n8930# 0.005987f
C2985 a_113110_13546# VDD 0.029536f
C2986 a_65117_n8035# a_65677_n8932# 0.0284f
C2987 a_66029_n8035# a_64243_n8932# 0.006457f
C2988 a_53145_n17803# a_54019_n17803# 0.006769f
C2989 a_84547_n8770# VDD 0.399226f
C2990 a_86903_n9675# a_87433_n8770# 0.012586f
C2991 a_100235_n18620# VDD 0.01295f
C2992 a_81205_n16810# a_81735_n14095# 0.012586f
C2993 a_113110_n34390# VDD 0.017204f
C2994 a_104527_n17715# a_103997_n21335# 0.035071f
C2995 a_96818_n29181# a_96818_n30339# 0.004047f
C2996 a_45797_n3548# a_46879_n3548# 0.011365f
C2997 a_46319_n2651# a_46319_n3548# 0.005987f
C2998 a_55601_7563# VDD 0.00658f
C2999 a_35781_n13316# a_35221_n13316# 0.0284f
C3000 a_75602_n3060# VDD 0.03531f
C3001 a_59411_n13318# a_59763_n14215# 0.053799f
C3002 a_57417_n13318# a_57977_n14215# 0.0284f
C3003 a_87433_n9675# VDD 0.150485f
C3004 a_93969_n2435# a_93969_n3340# 0.005903f
C3005 a_105365_n19525# VDD 0.016281f
C3006 a_81205_n19525# a_81735_n19525# 0.028522f
C3007 a_82573_n18620# a_83141_n18620# 0.027101f
C3008 a_81205_n21335# a_82573_n19525# 0.002134f
C3009 a_84547_n18620# a_84547_n20430# 0.011861f
C3010 a_109695_n16810# a_111063_n13190# 0.002563f
C3011 a_48313_n7136# a_48313_n8930# 0.005987f
C3012 a_45797_n8033# a_46319_n8033# 0.0284f
C3013 a_45445_n8033# a_46879_n8930# 1.57e-19
C3014 a_32353_n17801# a_32913_n18698# 0.0284f
C3015 a_56895_n17803# a_56895_n19597# 0.005987f
C3016 a_98829_n1530# VDD 0.150485f
C3017 a_94537_n7865# a_94537_n8770# 0.005903f
C3018 a_113037_n20430# VDD 0.392932f
C3019 a_63683_n16009# IBNOUT 0.004702f
C3020 a_86903_n16810# a_87433_n15905# 0.012586f
C3021 a_109695_n21335# a_110225_n18620# 0.012586f
C3022 a_71864_7563# OUT 0.003757f
C3023 a_66016_n34390# IBNOUT 5.91e-19
C3024 a_96818_7563# a_96818_6405# 0.004047f
C3025 a_52063_n3550# a_53145_n3550# 0.00117f
C3026 a_52585_n2653# a_52585_n3550# 0.005987f
C3027 a_40613_n13316# a_41487_n13316# 5.43e-19
C3028 a_66551_n12421# a_66551_n13318# 0.005987f
C3029 a_67111_n13318# a_66029_n14215# 5.37e-19
C3030 a_64243_n14215# a_64595_n14215# 0.210644f
C3031 a_106501_n1530# VDD 0.177586f
C3032 a_100235_n3340# a_100235_n4245# 0.005903f
C3033 a_87433_n19525# a_87433_n20430# 0.024773f
C3034 a_88839_n19525# a_89407_n19525# 0.027101f
C3035 a_53497_n8035# a_52585_n8035# 5.43e-19
C3036 a_40613_n17801# a_41487_n17801# 0.004425f
C3037 a_65677_n17803# a_65677_n19597# 0.01664f
C3038 a_75585_n8397# I1N 0.144473f
C3039 a_67111_n17803# a_66551_n17803# 0.0284f
C3040 a_111631_n2435# VDD 0.016652f
C3041 a_100235_n8770# a_100803_n8770# 0.027101f
C3042 a_34699_n3548# a_35221_n3548# 0.0284f
C3043 a_32913_n3548# a_32913_n6239# 0.008933f
C3044 a_35221_n2651# a_34347_n3548# 8.45e-19
C3045 a_59763_n3550# a_59411_n3550# 0.062551f
C3046 a_56895_n4447# a_57417_n3550# 0.0284f
C3047 a_36562_12380# VDD 0.009062f
C3048 a_93969_n14095# IBPOUT 0.003731f
C3049 a_46879_n13316# a_46319_n13316# 0.0284f
C3050 a_81735_n15000# VDD 0.121044f
C3051 a_105933_n4245# a_107339_n6960# 0.002302f
C3052 a_94537_n20430# a_95105_n20430# 0.027101f
C3053 VDD IBNOUT 1.55863f
C3054 a_33787_n7136# a_33787_n8033# 0.005987f
C3055 a_33265_n8033# a_34347_n8930# 5.37e-19
C3056 a_59763_n8035# a_60285_n8035# 0.0284f
C3057 a_57977_n8035# a_57977_n8932# 0.006457f
C3058 a_60109_11614# VDD 0.017204f
C3059 a_46879_n17801# a_46319_n17801# 0.037577f
C3060 a_44363_n17801# a_45445_n18698# 5.37e-19
C3061 a_47753_n16904# a_48313_n17801# 0.0284f
C3062 a_44885_n16904# a_44885_n17801# 0.005987f
C3063 a_81735_n6055# a_81735_n6960# 0.006141f
C3064 a_88271_n15905# VDD 0.023101f
C3065 a_105365_n9675# a_105933_n9675# 0.027101f
C3066 a_100235_n15905# a_101641_n18620# 0.002302f
C3067 a_42442_n36322# VDD 0.029536f
C3068 a_44608_24195# a_45706_24920# 1.81e-19
C3069 a_66029_n3550# a_67111_n4447# 5.37e-19
C3070 a_85089_10448# VDD 0.05812f
C3071 a_66551_n2653# a_66551_n3550# 0.005987f
C3072 a_53145_n13318# a_51711_n14215# 1.57e-19
C3073 a_88271_n1530# a_88271_n2435# 0.005903f
C3074 a_95943_n17715# VDD 0.509696f
C3075 a_110225_n6055# a_109695_n9675# 0.035071f
C3076 a_99667_n21335# a_100235_n21335# 0.027101f
C3077 a_79182_n34390# VDD 0.011958f
C3078 a_71896_10448# OUT 0.003436f
C3079 a_40965_n8033# a_41487_n7136# 0.0284f
C3080 a_53145_n17803# a_53497_n18700# 0.16936f
C3081 a_88271_n6960# a_88271_n7865# 0.005903f
C3082 a_83709_n7865# VDD 0.121044f
C3083 a_99667_n18620# VDD 0.023101f
C3084 a_84547_n6960# IN_POS 0.021832f
C3085 a_82573_n13190# a_83141_n13190# 0.027101f
C3086 a_114516_n33224# VDD 0.02294f
C3087 a_42442_11614# a_42442_10448# 0.004007f
C3088 a_48313_n2651# a_48313_n4445# 0.005987f
C3089 a_45445_n3548# a_46879_n3548# 9.78e-20
C3090 a_45797_n3548# a_46319_n3548# 0.0284f
C3091 a_35781_n13316# a_34699_n14213# 5.37e-19
C3092 a_32913_n14213# a_33265_n14213# 0.210644f
C3093 a_35221_n12419# a_35221_n13316# 0.005987f
C3094 a_59411_n13318# a_58851_n13318# 0.0284f
C3095 a_72596_n3060# VDD 0.03531f
C3096 a_95105_n2435# a_95943_n3340# 0.028522f
C3097 a_89407_n8770# VDD 0.121415f
C3098 a_104527_n19525# VDD 0.121044f
C3099 a_81205_n21335# a_81735_n19525# 0.012586f
C3100 a_87433_n6960# IN_POS 0.00603f
C3101 a_109695_n16810# a_110225_n13190# 0.044257f
C3102 a_79151_6405# a_79151_5639# 0.00778f
C3103 a_47231_n8033# a_47753_n7136# 0.0284f
C3104 a_57417_n17803# a_57977_n18700# 0.0284f
C3105 a_98299_n5150# VDD 1.40049f
C3106 a_112199_n19525# VDD 0.121044f
C3107 a_88271_n14095# a_88839_n14095# 0.027101f
C3108 a_109695_n21335# a_109695_n19525# 0.086339f
C3109 a_113037_n18620# a_112199_n18620# 0.032618f
C3110 a_52063_n3550# a_52585_n3550# 0.0284f
C3111 a_51711_n3550# a_53145_n3550# 5.12e-19
C3112 a_54579_n2653# a_54579_n4447# 0.005987f
C3113 a_40613_n13316# a_40965_n14213# 0.053799f
C3114 a_38619_n13316# a_39179_n14213# 0.0284f
C3115 a_65677_n13318# a_66551_n13318# 5.43e-19
C3116 a_105933_n1530# VDD 0.02546f
C3117 a_86903_n21335# a_88271_n21335# 0.002563f
C3118 a_30724_n27257# a_30724_n28415# 0.004047f
C3119 a_54229_n34390# a_54229_n35156# 0.00778f
C3120 a_52585_n7138# a_52585_n8035# 0.005987f
C3121 a_52063_n8035# a_53145_n8932# 5.37e-19
C3122 a_40613_n17801# a_40965_n18698# 0.062551f
C3123 a_38097_n17801# a_39531_n18698# 1.57e-19
C3124 a_67111_n17803# a_66029_n18700# 5.37e-19
C3125 a_66551_n16906# a_66551_n17803# 0.005987f
C3126 a_64243_n18700# a_64595_n18700# 0.210644f
C3127 a_72603_n8397# I1N 0.134725f
C3128 a_98829_n8770# a_98829_n9675# 0.024773f
C3129 a_111063_n2435# VDD 0.016652f
C3130 a_93131_n15000# a_93969_n15000# 0.027101f
C3131 a_95943_n15000# a_95105_n15000# 0.028522f
C3132 a_43817_n28415# a_43817_n29181# 0.00778f
C3133 a_32353_n19595# I1U 0.002649f
C3134 a_31831_n4445# a_32353_n3548# 0.0284f
C3135 a_34699_n3548# a_34347_n3548# 0.16936f
C3136 a_59763_n3550# a_58851_n3550# 5.43e-19
C3137 a_93131_n14095# IBPOUT 0.050612f
C3138 a_46319_n12419# a_46319_n13316# 0.005987f
C3139 a_46879_n13316# a_45797_n14213# 5.37e-19
C3140 a_44363_n13316# a_44363_n15110# 0.005987f
C3141 a_45445_n12419# a_47231_n14213# 0.006457f
C3142 a_105933_n4245# a_106501_n4245# 0.027101f
C3143 a_104527_n4245# a_104527_n6055# 0.006141f
C3144 a_81205_n15905# VDD 0.393432f
C3145 a_32913_n1754# I1U 2.01e-19
C3146 a_93131_n20430# a_93131_n21335# 0.024773f
C3147 a_33265_n8033# a_33787_n8033# 0.0284f
C3148 a_32913_n8033# a_34347_n8930# 1.57e-19
C3149 a_35781_n7136# a_35781_n8930# 0.005987f
C3150 a_56895_n8932# a_57417_n8035# 0.0284f
C3151 a_61515_12380# VDD 0.009062f
C3152 a_59763_n8035# a_59411_n8932# 0.053799f
C3153 a_44363_n17801# a_44885_n17801# 0.0284f
C3154 a_46879_n17801# a_45797_n18698# 0.00117f
C3155 a_106501_n8770# a_106501_n9675# 0.024773f
C3156 a_87433_n15905# VDD 0.113729f
C3157 a_43848_n35156# VDD 0.009062f
C3158 a_98829_n15905# a_98829_n17715# 0.006141f
C3159 a_100235_n15905# a_100803_n15905# 0.027101f
C3160 a_44608_24195# a_45138_24920# 0.017843f
C3161 a_39531_n3548# a_40613_n3548# 0.011365f
C3162 a_40053_n2651# a_40053_n3548# 0.005987f
C3163 a_83683_10448# VDD 0.073394f
C3164 a_64243_n3550# a_64243_n6241# 0.009307f
C3165 a_66029_n3550# a_66551_n3550# 0.0284f
C3166 a_54019_n12421# a_54579_n13318# 0.0284f
C3167 a_93131_n17715# VDD 0.41764f
C3168 a_77776_n34390# VDD 0.017204f
C3169 a_100803_n20430# a_100803_n21335# 0.024773f
C3170 a_30682_11614# a_30682_10448# 0.004007f
C3171 a_66058_n27257# IBNOUT 6.21e-20
C3172 a_39179_n8033# a_38619_n8033# 0.0284f
C3173 a_39531_n8033# a_38097_n8930# 1.57e-19
C3174 a_66029_n8035# a_67111_n8932# 5.37e-19
C3175 a_108636_10448# VDD 0.021515f
C3176 a_66551_n7138# a_66551_n8035# 0.005987f
C3177 a_53145_n17803# a_52585_n17803# 0.0284f
C3178 a_50629_n17803# a_52063_n18700# 1.57e-19
C3179 a_83141_n7865# VDD 0.016281f
C3180 a_88839_n6960# a_89407_n6960# 0.027101f
C3181 a_98829_n18620# VDD 0.113729f
C3182 a_107339_n18620# a_107339_n17715# 0.088786f
C3183 a_113110_n33224# VDD 0.029536f
C3184 a_95414_n29181# a_95414_n30339# 0.004047f
C3185 a_61484_5639# a_61484_4481# 0.004047f
C3186 a_47231_n3548# a_47753_n2651# 0.0284f
C3187 a_34347_n13316# a_35221_n13316# 5.43e-19
C3188 a_56895_n13318# a_56895_n15112# 0.005987f
C3189 a_59411_n13318# a_58329_n14215# 5.37e-19
C3190 a_58851_n12421# a_58851_n13318# 0.005987f
C3191 a_88839_n8770# VDD 0.016652f
C3192 a_93131_n2435# a_93131_n3340# 0.024773f
C3193 a_94537_n2435# a_95943_n3340# 2.31e-19
C3194 a_106501_n18620# VDD 0.138244f
C3195 a_81735_n18620# a_82573_n18620# 0.027101f
C3196 a_86903_n7865# IN_POS 0.001743f
C3197 a_45797_n8033# a_44363_n8930# 1.57e-19
C3198 a_45445_n8033# a_44885_n8033# 0.0284f
C3199 a_34347_n17801# a_35221_n17801# 0.004425f
C3200 a_59411_n17803# a_60285_n17803# 0.006769f
C3201 a_95105_n7865# a_95943_n8770# 0.028522f
C3202 a_95105_n9675# VDD 0.177586f
C3203 a_93969_n7865# a_93969_n8770# 0.005903f
C3204 a_111631_n19525# VDD 0.016281f
C3205 a_66029_n16906# IBNOUT 0.008853f
C3206 a_113037_n18620# a_111631_n18620# 7.35e-19
C3207 a_37968_n34390# a_37968_n35156# 0.00778f
C3208 a_66016_n33224# IBNOUT 5.91e-19
C3209 a_95414_7563# a_95414_6405# 0.004047f
C3210 a_53497_n3550# a_54019_n2653# 0.0284f
C3211 a_114485_4481# VDD 0.002225f
C3212 a_40613_n13316# a_40053_n13316# 0.0284f
C3213 a_63683_n13318# a_64243_n14215# 0.0284f
C3214 a_65677_n13318# a_66029_n14215# 0.053799f
C3215 a_101641_n3340# a_101641_n6960# 0.011861f
C3216 a_99667_n3340# a_99667_n4245# 0.005903f
C3217 a_105365_n1530# VDD 0.02546f
C3218 a_88271_n19525# a_88839_n19525# 0.027101f
C3219 a_86903_n21335# a_87433_n21335# 0.044257f
C3220 a_54579_n7138# a_54579_n8932# 0.005987f
C3221 a_51711_n8035# a_53145_n8932# 1.57e-19
C3222 a_52063_n8035# a_52585_n8035# 0.0284f
C3223 a_40613_n17801# a_40053_n17801# 0.037577f
C3224 a_38619_n16904# a_38619_n17801# 0.005987f
C3225 a_41487_n16904# a_42047_n17801# 0.0284f
C3226 a_38097_n17801# a_39179_n18698# 5.37e-19
C3227 a_63161_n17803# a_63161_n19597# 0.005987f
C3228 a_99667_n8770# a_100235_n8770# 0.027101f
C3229 a_110225_n2435# VDD 0.149203f
C3230 a_73268_n30339# VDD 0.00658f
C3231 a_95943_n15000# a_94537_n15000# 2.31e-19
C3232 a_92601_n15905# a_93969_n15000# 2.31e-19
C3233 a_95105_n14095# a_95105_n15000# 0.024773f
C3234 a_58329_n3550# a_59411_n3550# 0.00117f
C3235 a_58851_n2653# a_58851_n3550# 0.005987f
C3236 a_37968_13546# VDD 0.021314f
C3237 a_46879_n13316# a_45445_n14213# 1.57e-19
C3238 a_84547_n15000# VDD 0.392932f
C3239 a_32353_n1754# I1U 0.002649f
C3240 a_93969_n20430# a_94537_n20430# 0.027101f
C3241 a_34699_n8033# a_35221_n7136# 0.0284f
C3242 a_60109_12380# VDD 0.017204f
C3243 a_59763_n8035# a_58851_n8035# 5.43e-19
C3244 a_46879_n17801# a_45445_n18698# 5.12e-19
C3245 a_81735_n6055# a_81205_n9675# 0.03483f
C3246 a_89407_n15000# VDD 0.121044f
C3247 a_104527_n9675# a_105365_n9675# 0.027101f
C3248 a_42442_n35156# VDD 0.017204f
C3249 a_30724_7563# a_30724_6405# 0.004047f
C3250 a_42047_n2651# a_42047_n4445# 0.005987f
C3251 a_39179_n3548# a_40613_n3548# 9.78e-20
C3252 a_39531_n3548# a_40053_n3548# 0.0284f
C3253 a_85089_11614# VDD 0.046892f
C3254 a_63161_n4447# a_63683_n3550# 0.0284f
C3255 a_66029_n3550# a_65677_n3550# 0.062551f
C3256 a_53145_n13318# a_54579_n13318# 0.014106f
C3257 a_86903_n5150# a_88271_n2435# 0.002134f
C3258 a_87433_n1530# a_87433_n2435# 0.024773f
C3259 a_88839_n1530# a_89407_n1530# 0.027101f
C3260 a_113037_n6960# a_113037_n6055# 0.088786f
C3261 a_95943_n18620# VDD 1.25121f
C3262 a_79182_n33224# VDD 0.021515f
C3263 a_98829_n21335# a_99667_n21335# 0.027101f
C3264 a_71896_11614# OUT 0.001027f
C3265 a_39179_n8033# a_38097_n8930# 5.37e-19
C3266 a_38619_n7136# a_38619_n8033# 0.005987f
C3267 a_40053_n7136# a_40965_n8033# 5.43e-19
C3268 a_66029_n8035# a_66551_n8035# 0.0284f
C3269 a_107230_10448# VDD 0.021515f
C3270 a_64243_n8035# a_64243_n8932# 0.006457f
C3271 a_54019_n16906# a_54579_n17803# 0.0284f
C3272 a_53145_n17803# a_52063_n18700# 0.011365f
C3273 a_51151_n16906# a_51151_n17803# 0.005987f
C3274 a_50629_n17803# a_51711_n18700# 5.37e-19
C3275 a_87433_n6960# a_87433_n7865# 0.024773f
C3276 a_86903_n7865# a_88271_n7865# 2.31e-19
C3277 a_82573_n7865# VDD 0.016281f
C3278 a_81735_n13190# a_82573_n13190# 0.027101f
C3279 a_98299_n19525# VDD 0.393432f
C3280 a_108636_n36322# VDD 0.021314f
C3281 a_43848_12380# a_43848_11614# 0.00778f
C3282 a_45797_n3548# a_44363_n4445# 1.57e-19
C3283 a_45445_n3548# a_44885_n3548# 0.0284f
C3284 a_48313_n2651# a_46879_n3548# 0.018216f
C3285 a_32353_n13316# a_32913_n14213# 0.0284f
C3286 a_34347_n13316# a_34699_n14213# 0.053799f
C3287 a_59411_n13318# a_57977_n14215# 1.57e-19
C3288 a_92601_n5150# a_93969_n4245# 0.002134f
C3289 a_88271_n8770# VDD 0.016652f
C3290 a_94537_n2435# a_95105_n2435# 0.027101f
C3291 a_81205_n19525# a_82573_n18620# 2.31e-19
C3292 a_105933_n18620# VDD 0.01295f
C3293 a_86903_n9675# IN_POS 0.093087f
C3294 a_77747_6405# a_77747_5639# 0.00778f
C3295 a_46319_n7136# a_47231_n8033# 5.43e-19
C3296 a_44885_n7136# a_44885_n8033# 0.005987f
C3297 a_45445_n8033# a_44363_n8930# 5.37e-19
C3298 a_31831_n17801# a_33265_n18698# 1.57e-19
C3299 a_34347_n17801# a_34699_n18698# 0.062551f
C3300 a_59411_n17803# a_59763_n18700# 0.16936f
C3301 a_94537_n7865# a_95943_n8770# 2.31e-19
C3302 a_94537_n9675# VDD 0.02546f
C3303 a_86903_n16810# a_88271_n15000# 0.002134f
C3304 a_87433_n14095# a_88271_n14095# 0.027101f
C3305 a_89407_n13190# a_89407_n14095# 0.024773f
C3306 a_111063_n19525# VDD 0.016281f
C3307 a_64243_n16906# IBNOUT 0.239585f
C3308 a_110225_n17715# a_110225_n18620# 0.006141f
C3309 a_51711_n3550# a_51151_n3550# 0.0284f
C3310 a_52063_n3550# a_50629_n4447# 1.57e-19
C3311 a_40053_n12419# a_40053_n13316# 0.005987f
C3312 a_39179_n12419# a_40965_n14213# 0.006457f
C3313 a_38097_n13316# a_38097_n15110# 0.005987f
C3314 a_40613_n13316# a_39531_n14213# 5.37e-19
C3315 a_65677_n13318# a_65117_n13318# 0.0284f
C3316 a_104527_n1530# VDD 0.150485f
C3317 a_100235_n3340# a_100803_n3340# 0.027101f
C3318 a_89407_n18620# a_89407_n19525# 0.024773f
C3319 a_77747_n30339# VCM 0.003538f
C3320 a_53497_n8035# a_54019_n7138# 0.0284f
C3321 a_40613_n17801# a_39531_n18698# 0.00117f
C3322 a_38097_n17801# a_38619_n17801# 0.0284f
C3323 a_63683_n17803# a_64243_n18700# 0.0284f
C3324 a_112199_n1530# VDD 0.177586f
C3325 a_92601_n15905# a_93131_n15000# 0.028522f
C3326 a_92601_n16810# a_92601_n21335# 0.032645f
C3327 a_42413_n28415# a_42413_n29181# 0.00778f
C3328 a_33787_n2651# a_33787_n3548# 0.005987f
C3329 a_33265_n3548# a_34347_n3548# 0.011365f
C3330 a_60845_n2653# a_60845_n4447# 0.005987f
C3331 a_58329_n3550# a_58851_n3550# 0.0284f
C3332 a_57977_n3550# a_59411_n3550# 5.12e-19
C3333 a_47753_n12419# a_48313_n13316# 0.0284f
C3334 a_75585_n10073# a_75585_n10973# 0.005955f
C3335 a_83709_n14095# VDD 0.121415f
C3336 a_105365_n4245# a_105933_n4245# 0.027101f
C3337 a_31831_n2651# I1U 0.008518f
C3338 a_95943_n20430# a_95105_n20430# 0.028522f
C3339 a_33265_n8033# a_31831_n8930# 1.57e-19
C3340 a_32913_n8033# a_32353_n8033# 0.0284f
C3341 a_58851_n7138# a_58851_n8035# 0.005987f
C3342 a_58329_n8035# a_59411_n8932# 5.37e-19
C3343 a_88839_n15000# VDD 0.016281f
C3344 a_105933_n8770# a_105933_n9675# 0.005903f
C3345 a_43848_n34390# VDD 0.011958f
C3346 a_99667_n15905# a_100235_n15905# 0.027101f
C3347 a_40965_n3548# a_41487_n2651# 0.0284f
C3348 a_83683_11614# VDD 0.062166f
C3349 a_66029_n3550# a_65117_n3550# 5.43e-19
C3350 a_53145_n13318# a_54019_n12421# 5.43e-19
C3351 a_50629_n13318# a_52063_n14215# 1.57e-19
C3352 a_86903_n5150# a_87433_n2435# 0.012586f
C3353 a_95105_n15905# VDD 0.201f
C3354 a_77776_n33224# VDD 0.029536f
C3355 a_100235_n20430# a_100235_n21335# 0.005903f
C3356 a_32088_12380# a_32088_11614# 0.00778f
C3357 a_83725_n27257# a_83725_n28415# 0.004047f
C3358 OUT I1N 0.272652f
C3359 a_39531_n8033# a_40965_n8033# 0.014106f
C3360 VDD IBPOUT 3.44382f
C3361 a_63161_n8932# a_63683_n8035# 0.0284f
C3362 a_108636_11614# VDD 0.009062f
C3363 a_66029_n8035# a_65677_n8932# 0.053799f
C3364 a_53145_n17803# a_51711_n18700# 9.78e-20
C3365 a_50629_n17803# a_51151_n17803# 0.0284f
C3366 a_86903_n9675# a_88271_n7865# 0.002134f
C3367 a_90245_n6960# a_90245_n8770# 0.011861f
C3368 a_81735_n7865# VDD 0.121044f
C3369 a_86903_n7865# a_87433_n7865# 0.028522f
C3370 a_88271_n6960# a_88839_n6960# 0.027101f
C3371 a_81205_n16810# a_82573_n13190# 7.4e-19
C3372 a_107230_n36322# VDD 0.021314f
C3373 a_96818_n28415# a_96818_n29181# 0.00778f
C3374 a_60080_5639# a_60080_4481# 0.004047f
C3375 a_46319_n2651# a_47231_n3548# 5.43e-19
C3376 a_44885_n2651# a_44885_n3548# 0.005987f
C3377 a_45445_n3548# a_44363_n4445# 5.37e-19
C3378 a_34347_n13316# a_33787_n13316# 0.0284f
C3379 a_60285_n12421# a_60845_n13318# 0.0284f
C3380 a_87433_n8770# VDD 0.149203f
C3381 a_92601_n5150# a_93131_n4245# 0.012586f
C3382 a_81205_n21335# a_82573_n18620# 0.002134f
C3383 a_105365_n18620# VDD 0.023101f
C3384 a_81205_n19525# a_81735_n18620# 0.028522f
C3385 a_55635_12380# a_55635_11614# 0.00778f
C3386 a_45797_n8033# a_47231_n8033# 0.014106f
C3387 a_35221_n16904# a_35781_n17801# 0.0284f
C3388 a_32353_n16904# a_32353_n17801# 0.005987f
C3389 a_34347_n17801# a_33787_n17801# 0.037577f
C3390 a_31831_n17801# a_32913_n18698# 5.37e-19
C3391 a_59411_n17803# a_58851_n17803# 0.0284f
C3392 a_56895_n17803# a_58329_n18700# 1.57e-19
C3393 a_93969_n9675# VDD 0.02546f
C3394 a_94537_n7865# a_95105_n7865# 0.027101f
C3395 a_93131_n7865# a_93131_n8770# 0.024773f
C3396 a_86903_n16810# a_87433_n15000# 0.012586f
C3397 a_110225_n19525# VDD 0.121044f
C3398 a_63683_n15112# IBNOUT 0.004735f
C3399 a_36562_n34390# a_36562_n35156# 0.00778f
C3400 a_51151_n2653# a_51151_n3550# 0.005987f
C3401 a_52585_n2653# a_53497_n3550# 5.43e-19
C3402 a_51711_n3550# a_50629_n4447# 5.37e-19
C3403 a_114485_5639# VDD 0.002225f
C3404 a_40613_n13316# a_39179_n14213# 1.57e-19
C3405 a_65677_n13318# a_64595_n14215# 5.37e-19
C3406 a_65117_n12421# a_65117_n13318# 0.005987f
C3407 a_63161_n13318# a_63161_n15112# 0.005987f
C3408 a_98299_n4245# a_99667_n4245# 2.31e-19
C3409 a_103997_n5150# VDD 1.40049f
C3410 a_98829_n3340# a_98829_n4245# 0.024773f
C3411 a_87433_n19525# a_88271_n19525# 0.027101f
C3412 a_52063_n8035# a_50629_n8932# 1.57e-19
C3413 w_27790_n38888# VDD 96.053f
C3414 a_51711_n8035# a_51151_n8035# 0.0284f
C3415 a_40613_n17801# a_39179_n18698# 5.12e-19
C3416 a_65677_n17803# a_66551_n17803# 0.006769f
C3417 a_101641_n8770# a_100803_n8770# 0.028522f
C3418 a_111631_n1530# VDD 0.02546f
C3419 a_98829_n8770# a_99667_n8770# 0.027101f
C3420 a_94537_n14095# a_94537_n15000# 0.005903f
C3421 a_73268_n29181# VDD 0.034176f
C3422 a_33265_n3548# a_33787_n3548# 0.0284f
C3423 a_35781_n2651# a_35781_n4445# 0.005987f
C3424 a_32913_n3548# a_34347_n3548# 9.78e-20
C3425 a_59763_n3550# a_60285_n2653# 0.0284f
C3426 a_45445_n12419# a_45445_n14213# 0.006457f
C3427 a_46879_n13316# a_48313_n13316# 0.014106f
C3428 a_94537_n13190# IBPOUT 0.00243f
C3429 a_106501_n3340# a_106501_n4245# 0.024773f
C3430 a_83141_n14095# VDD 0.016652f
C3431 a_95105_n19525# a_95105_n20430# 0.024773f
C3432 a_93131_n20430# a_93969_n20430# 0.027101f
C3433 a_95943_n20430# a_94537_n20430# 2.31e-19
C3434 a_32353_n7136# a_32353_n8033# 0.005987f
C3435 a_33787_n7136# a_34699_n8033# 5.43e-19
C3436 a_32913_n8033# a_31831_n8930# 5.37e-19
C3437 a_57977_n8035# a_59411_n8932# 1.57e-19
C3438 a_58329_n8035# a_58851_n8035# 0.0284f
C3439 a_60845_n7138# a_60845_n8932# 0.005987f
C3440 a_61515_13546# VDD 0.024605f
C3441 a_46879_n17801# a_48313_n17801# 0.003256f
C3442 a_44363_n17801# a_44885_n16904# 0.0284f
C3443 a_47753_n16007# a_47753_n16904# 0.005987f
C3444 a_47231_n16904# a_47231_n18698# 0.009483f
C3445 a_84547_n6960# a_84547_n6055# 0.088786f
C3446 a_88271_n15000# VDD 0.016281f
C3447 a_42442_n34390# VDD 0.017204f
C3448 a_100803_n15000# a_100803_n15905# 0.024773f
C3449 a_87433_n13190# IN_POS 0.004984f
C3450 a_102756_n35156# a_102756_n36322# 0.004007f
C3451 a_39179_n3548# a_38619_n3548# 0.0284f
C3452 a_39531_n3548# a_38097_n4445# 1.57e-19
C3453 a_42047_n2651# a_40613_n3548# 0.018216f
C3454 a_85089_12380# VDD 0.061113f
C3455 a_64595_n3550# a_65677_n3550# 0.00117f
C3456 a_65117_n2653# a_65117_n3550# 0.005987f
C3457 a_51151_n12421# a_51151_n13318# 0.005987f
C3458 a_50629_n13318# a_51711_n14215# 5.37e-19
C3459 a_88271_n1530# a_88839_n1530# 0.027101f
C3460 a_94537_n15905# VDD 0.01901f
C3461 a_73302_n36322# VDD 0.021314f
C3462 a_71896_12380# OUT 0.001027f
C3463 a_39531_n8033# a_40053_n7136# 0.0284f
C3464 a_66029_n8035# a_65117_n8035# 5.43e-19
C3465 a_107230_11614# VDD 0.009062f
C3466 a_53497_n16906# a_53497_n18700# 0.0089f
C3467 a_83709_n6960# VDD 0.112244f
C3468 a_86903_n9675# a_87433_n7865# 0.012586f
C3469 a_81205_n16810# a_81735_n13190# 0.032766f
C3470 a_98299_n21335# VDD 0.921963f
C3471 a_108636_n35156# VDD 0.009062f
C3472 a_42442_12380# a_42442_11614# 0.00778f
C3473 a_46879_n2651# a_46879_n3548# 0.01664f
C3474 a_45797_n3548# a_47231_n3548# 0.005986f
C3475 a_34347_n13316# a_33265_n14213# 5.37e-19
C3476 a_33787_n12419# a_33787_n13316# 0.005987f
C3477 a_31831_n13316# a_31831_n15110# 0.005987f
C3478 a_32913_n12419# a_34699_n14213# 0.006457f
C3479 a_59411_n13318# a_60845_n13318# 0.014106f
C3480 a_93969_n2435# a_94537_n2435# 0.027101f
C3481 a_90245_n8770# VDD 0.399226f
C3482 a_104527_n18620# VDD 0.113729f
C3483 a_84547_n18620# a_83709_n18620# 0.042385f
C3484 a_81205_n21335# a_81735_n18620# 0.012586f
C3485 a_87433_n6055# IN_POS 0.005369f
C3486 a_105933_n21335# a_106501_n21335# 0.027101f
C3487 a_79151_7563# a_79151_6405# 0.004047f
C3488 a_45797_n8033# a_46319_n7136# 0.0284f
C3489 a_34347_n17801# a_33265_n18698# 0.00117f
C3490 a_31831_n17801# a_32353_n17801# 0.0284f
C3491 a_59411_n17803# a_58329_n18700# 0.011365f
C3492 a_57417_n16906# a_57417_n17803# 0.005987f
C3493 a_60285_n16906# a_60845_n17803# 0.0284f
C3494 a_56895_n17803# a_57977_n18700# 5.37e-19
C3495 a_93131_n9675# VDD 0.150485f
C3496 a_92601_n9675# a_93969_n9675# 0.002563f
C3497 a_112199_n18620# VDD 0.138244f
C3498 a_88839_n13190# a_88839_n14095# 0.005903f
C3499 a_86903_n16810# a_86903_n15905# 0.086339f
C3500 a_67422_11614# a_67422_10448# 0.004007f
C3501 a_52063_n3550# a_53497_n3550# 0.014106f
C3502 a_53145_n2653# a_53145_n3550# 0.011408f
C3503 a_41487_n12419# a_42047_n13316# 0.0284f
C3504 a_65677_n13318# a_64243_n14215# 1.57e-19
C3505 a_98299_n4245# a_98829_n4245# 0.028522f
C3506 a_99667_n3340# a_100235_n3340# 0.027101f
C3507 a_100803_n9675# VDD 0.150485f
C3508 a_88839_n18620# a_88839_n19525# 0.005903f
C3509 a_86903_n21335# a_88271_n20430# 0.002134f
C3510 a_77747_n29181# VCM 0.003538f
C3511 a_51151_n7138# a_51151_n8035# 0.005987f
C3512 a_51711_n8035# a_50629_n8932# 5.37e-19
C3513 a_65677_n17803# a_66029_n18700# 0.16936f
C3514 a_111063_n1530# VDD 0.02546f
C3515 a_101641_n8770# a_100235_n8770# 2.31e-19
C3516 a_100803_n7865# a_100803_n8770# 0.024773f
C3517 a_92601_n16810# a_93131_n17715# 0.035071f
C3518 a_71864_n29181# VDD 0.029136f
C3519 a_34699_n3548# a_35221_n2651# 0.0284f
C3520 a_36562_13546# VDD 0.021314f
C3521 a_58329_n3550# a_56895_n4447# 1.57e-19
C3522 a_57977_n3550# a_57417_n3550# 0.0284f
C3523 a_46879_n13316# a_47753_n12419# 5.43e-19
C3524 a_93969_n13190# IBPOUT 0.007416f
C3525 a_44363_n13316# a_45797_n14213# 1.57e-19
C3526 a_72603_n10073# a_72603_n10973# 0.005955f
C3527 a_104527_n4245# a_105365_n4245# 0.027101f
C3528 a_82573_n14095# VDD 0.016652f
C3529 a_33265_n8033# a_34699_n8033# 0.014106f
C3530 a_59763_n8035# a_60285_n7138# 0.0284f
C3531 a_46879_n17801# a_47753_n16904# 4.96e-19
C3532 a_105365_n8770# a_105365_n9675# 0.005903f
C3533 a_87433_n15000# VDD 0.121044f
C3534 a_98829_n15905# a_99667_n15905# 0.027101f
C3535 a_43848_n33224# VDD 0.021515f
C3536 a_86903_n16810# IN_POS 0.156237f
C3537 a_38619_n2651# a_38619_n3548# 0.005987f
C3538 a_39179_n3548# a_38097_n4445# 5.37e-19
C3539 a_40053_n2651# a_40965_n3548# 5.43e-19
C3540 a_67111_n2653# a_67111_n4447# 0.005987f
C3541 a_64595_n3550# a_65117_n3550# 0.0284f
C3542 a_64243_n3550# a_65677_n3550# 5.12e-19
C3543 a_83683_12380# VDD 0.076387f
C3544 a_50629_n13318# a_51151_n13318# 0.0284f
C3545 a_52585_n12421# a_53145_n13318# 0.0284f
C3546 a_93969_n15905# VDD 0.023101f
C3547 a_112199_n4245# a_113037_n6960# 0.042385f
C3548 a_99667_n20430# a_99667_n21335# 0.005903f
C3549 a_71896_n36322# VDD 0.021314f
C3550 a_30682_12380# a_30682_11614# 0.00778f
C3551 a_42047_n7136# a_41487_n7136# 0.0284f
C3552 a_108636_12380# VDD 0.009062f
C3553 a_65117_n7138# a_65117_n8035# 0.005987f
C3554 a_64595_n8035# a_65677_n8932# 5.37e-19
C3555 a_53145_n17803# a_54579_n17803# 0.08885f
C3556 a_83141_n6960# VDD 0.023105f
C3557 a_87433_n6960# a_88271_n6960# 0.027101f
C3558 a_101641_n17715# VDD 0.472471f
C3559 a_107230_n35156# VDD 0.009062f
C3560 a_106501_n15905# a_107339_n18620# 0.042385f
C3561 a_95414_n28415# a_95414_n29181# 0.00778f
C3562 a_61484_6405# a_61484_5639# 0.00778f
C3563 a_45797_n3548# a_46319_n2651# 0.0284f
C3564 a_34347_n13316# a_32913_n14213# 1.57e-19
C3565 a_56895_n13318# a_58329_n14215# 1.57e-19
C3566 a_59411_n13318# a_60285_n12421# 5.43e-19
C3567 a_89407_n7865# VDD 0.121044f
C3568 a_81205_n21335# a_81205_n19525# 0.086469f
C3569 a_84547_n18620# a_83141_n18620# 0.002302f
C3570 a_103997_n19525# VDD 0.393432f
C3571 a_54229_12380# a_54229_11614# 0.00778f
C3572 a_48313_n7136# a_47753_n7136# 0.0284f
C3573 a_34347_n17801# a_32913_n18698# 5.12e-19
C3574 a_59411_n17803# a_57977_n18700# 9.78e-20
C3575 a_56895_n17803# a_57417_n17803# 0.0284f
C3576 a_92601_n9675# a_93131_n9675# 0.044257f
C3577 a_95105_n8770# VDD 0.121415f
C3578 a_93969_n7865# a_94537_n7865# 0.027101f
C3579 a_111631_n18620# VDD 0.01295f
C3580 a_110225_n17715# a_109695_n21335# 0.035071f
C3581 a_52063_n3550# a_52585_n2653# 0.0284f
C3582 a_40613_n13316# a_42047_n13316# 0.014106f
C3583 a_114485_6405# VDD 0.002225f
C3584 a_39179_n12419# a_39179_n14213# 0.006457f
C3585 a_66551_n12421# a_67111_n13318# 0.0284f
C3586 a_100235_n9675# VDD 0.02546f
C3587 a_86903_n21335# a_87433_n20430# 0.012586f
C3588 a_77776_11614# a_77776_10448# 0.004007f
C3589 a_53145_n7138# a_54579_n8932# 0.018216f
C3590 a_52063_n8035# a_53497_n8035# 0.005986f
C3591 a_41487_n16007# a_41487_n16904# 0.005987f
C3592 a_38097_n17801# a_38619_n16904# 0.0284f
C3593 a_40613_n17801# a_42047_n17801# 0.003256f
C3594 a_40965_n16904# a_40965_n18698# 0.009483f
C3595 a_63161_n17803# a_64595_n18700# 1.57e-19
C3596 a_65677_n17803# a_65117_n17803# 0.0284f
C3597 a_110225_n1530# VDD 0.150485f
C3598 a_73268_n28415# VDD 0.042519f
C3599 a_93969_n14095# a_93969_n15000# 0.005903f
C3600 a_43817_n27257# a_43817_n28415# 0.004047f
C3601 a_32353_n18698# I1U 0.002649f
C3602 a_33265_n3548# a_31831_n4445# 1.57e-19
C3603 a_35781_n2651# a_34347_n3548# 0.018216f
C3604 a_32913_n3548# a_32353_n3548# 0.0284f
C3605 a_57977_n3550# a_56895_n4447# 5.37e-19
C3606 a_57417_n2653# a_57417_n3550# 0.005987f
C3607 a_58851_n2653# a_59763_n3550# 5.43e-19
C3608 a_93131_n13190# IBPOUT 0.054237f
C3609 a_45445_n12419# a_48313_n13316# 5.37e-19
C3610 a_44885_n12419# a_44885_n13316# 0.005987f
C3611 a_44363_n13316# a_45445_n14213# 5.37e-19
C3612 a_81735_n14095# VDD 0.121415f
C3613 a_105933_n3340# a_105933_n4245# 0.005903f
C3614 a_94537_n19525# a_94537_n20430# 0.005903f
C3615 a_55601_n28415# a_55601_n29181# 0.00778f
C3616 a_33265_n8033# a_33787_n7136# 0.0284f
C3617 a_58329_n8035# a_56895_n8932# 1.57e-19
C3618 a_57977_n8035# a_57417_n8035# 0.0284f
C3619 a_60109_13546# VDD 0.029536f
C3620 a_105933_n8770# a_106501_n8770# 0.027101f
C3621 a_86903_n15905# VDD 0.393432f
C3622 a_42442_n33224# VDD 0.029536f
C3623 a_100235_n15000# a_100235_n15905# 0.005903f
C3624 a_32353_n8930# I1U 0.002649f
C3625 a_101350_n35156# a_101350_n36322# 0.004007f
C3626 a_39531_n3548# a_40965_n3548# 0.005986f
C3627 a_40613_n2651# a_40613_n3548# 0.01664f
C3628 a_79182_n36322# VCM 0.001273f
C3629 a_85089_13546# VDD 0.05845f
C3630 a_66029_n3550# a_66551_n2653# 0.0284f
C3631 a_87433_n1530# a_88271_n1530# 0.027101f
C3632 a_93131_n15905# VDD 0.113729f
C3633 a_111631_n4245# a_113037_n6960# 0.002302f
C3634 a_100235_n20430# a_100803_n20430# 0.027101f
C3635 a_73302_n35156# VDD 0.009062f
C3636 a_43817_5639# a_43817_4481# 0.004047f
C3637 a_39179_n8033# a_39531_n8033# 0.210644f
C3638 a_40613_n7136# a_40613_n8930# 0.011408f
C3639 a_42047_n7136# a_40965_n8033# 5.37e-19
C3640 a_41487_n6239# a_41487_n7136# 0.005987f
C3641 a_64595_n8035# a_65117_n8035# 0.0284f
C3642 a_64243_n8035# a_65677_n8932# 1.57e-19
C3643 a_67111_n7138# a_67111_n8932# 0.005987f
C3644 a_107230_12380# VDD 0.009062f
C3645 a_50629_n17803# a_51151_n16906# 0.0284f
C3646 a_53145_n17803# a_54019_n16906# 0.005903f
C3647 a_82573_n6960# VDD 0.012916f
C3648 a_86903_n7865# a_88271_n6960# 2.31e-19
C3649 a_105933_n15905# a_107339_n18620# 0.002302f
C3650 a_108636_n34390# VDD 0.009062f
C3651 a_48313_n2651# a_47753_n2651# 0.0284f
C3652 a_35221_n12419# a_35781_n13316# 0.0284f
C3653 a_56895_n13318# a_57977_n14215# 5.37e-19
C3654 a_57417_n12421# a_57417_n13318# 0.005987f
C3655 a_88839_n7865# VDD 0.016281f
C3656 a_93131_n2435# a_93969_n2435# 0.027101f
C3657 a_95105_n1530# a_95105_n2435# 0.024773f
C3658 a_92601_n5150# a_93969_n3340# 0.002134f
C3659 a_81735_n17715# a_81735_n18620# 0.006141f
C3660 a_105365_n21335# a_105933_n21335# 0.027101f
C3661 a_77747_7563# a_77747_6405# 0.004047f
C3662 a_46879_n7136# a_46879_n8930# 0.011408f
C3663 a_45445_n8033# a_45797_n8033# 0.210644f
C3664 a_47753_n6239# a_47753_n7136# 0.005987f
C3665 a_48313_n7136# a_47231_n8033# 5.37e-19
C3666 a_59763_n16906# a_59763_n18700# 0.0089f
C3667 a_94537_n8770# VDD 0.016652f
C3668 a_95105_n6960# a_95105_n7865# 0.024773f
C3669 VDD IN_POS 6.65925f
C3670 a_88271_n13190# a_88271_n14095# 0.005903f
C3671 a_111063_n18620# VDD 0.023101f
C3672 a_65677_n14215# IBNOUT 0.0169f
C3673 a_66016_11614# a_66016_10448# 0.004007f
C3674 a_54579_n2653# a_54019_n2653# 0.0284f
C3675 a_38097_n13316# a_39531_n14213# 1.57e-19
C3676 a_40613_n13316# a_41487_n12419# 5.43e-19
C3677 a_65677_n13318# a_67111_n13318# 0.014106f
C3678 a_99667_n9675# VDD 0.02546f
C3679 a_98829_n3340# a_99667_n3340# 0.027101f
C3680 a_98299_n5150# a_98299_n9675# 0.032645f
C3681 a_101641_n3340# a_100803_n3340# 0.028522f
C3682 a_88271_n18620# a_88271_n19525# 0.005903f
C3683 a_108602_6405# a_108602_5639# 0.00778f
C3684 a_77747_n28415# VCM 0.003538f
C3685 a_53145_n7138# a_54019_n8035# 8.45e-19
C3686 a_52063_n8035# a_52585_n7138# 0.0284f
C3687 a_40613_n17801# a_41487_n16904# 4.96e-19
C3688 a_63161_n17803# a_64243_n18700# 5.37e-19
C3689 a_63683_n16906# a_63683_n17803# 0.005987f
C3690 a_66551_n16906# a_67111_n17803# 0.0284f
C3691 a_65677_n17803# a_64595_n18700# 0.011365f
C3692 a_109695_n5150# VDD 1.40049f
C3693 a_100235_n7865# a_100235_n8770# 0.005903f
C3694 a_71864_n28415# VDD 0.042519f
C3695 a_95105_n14095# a_95943_n15000# 0.028522f
C3696 a_31831_n19595# I1U 1.79e-35
C3697 a_32353_n2651# a_32353_n3548# 0.005987f
C3698 a_33787_n2651# a_34699_n3548# 5.43e-19
C3699 a_32913_n3548# a_31831_n4445# 5.37e-19
C3700 a_58329_n3550# a_59763_n3550# 0.014106f
C3701 a_59411_n2653# a_59411_n3550# 0.011408f
C3702 a_46319_n12419# a_46879_n13316# 0.0284f
C3703 a_45445_n12419# a_47753_n12419# 0.0284f
C3704 a_92601_n16810# IBPOUT 0.531205f
C3705 a_44363_n13316# a_44885_n13316# 0.0284f
C3706 a_85089_n35156# a_85089_n36322# 0.004007f
C3707 a_35781_n7136# a_35221_n7136# 0.0284f
C3708 a_57417_n7138# a_57417_n8035# 0.005987f
C3709 a_57977_n8035# a_56895_n8932# 5.37e-19
C3710 a_83709_n4245# a_84547_n6960# 0.032618f
C3711 a_90245_n15000# VDD 0.392932f
C3712 w_27790_n38888# I1U 0.020177f
C3713 a_104527_n8770# a_104527_n9675# 0.024773f
C3714 a_37968_n36322# VDD 0.021314f
C3715 a_39531_n3548# a_40053_n2651# 0.0284f
C3716 a_77776_n36322# VCM 0.003755f
C3717 a_83683_13546# VDD 0.073724f
C3718 a_64243_n3550# a_63683_n3550# 0.0284f
C3719 a_64595_n3550# a_63161_n4447# 1.57e-19
C3720 a_86903_n5150# a_88271_n1530# 7.4e-19
C3721 a_111631_n4245# a_112199_n4245# 0.027101f
C3722 a_95105_n15000# VDD 0.180258f
C3723 a_110225_n4245# a_110225_n6055# 0.006141f
C3724 a_98829_n20430# a_98829_n21335# 0.024773f
C3725 a_71896_n35156# VDD 0.009062f
C3726 a_32088_13546# a_32088_12380# 0.004007f
C3727 a_38097_n7136# a_38097_n8930# 0.005987f
C3728 a_66029_n8035# a_66551_n7138# 0.0284f
C3729 a_54019_n16009# a_54019_n16906# 0.005987f
C3730 a_81735_n6960# VDD 0.137705f
C3731 a_86903_n7865# a_87433_n6960# 0.028522f
C3732 a_86903_n9675# a_88271_n6960# 0.002134f
C3733 a_98829_n17715# VDD 0.41764f
C3734 a_107230_n34390# VDD 0.009062f
C3735 a_104527_n15905# a_104527_n17715# 0.006141f
C3736 a_105933_n15905# a_106501_n15905# 0.027101f
C3737 a_60080_6405# a_60080_5639# 0.00778f
C3738 a_45445_n3548# a_45797_n3548# 0.210644f
C3739 a_47753_n1754# a_47753_n2651# 0.005987f
C3740 a_48313_n2651# a_47231_n3548# 5.37e-19
C3741 a_34347_n13316# a_35781_n13316# 0.014106f
C3742 a_32913_n12419# a_32913_n14213# 0.006457f
C3743 a_58851_n12421# a_59411_n13318# 0.0284f
C3744 a_56895_n13318# a_57417_n13318# 0.0284f
C3745 a_88271_n7865# VDD 0.016281f
C3746 a_92601_n5150# a_93131_n3340# 0.012586f
C3747 a_103997_n21335# VDD 0.926275f
C3748 a_106501_n20430# a_106501_n21335# 0.024773f
C3749 a_44363_n7136# a_44363_n8930# 0.005987f
C3750 a_34347_n17801# a_35781_n17801# 0.003256f
C3751 a_35221_n16007# a_35221_n16904# 0.005987f
C3752 a_34699_n16904# a_34699_n18698# 0.009483f
C3753 a_31831_n17801# a_32353_n16904# 0.0284f
C3754 a_59411_n17803# a_60845_n17803# 0.08885f
C3755 a_93969_n8770# VDD 0.016652f
C3756 a_93131_n7865# a_93969_n7865# 0.027101f
C3757 a_65117_n14215# IBNOUT -2.98e-34
C3758 a_110225_n18620# VDD 0.113729f
C3759 a_113037_n18620# a_113037_n17715# 0.088786f
C3760 a_54019_n1756# a_54019_n2653# 0.005987f
C3761 a_54579_n2653# a_53497_n3550# 5.37e-19
C3762 a_51711_n3550# a_52063_n3550# 0.210644f
C3763 a_39179_n12419# a_42047_n13316# 5.37e-19
C3764 a_114485_7563# VDD 0.002225f
C3765 a_38097_n13316# a_39179_n14213# 5.37e-19
C3766 a_38619_n12419# a_38619_n13316# 0.005987f
C3767 a_63161_n13318# a_64595_n14215# 1.57e-19
C3768 a_65677_n13318# a_66551_n12421# 5.43e-19
C3769 a_98829_n9675# VDD 0.150485f
C3770 a_98299_n4245# a_99667_n3340# 2.31e-19
C3771 a_100803_n2435# a_100803_n3340# 0.024773f
C3772 a_101641_n3340# a_100235_n3340# 2.31e-19
C3773 a_88839_n18620# a_89407_n18620# 0.027101f
C3774 a_79182_12380# a_79182_11614# 0.00778f
C3775 a_53145_n7138# a_53145_n8932# 0.01664f
C3776 a_54579_n7138# a_54019_n7138# 0.0284f
C3777 a_63161_n17803# a_63683_n17803# 0.0284f
C3778 a_65677_n17803# a_64243_n18700# 9.78e-20
C3779 a_106501_n9675# VDD 0.150485f
C3780 a_94537_n14095# a_95943_n15000# 2.31e-19
C3781 a_93131_n14095# a_93131_n15000# 0.024773f
C3782 a_42413_n27257# a_42413_n28415# 0.004047f
C3783 a_33265_n3548# a_34699_n3548# 0.005986f
C3784 a_34347_n2651# a_34347_n3548# 0.01664f
C3785 a_32088_10448# VDD 0.05812f
C3786 a_58329_n3550# a_58851_n2653# 0.0284f
C3787 a_45445_n12419# a_46879_n13316# 0.054819f
C3788 a_83709_n13190# VDD 0.150485f
C3789 a_107339_n3340# a_107339_n6960# 0.011861f
C3790 a_105365_n3340# a_105365_n4245# 0.005903f
C3791 a_95105_n19525# a_95943_n20430# 0.028522f
C3792 a_93969_n19525# a_93969_n20430# 0.005903f
C3793 a_54197_n28415# a_54197_n29181# 0.00778f
C3794 a_35221_n6239# a_35221_n7136# 0.005987f
C3795 a_35781_n7136# a_34699_n8033# 5.37e-19
C3796 a_32913_n8033# a_33265_n8033# 0.210644f
C3797 a_34347_n7136# a_34347_n8930# 0.011408f
C3798 a_55635_10448# VDD 0.021515f
C3799 a_58329_n8035# a_59763_n8035# 0.005986f
C3800 a_59411_n7138# a_60845_n8932# 0.018216f
C3801 a_46879_n17801# a_47753_n16007# 0.030444f
C3802 a_44885_n16007# a_44885_n16904# 0.005987f
C3803 a_45445_n16904# a_45445_n18698# 0.009307f
C3804 a_83141_n4245# a_84547_n6960# 7.35e-19
C3805 a_89407_n14095# VDD 0.121415f
C3806 a_105365_n8770# a_105933_n8770# 0.027101f
C3807 a_36562_n36322# VDD 0.021314f
C3808 a_99667_n15000# a_99667_n15905# 0.005903f
C3809 a_101641_n15000# a_101641_n18620# 0.011861f
C3810 a_102756_n34390# a_102756_n35156# 0.00778f
C3811 a_42047_n2651# a_41487_n2651# 0.0284f
C3812 a_65117_n2653# a_66029_n3550# 5.43e-19
C3813 a_63683_n2653# a_63683_n3550# 0.005987f
C3814 a_64243_n3550# a_63161_n4447# 5.37e-19
C3815 a_86903_n5150# a_87433_n1530# 0.032766f
C3816 a_94537_n15000# VDD 0.02234f
C3817 a_73302_n34390# VDD 0.009062f
C3818 a_99667_n20430# a_100235_n20430# 0.027101f
C3819 a_42413_5639# a_42413_4481# 0.004047f
C3820 a_38619_n7136# a_39179_n8033# 0.0284f
C3821 a_108636_13546# VDD 0.021314f
C3822 a_64243_n8035# a_63683_n8035# 0.0284f
C3823 a_64595_n8035# a_63161_n8932# 1.57e-19
C3824 a_51711_n16906# a_51711_n18700# 0.008933f
C3825 a_81205_n7865# VDD 0.399575f
C3826 a_86903_n9675# a_87433_n6960# 0.012586f
C3827 a_90245_n6960# a_89407_n6960# 0.042385f
C3828 a_101641_n18620# VDD 1.15407f
C3829 a_111631_n9675# a_112199_n9675# 0.027101f
C3830 a_108636_n33224# VDD 0.021515f
C3831 a_96818_n27257# a_96818_n28415# 0.004047f
C3832 a_46879_n2651# a_47753_n2651# 5.43e-19
C3833 a_34347_n13316# a_35221_n12419# 5.43e-19
C3834 a_31831_n13316# a_33265_n14213# 1.57e-19
C3835 a_87433_n7865# VDD 0.121044f
C3836 a_94537_n1530# a_94537_n2435# 0.005903f
C3837 a_92601_n5150# a_92601_n4245# 0.086339f
C3838 a_81735_n17715# a_81205_n21335# 0.03483f
C3839 a_73268_n30339# I1N 0.003619f
C3840 a_107339_n17715# VDD 0.472471f
C3841 a_104527_n21335# a_105365_n21335# 0.027101f
C3842 a_108602_n28415# a_108602_n29181# 0.00778f
C3843 a_44885_n7136# a_45445_n8033# 0.0284f
C3844 a_34347_n17801# a_35221_n16904# 4.96e-19
C3845 a_56895_n17803# a_57417_n16906# 0.0284f
C3846 a_59411_n17803# a_60285_n16906# 0.005903f
C3847 a_93131_n8770# VDD 0.149203f
C3848 a_94537_n6960# a_94537_n7865# 0.005903f
C3849 a_92601_n9675# a_93969_n8770# 0.002134f
C3850 a_86903_n16810# a_88271_n14095# 0.002134f
C3851 a_87433_n13190# a_87433_n14095# 0.024773f
C3852 a_63683_n14215# IBNOUT 0.004735f
C3853 a_88839_n13190# a_89407_n13190# 0.027101f
C3854 a_109695_n19525# VDD 0.393432f
C3855 a_67422_12380# a_67422_11614# 0.00778f
C3856 a_53145_n2653# a_54019_n2653# 5.43e-19
C3857 a_38097_n13316# a_38619_n13316# 0.0284f
C3858 a_40053_n12419# a_40613_n13316# 0.0284f
C3859 a_39179_n12419# a_41487_n12419# 0.0284f
C3860 a_63161_n13318# a_64243_n14215# 5.37e-19
C3861 a_63683_n12421# a_63683_n13318# 0.005987f
C3862 a_100803_n8770# VDD 0.121415f
C3863 a_98299_n4245# a_98829_n3340# 0.028522f
C3864 a_87433_n18620# a_87433_n19525# 0.024773f
C3865 a_86903_n19525# a_88271_n19525# 2.31e-19
C3866 a_107198_6405# a_107198_5639# 0.00778f
C3867 a_54579_n7138# a_53497_n8035# 5.37e-19
C3868 a_51711_n8035# a_52063_n8035# 0.210644f
C3869 a_54019_n6241# a_54019_n7138# 0.005987f
C3870 a_66029_n16906# a_66029_n18700# 0.0089f
C3871 a_105933_n9675# VDD 0.02546f
C3872 a_99667_n7865# a_99667_n8770# 0.005903f
C3873 a_94537_n14095# a_95105_n14095# 0.027101f
C3874 a_92601_n16810# a_93969_n15905# 0.002134f
C3875 a_90969_12380# a_90969_11614# 0.00778f
C3876 a_33265_n3548# a_33787_n2651# 0.0284f
C3877 a_30682_10448# VDD 0.073394f
C3878 a_60845_n2653# a_60285_n2653# 0.0284f
C3879 a_45445_n12419# a_46319_n12419# 0.001405f
C3880 a_83141_n13190# VDD 0.02546f
C3881 a_105933_n3340# a_106501_n3340# 0.027101f
C3882 a_94537_n19525# a_95943_n20430# 2.31e-19
C3883 a_83683_n35156# a_83683_n36322# 0.004007f
C3884 a_31831_n7136# a_31831_n8930# 0.005987f
C3885 a_54229_10448# VDD 0.021515f
C3886 a_59411_n7138# a_60285_n8035# 8.45e-19
C3887 a_58329_n8035# a_58851_n7138# 0.0284f
C3888 a_47231_n16904# a_48313_n17801# 0.002917f
C3889 a_81735_n4245# a_81735_n6055# 0.006141f
C3890 a_83141_n4245# a_83709_n4245# 0.027101f
C3891 a_88839_n14095# VDD 0.016652f
C3892 a_37968_n35156# VDD 0.009062f
C3893 a_100235_n15000# a_100803_n15000# 0.027101f
C3894 a_66058_n29181# a_66058_n30339# 0.004047f
C3895 a_30377_18342# a_31699_17542# 0.009898f
C3896 a_41487_n1754# a_41487_n2651# 0.005987f
C3897 a_42047_n2651# a_40965_n3548# 5.37e-19
C3898 a_39179_n3548# a_39531_n3548# 0.210644f
C3899 a_77776_n35156# VCM 0.002508f
C3900 a_64595_n3550# a_66029_n3550# 0.014106f
C3901 a_65677_n2653# a_65677_n3550# 0.011408f
C3902 a_93969_n15000# VDD 0.016281f
C3903 a_111063_n4245# a_111631_n4245# 0.027101f
C3904 a_71896_n34390# VDD 0.009062f
C3905 a_71896_13546# OUT 0.001027f
C3906 a_30682_13546# a_30682_12380# 0.004007f
C3907 a_64243_n8035# a_63161_n8932# 5.37e-19
C3908 a_63683_n7138# a_63683_n8035# 0.005987f
C3909 a_51151_n16009# a_51151_n16906# 0.005987f
C3910 a_53497_n16906# a_54579_n17803# 0.001641f
C3911 a_90245_n6960# a_88839_n6960# 0.002302f
C3912 a_86903_n9675# a_86903_n7865# 0.086469f
C3913 a_81205_n9675# VDD 1.03081f
C3914 a_100803_n15905# VDD 0.112244f
C3915 a_105365_n15905# a_105933_n15905# 0.027101f
C3916 a_107230_n33224# VDD 0.021515f
C3917 a_61484_7563# a_61484_6405# 0.004047f
C3918 a_44885_n2651# a_45445_n3548# 0.0284f
C3919 a_46879_n2651# a_47231_n3548# 0.053799f
C3920 a_32913_n12419# a_35781_n13316# 5.37e-19
C3921 a_32353_n12419# a_32353_n13316# 0.005987f
C3922 a_31831_n13316# a_32913_n14213# 5.37e-19
C3923 a_89407_n6960# VDD 0.112244f
C3924 a_87433_n4245# IN_POS 0.00603f
C3925 a_105933_n20430# a_105933_n21335# 0.005903f
C3926 a_60285_n16009# a_60285_n16906# 0.005987f
C3927 a_95943_n8770# VDD 0.399226f
C3928 a_92601_n9675# a_93131_n8770# 0.012586f
C3929 a_63161_n15112# IBNOUT 0.001834f
C3930 a_86903_n16810# a_87433_n14095# 0.012586f
C3931 a_53145_n2653# a_53497_n3550# 0.053799f
C3932 a_51151_n2653# a_51711_n3550# 0.0284f
C3933 a_39179_n12419# a_40613_n13316# 0.054819f
C3934 a_63161_n13318# a_63683_n13318# 0.0284f
C3935 a_65117_n12421# a_65677_n13318# 0.0284f
C3936 a_100235_n8770# VDD 0.016652f
C3937 a_100235_n2435# a_100235_n3340# 0.005903f
C3938 a_98299_n5150# a_98829_n6055# 0.03483f
C3939 a_86903_n21335# a_88271_n19525# 0.002134f
C3940 a_90245_n18620# a_90245_n20430# 0.011861f
C3941 a_86903_n19525# a_87433_n19525# 0.028522f
C3942 a_88271_n18620# a_88839_n18620# 0.027101f
C3943 a_77776_12380# a_77776_11614# 0.00778f
C3944 a_77747_n27257# VCM 0.003538f
C3945 a_50629_n7138# a_50629_n8932# 0.005987f
C3946 a_39179_n16904# a_39179_n18698# 0.009307f
C3947 a_40613_n17801# a_41487_n16007# 0.030444f
C3948 a_38619_n16007# a_38619_n16904# 0.005987f
C3949 a_65677_n17803# a_67111_n17803# 0.08885f
C3950 a_105365_n9675# VDD 0.02546f
C3951 a_100803_n7865# a_101641_n8770# 0.028522f
C3952 a_92601_n16810# a_93131_n15905# 0.012586f
C3953 a_67422_n35156# a_67422_n36322# 0.004007f
C3954 a_35781_n2651# a_35221_n2651# 0.0284f
C3955 a_57977_n3550# a_58329_n3550# 0.210644f
C3956 a_60845_n2653# a_59763_n3550# 5.37e-19
C3957 a_60285_n1756# a_60285_n2653# 0.005987f
C3958 a_32088_11614# VDD 0.046892f
C3959 a_82573_n13190# VDD 0.02546f
C3960 a_104527_n3340# a_104527_n4245# 0.024773f
C3961 a_103997_n4245# a_105365_n4245# 2.31e-19
C3962 a_93131_n19525# a_93131_n20430# 0.024773f
C3963 a_94537_n19525# a_95105_n19525# 0.027101f
C3964 a_102756_11614# a_102756_10448# 0.004007f
C3965 a_32353_n7136# a_32913_n8033# 0.0284f
C3966 a_55635_11614# VDD 0.009062f
C3967 a_59411_n7138# a_59411_n8932# 0.01664f
C3968 a_60845_n7138# a_60285_n7138# 0.0284f
C3969 a_47231_n16904# a_47753_n16904# 0.035574f
C3970 a_88271_n14095# VDD 0.016652f
C3971 a_107339_n8770# a_106501_n8770# 0.028522f
C3972 a_104527_n8770# a_105365_n8770# 0.027101f
C3973 a_98829_n15000# a_98829_n15905# 0.024773f
C3974 a_98299_n15905# a_99667_n15905# 2.31e-19
C3975 a_36562_n35156# VDD 0.009062f
C3976 a_31699_19142# a_31699_17542# 0.007227f
C3977 a_101350_n34390# a_101350_n35156# 0.00778f
C3978 a_40613_n2651# a_41487_n2651# 5.43e-19
C3979 a_79182_10448# VDD 0.021515f
C3980 a_64595_n3550# a_65117_n2653# 0.0284f
C3981 a_93131_n15000# VDD 0.121044f
C3982 a_112199_n3340# a_112199_n4245# 0.024773f
C3983 a_101641_n20430# a_100803_n20430# 0.028522f
C3984 a_98829_n20430# a_99667_n20430# 0.027101f
C3985 a_43817_6405# a_43817_5639# 0.00778f
C3986 a_40613_n7136# a_41487_n7136# 0.004425f
C3987 a_65677_n7138# a_67111_n8932# 0.018216f
C3988 a_64595_n8035# a_66029_n8035# 0.005986f
C3989 a_54019_n16009# a_53145_n17803# 0.034652f
C3990 a_53497_n16906# a_54019_n16906# 0.034714f
C3991 a_84547_n6055# VDD 0.472471f
C3992 a_87433_n6055# a_87433_n6960# 0.006141f
C3993 a_100235_n15905# VDD 0.023105f
C3994 a_111063_n9675# a_111631_n9675# 0.027101f
C3995 a_84547_n3340# IN_POS 0.004986f
C3996 a_102756_n36322# VDD 0.05845f
C3997 a_106501_n15000# a_106501_n15905# 0.024773f
C3998 a_42442_13546# a_42442_12380# 0.004007f
C3999 a_95414_n27257# a_95414_n28415# 0.004047f
C4000 a_46879_n2651# a_46319_n2651# 0.0284f
C4001 w_27790_n38888# I1N 0.020706f
C4002 a_31831_n13316# a_32353_n13316# 0.0284f
C4003 a_32913_n12419# a_35221_n12419# 0.0284f
C4004 a_33787_n12419# a_34347_n13316# 0.0284f
C4005 a_88839_n6960# VDD 0.023105f
C4006 a_93969_n1530# a_93969_n2435# 0.005903f
C4007 a_104527_n17715# VDD 0.41764f
C4008 a_73268_n29181# I1N 0.002701f
C4009 a_84547_n18620# a_84547_n17715# 0.088786f
C4010 a_107198_n28415# a_107198_n29181# 0.00778f
C4011 a_46879_n7136# a_47753_n7136# 0.004425f
C4012 a_57977_n16906# a_57977_n18700# 0.008933f
C4013 a_93969_n6960# a_93969_n7865# 0.005903f
C4014 a_95105_n7865# VDD 0.121044f
C4015 a_109695_n21335# VDD 1.27413f
C4016 a_88271_n13190# a_88839_n13190# 0.027101f
C4017 a_66016_12380# a_66016_11614# 0.00778f
C4018 a_53145_n2653# a_52585_n2653# 0.0284f
C4019 a_39179_n12419# a_40053_n12419# 0.001405f
C4020 a_99667_n8770# VDD 0.016652f
C4021 a_86903_n21335# a_87433_n19525# 0.012586f
C4022 a_111631_n21335# a_112199_n21335# 0.027101f
C4023 a_51151_n7138# a_51711_n8035# 0.0284f
C4024 a_40965_n16904# a_42047_n17801# 0.002917f
C4025 a_63161_n17803# a_63683_n16906# 0.0284f
C4026 a_65677_n17803# a_66551_n16906# 0.005903f
C4027 a_100235_n7865# a_101641_n8770# 2.31e-19
C4028 a_104527_n9675# VDD 0.150485f
C4029 a_98829_n7865# a_98829_n8770# 0.024773f
C4030 a_93969_n14095# a_94537_n14095# 0.027101f
C4031 a_73302_n36322# I1N 0.002533f
C4032 a_89563_12380# a_89563_11614# 0.00778f
C4033 a_32913_n3548# a_33265_n3548# 0.210644f
C4034 a_35781_n2651# a_34699_n3548# 5.37e-19
C4035 a_35221_n1754# a_35221_n2651# 0.005987f
C4036 a_59411_n2653# a_60285_n2653# 5.43e-19
C4037 a_30682_11614# VDD 0.062166f
C4038 a_44885_n12419# a_45445_n12419# 0.0284f
C4039 a_81735_n13190# VDD 0.150485f
C4040 a_105365_n3340# a_105933_n3340# 0.027101f
C4041 a_103997_n4245# a_104527_n4245# 0.028522f
C4042 a_92601_n21335# a_93969_n21335# 0.002563f
C4043 a_85089_n34390# a_85089_n35156# 0.00778f
C4044 a_60285_n6241# a_60285_n7138# 0.005987f
C4045 a_60845_n7138# a_59763_n8035# 5.37e-19
C4046 a_57977_n8035# a_58329_n8035# 0.210644f
C4047 a_54229_11614# VDD 0.009062f
C4048 a_82573_n4245# a_83141_n4245# 0.027101f
C4049 a_87433_n14095# VDD 0.121415f
C4050 a_106501_n7865# a_106501_n8770# 0.024773f
C4051 a_107339_n8770# a_105933_n8770# 2.31e-19
C4052 a_98299_n15905# a_98829_n15905# 0.028522f
C4053 a_99667_n15000# a_100235_n15000# 0.027101f
C4054 a_32353_n8033# I1U 0.002649f
C4055 a_37968_n34390# VDD 0.009062f
C4056 a_31699_19142# a_30377_18342# 0.009898f
C4057 a_67462_n28415# a_67462_n29181# 0.00778f
C4058 a_38619_n2651# a_39179_n3548# 0.0284f
C4059 a_40613_n2651# a_40965_n3548# 0.053799f
C4060 a_77776_10448# VDD 0.029536f
C4061 a_67111_n2653# a_66551_n2653# 0.0284f
C4062 a_77776_n34390# VCM 0.002508f
C4063 a_50629_n13318# a_51151_n12421# 0.0284f
C4064 a_92601_n15905# VDD 0.393432f
C4065 a_32088_10448# I1U 0.003282f
C4066 a_110225_n4245# a_111063_n4245# 0.027101f
C4067 a_100803_n19525# a_100803_n20430# 0.024773f
C4068 a_101641_n20430# a_100235_n20430# 2.31e-19
C4069 a_73302_n33224# VDD 0.021515f
C4070 a_38097_n7136# a_39531_n8033# 1.57e-19
C4071 a_40613_n7136# a_40965_n8033# 0.062551f
C4072 a_64595_n8035# a_65117_n7138# 0.0284f
C4073 a_65677_n7138# a_66551_n8035# 8.45e-19
C4074 a_107230_13546# VDD 0.021314f
C4075 a_81735_n6055# VDD 0.41764f
C4076 a_99667_n15905# VDD 0.012916f
C4077 a_112199_n8770# a_112199_n9675# 0.024773f
C4078 a_104527_n15905# a_105365_n15905# 0.027101f
C4079 a_101350_n36322# VDD 0.073724f
C4080 a_60080_7563# a_60080_6405# 0.004047f
C4081 a_46879_n2651# a_45797_n3548# 5.37e-19
C4082 a_45445_n1754# a_47231_n3548# 0.006457f
C4083 a_46319_n1754# a_46319_n2651# 0.005987f
C4084 a_44363_n2651# a_44363_n4445# 0.005987f
C4085 a_32913_n12419# a_34347_n13316# 0.054819f
C4086 a_88271_n6960# VDD 0.012916f
C4087 a_107339_n18620# VDD 1.18674f
C4088 a_105365_n20430# a_105365_n21335# 0.005903f
C4089 a_46879_n7136# a_47231_n8033# 0.062551f
C4090 a_44363_n7136# a_45797_n8033# 1.57e-19
C4091 a_32353_n16007# a_32353_n16904# 0.005987f
C4092 a_32913_n16904# a_32913_n18698# 0.009307f
C4093 a_34347_n17801# a_35221_n16007# 0.030444f
C4094 a_57417_n16009# a_57417_n16906# 0.005987f
C4095 a_59763_n16906# a_60845_n17803# 0.001641f
C4096 a_94537_n6960# a_95105_n6960# 0.027101f
C4097 a_94537_n7865# VDD 0.016281f
C4098 a_113037_n17715# VDD 0.472471f
C4099 a_66029_n14215# IBNOUT 0.001202f
C4100 a_112199_n15905# a_113037_n18620# 0.042385f
C4101 a_90935_6405# a_90935_5639# 0.00778f
C4102 a_50629_n2653# a_50629_n4447# 0.005987f
C4103 a_53145_n2653# a_52063_n3550# 5.37e-19
C4104 a_52585_n1756# a_52585_n2653# 0.005987f
C4105 a_108602_5639# VDD 0.042519f
C4106 a_99667_n2435# a_99667_n3340# 0.005903f
C4107 a_98829_n8770# VDD 0.121415f
C4108 a_87433_n18620# a_88271_n18620# 0.027101f
C4109 a_53145_n7138# a_54019_n7138# 0.006769f
C4110 a_40965_n16904# a_41487_n16904# 0.035574f
C4111 a_66551_n16009# a_66551_n16906# 0.005987f
C4112 a_106501_n8770# VDD 0.121415f
C4113 a_100235_n7865# a_100803_n7865# 0.027101f
C4114 IN_NEG VSS 50.44224f
C4115 IN_POS VSS 38.26637f
C4116 VCM VSS 16.767963f
C4117 IBPOUT VSS 11.58886f
C4118 I1N VSS 53.45688f
C4119 IBNOUT VSS 9.23631f
C4120 I1U VSS 33.7696f
C4121 OUT VSS 44.56392f
C4122 VDD VSS 10.164393p
C4123 a_108636_n35156# VSS 0.04473f
C4124 a_107230_n35156# VSS 0.04473f
C4125 a_108636_n34390# VSS 0.04492f
C4126 a_107230_n34390# VSS 0.028915f
C4127 a_108636_n33224# VSS 0.016627f
C4128 a_90969_n35156# VSS 0.04473f
C4129 a_89563_n35156# VSS 0.04473f
C4130 a_90969_n34390# VSS 0.04492f
C4131 a_89563_n34390# VSS 0.028915f
C4132 a_90969_n33224# VSS 0.016627f
C4133 a_73302_n35156# VSS 0.04473f
C4134 a_71896_n35156# VSS 0.04473f
C4135 a_73302_n34390# VSS 0.04492f
C4136 a_71896_n34390# VSS 0.028915f
C4137 a_73302_n33224# VSS 0.016627f
C4138 a_55635_n35156# VSS 0.04473f
C4139 a_54229_n35156# VSS 0.04473f
C4140 a_55635_n34390# VSS 0.04492f
C4141 a_54229_n34390# VSS 0.028915f
C4142 a_55635_n33224# VSS 0.016627f
C4143 a_37968_n35156# VSS 0.04473f
C4144 a_36562_n35156# VSS 0.04473f
C4145 a_37968_n34390# VSS 0.04492f
C4146 a_36562_n34390# VSS 0.028915f
C4147 a_37968_n33224# VSS 0.016627f
C4148 a_114485_n30339# VSS 0.058211f
C4149 a_113081_n30339# VSS 0.070508f
C4150 a_114485_n29181# VSS 0.059789f
C4151 a_113081_n29181# VSS 0.072086f
C4152 a_114485_n28415# VSS 0.04696f
C4153 a_113081_n28415# VSS 0.059257f
C4154 a_114485_n27257# VSS 0.057864f
C4155 a_113081_n27257# VSS 0.070162f
C4156 a_108602_n30339# VSS 0.021386f
C4157 a_107198_n30339# VSS 0.02113f
C4158 a_108602_n29181# VSS 0.009003f
C4159 a_107198_n29181# VSS 0.009003f
C4160 a_108602_n28415# VSS 0.009003f
C4161 a_107198_n28415# VSS 0.009003f
C4162 a_108602_n27257# VSS 0.02113f
C4163 a_107198_n27257# VSS 0.02113f
C4164 a_102796_n30339# VSS 0.024094f
C4165 a_101392_n30339# VSS 0.029168f
C4166 a_102796_n29181# VSS 0.009003f
C4167 a_101392_n29181# VSS 0.017167f
C4168 a_102796_n28415# VSS 0.01202f
C4169 a_101392_n28415# VSS 0.017167f
C4170 a_102796_n27257# VSS 0.02113f
C4171 a_101392_n27257# VSS 0.029168f
C4172 a_96818_n30339# VSS 0.058211f
C4173 a_95414_n30339# VSS 0.070508f
C4174 a_96818_n29181# VSS 0.059789f
C4175 a_95414_n29181# VSS 0.072086f
C4176 a_96818_n28415# VSS 0.04696f
C4177 a_95414_n28415# VSS 0.059257f
C4178 a_96818_n27257# VSS 0.057864f
C4179 a_95414_n27257# VSS 0.070162f
C4180 a_90935_n30339# VSS 0.021386f
C4181 a_89531_n30339# VSS 0.02113f
C4182 a_90935_n29181# VSS 0.009003f
C4183 a_89531_n29181# VSS 0.009003f
C4184 a_90935_n28415# VSS 0.009003f
C4185 a_89531_n28415# VSS 0.009003f
C4186 a_90935_n27257# VSS 0.02113f
C4187 a_89531_n27257# VSS 0.02113f
C4188 a_85129_n30339# VSS 0.024094f
C4189 a_83725_n30339# VSS 0.029168f
C4190 a_85129_n29181# VSS 0.009003f
C4191 a_83725_n29181# VSS 0.017167f
C4192 a_85129_n28415# VSS 0.01202f
C4193 a_83725_n28415# VSS 0.017167f
C4194 a_85129_n27257# VSS 0.02113f
C4195 a_83725_n27257# VSS 0.029168f
C4196 a_79151_n30339# VSS 0.058211f
C4197 a_77747_n30339# VSS 0.070508f
C4198 a_79151_n29181# VSS 0.059789f
C4199 a_77747_n29181# VSS 0.072086f
C4200 a_79151_n28415# VSS 0.04696f
C4201 a_77747_n28415# VSS 0.059257f
C4202 a_79151_n27257# VSS 0.057864f
C4203 a_77747_n27257# VSS 0.070162f
C4204 a_73268_n30339# VSS 0.021386f
C4205 a_71864_n30339# VSS 0.02113f
C4206 a_73268_n29181# VSS 0.009003f
C4207 a_71864_n29181# VSS 0.009003f
C4208 a_73268_n28415# VSS 0.009003f
C4209 a_71864_n28415# VSS 0.009003f
C4210 a_73268_n27257# VSS 0.02113f
C4211 a_71864_n27257# VSS 0.02113f
C4212 a_67462_n30339# VSS 0.024094f
C4213 a_66058_n30339# VSS 0.029168f
C4214 a_67462_n29181# VSS 0.009003f
C4215 a_66058_n29181# VSS 0.017167f
C4216 a_67462_n28415# VSS 0.01202f
C4217 a_66058_n28415# VSS 0.017167f
C4218 a_67462_n27257# VSS 0.02113f
C4219 a_66058_n27257# VSS 0.029168f
C4220 a_61484_n30339# VSS 0.058211f
C4221 a_60080_n30339# VSS 0.070508f
C4222 a_61484_n29181# VSS 0.059789f
C4223 a_60080_n29181# VSS 0.072086f
C4224 a_61484_n28415# VSS 0.04696f
C4225 a_60080_n28415# VSS 0.059257f
C4226 a_61484_n27257# VSS 0.057864f
C4227 a_60080_n27257# VSS 0.070162f
C4228 a_55601_n30339# VSS 0.021386f
C4229 a_54197_n30339# VSS 0.02113f
C4230 a_55601_n29181# VSS 0.009003f
C4231 a_54197_n29181# VSS 0.009003f
C4232 a_55601_n28415# VSS 0.009003f
C4233 a_54197_n28415# VSS 0.009003f
C4234 a_55601_n27257# VSS 0.02113f
C4235 a_54197_n27257# VSS 0.02113f
C4236 a_49795_n30339# VSS 0.024094f
C4237 a_48391_n30339# VSS 0.029168f
C4238 a_49795_n29181# VSS 0.009003f
C4239 a_48391_n29181# VSS 0.017167f
C4240 a_49795_n28415# VSS 0.01202f
C4241 a_48391_n28415# VSS 0.017167f
C4242 a_49795_n27257# VSS 0.02113f
C4243 a_48391_n27257# VSS 0.029168f
C4244 a_43817_n30339# VSS 0.058211f
C4245 a_42413_n30339# VSS 0.070508f
C4246 a_43817_n29181# VSS 0.059789f
C4247 a_42413_n29181# VSS 0.072086f
C4248 a_43817_n28415# VSS 0.04696f
C4249 a_42413_n28415# VSS 0.059257f
C4250 a_43817_n27257# VSS 0.057864f
C4251 a_42413_n27257# VSS 0.070162f
C4252 a_37934_n30339# VSS 0.021386f
C4253 a_36530_n30339# VSS 0.02113f
C4254 a_37934_n29181# VSS 0.009003f
C4255 a_36530_n29181# VSS 0.009003f
C4256 a_37934_n28415# VSS 0.009003f
C4257 a_36530_n28415# VSS 0.009003f
C4258 a_37934_n27257# VSS 0.02113f
C4259 a_36530_n27257# VSS 0.02113f
C4260 a_32128_n30339# VSS 0.024094f
C4261 a_30724_n30339# VSS 0.029168f
C4262 a_32128_n29181# VSS 0.009003f
C4263 a_30724_n29181# VSS 0.017167f
C4264 a_32128_n28415# VSS 0.01202f
C4265 a_30724_n28415# VSS 0.017167f
C4266 a_32128_n27257# VSS 0.02113f
C4267 a_30724_n27257# VSS 0.029168f
C4268 a_113037_n20430# VSS 0.012478f
C4269 a_110225_n18620# VSS 0.001741f
C4270 a_109695_n19525# VSS 0.012478f
C4271 a_109695_n21335# VSS 0.246948f
C4272 a_110225_n17715# VSS 2.3e-25
C4273 a_113037_n18620# VSS 0.233537f
C4274 a_110225_n15905# VSS 0.001741f
C4275 a_109695_n15905# VSS 0.012478f
C4276 a_113037_n15000# VSS 0.012478f
C4277 a_109695_n16810# VSS 0.265878f
C4278 a_107339_n20430# VSS 0.012478f
C4279 a_104527_n18620# VSS 0.001741f
C4280 a_103997_n19525# VSS 0.012478f
C4281 a_103997_n21335# VSS 0.059722f
C4282 a_104527_n17715# VSS 2.3e-25
C4283 a_107339_n18620# VSS 0.233537f
C4284 a_104527_n15905# VSS 0.001741f
C4285 a_103997_n15905# VSS 0.012478f
C4286 a_107339_n15000# VSS 0.012478f
C4287 a_103997_n16810# VSS 0.059409f
C4288 a_101641_n20430# VSS 0.012478f
C4289 a_98829_n18620# VSS 0.001741f
C4290 a_98299_n19525# VSS 0.012478f
C4291 a_98299_n21335# VSS 0.059721f
C4292 a_98829_n17715# VSS 2.3e-25
C4293 a_101641_n18620# VSS 0.077718f
C4294 a_98829_n15905# VSS 0.001741f
C4295 a_98299_n15905# VSS 0.012478f
C4296 a_101641_n15000# VSS 0.012478f
C4297 a_98299_n16810# VSS 0.059409f
C4298 a_95943_n20430# VSS 0.012478f
C4299 a_93131_n18620# VSS 0.001741f
C4300 a_92601_n19525# VSS 0.012478f
C4301 a_92601_n21335# VSS 0.274655f
C4302 a_93131_n17715# VSS 2.3e-25
C4303 a_95943_n18620# VSS 0.077718f
C4304 a_93131_n15905# VSS 0.001741f
C4305 a_92601_n15905# VSS 0.012478f
C4306 a_95943_n15000# VSS 0.012478f
C4307 a_92601_n16810# VSS 0.255977f
C4308 a_90245_n20430# VSS 0.012478f
C4309 a_87433_n18620# VSS 0.001741f
C4310 a_86903_n19525# VSS 0.012478f
C4311 a_86903_n21335# VSS 0.274655f
C4312 a_87433_n17715# VSS 2.3e-25
C4313 a_90245_n18620# VSS 0.233537f
C4314 a_87433_n15905# VSS 0.001741f
C4315 a_86903_n15905# VSS 0.012478f
C4316 a_90245_n15000# VSS 0.012478f
C4317 a_86903_n16810# VSS 0.255977f
C4318 a_84547_n20430# VSS 0.012478f
C4319 a_81735_n18620# VSS 0.001741f
C4320 a_81205_n19525# VSS 0.012478f
C4321 a_81205_n21335# VSS 0.361326f
C4322 a_81735_n17715# VSS 2.3e-25
C4323 a_84547_n18620# VSS 0.233537f
C4324 a_81735_n15905# VSS 0.001741f
C4325 a_81205_n15905# VSS 0.012478f
C4326 a_84547_n15000# VSS 0.012478f
C4327 a_81205_n16810# VSS 0.341999f
C4328 a_113037_n8770# VSS 0.012478f
C4329 a_110225_n6960# VSS 0.001741f
C4330 a_109695_n7865# VSS 0.012478f
C4331 a_109695_n9675# VSS 0.255977f
C4332 a_110225_n6055# VSS 2.3e-25
C4333 a_113037_n6960# VSS 0.233537f
C4334 a_110225_n4245# VSS 0.001741f
C4335 a_109695_n4245# VSS 0.012478f
C4336 a_113037_n3340# VSS 0.012478f
C4337 a_109695_n5150# VSS 0.274655f
C4338 a_107339_n8770# VSS 0.012478f
C4339 a_104527_n6960# VSS 0.001741f
C4340 a_103997_n7865# VSS 0.012478f
C4341 a_103997_n9675# VSS 0.255977f
C4342 a_104527_n6055# VSS 2.3e-25
C4343 a_107339_n6960# VSS 0.233537f
C4344 a_104527_n4245# VSS 0.001741f
C4345 a_103997_n4245# VSS 0.012478f
C4346 a_107339_n3340# VSS 0.012478f
C4347 a_103997_n5150# VSS 0.274655f
C4348 a_101641_n8770# VSS 0.012478f
C4349 a_98829_n6960# VSS 0.001741f
C4350 a_98299_n7865# VSS 0.012478f
C4351 a_98299_n9675# VSS 0.255977f
C4352 a_98829_n6055# VSS 2.3e-25
C4353 a_101641_n6960# VSS 0.233537f
C4354 a_98829_n4245# VSS 0.001741f
C4355 a_98299_n4245# VSS 0.012478f
C4356 a_101641_n3340# VSS 0.012478f
C4357 a_98299_n5150# VSS 0.274655f
C4358 a_95943_n8770# VSS 0.012478f
C4359 a_93131_n6960# VSS 0.001741f
C4360 a_92601_n7865# VSS 0.012478f
C4361 a_92601_n9675# VSS 0.265878f
C4362 a_93131_n6055# VSS 2.3e-25
C4363 a_95943_n6960# VSS 0.233537f
C4364 a_93131_n4245# VSS 0.001741f
C4365 a_92601_n4245# VSS 0.012478f
C4366 a_95943_n3340# VSS 0.012478f
C4367 a_92601_n5150# VSS 0.264496f
C4368 a_90245_n8770# VSS 0.012478f
C4369 a_87433_n6960# VSS 0.001741f
C4370 a_86903_n7865# VSS 0.012478f
C4371 a_86903_n9675# VSS 0.059409f
C4372 a_87433_n6055# VSS 2.3e-25
C4373 a_90245_n6960# VSS 0.233537f
C4374 a_87433_n4245# VSS 0.001741f
C4375 a_86903_n4245# VSS 0.012478f
C4376 a_90245_n3340# VSS 0.012478f
C4377 a_86903_n5150# VSS 0.059721f
C4378 a_84547_n8770# VSS 0.012478f
C4379 a_81735_n6960# VSS 0.001741f
C4380 a_81205_n7865# VSS 0.012478f
C4381 a_81205_n9675# VSS 0.063176f
C4382 a_81735_n6055# VSS 2.3e-25
C4383 a_84547_n6960# VSS 0.077718f
C4384 a_81735_n4245# VSS 0.001741f
C4385 a_81205_n4245# VSS 0.012478f
C4386 a_84547_n3340# VSS 0.012478f
C4387 a_81205_n5150# VSS 0.059721f
C4388 a_75585_n10973# VSS 0.036472f
C4389 a_72603_n10973# VSS 0.036472f
C4390 a_75585_n10073# VSS 0.02091f
C4391 a_72603_n10073# VSS 0.02091f
C4392 a_75585_n9297# VSS 0.020886f
C4393 a_72603_n9297# VSS 0.02091f
C4394 a_75585_n8397# VSS 0.036472f
C4395 a_72603_n8397# VSS 0.036472f
C4396 a_66551_n19597# VSS 0.025764f
C4397 a_65117_n19597# VSS 0.053627f
C4398 a_64243_n19597# VSS 1.20649f
C4399 a_63683_n19597# VSS 0.025764f
C4400 a_67111_n19597# VSS 0.398427f
C4401 a_66551_n18700# VSS 0.017066f
C4402 a_65677_n19597# VSS 0.225452f
C4403 a_65117_n18700# VSS 0.016529f
C4404 a_63683_n18700# VSS 0.017066f
C4405 a_63161_n19597# VSS 0.412143f
C4406 a_66551_n17803# VSS 0.016697f
C4407 a_66029_n18700# VSS 0.200377f
C4408 a_65117_n17803# VSS 0.023002f
C4409 a_64595_n18700# VSS 0.178599f
C4410 a_64243_n18700# VSS 0.192438f
C4411 a_63683_n17803# VSS 0.016697f
C4412 a_67111_n17803# VSS 0.405499f
C4413 a_66551_n16906# VSS 0.017551f
C4414 a_63683_n16906# VSS 0.017551f
C4415 a_63161_n17803# VSS 0.417122f
C4416 a_65677_n17803# VSS 1.46283f
C4417 a_66551_n16009# VSS 0.018938f
C4418 a_63683_n16009# VSS 0.056084f
C4419 a_66551_n15112# VSS 0.017564f
C4420 a_66029_n16906# VSS 0.550027f
C4421 a_64243_n16906# VSS 0.622493f
C4422 a_63683_n15112# VSS 0.024755f
C4423 a_67111_n15112# VSS 0.405615f
C4424 a_66551_n14215# VSS 0.016697f
C4425 a_65677_n14215# VSS 0.385498f
C4426 a_65117_n14215# VSS 0.023005f
C4427 a_63683_n14215# VSS 0.023888f
C4428 a_63161_n15112# VSS 0.490894f
C4429 a_66551_n13318# VSS 0.017062f
C4430 a_66029_n14215# VSS 0.227033f
C4431 a_65117_n13318# VSS 0.016525f
C4432 a_64595_n14215# VSS 0.175025f
C4433 a_64243_n14215# VSS 0.199765f
C4434 a_63683_n13318# VSS 0.024253f
C4435 a_67111_n13318# VSS 0.398946f
C4436 a_66551_n12421# VSS 0.054141f
C4437 a_65677_n13318# VSS 0.298391f
C4438 a_65117_n12421# VSS 0.025832f
C4439 a_63683_n12421# VSS 0.032931f
C4440 a_63161_n13318# VSS 0.491582f
C4441 a_60285_n19597# VSS 0.025764f
C4442 a_58851_n19597# VSS 0.053627f
C4443 a_57977_n19597# VSS 1.20649f
C4444 a_57417_n19597# VSS 0.025764f
C4445 a_60845_n19597# VSS 0.398427f
C4446 a_60285_n18700# VSS 0.017066f
C4447 a_59411_n19597# VSS 0.225452f
C4448 a_58851_n18700# VSS 0.016529f
C4449 a_57417_n18700# VSS 0.017066f
C4450 a_56895_n19597# VSS 0.412143f
C4451 a_60285_n17803# VSS 0.016697f
C4452 a_59763_n18700# VSS 0.200377f
C4453 a_58851_n17803# VSS 0.023002f
C4454 a_58329_n18700# VSS 0.178599f
C4455 a_57977_n18700# VSS 0.192438f
C4456 a_57417_n17803# VSS 0.016697f
C4457 a_60845_n17803# VSS 0.405499f
C4458 a_60285_n16906# VSS 0.017551f
C4459 a_57417_n16906# VSS 0.017551f
C4460 a_56895_n17803# VSS 0.405047f
C4461 a_59411_n17803# VSS 1.45216f
C4462 a_60285_n16009# VSS 0.018938f
C4463 a_57417_n16009# VSS 0.018938f
C4464 a_60285_n15112# VSS 0.017564f
C4465 a_59763_n16906# VSS 0.550027f
C4466 a_57977_n16906# VSS 0.546597f
C4467 a_57417_n15112# VSS 0.017564f
C4468 a_60845_n15112# VSS 0.405615f
C4469 a_60285_n14215# VSS 0.016697f
C4470 a_59411_n14215# VSS 0.385498f
C4471 a_58851_n14215# VSS 0.023005f
C4472 a_57417_n14215# VSS 0.016697f
C4473 a_56895_n15112# VSS 0.405161f
C4474 a_60285_n13318# VSS 0.017062f
C4475 a_59763_n14215# VSS 0.227033f
C4476 a_58851_n13318# VSS 0.016525f
C4477 a_58329_n14215# VSS 0.174939f
C4478 a_57977_n14215# VSS 0.192438f
C4479 a_57417_n13318# VSS 0.017062f
C4480 a_60845_n13318# VSS 0.398946f
C4481 a_60285_n12421# VSS 0.054141f
C4482 a_59411_n13318# VSS 0.298391f
C4483 a_58851_n12421# VSS 0.025832f
C4484 a_57417_n12421# VSS 0.025741f
C4485 a_56895_n13318# VSS 0.411967f
C4486 a_54019_n19597# VSS 0.025764f
C4487 a_52585_n19597# VSS 0.053627f
C4488 a_51711_n19597# VSS 1.20649f
C4489 a_51151_n19597# VSS 0.025764f
C4490 a_54579_n19597# VSS 0.398427f
C4491 a_54019_n18700# VSS 0.017066f
C4492 a_53145_n19597# VSS 0.225452f
C4493 a_52585_n18700# VSS 0.016529f
C4494 a_51151_n18700# VSS 0.017066f
C4495 a_50629_n19597# VSS 0.412149f
C4496 a_54019_n17803# VSS 0.016697f
C4497 a_53497_n18700# VSS 0.200377f
C4498 a_52585_n17803# VSS 0.023002f
C4499 a_52063_n18700# VSS 0.178599f
C4500 a_51711_n18700# VSS 0.192438f
C4501 a_51151_n17803# VSS 0.016697f
C4502 a_54579_n17803# VSS 0.405499f
C4503 a_54019_n16906# VSS 0.017551f
C4504 a_51151_n16906# VSS 0.017551f
C4505 a_50629_n17803# VSS 0.405053f
C4506 a_53145_n17803# VSS 1.45216f
C4507 a_54019_n16009# VSS 0.018938f
C4508 a_51151_n16009# VSS 0.018938f
C4509 a_54019_n15112# VSS 0.017564f
C4510 a_53497_n16906# VSS 0.550027f
C4511 a_51711_n16906# VSS 0.546597f
C4512 a_51151_n15112# VSS 0.017564f
C4513 a_54579_n15112# VSS 0.405615f
C4514 a_54019_n14215# VSS 0.016697f
C4515 a_53145_n14215# VSS 0.385498f
C4516 a_52585_n14215# VSS 0.023005f
C4517 a_51151_n14215# VSS 0.016697f
C4518 a_50629_n15112# VSS 0.405167f
C4519 a_54019_n13318# VSS 0.017062f
C4520 a_53497_n14215# VSS 0.227033f
C4521 a_52585_n13318# VSS 0.016525f
C4522 a_52063_n14215# VSS 0.174939f
C4523 a_51711_n14215# VSS 0.192438f
C4524 a_51151_n13318# VSS 0.017062f
C4525 a_54579_n13318# VSS 0.398946f
C4526 a_54019_n12421# VSS 0.054141f
C4527 a_53145_n13318# VSS 0.298391f
C4528 a_52585_n12421# VSS 0.025832f
C4529 a_51151_n12421# VSS 0.025741f
C4530 a_50629_n13318# VSS 0.411972f
C4531 a_47753_n19595# VSS 0.054141f
C4532 a_46319_n19595# VSS 0.025832f
C4533 a_44885_n19595# VSS 0.025741f
C4534 a_48313_n19595# VSS 0.398952f
C4535 a_47753_n18698# VSS 0.017062f
C4536 a_46879_n19595# VSS 0.298391f
C4537 a_46319_n18698# VSS 0.016525f
C4538 a_44885_n18698# VSS 0.017062f
C4539 a_44363_n19595# VSS 0.411967f
C4540 a_47753_n17801# VSS 0.016697f
C4541 a_47231_n18698# VSS 0.227033f
C4542 a_46319_n17801# VSS 0.023005f
C4543 a_45797_n18698# VSS 0.174939f
C4544 a_45445_n18698# VSS 0.192438f
C4545 a_44885_n17801# VSS 0.016697f
C4546 a_48313_n17801# VSS 0.40562f
C4547 a_47753_n16904# VSS 0.017564f
C4548 a_44885_n16904# VSS 0.017564f
C4549 a_44363_n17801# VSS 0.405161f
C4550 a_47753_n16007# VSS 0.018938f
C4551 a_46879_n17801# VSS 0.385498f
C4552 a_44885_n16007# VSS 0.018938f
C4553 a_47753_n15110# VSS 0.017551f
C4554 a_47231_n16904# VSS 0.550027f
C4555 a_45445_n16904# VSS 0.546597f
C4556 a_44885_n15110# VSS 0.017551f
C4557 a_48313_n15110# VSS 0.405505f
C4558 a_47753_n14213# VSS 0.016697f
C4559 a_46879_n14213# VSS 1.45219f
C4560 a_46319_n14213# VSS 0.023002f
C4561 a_44885_n14213# VSS 0.016697f
C4562 a_44363_n15110# VSS 0.405047f
C4563 a_47753_n13316# VSS 0.017066f
C4564 a_47231_n14213# VSS 0.200377f
C4565 a_46319_n13316# VSS 0.016529f
C4566 a_45797_n14213# VSS 0.178599f
C4567 a_45445_n14213# VSS 0.192438f
C4568 a_44885_n13316# VSS 0.017066f
C4569 a_48313_n13316# VSS 0.398433f
C4570 a_47753_n12419# VSS 0.025764f
C4571 a_46879_n13316# VSS 0.225452f
C4572 a_46319_n12419# VSS 0.053627f
C4573 a_45445_n12419# VSS 1.14257f
C4574 a_44885_n12419# VSS 0.025764f
C4575 a_44363_n13316# VSS 0.412143f
C4576 a_41487_n19595# VSS 0.054141f
C4577 a_40053_n19595# VSS 0.025832f
C4578 a_38619_n19595# VSS 0.025741f
C4579 a_42047_n19595# VSS 0.398946f
C4580 a_41487_n18698# VSS 0.017062f
C4581 a_40613_n19595# VSS 0.298391f
C4582 a_40053_n18698# VSS 0.016525f
C4583 a_38619_n18698# VSS 0.017062f
C4584 a_38097_n19595# VSS 0.411967f
C4585 a_41487_n17801# VSS 0.016697f
C4586 a_40965_n18698# VSS 0.227033f
C4587 a_40053_n17801# VSS 0.023005f
C4588 a_39531_n18698# VSS 0.174939f
C4589 a_39179_n18698# VSS 0.192438f
C4590 a_38619_n17801# VSS 0.016697f
C4591 a_42047_n17801# VSS 0.405615f
C4592 a_41487_n16904# VSS 0.017564f
C4593 a_38619_n16904# VSS 0.017564f
C4594 a_38097_n17801# VSS 0.405161f
C4595 a_41487_n16007# VSS 0.018938f
C4596 a_40613_n17801# VSS 0.385498f
C4597 a_38619_n16007# VSS 0.018938f
C4598 a_41487_n15110# VSS 0.017551f
C4599 a_40965_n16904# VSS 0.550027f
C4600 a_39179_n16904# VSS 0.497514f
C4601 a_38619_n15110# VSS 0.017551f
C4602 a_42047_n15110# VSS 0.405499f
C4603 a_41487_n14213# VSS 0.016697f
C4604 a_40613_n14213# VSS 1.45216f
C4605 a_40053_n14213# VSS 0.023002f
C4606 a_38619_n14213# VSS 0.016697f
C4607 a_38097_n15110# VSS 0.405047f
C4608 a_41487_n13316# VSS 0.017066f
C4609 a_40965_n14213# VSS 0.200377f
C4610 a_40053_n13316# VSS 0.016529f
C4611 a_39531_n14213# VSS 0.178599f
C4612 a_39179_n14213# VSS 0.192438f
C4613 a_38619_n13316# VSS 0.017066f
C4614 a_42047_n13316# VSS 0.398427f
C4615 a_41487_n12419# VSS 0.025764f
C4616 a_40613_n13316# VSS 0.225452f
C4617 a_40053_n12419# VSS 0.053627f
C4618 a_39179_n12419# VSS 1.10481f
C4619 a_38619_n12419# VSS 0.025764f
C4620 a_38097_n13316# VSS 0.412143f
C4621 a_35221_n19595# VSS 0.054141f
C4622 a_33787_n19595# VSS 0.025832f
C4623 a_32353_n19595# VSS 0.025741f
C4624 a_35781_n19595# VSS 0.398946f
C4625 a_35221_n18698# VSS 0.017062f
C4626 a_34347_n19595# VSS 0.298391f
C4627 a_33787_n18698# VSS 0.016525f
C4628 a_32353_n18698# VSS 0.017062f
C4629 a_31831_n19595# VSS 0.411967f
C4630 a_35221_n17801# VSS 0.016697f
C4631 a_34699_n18698# VSS 0.227033f
C4632 a_33787_n17801# VSS 0.023005f
C4633 a_33265_n18698# VSS 0.174939f
C4634 a_32913_n18698# VSS 0.192438f
C4635 a_32353_n17801# VSS 0.016697f
C4636 a_35781_n17801# VSS 0.405615f
C4637 a_35221_n16904# VSS 0.017564f
C4638 a_32353_n16904# VSS 0.017564f
C4639 a_31831_n17801# VSS 0.405161f
C4640 a_35221_n16007# VSS 0.018938f
C4641 a_34347_n17801# VSS 0.385498f
C4642 a_32353_n16007# VSS 0.018938f
C4643 a_35221_n15110# VSS 0.017551f
C4644 a_34699_n16904# VSS 0.550027f
C4645 a_32913_n16904# VSS 0.497494f
C4646 a_32353_n15110# VSS 0.017551f
C4647 a_35781_n15110# VSS 0.405499f
C4648 a_35221_n14213# VSS 0.016697f
C4649 a_34347_n14213# VSS 1.29606f
C4650 a_33787_n14213# VSS 0.023002f
C4651 a_32353_n14213# VSS 0.016697f
C4652 a_31831_n15110# VSS 0.405047f
C4653 a_35221_n13316# VSS 0.017066f
C4654 a_34699_n14213# VSS 0.200377f
C4655 a_33787_n13316# VSS 0.016529f
C4656 a_33265_n14213# VSS 0.178599f
C4657 a_32913_n14213# VSS 0.192438f
C4658 a_32353_n13316# VSS 0.017066f
C4659 a_35781_n13316# VSS 0.398427f
C4660 a_35221_n12419# VSS 0.025764f
C4661 a_34347_n13316# VSS 0.225452f
C4662 a_33787_n12419# VSS 0.053627f
C4663 a_32913_n12419# VSS 1.14404f
C4664 a_32353_n12419# VSS 0.025764f
C4665 a_31831_n13316# VSS 0.412143f
C4666 a_66551_n8932# VSS 0.025764f
C4667 a_65117_n8932# VSS 0.053627f
C4668 a_64243_n8932# VSS 1.10481f
C4669 a_63683_n8932# VSS 0.025764f
C4670 a_67111_n8932# VSS 0.398427f
C4671 a_66551_n8035# VSS 0.017066f
C4672 a_65677_n8932# VSS 0.225452f
C4673 a_65117_n8035# VSS 0.016529f
C4674 a_63683_n8035# VSS 0.017066f
C4675 a_63161_n8932# VSS 0.412143f
C4676 a_66551_n7138# VSS 0.016697f
C4677 a_66029_n8035# VSS 0.200377f
C4678 a_65117_n7138# VSS 0.023002f
C4679 a_64595_n8035# VSS 0.178599f
C4680 a_64243_n8035# VSS 0.192438f
C4681 a_63683_n7138# VSS 0.016697f
C4682 a_67111_n7138# VSS 0.405499f
C4683 a_66551_n6241# VSS 0.017551f
C4684 a_63683_n6241# VSS 0.017551f
C4685 a_63161_n7138# VSS 0.405047f
C4686 a_65677_n7138# VSS 1.28647f
C4687 a_66551_n5344# VSS 0.018938f
C4688 a_63683_n5344# VSS 0.018938f
C4689 a_66551_n4447# VSS 0.017564f
C4690 a_66029_n6241# VSS 0.550027f
C4691 a_64243_n6241# VSS 0.546597f
C4692 a_63683_n4447# VSS 0.017564f
C4693 a_67111_n4447# VSS 0.405615f
C4694 a_66551_n3550# VSS 0.016697f
C4695 a_65677_n3550# VSS 0.385498f
C4696 a_65117_n3550# VSS 0.023005f
C4697 a_63683_n3550# VSS 0.016697f
C4698 a_63161_n4447# VSS 0.405161f
C4699 a_66551_n2653# VSS 0.017062f
C4700 a_66029_n3550# VSS 0.227033f
C4701 a_65117_n2653# VSS 0.016525f
C4702 a_64595_n3550# VSS 0.174939f
C4703 a_64243_n3550# VSS 0.192438f
C4704 a_63683_n2653# VSS 0.017062f
C4705 a_67111_n2653# VSS 0.398946f
C4706 a_66551_n1756# VSS 0.054141f
C4707 a_65677_n2653# VSS 0.298391f
C4708 a_65117_n1756# VSS 0.025832f
C4709 a_63683_n1756# VSS 0.025741f
C4710 a_63161_n2653# VSS 0.411967f
C4711 a_60285_n8932# VSS 0.025764f
C4712 a_58851_n8932# VSS 0.053627f
C4713 a_57977_n8932# VSS 1.10481f
C4714 a_57417_n8932# VSS 0.025764f
C4715 a_60845_n8932# VSS 0.398427f
C4716 a_60285_n8035# VSS 0.017066f
C4717 a_59411_n8932# VSS 0.225452f
C4718 a_58851_n8035# VSS 0.016529f
C4719 a_57417_n8035# VSS 0.017066f
C4720 a_56895_n8932# VSS 0.412143f
C4721 a_60285_n7138# VSS 0.016697f
C4722 a_59763_n8035# VSS 0.200377f
C4723 a_58851_n7138# VSS 0.023002f
C4724 a_58329_n8035# VSS 0.178599f
C4725 a_57977_n8035# VSS 0.192438f
C4726 a_57417_n7138# VSS 0.016697f
C4727 a_60845_n7138# VSS 0.405499f
C4728 a_60285_n6241# VSS 0.017551f
C4729 a_57417_n6241# VSS 0.017551f
C4730 a_56895_n7138# VSS 0.405047f
C4731 a_59411_n7138# VSS 1.45216f
C4732 a_60285_n5344# VSS 0.018938f
C4733 a_57417_n5344# VSS 0.018938f
C4734 a_60285_n4447# VSS 0.017564f
C4735 a_59763_n6241# VSS 0.550027f
C4736 a_57977_n6241# VSS 0.546597f
C4737 a_57417_n4447# VSS 0.017564f
C4738 a_60845_n4447# VSS 0.405615f
C4739 a_60285_n3550# VSS 0.016697f
C4740 a_59411_n3550# VSS 0.385498f
C4741 a_58851_n3550# VSS 0.023005f
C4742 a_57417_n3550# VSS 0.016697f
C4743 a_56895_n4447# VSS 0.405161f
C4744 a_60285_n2653# VSS 0.017062f
C4745 a_59763_n3550# VSS 0.227033f
C4746 a_58851_n2653# VSS 0.016525f
C4747 a_58329_n3550# VSS 0.174939f
C4748 a_57977_n3550# VSS 0.192438f
C4749 a_57417_n2653# VSS 0.017062f
C4750 a_60845_n2653# VSS 0.398946f
C4751 a_60285_n1756# VSS 0.054141f
C4752 a_59411_n2653# VSS 0.298391f
C4753 a_58851_n1756# VSS 0.025832f
C4754 a_57417_n1756# VSS 0.025741f
C4755 a_56895_n2653# VSS 0.411967f
C4756 a_54019_n8932# VSS 0.025764f
C4757 a_52585_n8932# VSS 0.053627f
C4758 a_51711_n8932# VSS 1.13141f
C4759 a_51151_n8932# VSS 0.025764f
C4760 a_54579_n8932# VSS 0.398427f
C4761 a_54019_n8035# VSS 0.017066f
C4762 a_53145_n8932# VSS 0.225452f
C4763 a_52585_n8035# VSS 0.016529f
C4764 a_51151_n8035# VSS 0.017066f
C4765 a_50629_n8932# VSS 0.412149f
C4766 a_54019_n7138# VSS 0.016697f
C4767 a_53497_n8035# VSS 0.200377f
C4768 a_52585_n7138# VSS 0.023002f
C4769 a_52063_n8035# VSS 0.178599f
C4770 a_51711_n8035# VSS 0.192438f
C4771 a_51151_n7138# VSS 0.016697f
C4772 a_54579_n7138# VSS 0.405499f
C4773 a_54019_n6241# VSS 0.017551f
C4774 a_51151_n6241# VSS 0.017551f
C4775 a_50629_n7138# VSS 0.405053f
C4776 a_53145_n7138# VSS 1.28672f
C4777 a_54019_n5344# VSS 0.018938f
C4778 a_51151_n5344# VSS 0.018938f
C4779 a_54019_n4447# VSS 0.017564f
C4780 a_53497_n6241# VSS 0.550027f
C4781 a_51711_n6241# VSS 0.546597f
C4782 a_51151_n4447# VSS 0.017564f
C4783 a_54579_n4447# VSS 0.405615f
C4784 a_54019_n3550# VSS 0.016697f
C4785 a_53145_n3550# VSS 0.385498f
C4786 a_52585_n3550# VSS 0.023005f
C4787 a_51151_n3550# VSS 0.016697f
C4788 a_50629_n4447# VSS 0.405167f
C4789 a_54019_n2653# VSS 0.017062f
C4790 a_53497_n3550# VSS 0.227033f
C4791 a_52585_n2653# VSS 0.016525f
C4792 a_52063_n3550# VSS 0.174939f
C4793 a_51711_n3550# VSS 0.192438f
C4794 a_51151_n2653# VSS 0.017062f
C4795 a_54579_n2653# VSS 0.398946f
C4796 a_54019_n1756# VSS 0.054141f
C4797 a_53145_n2653# VSS 0.298391f
C4798 a_52585_n1756# VSS 0.025832f
C4799 a_51151_n1756# VSS 0.025741f
C4800 a_50629_n2653# VSS 0.411972f
C4801 a_47753_n8930# VSS 0.054141f
C4802 a_46319_n8930# VSS 0.025832f
C4803 a_44885_n8930# VSS 0.070369f
C4804 a_48313_n8930# VSS 0.398952f
C4805 a_47753_n8033# VSS 0.017062f
C4806 a_46879_n8930# VSS 0.298549f
C4807 a_46319_n8033# VSS 0.016525f
C4808 a_44885_n8033# VSS 0.024253f
C4809 a_44363_n8930# VSS 0.49306f
C4810 a_47753_n7136# VSS 0.016697f
C4811 a_47231_n8033# VSS 0.227033f
C4812 a_46319_n7136# VSS 0.023005f
C4813 a_45797_n8033# VSS 0.175025f
C4814 a_45445_n8033# VSS 0.211553f
C4815 a_44885_n7136# VSS 0.023888f
C4816 a_48313_n7136# VSS 0.40562f
C4817 a_47753_n6239# VSS 0.017564f
C4818 a_44885_n6239# VSS 0.024755f
C4819 a_44363_n7136# VSS 0.490894f
C4820 a_47753_n5342# VSS 0.018938f
C4821 a_46879_n7136# VSS 0.385498f
C4822 a_44885_n5342# VSS 0.056084f
C4823 a_47753_n4445# VSS 0.017551f
C4824 a_47231_n6239# VSS 0.550027f
C4825 a_45445_n6239# VSS 0.622493f
C4826 a_44885_n4445# VSS 0.017551f
C4827 a_48313_n4445# VSS 0.405505f
C4828 a_47753_n3548# VSS 0.016697f
C4829 a_46879_n3548# VSS 1.28675f
C4830 a_46319_n3548# VSS 0.023002f
C4831 a_44885_n3548# VSS 0.016697f
C4832 a_44363_n4445# VSS 0.417122f
C4833 a_47753_n2651# VSS 0.017066f
C4834 a_47231_n3548# VSS 0.200377f
C4835 a_46319_n2651# VSS 0.016529f
C4836 a_45797_n3548# VSS 0.178599f
C4837 a_45445_n3548# VSS 0.192438f
C4838 a_44885_n2651# VSS 0.017066f
C4839 a_48313_n2651# VSS 0.398433f
C4840 a_47753_n1754# VSS 0.025764f
C4841 a_46879_n2651# VSS 0.225452f
C4842 a_46319_n1754# VSS 0.053627f
C4843 a_45445_n1754# VSS 1.20649f
C4844 a_44885_n1754# VSS 0.025764f
C4845 a_44363_n2651# VSS 0.412143f
C4846 a_41487_n8930# VSS 0.054141f
C4847 a_40053_n8930# VSS 0.025832f
C4848 a_38619_n8930# VSS 0.025741f
C4849 a_42047_n8930# VSS 0.398946f
C4850 a_41487_n8033# VSS 0.017062f
C4851 a_40613_n8930# VSS 0.298391f
C4852 a_40053_n8033# VSS 0.016525f
C4853 a_38619_n8033# VSS 0.017062f
C4854 a_38097_n8930# VSS 0.411967f
C4855 a_41487_n7136# VSS 0.016697f
C4856 a_40965_n8033# VSS 0.227033f
C4857 a_40053_n7136# VSS 0.023005f
C4858 a_39531_n8033# VSS 0.174939f
C4859 a_39179_n8033# VSS 0.192438f
C4860 a_38619_n7136# VSS 0.016697f
C4861 a_42047_n7136# VSS 0.405615f
C4862 a_41487_n6239# VSS 0.017564f
C4863 a_38619_n6239# VSS 0.017564f
C4864 a_38097_n7136# VSS 0.405161f
C4865 a_41487_n5342# VSS 0.018938f
C4866 a_40613_n7136# VSS 0.385498f
C4867 a_38619_n5342# VSS 0.018938f
C4868 a_41487_n4445# VSS 0.017551f
C4869 a_40965_n6239# VSS 0.550027f
C4870 a_39179_n6239# VSS 0.546597f
C4871 a_38619_n4445# VSS 0.017551f
C4872 a_42047_n4445# VSS 0.405499f
C4873 a_41487_n3548# VSS 0.016697f
C4874 a_40613_n3548# VSS 1.45216f
C4875 a_40053_n3548# VSS 0.023002f
C4876 a_38619_n3548# VSS 0.016697f
C4877 a_38097_n4445# VSS 0.405047f
C4878 a_41487_n2651# VSS 0.017066f
C4879 a_40965_n3548# VSS 0.200377f
C4880 a_40053_n2651# VSS 0.016529f
C4881 a_39531_n3548# VSS 0.178599f
C4882 a_39179_n3548# VSS 0.192438f
C4883 a_38619_n2651# VSS 0.017066f
C4884 a_42047_n2651# VSS 0.398427f
C4885 a_41487_n1754# VSS 0.025764f
C4886 a_40613_n2651# VSS 0.225452f
C4887 a_40053_n1754# VSS 0.053627f
C4888 a_39179_n1754# VSS 1.20649f
C4889 a_38619_n1754# VSS 0.025764f
C4890 a_38097_n2651# VSS 0.412143f
C4891 a_35221_n8930# VSS 0.054141f
C4892 a_33787_n8930# VSS 0.025832f
C4893 a_32353_n8930# VSS 0.025741f
C4894 a_35781_n8930# VSS 0.398946f
C4895 a_35221_n8033# VSS 0.017062f
C4896 a_34347_n8930# VSS 0.298391f
C4897 a_33787_n8033# VSS 0.016525f
C4898 a_32353_n8033# VSS 0.017062f
C4899 a_31831_n8930# VSS 0.411967f
C4900 a_35221_n7136# VSS 0.016697f
C4901 a_34699_n8033# VSS 0.227033f
C4902 a_33787_n7136# VSS 0.023005f
C4903 a_33265_n8033# VSS 0.174939f
C4904 a_32913_n8033# VSS 0.192438f
C4905 a_32353_n7136# VSS 0.016697f
C4906 a_35781_n7136# VSS 0.405615f
C4907 a_35221_n6239# VSS 0.017564f
C4908 a_32353_n6239# VSS 0.017564f
C4909 a_31831_n7136# VSS 0.405161f
C4910 a_35221_n5342# VSS 0.018938f
C4911 a_34347_n7136# VSS 0.385498f
C4912 a_32353_n5342# VSS 0.018938f
C4913 a_35221_n4445# VSS 0.017551f
C4914 a_34699_n6239# VSS 0.550027f
C4915 a_32913_n6239# VSS 0.546597f
C4916 a_32353_n4445# VSS 0.017551f
C4917 a_35781_n4445# VSS 0.405499f
C4918 a_35221_n3548# VSS 0.016697f
C4919 a_34347_n3548# VSS 1.45216f
C4920 a_33787_n3548# VSS 0.023002f
C4921 a_32353_n3548# VSS 0.016697f
C4922 a_31831_n4445# VSS 0.405047f
C4923 a_35221_n2651# VSS 0.017066f
C4924 a_34699_n3548# VSS 0.200377f
C4925 a_33787_n2651# VSS 0.016529f
C4926 a_33265_n3548# VSS 0.178599f
C4927 a_32913_n3548# VSS 0.192438f
C4928 a_32353_n2651# VSS 0.017066f
C4929 a_35781_n2651# VSS 0.398427f
C4930 a_35221_n1754# VSS 0.025764f
C4931 a_34347_n2651# VSS 0.225452f
C4932 a_33787_n1754# VSS 0.053627f
C4933 a_32913_n1754# VSS 1.20649f
C4934 a_32353_n1754# VSS 0.025764f
C4935 a_31831_n2651# VSS 0.412143f
C4936 a_114485_4481# VSS 0.057864f
C4937 a_113081_4481# VSS 0.070162f
C4938 a_114485_5639# VSS 0.04696f
C4939 a_113081_5639# VSS 0.059257f
C4940 a_114485_6405# VSS 0.059789f
C4941 a_113081_6405# VSS 0.072086f
C4942 a_114485_7563# VSS 0.058211f
C4943 a_113081_7563# VSS 0.070508f
C4944 a_108602_4481# VSS 0.02113f
C4945 a_107198_4481# VSS 0.02113f
C4946 a_108602_5639# VSS 0.009003f
C4947 a_107198_5639# VSS 0.009003f
C4948 a_108602_6405# VSS 0.009003f
C4949 a_107198_6405# VSS 0.009003f
C4950 a_108602_7563# VSS 0.021386f
C4951 a_107198_7563# VSS 0.02113f
C4952 a_102796_4481# VSS 0.02113f
C4953 a_101392_4481# VSS 0.029168f
C4954 a_102796_5639# VSS 0.01202f
C4955 a_101392_5639# VSS 0.017167f
C4956 a_102796_6405# VSS 0.009003f
C4957 a_101392_6405# VSS 0.017167f
C4958 a_102796_7563# VSS 0.024094f
C4959 a_101392_7563# VSS 0.029168f
C4960 a_96818_4481# VSS 0.057864f
C4961 a_95414_4481# VSS 0.070162f
C4962 a_96818_5639# VSS 0.04696f
C4963 a_95414_5639# VSS 0.059257f
C4964 a_96818_6405# VSS 0.059789f
C4965 a_95414_6405# VSS 0.072086f
C4966 a_96818_7563# VSS 0.058211f
C4967 a_95414_7563# VSS 0.070508f
C4968 a_90935_4481# VSS 0.02113f
C4969 a_89531_4481# VSS 0.02113f
C4970 a_90935_5639# VSS 0.009003f
C4971 a_89531_5639# VSS 0.009003f
C4972 a_90935_6405# VSS 0.009003f
C4973 a_89531_6405# VSS 0.009003f
C4974 a_90935_7563# VSS 0.021386f
C4975 a_89531_7563# VSS 0.02113f
C4976 a_85129_4481# VSS 0.02113f
C4977 a_83725_4481# VSS 0.029168f
C4978 a_85129_5639# VSS 0.01202f
C4979 a_83725_5639# VSS 0.017167f
C4980 a_85129_6405# VSS 0.009003f
C4981 a_83725_6405# VSS 0.017167f
C4982 a_85129_7563# VSS 0.024094f
C4983 a_83725_7563# VSS 0.029168f
C4984 a_79151_4481# VSS 0.057864f
C4985 a_77747_4481# VSS 0.070162f
C4986 a_79151_5639# VSS 0.04696f
C4987 a_77747_5639# VSS 0.059257f
C4988 a_79151_6405# VSS 0.059789f
C4989 a_77747_6405# VSS 0.072086f
C4990 a_79151_7563# VSS 0.058211f
C4991 a_77747_7563# VSS 0.070508f
C4992 a_73268_4481# VSS 0.02113f
C4993 a_71864_4481# VSS 0.02113f
C4994 a_73268_5639# VSS 0.009003f
C4995 a_71864_5639# VSS 0.009003f
C4996 a_73268_6405# VSS 0.009003f
C4997 a_71864_6405# VSS 0.009003f
C4998 a_73268_7563# VSS 0.021386f
C4999 a_71864_7563# VSS 0.02113f
C5000 a_67462_4481# VSS 0.02113f
C5001 a_66058_4481# VSS 0.029168f
C5002 a_67462_5639# VSS 0.01202f
C5003 a_66058_5639# VSS 0.017167f
C5004 a_67462_6405# VSS 0.009003f
C5005 a_66058_6405# VSS 0.017167f
C5006 a_67462_7563# VSS 0.024094f
C5007 a_66058_7563# VSS 0.029168f
C5008 a_61484_4481# VSS 0.057864f
C5009 a_60080_4481# VSS 0.070162f
C5010 a_61484_5639# VSS 0.04696f
C5011 a_60080_5639# VSS 0.059257f
C5012 a_61484_6405# VSS 0.059789f
C5013 a_60080_6405# VSS 0.072086f
C5014 a_61484_7563# VSS 0.058211f
C5015 a_60080_7563# VSS 0.070508f
C5016 a_55601_4481# VSS 0.02113f
C5017 a_54197_4481# VSS 0.02113f
C5018 a_55601_5639# VSS 0.009003f
C5019 a_54197_5639# VSS 0.009003f
C5020 a_55601_6405# VSS 0.009003f
C5021 a_54197_6405# VSS 0.009003f
C5022 a_55601_7563# VSS 0.021386f
C5023 a_54197_7563# VSS 0.02113f
C5024 a_49795_4481# VSS 0.02113f
C5025 a_48391_4481# VSS 0.029168f
C5026 a_49795_5639# VSS 0.01202f
C5027 a_48391_5639# VSS 0.017167f
C5028 a_49795_6405# VSS 0.009003f
C5029 a_48391_6405# VSS 0.017167f
C5030 a_49795_7563# VSS 0.024094f
C5031 a_48391_7563# VSS 0.029168f
C5032 a_43817_4481# VSS 0.057864f
C5033 a_42413_4481# VSS 0.070162f
C5034 a_43817_5639# VSS 0.04696f
C5035 a_42413_5639# VSS 0.059257f
C5036 a_43817_6405# VSS 0.059789f
C5037 a_42413_6405# VSS 0.072086f
C5038 a_43817_7563# VSS 0.058211f
C5039 a_42413_7563# VSS 0.070508f
C5040 a_37934_4481# VSS 0.02113f
C5041 a_36530_4481# VSS 0.02113f
C5042 a_37934_5639# VSS 0.009003f
C5043 a_36530_5639# VSS 0.009003f
C5044 a_37934_6405# VSS 0.009003f
C5045 a_36530_6405# VSS 0.009003f
C5046 a_37934_7563# VSS 0.021386f
C5047 a_36530_7563# VSS 0.02113f
C5048 a_32128_4481# VSS 0.02113f
C5049 a_30724_4481# VSS 0.029168f
C5050 a_32128_5639# VSS 0.01202f
C5051 a_30724_5639# VSS 0.017167f
C5052 a_32128_6405# VSS 0.009003f
C5053 a_30724_6405# VSS 0.017167f
C5054 a_32128_7563# VSS 0.024094f
C5055 a_30724_7563# VSS 0.029168f
C5056 a_108636_10448# VSS 0.016627f
C5057 a_108636_11614# VSS 0.04492f
C5058 a_107230_11614# VSS 0.028915f
C5059 a_108636_12380# VSS 0.04473f
C5060 a_107230_12380# VSS 0.04473f
C5061 a_90969_10448# VSS 0.016627f
C5062 a_90969_11614# VSS 0.04492f
C5063 a_89563_11614# VSS 0.028915f
C5064 a_90969_12380# VSS 0.04473f
C5065 a_89563_12380# VSS 0.04473f
C5066 a_73302_10448# VSS 0.016627f
C5067 a_73302_11614# VSS 0.04492f
C5068 a_71896_11614# VSS 0.028915f
C5069 a_73302_12380# VSS 0.04473f
C5070 a_71896_12380# VSS 0.04473f
C5071 a_55635_10448# VSS 0.016627f
C5072 a_55635_11614# VSS 0.04492f
C5073 a_54229_11614# VSS 0.028915f
C5074 a_55635_12380# VSS 0.04473f
C5075 a_54229_12380# VSS 0.04473f
C5076 a_37968_10448# VSS 0.016627f
C5077 a_37968_11614# VSS 0.04492f
C5078 a_36562_11614# VSS 0.028915f
C5079 a_37968_12380# VSS 0.04473f
C5080 a_36562_12380# VSS 0.04473f
C5081 a_41100_19075# VSS 0.05176f
C5082 a_41100_19698# VSS 0.017025f
C5083 a_40578_19075# VSS 0.399052f
C5084 a_41660_19698# VSS 0.376201f
C5085 a_41100_20251# VSS 0.033958f
C5086 a_44608_22884# VSS 0.01042f
C5087 a_46274_23609# VSS 0.010763f
C5088 a_46274_24920# VSS 0.005065f
C5089 a_44608_24195# VSS 0.01042f
C5090 a_31699_17542# VSS 0.405869f
C5091 a_30377_18342# VSS 0.415926f
C5092 a_31699_19142# VSS 0.395971f
C5093 a_30377_19942# VSS 0.420382f
C5094 w_27790_n38888# VSS 0.430923p $ **FLOATING
C5095 a_101111_n17715.t1 VSS 0.995519f
C5096 a_101111_n17715.t0 VSS 1.00448f
C5097 IN_NEG.n0 VSS 2.14417f
C5098 IN_NEG.n1 VSS 0.167353f
C5099 IN_NEG.n2 VSS 0.124262f
C5100 IN_NEG.n3 VSS 0.046483f
C5101 IN_NEG.n4 VSS 0.051882f
C5102 IN_NEG.n5 VSS 0.122693f
C5103 IN_NEG.n6 VSS 0.17532f
C5104 IN_NEG.n7 VSS 3.88312f
C5105 IN_NEG.t1 VSS -11.2283f
C5106 IN_NEG.n8 VSS 3.9473f
C5107 IN_NEG.n9 VSS 1.12359f
C5108 IN_NEG.n10 VSS 2.68065f
C5109 IN_NEG.n11 VSS 0.173712f
C5110 IN_NEG.n12 VSS 0.840066f
C5111 IN_NEG.n13 VSS 1.8676f
C5112 IN_NEG.n14 VSS 0.138196f
C5113 IN_NEG.n15 VSS 0.604481f
C5114 IN_NEG.n16 VSS 1.08259f
C5115 IN_NEG.n17 VSS 0.10963f
C5116 IN_NEG.n18 VSS 0.434304f
C5117 IN_NEG.n19 VSS 0.401753f
C5118 IN_NEG.n20 VSS 0.09853f
C5119 IN_NEG.n21 VSS 0.591504f
C5120 IN_NEG.n22 VSS 1.06551f
C5121 IN_NEG.n23 VSS 0.135608f
C5122 IN_NEG.n24 VSS 0.839584f
C5123 IN_NEG.n25 VSS 1.87274f
C5124 IN_NEG.n26 VSS 0.177873f
C5125 IN_NEG.n27 VSS 2.63138f
C5126 IN_NEG.n28 VSS 1.09392f
C5127 IN_NEG.n29 VSS 2.1073f
C5128 IN_NEG.t0 VSS 12.679f
C5129 IN_NEG.n30 VSS 7.87284f
C5130 a_84017_n16810.t1 VSS 0.995519f
C5131 a_84017_n16810.t0 VSS 1.00448f
C5132 IBPOUT.t0 VSS 0.154788f
C5133 a_45445_n16007.t1 VSS 1.26793f
C5134 a_45445_n16007.t0 VSS 1.23207f
C5135 a_32913_n16007.t1 VSS 1.23207f
C5136 a_32913_n16007.t0 VSS 1.26793f
C5137 a_95413_n16810.t1 VSS 0.995519f
C5138 a_95413_n16810.t0 VSS 1.00448f
C5139 a_112507_n6055.t1 VSS 0.995519f
C5140 a_112507_n6055.t0 VSS 1.00448f
C5141 a_95413_n5150.t1 VSS 0.995519f
C5142 a_95413_n5150.t0 VSS 1.00448f
C5143 a_106676_n27257.n0 VSS 9.95669f
C5144 a_106676_n27257.t0 VSS 0.704006f
C5145 a_106676_n27257.t1 VSS 0.606767f
C5146 a_106676_n27257.t3 VSS 0.922584f
C5147 a_106676_n27257.t2 VSS 0.509953f
C5148 a_84017_n5150.t1 VSS 0.995519f
C5149 a_84017_n5150.t0 VSS 1.00448f
C5150 a_71266_n4019.t0 VSS 19.538f
C5151 a_71266_n4019.t1 VSS 16.362f
C5152 a_36008_n27257.n0 VSS 9.956639f
C5153 a_36008_n27257.t2 VSS 0.704006f
C5154 a_36008_n27257.t3 VSS 0.606767f
C5155 a_36008_n27257.t1 VSS 0.509953f
C5156 a_36008_n27257.t0 VSS 0.922634f
C5157 a_57977_n16009.t1 VSS 1.26787f
C5158 a_57977_n16009.t0 VSS 1.23213f
C5159 a_64243_n16009.t1 VSS 1.26787f
C5160 a_64243_n16009.t0 VSS 1.23213f
C5161 a_43010_n36322.t0 VSS 3.08334f
C5162 a_43010_n36322.t2 VSS 51.9827f
C5163 a_43010_n36322.t1 VSS 1.84861f
C5164 a_43010_n36322.t3 VSS 33.885303f
C5165 a_45445_n5342.t1 VSS 1.26793f
C5166 a_45445_n5342.t0 VSS 1.23207f
C5167 a_53675_7563.n0 VSS 10.6245f
C5168 a_53675_7563.t3 VSS 0.812605f
C5169 a_53675_7563.t0 VSS 0.843931f
C5170 a_53675_7563.t1 VSS 0.685986f
C5171 a_53675_7563.t2 VSS 0.632999f
C5172 a_112507_n17715.t1 VSS 0.995519f
C5173 a_112507_n17715.t0 VSS 1.00448f
C5174 a_89009_n30339.n0 VSS 10.6245f
C5175 a_89009_n30339.t1 VSS 0.843931f
C5176 a_89009_n30339.t0 VSS 0.685986f
C5177 a_89009_n30339.t3 VSS 0.812605f
C5178 a_89009_n30339.t2 VSS 0.632986f
C5179 a_36008_n30339.n0 VSS 10.6245f
C5180 a_36008_n30339.t2 VSS 0.843931f
C5181 a_36008_n30339.t3 VSS 0.685986f
C5182 a_36008_n30339.t1 VSS 0.812605f
C5183 a_36008_n30339.t0 VSS 0.632986f
C5184 VCM.t2 VSS 3.82305f
C5185 VCM.t3 VSS 2.11966f
C5186 VCM.n0 VSS 4.64613f
C5187 VCM.t0 VSS 0.091648f
C5188 VCM.t1 VSS 0.088287f
C5189 VCM.n1 VSS 3.62553f
C5190 VCM.n2 VSS 5.40563f
C5191 a_106809_n6055.t1 VSS 0.995519f
C5192 a_106809_n6055.t0 VSS 1.00448f
C5193 a_39179_n5342.t1 VSS 1.26793f
C5194 a_39179_n5342.t0 VSS 1.23207f
C5195 a_89009_4481.n0 VSS 9.956611f
C5196 a_89009_4481.t0 VSS 0.704006f
C5197 a_89009_4481.t1 VSS 0.606767f
C5198 a_89009_4481.t3 VSS 0.509963f
C5199 a_89009_4481.t2 VSS 0.92265f
C5200 a_64243_n5344.t1 VSS 1.26787f
C5201 a_64243_n5344.t0 VSS 1.23213f
C5202 a_89715_n5150.t1 VSS 1.00453f
C5203 a_89715_n5150.t0 VSS 0.995467f
C5204 a_51711_n16009.t1 VSS 1.26787f
C5205 a_51711_n16009.t0 VSS 1.23213f
C5206 a_53675_n27257.n0 VSS 9.956639f
C5207 a_53675_n27257.t1 VSS 0.704006f
C5208 a_53675_n27257.t0 VSS 0.606767f
C5209 a_53675_n27257.t3 VSS 0.509953f
C5210 a_53675_n27257.t2 VSS 0.922634f
C5211 a_89033_n36322.t2 VSS 0.781529f
C5212 a_89033_n36322.t3 VSS 0.752866f
C5213 a_89033_n36322.n0 VSS 8.139339f
C5214 a_89033_n36322.t1 VSS 0.676033f
C5215 a_89033_n36322.n1 VSS 8.25763f
C5216 a_89033_n36322.t0 VSS 0.792603f
C5217 a_94892_4481.t8 VSS 3.64456f
C5218 a_94892_4481.n0 VSS 0.449404f
C5219 a_94892_4481.n1 VSS 7.74464f
C5220 a_94892_4481.t9 VSS 0.182047f
C5221 a_94892_4481.t5 VSS 0.177333f
C5222 a_94892_4481.t7 VSS 0.152849f
C5223 a_94892_4481.t4 VSS 0.296925f
C5224 a_94892_4481.t17 VSS 0.284336f
C5225 a_94892_4481.t19 VSS 0.293711f
C5226 a_94892_4481.t14 VSS 0.296925f
C5227 a_94892_4481.t15 VSS 0.284336f
C5228 a_94892_4481.t20 VSS 0.296925f
C5229 a_94892_4481.t21 VSS 0.284336f
C5230 a_94892_4481.t2 VSS 0.294005f
C5231 a_94892_4481.t22 VSS 0.284359f
C5232 a_94892_4481.t1 VSS 0.177256f
C5233 a_94892_4481.t3 VSS 0.152918f
C5234 a_94892_4481.t0 VSS 0.296925f
C5235 a_94892_4481.t11 VSS 0.284336f
C5236 a_94892_4481.t13 VSS 0.293956f
C5237 a_94892_4481.t12 VSS 0.284359f
C5238 a_94892_4481.t16 VSS 0.284359f
C5239 a_94892_4481.t6 VSS 0.293809f
C5240 a_94892_4481.t18 VSS 0.284359f
C5241 a_94892_4481.t10 VSS 0.181041f
C5242 IN_POS.n0 VSS 4.48494f
C5243 IN_POS.n1 VSS 4.29823f
C5244 IN_POS.n2 VSS 0.112587f
C5245 IN_POS.n3 VSS 0.150651f
C5246 IN_POS.n4 VSS 0.197583f
C5247 IN_POS.n5 VSS 0.109064f
C5248 IN_POS.n6 VSS 0.152994f
C5249 IN_POS.n7 VSS 0.192313f
C5250 IN_POS.n8 VSS 0.185273f
C5251 IN_POS.n9 VSS 0.278197f
C5252 IN_POS.n10 VSS 1.21126f
C5253 IN_POS.n11 VSS 0.442472f
C5254 IN_POS.n12 VSS 2.06759f
C5255 IN_POS.n13 VSS 0.930021f
C5256 IN_POS.n14 VSS 0.137568f
C5257 IN_POS.n15 VSS 2.3333f
C5258 IN_POS.n16 VSS 2.91269f
C5259 IN_POS.n17 VSS 1.21105f
C5260 IN_POS.n18 VSS 0.194093f
C5261 IN_POS.n19 VSS 2.07287f
C5262 IN_POS.n20 VSS 0.929487f
C5263 IN_POS.n21 VSS 0.135831f
C5264 IN_POS.n22 VSS 0.441933f
C5265 IN_POS.n23 VSS 0.480809f
C5266 IN_POS.n24 VSS 1.17853f
C5267 IN_POS.n25 VSS 0.658594f
C5268 IN_POS.n26 VSS 0.053687f
C5269 IN_POS.t0 VSS -0.890219f
C5270 IN_POS.n27 VSS 1.94474f
C5271 IN_POS.n28 VSS 1.2439f
C5272 IN_POS.n29 VSS 2.94329f
C5273 IN_POS.n30 VSS 0.229628f
C5274 IN_POS.t1 VSS -14.683901f
C5275 IN_POS.n31 VSS 12.7299f
C5276 IN_POS.n32 VSS 5.28104f
C5277 a_101111_n6055.t1 VSS 1.00453f
C5278 a_101111_n6055.t0 VSS 0.995467f
C5279 a_36032_13546.t2 VSS 0.77626f
C5280 a_36032_13546.t3 VSS 0.662094f
C5281 a_36032_13546.n0 VSS 8.089789f
C5282 a_36032_13546.t1 VSS 0.737343f
C5283 a_36032_13546.n1 VSS 7.9691f
C5284 a_36032_13546.t0 VSS 0.765415f
C5285 a_89009_7563.n0 VSS 10.6245f
C5286 a_89009_7563.t0 VSS 0.843931f
C5287 a_89009_7563.t1 VSS 0.685986f
C5288 a_89009_7563.t3 VSS 0.632998f
C5289 a_89009_7563.t2 VSS 0.812605f
C5290 a_36008_7563.n0 VSS 10.6245f
C5291 a_36008_7563.t1 VSS 0.812605f
C5292 a_36008_7563.t2 VSS 0.843931f
C5293 a_36008_7563.t3 VSS 0.685986f
C5294 a_36008_7563.t0 VSS 0.632999f
C5295 a_106830_n36382.n0 VSS 2.51436f
C5296 a_106830_n36382.n1 VSS 9.83545f
C5297 a_106830_n36382.n2 VSS 0.932965f
C5298 a_106830_n36382.n3 VSS 1.58916f
C5299 a_106830_n36382.n4 VSS 5.82997f
C5300 a_106830_n36382.n5 VSS 7.8766f
C5301 a_106830_n36382.n6 VSS 0.903342f
C5302 a_106830_n36382.t11 VSS 0.56727f
C5303 a_106830_n36382.t12 VSS 0.600109f
C5304 a_106830_n36382.t8 VSS 0.567069f
C5305 a_106830_n36382.t6 VSS 0.343871f
C5306 a_106830_n36382.t2 VSS 0.593475f
C5307 a_106830_n36382.t0 VSS 0.31856f
C5308 a_106830_n36382.t3 VSS 0.323606f
C5309 a_106830_n36382.t1 VSS 0.493914f
C5310 a_106830_n36382.t7 VSS 0.521169f
C5311 a_106830_n36382.t16 VSS 0.558714f
C5312 a_106830_n36382.t21 VSS 0.558674f
C5313 a_106830_n36382.t15 VSS 0.556508f
C5314 a_106830_n36382.t10 VSS 0.556508f
C5315 a_106830_n36382.t18 VSS 0.556508f
C5316 a_106830_n36382.t23 VSS 0.556508f
C5317 a_106830_n36382.t17 VSS 0.558581f
C5318 a_106830_n36382.t20 VSS 0.558735f
C5319 a_106830_n36382.t14 VSS 0.556508f
C5320 a_106830_n36382.t13 VSS 0.556508f
C5321 a_106830_n36382.t19 VSS 0.556508f
C5322 a_106830_n36382.t9 VSS 0.566653f
C5323 a_106830_n36382.t22 VSS 0.556508f
C5324 a_106830_n36382.t5 VSS 0.51848f
C5325 a_106830_n36382.n7 VSS 0.904225f
C5326 a_106830_n36382.t4 VSS 0.312958f
C5327 a_106676_7563.n0 VSS 10.6245f
C5328 a_106676_7563.t3 VSS 0.812605f
C5329 a_106676_7563.t1 VSS 0.843931f
C5330 a_106676_7563.t0 VSS 0.685986f
C5331 a_106676_7563.t2 VSS 0.632999f
C5332 a_39179_n8930.t1 VSS 59.5026f
C5333 a_39179_n8930.t2 VSS 2.36783f
C5334 a_39179_n8930.t0 VSS 30.229502f
C5335 a_50629_n16009.t1 VSS 48.396698f
C5336 a_50629_n16009.t0 VSS 6.29607f
C5337 a_50629_n16009.t2 VSS 33.0072f
C5338 a_71342_n27257.n0 VSS 9.95669f
C5339 a_71342_n27257.t0 VSS 0.704006f
C5340 a_71342_n27257.t1 VSS 0.606767f
C5341 a_71342_n27257.t3 VSS 0.922584f
C5342 a_71342_n27257.t2 VSS 0.509952f
C5343 a_30324_5507.t1 VSS 34.531998f
C5344 a_30324_5507.t2 VSS 1.63453f
C5345 a_30324_5507.t0 VSS 16.5335f
C5346 a_71366_n36322.t3 VSS 0.793614f
C5347 a_71366_n36322.t2 VSS 0.764508f
C5348 a_71366_n36322.n0 VSS 8.26458f
C5349 a_71366_n36322.t1 VSS 0.686487f
C5350 a_71366_n36322.n1 VSS 8.385951f
C5351 a_71366_n36322.t0 VSS 0.804859f
C5352 a_39179_n16007.t1 VSS 1.23207f
C5353 a_39179_n16007.t0 VSS 1.26793f
C5354 a_65658_n29313.t0 VSS 23.122198f
C5355 a_65658_n29313.t1 VSS 8.80583f
C5356 a_65658_n29313.t2 VSS 7.57194f
C5357 a_32913_n5342.t1 VSS 1.23207f
C5358 a_32913_n5342.t0 VSS 1.26793f
C5359 a_36162_10388.n0 VSS 2.54961f
C5360 a_36162_10388.n1 VSS 9.97333f
C5361 a_36162_10388.n2 VSS 0.946045f
C5362 a_36162_10388.n3 VSS 1.61144f
C5363 a_36162_10388.n4 VSS 5.9117f
C5364 a_36162_10388.n5 VSS 7.98701f
C5365 a_36162_10388.n6 VSS 0.915998f
C5366 a_36162_10388.t22 VSS 0.575018f
C5367 a_36162_10388.t12 VSS 0.575223f
C5368 a_36162_10388.t23 VSS 0.608523f
C5369 a_36162_10388.t21 VSS 0.574597f
C5370 a_36162_10388.t6 VSS 0.348688f
C5371 a_36162_10388.t16 VSS 0.566547f
C5372 a_36162_10388.t17 VSS 0.566506f
C5373 a_36162_10388.t13 VSS 0.56431f
C5374 a_36162_10388.t14 VSS 0.56431f
C5375 a_36162_10388.t11 VSS 0.56431f
C5376 a_36162_10388.t9 VSS 0.56431f
C5377 a_36162_10388.t15 VSS 0.566411f
C5378 a_36162_10388.t20 VSS 0.566568f
C5379 a_36162_10388.t8 VSS 0.56431f
C5380 a_36162_10388.t10 VSS 0.56431f
C5381 a_36162_10388.t19 VSS 0.56431f
C5382 a_36162_10388.t18 VSS 0.56431f
C5383 a_36162_10388.t5 VSS 0.525765f
C5384 a_36162_10388.t2 VSS 0.601787f
C5385 a_36162_10388.t0 VSS 0.323035f
C5386 a_36162_10388.t1 VSS 0.328142f
C5387 a_36162_10388.t3 VSS 0.500853f
C5388 a_36162_10388.t7 VSS 0.528477f
C5389 a_36162_10388.n7 VSS 0.916908f
C5390 a_36162_10388.t4 VSS 0.317345f
C5391 a_53675_4481.n0 VSS 9.95668f
C5392 a_53675_4481.t3 VSS 0.922601f
C5393 a_53675_4481.t0 VSS 0.704006f
C5394 a_53675_4481.t1 VSS 0.606767f
C5395 a_53675_4481.t2 VSS 0.50995f
C5396 a_38097_n16007.t1 VSS 6.98815f
C5397 a_38097_n16007.t2 VSS 51.744198f
C5398 a_38097_n16007.t0 VSS 24.7676f
C5399 a_78344_10448.t0 VSS 61.014305f
C5400 a_78344_10448.t3 VSS 0.47299f
C5401 a_78344_10448.t1 VSS 0.931156f
C5402 a_78344_10448.t2 VSS 0.7853f
C5403 a_78344_10448.t4 VSS 27.6962f
C5404 a_71366_11614.n0 VSS 11.663199f
C5405 a_71366_11614.n1 VSS 55.209698f
C5406 a_71366_11614.t1 VSS 3.83162f
C5407 a_71366_11614.t8 VSS 0.958145f
C5408 a_71366_11614.n2 VSS 4.27801f
C5409 a_71366_11614.t9 VSS 0.97727f
C5410 a_71366_11614.t10 VSS 0.876653f
C5411 a_71366_11614.t4 VSS 0.876653f
C5412 a_71366_11614.t6 VSS 0.930598f
C5413 a_71366_11614.t3 VSS 0.876653f
C5414 a_71366_11614.t7 VSS 0.876653f
C5415 a_71366_11614.t5 VSS 0.859167f
C5416 a_71366_11614.t2 VSS 19.8418f
C5417 a_71366_11614.t0 VSS 0.243962f
C5418 a_71342_7563.n0 VSS 10.6245f
C5419 a_71342_7563.t3 VSS 0.812605f
C5420 a_71342_7563.t1 VSS 0.843931f
C5421 a_71342_7563.t0 VSS 0.685986f
C5422 a_71342_7563.t2 VSS 0.632999f
C5423 a_36162_n36382.n0 VSS 2.54373f
C5424 a_36162_n36382.n1 VSS 9.950349f
C5425 a_36162_n36382.n2 VSS 0.943864f
C5426 a_36162_n36382.n3 VSS 1.60773f
C5427 a_36162_n36382.n4 VSS 0.914774f
C5428 a_36162_n36382.n5 VSS 5.89808f
C5429 a_36162_n36382.n6 VSS 7.968601f
C5430 a_36162_n36382.n7 VSS 0.913895f
C5431 a_36162_n36382.t18 VSS 0.573897f
C5432 a_36162_n36382.t19 VSS 0.60712f
C5433 a_36162_n36382.t11 VSS 0.573693f
C5434 a_36162_n36382.t7 VSS 0.600409f
C5435 a_36162_n36382.t6 VSS 0.322282f
C5436 a_36162_n36382.t4 VSS 0.327386f
C5437 a_36162_n36382.t5 VSS 0.499684f
C5438 a_36162_n36382.t3 VSS 0.527258f
C5439 a_36162_n36382.t1 VSS 0.316629f
C5440 a_36162_n36382.t2 VSS 0.347889f
C5441 a_36162_n36382.t20 VSS 0.565241f
C5442 a_36162_n36382.t23 VSS 0.5652f
C5443 a_36162_n36382.t15 VSS 0.56301f
C5444 a_36162_n36382.t8 VSS 0.56301f
C5445 a_36162_n36382.t9 VSS 0.56301f
C5446 a_36162_n36382.t17 VSS 0.56301f
C5447 a_36162_n36382.t21 VSS 0.565106f
C5448 a_36162_n36382.t22 VSS 0.565262f
C5449 a_36162_n36382.t14 VSS 0.56301f
C5450 a_36162_n36382.t10 VSS 0.56301f
C5451 a_36162_n36382.t12 VSS 0.56301f
C5452 a_36162_n36382.t13 VSS 0.573273f
C5453 a_36162_n36382.t16 VSS 0.56301f
C5454 a_36162_n36382.t0 VSS 0.524551f
C5455 a_71366_13546.t2 VSS 0.753329f
C5456 a_71366_13546.t3 VSS 0.725701f
C5457 a_71366_13546.n0 VSS 7.84506f
C5458 a_71366_13546.t1 VSS 0.764004f
C5459 a_71366_13546.n1 VSS 7.96027f
C5460 a_71366_13546.t0 VSS 0.65164f
C5461 a_89715_n16810.t1 VSS 1.00453f
C5462 a_89715_n16810.t0 VSS 0.995467f
C5463 I1N.t3 VSS 0.039015f
C5464 I1N.n0 VSS 0.185846f
C5465 I1N.n1 VSS 0.459261f
C5466 I1N.t4 VSS 0.569267f
C5467 I1N.n2 VSS 0.129935f
C5468 I1N.t12 VSS 0.567877f
C5469 I1N.t17 VSS 0.567877f
C5470 I1N.n3 VSS 0.620332f
C5471 I1N.n4 VSS 0.093095f
C5472 I1N.n5 VSS 0.130474f
C5473 I1N.t8 VSS 0.472566f
C5474 I1N.n6 VSS 0.519707f
C5475 I1N.t5 VSS 0.472566f
C5476 I1N.n7 VSS 0.459261f
C5477 I1N.t1 VSS 0.181106f
C5478 I1N.n8 VSS 0.486982f
C5479 I1N.n9 VSS 0.459261f
C5480 I1N.t7 VSS 0.696518f
C5481 I1N.t0 VSS 0.693737f
C5482 I1N.t14 VSS 0.503115f
C5483 I1N.n10 VSS 0.459261f
C5484 I1N.n11 VSS 0.065378f
C5485 I1N.n12 VSS 0.461407f
C5486 I1N.t9 VSS 0.503115f
C5487 I1N.n13 VSS 0.461407f
C5488 I1N.n14 VSS 0.065378f
C5489 I1N.n15 VSS 0.12141f
C5490 I1N.n16 VSS 0.135111f
C5491 I1N.n17 VSS 0.065378f
C5492 I1N.n18 VSS 0.619862f
C5493 I1N.t10 VSS 0.569267f
C5494 I1N.n19 VSS 0.461407f
C5495 I1N.t15 VSS 0.472566f
C5496 I1N.n20 VSS 0.519667f
C5497 I1N.t11 VSS 0.472566f
C5498 I1N.n21 VSS 0.461407f
C5499 I1N.n22 VSS 0.065378f
C5500 I1N.n23 VSS 0.133755f
C5501 I1N.n24 VSS 0.121817f
C5502 I1N.n25 VSS 0.459261f
C5503 I1N.t2 VSS 0.689458f
C5504 I1N.t6 VSS 0.687983f
C5505 I1N.t13 VSS 0.503115f
C5506 I1N.n26 VSS 0.447321f
C5507 I1N.n27 VSS 0.065378f
C5508 I1N.n28 VSS 0.461407f
C5509 I1N.t16 VSS 0.503115f
C5510 I1N.n29 VSS 0.446733f
C5511 I1N.n30 VSS 0.065378f
C5512 I1N.n31 VSS -6.14373f
C5513 I1N.n32 VSS 0.167762f
C5514 a_65658_4421.t0 VSS 25.151001f
C5515 a_65658_4421.t2 VSS 13.2043f
C5516 a_65658_4421.t1 VSS 1.14464f
C5517 a_53699_11614.n0 VSS 11.7253f
C5518 a_53699_11614.t0 VSS 54.606003f
C5519 a_53699_11614.t7 VSS 0.963247f
C5520 a_53699_11614.n1 VSS 4.30079f
C5521 a_53699_11614.t1 VSS 0.937962f
C5522 a_53699_11614.t8 VSS 0.982475f
C5523 a_53699_11614.t10 VSS 0.881321f
C5524 a_53699_11614.t6 VSS 0.881321f
C5525 a_53699_11614.t5 VSS 0.935554f
C5526 a_53699_11614.t3 VSS 0.881321f
C5527 a_53699_11614.t9 VSS 0.881321f
C5528 a_53699_11614.t4 VSS 0.863743f
C5529 a_53699_11614.t2 VSS 23.3596f
C5530 a_53699_13546.t2 VSS 0.77626f
C5531 a_53699_13546.t3 VSS 0.662094f
C5532 a_53699_13546.n0 VSS 8.0887f
C5533 a_53699_13546.t1 VSS 0.737343f
C5534 a_53699_13546.n1 VSS 7.97019f
C5535 a_53699_13546.t0 VSS 0.765415f
C5536 a_53829_10388.n0 VSS 2.53786f
C5537 a_53829_10388.n1 VSS 9.92737f
C5538 a_53829_10388.n2 VSS 0.941685f
C5539 a_53829_10388.n3 VSS 1.60401f
C5540 a_53829_10388.n4 VSS 5.88445f
C5541 a_53829_10388.n5 VSS 7.950201f
C5542 a_53829_10388.n6 VSS 0.911776f
C5543 a_53829_10388.t12 VSS 0.572368f
C5544 a_53829_10388.t21 VSS 0.572572f
C5545 a_53829_10388.t14 VSS 0.605719f
C5546 a_53829_10388.t11 VSS 0.571949f
C5547 a_53829_10388.t6 VSS 0.315882f
C5548 a_53829_10388.t9 VSS 0.563936f
C5549 a_53829_10388.t10 VSS 0.563895f
C5550 a_53829_10388.t17 VSS 0.561709f
C5551 a_53829_10388.t20 VSS 0.561709f
C5552 a_53829_10388.t19 VSS 0.561709f
C5553 a_53829_10388.t15 VSS 0.561709f
C5554 a_53829_10388.t8 VSS 0.563801f
C5555 a_53829_10388.t16 VSS 0.563957f
C5556 a_53829_10388.t13 VSS 0.561709f
C5557 a_53829_10388.t18 VSS 0.561709f
C5558 a_53829_10388.t23 VSS 0.561709f
C5559 a_53829_10388.t22 VSS 0.561709f
C5560 a_53829_10388.t7 VSS 0.523342f
C5561 a_53829_10388.t3 VSS 0.599013f
C5562 a_53829_10388.t0 VSS 0.321546f
C5563 a_53829_10388.t2 VSS 0.32663f
C5564 a_53829_10388.t1 VSS 0.498545f
C5565 a_53829_10388.t5 VSS 0.526042f
C5566 a_53829_10388.n7 VSS 0.912681f
C5567 a_53829_10388.t4 VSS 0.347081f
C5568 a_65486_11614.n0 VSS 0.727613f
C5569 a_65486_11614.n1 VSS 11.477901f
C5570 a_65486_11614.n2 VSS 11.550099f
C5571 a_65486_11614.t17 VSS 0.458761f
C5572 a_65486_11614.t9 VSS 0.458717f
C5573 a_65486_11614.t1 VSS 0.509737f
C5574 a_65486_11614.t3 VSS 0.260912f
C5575 a_65486_11614.t2 VSS 0.278471f
C5576 a_65486_11614.t14 VSS 0.452124f
C5577 a_65486_11614.t18 VSS 0.452124f
C5578 a_65486_11614.t20 VSS 0.450255f
C5579 a_65486_11614.t16 VSS 0.450255f
C5580 a_65486_11614.t11 VSS 0.450255f
C5581 a_65486_11614.t13 VSS 0.458761f
C5582 a_65486_11614.t15 VSS 0.450255f
C5583 a_65486_11614.t22 VSS 0.452124f
C5584 a_65486_11614.t10 VSS 0.452124f
C5585 a_65486_11614.t12 VSS 0.450255f
C5586 a_65486_11614.t23 VSS 0.450255f
C5587 a_65486_11614.t19 VSS 0.450255f
C5588 a_65486_11614.t21 VSS 0.458717f
C5589 a_65486_11614.t8 VSS 0.450255f
C5590 a_65486_11614.t4 VSS 0.410824f
C5591 a_65486_11614.t5 VSS 0.242329f
C5592 a_65486_11614.t7 VSS 0.273794f
C5593 a_65486_11614.t6 VSS 0.423369f
C5594 a_65486_11614.t0 VSS 0.399525f
C5595 a_60677_n36322.t2 VSS 3.06439f
C5596 a_60677_n36322.t1 VSS 57.1458f
C5597 a_60677_n36322.t3 VSS 1.83725f
C5598 a_60677_n36322.t0 VSS 28.752499f
C5599 a_53675_n30339.n0 VSS 10.6245f
C5600 a_53675_n30339.t0 VSS 0.843931f
C5601 a_53675_n30339.t1 VSS 0.685986f
C5602 a_53675_n30339.t3 VSS 0.632984f
C5603 a_53675_n30339.t2 VSS 0.812605f
C5604 a_59558_n29181.t8 VSS 3.64456f
C5605 a_59558_n29181.n0 VSS 4.17871f
C5606 a_59558_n29181.n1 VSS 4.01532f
C5607 a_59558_n29181.t1 VSS 0.177332f
C5608 a_59558_n29181.t7 VSS 0.152852f
C5609 a_59558_n29181.t0 VSS 0.296925f
C5610 a_59558_n29181.t15 VSS 0.284336f
C5611 a_59558_n29181.t12 VSS 0.293711f
C5612 a_59558_n29181.t17 VSS 0.296925f
C5613 a_59558_n29181.t13 VSS 0.284336f
C5614 a_59558_n29181.t11 VSS 0.296925f
C5615 a_59558_n29181.t21 VSS 0.284336f
C5616 a_59558_n29181.t4 VSS 0.294005f
C5617 a_59558_n29181.t22 VSS 0.284359f
C5618 a_59558_n29181.t3 VSS 0.177255f
C5619 a_59558_n29181.t5 VSS 0.152921f
C5620 a_59558_n29181.t2 VSS 0.296925f
C5621 a_59558_n29181.t19 VSS 0.284336f
C5622 a_59558_n29181.t18 VSS 0.293956f
C5623 a_59558_n29181.t20 VSS 0.284359f
C5624 a_59558_n29181.t14 VSS 0.284359f
C5625 a_59558_n29181.t6 VSS 0.293809f
C5626 a_59558_n29181.t16 VSS 0.284359f
C5627 a_59558_n29181.t10 VSS 0.182045f
C5628 a_59558_n29181.t9 VSS 0.181038f
C5629 a_47991_n29313.t0 VSS 23.122198f
C5630 a_47991_n29313.t1 VSS 8.80583f
C5631 a_47991_n29313.t2 VSS 7.57194f
C5632 a_48951_4481.t2 VSS 5.00668f
C5633 a_48951_4481.t1 VSS 46.7297f
C5634 a_48951_4481.t0 VSS 31.663698f
C5635 a_47991_5507.t0 VSS 71.2991f
C5636 a_47991_5507.t2 VSS 2.73325f
C5637 a_47991_5507.t1 VSS 14.967599f
C5638 a_103997_n8770.t10 VSS 0.90388f
C5639 a_103997_n8770.n0 VSS 11.0025f
C5640 a_103997_n8770.n1 VSS 4.03565f
C5641 a_103997_n8770.t9 VSS 0.921926f
C5642 a_103997_n8770.t8 VSS 0.82699f
C5643 a_103997_n8770.t12 VSS 0.82699f
C5644 a_103997_n8770.t5 VSS 0.877864f
C5645 a_103997_n8770.t7 VSS 0.82699f
C5646 a_103997_n8770.t11 VSS 0.82699f
C5647 a_103997_n8770.t6 VSS 0.810495f
C5648 a_103997_n8770.t2 VSS 0.62174f
C5649 a_103997_n8770.n2 VSS 0.898369f
C5650 a_103997_n8770.t1 VSS 3.70434f
C5651 a_103997_n8770.t4 VSS 0.236575f
C5652 a_103997_n8770.t3 VSS 0.230142f
C5653 a_103997_n8770.n3 VSS 57.1449f
C5654 a_103997_n8770.t0 VSS 25.2037f
C5655 a_57977_n5344.t1 VSS 1.23213f
C5656 a_57977_n5344.t0 VSS 1.26787f
C5657 a_47991_4421.t0 VSS 25.151001f
C5658 a_47991_4421.t1 VSS 13.2043f
C5659 a_47991_4421.t2 VSS 1.14464f
C5660 a_47819_11614.n0 VSS 0.727613f
C5661 a_47819_11614.n1 VSS 11.477901f
C5662 a_47819_11614.n2 VSS 11.550099f
C5663 a_47819_11614.t13 VSS 0.458761f
C5664 a_47819_11614.t21 VSS 0.458717f
C5665 a_47819_11614.t19 VSS 0.452124f
C5666 a_47819_11614.t23 VSS 0.452124f
C5667 a_47819_11614.t8 VSS 0.450255f
C5668 a_47819_11614.t20 VSS 0.450255f
C5669 a_47819_11614.t11 VSS 0.450255f
C5670 a_47819_11614.t9 VSS 0.458761f
C5671 a_47819_11614.t14 VSS 0.450255f
C5672 a_47819_11614.t10 VSS 0.452124f
C5673 a_47819_11614.t17 VSS 0.452124f
C5674 a_47819_11614.t18 VSS 0.450255f
C5675 a_47819_11614.t12 VSS 0.450255f
C5676 a_47819_11614.t16 VSS 0.450255f
C5677 a_47819_11614.t15 VSS 0.458717f
C5678 a_47819_11614.t22 VSS 0.450255f
C5679 a_47819_11614.t6 VSS 0.410823f
C5680 a_47819_11614.t5 VSS 0.242329f
C5681 a_47819_11614.t7 VSS 0.273794f
C5682 a_47819_11614.t4 VSS 0.423369f
C5683 a_47819_11614.t3 VSS 0.399525f
C5684 a_47819_11614.t2 VSS 0.260912f
C5685 a_47819_11614.t1 VSS 0.278471f
C5686 a_47819_11614.t0 VSS 0.509737f
C5687 a_83153_10448.t1 VSS 20.5853f
C5688 a_83153_10448.t2 VSS 1.77451f
C5689 a_83153_10448.t11 VSS 0.34777f
C5690 a_83153_10448.t3 VSS 0.330207f
C5691 a_83153_10448.t0 VSS 0.329925f
C5692 a_83153_10448.t12 VSS 0.568066f
C5693 a_83153_10448.t19 VSS 0.544019f
C5694 a_83153_10448.t18 VSS 0.544019f
C5695 a_83153_10448.t4 VSS 0.562597f
C5696 a_83153_10448.t17 VSS 0.568066f
C5697 a_83153_10448.t23 VSS 0.544019f
C5698 a_83153_10448.t8 VSS 0.568066f
C5699 a_83153_10448.t15 VSS 0.544019f
C5700 a_83153_10448.t13 VSS 0.544019f
C5701 a_83153_10448.t20 VSS 0.562597f
C5702 a_83153_10448.t9 VSS 0.34777f
C5703 a_83153_10448.t7 VSS 0.30485f
C5704 a_83153_10448.t6 VSS 0.562597f
C5705 a_83153_10448.t22 VSS 0.544019f
C5706 a_83153_10448.t10 VSS 0.568066f
C5707 a_83153_10448.t16 VSS 0.544019f
C5708 a_83153_10448.t21 VSS 0.562597f
C5709 a_83153_10448.t14 VSS 0.544019f
C5710 a_83153_10448.t5 VSS 0.30485f
C5711 a_83153_n36322.n0 VSS 11.550099f
C5712 a_83153_n36322.n1 VSS 0.727597f
C5713 a_83153_n36322.n2 VSS 11.477901f
C5714 a_83153_n36322.t14 VSS 0.458717f
C5715 a_83153_n36322.t19 VSS 0.45876f
C5716 a_83153_n36322.t7 VSS 0.260911f
C5717 a_83153_n36322.t10 VSS 0.452124f
C5718 a_83153_n36322.t13 VSS 0.452124f
C5719 a_83153_n36322.t18 VSS 0.450255f
C5720 a_83153_n36322.t8 VSS 0.450255f
C5721 a_83153_n36322.t21 VSS 0.45876f
C5722 a_83153_n36322.t23 VSS 0.450255f
C5723 a_83153_n36322.t15 VSS 0.450255f
C5724 a_83153_n36322.t22 VSS 0.452124f
C5725 a_83153_n36322.t9 VSS 0.450255f
C5726 a_83153_n36322.t20 VSS 0.452124f
C5727 a_83153_n36322.t16 VSS 0.450255f
C5728 a_83153_n36322.t12 VSS 0.458717f
C5729 a_83153_n36322.t17 VSS 0.450255f
C5730 a_83153_n36322.t11 VSS 0.450255f
C5731 a_83153_n36322.t3 VSS 0.410822f
C5732 a_83153_n36322.t1 VSS 0.242341f
C5733 a_83153_n36322.t0 VSS 0.273797f
C5734 a_83153_n36322.t2 VSS 0.423358f
C5735 a_83153_n36322.t6 VSS 0.39953f
C5736 a_83153_n36322.t5 VSS 0.50972f
C5737 a_83153_n36322.t4 VSS 0.278471f
C5738 a_84017_n17715.t2 VSS 62.4781f
C5739 a_84017_n17715.t3 VSS 0.430693f
C5740 a_84017_n17715.t0 VSS 0.847888f
C5741 a_84017_n17715.t1 VSS 0.715074f
C5742 a_84017_n17715.t4 VSS 34.528202f
C5743 a_83325_4421.t0 VSS 25.151001f
C5744 a_83325_4421.t1 VSS 13.2043f
C5745 a_83325_4421.t2 VSS 1.14464f
C5746 a_47819_n36322.n0 VSS 11.550099f
C5747 a_47819_n36322.n1 VSS 0.727598f
C5748 a_47819_n36322.n2 VSS 11.477901f
C5749 a_47819_n36322.t21 VSS 0.458717f
C5750 a_47819_n36322.t9 VSS 0.458761f
C5751 a_47819_n36322.t23 VSS 0.452124f
C5752 a_47819_n36322.t8 VSS 0.452124f
C5753 a_47819_n36322.t19 VSS 0.450255f
C5754 a_47819_n36322.t22 VSS 0.450255f
C5755 a_47819_n36322.t10 VSS 0.458761f
C5756 a_47819_n36322.t20 VSS 0.450255f
C5757 a_47819_n36322.t16 VSS 0.450255f
C5758 a_47819_n36322.t17 VSS 0.452124f
C5759 a_47819_n36322.t11 VSS 0.450255f
C5760 a_47819_n36322.t15 VSS 0.452124f
C5761 a_47819_n36322.t13 VSS 0.450255f
C5762 a_47819_n36322.t18 VSS 0.458717f
C5763 a_47819_n36322.t14 VSS 0.450255f
C5764 a_47819_n36322.t12 VSS 0.450255f
C5765 a_47819_n36322.t5 VSS 0.410822f
C5766 a_47819_n36322.t4 VSS 0.242342f
C5767 a_47819_n36322.t6 VSS 0.273797f
C5768 a_47819_n36322.t7 VSS 0.423358f
C5769 a_47819_n36322.t2 VSS 0.39953f
C5770 a_47819_n36322.t3 VSS 0.260911f
C5771 a_47819_n36322.t1 VSS 0.278471f
C5772 a_47819_n36322.t0 VSS 0.50972f
C5773 a_47819_10448.n0 VSS 7.87162f
C5774 a_47819_10448.n1 VSS 0.865678f
C5775 a_47819_10448.t1 VSS 13.622499f
C5776 a_47819_10448.t10 VSS 0.30485f
C5777 a_47819_10448.t3 VSS 0.568066f
C5778 a_47819_10448.t16 VSS 0.544019f
C5779 a_47819_10448.t19 VSS 0.568066f
C5780 a_47819_10448.t11 VSS 0.544019f
C5781 a_47819_10448.t14 VSS 0.544019f
C5782 a_47819_10448.t9 VSS 0.562597f
C5783 a_47819_10448.t12 VSS 0.562597f
C5784 a_47819_10448.t20 VSS 0.544019f
C5785 a_47819_10448.t15 VSS 0.568066f
C5786 a_47819_10448.t18 VSS 0.544019f
C5787 a_47819_10448.t6 VSS 0.34777f
C5788 a_47819_10448.t8 VSS 0.30485f
C5789 a_47819_10448.t2 VSS 0.330207f
C5790 a_47819_10448.t0 VSS 0.329925f
C5791 a_47819_10448.t7 VSS 0.562597f
C5792 a_47819_10448.t22 VSS 0.544019f
C5793 a_47819_10448.t5 VSS 0.568066f
C5794 a_47819_10448.t17 VSS 0.544019f
C5795 a_47819_10448.t13 VSS 0.562597f
C5796 a_47819_10448.t21 VSS 0.544019f
C5797 a_47819_10448.t4 VSS 0.34777f
C5798 a_112559_n29181.n0 VSS 4.20259f
C5799 a_112559_n29181.n1 VSS 4.03827f
C5800 a_112559_n29181.t1 VSS 3.66539f
C5801 a_112559_n29181.t4 VSS 0.178345f
C5802 a_112559_n29181.t6 VSS 0.153725f
C5803 a_112559_n29181.t3 VSS 0.298622f
C5804 a_112559_n29181.t18 VSS 0.285961f
C5805 a_112559_n29181.t21 VSS 0.295389f
C5806 a_112559_n29181.t20 VSS 0.298622f
C5807 a_112559_n29181.t15 VSS 0.285961f
C5808 a_112559_n29181.t14 VSS 0.298622f
C5809 a_112559_n29181.t12 VSS 0.285961f
C5810 a_112559_n29181.t7 VSS 0.295686f
C5811 a_112559_n29181.t13 VSS 0.285983f
C5812 a_112559_n29181.t10 VSS 0.178268f
C5813 a_112559_n29181.t8 VSS 0.153794f
C5814 a_112559_n29181.t9 VSS 0.298622f
C5815 a_112559_n29181.t22 VSS 0.285961f
C5816 a_112559_n29181.t16 VSS 0.295636f
C5817 a_112559_n29181.t11 VSS 0.285983f
C5818 a_112559_n29181.t17 VSS 0.285983f
C5819 a_112559_n29181.t5 VSS 0.295488f
C5820 a_112559_n29181.t19 VSS 0.285983f
C5821 a_112559_n29181.t2 VSS 0.182073f
C5822 a_112559_n29181.t0 VSS 0.183085f
C5823 a_30324_n29313.t0 VSS 23.414902f
C5824 a_30324_n29313.t2 VSS 8.917299f
C5825 a_30324_n29313.t1 VSS 7.66778f
C5826 a_56895_n16009.t0 VSS 50.790398f
C5827 a_56895_n16009.t1 VSS 36.409603f
C5828 a_83153_n35156.t10 VSS 20.5853f
C5829 a_83153_n35156.t11 VSS 1.77452f
C5830 a_83153_n35156.t5 VSS 0.304855f
C5831 a_83153_n35156.t8 VSS 0.330202f
C5832 a_83153_n35156.t9 VSS 0.329919f
C5833 a_83153_n35156.t0 VSS 0.568066f
C5834 a_83153_n35156.t13 VSS 0.544019f
C5835 a_83153_n35156.t12 VSS 0.544019f
C5836 a_83153_n35156.t22 VSS 0.562597f
C5837 a_83153_n35156.t21 VSS 0.568066f
C5838 a_83153_n35156.t19 VSS 0.544019f
C5839 a_83153_n35156.t4 VSS 0.562597f
C5840 a_83153_n35156.t17 VSS 0.544019f
C5841 a_83153_n35156.t6 VSS 0.568066f
C5842 a_83153_n35156.t15 VSS 0.544019f
C5843 a_83153_n35156.t7 VSS 0.347769f
C5844 a_83153_n35156.t3 VSS 0.304855f
C5845 a_83153_n35156.t23 VSS 0.562597f
C5846 a_83153_n35156.t14 VSS 0.544019f
C5847 a_83153_n35156.t20 VSS 0.568066f
C5848 a_83153_n35156.t18 VSS 0.544019f
C5849 a_83153_n35156.t2 VSS 0.562597f
C5850 a_83153_n35156.t16 VSS 0.544019f
C5851 a_83153_n35156.t1 VSS 0.347769f
C5852 a_89033_n35156.t10 VSS 0.906416f
C5853 a_89033_n35156.n0 VSS 11.033299f
C5854 a_89033_n35156.n1 VSS 4.04697f
C5855 a_89033_n35156.t9 VSS 0.924513f
C5856 a_89033_n35156.t8 VSS 0.829311f
C5857 a_89033_n35156.t6 VSS 0.829311f
C5858 a_89033_n35156.t11 VSS 0.880327f
C5859 a_89033_n35156.t7 VSS 0.829311f
C5860 a_89033_n35156.t5 VSS 0.829311f
C5861 a_89033_n35156.t12 VSS 0.81277f
C5862 a_89033_n35156.t3 VSS 0.623484f
C5863 a_89033_n35156.n2 VSS 0.90089f
C5864 a_89033_n35156.t4 VSS 3.71473f
C5865 a_89033_n35156.t2 VSS 0.237239f
C5866 a_89033_n35156.t1 VSS 0.230787f
C5867 a_89033_n35156.n3 VSS 62.454002f
C5868 a_89033_n35156.t0 VSS 19.6173f
C5869 a_96011_n36322.t2 VSS 2.81139f
C5870 a_96011_n36322.t1 VSS 67.4611f
C5871 a_96011_n36322.t3 VSS 1.68557f
C5872 a_96011_n36322.t0 VSS 27.042f
C5873 a_36008_4481.n0 VSS 9.956611f
C5874 a_36008_4481.t1 VSS 0.704006f
C5875 a_36008_4481.t0 VSS 0.606767f
C5876 a_36008_4481.t3 VSS 0.509963f
C5877 a_36008_4481.t2 VSS 0.92265f
C5878 a_30152_11614.n0 VSS 0.729765f
C5879 a_30152_11614.n1 VSS 11.5118f
C5880 a_30152_11614.n2 VSS 11.584201f
C5881 a_30152_11614.t8 VSS 0.460118f
C5882 a_30152_11614.t17 VSS 0.460074f
C5883 a_30152_11614.t15 VSS 0.453462f
C5884 a_30152_11614.t19 VSS 0.453462f
C5885 a_30152_11614.t18 VSS 0.451587f
C5886 a_30152_11614.t14 VSS 0.451587f
C5887 a_30152_11614.t13 VSS 0.451587f
C5888 a_30152_11614.t21 VSS 0.460118f
C5889 a_30152_11614.t16 VSS 0.451587f
C5890 a_30152_11614.t23 VSS 0.453462f
C5891 a_30152_11614.t12 VSS 0.453462f
C5892 a_30152_11614.t11 VSS 0.451587f
C5893 a_30152_11614.t22 VSS 0.451587f
C5894 a_30152_11614.t20 VSS 0.451587f
C5895 a_30152_11614.t9 VSS 0.460074f
C5896 a_30152_11614.t10 VSS 0.451587f
C5897 a_30152_11614.t0 VSS 0.412039f
C5898 a_30152_11614.t3 VSS 0.243046f
C5899 a_30152_11614.t2 VSS 0.274604f
C5900 a_30152_11614.t1 VSS 0.424622f
C5901 a_30152_11614.t7 VSS 0.400707f
C5902 a_30152_11614.t5 VSS 0.261684f
C5903 a_30152_11614.t6 VSS 0.279295f
C5904 a_30152_11614.t4 VSS 0.511245f
C5905 a_63161_n5344.t2 VSS 4.9628f
C5906 a_63161_n5344.t1 VSS 49.1395f
C5907 a_63161_n5344.t0 VSS 29.1977f
C5908 a_64243_n1756.t1 VSS 69.347206f
C5909 a_64243_n1756.t2 VSS 2.72276f
C5910 a_64243_n1756.t0 VSS 16.93f
C5911 a_77225_n29181.n0 VSS 4.17871f
C5912 a_77225_n29181.n1 VSS 4.01532f
C5913 a_77225_n29181.t9 VSS 3.64456f
C5914 a_77225_n29181.t5 VSS 0.177332f
C5915 a_77225_n29181.t1 VSS 0.152852f
C5916 a_77225_n29181.t4 VSS 0.296925f
C5917 a_77225_n29181.t12 VSS 0.284336f
C5918 a_77225_n29181.t18 VSS 0.293711f
C5919 a_77225_n29181.t19 VSS 0.296925f
C5920 a_77225_n29181.t11 VSS 0.284336f
C5921 a_77225_n29181.t15 VSS 0.296925f
C5922 a_77225_n29181.t20 VSS 0.284336f
C5923 a_77225_n29181.t2 VSS 0.294005f
C5924 a_77225_n29181.t16 VSS 0.284359f
C5925 a_77225_n29181.t7 VSS 0.177255f
C5926 a_77225_n29181.t3 VSS 0.152921f
C5927 a_77225_n29181.t6 VSS 0.296925f
C5928 a_77225_n29181.t17 VSS 0.284336f
C5929 a_77225_n29181.t13 VSS 0.293956f
C5930 a_77225_n29181.t14 VSS 0.284359f
C5931 a_77225_n29181.t21 VSS 0.284359f
C5932 a_77225_n29181.t0 VSS 0.293809f
C5933 a_77225_n29181.t22 VSS 0.284359f
C5934 a_77225_n29181.t10 VSS 0.181038f
C5935 a_77225_n29181.t8 VSS 0.182045f
C5936 a_94892_n29181.n0 VSS 4.17871f
C5937 a_94892_n29181.n1 VSS 4.01532f
C5938 a_94892_n29181.t9 VSS 3.64456f
C5939 a_94892_n29181.t3 VSS 0.177332f
C5940 a_94892_n29181.t7 VSS 0.152852f
C5941 a_94892_n29181.t2 VSS 0.296925f
C5942 a_94892_n29181.t19 VSS 0.284336f
C5943 a_94892_n29181.t16 VSS 0.293711f
C5944 a_94892_n29181.t22 VSS 0.296925f
C5945 a_94892_n29181.t17 VSS 0.284336f
C5946 a_94892_n29181.t18 VSS 0.296925f
C5947 a_94892_n29181.t13 VSS 0.284336f
C5948 a_94892_n29181.t4 VSS 0.294005f
C5949 a_94892_n29181.t15 VSS 0.284359f
C5950 a_94892_n29181.t1 VSS 0.177255f
C5951 a_94892_n29181.t5 VSS 0.152921f
C5952 a_94892_n29181.t0 VSS 0.296925f
C5953 a_94892_n29181.t12 VSS 0.284336f
C5954 a_94892_n29181.t11 VSS 0.293956f
C5955 a_94892_n29181.t14 VSS 0.284359f
C5956 a_94892_n29181.t20 VSS 0.284359f
C5957 a_94892_n29181.t6 VSS 0.293809f
C5958 a_94892_n29181.t21 VSS 0.284359f
C5959 a_94892_n29181.t10 VSS 0.182045f
C5960 a_94892_n29181.t8 VSS 0.181038f
C5961 a_83325_n29313.t0 VSS 23.122198f
C5962 a_83325_n29313.t1 VSS 8.80583f
C5963 a_83325_n29313.t2 VSS 7.57194f
C5964 a_53699_n35156.t10 VSS 0.964284f
C5965 a_53699_n35156.n0 VSS 11.7377f
C5966 a_53699_n35156.n1 VSS 4.30534f
C5967 a_53699_n35156.t9 VSS 0.983536f
C5968 a_53699_n35156.t8 VSS 0.882256f
C5969 a_53699_n35156.t12 VSS 0.882256f
C5970 a_53699_n35156.t5 VSS 0.936529f
C5971 a_53699_n35156.t7 VSS 0.882256f
C5972 a_53699_n35156.t11 VSS 0.882256f
C5973 a_53699_n35156.t6 VSS 0.864658f
C5974 a_53699_n35156.t4 VSS 0.663289f
C5975 a_53699_n35156.n2 VSS 0.958405f
C5976 a_53699_n35156.t3 VSS 3.95189f
C5977 a_53699_n35156.t1 VSS 0.252384f
C5978 a_53699_n35156.t2 VSS 0.245521f
C5979 a_53699_n35156.n3 VSS 51.853f
C5980 a_53699_n35156.t0 VSS 20.954401f
C5981 a_59558_4481.n0 VSS 0.449404f
C5982 a_59558_4481.n1 VSS 7.74464f
C5983 a_59558_4481.t2 VSS 3.64456f
C5984 a_59558_4481.t6 VSS 0.177333f
C5985 a_59558_4481.t4 VSS 0.152849f
C5986 a_59558_4481.t5 VSS 0.296925f
C5987 a_59558_4481.t22 VSS 0.284336f
C5988 a_59558_4481.t18 VSS 0.293711f
C5989 a_59558_4481.t14 VSS 0.296925f
C5990 a_59558_4481.t20 VSS 0.284336f
C5991 a_59558_4481.t19 VSS 0.296925f
C5992 a_59558_4481.t11 VSS 0.284336f
C5993 a_59558_4481.t9 VSS 0.294005f
C5994 a_59558_4481.t21 VSS 0.284359f
C5995 a_59558_4481.t8 VSS 0.177256f
C5996 a_59558_4481.t10 VSS 0.152918f
C5997 a_59558_4481.t7 VSS 0.296925f
C5998 a_59558_4481.t16 VSS 0.284336f
C5999 a_59558_4481.t13 VSS 0.293956f
C6000 a_59558_4481.t12 VSS 0.284359f
C6001 a_59558_4481.t15 VSS 0.284359f
C6002 a_59558_4481.t3 VSS 0.293809f
C6003 a_59558_4481.t17 VSS 0.284359f
C6004 a_59558_4481.t1 VSS 0.181041f
C6005 a_59558_4481.t0 VSS 0.182047f
C6006 a_39179_n19595.t0 VSS 72.542206f
C6007 a_39179_n19595.t2 VSS 2.69368f
C6008 a_39179_n19595.t1 VSS 13.8641f
C6009 a_78344_n36322.t3 VSS 3.04902f
C6010 a_78344_n36322.t2 VSS 61.7295f
C6011 a_78344_n36322.t1 VSS 1.82803f
C6012 a_78344_n36322.t0 VSS 24.293499f
C6013 a_71366_n35156.t7 VSS 0.960498f
C6014 a_71366_n35156.n0 VSS 11.6917f
C6015 a_71366_n35156.n1 VSS 4.28844f
C6016 a_71366_n35156.t6 VSS 0.979675f
C6017 a_71366_n35156.t11 VSS 0.878792f
C6018 a_71366_n35156.t9 VSS 0.878792f
C6019 a_71366_n35156.t12 VSS 0.932853f
C6020 a_71366_n35156.t10 VSS 0.878792f
C6021 a_71366_n35156.t8 VSS 0.878792f
C6022 a_71366_n35156.t5 VSS 0.861264f
C6023 a_71366_n35156.t2 VSS 0.660685f
C6024 a_71366_n35156.n2 VSS 0.954642f
C6025 a_71366_n35156.t4 VSS 3.93638f
C6026 a_71366_n35156.t3 VSS 0.251394f
C6027 a_71366_n35156.t1 VSS 0.244558f
C6028 a_71366_n35156.n3 VSS 57.0977f
C6029 a_71366_n35156.t0 VSS 16.425098f
C6030 a_44363_n16007.t1 VSS 6.93736f
C6031 a_44363_n16007.t2 VSS 50.117397f
C6032 a_44363_n16007.t0 VSS 26.445198f
C6033 a_53699_n36322.t3 VSS 0.781529f
C6034 a_53699_n36322.t2 VSS 0.752866f
C6035 a_53699_n36322.n0 VSS 8.13798f
C6036 a_53699_n36322.t1 VSS 0.676033f
C6037 a_53699_n36322.n1 VSS 8.25899f
C6038 a_53699_n36322.t0 VSS 0.792603f
C6039 a_71496_n36382.n0 VSS 2.53786f
C6040 a_71496_n36382.n1 VSS 9.92737f
C6041 a_71496_n36382.n2 VSS 0.941684f
C6042 a_71496_n36382.n3 VSS 1.60401f
C6043 a_71496_n36382.n4 VSS 5.88446f
C6044 a_71496_n36382.n5 VSS 7.95021f
C6045 a_71496_n36382.n6 VSS 0.911784f
C6046 a_71496_n36382.t12 VSS 0.572572f
C6047 a_71496_n36382.t13 VSS 0.605718f
C6048 a_71496_n36382.t21 VSS 0.572368f
C6049 a_71496_n36382.t6 VSS 0.315898f
C6050 a_71496_n36382.t1 VSS 0.599022f
C6051 a_71496_n36382.t3 VSS 0.321538f
C6052 a_71496_n36382.t0 VSS 0.32663f
C6053 a_71496_n36382.t2 VSS 0.49853f
C6054 a_71496_n36382.t7 VSS 0.52604f
C6055 a_71496_n36382.t18 VSS 0.563936f
C6056 a_71496_n36382.t11 VSS 0.563895f
C6057 a_71496_n36382.t15 VSS 0.561709f
C6058 a_71496_n36382.t22 VSS 0.561709f
C6059 a_71496_n36382.t16 VSS 0.561709f
C6060 a_71496_n36382.t20 VSS 0.561709f
C6061 a_71496_n36382.t23 VSS 0.563801f
C6062 a_71496_n36382.t10 VSS 0.563957f
C6063 a_71496_n36382.t14 VSS 0.561709f
C6064 a_71496_n36382.t9 VSS 0.561709f
C6065 a_71496_n36382.t17 VSS 0.561709f
C6066 a_71496_n36382.t8 VSS 0.571948f
C6067 a_71496_n36382.t19 VSS 0.561709f
C6068 a_71496_n36382.t5 VSS 0.523325f
C6069 a_71496_n36382.n7 VSS 0.912668f
C6070 a_71496_n36382.t4 VSS 0.347078f
C6071 a_89009_n27257.n0 VSS 9.95669f
C6072 a_89009_n27257.t3 VSS 0.704006f
C6073 a_89009_n27257.t2 VSS 0.606767f
C6074 a_89009_n27257.t1 VSS 0.922584f
C6075 a_89009_n27257.t0 VSS 0.509953f
C6076 a_41891_n29181.t0 VSS 3.64456f
C6077 a_41891_n29181.n0 VSS 4.17871f
C6078 a_41891_n29181.n1 VSS 4.01532f
C6079 a_41891_n29181.t8 VSS 0.177332f
C6080 a_41891_n29181.t6 VSS 0.152852f
C6081 a_41891_n29181.t7 VSS 0.296925f
C6082 a_41891_n29181.t15 VSS 0.284336f
C6083 a_41891_n29181.t12 VSS 0.293711f
C6084 a_41891_n29181.t18 VSS 0.296925f
C6085 a_41891_n29181.t13 VSS 0.284336f
C6086 a_41891_n29181.t14 VSS 0.296925f
C6087 a_41891_n29181.t21 VSS 0.284336f
C6088 a_41891_n29181.t3 VSS 0.294005f
C6089 a_41891_n29181.t11 VSS 0.284359f
C6090 a_41891_n29181.t10 VSS 0.177255f
C6091 a_41891_n29181.t4 VSS 0.152921f
C6092 a_41891_n29181.t9 VSS 0.296925f
C6093 a_41891_n29181.t20 VSS 0.284336f
C6094 a_41891_n29181.t19 VSS 0.293956f
C6095 a_41891_n29181.t22 VSS 0.284359f
C6096 a_41891_n29181.t16 VSS 0.284359f
C6097 a_41891_n29181.t5 VSS 0.293809f
C6098 a_41891_n29181.t17 VSS 0.284359f
C6099 a_41891_n29181.t1 VSS 0.182045f
C6100 a_41891_n29181.t2 VSS 0.181038f
C6101 a_106809_n5150.t1 VSS 1.82106f
C6102 a_106809_n5150.t2 VSS 39.9196f
C6103 a_106809_n5150.t3 VSS 1.09181f
C6104 a_106809_n5150.t0 VSS 21.667599f
C6105 a_89163_n36382.n0 VSS 2.53786f
C6106 a_89163_n36382.n1 VSS 9.92737f
C6107 a_89163_n36382.n2 VSS 0.941685f
C6108 a_89163_n36382.n3 VSS 1.60401f
C6109 a_89163_n36382.n4 VSS 5.88446f
C6110 a_89163_n36382.n5 VSS 7.95021f
C6111 a_89163_n36382.n6 VSS 0.911784f
C6112 a_89163_n36382.t20 VSS 0.572572f
C6113 a_89163_n36382.t21 VSS 0.605718f
C6114 a_89163_n36382.t15 VSS 0.572369f
C6115 a_89163_n36382.t2 VSS 0.315898f
C6116 a_89163_n36382.t6 VSS 0.599022f
C6117 a_89163_n36382.t7 VSS 0.321538f
C6118 a_89163_n36382.t4 VSS 0.32663f
C6119 a_89163_n36382.t5 VSS 0.49853f
C6120 a_89163_n36382.t3 VSS 0.52604f
C6121 a_89163_n36382.t10 VSS 0.563936f
C6122 a_89163_n36382.t13 VSS 0.563895f
C6123 a_89163_n36382.t9 VSS 0.561709f
C6124 a_89163_n36382.t22 VSS 0.561709f
C6125 a_89163_n36382.t14 VSS 0.561709f
C6126 a_89163_n36382.t19 VSS 0.561709f
C6127 a_89163_n36382.t11 VSS 0.563801f
C6128 a_89163_n36382.t12 VSS 0.563957f
C6129 a_89163_n36382.t8 VSS 0.561709f
C6130 a_89163_n36382.t23 VSS 0.561709f
C6131 a_89163_n36382.t16 VSS 0.561709f
C6132 a_89163_n36382.t17 VSS 0.571948f
C6133 a_89163_n36382.t18 VSS 0.561709f
C6134 a_89163_n36382.t1 VSS 0.523326f
C6135 a_89163_n36382.n7 VSS 0.912668f
C6136 a_89163_n36382.t0 VSS 0.347078f
C6137 a_81205_n14095.n0 VSS 10.8627f
C6138 a_81205_n14095.t0 VSS 60.3566f
C6139 a_81205_n14095.t9 VSS 0.892387f
C6140 a_81205_n14095.n1 VSS 3.98441f
C6141 a_81205_n14095.t1 VSS 0.868961f
C6142 a_81205_n14095.t10 VSS 0.9102f
C6143 a_81205_n14095.t4 VSS 0.816488f
C6144 a_81205_n14095.t8 VSS 0.816488f
C6145 a_81205_n14095.t6 VSS 0.866731f
C6146 a_81205_n14095.t7 VSS 0.816488f
C6147 a_81205_n14095.t3 VSS 0.816488f
C6148 a_81205_n14095.t5 VSS 0.800202f
C6149 a_81205_n14095.t2 VSS 26.191801f
C6150 a_43010_10448.t2 VSS 3.0792f
C6151 a_43010_10448.t0 VSS 49.849697f
C6152 a_43010_10448.t1 VSS 0.941624f
C6153 a_43010_10448.t3 VSS 0.280444f
C6154 a_43010_10448.t4 VSS 36.6491f
C6155 a_36032_11614.n0 VSS 11.817201f
C6156 a_36032_11614.t0 VSS 50.134502f
C6157 a_36032_11614.t7 VSS 0.970796f
C6158 a_36032_11614.n1 VSS 4.3345f
C6159 a_36032_11614.t1 VSS 0.945312f
C6160 a_36032_11614.t8 VSS 0.990174f
C6161 a_36032_11614.t10 VSS 0.888228f
C6162 a_36032_11614.t6 VSS 0.888228f
C6163 a_36032_11614.t4 VSS 0.942885f
C6164 a_36032_11614.t5 VSS 0.888228f
C6165 a_36032_11614.t9 VSS 0.888228f
C6166 a_36032_11614.t3 VSS 0.870512f
C6167 a_36032_11614.t2 VSS 27.941301f
C6168 a_65486_10448.n0 VSS 7.87162f
C6169 a_65486_10448.n1 VSS 0.865678f
C6170 a_65486_10448.t10 VSS 13.622499f
C6171 a_65486_10448.t3 VSS 0.34777f
C6172 a_65486_10448.t2 VSS 0.568066f
C6173 a_65486_10448.t11 VSS 0.544019f
C6174 a_65486_10448.t19 VSS 0.568066f
C6175 a_65486_10448.t15 VSS 0.544019f
C6176 a_65486_10448.t14 VSS 0.544019f
C6177 a_65486_10448.t0 VSS 0.562597f
C6178 a_65486_10448.t17 VSS 0.562597f
C6179 a_65486_10448.t20 VSS 0.544019f
C6180 a_65486_10448.t16 VSS 0.568066f
C6181 a_65486_10448.t13 VSS 0.544019f
C6182 a_65486_10448.t7 VSS 0.34777f
C6183 a_65486_10448.t5 VSS 0.30485f
C6184 a_65486_10448.t9 VSS 0.330207f
C6185 a_65486_10448.t8 VSS 0.329925f
C6186 a_65486_10448.t4 VSS 0.562597f
C6187 a_65486_10448.t22 VSS 0.544019f
C6188 a_65486_10448.t6 VSS 0.568066f
C6189 a_65486_10448.t12 VSS 0.544019f
C6190 a_65486_10448.t18 VSS 0.562597f
C6191 a_65486_10448.t21 VSS 0.544019f
C6192 a_65486_10448.t1 VSS 0.30485f
C6193 a_89033_13546.t2 VSS 0.764004f
C6194 a_89033_13546.t3 VSS 0.65164f
C6195 a_89033_13546.n0 VSS 7.959681f
C6196 a_89033_13546.t1 VSS 0.753329f
C6197 a_89033_13546.n1 VSS 7.84565f
C6198 a_89033_13546.t0 VSS 0.725701f
C6199 a_89163_10388.n0 VSS 2.53786f
C6200 a_89163_10388.n1 VSS 9.92737f
C6201 a_89163_10388.n2 VSS 0.941685f
C6202 a_89163_10388.n3 VSS 1.60401f
C6203 a_89163_10388.n4 VSS 0.912682f
C6204 a_89163_10388.n5 VSS 5.88445f
C6205 a_89163_10388.n6 VSS 7.950201f
C6206 a_89163_10388.n7 VSS 0.911776f
C6207 a_89163_10388.t23 VSS 0.572368f
C6208 a_89163_10388.t15 VSS 0.572572f
C6209 a_89163_10388.t10 VSS 0.605719f
C6210 a_89163_10388.t22 VSS 0.571949f
C6211 a_89163_10388.t9 VSS 0.563936f
C6212 a_89163_10388.t11 VSS 0.563895f
C6213 a_89163_10388.t21 VSS 0.561709f
C6214 a_89163_10388.t16 VSS 0.561709f
C6215 a_89163_10388.t14 VSS 0.561709f
C6216 a_89163_10388.t20 VSS 0.561709f
C6217 a_89163_10388.t8 VSS 0.563801f
C6218 a_89163_10388.t17 VSS 0.563957f
C6219 a_89163_10388.t19 VSS 0.561709f
C6220 a_89163_10388.t13 VSS 0.561709f
C6221 a_89163_10388.t18 VSS 0.561709f
C6222 a_89163_10388.t12 VSS 0.561709f
C6223 a_89163_10388.t6 VSS 0.523342f
C6224 a_89163_10388.t5 VSS 0.315882f
C6225 a_89163_10388.t7 VSS 0.347081f
C6226 a_89163_10388.t3 VSS 0.599013f
C6227 a_89163_10388.t1 VSS 0.321546f
C6228 a_89163_10388.t0 VSS 0.32663f
C6229 a_89163_10388.t2 VSS 0.498545f
C6230 a_89163_10388.t4 VSS 0.526042f
C6231 a_30152_n35156.t8 VSS 20.5853f
C6232 a_30152_n35156.t11 VSS 1.77452f
C6233 a_30152_n35156.t3 VSS 0.304855f
C6234 a_30152_n35156.t9 VSS 0.330202f
C6235 a_30152_n35156.t10 VSS 0.329919f
C6236 a_30152_n35156.t0 VSS 0.568066f
C6237 a_30152_n35156.t22 VSS 0.544019f
C6238 a_30152_n35156.t21 VSS 0.544019f
C6239 a_30152_n35156.t19 VSS 0.562597f
C6240 a_30152_n35156.t18 VSS 0.568066f
C6241 a_30152_n35156.t16 VSS 0.544019f
C6242 a_30152_n35156.t2 VSS 0.562597f
C6243 a_30152_n35156.t14 VSS 0.544019f
C6244 a_30152_n35156.t6 VSS 0.568066f
C6245 a_30152_n35156.t12 VSS 0.544019f
C6246 a_30152_n35156.t7 VSS 0.347769f
C6247 a_30152_n35156.t5 VSS 0.304855f
C6248 a_30152_n35156.t20 VSS 0.562597f
C6249 a_30152_n35156.t23 VSS 0.544019f
C6250 a_30152_n35156.t17 VSS 0.568066f
C6251 a_30152_n35156.t15 VSS 0.544019f
C6252 a_30152_n35156.t4 VSS 0.562597f
C6253 a_30152_n35156.t13 VSS 0.544019f
C6254 a_30152_n35156.t1 VSS 0.347769f
C6255 a_36032_n35156.t12 VSS 0.968935f
C6256 a_36032_n35156.n0 VSS 11.7943f
C6257 a_36032_n35156.n1 VSS 4.3261f
C6258 a_36032_n35156.t11 VSS 0.98828f
C6259 a_36032_n35156.t10 VSS 0.886511f
C6260 a_36032_n35156.t8 VSS 0.886511f
C6261 a_36032_n35156.t5 VSS 0.941046f
C6262 a_36032_n35156.t9 VSS 0.886511f
C6263 a_36032_n35156.t7 VSS 0.886511f
C6264 a_36032_n35156.t6 VSS 0.868829f
C6265 a_36032_n35156.t2 VSS 0.666488f
C6266 a_36032_n35156.n2 VSS 0.963028f
C6267 a_36032_n35156.t1 VSS 3.97095f
C6268 a_36032_n35156.t4 VSS 0.253602f
C6269 a_36032_n35156.t3 VSS 0.246706f
C6270 a_36032_n35156.n3 VSS 47.1512f
C6271 a_36032_n35156.t0 VSS 25.5144f
C6272 a_106676_4481.n0 VSS 9.95668f
C6273 a_106676_4481.t3 VSS 0.922601f
C6274 a_106676_4481.t1 VSS 0.704006f
C6275 a_106676_4481.t0 VSS 0.606767f
C6276 a_106676_4481.t2 VSS 0.50995f
C6277 a_106830_10388.n0 VSS 2.51436f
C6278 a_106830_10388.n1 VSS 9.83545f
C6279 a_106830_10388.n2 VSS 0.932966f
C6280 a_106830_10388.n3 VSS 1.58916f
C6281 a_106830_10388.n4 VSS 0.904231f
C6282 a_106830_10388.n5 VSS 5.82997f
C6283 a_106830_10388.n6 VSS 7.87659f
C6284 a_106830_10388.n7 VSS 0.903334f
C6285 a_106830_10388.t20 VSS 0.567068f
C6286 a_106830_10388.t12 VSS 0.567271f
C6287 a_106830_10388.t22 VSS 0.60011f
C6288 a_106830_10388.t19 VSS 0.566653f
C6289 a_106830_10388.t15 VSS 0.558714f
C6290 a_106830_10388.t17 VSS 0.558674f
C6291 a_106830_10388.t8 VSS 0.556508f
C6292 a_106830_10388.t11 VSS 0.556508f
C6293 a_106830_10388.t10 VSS 0.556508f
C6294 a_106830_10388.t23 VSS 0.556508f
C6295 a_106830_10388.t14 VSS 0.558581f
C6296 a_106830_10388.t18 VSS 0.558735f
C6297 a_106830_10388.t21 VSS 0.556508f
C6298 a_106830_10388.t9 VSS 0.556508f
C6299 a_106830_10388.t16 VSS 0.556508f
C6300 a_106830_10388.t13 VSS 0.556508f
C6301 a_106830_10388.t7 VSS 0.593467f
C6302 a_106830_10388.t6 VSS 0.318569f
C6303 a_106830_10388.t5 VSS 0.323606f
C6304 a_106830_10388.t4 VSS 0.493929f
C6305 a_106830_10388.t2 VSS 0.521171f
C6306 a_106830_10388.t3 VSS 0.312957f
C6307 a_106830_10388.t1 VSS 0.343867f
C6308 a_106830_10388.t0 VSS 0.518497f
C6309 a_77225_4481.t8 VSS 3.64456f
C6310 a_77225_4481.n0 VSS 0.449404f
C6311 a_77225_4481.n1 VSS 7.74464f
C6312 a_77225_4481.t10 VSS 0.182047f
C6313 a_77225_4481.t7 VSS 0.177333f
C6314 a_77225_4481.t5 VSS 0.152849f
C6315 a_77225_4481.t6 VSS 0.296925f
C6316 a_77225_4481.t14 VSS 0.284336f
C6317 a_77225_4481.t11 VSS 0.293711f
C6318 a_77225_4481.t13 VSS 0.296925f
C6319 a_77225_4481.t12 VSS 0.284336f
C6320 a_77225_4481.t16 VSS 0.296925f
C6321 a_77225_4481.t15 VSS 0.284336f
C6322 a_77225_4481.t2 VSS 0.294005f
C6323 a_77225_4481.t21 VSS 0.284359f
C6324 a_77225_4481.t1 VSS 0.177256f
C6325 a_77225_4481.t3 VSS 0.152918f
C6326 a_77225_4481.t0 VSS 0.296925f
C6327 a_77225_4481.t22 VSS 0.284336f
C6328 a_77225_4481.t19 VSS 0.293956f
C6329 a_77225_4481.t17 VSS 0.284359f
C6330 a_77225_4481.t18 VSS 0.284359f
C6331 a_77225_4481.t4 VSS 0.293809f
C6332 a_77225_4481.t20 VSS 0.284359f
C6333 a_77225_4481.t9 VSS 0.181041f
C6334 a_100820_n35156.n0 VSS 7.87162f
C6335 a_100820_n35156.n1 VSS 0.865673f
C6336 a_100820_n35156.t1 VSS 13.622499f
C6337 a_100820_n35156.t6 VSS 0.304855f
C6338 a_100820_n35156.t3 VSS 0.568066f
C6339 a_100820_n35156.t14 VSS 0.544019f
C6340 a_100820_n35156.t18 VSS 0.544019f
C6341 a_100820_n35156.t12 VSS 0.562597f
C6342 a_100820_n35156.t7 VSS 0.568066f
C6343 a_100820_n35156.t13 VSS 0.544019f
C6344 a_100820_n35156.t0 VSS 0.330202f
C6345 a_100820_n35156.t2 VSS 0.329919f
C6346 a_100820_n35156.t20 VSS 0.568066f
C6347 a_100820_n35156.t16 VSS 0.544019f
C6348 a_100820_n35156.t22 VSS 0.544019f
C6349 a_100820_n35156.t9 VSS 0.562597f
C6350 a_100820_n35156.t8 VSS 0.347769f
C6351 a_100820_n35156.t10 VSS 0.304855f
C6352 a_100820_n35156.t11 VSS 0.562597f
C6353 a_100820_n35156.t17 VSS 0.544019f
C6354 a_100820_n35156.t19 VSS 0.568066f
C6355 a_100820_n35156.t15 VSS 0.544019f
C6356 a_100820_n35156.t5 VSS 0.562597f
C6357 a_100820_n35156.t21 VSS 0.544019f
C6358 a_100820_n35156.t4 VSS 0.347769f
C6359 a_51711_n12421.t0 VSS 63.9549f
C6360 a_51711_n12421.t2 VSS 2.46089f
C6361 a_51711_n12421.t1 VSS 26.9842f
C6362 a_47819_n35156.n0 VSS 7.87162f
C6363 a_47819_n35156.n1 VSS 0.865673f
C6364 a_47819_n35156.t8 VSS 13.622499f
C6365 a_47819_n35156.t3 VSS 0.304855f
C6366 a_47819_n35156.t0 VSS 0.568066f
C6367 a_47819_n35156.t16 VSS 0.544019f
C6368 a_47819_n35156.t22 VSS 0.544019f
C6369 a_47819_n35156.t21 VSS 0.562597f
C6370 a_47819_n35156.t4 VSS 0.568066f
C6371 a_47819_n35156.t15 VSS 0.544019f
C6372 a_47819_n35156.t9 VSS 0.330202f
C6373 a_47819_n35156.t10 VSS 0.329919f
C6374 a_47819_n35156.t12 VSS 0.568066f
C6375 a_47819_n35156.t18 VSS 0.544019f
C6376 a_47819_n35156.t14 VSS 0.544019f
C6377 a_47819_n35156.t6 VSS 0.562597f
C6378 a_47819_n35156.t5 VSS 0.347769f
C6379 a_47819_n35156.t7 VSS 0.304855f
C6380 a_47819_n35156.t19 VSS 0.562597f
C6381 a_47819_n35156.t20 VSS 0.544019f
C6382 a_47819_n35156.t11 VSS 0.568066f
C6383 a_47819_n35156.t17 VSS 0.544019f
C6384 a_47819_n35156.t2 VSS 0.562597f
C6385 a_47819_n35156.t13 VSS 0.544019f
C6386 a_47819_n35156.t1 VSS 0.347769f
C6387 a_30152_n36322.n0 VSS 11.584201f
C6388 a_30152_n36322.n1 VSS 0.72975f
C6389 a_30152_n36322.n2 VSS 11.5119f
C6390 a_30152_n36322.t12 VSS 0.460074f
C6391 a_30152_n36322.t16 VSS 0.460118f
C6392 a_30152_n36322.t7 VSS 0.279295f
C6393 a_30152_n36322.t18 VSS 0.453462f
C6394 a_30152_n36322.t21 VSS 0.453462f
C6395 a_30152_n36322.t9 VSS 0.451587f
C6396 a_30152_n36322.t23 VSS 0.451587f
C6397 a_30152_n36322.t19 VSS 0.460118f
C6398 a_30152_n36322.t22 VSS 0.451587f
C6399 a_30152_n36322.t8 VSS 0.451587f
C6400 a_30152_n36322.t13 VSS 0.453462f
C6401 a_30152_n36322.t17 VSS 0.451587f
C6402 a_30152_n36322.t11 VSS 0.453462f
C6403 a_30152_n36322.t14 VSS 0.451587f
C6404 a_30152_n36322.t10 VSS 0.460074f
C6405 a_30152_n36322.t15 VSS 0.451587f
C6406 a_30152_n36322.t20 VSS 0.451587f
C6407 a_30152_n36322.t4 VSS 0.412038f
C6408 a_30152_n36322.t1 VSS 0.243058f
C6409 a_30152_n36322.t2 VSS 0.274607f
C6410 a_30152_n36322.t3 VSS 0.42461f
C6411 a_30152_n36322.t6 VSS 0.400712f
C6412 a_30152_n36322.t5 VSS 0.511228f
C6413 a_30152_n36322.t0 VSS 0.261683f
C6414 a_112559_4481.n0 VSS 0.451972f
C6415 a_112559_4481.n1 VSS 7.78889f
C6416 a_112559_4481.t1 VSS 3.66538f
C6417 a_112559_4481.t2 VSS 0.183088f
C6418 a_112559_4481.t8 VSS 0.178346f
C6419 a_112559_4481.t10 VSS 0.153723f
C6420 a_112559_4481.t7 VSS 0.298622f
C6421 a_112559_4481.t20 VSS 0.285961f
C6422 a_112559_4481.t15 VSS 0.295389f
C6423 a_112559_4481.t12 VSS 0.298622f
C6424 a_112559_4481.t18 VSS 0.285961f
C6425 a_112559_4481.t17 VSS 0.298622f
C6426 a_112559_4481.t21 VSS 0.285961f
C6427 a_112559_4481.t3 VSS 0.295686f
C6428 a_112559_4481.t19 VSS 0.285983f
C6429 a_112559_4481.t6 VSS 0.178268f
C6430 a_112559_4481.t4 VSS 0.153791f
C6431 a_112559_4481.t5 VSS 0.298622f
C6432 a_112559_4481.t14 VSS 0.285961f
C6433 a_112559_4481.t22 VSS 0.295636f
C6434 a_112559_4481.t11 VSS 0.285983f
C6435 a_112559_4481.t13 VSS 0.285983f
C6436 a_112559_4481.t9 VSS 0.295488f
C6437 a_112559_4481.t16 VSS 0.285983f
C6438 a_112559_4481.t0 VSS 0.182075f
C6439 a_89715_n17715.t3 VSS 0.546172f
C6440 a_89715_n17715.t4 VSS 0.322785f
C6441 a_89715_n17715.t1 VSS 36.1967f
C6442 a_89715_n17715.t2 VSS 0.460619f
C6443 a_89715_n17715.t5 VSS 26.2963f
C6444 a_89715_n17715.t0 VSS 0.277433f
C6445 a_86903_n14095.n0 VSS 10.9263f
C6446 a_86903_n14095.t0 VSS 55.2877f
C6447 a_86903_n14095.t4 VSS 0.897611f
C6448 a_86903_n14095.n1 VSS 4.00774f
C6449 a_86903_n14095.t1 VSS 0.874049f
C6450 a_86903_n14095.t5 VSS 0.915529f
C6451 a_86903_n14095.t7 VSS 0.821268f
C6452 a_86903_n14095.t3 VSS 0.821268f
C6453 a_86903_n14095.t10 VSS 0.871805f
C6454 a_86903_n14095.t8 VSS 0.821268f
C6455 a_86903_n14095.t6 VSS 0.821268f
C6456 a_86903_n14095.t9 VSS 0.804887f
C6457 a_86903_n14095.t2 VSS 32.2293f
C6458 a_83153_11614.n0 VSS 0.727613f
C6459 a_83153_11614.n1 VSS 11.477901f
C6460 a_83153_11614.n2 VSS 11.550099f
C6461 a_83153_11614.t17 VSS 0.458761f
C6462 a_83153_11614.t8 VSS 0.458717f
C6463 a_83153_11614.t6 VSS 0.509737f
C6464 a_83153_11614.t5 VSS 0.260912f
C6465 a_83153_11614.t7 VSS 0.278471f
C6466 a_83153_11614.t10 VSS 0.452124f
C6467 a_83153_11614.t14 VSS 0.452124f
C6468 a_83153_11614.t12 VSS 0.450255f
C6469 a_83153_11614.t9 VSS 0.450255f
C6470 a_83153_11614.t20 VSS 0.450255f
C6471 a_83153_11614.t13 VSS 0.458761f
C6472 a_83153_11614.t23 VSS 0.450255f
C6473 a_83153_11614.t16 VSS 0.452124f
C6474 a_83153_11614.t22 VSS 0.452124f
C6475 a_83153_11614.t21 VSS 0.450255f
C6476 a_83153_11614.t15 VSS 0.450255f
C6477 a_83153_11614.t11 VSS 0.450255f
C6478 a_83153_11614.t18 VSS 0.458717f
C6479 a_83153_11614.t19 VSS 0.450255f
C6480 a_83153_11614.t0 VSS 0.410824f
C6481 a_83153_11614.t1 VSS 0.242329f
C6482 a_83153_11614.t3 VSS 0.273794f
C6483 a_83153_11614.t2 VSS 0.423369f
C6484 a_83153_11614.t4 VSS 0.399525f
C6485 a_106676_n30339.n0 VSS 10.6245f
C6486 a_106676_n30339.t1 VSS 0.843931f
C6487 a_106676_n30339.t0 VSS 0.685986f
C6488 a_106676_n30339.t3 VSS 0.812605f
C6489 a_106676_n30339.t2 VSS 0.632986f
C6490 a_100820_n36322.n0 VSS 11.550099f
C6491 a_100820_n36322.n1 VSS 0.727597f
C6492 a_100820_n36322.n2 VSS 11.477901f
C6493 a_100820_n36322.t8 VSS 0.458717f
C6494 a_100820_n36322.t12 VSS 0.45876f
C6495 a_100820_n36322.t2 VSS 0.260911f
C6496 a_100820_n36322.t10 VSS 0.452124f
C6497 a_100820_n36322.t11 VSS 0.452124f
C6498 a_100820_n36322.t22 VSS 0.450255f
C6499 a_100820_n36322.t9 VSS 0.450255f
C6500 a_100820_n36322.t13 VSS 0.45876f
C6501 a_100820_n36322.t23 VSS 0.450255f
C6502 a_100820_n36322.t19 VSS 0.450255f
C6503 a_100820_n36322.t20 VSS 0.452124f
C6504 a_100820_n36322.t14 VSS 0.450255f
C6505 a_100820_n36322.t18 VSS 0.452124f
C6506 a_100820_n36322.t16 VSS 0.450255f
C6507 a_100820_n36322.t21 VSS 0.458717f
C6508 a_100820_n36322.t17 VSS 0.450255f
C6509 a_100820_n36322.t15 VSS 0.450255f
C6510 a_100820_n36322.t5 VSS 0.410822f
C6511 a_100820_n36322.t6 VSS 0.242341f
C6512 a_100820_n36322.t4 VSS 0.273797f
C6513 a_100820_n36322.t7 VSS 0.423358f
C6514 a_100820_n36322.t3 VSS 0.39953f
C6515 a_100820_n36322.t1 VSS 0.50972f
C6516 a_100820_n36322.t0 VSS 0.278471f
C6517 a_65486_n35156.t8 VSS 20.5853f
C6518 a_65486_n35156.t11 VSS 1.77452f
C6519 a_65486_n35156.t7 VSS 0.304855f
C6520 a_65486_n35156.t10 VSS 0.330202f
C6521 a_65486_n35156.t9 VSS 0.329919f
C6522 a_65486_n35156.t0 VSS 0.568066f
C6523 a_65486_n35156.t17 VSS 0.544019f
C6524 a_65486_n35156.t23 VSS 0.544019f
C6525 a_65486_n35156.t21 VSS 0.562597f
C6526 a_65486_n35156.t14 VSS 0.568066f
C6527 a_65486_n35156.t20 VSS 0.544019f
C6528 a_65486_n35156.t6 VSS 0.562597f
C6529 a_65486_n35156.t16 VSS 0.544019f
C6530 a_65486_n35156.t2 VSS 0.568066f
C6531 a_65486_n35156.t18 VSS 0.544019f
C6532 a_65486_n35156.t3 VSS 0.347769f
C6533 a_65486_n35156.t5 VSS 0.304855f
C6534 a_65486_n35156.t22 VSS 0.562597f
C6535 a_65486_n35156.t12 VSS 0.544019f
C6536 a_65486_n35156.t13 VSS 0.568066f
C6537 a_65486_n35156.t19 VSS 0.544019f
C6538 a_65486_n35156.t4 VSS 0.562597f
C6539 a_65486_n35156.t15 VSS 0.544019f
C6540 a_65486_n35156.t1 VSS 0.347769f
C6541 a_33249_34067.n0 VSS 0.97453f
C6542 a_33249_34067.n1 VSS 0.846499f
C6543 a_33249_34067.n2 VSS 0.928454f
C6544 a_33249_34067.n3 VSS 0.634254f
C6545 a_33249_34067.n4 VSS 0.942033f
C6546 a_33249_34067.n5 VSS 0.942032f
C6547 a_33249_34067.n6 VSS 0.500233f
C6548 a_33249_34067.n7 VSS 0.846499f
C6549 a_33249_34067.n8 VSS 0.928454f
C6550 a_33249_34067.n9 VSS 1.10607f
C6551 a_33249_34067.n10 VSS 0.97453f
C6552 a_33249_34067.n11 VSS 0.846499f
C6553 a_33249_34067.n12 VSS 0.928454f
C6554 a_33249_34067.n13 VSS 0.634254f
C6555 a_33249_34067.n14 VSS 0.942033f
C6556 a_33249_34067.n15 VSS 0.942032f
C6557 a_33249_34067.n16 VSS 0.500233f
C6558 a_33249_34067.n17 VSS 0.846499f
C6559 a_33249_34067.n18 VSS 0.928454f
C6560 a_33249_34067.n19 VSS 1.10607f
C6561 a_33249_34067.n20 VSS 0.559204f
C6562 a_33249_34067.n21 VSS 0.892947f
C6563 a_33249_34067.n22 VSS 1.4803f
C6564 a_33249_34067.n23 VSS 0.957103f
C6565 a_33249_34067.n24 VSS 0.829503f
C6566 a_33249_34067.n25 VSS 1.47288f
C6567 a_33249_34067.t55 VSS 0.07705f
C6568 a_33249_34067.t38 VSS 0.189907f
C6569 a_33249_34067.t43 VSS 0.231711f
C6570 a_33249_34067.n26 VSS 1.24188f
C6571 a_33249_34067.t47 VSS 0.189907f
C6572 a_33249_34067.t52 VSS 0.231711f
C6573 a_33249_34067.n27 VSS 0.679056f
C6574 a_33249_34067.n28 VSS 1.38796f
C6575 a_33249_34067.t23 VSS 0.431389f
C6576 a_33249_34067.t88 VSS 0.07705f
C6577 a_33249_34067.t63 VSS 0.07705f
C6578 a_33249_34067.n29 VSS 0.333558f
C6579 a_33249_34067.n30 VSS 1.09797f
C6580 a_33249_34067.t36 VSS 0.326996f
C6581 a_33249_34067.n31 VSS 0.929305f
C6582 a_33249_34067.t69 VSS 0.324197f
C6583 a_33249_34067.n32 VSS 0.842019f
C6584 a_33249_34067.n33 VSS 0.750688f
C6585 a_33249_34067.n34 VSS 2.82575f
C6586 a_33249_34067.t101 VSS 0.435448f
C6587 a_33249_34067.t81 VSS 0.07705f
C6588 a_33249_34067.t53 VSS 0.07705f
C6589 a_33249_34067.n35 VSS 0.33288f
C6590 a_33249_34067.t26 VSS 0.326332f
C6591 a_33249_34067.t57 VSS 0.325909f
C6592 a_33249_34067.t22 VSS 0.07705f
C6593 a_33249_34067.t87 VSS 0.07705f
C6594 a_33249_34067.n36 VSS 0.33288f
C6595 a_33249_34067.t61 VSS 0.326332f
C6596 a_33249_34067.t50 VSS 0.326332f
C6597 a_33249_34067.t25 VSS 0.07705f
C6598 a_33249_34067.t82 VSS 0.07705f
C6599 a_33249_34067.n37 VSS 0.33288f
C6600 a_33249_34067.t54 VSS 0.326332f
C6601 a_33249_34067.t84 VSS 0.325909f
C6602 a_33249_34067.t28 VSS 0.07705f
C6603 a_33249_34067.t83 VSS 0.07705f
C6604 a_33249_34067.n38 VSS 0.33288f
C6605 a_33249_34067.t70 VSS 0.436032f
C6606 a_33249_34067.t30 VSS 0.07705f
C6607 a_33249_34067.t99 VSS 0.07705f
C6608 a_33249_34067.n39 VSS 0.333558f
C6609 a_33249_34067.n40 VSS 0.500562f
C6610 a_33249_34067.t72 VSS 0.326905f
C6611 a_33249_34067.n41 VSS 0.942835f
C6612 a_33249_34067.t62 VSS 0.324197f
C6613 a_33249_34067.n42 VSS 0.93517f
C6614 a_33249_34067.t32 VSS 0.07705f
C6615 a_33249_34067.t90 VSS 0.07705f
C6616 a_33249_34067.n43 VSS 0.333558f
C6617 a_33249_34067.n44 VSS 0.634013f
C6618 a_33249_34067.t65 VSS 0.326996f
C6619 a_33249_34067.n45 VSS 0.929305f
C6620 a_33249_34067.t97 VSS 0.324197f
C6621 a_33249_34067.n46 VSS 0.842019f
C6622 a_33249_34067.t77 VSS 0.437465f
C6623 a_33249_34067.t37 VSS 0.07705f
C6624 a_33249_34067.t96 VSS 0.07705f
C6625 a_33249_34067.n47 VSS 0.333558f
C6626 a_33249_34067.n48 VSS 0.979186f
C6627 a_33249_34067.n49 VSS 0.750687f
C6628 a_33249_34067.t19 VSS 0.07705f
C6629 a_33249_34067.t71 VSS 0.07705f
C6630 a_33249_34067.n50 VSS 0.180326f
C6631 a_33249_34067.t24 VSS 0.07705f
C6632 a_33249_34067.t76 VSS 0.07705f
C6633 a_33249_34067.n51 VSS 0.229413f
C6634 a_33249_34067.n52 VSS 0.522158f
C6635 a_33249_34067.n53 VSS 0.907551f
C6636 a_33249_34067.n54 VSS 4.90658f
C6637 a_33249_34067.n55 VSS 7.56734f
C6638 a_33249_34067.t34 VSS 0.189907f
C6639 a_33249_34067.t35 VSS 0.231711f
C6640 a_33249_34067.n56 VSS 1.24177f
C6641 a_33249_34067.t93 VSS 0.07705f
C6642 a_33249_34067.t44 VSS 0.07705f
C6643 a_33249_34067.n57 VSS 0.180326f
C6644 a_33249_34067.t94 VSS 0.07705f
C6645 a_33249_34067.t46 VSS 0.07705f
C6646 a_33249_34067.n58 VSS 0.229413f
C6647 a_33249_34067.n59 VSS 0.522158f
C6648 a_33249_34067.n60 VSS 1.14141f
C6649 a_33249_34067.n61 VSS 5.40296f
C6650 a_33249_34067.t106 VSS 0.073381f
C6651 a_33249_34067.t120 VSS 0.073381f
C6652 a_33249_34067.n62 VSS 0.375103f
C6653 a_33249_34067.n63 VSS 1.62793f
C6654 a_33249_34067.t129 VSS 0.189776f
C6655 a_33249_34067.t125 VSS 0.22852f
C6656 a_33249_34067.n64 VSS 1.13624f
C6657 a_33249_34067.t128 VSS 0.073381f
C6658 a_33249_34067.t140 VSS 0.073381f
C6659 a_33249_34067.n65 VSS 0.169422f
C6660 a_33249_34067.t121 VSS 0.073381f
C6661 a_33249_34067.t134 VSS 0.073381f
C6662 a_33249_34067.n66 VSS 0.213704f
C6663 a_33249_34067.n67 VSS 0.536186f
C6664 a_33249_34067.n68 VSS 1.05092f
C6665 a_33249_34067.t133 VSS 0.43417f
C6666 a_33249_34067.t110 VSS 0.073381f
C6667 a_33249_34067.t108 VSS 0.073381f
C6668 a_33249_34067.n69 VSS 0.310987f
C6669 a_33249_34067.t114 VSS 0.319326f
C6670 a_33249_34067.n70 VSS 0.954758f
C6671 a_33249_34067.t123 VSS 0.073381f
C6672 a_33249_34067.t135 VSS 0.073381f
C6673 a_33249_34067.n71 VSS 0.310987f
C6674 a_33249_34067.t118 VSS 0.073381f
C6675 a_33249_34067.t122 VSS 0.073381f
C6676 a_33249_34067.n72 VSS 0.310987f
C6677 a_33249_34067.t130 VSS 0.319326f
C6678 a_33249_34067.n73 VSS 0.954758f
C6679 a_33249_34067.t109 VSS 0.319326f
C6680 a_33249_34067.n74 VSS 1.03839f
C6681 a_33249_34067.n75 VSS 1.04549f
C6682 a_33249_34067.n76 VSS 4.76973f
C6683 a_33249_34067.n77 VSS 1.24553f
C6684 a_33249_34067.t141 VSS 0.189776f
C6685 a_33249_34067.t136 VSS 0.22852f
C6686 a_33249_34067.n78 VSS 0.655117f
C6687 a_33249_34067.n79 VSS 1.16921f
C6688 a_33249_34067.t139 VSS 0.073381f
C6689 a_33249_34067.t117 VSS 0.073381f
C6690 a_33249_34067.n80 VSS 0.169422f
C6691 a_33249_34067.t132 VSS 0.073381f
C6692 a_33249_34067.t115 VSS 0.073381f
C6693 a_33249_34067.n81 VSS 0.213704f
C6694 a_33249_34067.n82 VSS 0.536186f
C6695 a_33249_34067.n83 VSS 0.85096f
C6696 a_33249_34067.n84 VSS 5.1877f
C6697 a_33249_34067.t137 VSS 0.073381f
C6698 a_33249_34067.t113 VSS 0.073381f
C6699 a_33249_34067.n85 VSS 0.478627f
C6700 a_33249_34067.t111 VSS 0.318572f
C6701 a_33249_34067.n86 VSS 1.51427f
C6702 a_33249_34067.t116 VSS 0.315853f
C6703 a_33249_34067.n87 VSS 0.836289f
C6704 a_33249_34067.n88 VSS 0.21186f
C6705 a_33249_34067.t127 VSS 0.073381f
C6706 a_33249_34067.t138 VSS 0.073381f
C6707 a_33249_34067.n89 VSS 0.31157f
C6708 a_33249_34067.n90 VSS 0.93242f
C6709 a_33249_34067.t112 VSS 0.073381f
C6710 a_33249_34067.t119 VSS 0.073381f
C6711 a_33249_34067.n91 VSS 0.31157f
C6712 a_33249_34067.n92 VSS 1.06142f
C6713 a_33249_34067.t126 VSS 0.318572f
C6714 a_33249_34067.n93 VSS 0.925218f
C6715 a_33249_34067.t131 VSS 0.315853f
C6716 a_33249_34067.n94 VSS 0.836289f
C6717 a_33249_34067.t107 VSS 0.073381f
C6718 a_33249_34067.t124 VSS 0.073381f
C6719 a_33249_34067.n95 VSS 0.375696f
C6720 a_33249_34067.n96 VSS 0.794745f
C6721 a_33249_34067.n97 VSS 4.38744f
C6722 a_33249_34067.n98 VSS 5.63217f
C6723 a_33249_34067.t17 VSS 0.073381f
C6724 a_33249_34067.t4 VSS 0.073381f
C6725 a_33249_34067.n99 VSS 0.428777f
C6726 a_33249_34067.t10 VSS 0.276508f
C6727 a_33249_34067.t6 VSS 0.073381f
C6728 a_33249_34067.t5 VSS 0.073381f
C6729 a_33249_34067.n100 VSS 0.263142f
C6730 a_33249_34067.t11 VSS 0.276508f
C6731 a_33249_34067.n101 VSS 3.23788f
C6732 a_33249_34067.t8 VSS 0.073381f
C6733 a_33249_34067.t13 VSS 0.073381f
C6734 a_33249_34067.n102 VSS 0.198194f
C6735 a_33249_34067.t16 VSS 0.073381f
C6736 a_33249_34067.t2 VSS 0.073381f
C6737 a_33249_34067.n103 VSS 0.181808f
C6738 a_33249_34067.n104 VSS 1.12528f
C6739 a_33249_34067.t3 VSS 0.215053f
C6740 a_33249_34067.t9 VSS 0.200752f
C6741 a_33249_34067.n105 VSS 0.667789f
C6742 a_33249_34067.n106 VSS 1.45399f
C6743 a_33249_34067.n107 VSS 3.01461f
C6744 a_33249_34067.t7 VSS 0.383044f
C6745 a_33249_34067.t12 VSS 0.073381f
C6746 a_33249_34067.t0 VSS 0.073381f
C6747 a_33249_34067.n108 VSS 0.263908f
C6748 a_33249_34067.n109 VSS 1.44297f
C6749 a_33249_34067.t15 VSS 0.073381f
C6750 a_33249_34067.t14 VSS 0.073381f
C6751 a_33249_34067.n110 VSS 0.263908f
C6752 a_33249_34067.n111 VSS 0.996653f
C6753 a_33249_34067.t1 VSS 0.277157f
C6754 a_33249_34067.n112 VSS 0.556872f
C6755 a_33249_34067.n113 VSS 8.876969f
C6756 a_33249_34067.n114 VSS 12.1615f
C6757 a_33249_34067.t89 VSS 0.435448f
C6758 a_33249_34067.t73 VSS 0.07705f
C6759 a_33249_34067.t42 VSS 0.07705f
C6760 a_33249_34067.n115 VSS 0.33288f
C6761 a_33249_34067.t18 VSS 0.326332f
C6762 a_33249_34067.t48 VSS 0.325909f
C6763 a_33249_34067.t100 VSS 0.07705f
C6764 a_33249_34067.t80 VSS 0.07705f
C6765 a_33249_34067.n116 VSS 0.33288f
C6766 a_33249_34067.t51 VSS 0.326332f
C6767 a_33249_34067.t39 VSS 0.326332f
C6768 a_33249_34067.t104 VSS 0.07705f
C6769 a_33249_34067.t75 VSS 0.07705f
C6770 a_33249_34067.n117 VSS 0.33288f
C6771 a_33249_34067.t45 VSS 0.326332f
C6772 a_33249_34067.t79 VSS 0.325909f
C6773 a_33249_34067.t21 VSS 0.07705f
C6774 a_33249_34067.t78 VSS 0.07705f
C6775 a_33249_34067.n118 VSS 0.33288f
C6776 a_33249_34067.t60 VSS 0.436032f
C6777 a_33249_34067.n119 VSS 0.214777f
C6778 a_33249_34067.n120 VSS 0.214777f
C6779 a_33249_34067.n121 VSS 3.96945f
C6780 a_33249_34067.n122 VSS 3.16582f
C6781 a_33249_34067.n123 VSS 1.46267f
C6782 a_33249_34067.t40 VSS 0.189907f
C6783 a_33249_34067.t41 VSS 0.231711f
C6784 a_33249_34067.n124 VSS 0.679056f
C6785 a_33249_34067.n125 VSS 1.38796f
C6786 a_33249_34067.t102 VSS 0.07705f
C6787 a_33249_34067.t66 VSS 0.07705f
C6788 a_33249_34067.n126 VSS 0.180326f
C6789 a_33249_34067.t103 VSS 0.07705f
C6790 a_33249_34067.t67 VSS 0.07705f
C6791 a_33249_34067.n127 VSS 0.229413f
C6792 a_33249_34067.n128 VSS 0.522158f
C6793 a_33249_34067.n129 VSS 0.907551f
C6794 a_33249_34067.n130 VSS 3.64644f
C6795 a_33249_34067.t20 VSS 0.431389f
C6796 a_33249_34067.t85 VSS 0.07705f
C6797 a_33249_34067.t58 VSS 0.07705f
C6798 a_33249_34067.n131 VSS 0.333558f
C6799 a_33249_34067.n132 VSS 1.09797f
C6800 a_33249_34067.t31 VSS 0.326996f
C6801 a_33249_34067.n133 VSS 0.929305f
C6802 a_33249_34067.t64 VSS 0.324197f
C6803 a_33249_34067.n134 VSS 0.842019f
C6804 a_33249_34067.n135 VSS 0.214786f
C6805 a_33249_34067.t27 VSS 0.07705f
C6806 a_33249_34067.t95 VSS 0.07705f
C6807 a_33249_34067.n136 VSS 0.333558f
C6808 a_33249_34067.n137 VSS 0.500562f
C6809 a_33249_34067.t68 VSS 0.326905f
C6810 a_33249_34067.n138 VSS 0.942835f
C6811 a_33249_34067.t56 VSS 0.324197f
C6812 a_33249_34067.n139 VSS 0.93517f
C6813 a_33249_34067.t29 VSS 0.07705f
C6814 a_33249_34067.t86 VSS 0.07705f
C6815 a_33249_34067.n140 VSS 0.333558f
C6816 a_33249_34067.n141 VSS 0.634013f
C6817 a_33249_34067.t59 VSS 0.326996f
C6818 a_33249_34067.n142 VSS 0.929305f
C6819 a_33249_34067.t92 VSS 0.324197f
C6820 a_33249_34067.n143 VSS 0.842019f
C6821 a_33249_34067.t74 VSS 0.437465f
C6822 a_33249_34067.t33 VSS 0.07705f
C6823 a_33249_34067.t91 VSS 0.07705f
C6824 a_33249_34067.n144 VSS 0.333558f
C6825 a_33249_34067.n145 VSS 0.979186f
C6826 a_33249_34067.n146 VSS 0.214786f
C6827 a_33249_34067.n147 VSS 2.82575f
C6828 a_33249_34067.n148 VSS 3.14342f
C6829 a_33249_34067.n149 VSS 0.214777f
C6830 a_33249_34067.n150 VSS 0.214777f
C6831 a_33249_34067.n151 VSS 3.14342f
C6832 a_33249_34067.n152 VSS 4.42596f
C6833 a_33249_34067.n153 VSS 1.46262f
C6834 a_33249_34067.n154 VSS 1.14136f
C6835 a_33249_34067.t98 VSS 0.07705f
C6836 a_33249_34067.t49 VSS 0.07705f
C6837 a_33249_34067.n155 VSS 0.180326f
C6838 a_33249_34067.n156 VSS 0.522158f
C6839 a_33249_34067.n157 VSS 0.229413f
C6840 a_33249_34067.t105 VSS 0.07705f
C6841 a_33379_34007.n0 VSS 1.38521f
C6842 a_33379_34007.t1 VSS 0.192333f
C6843 a_33379_34007.n1 VSS 0.669724f
C6844 a_33379_34007.t0 VSS 0.199152f
C6845 a_33379_34007.n2 VSS 0.002305f
C6846 a_33379_34007.n3 VSS 0.008055f
C6847 a_33379_34007.n4 VSS 0.002305f
C6848 a_33379_34007.n5 VSS 0.002109f
C6849 a_33379_34007.n6 VSS 0.008055f
C6850 a_33379_34007.n7 VSS 0.002305f
C6851 a_33379_34007.n8 VSS 0.002109f
C6852 a_33379_34007.n9 VSS 0.008055f
C6853 a_33379_34007.t87 VSS 0.019031f
C6854 a_33379_34007.n10 VSS 0.013755f
C6855 a_33379_34007.n11 VSS 0.002305f
C6856 a_33379_34007.n12 VSS 0.009971f
C6857 a_33379_34007.n13 VSS 0.002305f
C6858 a_33379_34007.n14 VSS 0.002109f
C6859 a_33379_34007.n15 VSS 0.008055f
C6860 a_33379_34007.n16 VSS 0.002305f
C6861 a_33379_34007.n17 VSS 0.002109f
C6862 a_33379_34007.n18 VSS 0.008055f
C6863 a_33379_34007.n19 VSS 0.008055f
C6864 a_33379_34007.n20 VSS 0.009971f
C6865 a_33379_34007.n21 VSS 0.013755f
C6866 a_33379_34007.n22 VSS 0.00225f
C6867 a_33379_34007.n23 VSS 0.008045f
C6868 a_33379_34007.n24 VSS 0.00225f
C6869 a_33379_34007.n25 VSS 0.00894f
C6870 a_33379_34007.n26 VSS 0.015839f
C6871 a_33379_34007.n27 VSS 0.001317f
C6872 a_33379_34007.n28 VSS 0.00225f
C6873 a_33379_34007.n29 VSS 0.008045f
C6874 a_33379_34007.n30 VSS 0.001317f
C6875 a_33379_34007.n31 VSS 0.00225f
C6876 a_33379_34007.n32 VSS 0.008045f
C6877 a_33379_34007.n33 VSS 0.00894f
C6878 a_33379_34007.n34 VSS 0.015839f
C6879 a_33379_34007.n35 VSS 0.001317f
C6880 a_33379_34007.n36 VSS 0.008045f
C6881 a_33379_34007.n37 VSS 0.008035f
C6882 a_33379_34007.n38 VSS 0.009116f
C6883 a_33379_34007.n39 VSS 0.015844f
C6884 a_33379_34007.n40 VSS 0.001317f
C6885 a_33379_34007.n41 VSS 0.001912f
C6886 a_33379_34007.n42 VSS 0.008035f
C6887 a_33379_34007.n43 VSS 0.001317f
C6888 a_33379_34007.n44 VSS 0.001912f
C6889 a_33379_34007.n45 VSS 0.008035f
C6890 a_33379_34007.n46 VSS 0.001912f
C6891 a_33379_34007.n47 VSS 0.009116f
C6892 a_33379_34007.n48 VSS 0.015844f
C6893 a_33379_34007.n49 VSS 0.001912f
C6894 a_33379_34007.n50 VSS 0.008035f
C6895 a_33379_34007.n51 VSS 0.007934f
C6896 a_33379_34007.n52 VSS 0.001317f
C6897 a_33379_34007.n53 VSS 0.007934f
C6898 a_33379_34007.n54 VSS 0.009766f
C6899 a_33379_34007.n55 VSS 0.01388f
C6900 a_33379_34007.n56 VSS 0.007934f
C6901 a_33379_34007.n57 VSS 0.001317f
C6902 a_33379_34007.n58 VSS 0.007934f
C6903 a_33379_34007.n59 VSS 0.001317f
C6904 a_33379_34007.n60 VSS 0.007934f
C6905 a_33379_34007.n61 VSS 0.001317f
C6906 a_33379_34007.n62 VSS 0.00222f
C6907 a_33379_34007.n63 VSS 0.007934f
C6908 a_33379_34007.n64 VSS 0.00224f
C6909 a_33379_34007.n65 VSS 0.00222f
C6910 a_33379_34007.n66 VSS 0.007934f
C6911 a_33379_34007.n67 VSS 0.007934f
C6912 a_33379_34007.n68 VSS 0.008912f
C6913 a_33379_34007.n69 VSS 0.015582f
C6914 a_33379_34007.n70 VSS 0.001317f
C6915 a_33379_34007.n71 VSS 0.00224f
C6916 a_33379_34007.n72 VSS 0.007934f
C6917 a_33379_34007.n73 VSS 0.001317f
C6918 a_33379_34007.n74 VSS 0.00224f
C6919 a_33379_34007.n75 VSS 0.007934f
C6920 a_33379_34007.n76 VSS 0.001317f
C6921 a_33379_34007.n77 VSS 0.00222f
C6922 a_33379_34007.n78 VSS 0.007934f
C6923 a_33379_34007.n79 VSS 0.00224f
C6924 a_33379_34007.n80 VSS 0.00222f
C6925 a_33379_34007.n81 VSS 0.007934f
C6926 a_33379_34007.n82 VSS 0.009766f
C6927 a_33379_34007.n83 VSS 0.01388f
C6928 a_33379_34007.n84 VSS 0.00224f
C6929 a_33379_34007.n85 VSS 0.00222f
C6930 a_33379_34007.n86 VSS 0.007934f
C6931 a_33379_34007.n87 VSS 0.001317f
C6932 a_33379_34007.n88 VSS 0.00224f
C6933 a_33379_34007.n89 VSS 0.007934f
C6934 a_33379_34007.n90 VSS 0.001317f
C6935 a_33379_34007.n91 VSS 0.00224f
C6936 a_33379_34007.n92 VSS 0.007934f
C6937 a_33379_34007.n93 VSS 0.006222f
C6938 a_33379_34007.n94 VSS 0.007934f
C6939 a_33379_34007.n95 VSS 0.00224f
C6940 a_33379_34007.n96 VSS 0.007934f
C6941 a_33379_34007.n97 VSS 0.00224f
C6942 a_33379_34007.n98 VSS 0.00222f
C6943 a_33379_34007.n99 VSS 0.007934f
C6944 a_33379_34007.n100 VSS 0.00224f
C6945 a_33379_34007.n101 VSS 0.008912f
C6946 a_33379_34007.n102 VSS 0.015582f
C6947 a_33379_34007.n103 VSS 0.00224f
C6948 a_33379_34007.n104 VSS 0.007934f
C6949 a_33379_34007.n105 VSS 0.00224f
C6950 a_33379_34007.n106 VSS 0.007934f
C6951 a_33379_34007.t27 VSS 0.215533p
C6952 a_33379_34007.t3 VSS 0.022362f
C6953 a_33379_34007.n107 VSS 0.094108f
C6954 a_33379_34007.n108 VSS 0.198968f
C6955 a_33379_34007.n109 VSS 0.010991f
C6956 a_33379_34007.n110 VSS 0.001317f
C6957 a_33379_34007.n111 VSS 0.002368f
C6958 a_33379_34007.n112 VSS 0.001912f
C6959 a_33379_34007.n113 VSS 0.002427f
C6960 a_33379_34007.n114 VSS 0.002368f
C6961 a_33379_34007.t46 VSS 0.018613f
C6962 a_33379_34007.n115 VSS 0.010991f
C6963 a_33379_34007.n116 VSS 0.001317f
C6964 a_33379_34007.t21 VSS 0.018613f
C6965 a_33379_34007.n117 VSS 0.008803f
C6966 a_33379_34007.n118 VSS 0.002427f
C6967 a_33379_34007.n119 VSS 0.002098f
C6968 a_33379_34007.t47 VSS 0.018613f
C6969 a_33379_34007.n120 VSS 0.007288f
C6970 a_33379_34007.n121 VSS 8.32e-19
C6971 a_33379_34007.n122 VSS 0.001912f
C6972 a_33379_34007.n123 VSS 0.002012f
C6973 a_33379_34007.n124 VSS 0.002012f
C6974 a_33379_34007.t74 VSS 0.018613f
C6975 a_33379_34007.n125 VSS 0.006231f
C6976 a_33379_34007.t72 VSS 0.018613f
C6977 a_33379_34007.n126 VSS 0.015182f
C6978 a_33379_34007.t11 VSS 0.018613f
C6979 a_33379_34007.n127 VSS 0.012393f
C6980 a_33379_34007.t61 VSS 0.018613f
C6981 a_33379_34007.n128 VSS 0.015194f
C6982 a_33379_34007.n129 VSS 0.002427f
C6983 a_33379_34007.t80 VSS 0.018613f
C6984 a_33379_34007.t10 VSS 0.018613f
C6985 a_33379_34007.n130 VSS 0.007288f
C6986 a_33379_34007.n131 VSS 0.002012f
C6987 a_33379_34007.n132 VSS 0.002427f
C6988 a_33379_34007.t78 VSS 0.018613f
C6989 a_33379_34007.t19 VSS 0.018613f
C6990 a_33379_34007.n133 VSS 0.007288f
C6991 a_33379_34007.n134 VSS 0.002012f
C6992 a_33379_34007.n135 VSS 0.049906f
C6993 a_33379_34007.t45 VSS 0.018613f
C6994 a_33379_34007.t12 VSS 0.018613f
C6995 a_33379_34007.n136 VSS 0.002368f
C6996 a_33379_34007.t73 VSS 0.018613f
C6997 a_33379_34007.n137 VSS 0.002427f
C6998 a_33379_34007.t13 VSS 0.018613f
C6999 a_33379_34007.n138 VSS 0.00935f
C7000 a_33379_34007.t33 VSS 0.018984f
C7001 a_33379_34007.n139 VSS 0.013868f
C7002 a_33379_34007.n140 VSS 0.008496f
C7003 a_33379_34007.n141 VSS 0.002098f
C7004 a_33379_34007.n142 VSS 0.001317f
C7005 a_33379_34007.n143 VSS 0.002368f
C7006 a_33379_34007.n144 VSS 0.002109f
C7007 a_33379_34007.n145 VSS 0.001317f
C7008 a_33379_34007.n146 VSS 0.004205f
C7009 a_33379_34007.n147 VSS 0.006229f
C7010 a_33379_34007.t39 VSS 0.018613f
C7011 a_33379_34007.n148 VSS 0.015194f
C7012 a_33379_34007.t91 VSS 0.018613f
C7013 a_33379_34007.n149 VSS 0.012393f
C7014 a_33379_34007.t63 VSS 0.018613f
C7015 a_33379_34007.n150 VSS 0.015182f
C7016 a_33379_34007.n151 VSS 0.006231f
C7017 a_33379_34007.n152 VSS 0.010991f
C7018 a_33379_34007.n153 VSS 0.001317f
C7019 a_33379_34007.n154 VSS 0.002012f
C7020 a_33379_34007.n155 VSS 0.001912f
C7021 a_33379_34007.n156 VSS 0.001912f
C7022 a_33379_34007.n157 VSS 8.32e-19
C7023 a_33379_34007.n158 VSS 0.001317f
C7024 a_33379_34007.n159 VSS 0.002427f
C7025 a_33379_34007.n160 VSS 0.002098f
C7026 a_33379_34007.n161 VSS 0.001317f
C7027 a_33379_34007.n162 VSS 0.002368f
C7028 a_33379_34007.n163 VSS 0.002801f
C7029 a_33379_34007.t48 VSS 0.018613f
C7030 a_33379_34007.t38 VSS 0.018613f
C7031 a_33379_34007.n164 VSS 0.002445f
C7032 a_33379_34007.n165 VSS 0.001912f
C7033 a_33379_34007.n166 VSS 0.001912f
C7034 a_33379_34007.n167 VSS 8.32e-19
C7035 a_33379_34007.n168 VSS 0.001317f
C7036 a_33379_34007.n169 VSS 0.002427f
C7037 a_33379_34007.n170 VSS 0.002098f
C7038 a_33379_34007.n171 VSS 0.001317f
C7039 a_33379_34007.n172 VSS 0.002368f
C7040 a_33379_34007.n173 VSS 0.002368f
C7041 a_33379_34007.t41 VSS 0.018613f
C7042 a_33379_34007.n174 VSS 0.006229f
C7043 a_33379_34007.n175 VSS 0.004205f
C7044 a_33379_34007.n176 VSS 0.049906f
C7045 a_33379_34007.n177 VSS 0.010885f
C7046 a_33379_34007.n178 VSS 0.00222f
C7047 a_33379_34007.t29 VSS 0.018613f
C7048 a_33379_34007.n179 VSS 0.009703f
C7049 a_33379_34007.t8 VSS 0.019013f
C7050 a_33379_34007.n180 VSS 0.01388f
C7051 a_33379_34007.n181 VSS 0.008554f
C7052 a_33379_34007.n182 VSS 0.002358f
C7053 a_33379_34007.t57 VSS 0.018613f
C7054 a_33379_34007.n183 VSS 0.00222f
C7055 a_33379_34007.n184 VSS 0.002358f
C7056 a_33379_34007.n185 VSS 0.002358f
C7057 a_33379_34007.t84 VSS 0.018613f
C7058 a_33379_34007.n186 VSS 0.006239f
C7059 a_33379_34007.t67 VSS 0.018613f
C7060 a_33379_34007.n187 VSS 0.015072f
C7061 a_33379_34007.t4 VSS 0.018613f
C7062 a_33379_34007.n188 VSS 0.012393f
C7063 a_33379_34007.t55 VSS 0.018613f
C7064 a_33379_34007.n189 VSS 0.015029f
C7065 a_33379_34007.n190 VSS 0.002358f
C7066 a_33379_34007.n191 VSS 0.00279f
C7067 a_33379_34007.t22 VSS 0.018613f
C7068 a_33379_34007.t49 VSS 0.018613f
C7069 a_33379_34007.n192 VSS 0.00279f
C7070 a_33379_34007.n193 VSS 0.002358f
C7071 a_33379_34007.t85 VSS 0.018613f
C7072 a_33379_34007.t28 VSS 0.018613f
C7073 a_33379_34007.n194 VSS 0.002358f
C7074 a_33379_34007.t56 VSS 0.018613f
C7075 a_33379_34007.n195 VSS 0.013615f
C7076 a_33379_34007.n196 VSS 0.002358f
C7077 a_33379_34007.t25 VSS 0.018613f
C7078 a_33379_34007.t82 VSS 0.018613f
C7079 a_33379_34007.n197 VSS 0.008689f
C7080 a_33379_34007.t26 VSS 0.018613f
C7081 a_33379_34007.t40 VSS 0.019019f
C7082 a_33379_34007.n198 VSS 0.00224f
C7083 a_33379_34007.n199 VSS 0.00222f
C7084 a_33379_34007.n200 VSS 0.002358f
C7085 a_33379_34007.n201 VSS 0.00224f
C7086 a_33379_34007.n202 VSS 0.00222f
C7087 a_33379_34007.n203 VSS 0.002358f
C7088 a_33379_34007.n204 VSS 0.001317f
C7089 a_33379_34007.n205 VSS 0.004046f
C7090 a_33379_34007.n206 VSS 0.006222f
C7091 a_33379_34007.t34 VSS 0.018613f
C7092 a_33379_34007.n207 VSS 0.015029f
C7093 a_33379_34007.t86 VSS 0.018613f
C7094 a_33379_34007.n208 VSS 0.012393f
C7095 a_33379_34007.t58 VSS 0.018613f
C7096 a_33379_34007.n209 VSS 0.015072f
C7097 a_33379_34007.n210 VSS 0.006239f
C7098 a_33379_34007.n211 VSS 0.010885f
C7099 a_33379_34007.n212 VSS 0.00224f
C7100 a_33379_34007.n213 VSS 0.00222f
C7101 a_33379_34007.n214 VSS 0.002358f
C7102 a_33379_34007.n215 VSS 0.00224f
C7103 a_33379_34007.n216 VSS 0.00222f
C7104 a_33379_34007.n217 VSS 0.002358f
C7105 a_33379_34007.n218 VSS 0.001317f
C7106 a_33379_34007.n219 VSS 0.002358f
C7107 a_33379_34007.n220 VSS 0.00224f
C7108 a_33379_34007.n221 VSS 0.00222f
C7109 a_33379_34007.t60 VSS 0.018613f
C7110 a_33379_34007.n222 VSS 0.008946f
C7111 a_33379_34007.n223 VSS 0.015587f
C7112 a_33379_34007.n224 VSS 0.00224f
C7113 a_33379_34007.n225 VSS 0.00222f
C7114 a_33379_34007.n226 VSS 0.002358f
C7115 a_33379_34007.n227 VSS 0.001317f
C7116 a_33379_34007.n228 VSS 0.002358f
C7117 a_33379_34007.n229 VSS 0.00224f
C7118 a_33379_34007.t88 VSS 0.018613f
C7119 a_33379_34007.n230 VSS 0.001317f
C7120 a_33379_34007.n231 VSS 0.002358f
C7121 a_33379_34007.n232 VSS 0.002358f
C7122 a_33379_34007.t53 VSS 0.018613f
C7123 a_33379_34007.n233 VSS 0.006222f
C7124 a_33379_34007.n234 VSS 0.004046f
C7125 a_33379_34007.n235 VSS 0.013615f
C7126 a_33379_34007.n236 VSS 0.198968f
C7127 a_33379_34007.n237 VSS 0.132203f
C7128 a_33379_34007.n238 VSS 0.01388f
C7129 a_33379_34007.t79 VSS 0.018613f
C7130 a_33379_34007.n239 VSS 0.002012f
C7131 a_33379_34007.n240 VSS 8.32e-19
C7132 a_33379_34007.n241 VSS 0.008803f
C7133 a_33379_34007.t24 VSS 0.018613f
C7134 a_33379_34007.t90 VSS 0.019031f
C7135 a_33379_34007.n242 VSS 0.002305f
C7136 a_33379_34007.t52 VSS 0.018613f
C7137 a_33379_34007.n243 VSS 0.007288f
C7138 a_33379_34007.n244 VSS 0.002098f
C7139 a_33379_34007.n245 VSS 0.002427f
C7140 a_33379_34007.n246 VSS 0.001317f
C7141 a_33379_34007.n247 VSS 0.002012f
C7142 a_33379_34007.n248 VSS 0.001912f
C7143 a_33379_34007.n249 VSS 0.001317f
C7144 a_33379_34007.n250 VSS 0.010991f
C7145 a_33379_34007.n251 VSS 0.006231f
C7146 a_33379_34007.t76 VSS 0.018613f
C7147 a_33379_34007.n252 VSS 0.015182f
C7148 a_33379_34007.t16 VSS 0.018613f
C7149 a_33379_34007.n253 VSS 0.012393f
C7150 a_33379_34007.t66 VSS 0.018613f
C7151 a_33379_34007.n254 VSS 0.015194f
C7152 a_33379_34007.n255 VSS 0.006229f
C7153 a_33379_34007.n256 VSS 0.004205f
C7154 a_33379_34007.n257 VSS 0.00225f
C7155 a_33379_34007.t83 VSS 0.018613f
C7156 a_33379_34007.n258 VSS 0.002109f
C7157 a_33379_34007.n259 VSS 0.002368f
C7158 a_33379_34007.n260 VSS 0.001317f
C7159 a_33379_34007.n261 VSS 0.002427f
C7160 a_33379_34007.n262 VSS 0.002305f
C7161 a_33379_34007.n263 VSS 0.002098f
C7162 a_33379_34007.t14 VSS 0.018613f
C7163 a_33379_34007.n264 VSS 0.007288f
C7164 a_33379_34007.n265 VSS 8.32e-19
C7165 a_33379_34007.n266 VSS 0.001317f
C7166 a_33379_34007.n267 VSS 0.002012f
C7167 a_33379_34007.n268 VSS 0.002445f
C7168 a_33379_34007.t42 VSS 0.018613f
C7169 a_33379_34007.t54 VSS 0.018613f
C7170 a_33379_34007.n269 VSS 0.002801f
C7171 a_33379_34007.n270 VSS 0.00225f
C7172 a_33379_34007.t81 VSS 0.018613f
C7173 a_33379_34007.n271 VSS 0.001317f
C7174 a_33379_34007.n272 VSS 0.002427f
C7175 a_33379_34007.n273 VSS 0.002427f
C7176 a_33379_34007.n274 VSS 0.002098f
C7177 a_33379_34007.t23 VSS 0.018613f
C7178 a_33379_34007.n275 VSS 0.007288f
C7179 a_33379_34007.n276 VSS 8.32e-19
C7180 a_33379_34007.n277 VSS 0.001912f
C7181 a_33379_34007.n278 VSS 0.002012f
C7182 a_33379_34007.n279 VSS 0.002012f
C7183 a_33379_34007.t51 VSS 0.018613f
C7184 a_33379_34007.n280 VSS 0.006231f
C7185 a_33379_34007.t70 VSS 0.018613f
C7186 a_33379_34007.n281 VSS 0.015182f
C7187 a_33379_34007.t7 VSS 0.018613f
C7188 a_33379_34007.n282 VSS 0.012393f
C7189 a_33379_34007.t44 VSS 0.018613f
C7190 a_33379_34007.n283 VSS 0.015194f
C7191 a_33379_34007.n284 VSS 0.002427f
C7192 a_33379_34007.t77 VSS 0.018613f
C7193 a_33379_34007.t18 VSS 0.018613f
C7194 a_33379_34007.n285 VSS 0.00935f
C7195 a_33379_34007.t36 VSS 0.018984f
C7196 a_33379_34007.n286 VSS 0.013868f
C7197 a_33379_34007.n287 VSS 0.008496f
C7198 a_33379_34007.n288 VSS 0.002098f
C7199 a_33379_34007.n289 VSS 0.001317f
C7200 a_33379_34007.n290 VSS 0.002368f
C7201 a_33379_34007.n291 VSS 0.002368f
C7202 a_33379_34007.t17 VSS 0.018613f
C7203 a_33379_34007.n292 VSS 0.006229f
C7204 a_33379_34007.n293 VSS 0.004205f
C7205 a_33379_34007.n294 VSS 0.01388f
C7206 a_33379_34007.n295 VSS 0.132203f
C7207 a_33379_34007.n296 VSS 0.010885f
C7208 a_33379_34007.n297 VSS 0.002358f
C7209 a_33379_34007.t71 VSS 0.018613f
C7210 a_33379_34007.n298 VSS 0.008946f
C7211 a_33379_34007.n299 VSS 0.002358f
C7212 a_33379_34007.t9 VSS 0.018613f
C7213 a_33379_34007.n300 VSS 0.002358f
C7214 a_33379_34007.t62 VSS 0.018613f
C7215 a_33379_34007.n301 VSS 0.004046f
C7216 a_33379_34007.t92 VSS 0.018613f
C7217 a_33379_34007.n302 VSS 0.002358f
C7218 a_33379_34007.t68 VSS 0.018613f
C7219 a_33379_34007.n303 VSS 0.002358f
C7220 a_33379_34007.t37 VSS 0.018613f
C7221 a_33379_34007.n304 VSS 0.009703f
C7222 a_33379_34007.t20 VSS 0.019013f
C7223 a_33379_34007.n305 VSS 0.01388f
C7224 a_33379_34007.n306 VSS 0.008554f
C7225 a_33379_34007.n307 VSS 0.00222f
C7226 a_33379_34007.n308 VSS 0.001317f
C7227 a_33379_34007.n309 VSS 0.002358f
C7228 a_33379_34007.n310 VSS 0.00222f
C7229 a_33379_34007.n311 VSS 0.001317f
C7230 a_33379_34007.n312 VSS 0.013615f
C7231 a_33379_34007.n313 VSS 0.010885f
C7232 a_33379_34007.n314 VSS 0.006239f
C7233 a_33379_34007.t75 VSS 0.018613f
C7234 a_33379_34007.n315 VSS 0.015072f
C7235 a_33379_34007.t15 VSS 0.018613f
C7236 a_33379_34007.n316 VSS 0.012393f
C7237 a_33379_34007.t64 VSS 0.018613f
C7238 a_33379_34007.n317 VSS 0.015029f
C7239 a_33379_34007.n318 VSS 0.001317f
C7240 a_33379_34007.n319 VSS 0.002358f
C7241 a_33379_34007.n320 VSS 0.00222f
C7242 a_33379_34007.n321 VSS 0.001317f
C7243 a_33379_34007.n322 VSS 0.002358f
C7244 a_33379_34007.n323 VSS 0.00222f
C7245 a_33379_34007.t30 VSS 0.018613f
C7246 a_33379_34007.n324 VSS 0.001317f
C7247 a_33379_34007.n325 VSS 0.002358f
C7248 a_33379_34007.n326 VSS 0.00279f
C7249 a_33379_34007.t59 VSS 0.018613f
C7250 a_33379_34007.n327 VSS 0.015587f
C7251 a_33379_34007.n328 VSS 0.00279f
C7252 a_33379_34007.n329 VSS 0.00222f
C7253 a_33379_34007.t5 VSS 0.018613f
C7254 a_33379_34007.n330 VSS 0.001317f
C7255 a_33379_34007.n331 VSS 0.002358f
C7256 a_33379_34007.n332 VSS 0.002358f
C7257 a_33379_34007.t35 VSS 0.018613f
C7258 a_33379_34007.n333 VSS 0.00222f
C7259 a_33379_34007.n334 VSS 0.002358f
C7260 a_33379_34007.n335 VSS 0.002358f
C7261 a_33379_34007.t65 VSS 0.018613f
C7262 a_33379_34007.n336 VSS 0.006239f
C7263 a_33379_34007.t69 VSS 0.018613f
C7264 a_33379_34007.n337 VSS 0.015072f
C7265 a_33379_34007.t6 VSS 0.018613f
C7266 a_33379_34007.n338 VSS 0.012393f
C7267 a_33379_34007.t43 VSS 0.018613f
C7268 a_33379_34007.n339 VSS 0.015029f
C7269 a_33379_34007.n340 VSS 0.002358f
C7270 a_33379_34007.t50 VSS 0.019019f
C7271 a_33379_34007.t32 VSS 0.018613f
C7272 a_33379_34007.n341 VSS 0.008689f
C7273 a_33379_34007.n342 VSS 0.00224f
C7274 a_33379_34007.t89 VSS 0.018613f
C7275 a_33379_34007.n343 VSS 0.001317f
C7276 a_33379_34007.n344 VSS 0.002358f
C7277 a_33379_34007.n345 VSS 0.002358f
C7278 a_33379_34007.t31 VSS 0.018613f
C7279 a_33379_34007.n346 VSS 0.006222f
C7280 a_33379_34007.n347 VSS 0.004046f
C7281 a_33379_34007.n348 VSS 0.013615f
C7282 a_33379_34007.n349 VSS 0.236716f
C7283 a_33379_34007.n350 VSS 0.962583f
C7284 a_33379_34007.n351 VSS 1.46779f
C7285 a_33379_34007.t2 VSS 0.019073f
C7286 a_60677_10448.t1 VSS 0.935952f
C7287 a_60677_10448.t2 VSS 56.413002f
C7288 a_60677_10448.t5 VSS 0.475426f
C7289 a_60677_10448.t3 VSS 0.789344f
C7290 a_60677_10448.t4 VSS 31.633099f
C7291 a_60677_10448.t0 VSS 0.553147f
C7292 a_71281_n10073.n0 VSS 3.63047f
C7293 a_71281_n10073.t63 VSS 0.033171f
C7294 a_71281_n10073.t45 VSS 0.157501f
C7295 a_71281_n10073.n1 VSS 0.051957f
C7296 a_71281_n10073.n2 VSS 0.046844f
C7297 a_71281_n10073.n3 VSS 0.431228f
C7298 a_71281_n10073.t174 VSS 0.41704f
C7299 a_71281_n10073.n4 VSS 0.425799f
C7300 a_71281_n10073.t228 VSS 0.377955f
C7301 a_71281_n10073.n5 VSS 0.425799f
C7302 a_71281_n10073.n6 VSS 0.046844f
C7303 a_71281_n10073.t108 VSS 0.417015f
C7304 a_71281_n10073.t322 VSS 0.377866f
C7305 a_71281_n10073.n7 VSS 0.431228f
C7306 a_71281_n10073.n8 VSS 0.041724f
C7307 a_71281_n10073.n9 VSS 0.147642f
C7308 a_71281_n10073.t261 VSS 0.332539f
C7309 a_71281_n10073.n10 VSS 0.147642f
C7310 a_71281_n10073.n11 VSS 0.041724f
C7311 a_71281_n10073.n12 VSS 0.01935f
C7312 a_71281_n10073.n13 VSS 0.536641f
C7313 a_71281_n10073.n14 VSS 0.265045f
C7314 a_71281_n10073.n15 VSS 0.046844f
C7315 a_71281_n10073.n16 VSS 0.431228f
C7316 a_71281_n10073.t254 VSS 0.41704f
C7317 a_71281_n10073.n17 VSS 0.425799f
C7318 a_71281_n10073.t313 VSS 0.377955f
C7319 a_71281_n10073.n18 VSS 0.425799f
C7320 a_71281_n10073.n19 VSS 0.046844f
C7321 a_71281_n10073.n20 VSS 0.01935f
C7322 a_71281_n10073.t173 VSS 0.417015f
C7323 a_71281_n10073.t121 VSS 0.377866f
C7324 a_71281_n10073.n21 VSS 0.431228f
C7325 a_71281_n10073.n22 VSS 0.041724f
C7326 a_71281_n10073.n23 VSS 0.147642f
C7327 a_71281_n10073.t337 VSS 0.332539f
C7328 a_71281_n10073.n24 VSS 0.147642f
C7329 a_71281_n10073.n25 VSS 0.041724f
C7330 a_71281_n10073.n26 VSS 0.01935f
C7331 a_71281_n10073.n27 VSS 0.265045f
C7332 a_71281_n10073.n28 VSS 0.264461f
C7333 a_71281_n10073.n29 VSS 0.046844f
C7334 a_71281_n10073.n30 VSS 0.431228f
C7335 a_71281_n10073.t241 VSS 0.41704f
C7336 a_71281_n10073.n31 VSS 0.425799f
C7337 a_71281_n10073.t299 VSS 0.377955f
C7338 a_71281_n10073.n32 VSS 0.425799f
C7339 a_71281_n10073.n33 VSS 0.046844f
C7340 a_71281_n10073.n34 VSS 0.01935f
C7341 a_71281_n10073.t168 VSS 0.417015f
C7342 a_71281_n10073.t116 VSS 0.377866f
C7343 a_71281_n10073.n35 VSS 0.431228f
C7344 a_71281_n10073.n36 VSS 0.041724f
C7345 a_71281_n10073.n37 VSS 0.147642f
C7346 a_71281_n10073.t332 VSS 0.332539f
C7347 a_71281_n10073.n38 VSS 0.147642f
C7348 a_71281_n10073.n39 VSS 0.041724f
C7349 a_71281_n10073.n40 VSS 0.01935f
C7350 a_71281_n10073.n41 VSS 0.264461f
C7351 a_71281_n10073.n42 VSS 0.264168f
C7352 a_71281_n10073.n43 VSS 0.046844f
C7353 a_71281_n10073.n44 VSS 0.431228f
C7354 a_71281_n10073.t321 VSS 0.41704f
C7355 a_71281_n10073.n45 VSS 0.425799f
C7356 a_71281_n10073.t105 VSS 0.377955f
C7357 a_71281_n10073.n46 VSS 0.425799f
C7358 a_71281_n10073.n47 VSS 0.046844f
C7359 a_71281_n10073.n48 VSS 0.01935f
C7360 a_71281_n10073.t239 VSS 0.417015f
C7361 a_71281_n10073.t180 VSS 0.377866f
C7362 a_71281_n10073.n49 VSS 0.431228f
C7363 a_71281_n10073.n50 VSS 0.041724f
C7364 a_71281_n10073.n51 VSS 0.147642f
C7365 a_71281_n10073.t125 VSS 0.332539f
C7366 a_71281_n10073.n52 VSS 0.147642f
C7367 a_71281_n10073.n53 VSS 0.041724f
C7368 a_71281_n10073.n54 VSS 0.01935f
C7369 a_71281_n10073.n55 VSS 0.21829f
C7370 a_71281_n10073.n56 VSS 0.050894f
C7371 a_71281_n10073.n57 VSS 0.046844f
C7372 a_71281_n10073.n58 VSS 0.431228f
C7373 a_71281_n10073.t126 VSS 0.413932f
C7374 a_71281_n10073.n59 VSS 0.415054f
C7375 a_71281_n10073.t288 VSS 0.377955f
C7376 a_71281_n10073.n60 VSS 0.425799f
C7377 a_71281_n10073.n61 VSS 0.046844f
C7378 a_71281_n10073.t106 VSS 0.417015f
C7379 a_71281_n10073.t190 VSS 0.377866f
C7380 a_71281_n10073.n62 VSS 0.431228f
C7381 a_71281_n10073.n63 VSS 0.041724f
C7382 a_71281_n10073.n64 VSS 0.147642f
C7383 a_71281_n10073.t104 VSS 0.332539f
C7384 a_71281_n10073.n65 VSS 0.147642f
C7385 a_71281_n10073.n66 VSS 0.041724f
C7386 a_71281_n10073.n67 VSS 0.01935f
C7387 a_71281_n10073.n68 VSS 0.527768f
C7388 a_71281_n10073.n69 VSS 0.264168f
C7389 a_71281_n10073.n70 VSS 0.046844f
C7390 a_71281_n10073.n71 VSS 0.431228f
C7391 a_71281_n10073.t333 VSS 0.41704f
C7392 a_71281_n10073.n72 VSS 0.425799f
C7393 a_71281_n10073.t210 VSS 0.377955f
C7394 a_71281_n10073.n73 VSS 0.425799f
C7395 a_71281_n10073.n74 VSS 0.046844f
C7396 a_71281_n10073.t300 VSS 0.417015f
C7397 a_71281_n10073.t128 VSS 0.377866f
C7398 a_71281_n10073.n75 VSS 0.431228f
C7399 a_71281_n10073.n76 VSS 0.01935f
C7400 a_71281_n10073.n77 VSS 0.041724f
C7401 a_71281_n10073.n78 VSS 0.147642f
C7402 a_71281_n10073.t298 VSS 0.332539f
C7403 a_71281_n10073.n79 VSS 0.147642f
C7404 a_71281_n10073.n80 VSS 0.041724f
C7405 a_71281_n10073.n81 VSS 0.01935f
C7406 a_71281_n10073.n82 VSS 0.264168f
C7407 a_71281_n10073.n83 VSS 0.264461f
C7408 a_71281_n10073.n84 VSS 0.046844f
C7409 a_71281_n10073.n85 VSS 0.431228f
C7410 a_71281_n10073.t183 VSS 0.41704f
C7411 a_71281_n10073.n86 VSS 0.425799f
C7412 a_71281_n10073.t84 VSS 0.377955f
C7413 a_71281_n10073.n87 VSS 0.425799f
C7414 a_71281_n10073.n88 VSS 0.046844f
C7415 a_71281_n10073.t161 VSS 0.417015f
C7416 a_71281_n10073.t265 VSS 0.377866f
C7417 a_71281_n10073.n89 VSS 0.431228f
C7418 a_71281_n10073.n90 VSS 0.01935f
C7419 a_71281_n10073.n91 VSS 0.041724f
C7420 a_71281_n10073.n92 VSS 0.147642f
C7421 a_71281_n10073.t155 VSS 0.332539f
C7422 a_71281_n10073.n93 VSS 0.147642f
C7423 a_71281_n10073.n94 VSS 0.041724f
C7424 a_71281_n10073.n95 VSS 0.01935f
C7425 a_71281_n10073.n96 VSS 0.264461f
C7426 a_71281_n10073.n97 VSS 0.265045f
C7427 a_71281_n10073.n98 VSS 0.046844f
C7428 a_71281_n10073.n99 VSS 0.431228f
C7429 a_71281_n10073.t119 VSS 0.41704f
C7430 a_71281_n10073.n100 VSS 0.425799f
C7431 a_71281_n10073.t278 VSS 0.377955f
C7432 a_71281_n10073.n101 VSS 0.425799f
C7433 a_71281_n10073.n102 VSS 0.046844f
C7434 a_71281_n10073.t94 VSS 0.417015f
C7435 a_71281_n10073.t187 VSS 0.377866f
C7436 a_71281_n10073.n103 VSS 0.431228f
C7437 a_71281_n10073.n104 VSS 0.01935f
C7438 a_71281_n10073.n105 VSS 0.041724f
C7439 a_71281_n10073.n106 VSS 0.147642f
C7440 a_71281_n10073.t90 VSS 0.332539f
C7441 a_71281_n10073.n107 VSS 0.147642f
C7442 a_71281_n10073.n108 VSS 0.041724f
C7443 a_71281_n10073.n109 VSS 0.01935f
C7444 a_71281_n10073.n110 VSS 0.218874f
C7445 a_71281_n10073.t15 VSS 0.157278f
C7446 a_71281_n10073.t67 VSS 0.033171f
C7447 a_71281_n10073.t39 VSS 0.033171f
C7448 a_71281_n10073.n111 VSS 0.135406f
C7449 a_71281_n10073.n112 VSS 0.378573f
C7450 a_71281_n10073.n113 VSS 0.091758f
C7451 a_71281_n10073.n114 VSS 0.218874f
C7452 a_71281_n10073.n115 VSS 0.046844f
C7453 a_71281_n10073.n116 VSS 0.431228f
C7454 a_71281_n10073.t124 VSS 0.41704f
C7455 a_71281_n10073.n117 VSS 0.425799f
C7456 a_71281_n10073.t14 VSS 0.377955f
C7457 a_71281_n10073.n118 VSS 0.425799f
C7458 a_71281_n10073.n119 VSS 0.046844f
C7459 a_71281_n10073.t101 VSS 0.417015f
C7460 a_71281_n10073.t38 VSS 0.377866f
C7461 a_71281_n10073.n120 VSS 0.431228f
C7462 a_71281_n10073.n121 VSS 0.01935f
C7463 a_71281_n10073.n122 VSS 0.041724f
C7464 a_71281_n10073.n123 VSS 0.147642f
C7465 a_71281_n10073.t66 VSS 0.332539f
C7466 a_71281_n10073.n124 VSS 0.147642f
C7467 a_71281_n10073.n125 VSS 0.041724f
C7468 a_71281_n10073.n126 VSS 0.01935f
C7469 a_71281_n10073.n127 VSS 0.264461f
C7470 a_71281_n10073.n128 VSS 0.264461f
C7471 a_71281_n10073.n129 VSS 0.046844f
C7472 a_71281_n10073.n130 VSS 0.431228f
C7473 a_71281_n10073.t328 VSS 0.41704f
C7474 a_71281_n10073.n131 VSS 0.425799f
C7475 a_71281_n10073.t30 VSS 0.377955f
C7476 a_71281_n10073.n132 VSS 0.425799f
C7477 a_71281_n10073.n133 VSS 0.046844f
C7478 a_71281_n10073.t293 VSS 0.417015f
C7479 a_71281_n10073.t60 VSS 0.377866f
C7480 a_71281_n10073.n134 VSS 0.431228f
C7481 a_71281_n10073.n135 VSS 0.01935f
C7482 a_71281_n10073.n136 VSS 0.041724f
C7483 a_71281_n10073.n137 VSS 0.147642f
C7484 a_71281_n10073.t8 VSS 0.332539f
C7485 a_71281_n10073.n138 VSS 0.147642f
C7486 a_71281_n10073.n139 VSS 0.041724f
C7487 a_71281_n10073.n140 VSS 0.01935f
C7488 a_71281_n10073.n141 VSS 0.218582f
C7489 a_71281_n10073.t31 VSS 0.033171f
C7490 a_71281_n10073.t9 VSS 0.033171f
C7491 a_71281_n10073.n142 VSS 0.135177f
C7492 a_71281_n10073.t61 VSS 0.157501f
C7493 a_71281_n10073.n143 VSS 0.380031f
C7494 a_71281_n10073.n144 VSS 0.091758f
C7495 a_71281_n10073.n145 VSS 0.21829f
C7496 a_71281_n10073.n146 VSS 0.046844f
C7497 a_71281_n10073.n147 VSS 0.431228f
C7498 a_71281_n10073.t336 VSS 0.41704f
C7499 a_71281_n10073.n148 VSS 0.425799f
C7500 a_71281_n10073.t216 VSS 0.377955f
C7501 a_71281_n10073.n149 VSS 0.425799f
C7502 a_71281_n10073.n150 VSS 0.046844f
C7503 a_71281_n10073.t309 VSS 0.417015f
C7504 a_71281_n10073.t129 VSS 0.377866f
C7505 a_71281_n10073.n151 VSS 0.431228f
C7506 a_71281_n10073.n152 VSS 0.01935f
C7507 a_71281_n10073.n153 VSS 0.041724f
C7508 a_71281_n10073.n154 VSS 0.147642f
C7509 a_71281_n10073.t306 VSS 0.332539f
C7510 a_71281_n10073.n155 VSS 0.147642f
C7511 a_71281_n10073.n156 VSS 0.041724f
C7512 a_71281_n10073.n157 VSS 0.01935f
C7513 a_71281_n10073.n158 VSS 0.264168f
C7514 a_71281_n10073.n159 VSS 0.264461f
C7515 a_71281_n10073.n160 VSS 0.046844f
C7516 a_71281_n10073.n161 VSS 0.431228f
C7517 a_71281_n10073.t329 VSS 0.41704f
C7518 a_71281_n10073.n162 VSS 0.425799f
C7519 a_71281_n10073.t204 VSS 0.377955f
C7520 a_71281_n10073.n163 VSS 0.425799f
C7521 a_71281_n10073.n164 VSS 0.046844f
C7522 a_71281_n10073.t294 VSS 0.417015f
C7523 a_71281_n10073.t127 VSS 0.377866f
C7524 a_71281_n10073.n165 VSS 0.431228f
C7525 a_71281_n10073.n166 VSS 0.01935f
C7526 a_71281_n10073.n167 VSS 0.041724f
C7527 a_71281_n10073.n168 VSS 0.147642f
C7528 a_71281_n10073.t290 VSS 0.332539f
C7529 a_71281_n10073.n169 VSS 0.147642f
C7530 a_71281_n10073.n170 VSS 0.041724f
C7531 a_71281_n10073.n171 VSS 0.01935f
C7532 a_71281_n10073.n172 VSS 0.264461f
C7533 a_71281_n10073.n173 VSS 0.265045f
C7534 a_71281_n10073.n174 VSS 0.046844f
C7535 a_71281_n10073.n175 VSS 0.431228f
C7536 a_71281_n10073.t76 VSS 0.41704f
C7537 a_71281_n10073.n176 VSS 0.425799f
C7538 a_71281_n10073.t238 VSS 0.377955f
C7539 a_71281_n10073.n177 VSS 0.425799f
C7540 a_71281_n10073.n178 VSS 0.046844f
C7541 a_71281_n10073.t330 VSS 0.417015f
C7542 a_71281_n10073.t142 VSS 0.377866f
C7543 a_71281_n10073.n179 VSS 0.431228f
C7544 a_71281_n10073.n180 VSS 0.01935f
C7545 a_71281_n10073.n181 VSS 0.041724f
C7546 a_71281_n10073.n182 VSS 0.147642f
C7547 a_71281_n10073.t324 VSS 0.332539f
C7548 a_71281_n10073.n183 VSS 0.147642f
C7549 a_71281_n10073.n184 VSS 0.041724f
C7550 a_71281_n10073.n185 VSS 0.01935f
C7551 a_71281_n10073.n186 VSS 0.265045f
C7552 a_71281_n10073.n187 VSS 0.264461f
C7553 a_71281_n10073.n188 VSS 0.046844f
C7554 a_71281_n10073.n189 VSS 0.431228f
C7555 a_71281_n10073.t268 VSS 0.41704f
C7556 a_71281_n10073.n190 VSS 0.425799f
C7557 a_71281_n10073.t167 VSS 0.377955f
C7558 a_71281_n10073.n191 VSS 0.425799f
C7559 a_71281_n10073.n192 VSS 0.046844f
C7560 a_71281_n10073.n193 VSS 0.01935f
C7561 a_71281_n10073.t251 VSS 0.417015f
C7562 a_71281_n10073.t79 VSS 0.377866f
C7563 a_71281_n10073.n194 VSS 0.431228f
C7564 a_71281_n10073.n195 VSS 0.041724f
C7565 a_71281_n10073.n196 VSS 0.147642f
C7566 a_71281_n10073.t248 VSS 0.332539f
C7567 a_71281_n10073.n197 VSS 0.147642f
C7568 a_71281_n10073.n198 VSS 0.041724f
C7569 a_71281_n10073.n199 VSS 0.01935f
C7570 a_71281_n10073.n200 VSS 0.59847f
C7571 a_71281_n10073.n201 VSS 0.051957f
C7572 a_71281_n10073.n202 VSS 0.046844f
C7573 a_71281_n10073.n203 VSS 0.431228f
C7574 a_71281_n10073.t178 VSS 0.41704f
C7575 a_71281_n10073.n204 VSS 0.425799f
C7576 a_71281_n10073.t235 VSS 0.377955f
C7577 a_71281_n10073.n205 VSS 0.425799f
C7578 a_71281_n10073.n206 VSS 0.046844f
C7579 a_71281_n10073.t112 VSS 0.417015f
C7580 a_71281_n10073.t120 VSS 0.377866f
C7581 a_71281_n10073.n207 VSS 0.431228f
C7582 a_71281_n10073.n208 VSS 0.041724f
C7583 a_71281_n10073.n209 VSS 0.147642f
C7584 a_71281_n10073.t296 VSS 0.332539f
C7585 a_71281_n10073.n210 VSS 0.147642f
C7586 a_71281_n10073.n211 VSS 0.041724f
C7587 a_71281_n10073.n212 VSS 0.01935f
C7588 a_71281_n10073.n213 VSS 0.536641f
C7589 a_71281_n10073.n214 VSS 0.265045f
C7590 a_71281_n10073.n215 VSS 0.046844f
C7591 a_71281_n10073.n216 VSS 0.431228f
C7592 a_71281_n10073.t259 VSS 0.41704f
C7593 a_71281_n10073.n217 VSS 0.425799f
C7594 a_71281_n10073.t318 VSS 0.377955f
C7595 a_71281_n10073.n218 VSS 0.425799f
C7596 a_71281_n10073.n219 VSS 0.046844f
C7597 a_71281_n10073.n220 VSS 0.01935f
C7598 a_71281_n10073.t177 VSS 0.417015f
C7599 a_71281_n10073.t185 VSS 0.377866f
C7600 a_71281_n10073.n221 VSS 0.431228f
C7601 a_71281_n10073.n222 VSS 0.041724f
C7602 a_71281_n10073.n223 VSS 0.147642f
C7603 a_71281_n10073.t103 VSS 0.332539f
C7604 a_71281_n10073.n224 VSS 0.147642f
C7605 a_71281_n10073.n225 VSS 0.041724f
C7606 a_71281_n10073.n226 VSS 0.01935f
C7607 a_71281_n10073.n227 VSS 0.265045f
C7608 a_71281_n10073.n228 VSS 0.264461f
C7609 a_71281_n10073.n229 VSS 0.046844f
C7610 a_71281_n10073.n230 VSS 0.431228f
C7611 a_71281_n10073.t250 VSS 0.41704f
C7612 a_71281_n10073.n231 VSS 0.425799f
C7613 a_71281_n10073.t305 VSS 0.377955f
C7614 a_71281_n10073.n232 VSS 0.425799f
C7615 a_71281_n10073.n233 VSS 0.046844f
C7616 a_71281_n10073.n234 VSS 0.01935f
C7617 a_71281_n10073.t172 VSS 0.417015f
C7618 a_71281_n10073.t179 VSS 0.377866f
C7619 a_71281_n10073.n235 VSS 0.431228f
C7620 a_71281_n10073.n236 VSS 0.041724f
C7621 a_71281_n10073.n237 VSS 0.147642f
C7622 a_71281_n10073.t96 VSS 0.332539f
C7623 a_71281_n10073.n238 VSS 0.147642f
C7624 a_71281_n10073.n239 VSS 0.041724f
C7625 a_71281_n10073.n240 VSS 0.01935f
C7626 a_71281_n10073.n241 VSS 0.264461f
C7627 a_71281_n10073.n242 VSS 0.264168f
C7628 a_71281_n10073.n243 VSS 0.046844f
C7629 a_71281_n10073.n244 VSS 0.431228f
C7630 a_71281_n10073.t327 VSS 0.41704f
C7631 a_71281_n10073.n245 VSS 0.425799f
C7632 a_71281_n10073.t110 VSS 0.377955f
C7633 a_71281_n10073.n246 VSS 0.425799f
C7634 a_71281_n10073.n247 VSS 0.046844f
C7635 a_71281_n10073.n248 VSS 0.01935f
C7636 a_71281_n10073.t247 VSS 0.417015f
C7637 a_71281_n10073.t260 VSS 0.377866f
C7638 a_71281_n10073.n249 VSS 0.431228f
C7639 a_71281_n10073.n250 VSS 0.041724f
C7640 a_71281_n10073.n251 VSS 0.147642f
C7641 a_71281_n10073.t163 VSS 0.332539f
C7642 a_71281_n10073.n252 VSS 0.147642f
C7643 a_71281_n10073.n253 VSS 0.041724f
C7644 a_71281_n10073.n254 VSS 0.01935f
C7645 a_71281_n10073.n255 VSS 0.21829f
C7646 a_71281_n10073.t69 VSS 0.033171f
C7647 a_71281_n10073.t53 VSS 0.033171f
C7648 a_71281_n10073.n256 VSS 0.135177f
C7649 a_71281_n10073.t19 VSS 0.157501f
C7650 a_71281_n10073.n257 VSS 0.380031f
C7651 a_71281_n10073.n258 VSS 0.091758f
C7652 a_71281_n10073.n259 VSS 0.218582f
C7653 a_71281_n10073.n260 VSS 0.046844f
C7654 a_71281_n10073.n261 VSS 0.431228f
C7655 a_71281_n10073.t317 VSS 0.41704f
C7656 a_71281_n10073.n262 VSS 0.425799f
C7657 a_71281_n10073.t68 VSS 0.377955f
C7658 a_71281_n10073.n263 VSS 0.425799f
C7659 a_71281_n10073.n264 VSS 0.046844f
C7660 a_71281_n10073.n265 VSS 0.01935f
C7661 a_71281_n10073.t231 VSS 0.417015f
C7662 a_71281_n10073.t18 VSS 0.377866f
C7663 a_71281_n10073.n266 VSS 0.431228f
C7664 a_71281_n10073.n267 VSS 0.041724f
C7665 a_71281_n10073.n268 VSS 0.147642f
C7666 a_71281_n10073.t52 VSS 0.332539f
C7667 a_71281_n10073.n269 VSS 0.147642f
C7668 a_71281_n10073.n270 VSS 0.041724f
C7669 a_71281_n10073.n271 VSS 0.01935f
C7670 a_71281_n10073.n272 VSS 0.264461f
C7671 a_71281_n10073.n273 VSS 0.264461f
C7672 a_71281_n10073.n274 VSS 0.046844f
C7673 a_71281_n10073.n275 VSS 0.431228f
C7674 a_71281_n10073.t118 VSS 0.41704f
C7675 a_71281_n10073.n276 VSS 0.425799f
C7676 a_71281_n10073.t46 VSS 0.377955f
C7677 a_71281_n10073.n277 VSS 0.425799f
C7678 a_71281_n10073.n278 VSS 0.046844f
C7679 a_71281_n10073.n279 VSS 0.01935f
C7680 a_71281_n10073.t316 VSS 0.417015f
C7681 a_71281_n10073.t2 VSS 0.377866f
C7682 a_71281_n10073.n280 VSS 0.431228f
C7683 a_71281_n10073.n281 VSS 0.041724f
C7684 a_71281_n10073.n282 VSS 0.147642f
C7685 a_71281_n10073.t24 VSS 0.332539f
C7686 a_71281_n10073.n283 VSS 0.147642f
C7687 a_71281_n10073.n284 VSS 0.041724f
C7688 a_71281_n10073.n285 VSS 0.01935f
C7689 a_71281_n10073.n286 VSS 0.218874f
C7690 a_71281_n10073.t47 VSS 0.157278f
C7691 a_71281_n10073.t25 VSS 0.033171f
C7692 a_71281_n10073.t3 VSS 0.033171f
C7693 a_71281_n10073.n287 VSS 0.135406f
C7694 a_71281_n10073.n288 VSS 0.378573f
C7695 a_71281_n10073.n289 VSS 0.091758f
C7696 a_71281_n10073.n290 VSS 0.218874f
C7697 a_71281_n10073.n291 VSS 0.046844f
C7698 a_71281_n10073.n292 VSS 0.431228f
C7699 a_71281_n10073.t93 VSS 0.41704f
C7700 a_71281_n10073.n293 VSS 0.425799f
C7701 a_71281_n10073.t143 VSS 0.377955f
C7702 a_71281_n10073.n294 VSS 0.425799f
C7703 a_71281_n10073.n295 VSS 0.046844f
C7704 a_71281_n10073.n296 VSS 0.01935f
C7705 a_71281_n10073.t284 VSS 0.417015f
C7706 a_71281_n10073.t295 VSS 0.377866f
C7707 a_71281_n10073.n297 VSS 0.431228f
C7708 a_71281_n10073.n298 VSS 0.041724f
C7709 a_71281_n10073.n299 VSS 0.147642f
C7710 a_71281_n10073.t194 VSS 0.332539f
C7711 a_71281_n10073.n300 VSS 0.147642f
C7712 a_71281_n10073.n301 VSS 0.041724f
C7713 a_71281_n10073.n302 VSS 0.01935f
C7714 a_71281_n10073.n303 VSS 0.265045f
C7715 a_71281_n10073.n304 VSS 0.264461f
C7716 a_71281_n10073.n305 VSS 0.046844f
C7717 a_71281_n10073.n306 VSS 0.431228f
C7718 a_71281_n10073.t159 VSS 0.41704f
C7719 a_71281_n10073.n307 VSS 0.425799f
C7720 a_71281_n10073.t209 VSS 0.377955f
C7721 a_71281_n10073.n308 VSS 0.425799f
C7722 a_71281_n10073.n309 VSS 0.046844f
C7723 a_71281_n10073.n310 VSS 0.01935f
C7724 a_71281_n10073.t89 VSS 0.417015f
C7725 a_71281_n10073.t102 VSS 0.377866f
C7726 a_71281_n10073.n311 VSS 0.431228f
C7727 a_71281_n10073.n312 VSS 0.041724f
C7728 a_71281_n10073.n313 VSS 0.147642f
C7729 a_71281_n10073.t276 VSS 0.332539f
C7730 a_71281_n10073.n314 VSS 0.147642f
C7731 a_71281_n10073.n315 VSS 0.041724f
C7732 a_71281_n10073.n316 VSS 0.01935f
C7733 a_71281_n10073.n317 VSS 0.264461f
C7734 a_71281_n10073.n318 VSS 0.264168f
C7735 a_71281_n10073.n319 VSS 0.046844f
C7736 a_71281_n10073.n320 VSS 0.431228f
C7737 a_71281_n10073.t150 VSS 0.41704f
C7738 a_71281_n10073.n321 VSS 0.425799f
C7739 a_71281_n10073.t199 VSS 0.377955f
C7740 a_71281_n10073.n322 VSS 0.425799f
C7741 a_71281_n10073.n323 VSS 0.046844f
C7742 a_71281_n10073.n324 VSS 0.01935f
C7743 a_71281_n10073.t83 VSS 0.417015f
C7744 a_71281_n10073.t95 VSS 0.377866f
C7745 a_71281_n10073.n325 VSS 0.431228f
C7746 a_71281_n10073.n326 VSS 0.041724f
C7747 a_71281_n10073.n327 VSS 0.147642f
C7748 a_71281_n10073.t269 VSS 0.332539f
C7749 a_71281_n10073.n328 VSS 0.147642f
C7750 a_71281_n10073.n329 VSS 0.041724f
C7751 a_71281_n10073.n330 VSS 0.01935f
C7752 a_71281_n10073.n331 VSS 0.264168f
C7753 a_71281_n10073.n332 VSS 0.264461f
C7754 a_71281_n10073.n333 VSS 0.046844f
C7755 a_71281_n10073.n334 VSS 0.431228f
C7756 a_71281_n10073.t218 VSS 0.413932f
C7757 a_71281_n10073.n335 VSS 0.425799f
C7758 a_71281_n10073.t283 VSS 0.377955f
C7759 a_71281_n10073.n336 VSS 0.415054f
C7760 a_71281_n10073.n337 VSS 0.046844f
C7761 a_71281_n10073.n338 VSS 0.01935f
C7762 a_71281_n10073.t149 VSS 0.417015f
C7763 a_71281_n10073.t162 VSS 0.377866f
C7764 a_71281_n10073.n339 VSS 0.431228f
C7765 a_71281_n10073.n340 VSS 0.041724f
C7766 a_71281_n10073.n341 VSS 0.147642f
C7767 a_71281_n10073.t78 VSS 0.332539f
C7768 a_71281_n10073.n342 VSS 0.147642f
C7769 a_71281_n10073.n343 VSS 0.041724f
C7770 a_71281_n10073.n344 VSS 0.01935f
C7771 a_71281_n10073.n345 VSS 0.600807f
C7772 a_71281_n10073.n346 VSS 0.050894f
C7773 a_71281_n10073.n347 VSS 0.046844f
C7774 a_71281_n10073.n348 VSS 0.431228f
C7775 a_71281_n10073.t325 VSS 0.413932f
C7776 a_71281_n10073.n349 VSS 0.415054f
C7777 a_71281_n10073.t201 VSS 0.377955f
C7778 a_71281_n10073.n350 VSS 0.425799f
C7779 a_71281_n10073.n351 VSS 0.046844f
C7780 a_71281_n10073.t291 VSS 0.417015f
C7781 a_71281_n10073.t308 VSS 0.377866f
C7782 a_71281_n10073.n352 VSS 0.431228f
C7783 a_71281_n10073.n353 VSS 0.041724f
C7784 a_71281_n10073.n354 VSS 0.147642f
C7785 a_71281_n10073.t331 VSS 0.332539f
C7786 a_71281_n10073.n355 VSS 0.147642f
C7787 a_71281_n10073.n356 VSS 0.041724f
C7788 a_71281_n10073.n357 VSS 0.01935f
C7789 a_71281_n10073.n358 VSS 0.527768f
C7790 a_71281_n10073.n359 VSS 0.264168f
C7791 a_71281_n10073.n360 VSS 0.046844f
C7792 a_71281_n10073.n361 VSS 0.431228f
C7793 a_71281_n10073.t249 VSS 0.41704f
C7794 a_71281_n10073.n362 VSS 0.425799f
C7795 a_71281_n10073.t137 VSS 0.377955f
C7796 a_71281_n10073.n363 VSS 0.425799f
C7797 a_71281_n10073.n364 VSS 0.046844f
C7798 a_71281_n10073.t212 VSS 0.417015f
C7799 a_71281_n10073.t224 VSS 0.377866f
C7800 a_71281_n10073.n365 VSS 0.431228f
C7801 a_71281_n10073.n366 VSS 0.01935f
C7802 a_71281_n10073.n367 VSS 0.041724f
C7803 a_71281_n10073.n368 VSS 0.147642f
C7804 a_71281_n10073.t252 VSS 0.332539f
C7805 a_71281_n10073.n369 VSS 0.147642f
C7806 a_71281_n10073.n370 VSS 0.041724f
C7807 a_71281_n10073.n371 VSS 0.01935f
C7808 a_71281_n10073.n372 VSS 0.264168f
C7809 a_71281_n10073.n373 VSS 0.264461f
C7810 a_71281_n10073.n374 VSS 0.046844f
C7811 a_71281_n10073.n375 VSS 0.431228f
C7812 a_71281_n10073.t113 VSS 0.41704f
C7813 a_71281_n10073.n376 VSS 0.425799f
C7814 a_71281_n10073.t273 VSS 0.377955f
C7815 a_71281_n10073.n377 VSS 0.425799f
C7816 a_71281_n10073.n378 VSS 0.046844f
C7817 a_71281_n10073.t87 VSS 0.417015f
C7818 a_71281_n10073.t99 VSS 0.377866f
C7819 a_71281_n10073.n379 VSS 0.431228f
C7820 a_71281_n10073.n380 VSS 0.01935f
C7821 a_71281_n10073.n381 VSS 0.041724f
C7822 a_71281_n10073.n382 VSS 0.147642f
C7823 a_71281_n10073.t115 VSS 0.332539f
C7824 a_71281_n10073.n383 VSS 0.147642f
C7825 a_71281_n10073.n384 VSS 0.041724f
C7826 a_71281_n10073.n385 VSS 0.01935f
C7827 a_71281_n10073.n386 VSS 0.264461f
C7828 a_71281_n10073.n387 VSS 0.265045f
C7829 a_71281_n10073.n388 VSS 0.046844f
C7830 a_71281_n10073.n389 VSS 0.431228f
C7831 a_71281_n10073.t311 VSS 0.41704f
C7832 a_71281_n10073.n390 VSS 0.425799f
C7833 a_71281_n10073.t191 VSS 0.377955f
C7834 a_71281_n10073.n391 VSS 0.425799f
C7835 a_71281_n10073.n392 VSS 0.046844f
C7836 a_71281_n10073.t280 VSS 0.417015f
C7837 a_71281_n10073.t287 VSS 0.377866f
C7838 a_71281_n10073.n393 VSS 0.431228f
C7839 a_71281_n10073.n394 VSS 0.01935f
C7840 a_71281_n10073.n395 VSS 0.041724f
C7841 a_71281_n10073.n396 VSS 0.147642f
C7842 a_71281_n10073.t314 VSS 0.332539f
C7843 a_71281_n10073.n397 VSS 0.147642f
C7844 a_71281_n10073.n398 VSS 0.041724f
C7845 a_71281_n10073.n399 VSS 0.01935f
C7846 a_71281_n10073.n400 VSS 0.218874f
C7847 a_71281_n10073.t35 VSS 0.157278f
C7848 a_71281_n10073.t5 VSS 0.033171f
C7849 a_71281_n10073.t7 VSS 0.033171f
C7850 a_71281_n10073.n401 VSS 0.135406f
C7851 a_71281_n10073.n402 VSS 0.378573f
C7852 a_71281_n10073.n403 VSS 0.091758f
C7853 a_71281_n10073.n404 VSS 0.218874f
C7854 a_71281_n10073.n405 VSS 0.046844f
C7855 a_71281_n10073.n406 VSS 0.431228f
C7856 a_71281_n10073.t320 VSS 0.41704f
C7857 a_71281_n10073.n407 VSS 0.425799f
C7858 a_71281_n10073.t34 VSS 0.377955f
C7859 a_71281_n10073.n408 VSS 0.425799f
C7860 a_71281_n10073.n409 VSS 0.046844f
C7861 a_71281_n10073.t286 VSS 0.417015f
C7862 a_71281_n10073.t6 VSS 0.377866f
C7863 a_71281_n10073.n410 VSS 0.431228f
C7864 a_71281_n10073.n411 VSS 0.01935f
C7865 a_71281_n10073.n412 VSS 0.041724f
C7866 a_71281_n10073.n413 VSS 0.147642f
C7867 a_71281_n10073.t4 VSS 0.332539f
C7868 a_71281_n10073.n414 VSS 0.147642f
C7869 a_71281_n10073.n415 VSS 0.041724f
C7870 a_71281_n10073.n416 VSS 0.01935f
C7871 a_71281_n10073.n417 VSS 0.264461f
C7872 a_71281_n10073.n418 VSS 0.264461f
C7873 a_71281_n10073.n419 VSS 0.046844f
C7874 a_71281_n10073.n420 VSS 0.431228f
C7875 a_71281_n10073.t240 VSS 0.41704f
C7876 a_71281_n10073.n421 VSS 0.425799f
C7877 a_71281_n10073.t56 VSS 0.377955f
C7878 a_71281_n10073.n422 VSS 0.425799f
C7879 a_71281_n10073.n423 VSS 0.046844f
C7880 a_71281_n10073.t206 VSS 0.417015f
C7881 a_71281_n10073.t26 VSS 0.377866f
C7882 a_71281_n10073.n424 VSS 0.431228f
C7883 a_71281_n10073.n425 VSS 0.01935f
C7884 a_71281_n10073.n426 VSS 0.041724f
C7885 a_71281_n10073.n427 VSS 0.147642f
C7886 a_71281_n10073.t20 VSS 0.332539f
C7887 a_71281_n10073.n428 VSS 0.147642f
C7888 a_71281_n10073.n429 VSS 0.041724f
C7889 a_71281_n10073.n430 VSS 0.01935f
C7890 a_71281_n10073.n431 VSS 0.218582f
C7891 a_71281_n10073.t57 VSS 0.033171f
C7892 a_71281_n10073.t21 VSS 0.033171f
C7893 a_71281_n10073.n432 VSS 0.135177f
C7894 a_71281_n10073.t27 VSS 0.157501f
C7895 a_71281_n10073.n433 VSS 0.380031f
C7896 a_71281_n10073.n434 VSS 0.091758f
C7897 a_71281_n10073.n435 VSS 0.21829f
C7898 a_71281_n10073.n436 VSS 0.046844f
C7899 a_71281_n10073.n437 VSS 0.431228f
C7900 a_71281_n10073.t253 VSS 0.41704f
C7901 a_71281_n10073.n438 VSS 0.425799f
C7902 a_71281_n10073.t144 VSS 0.377955f
C7903 a_71281_n10073.n439 VSS 0.425799f
C7904 a_71281_n10073.n440 VSS 0.046844f
C7905 a_71281_n10073.t219 VSS 0.417015f
C7906 a_71281_n10073.t234 VSS 0.377866f
C7907 a_71281_n10073.n441 VSS 0.431228f
C7908 a_71281_n10073.n442 VSS 0.01935f
C7909 a_71281_n10073.n443 VSS 0.041724f
C7910 a_71281_n10073.n444 VSS 0.147642f
C7911 a_71281_n10073.t257 VSS 0.332539f
C7912 a_71281_n10073.n445 VSS 0.147642f
C7913 a_71281_n10073.n446 VSS 0.041724f
C7914 a_71281_n10073.n447 VSS 0.01935f
C7915 a_71281_n10073.n448 VSS 0.264168f
C7916 a_71281_n10073.n449 VSS 0.264461f
C7917 a_71281_n10073.n450 VSS 0.046844f
C7918 a_71281_n10073.n451 VSS 0.431228f
C7919 a_71281_n10073.t242 VSS 0.41704f
C7920 a_71281_n10073.n452 VSS 0.425799f
C7921 a_71281_n10073.t133 VSS 0.377955f
C7922 a_71281_n10073.n453 VSS 0.425799f
C7923 a_71281_n10073.n454 VSS 0.046844f
C7924 a_71281_n10073.t207 VSS 0.417015f
C7925 a_71281_n10073.t222 VSS 0.377866f
C7926 a_71281_n10073.n455 VSS 0.431228f
C7927 a_71281_n10073.n456 VSS 0.01935f
C7928 a_71281_n10073.n457 VSS 0.041724f
C7929 a_71281_n10073.n458 VSS 0.147642f
C7930 a_71281_n10073.t245 VSS 0.332539f
C7931 a_71281_n10073.n459 VSS 0.147642f
C7932 a_71281_n10073.n460 VSS 0.041724f
C7933 a_71281_n10073.n461 VSS 0.01935f
C7934 a_71281_n10073.n462 VSS 0.264461f
C7935 a_71281_n10073.n463 VSS 0.265045f
C7936 a_71281_n10073.n464 VSS 0.046844f
C7937 a_71281_n10073.n465 VSS 0.431228f
C7938 a_71281_n10073.t264 VSS 0.41704f
C7939 a_71281_n10073.n466 VSS 0.425799f
C7940 a_71281_n10073.t156 VSS 0.377955f
C7941 a_71281_n10073.n467 VSS 0.425799f
C7942 a_71281_n10073.n468 VSS 0.046844f
C7943 a_71281_n10073.t243 VSS 0.417015f
C7944 a_71281_n10073.t256 VSS 0.377866f
C7945 a_71281_n10073.n469 VSS 0.431228f
C7946 a_71281_n10073.n470 VSS 0.01935f
C7947 a_71281_n10073.n471 VSS 0.041724f
C7948 a_71281_n10073.n472 VSS 0.147642f
C7949 a_71281_n10073.t266 VSS 0.332539f
C7950 a_71281_n10073.n473 VSS 0.147642f
C7951 a_71281_n10073.n474 VSS 0.041724f
C7952 a_71281_n10073.n475 VSS 0.01935f
C7953 a_71281_n10073.n476 VSS 0.265045f
C7954 a_71281_n10073.n477 VSS 0.264461f
C7955 a_71281_n10073.n478 VSS 0.046844f
C7956 a_71281_n10073.n479 VSS 0.431228f
C7957 a_71281_n10073.t186 VSS 0.41704f
C7958 a_71281_n10073.n480 VSS 0.425799f
C7959 a_71281_n10073.t91 VSS 0.377955f
C7960 a_71281_n10073.n481 VSS 0.425799f
C7961 a_71281_n10073.n482 VSS 0.046844f
C7962 a_71281_n10073.n483 VSS 0.01935f
C7963 a_71281_n10073.t170 VSS 0.417015f
C7964 a_71281_n10073.t175 VSS 0.377866f
C7965 a_71281_n10073.n484 VSS 0.431228f
C7966 a_71281_n10073.n485 VSS 0.041724f
C7967 a_71281_n10073.n486 VSS 0.147642f
C7968 a_71281_n10073.t188 VSS 0.332539f
C7969 a_71281_n10073.n487 VSS 0.147642f
C7970 a_71281_n10073.n488 VSS 0.041724f
C7971 a_71281_n10073.n489 VSS 0.01935f
C7972 a_71281_n10073.n490 VSS 0.59847f
C7973 a_71281_n10073.n491 VSS 2.21256f
C7974 a_71281_n10073.n492 VSS 0.051957f
C7975 a_71281_n10073.n493 VSS 0.046844f
C7976 a_71281_n10073.n494 VSS 0.431228f
C7977 a_71281_n10073.t130 VSS 0.41704f
C7978 a_71281_n10073.n495 VSS 0.425799f
C7979 a_71281_n10073.t160 VSS 0.377955f
C7980 a_71281_n10073.n496 VSS 0.425799f
C7981 a_71281_n10073.n497 VSS 0.046844f
C7982 a_71281_n10073.t304 VSS 0.417015f
C7983 a_71281_n10073.t271 VSS 0.377866f
C7984 a_71281_n10073.n498 VSS 0.431228f
C7985 a_71281_n10073.n499 VSS 0.041724f
C7986 a_71281_n10073.n500 VSS 0.147642f
C7987 a_71281_n10073.t258 VSS 0.332539f
C7988 a_71281_n10073.n501 VSS 0.147642f
C7989 a_71281_n10073.n502 VSS 0.041724f
C7990 a_71281_n10073.n503 VSS 0.01935f
C7991 a_71281_n10073.n504 VSS 0.536641f
C7992 a_71281_n10073.n505 VSS 0.265045f
C7993 a_71281_n10073.n506 VSS 0.046844f
C7994 a_71281_n10073.n507 VSS 0.431228f
C7995 a_71281_n10073.t195 VSS 0.41704f
C7996 a_71281_n10073.n508 VSS 0.425799f
C7997 a_71281_n10073.t233 VSS 0.377955f
C7998 a_71281_n10073.n509 VSS 0.425799f
C7999 a_71281_n10073.n510 VSS 0.046844f
C8000 a_71281_n10073.n511 VSS 0.01935f
C8001 a_71281_n10073.t109 VSS 0.417015f
C8002 a_71281_n10073.t80 VSS 0.377866f
C8003 a_71281_n10073.n512 VSS 0.431228f
C8004 a_71281_n10073.n513 VSS 0.041724f
C8005 a_71281_n10073.n514 VSS 0.147642f
C8006 a_71281_n10073.t335 VSS 0.332539f
C8007 a_71281_n10073.n515 VSS 0.147642f
C8008 a_71281_n10073.n516 VSS 0.041724f
C8009 a_71281_n10073.n517 VSS 0.01935f
C8010 a_71281_n10073.n518 VSS 0.265045f
C8011 a_71281_n10073.n519 VSS 0.264461f
C8012 a_71281_n10073.n520 VSS 0.046844f
C8013 a_71281_n10073.n521 VSS 0.431228f
C8014 a_71281_n10073.t189 VSS 0.41704f
C8015 a_71281_n10073.n522 VSS 0.425799f
C8016 a_71281_n10073.t220 VSS 0.377955f
C8017 a_71281_n10073.n523 VSS 0.425799f
C8018 a_71281_n10073.n524 VSS 0.046844f
C8019 a_71281_n10073.n525 VSS 0.01935f
C8020 a_71281_n10073.t100 VSS 0.417015f
C8021 a_71281_n10073.t75 VSS 0.377866f
C8022 a_71281_n10073.n526 VSS 0.431228f
C8023 a_71281_n10073.n527 VSS 0.041724f
C8024 a_71281_n10073.n528 VSS 0.147642f
C8025 a_71281_n10073.t326 VSS 0.332539f
C8026 a_71281_n10073.n529 VSS 0.147642f
C8027 a_71281_n10073.n530 VSS 0.041724f
C8028 a_71281_n10073.n531 VSS 0.01935f
C8029 a_71281_n10073.n532 VSS 0.264461f
C8030 a_71281_n10073.n533 VSS 0.264168f
C8031 a_71281_n10073.n534 VSS 0.046844f
C8032 a_71281_n10073.n535 VSS 0.431228f
C8033 a_71281_n10073.t270 VSS 0.41704f
C8034 a_71281_n10073.n536 VSS 0.425799f
C8035 a_71281_n10073.t303 VSS 0.377955f
C8036 a_71281_n10073.n537 VSS 0.425799f
C8037 a_71281_n10073.n538 VSS 0.046844f
C8038 a_71281_n10073.n539 VSS 0.01935f
C8039 a_71281_n10073.t169 VSS 0.417015f
C8040 a_71281_n10073.t134 VSS 0.377866f
C8041 a_71281_n10073.n540 VSS 0.431228f
C8042 a_71281_n10073.n541 VSS 0.041724f
C8043 a_71281_n10073.n542 VSS 0.147642f
C8044 a_71281_n10073.t123 VSS 0.332539f
C8045 a_71281_n10073.n543 VSS 0.147642f
C8046 a_71281_n10073.n544 VSS 0.041724f
C8047 a_71281_n10073.n545 VSS 0.01935f
C8048 a_71281_n10073.n546 VSS 0.21829f
C8049 a_71281_n10073.t13 VSS 0.033171f
C8050 a_71281_n10073.t65 VSS 0.033171f
C8051 a_71281_n10073.n547 VSS 0.135177f
C8052 a_71281_n10073.t59 VSS 0.157501f
C8053 a_71281_n10073.n548 VSS 0.380031f
C8054 a_71281_n10073.n549 VSS 0.091758f
C8055 a_71281_n10073.n550 VSS 0.218582f
C8056 a_71281_n10073.n551 VSS 0.046844f
C8057 a_71281_n10073.n552 VSS 0.431228f
C8058 a_71281_n10073.t267 VSS 0.41704f
C8059 a_71281_n10073.n553 VSS 0.425799f
C8060 a_71281_n10073.t12 VSS 0.377955f
C8061 a_71281_n10073.n554 VSS 0.425799f
C8062 a_71281_n10073.n555 VSS 0.046844f
C8063 a_71281_n10073.n556 VSS 0.01935f
C8064 a_71281_n10073.t154 VSS 0.417015f
C8065 a_71281_n10073.t58 VSS 0.377866f
C8066 a_71281_n10073.n557 VSS 0.431228f
C8067 a_71281_n10073.n558 VSS 0.041724f
C8068 a_71281_n10073.n559 VSS 0.147642f
C8069 a_71281_n10073.t64 VSS 0.332539f
C8070 a_71281_n10073.n560 VSS 0.147642f
C8071 a_71281_n10073.n561 VSS 0.041724f
C8072 a_71281_n10073.n562 VSS 0.01935f
C8073 a_71281_n10073.n563 VSS 0.264461f
C8074 a_71281_n10073.n564 VSS 0.264461f
C8075 a_71281_n10073.n565 VSS 0.046844f
C8076 a_71281_n10073.n566 VSS 0.431228f
C8077 a_71281_n10073.t74 VSS 0.41704f
C8078 a_71281_n10073.n567 VSS 0.425799f
C8079 a_71281_n10073.t70 VSS 0.377955f
C8080 a_71281_n10073.n568 VSS 0.425799f
C8081 a_71281_n10073.n569 VSS 0.046844f
C8082 a_71281_n10073.n570 VSS 0.01935f
C8083 a_71281_n10073.t227 VSS 0.417015f
C8084 a_71281_n10073.t36 VSS 0.377866f
C8085 a_71281_n10073.n571 VSS 0.431228f
C8086 a_71281_n10073.n572 VSS 0.041724f
C8087 a_71281_n10073.n573 VSS 0.147642f
C8088 a_71281_n10073.t42 VSS 0.332539f
C8089 a_71281_n10073.n574 VSS 0.147642f
C8090 a_71281_n10073.n575 VSS 0.041724f
C8091 a_71281_n10073.n576 VSS 0.01935f
C8092 a_71281_n10073.n577 VSS 0.218874f
C8093 a_71281_n10073.t71 VSS 0.157278f
C8094 a_71281_n10073.t43 VSS 0.033171f
C8095 a_71281_n10073.t37 VSS 0.033171f
C8096 a_71281_n10073.n578 VSS 0.135406f
C8097 a_71281_n10073.n579 VSS 0.378573f
C8098 a_71281_n10073.n580 VSS 0.091758f
C8099 a_71281_n10073.n581 VSS 0.218874f
C8100 a_71281_n10073.n582 VSS 0.046844f
C8101 a_71281_n10073.n583 VSS 0.431228f
C8102 a_71281_n10073.t323 VSS 0.41704f
C8103 a_71281_n10073.n584 VSS 0.425799f
C8104 a_71281_n10073.t77 VSS 0.377955f
C8105 a_71281_n10073.n585 VSS 0.425799f
C8106 a_71281_n10073.n586 VSS 0.046844f
C8107 a_71281_n10073.n587 VSS 0.01935f
C8108 a_71281_n10073.t198 VSS 0.417015f
C8109 a_71281_n10073.t182 VSS 0.377866f
C8110 a_71281_n10073.n588 VSS 0.431228f
C8111 a_71281_n10073.n589 VSS 0.041724f
C8112 a_71281_n10073.n590 VSS 0.147642f
C8113 a_71281_n10073.t158 VSS 0.332539f
C8114 a_71281_n10073.n591 VSS 0.147642f
C8115 a_71281_n10073.n592 VSS 0.041724f
C8116 a_71281_n10073.n593 VSS 0.01935f
C8117 a_71281_n10073.n594 VSS 0.265045f
C8118 a_71281_n10073.n595 VSS 0.264461f
C8119 a_71281_n10073.n596 VSS 0.046844f
C8120 a_71281_n10073.n597 VSS 0.431228f
C8121 a_71281_n10073.t122 VSS 0.41704f
C8122 a_71281_n10073.n598 VSS 0.425799f
C8123 a_71281_n10073.t141 VSS 0.377955f
C8124 a_71281_n10073.n599 VSS 0.425799f
C8125 a_71281_n10073.n600 VSS 0.046844f
C8126 a_71281_n10073.n601 VSS 0.01935f
C8127 a_71281_n10073.t281 VSS 0.417015f
C8128 a_71281_n10073.t262 VSS 0.377866f
C8129 a_71281_n10073.n602 VSS 0.431228f
C8130 a_71281_n10073.n603 VSS 0.041724f
C8131 a_71281_n10073.n604 VSS 0.147642f
C8132 a_71281_n10073.t229 VSS 0.332539f
C8133 a_71281_n10073.n605 VSS 0.147642f
C8134 a_71281_n10073.n606 VSS 0.041724f
C8135 a_71281_n10073.n607 VSS 0.01935f
C8136 a_71281_n10073.n608 VSS 0.264461f
C8137 a_71281_n10073.n609 VSS 0.264168f
C8138 a_71281_n10073.n610 VSS 0.046844f
C8139 a_71281_n10073.n611 VSS 0.431228f
C8140 a_71281_n10073.t117 VSS 0.41704f
C8141 a_71281_n10073.n612 VSS 0.425799f
C8142 a_71281_n10073.t131 VSS 0.377955f
C8143 a_71281_n10073.n613 VSS 0.425799f
C8144 a_71281_n10073.n614 VSS 0.046844f
C8145 a_71281_n10073.n615 VSS 0.01935f
C8146 a_71281_n10073.t272 VSS 0.417015f
C8147 a_71281_n10073.t255 VSS 0.377866f
C8148 a_71281_n10073.n616 VSS 0.431228f
C8149 a_71281_n10073.n617 VSS 0.041724f
C8150 a_71281_n10073.n618 VSS 0.147642f
C8151 a_71281_n10073.t217 VSS 0.332539f
C8152 a_71281_n10073.n619 VSS 0.147642f
C8153 a_71281_n10073.n620 VSS 0.041724f
C8154 a_71281_n10073.n621 VSS 0.01935f
C8155 a_71281_n10073.n622 VSS 0.264168f
C8156 a_71281_n10073.n623 VSS 0.264461f
C8157 a_71281_n10073.n624 VSS 0.046844f
C8158 a_71281_n10073.n625 VSS 0.431228f
C8159 a_71281_n10073.t181 VSS 0.413932f
C8160 a_71281_n10073.n626 VSS 0.425799f
C8161 a_71281_n10073.t197 VSS 0.377955f
C8162 a_71281_n10073.n627 VSS 0.415054f
C8163 a_71281_n10073.n628 VSS 0.046844f
C8164 a_71281_n10073.n629 VSS 0.01935f
C8165 a_71281_n10073.t82 VSS 0.417015f
C8166 a_71281_n10073.t334 VSS 0.377866f
C8167 a_71281_n10073.n630 VSS 0.431228f
C8168 a_71281_n10073.n631 VSS 0.041724f
C8169 a_71281_n10073.n632 VSS 0.147642f
C8170 a_71281_n10073.t301 VSS 0.332539f
C8171 a_71281_n10073.n633 VSS 0.147642f
C8172 a_71281_n10073.n634 VSS 0.041724f
C8173 a_71281_n10073.n635 VSS 0.01935f
C8174 a_71281_n10073.n636 VSS 0.600807f
C8175 a_71281_n10073.n637 VSS 0.050894f
C8176 a_71281_n10073.n638 VSS 0.046844f
C8177 a_71281_n10073.n639 VSS 0.431228f
C8178 a_71281_n10073.t202 VSS 0.413932f
C8179 a_71281_n10073.n640 VSS 0.415054f
C8180 a_71281_n10073.t226 VSS 0.377955f
C8181 a_71281_n10073.n641 VSS 0.425799f
C8182 a_71281_n10073.n642 VSS 0.046844f
C8183 a_71281_n10073.t319 VSS 0.417015f
C8184 a_71281_n10073.t292 VSS 0.377866f
C8185 a_71281_n10073.n643 VSS 0.431228f
C8186 a_71281_n10073.n644 VSS 0.041724f
C8187 a_71281_n10073.n645 VSS 0.147642f
C8188 a_71281_n10073.t205 VSS 0.332539f
C8189 a_71281_n10073.n646 VSS 0.147642f
C8190 a_71281_n10073.n647 VSS 0.041724f
C8191 a_71281_n10073.n648 VSS 0.01935f
C8192 a_71281_n10073.n649 VSS 0.527768f
C8193 a_71281_n10073.n650 VSS 0.264168f
C8194 a_71281_n10073.n651 VSS 0.046844f
C8195 a_71281_n10073.n652 VSS 0.431228f
C8196 a_71281_n10073.t138 VSS 0.41704f
C8197 a_71281_n10073.n653 VSS 0.425799f
C8198 a_71281_n10073.t153 VSS 0.377955f
C8199 a_71281_n10073.n654 VSS 0.425799f
C8200 a_71281_n10073.n655 VSS 0.046844f
C8201 a_71281_n10073.t237 VSS 0.417015f
C8202 a_71281_n10073.t213 VSS 0.377866f
C8203 a_71281_n10073.n656 VSS 0.431228f
C8204 a_71281_n10073.n657 VSS 0.01935f
C8205 a_71281_n10073.n658 VSS 0.041724f
C8206 a_71281_n10073.n659 VSS 0.147642f
C8207 a_71281_n10073.t140 VSS 0.332539f
C8208 a_71281_n10073.n660 VSS 0.147642f
C8209 a_71281_n10073.n661 VSS 0.041724f
C8210 a_71281_n10073.n662 VSS 0.01935f
C8211 a_71281_n10073.n663 VSS 0.264168f
C8212 a_71281_n10073.n664 VSS 0.264461f
C8213 a_71281_n10073.n665 VSS 0.046844f
C8214 a_71281_n10073.n666 VSS 0.431228f
C8215 a_71281_n10073.t274 VSS 0.41704f
C8216 a_71281_n10073.n667 VSS 0.425799f
C8217 a_71281_n10073.t289 VSS 0.377955f
C8218 a_71281_n10073.n668 VSS 0.425799f
C8219 a_71281_n10073.n669 VSS 0.046844f
C8220 a_71281_n10073.t107 VSS 0.417015f
C8221 a_71281_n10073.t88 VSS 0.377866f
C8222 a_71281_n10073.n670 VSS 0.431228f
C8223 a_71281_n10073.n671 VSS 0.01935f
C8224 a_71281_n10073.n672 VSS 0.041724f
C8225 a_71281_n10073.n673 VSS 0.147642f
C8226 a_71281_n10073.t275 VSS 0.332539f
C8227 a_71281_n10073.n674 VSS 0.147642f
C8228 a_71281_n10073.n675 VSS 0.041724f
C8229 a_71281_n10073.n676 VSS 0.01935f
C8230 a_71281_n10073.n677 VSS 0.264461f
C8231 a_71281_n10073.n678 VSS 0.265045f
C8232 a_71281_n10073.n679 VSS 0.046844f
C8233 a_71281_n10073.n680 VSS 0.431228f
C8234 a_71281_n10073.t192 VSS 0.41704f
C8235 a_71281_n10073.n681 VSS 0.425799f
C8236 a_71281_n10073.t211 VSS 0.377955f
C8237 a_71281_n10073.n682 VSS 0.425799f
C8238 a_71281_n10073.n683 VSS 0.046844f
C8239 a_71281_n10073.t302 VSS 0.417015f
C8240 a_71281_n10073.t282 VSS 0.377866f
C8241 a_71281_n10073.n684 VSS 0.431228f
C8242 a_71281_n10073.n685 VSS 0.01935f
C8243 a_71281_n10073.n686 VSS 0.041724f
C8244 a_71281_n10073.n687 VSS 0.147642f
C8245 a_71281_n10073.t193 VSS 0.332539f
C8246 a_71281_n10073.n688 VSS 0.147642f
C8247 a_71281_n10073.n689 VSS 0.041724f
C8248 a_71281_n10073.n690 VSS 0.01935f
C8249 a_71281_n10073.n691 VSS 0.218874f
C8250 a_71281_n10073.t23 VSS 0.157278f
C8251 a_71281_n10073.t33 VSS 0.033171f
C8252 a_71281_n10073.t11 VSS 0.033171f
C8253 a_71281_n10073.n692 VSS 0.135406f
C8254 a_71281_n10073.n693 VSS 0.378573f
C8255 a_71281_n10073.n694 VSS 0.091758f
C8256 a_71281_n10073.n695 VSS 0.218874f
C8257 a_71281_n10073.n696 VSS 0.046844f
C8258 a_71281_n10073.n697 VSS 0.431228f
C8259 a_71281_n10073.t200 VSS 0.41704f
C8260 a_71281_n10073.n698 VSS 0.425799f
C8261 a_71281_n10073.t22 VSS 0.377955f
C8262 a_71281_n10073.n699 VSS 0.425799f
C8263 a_71281_n10073.n700 VSS 0.046844f
C8264 a_71281_n10073.t315 VSS 0.417015f
C8265 a_71281_n10073.t10 VSS 0.377866f
C8266 a_71281_n10073.n701 VSS 0.431228f
C8267 a_71281_n10073.n702 VSS 0.01935f
C8268 a_71281_n10073.n703 VSS 0.041724f
C8269 a_71281_n10073.n704 VSS 0.147642f
C8270 a_71281_n10073.t32 VSS 0.332539f
C8271 a_71281_n10073.n705 VSS 0.147642f
C8272 a_71281_n10073.n706 VSS 0.041724f
C8273 a_71281_n10073.n707 VSS 0.01935f
C8274 a_71281_n10073.n708 VSS 0.264461f
C8275 a_71281_n10073.n709 VSS 0.264461f
C8276 a_71281_n10073.n710 VSS 0.046844f
C8277 a_71281_n10073.n711 VSS 0.431228f
C8278 a_71281_n10073.t132 VSS 0.41704f
C8279 a_71281_n10073.n712 VSS 0.425799f
C8280 a_71281_n10073.t50 VSS 0.377955f
C8281 a_71281_n10073.n713 VSS 0.425799f
C8282 a_71281_n10073.n714 VSS 0.046844f
C8283 a_71281_n10073.t230 VSS 0.417015f
C8284 a_71281_n10073.t28 VSS 0.377866f
C8285 a_71281_n10073.n715 VSS 0.431228f
C8286 a_71281_n10073.n716 VSS 0.01935f
C8287 a_71281_n10073.n717 VSS 0.041724f
C8288 a_71281_n10073.n718 VSS 0.147642f
C8289 a_71281_n10073.t54 VSS 0.332539f
C8290 a_71281_n10073.n719 VSS 0.147642f
C8291 a_71281_n10073.n720 VSS 0.041724f
C8292 a_71281_n10073.n721 VSS 0.01935f
C8293 a_71281_n10073.n722 VSS 0.218582f
C8294 a_71281_n10073.t51 VSS 0.033171f
C8295 a_71281_n10073.t55 VSS 0.033171f
C8296 a_71281_n10073.n723 VSS 0.135177f
C8297 a_71281_n10073.t29 VSS 0.157501f
C8298 a_71281_n10073.n724 VSS 0.380031f
C8299 a_71281_n10073.n725 VSS 0.091758f
C8300 a_71281_n10073.n726 VSS 0.21829f
C8301 a_71281_n10073.n727 VSS 0.046844f
C8302 a_71281_n10073.n728 VSS 0.431228f
C8303 a_71281_n10073.t145 VSS 0.41704f
C8304 a_71281_n10073.n729 VSS 0.425799f
C8305 a_71281_n10073.t165 VSS 0.377955f
C8306 a_71281_n10073.n730 VSS 0.425799f
C8307 a_71281_n10073.n731 VSS 0.046844f
C8308 a_71281_n10073.t246 VSS 0.417015f
C8309 a_71281_n10073.t221 VSS 0.377866f
C8310 a_71281_n10073.n732 VSS 0.431228f
C8311 a_71281_n10073.n733 VSS 0.01935f
C8312 a_71281_n10073.n734 VSS 0.041724f
C8313 a_71281_n10073.n735 VSS 0.147642f
C8314 a_71281_n10073.t147 VSS 0.332539f
C8315 a_71281_n10073.n736 VSS 0.147642f
C8316 a_71281_n10073.n737 VSS 0.041724f
C8317 a_71281_n10073.n738 VSS 0.01935f
C8318 a_71281_n10073.n739 VSS 0.264168f
C8319 a_71281_n10073.n740 VSS 0.264461f
C8320 a_71281_n10073.n741 VSS 0.046844f
C8321 a_71281_n10073.n742 VSS 0.431228f
C8322 a_71281_n10073.t135 VSS 0.41704f
C8323 a_71281_n10073.n743 VSS 0.425799f
C8324 a_71281_n10073.t151 VSS 0.377955f
C8325 a_71281_n10073.n744 VSS 0.425799f
C8326 a_71281_n10073.n745 VSS 0.046844f
C8327 a_71281_n10073.t232 VSS 0.417015f
C8328 a_71281_n10073.t208 VSS 0.377866f
C8329 a_71281_n10073.n746 VSS 0.431228f
C8330 a_71281_n10073.n747 VSS 0.01935f
C8331 a_71281_n10073.n748 VSS 0.041724f
C8332 a_71281_n10073.n749 VSS 0.147642f
C8333 a_71281_n10073.t136 VSS 0.332539f
C8334 a_71281_n10073.n750 VSS 0.147642f
C8335 a_71281_n10073.n751 VSS 0.041724f
C8336 a_71281_n10073.n752 VSS 0.01935f
C8337 a_71281_n10073.n753 VSS 0.264461f
C8338 a_71281_n10073.n754 VSS 0.265045f
C8339 a_71281_n10073.n755 VSS 0.046844f
C8340 a_71281_n10073.n756 VSS 0.431228f
C8341 a_71281_n10073.t157 VSS 0.41704f
C8342 a_71281_n10073.n757 VSS 0.425799f
C8343 a_71281_n10073.t176 VSS 0.377955f
C8344 a_71281_n10073.n758 VSS 0.425799f
C8345 a_71281_n10073.n759 VSS 0.046844f
C8346 a_71281_n10073.t263 VSS 0.417015f
C8347 a_71281_n10073.t244 VSS 0.377866f
C8348 a_71281_n10073.n760 VSS 0.431228f
C8349 a_71281_n10073.n761 VSS 0.01935f
C8350 a_71281_n10073.n762 VSS 0.041724f
C8351 a_71281_n10073.n763 VSS 0.147642f
C8352 a_71281_n10073.t164 VSS 0.332539f
C8353 a_71281_n10073.n764 VSS 0.147642f
C8354 a_71281_n10073.n765 VSS 0.041724f
C8355 a_71281_n10073.n766 VSS 0.01935f
C8356 a_71281_n10073.n767 VSS 0.265045f
C8357 a_71281_n10073.n768 VSS 0.264461f
C8358 a_71281_n10073.n769 VSS 0.046844f
C8359 a_71281_n10073.n770 VSS 0.431228f
C8360 a_71281_n10073.t92 VSS 0.41704f
C8361 a_71281_n10073.n771 VSS 0.425799f
C8362 a_71281_n10073.t111 VSS 0.377955f
C8363 a_71281_n10073.n772 VSS 0.425799f
C8364 a_71281_n10073.n773 VSS 0.046844f
C8365 a_71281_n10073.n774 VSS 0.01935f
C8366 a_71281_n10073.t184 VSS 0.417015f
C8367 a_71281_n10073.t171 VSS 0.377866f
C8368 a_71281_n10073.n775 VSS 0.431228f
C8369 a_71281_n10073.n776 VSS 0.041724f
C8370 a_71281_n10073.n777 VSS 0.147642f
C8371 a_71281_n10073.t97 VSS 0.332539f
C8372 a_71281_n10073.n778 VSS 0.147642f
C8373 a_71281_n10073.n779 VSS 0.041724f
C8374 a_71281_n10073.n780 VSS 0.01935f
C8375 a_71281_n10073.n781 VSS 0.59847f
C8376 a_71281_n10073.n782 VSS 0.853871f
C8377 a_71281_n10073.n783 VSS 2.36947f
C8378 a_71281_n10073.t0 VSS 0.078987f
C8379 a_71281_n10073.t1 VSS 0.080021f
C8380 a_71281_n10073.n784 VSS 5.12344f
C8381 a_71281_n10073.n785 VSS 0.853871f
C8382 a_71281_n10073.n786 VSS 0.600807f
C8383 a_71281_n10073.n787 VSS 0.046844f
C8384 a_71281_n10073.n788 VSS 0.431228f
C8385 a_71281_n10073.t214 VSS 0.413932f
C8386 a_71281_n10073.n789 VSS 0.415054f
C8387 a_71281_n10073.t277 VSS 0.377955f
C8388 a_71281_n10073.n790 VSS 0.425799f
C8389 a_71281_n10073.n791 VSS 0.046844f
C8390 a_71281_n10073.t146 VSS 0.417015f
C8391 a_71281_n10073.t98 VSS 0.377866f
C8392 a_71281_n10073.n792 VSS 0.431228f
C8393 a_71281_n10073.n793 VSS 0.01935f
C8394 a_71281_n10073.n794 VSS 0.041724f
C8395 a_71281_n10073.n795 VSS 0.147642f
C8396 a_71281_n10073.t307 VSS 0.332539f
C8397 a_71281_n10073.n796 VSS 0.147642f
C8398 a_71281_n10073.n797 VSS 0.041724f
C8399 a_71281_n10073.n798 VSS 0.01935f
C8400 a_71281_n10073.n799 VSS 0.264461f
C8401 a_71281_n10073.n800 VSS 0.264168f
C8402 a_71281_n10073.n801 VSS 0.046844f
C8403 a_71281_n10073.n802 VSS 0.431228f
C8404 a_71281_n10073.t148 VSS 0.41704f
C8405 a_71281_n10073.n803 VSS 0.425799f
C8406 a_71281_n10073.t196 VSS 0.377955f
C8407 a_71281_n10073.n804 VSS 0.425799f
C8408 a_71281_n10073.n805 VSS 0.046844f
C8409 a_71281_n10073.t81 VSS 0.417015f
C8410 a_71281_n10073.t285 VSS 0.377866f
C8411 a_71281_n10073.n806 VSS 0.431228f
C8412 a_71281_n10073.n807 VSS 0.01935f
C8413 a_71281_n10073.n808 VSS 0.041724f
C8414 a_71281_n10073.n809 VSS 0.147642f
C8415 a_71281_n10073.t223 VSS 0.332539f
C8416 a_71281_n10073.n810 VSS 0.147642f
C8417 a_71281_n10073.n811 VSS 0.041724f
C8418 a_71281_n10073.n812 VSS 0.01935f
C8419 a_71281_n10073.n813 VSS 0.264168f
C8420 a_71281_n10073.n814 VSS 0.264461f
C8421 a_71281_n10073.n815 VSS 0.046844f
C8422 a_71281_n10073.n816 VSS 0.431228f
C8423 a_71281_n10073.t152 VSS 0.41704f
C8424 a_71281_n10073.n817 VSS 0.425799f
C8425 a_71281_n10073.t203 VSS 0.377955f
C8426 a_71281_n10073.n818 VSS 0.425799f
C8427 a_71281_n10073.n819 VSS 0.046844f
C8428 a_71281_n10073.t85 VSS 0.417015f
C8429 a_71281_n10073.t297 VSS 0.377866f
C8430 a_71281_n10073.n820 VSS 0.431228f
C8431 a_71281_n10073.n821 VSS 0.01935f
C8432 a_71281_n10073.n822 VSS 0.041724f
C8433 a_71281_n10073.n823 VSS 0.147642f
C8434 a_71281_n10073.t236 VSS 0.332539f
C8435 a_71281_n10073.n824 VSS 0.147642f
C8436 a_71281_n10073.n825 VSS 0.041724f
C8437 a_71281_n10073.n826 VSS 0.01935f
C8438 a_71281_n10073.n827 VSS 0.264461f
C8439 a_71281_n10073.n828 VSS 0.265045f
C8440 a_71281_n10073.n829 VSS 0.046844f
C8441 a_71281_n10073.n830 VSS 0.431228f
C8442 a_71281_n10073.t86 VSS 0.41704f
C8443 a_71281_n10073.n831 VSS 0.425799f
C8444 a_71281_n10073.t139 VSS 0.377955f
C8445 a_71281_n10073.n832 VSS 0.425799f
C8446 a_71281_n10073.n833 VSS 0.046844f
C8447 a_71281_n10073.t279 VSS 0.417015f
C8448 a_71281_n10073.t215 VSS 0.377866f
C8449 a_71281_n10073.n834 VSS 0.431228f
C8450 a_71281_n10073.n835 VSS 0.01935f
C8451 a_71281_n10073.n836 VSS 0.041724f
C8452 a_71281_n10073.n837 VSS 0.147642f
C8453 a_71281_n10073.t166 VSS 0.332539f
C8454 a_71281_n10073.n838 VSS 0.147642f
C8455 a_71281_n10073.n839 VSS 0.041724f
C8456 a_71281_n10073.n840 VSS 0.01935f
C8457 a_71281_n10073.n841 VSS 0.218874f
C8458 a_71281_n10073.t49 VSS 0.157278f
C8459 a_71281_n10073.t41 VSS 0.033171f
C8460 a_71281_n10073.t17 VSS 0.033171f
C8461 a_71281_n10073.n842 VSS 0.135406f
C8462 a_71281_n10073.n843 VSS 0.378573f
C8463 a_71281_n10073.n844 VSS 0.091758f
C8464 a_71281_n10073.n845 VSS 0.218874f
C8465 a_71281_n10073.n846 VSS 0.046844f
C8466 a_71281_n10073.n847 VSS 0.431228f
C8467 a_71281_n10073.t114 VSS 0.41704f
C8468 a_71281_n10073.n848 VSS 0.425799f
C8469 a_71281_n10073.t48 VSS 0.377955f
C8470 a_71281_n10073.n849 VSS 0.425799f
C8471 a_71281_n10073.n850 VSS 0.046844f
C8472 a_71281_n10073.t310 VSS 0.417015f
C8473 a_71281_n10073.t16 VSS 0.377866f
C8474 a_71281_n10073.n851 VSS 0.431228f
C8475 a_71281_n10073.n852 VSS 0.01935f
C8476 a_71281_n10073.n853 VSS 0.041724f
C8477 a_71281_n10073.n854 VSS 0.147642f
C8478 a_71281_n10073.t40 VSS 0.332539f
C8479 a_71281_n10073.n855 VSS 0.147642f
C8480 a_71281_n10073.n856 VSS 0.041724f
C8481 a_71281_n10073.n857 VSS 0.01935f
C8482 a_71281_n10073.n858 VSS 0.264461f
C8483 a_71281_n10073.n859 VSS 0.264461f
C8484 a_71281_n10073.n860 VSS 0.046844f
C8485 a_71281_n10073.n861 VSS 0.431228f
C8486 a_71281_n10073.t312 VSS 0.41704f
C8487 a_71281_n10073.n862 VSS 0.425799f
C8488 a_71281_n10073.t72 VSS 0.377955f
C8489 a_71281_n10073.n863 VSS 0.425799f
C8490 a_71281_n10073.n864 VSS 0.046844f
C8491 a_71281_n10073.t225 VSS 0.417015f
C8492 a_71281_n10073.t44 VSS 0.377866f
C8493 a_71281_n10073.n865 VSS 0.431228f
C8494 a_71281_n10073.n866 VSS 0.01935f
C8495 a_71281_n10073.n867 VSS 0.041724f
C8496 a_71281_n10073.n868 VSS 0.147642f
C8497 a_71281_n10073.t62 VSS 0.332539f
C8498 a_71281_n10073.n869 VSS 0.147642f
C8499 a_71281_n10073.n870 VSS 0.041724f
C8500 a_71281_n10073.n871 VSS 0.01935f
C8501 a_71281_n10073.n872 VSS 0.218582f
C8502 a_71281_n10073.n873 VSS 0.091758f
C8503 a_71281_n10073.n874 VSS 0.380031f
C8504 a_71281_n10073.n875 VSS 0.135177f
C8505 a_71281_n10073.t73 VSS 0.033171f
C8506 a_45445_n19595.t1 VSS 68.227104f
C8507 a_45445_n19595.t2 VSS 2.67562f
C8508 a_45445_n19595.t0 VSS 18.1973f
C8509 a_33379_34917.n0 VSS 3.81673f
C8510 a_33379_34917.n1 VSS 1.71606f
C8511 a_33379_34917.n2 VSS 0.239374f
C8512 a_33379_34917.n3 VSS 0.251463f
C8513 a_33379_34917.n4 VSS 0.363149f
C8514 a_33379_34917.n5 VSS 0.002078f
C8515 a_33379_34917.n6 VSS 0.177139f
C8516 a_33379_34917.t0 VSS 1.07595f
C8517 a_33379_34917.n7 VSS 0.151788f
C8518 a_33379_34917.n8 VSS 0.153725f
C8519 a_33379_34917.t68 VSS 0.221873p
C8520 a_33379_34917.t60 VSS 0.018975f
C8521 a_33379_34917.t46 VSS 0.018975f
C8522 a_33379_34917.t90 VSS 0.018975f
C8523 a_33379_34917.t51 VSS 0.018975f
C8524 a_33379_34917.t83 VSS 0.018975f
C8525 a_33379_34917.t30 VSS 0.018975f
C8526 a_33379_34917.t7 VSS 0.018975f
C8527 a_33379_34917.t59 VSS 0.018975f
C8528 a_33379_34917.t5 VSS 0.018975f
C8529 a_33379_34917.t56 VSS 0.018975f
C8530 a_33379_34917.t66 VSS 0.018975f
C8531 a_33379_34917.t63 VSS 0.018975f
C8532 a_33379_34917.t4 VSS 0.018975f
C8533 a_33379_34917.t26 VSS 0.018975f
C8534 a_33379_34917.t52 VSS 0.018975f
C8535 a_33379_34917.t76 VSS 0.018975f
C8536 a_33379_34917.t91 VSS 0.018975f
C8537 a_33379_34917.t48 VSS 0.018975f
C8538 a_33379_34917.t43 VSS 0.018975f
C8539 a_33379_34917.t84 VSS 0.018975f
C8540 a_33379_34917.t13 VSS 0.018975f
C8541 a_33379_34917.t40 VSS 0.018975f
C8542 a_33379_34917.t81 VSS 0.018975f
C8543 a_33379_34917.t31 VSS 0.018975f
C8544 a_33379_34917.t15 VSS 0.018975f
C8545 a_33379_34917.t74 VSS 0.018975f
C8546 a_33379_34917.t16 VSS 0.018975f
C8547 a_33379_34917.t34 VSS 0.018975f
C8548 a_33379_34917.t53 VSS 0.018975f
C8549 a_33379_34917.t50 VSS 0.018975f
C8550 a_33379_34917.t25 VSS 0.018975f
C8551 a_33379_34917.t80 VSS 0.018975f
C8552 a_33379_34917.t54 VSS 0.018975f
C8553 a_33379_34917.t69 VSS 0.018975f
C8554 a_33379_34917.t42 VSS 0.018975f
C8555 a_33379_34917.t17 VSS 0.018975f
C8556 a_33379_34917.t88 VSS 0.018975f
C8557 a_33379_34917.t72 VSS 0.018975f
C8558 a_33379_34917.t9 VSS 0.018975f
C8559 a_33379_34917.t64 VSS 0.018975f
C8560 a_33379_34917.t75 VSS 0.018975f
C8561 a_33379_34917.t8 VSS 0.018975f
C8562 a_33379_34917.t35 VSS 0.018975f
C8563 a_33379_34917.t14 VSS 0.018975f
C8564 a_33379_34917.t41 VSS 0.018975f
C8565 a_33379_34917.t3 VSS 0.018975f
C8566 a_33379_34917.t37 VSS 0.018975f
C8567 a_33379_34917.t10 VSS 0.018975f
C8568 a_33379_34917.t70 VSS 0.018975f
C8569 a_33379_34917.t11 VSS 0.018975f
C8570 a_33379_34917.t32 VSS 0.018975f
C8571 a_33379_34917.t65 VSS 0.018975f
C8572 a_33379_34917.t73 VSS 0.018975f
C8573 a_33379_34917.t45 VSS 0.018975f
C8574 a_33379_34917.t39 VSS 0.018975f
C8575 a_33379_34917.t19 VSS 0.018975f
C8576 a_33379_34917.t62 VSS 0.018975f
C8577 a_33379_34917.t86 VSS 0.018975f
C8578 a_33379_34917.t29 VSS 0.018975f
C8579 a_33379_34917.t58 VSS 0.018975f
C8580 a_33379_34917.t87 VSS 0.018975f
C8581 a_33379_34917.t33 VSS 0.018975f
C8582 a_33379_34917.t23 VSS 0.018975f
C8583 a_33379_34917.t79 VSS 0.018975f
C8584 a_33379_34917.t24 VSS 0.018975f
C8585 a_33379_34917.t38 VSS 0.018975f
C8586 a_33379_34917.t71 VSS 0.018975f
C8587 a_33379_34917.t27 VSS 0.018975f
C8588 a_33379_34917.t85 VSS 0.018975f
C8589 a_33379_34917.t18 VSS 0.018975f
C8590 a_33379_34917.t89 VSS 0.018975f
C8591 a_33379_34917.t77 VSS 0.018975f
C8592 a_33379_34917.t82 VSS 0.018975f
C8593 a_33379_34917.t57 VSS 0.018975f
C8594 a_33379_34917.t28 VSS 0.018975f
C8595 a_33379_34917.t6 VSS 0.018975f
C8596 a_33379_34917.t20 VSS 0.018975f
C8597 a_33379_34917.t67 VSS 0.018975f
C8598 a_33379_34917.t49 VSS 0.018975f
C8599 a_33379_34917.t44 VSS 0.018975f
C8600 a_33379_34917.t61 VSS 0.018975f
C8601 a_33379_34917.t55 VSS 0.018975f
C8602 a_33379_34917.t12 VSS 0.018975f
C8603 a_33379_34917.t47 VSS 0.018975f
C8604 a_33379_34917.t78 VSS 0.018975f
C8605 a_33379_34917.t22 VSS 0.018975f
C8606 a_33379_34917.t36 VSS 0.018975f
C8607 a_33379_34917.t21 VSS 0.018975f
C8608 a_33379_34917.t1 VSS 0.022797f
C8609 a_33379_34917.t2 VSS 0.019444f
C8610 a_33379_34917.n9 VSS 1.76731f
C8611 a_51711_n5344.t1 VSS 1.26787f
C8612 a_51711_n5344.t0 VSS 1.23213f
C8613 a_31831_n5342.t0 VSS 5.871891f
C8614 a_31831_n5342.t1 VSS 49.2433f
C8615 a_31831_n5342.t2 VSS 31.4848f
C8616 a_32913_n8930.t1 VSS 63.4564f
C8617 a_32913_n8930.t2 VSS 2.38382f
C8618 a_32913_n8930.t0 VSS 26.3598f
C8619 a_30152_10448.t3 VSS 20.5853f
C8620 a_30152_10448.t0 VSS 1.77451f
C8621 a_30152_10448.t9 VSS 0.34777f
C8622 a_30152_10448.t2 VSS 0.330207f
C8623 a_30152_10448.t1 VSS 0.329925f
C8624 a_30152_10448.t14 VSS 0.568066f
C8625 a_30152_10448.t21 VSS 0.544019f
C8626 a_30152_10448.t20 VSS 0.544019f
C8627 a_30152_10448.t4 VSS 0.562597f
C8628 a_30152_10448.t19 VSS 0.568066f
C8629 a_30152_10448.t13 VSS 0.544019f
C8630 a_30152_10448.t6 VSS 0.568066f
C8631 a_30152_10448.t17 VSS 0.544019f
C8632 a_30152_10448.t15 VSS 0.544019f
C8633 a_30152_10448.t22 VSS 0.562597f
C8634 a_30152_10448.t7 VSS 0.34777f
C8635 a_30152_10448.t11 VSS 0.30485f
C8636 a_30152_10448.t10 VSS 0.562597f
C8637 a_30152_10448.t12 VSS 0.544019f
C8638 a_30152_10448.t8 VSS 0.568066f
C8639 a_30152_10448.t18 VSS 0.544019f
C8640 a_30152_10448.t23 VSS 0.562597f
C8641 a_30152_10448.t16 VSS 0.544019f
C8642 a_30152_10448.t5 VSS 0.30485f
C8643 a_71342_4481.n0 VSS 9.95668f
C8644 a_71342_4481.t3 VSS 0.922601f
C8645 a_71342_4481.t1 VSS 0.704006f
C8646 a_71342_4481.t0 VSS 0.606767f
C8647 a_71342_4481.t2 VSS 0.50995f
C8648 a_71496_10388.n0 VSS 2.53786f
C8649 a_71496_10388.n1 VSS 9.92737f
C8650 a_71496_10388.n2 VSS 0.941685f
C8651 a_71496_10388.n3 VSS 1.60401f
C8652 a_71496_10388.n4 VSS 5.88445f
C8653 a_71496_10388.n5 VSS 7.950201f
C8654 a_71496_10388.n6 VSS 0.911776f
C8655 a_71496_10388.t16 VSS 0.572368f
C8656 a_71496_10388.t20 VSS 0.572572f
C8657 a_71496_10388.t18 VSS 0.605719f
C8658 a_71496_10388.t15 VSS 0.571949f
C8659 a_71496_10388.t6 VSS 0.347081f
C8660 a_71496_10388.t12 VSS 0.563936f
C8661 a_71496_10388.t14 VSS 0.563895f
C8662 a_71496_10388.t23 VSS 0.561709f
C8663 a_71496_10388.t11 VSS 0.561709f
C8664 a_71496_10388.t9 VSS 0.561709f
C8665 a_71496_10388.t22 VSS 0.561709f
C8666 a_71496_10388.t10 VSS 0.563801f
C8667 a_71496_10388.t19 VSS 0.563957f
C8668 a_71496_10388.t21 VSS 0.561709f
C8669 a_71496_10388.t8 VSS 0.561709f
C8670 a_71496_10388.t17 VSS 0.561709f
C8671 a_71496_10388.t13 VSS 0.561709f
C8672 a_71496_10388.t5 VSS 0.523342f
C8673 a_71496_10388.t2 VSS 0.599013f
C8674 a_71496_10388.t1 VSS 0.321546f
C8675 a_71496_10388.t3 VSS 0.32663f
C8676 a_71496_10388.t0 VSS 0.498545f
C8677 a_71496_10388.t7 VSS 0.526042f
C8678 a_71496_10388.n7 VSS 0.912682f
C8679 a_71496_10388.t4 VSS 0.315882f
C8680 a_100992_4421.t0 VSS 25.151001f
C8681 a_100992_4421.t1 VSS 13.2043f
C8682 a_100992_4421.t2 VSS 1.14464f
C8683 a_38097_n5342.t0 VSS 5.82902f
C8684 a_38097_n5342.t1 VSS 45.8437f
C8685 a_38097_n5342.t2 VSS 34.8273f
C8686 a_100992_n29313.t0 VSS 23.122198f
C8687 a_100992_n29313.t2 VSS 8.80583f
C8688 a_100992_n29313.t1 VSS 7.57194f
C8689 a_31284_n30339.t0 VSS 6.7139f
C8690 a_31284_n30339.t1 VSS 50.219196f
C8691 a_31284_n30339.t2 VSS 26.6669f
C8692 a_30324_n30399.t1 VSS 45.1766f
C8693 a_30324_n30399.t2 VSS 1.60691f
C8694 a_30324_n30399.t0 VSS 6.01645f
C8695 OUT.t50 VSS 0.043976f
C8696 OUT.t45 VSS 0.043976f
C8697 OUT.n0 VSS 0.096683f
C8698 OUT.n1 VSS 0.057699f
C8699 OUT.n2 VSS 0.386484f
C8700 OUT.n3 VSS 0.025967f
C8701 OUT.t78 VSS 0.131502f
C8702 OUT.n4 VSS 0.20405f
C8703 OUT.n5 VSS 0.025967f
C8704 OUT.t76 VSS 0.043976f
C8705 OUT.t52 VSS 0.043976f
C8706 OUT.n6 VSS 0.130054f
C8707 OUT.n7 VSS 0.157333f
C8708 OUT.t81 VSS 0.343659f
C8709 OUT.n8 VSS 0.845976f
C8710 OUT.n9 VSS 0.057699f
C8711 OUT.n10 VSS 0.154755f
C8712 OUT.n11 VSS 1.93161f
C8713 OUT.t109 VSS 7.241391f
C8714 OUT.t108 VSS 10.055799f
C8715 OUT.n12 VSS 21.947802f
C8716 OUT.t1 VSS 0.434784f
C8717 OUT.t0 VSS 0.418838f
C8718 OUT.n13 VSS 20.055302f
C8719 OUT.n14 VSS 40.5919f
C8720 OUT.n15 VSS 1.90125f
C8721 OUT.t67 VSS 0.043976f
C8722 OUT.t105 VSS 0.043976f
C8723 OUT.n16 VSS 0.422694f
C8724 OUT.t85 VSS 0.197725f
C8725 OUT.n17 VSS 1.13405f
C8726 OUT.t69 VSS 0.043976f
C8727 OUT.t26 VSS 0.043976f
C8728 OUT.n18 VSS 0.422694f
C8729 OUT.t93 VSS 0.197725f
C8730 OUT.n19 VSS 1.13405f
C8731 OUT.n20 VSS 1.17727f
C8732 OUT.t95 VSS 0.115858f
C8733 OUT.t107 VSS 0.123364f
C8734 OUT.n21 VSS 0.468341f
C8735 OUT.t44 VSS 0.043976f
C8736 OUT.t94 VSS 0.043976f
C8737 OUT.n22 VSS 0.111591f
C8738 OUT.t48 VSS 0.043976f
C8739 OUT.t106 VSS 0.043976f
C8740 OUT.n23 VSS 0.120432f
C8741 OUT.n24 VSS 0.305656f
C8742 OUT.n25 VSS 0.254719f
C8743 OUT.t65 VSS 0.043976f
C8744 OUT.t98 VSS 0.043976f
C8745 OUT.n26 VSS 0.20307f
C8746 OUT.n27 VSS 0.996211f
C8747 OUT.t68 VSS 0.197725f
C8748 OUT.n28 VSS 0.928666f
C8749 OUT.n29 VSS 2.86532f
C8750 OUT.n30 VSS 0.120993f
C8751 OUT.t75 VSS 0.115858f
C8752 OUT.t79 VSS 0.123364f
C8753 OUT.n31 VSS 0.390598f
C8754 OUT.n32 VSS 0.300976f
C8755 OUT.t104 VSS 0.115858f
C8756 OUT.t27 VSS 0.123364f
C8757 OUT.n33 VSS 0.388979f
C8758 OUT.n34 VSS 0.356044f
C8759 OUT.t58 VSS 0.043976f
C8760 OUT.t36 VSS 0.043976f
C8761 OUT.n35 VSS 0.111591f
C8762 OUT.t63 VSS 0.043976f
C8763 OUT.t40 VSS 0.043976f
C8764 OUT.n36 VSS 0.120432f
C8765 OUT.n37 VSS 0.305656f
C8766 OUT.n38 VSS 0.238723f
C8767 OUT.t22 VSS 0.115858f
C8768 OUT.t34 VSS 0.123364f
C8769 OUT.n39 VSS 0.394785f
C8770 OUT.n40 VSS 0.362483f
C8771 OUT.t91 VSS 0.115858f
C8772 OUT.t100 VSS 0.123364f
C8773 OUT.n41 VSS 0.394785f
C8774 OUT.n42 VSS 0.362496f
C8775 OUT.t49 VSS 0.043976f
C8776 OUT.t23 VSS 0.043976f
C8777 OUT.n43 VSS 0.111591f
C8778 OUT.t57 VSS 0.043976f
C8779 OUT.t35 VSS 0.043976f
C8780 OUT.n44 VSS 0.120432f
C8781 OUT.n45 VSS 0.305656f
C8782 OUT.n46 VSS 0.169975f
C8783 OUT.t37 VSS 0.115858f
C8784 OUT.t41 VSS 0.123364f
C8785 OUT.n47 VSS 0.467878f
C8786 OUT.t72 VSS 0.043976f
C8787 OUT.t59 VSS 0.043976f
C8788 OUT.n48 VSS 0.111591f
C8789 OUT.t77 VSS 0.043976f
C8790 OUT.t64 VSS 0.043976f
C8791 OUT.n49 VSS 0.120432f
C8792 OUT.n50 VSS 0.305656f
C8793 OUT.n51 VSS 0.322916f
C8794 OUT.t33 VSS 0.115858f
C8795 OUT.t39 VSS 0.123364f
C8796 OUT.n52 VSS 0.388979f
C8797 OUT.n53 VSS 0.356044f
C8798 OUT.t29 VSS 0.115858f
C8799 OUT.t38 VSS 0.123364f
C8800 OUT.n54 VSS 0.390598f
C8801 OUT.n55 VSS 0.300976f
C8802 OUT.n56 VSS 0.120993f
C8803 OUT.n57 VSS 2.62673f
C8804 OUT.n58 VSS 0.025967f
C8805 OUT.n59 VSS 0.025967f
C8806 OUT.n60 VSS 0.386484f
C8807 OUT.t61 VSS 0.043976f
C8808 OUT.t55 VSS 0.043976f
C8809 OUT.n61 VSS 0.130054f
C8810 OUT.n62 VSS 0.157333f
C8811 OUT.n63 VSS 0.057699f
C8812 OUT.n64 VSS 0.106379f
C8813 OUT.n65 VSS 0.106381f
C8814 OUT.t82 VSS 0.131502f
C8815 OUT.n66 VSS 0.20405f
C8816 OUT.n67 VSS 0.057699f
C8817 OUT.n68 VSS 0.680579f
C8818 OUT.n69 VSS 0.025967f
C8819 OUT.t80 VSS 0.043976f
C8820 OUT.t62 VSS 0.043976f
C8821 OUT.n70 VSS 0.130054f
C8822 OUT.n71 VSS 0.157333f
C8823 OUT.t92 VSS 0.343659f
C8824 OUT.n72 VSS 0.845976f
C8825 OUT.n73 VSS 0.057699f
C8826 OUT.n74 VSS 0.154755f
C8827 OUT.n75 VSS 0.808529f
C8828 OUT.n76 VSS 1.66662f
C8829 OUT.n77 VSS 1.61549f
C8830 OUT.n78 VSS 0.835304f
C8831 OUT.t60 VSS 0.043976f
C8832 OUT.t90 VSS 0.043976f
C8833 OUT.n79 VSS 0.20307f
C8834 OUT.n80 VSS 0.996211f
C8835 OUT.t66 VSS 0.197725f
C8836 OUT.n81 VSS 0.655054f
C8837 OUT.n82 VSS 1.78572f
C8838 OUT.t87 VSS 0.115858f
C8839 OUT.t89 VSS 0.123364f
C8840 OUT.n83 VSS 0.468341f
C8841 OUT.t42 VSS 0.043976f
C8842 OUT.t86 VSS 0.043976f
C8843 OUT.n84 VSS 0.111591f
C8844 OUT.t43 VSS 0.043976f
C8845 OUT.t88 VSS 0.043976f
C8846 OUT.n85 VSS 0.120432f
C8847 OUT.n86 VSS 0.305656f
C8848 OUT.n87 VSS 0.254719f
C8849 OUT.t30 VSS 0.115858f
C8850 OUT.t32 VSS 0.123364f
C8851 OUT.n88 VSS 0.467878f
C8852 OUT.t70 VSS 0.043976f
C8853 OUT.t53 VSS 0.043976f
C8854 OUT.n89 VSS 0.111591f
C8855 OUT.t71 VSS 0.043976f
C8856 OUT.t56 VSS 0.043976f
C8857 OUT.n90 VSS 0.120432f
C8858 OUT.n91 VSS 0.305656f
C8859 OUT.n92 VSS 0.322916f
C8860 OUT.t24 VSS 0.115858f
C8861 OUT.t25 VSS 0.123364f
C8862 OUT.n93 VSS 0.388979f
C8863 OUT.n94 VSS 0.356044f
C8864 OUT.t20 VSS 0.115858f
C8865 OUT.t21 VSS 0.123364f
C8866 OUT.n95 VSS 0.390598f
C8867 OUT.n96 VSS 0.300976f
C8868 OUT.n97 VSS 0.120993f
C8869 OUT.t46 VSS 0.043976f
C8870 OUT.t101 VSS 0.043976f
C8871 OUT.n98 VSS 0.111591f
C8872 OUT.t47 VSS 0.043976f
C8873 OUT.t103 VSS 0.043976f
C8874 OUT.n99 VSS 0.120432f
C8875 OUT.n100 VSS 0.305656f
C8876 OUT.n101 VSS 0.169975f
C8877 OUT.t83 VSS 0.115858f
C8878 OUT.t84 VSS 0.123364f
C8879 OUT.n102 VSS 0.394785f
C8880 OUT.n103 VSS 0.362496f
C8881 OUT.t99 VSS 0.115858f
C8882 OUT.t102 VSS 0.123364f
C8883 OUT.n104 VSS 0.394785f
C8884 OUT.n105 VSS 0.362483f
C8885 OUT.t51 VSS 0.043976f
C8886 OUT.t28 VSS 0.043976f
C8887 OUT.n106 VSS 0.111591f
C8888 OUT.t54 VSS 0.043976f
C8889 OUT.t31 VSS 0.043976f
C8890 OUT.n107 VSS 0.120432f
C8891 OUT.n108 VSS 0.305656f
C8892 OUT.n109 VSS 0.238723f
C8893 OUT.t96 VSS 0.115858f
C8894 OUT.t97 VSS 0.123364f
C8895 OUT.n110 VSS 0.388979f
C8896 OUT.n111 VSS 0.356044f
C8897 OUT.t73 VSS 0.115858f
C8898 OUT.t74 VSS 0.123364f
C8899 OUT.n112 VSS 0.390598f
C8900 OUT.n113 VSS 0.300976f
C8901 OUT.n114 VSS 0.120993f
C8902 OUT.n115 VSS 1.93161f
C8903 OUT.n116 VSS 2.24453f
C8904 OUT.n117 VSS 5.82271f
C8905 OUT.n118 VSS 0.025967f
C8906 OUT.t10 VSS 0.041882f
C8907 OUT.t16 VSS 0.041882f
C8908 OUT.n119 VSS 0.121043f
C8909 OUT.n120 VSS 0.162555f
C8910 OUT.t4 VSS 0.31957f
C8911 OUT.n121 VSS 0.777903f
C8912 OUT.n122 VSS 0.057699f
C8913 OUT.n123 VSS 0.668995f
C8914 OUT.t19 VSS 0.041882f
C8915 OUT.t6 VSS 0.041882f
C8916 OUT.n124 VSS 0.104381f
C8917 OUT.t8 VSS 0.041882f
C8918 OUT.t14 VSS 0.041882f
C8919 OUT.n125 VSS 0.11243f
C8920 OUT.n126 VSS 0.375749f
C8921 OUT.t7 VSS 0.041882f
C8922 OUT.t13 VSS 0.041882f
C8923 OUT.n127 VSS 0.104381f
C8924 OUT.t15 VSS 0.041882f
C8925 OUT.t3 VSS 0.041882f
C8926 OUT.n128 VSS 0.11243f
C8927 OUT.n129 VSS 0.457073f
C8928 OUT.t9 VSS 0.115118f
C8929 OUT.t17 VSS 0.122142f
C8930 OUT.n130 VSS 0.375382f
C8931 OUT.n131 VSS 0.524479f
C8932 OUT.t11 VSS 0.115118f
C8933 OUT.t2 VSS 0.122142f
C8934 OUT.n132 VSS 0.377001f
C8935 OUT.n133 VSS 0.303489f
C8936 OUT.n134 VSS 0.288151f
C8937 OUT.n135 VSS 3.11177f
C8938 OUT.t5 VSS 0.041882f
C8939 OUT.t12 VSS 0.041882f
C8940 OUT.n136 VSS 0.376498f
C8941 OUT.t18 VSS 0.192513f
C8942 OUT.n137 VSS 1.31092f
C8943 OUT.n138 VSS 2.17189f
C8944 OUT.n139 VSS 2.93552f
C8945 OUT.n140 VSS 2.98586f
C8946 OUT.n141 VSS 0.808529f
C8947 OUT.n142 VSS 0.680579f
C8948 OUT.n143 VSS 0.057699f
C8949 OUT.n144 VSS 0.106381f
C8950 OUT.n145 VSS 0.106379f
C8951 OUT.n146 VSS 0.025967f
C8952 OUT.n147 VSS 0.058488f
C8953 a_33249_48695.n0 VSS 0.833973f
C8954 a_33249_48695.n1 VSS 0.724408f
C8955 a_33249_48695.n2 VSS 0.794543f
C8956 a_33249_48695.n3 VSS 0.542775f
C8957 a_33249_48695.n4 VSS 0.806163f
C8958 a_33249_48695.n5 VSS 0.806162f
C8959 a_33249_48695.n6 VSS 0.428084f
C8960 a_33249_48695.n7 VSS 0.724408f
C8961 a_33249_48695.n8 VSS 0.794543f
C8962 a_33249_48695.n9 VSS 0.94654f
C8963 a_33249_48695.n10 VSS 0.833973f
C8964 a_33249_48695.n11 VSS 0.724408f
C8965 a_33249_48695.n12 VSS 0.794543f
C8966 a_33249_48695.n13 VSS 0.542775f
C8967 a_33249_48695.n14 VSS 0.806163f
C8968 a_33249_48695.n15 VSS 0.806162f
C8969 a_33249_48695.n16 VSS 0.428084f
C8970 a_33249_48695.n17 VSS 0.724408f
C8971 a_33249_48695.n18 VSS 0.794543f
C8972 a_33249_48695.n19 VSS 0.94654f
C8973 a_33249_48695.n20 VSS 1.77855f
C8974 a_33249_48695.n21 VSS 1.25797f
C8975 a_33249_48695.n22 VSS 1.19957f
C8976 a_33249_48695.n23 VSS 1.77855f
C8977 a_33249_48695.n24 VSS 1.25797f
C8978 a_33249_48695.n25 VSS 0.915081f
C8979 a_33249_48695.n26 VSS 1.70465f
C8980 a_33249_48695.n27 VSS 1.49105f
C8981 a_33249_48695.n28 VSS 0.962832f
C8982 a_33249_48695.n29 VSS 1.70465f
C8983 a_33249_48695.n30 VSS 1.49105f
C8984 a_33249_48695.n31 VSS 0.962832f
C8985 a_33249_48695.n32 VSS 0.523558f
C8986 a_33249_48695.n33 VSS 0.842989f
C8987 a_33249_48695.n34 VSS 0.842982f
C8988 a_33249_48695.n35 VSS 0.820906f
C8989 a_33249_48695.n36 VSS 0.338474f
C8990 a_33249_48695.n37 VSS 0.842989f
C8991 a_33249_48695.n38 VSS 1.18777f
C8992 a_33249_48695.n39 VSS 1.05609f
C8993 a_33249_48695.n40 VSS 0.842989f
C8994 a_33249_48695.n41 VSS 0.842982f
C8995 a_33249_48695.n42 VSS 0.820906f
C8996 a_33249_48695.n43 VSS 0.338474f
C8997 a_33249_48695.n44 VSS 0.842989f
C8998 a_33249_48695.n45 VSS 1.18777f
C8999 a_33249_48695.t242 VSS 0.36917f
C9000 a_33249_48695.t202 VSS 0.065937f
C9001 a_33249_48695.t322 VSS 0.065937f
C9002 a_33249_48695.n46 VSS 0.285449f
C9003 a_33249_48695.n47 VSS 0.93961f
C9004 a_33249_48695.t264 VSS 0.279833f
C9005 a_33249_48695.n48 VSS 0.795316f
C9006 a_33249_48695.t256 VSS 0.065937f
C9007 a_33249_48695.t219 VSS 0.065937f
C9008 a_33249_48695.n49 VSS 0.285449f
C9009 a_33249_48695.n50 VSS 0.428366f
C9010 a_33249_48695.n51 VSS 2.69004f
C9011 a_33249_48695.t272 VSS 0.162517f
C9012 a_33249_48695.t318 VSS 0.198291f
C9013 a_33249_48695.n52 VSS 1.06267f
C9014 a_33249_48695.t214 VSS 0.065937f
C9015 a_33249_48695.t294 VSS 0.065937f
C9016 a_33249_48695.n53 VSS 0.154318f
C9017 a_33249_48695.t258 VSS 0.065937f
C9018 a_33249_48695.t164 VSS 0.065937f
C9019 a_33249_48695.n54 VSS 0.196324f
C9020 a_33249_48695.n55 VSS 0.446847f
C9021 a_33249_48695.n56 VSS 0.976786f
C9022 a_33249_48695.t161 VSS 0.279755f
C9023 a_33249_48695.n57 VSS 0.806849f
C9024 a_33249_48695.t317 VSS 0.277438f
C9025 a_33249_48695.n58 VSS 0.80029f
C9026 a_33249_48695.t262 VSS 0.065937f
C9027 a_33249_48695.t206 VSS 0.065937f
C9028 a_33249_48695.n59 VSS 0.285449f
C9029 a_33249_48695.n60 VSS 0.542569f
C9030 a_33249_48695.t325 VSS 0.279833f
C9031 a_33249_48695.n61 VSS 0.795271f
C9032 a_33249_48695.t213 VSS 0.277438f
C9033 a_33249_48695.n62 VSS 0.720574f
C9034 a_33249_48695.t176 VSS 0.374369f
C9035 a_33249_48695.t271 VSS 0.065937f
C9036 a_33249_48695.t211 VSS 0.065937f
C9037 a_33249_48695.n63 VSS 0.285449f
C9038 a_33249_48695.n64 VSS 0.837958f
C9039 a_33249_48695.n65 VSS 0.642415f
C9040 a_33249_48695.n66 VSS 3.12051f
C9041 a_33249_48695.t315 VSS 0.36917f
C9042 a_33249_48695.t275 VSS 0.065937f
C9043 a_33249_48695.t217 VSS 0.065937f
C9044 a_33249_48695.n67 VSS 0.285449f
C9045 a_33249_48695.n68 VSS 0.93961f
C9046 a_33249_48695.t165 VSS 0.279833f
C9047 a_33249_48695.n69 VSS 0.795271f
C9048 a_33249_48695.t227 VSS 0.277438f
C9049 a_33249_48695.n70 VSS 0.720574f
C9050 a_33249_48695.n71 VSS 2.09974f
C9051 a_33249_48695.t203 VSS 0.372643f
C9052 a_33249_48695.t166 VSS 0.065937f
C9053 a_33249_48695.t281 VSS 0.065937f
C9054 a_33249_48695.n72 VSS 0.284868f
C9055 a_33249_48695.t229 VSS 0.279265f
C9056 a_33249_48695.t293 VSS 0.278903f
C9057 a_33249_48695.t220 VSS 0.065937f
C9058 a_33249_48695.t179 VSS 0.065937f
C9059 a_33249_48695.n73 VSS 0.284868f
C9060 a_33249_48695.t297 VSS 0.279265f
C9061 a_33249_48695.t278 VSS 0.279265f
C9062 a_33249_48695.t224 VSS 0.065937f
C9063 a_33249_48695.t167 VSS 0.065937f
C9064 a_33249_48695.n74 VSS 0.284868f
C9065 a_33249_48695.t282 VSS 0.279265f
C9066 a_33249_48695.t178 VSS 0.278903f
C9067 a_33249_48695.t239 VSS 0.065937f
C9068 a_33249_48695.t177 VSS 0.065937f
C9069 a_33249_48695.n75 VSS 0.284868f
C9070 a_33249_48695.t313 VSS 0.373143f
C9071 a_33249_48695.n76 VSS 2.10814f
C9072 a_33249_48695.n77 VSS 2.64144f
C9073 a_33249_48695.t151 VSS 0.065937f
C9074 a_33249_48695.t112 VSS 0.065937f
C9075 a_33249_48695.n78 VSS 0.362253f
C9076 a_33249_48695.t3 VSS 0.065937f
C9077 a_33249_48695.t138 VSS 0.065937f
C9078 a_33249_48695.n79 VSS 0.241904f
C9079 a_33249_48695.n80 VSS 1.18974f
C9080 a_33249_48695.t347 VSS 0.065937f
C9081 a_33249_48695.t144 VSS 0.065937f
C9082 a_33249_48695.n81 VSS 0.241904f
C9083 a_33249_48695.n82 VSS 0.843784f
C9084 a_33249_48695.t115 VSS 0.065937f
C9085 a_33249_48695.t344 VSS 0.065937f
C9086 a_33249_48695.n83 VSS 0.241904f
C9087 a_33249_48695.n84 VSS 0.338896f
C9088 a_33249_48695.n85 VSS 2.52449f
C9089 a_33249_48695.n86 VSS 2.89625f
C9090 a_33249_48695.t253 VSS 0.065937f
C9091 a_33249_48695.t193 VSS 0.065937f
C9092 a_33249_48695.n87 VSS 0.306918f
C9093 a_33249_48695.t268 VSS 0.298209f
C9094 a_33249_48695.t265 VSS 0.065937f
C9095 a_33249_48695.t209 VSS 0.065937f
C9096 a_33249_48695.n88 VSS 0.306918f
C9097 a_33249_48695.t311 VSS 0.5404f
C9098 a_33249_48695.n89 VSS 2.49893f
C9099 a_33249_48695.t289 VSS 0.296468f
C9100 a_33249_48695.n90 VSS 1.39244f
C9101 a_33249_48695.t225 VSS 0.173717f
C9102 a_33249_48695.t267 VSS 0.184972f
C9103 a_33249_48695.n91 VSS 0.702229f
C9104 a_33249_48695.t186 VSS 0.065937f
C9105 a_33249_48695.t307 VSS 0.065937f
C9106 a_33249_48695.n92 VSS 0.16732f
C9107 a_33249_48695.t234 VSS 0.065937f
C9108 a_33249_48695.t174 VSS 0.065937f
C9109 a_33249_48695.n93 VSS 0.180576f
C9110 a_33249_48695.n94 VSS 0.4583f
C9111 a_33249_48695.n95 VSS 0.381925f
C9112 a_33249_48695.t163 VSS 0.173717f
C9113 a_33249_48695.t205 VSS 0.184972f
C9114 a_33249_48695.n96 VSS 0.701535f
C9115 a_33249_48695.t257 VSS 0.065937f
C9116 a_33249_48695.t195 VSS 0.065937f
C9117 a_33249_48695.n97 VSS 0.16732f
C9118 a_33249_48695.t301 VSS 0.065937f
C9119 a_33249_48695.t243 VSS 0.065937f
C9120 a_33249_48695.n98 VSS 0.180576f
C9121 a_33249_48695.n99 VSS 0.4583f
C9122 a_33249_48695.n100 VSS 0.484179f
C9123 a_33249_48695.t197 VSS 0.173717f
C9124 a_33249_48695.t244 VSS 0.184972f
C9125 a_33249_48695.n101 VSS 0.583234f
C9126 a_33249_48695.n102 VSS 0.533851f
C9127 a_33249_48695.t308 VSS 0.173717f
C9128 a_33249_48695.t175 VSS 0.184972f
C9129 a_33249_48695.n103 VSS 0.585662f
C9130 a_33249_48695.n104 VSS 0.451283f
C9131 a_33249_48695.t231 VSS 0.065937f
C9132 a_33249_48695.t310 VSS 0.065937f
C9133 a_33249_48695.n105 VSS 0.304483f
C9134 a_33249_48695.n106 VSS 1.49372f
C9135 a_33249_48695.t248 VSS 0.065937f
C9136 a_33249_48695.t172 VSS 0.065937f
C9137 a_33249_48695.n107 VSS 0.633787f
C9138 a_33249_48695.t306 VSS 0.296468f
C9139 a_33249_48695.n108 VSS 1.70039f
C9140 a_33249_48695.n109 VSS 1.7652f
C9141 a_33249_48695.n110 VSS 3.93851f
C9142 a_33249_48695.n111 VSS 0.181417f
C9143 a_33249_48695.t250 VSS 0.065937f
C9144 a_33249_48695.t189 VSS 0.065937f
C9145 a_33249_48695.n112 VSS 0.16732f
C9146 a_33249_48695.t292 VSS 0.065937f
C9147 a_33249_48695.t236 VSS 0.065937f
C9148 a_33249_48695.n113 VSS 0.180576f
C9149 a_33249_48695.n114 VSS 0.4583f
C9150 a_33249_48695.n115 VSS 0.25486f
C9151 a_33249_48695.t302 VSS 0.173717f
C9152 a_33249_48695.t170 VSS 0.184972f
C9153 a_33249_48695.n116 VSS 0.59194f
C9154 a_33249_48695.n117 VSS 0.543525f
C9155 a_33249_48695.t321 VSS 0.173717f
C9156 a_33249_48695.t187 VSS 0.184972f
C9157 a_33249_48695.n118 VSS 0.59194f
C9158 a_33249_48695.n119 VSS 0.543507f
C9159 a_33249_48695.t241 VSS 0.065937f
C9160 a_33249_48695.t201 VSS 0.065937f
C9161 a_33249_48695.n120 VSS 0.16732f
C9162 a_33249_48695.t283 VSS 0.065937f
C9163 a_33249_48695.t249 VSS 0.065937f
C9164 a_33249_48695.n121 VSS 0.180576f
C9165 a_33249_48695.n122 VSS 0.4583f
C9166 a_33249_48695.n123 VSS 0.357941f
C9167 a_33249_48695.t316 VSS 0.173717f
C9168 a_33249_48695.t182 VSS 0.184972f
C9169 a_33249_48695.n124 VSS 0.583234f
C9170 a_33249_48695.n125 VSS 0.533851f
C9171 a_33249_48695.t254 VSS 0.173717f
C9172 a_33249_48695.t296 VSS 0.184972f
C9173 a_33249_48695.n126 VSS 0.585662f
C9174 a_33249_48695.n127 VSS 0.451283f
C9175 a_33249_48695.n128 VSS 0.181417f
C9176 a_33249_48695.n129 VSS 4.29625f
C9177 a_33249_48695.t303 VSS 0.065937f
C9178 a_33249_48695.t245 VSS 0.065937f
C9179 a_33249_48695.n130 VSS 0.306918f
C9180 a_33249_48695.t324 VSS 0.298209f
C9181 a_33249_48695.t319 VSS 0.065937f
C9182 a_33249_48695.t259 VSS 0.065937f
C9183 a_33249_48695.n131 VSS 0.306918f
C9184 a_33249_48695.t183 VSS 0.5404f
C9185 a_33249_48695.n132 VSS 1.25177f
C9186 a_33249_48695.n133 VSS 2.87631f
C9187 a_33249_48695.n134 VSS 2.6775f
C9188 a_33249_48695.t184 VSS 0.296468f
C9189 a_33249_48695.n135 VSS 0.982186f
C9190 a_33249_48695.t304 VSS 0.065937f
C9191 a_33249_48695.t207 VSS 0.065937f
C9192 a_33249_48695.n136 VSS 0.304483f
C9193 a_33249_48695.n137 VSS 1.49372f
C9194 a_33249_48695.t320 VSS 0.065937f
C9195 a_33249_48695.t247 VSS 0.065937f
C9196 a_33249_48695.n138 VSS 0.633787f
C9197 a_33249_48695.t199 VSS 0.296468f
C9198 a_33249_48695.n139 VSS 1.70039f
C9199 a_33249_48695.n140 VSS 1.25245f
C9200 a_33249_48695.n141 VSS 2.42226f
C9201 a_33249_48695.t299 VSS 0.173717f
C9202 a_33249_48695.t221 VSS 0.184972f
C9203 a_33249_48695.n142 VSS 0.702229f
C9204 a_33249_48695.t260 VSS 0.065937f
C9205 a_33249_48695.t200 VSS 0.065937f
C9206 a_33249_48695.n143 VSS 0.16732f
C9207 a_33249_48695.t180 VSS 0.065937f
C9208 a_33249_48695.t298 VSS 0.065937f
C9209 a_33249_48695.n144 VSS 0.180576f
C9210 a_33249_48695.n145 VSS 0.4583f
C9211 a_33249_48695.n146 VSS 0.381925f
C9212 a_33249_48695.n147 VSS 0.181417f
C9213 a_33249_48695.t326 VSS 0.173717f
C9214 a_33249_48695.t246 VSS 0.184972f
C9215 a_33249_48695.n148 VSS 0.585662f
C9216 a_33249_48695.n149 VSS 0.451283f
C9217 a_33249_48695.t210 VSS 0.173717f
C9218 a_33249_48695.t309 VSS 0.184972f
C9219 a_33249_48695.n150 VSS 0.583234f
C9220 a_33249_48695.n151 VSS 0.533851f
C9221 a_33249_48695.t314 VSS 0.065937f
C9222 a_33249_48695.t274 VSS 0.065937f
C9223 a_33249_48695.n152 VSS 0.16732f
C9224 a_33249_48695.t238 VSS 0.065937f
C9225 a_33249_48695.t194 VSS 0.065937f
C9226 a_33249_48695.n153 VSS 0.180576f
C9227 a_33249_48695.n154 VSS 0.4583f
C9228 a_33249_48695.n155 VSS 0.357941f
C9229 a_33249_48695.t216 VSS 0.173717f
C9230 a_33249_48695.t312 VSS 0.184972f
C9231 a_33249_48695.n156 VSS 0.59194f
C9232 a_33249_48695.n157 VSS 0.543507f
C9233 a_33249_48695.t196 VSS 0.173717f
C9234 a_33249_48695.t295 VSS 0.184972f
C9235 a_33249_48695.n158 VSS 0.59194f
C9236 a_33249_48695.n159 VSS 0.543525f
C9237 a_33249_48695.t323 VSS 0.065937f
C9238 a_33249_48695.t261 VSS 0.065937f
C9239 a_33249_48695.n160 VSS 0.16732f
C9240 a_33249_48695.t240 VSS 0.065937f
C9241 a_33249_48695.t181 VSS 0.065937f
C9242 a_33249_48695.n161 VSS 0.180576f
C9243 a_33249_48695.n162 VSS 0.4583f
C9244 a_33249_48695.n163 VSS 0.25486f
C9245 a_33249_48695.t237 VSS 0.173717f
C9246 a_33249_48695.t328 VSS 0.184972f
C9247 a_33249_48695.n164 VSS 0.701535f
C9248 a_33249_48695.t330 VSS 0.065937f
C9249 a_33249_48695.t269 VSS 0.065937f
C9250 a_33249_48695.n165 VSS 0.16732f
C9251 a_33249_48695.t252 VSS 0.065937f
C9252 a_33249_48695.t191 VSS 0.065937f
C9253 a_33249_48695.n166 VSS 0.180576f
C9254 a_33249_48695.n167 VSS 0.4583f
C9255 a_33249_48695.n168 VSS 0.484179f
C9256 a_33249_48695.t270 VSS 0.173717f
C9257 a_33249_48695.t192 VSS 0.184972f
C9258 a_33249_48695.n169 VSS 0.583234f
C9259 a_33249_48695.n170 VSS 0.533851f
C9260 a_33249_48695.t204 VSS 0.173717f
C9261 a_33249_48695.t300 VSS 0.184972f
C9262 a_33249_48695.n171 VSS 0.585662f
C9263 a_33249_48695.n172 VSS 0.451283f
C9264 a_33249_48695.n173 VSS 0.181417f
C9265 a_33249_48695.n174 VSS 2.89625f
C9266 a_33249_48695.n175 VSS 2.84854f
C9267 a_33249_48695.n176 VSS 1.25177f
C9268 a_33249_48695.n177 VSS 3.2993f
C9269 a_33249_48695.n178 VSS 2.73275f
C9270 a_33249_48695.n179 VSS 3.19912f
C9271 a_33249_48695.t83 VSS 0.260673f
C9272 a_33249_48695.t24 VSS 0.065937f
C9273 a_33249_48695.t79 VSS 0.065937f
C9274 a_33249_48695.n180 VSS 0.262999f
C9275 a_33249_48695.t80 VSS 0.260673f
C9276 a_33249_48695.t18 VSS 0.065937f
C9277 a_33249_48695.t52 VSS 0.065937f
C9278 a_33249_48695.n181 VSS 0.603414f
C9279 a_33249_48695.t85 VSS 0.260673f
C9280 a_33249_48695.t27 VSS 0.065937f
C9281 a_33249_48695.t62 VSS 0.065937f
C9282 a_33249_48695.n182 VSS 0.603414f
C9283 a_33249_48695.n183 VSS 1.78511f
C9284 a_33249_48695.t91 VSS 0.260673f
C9285 a_33249_48695.t35 VSS 0.065937f
C9286 a_33249_48695.t82 VSS 0.065937f
C9287 a_33249_48695.n184 VSS 0.262999f
C9288 a_33249_48695.n185 VSS 4.43096f
C9289 a_33249_48695.t22 VSS 0.065937f
C9290 a_33249_48695.t45 VSS 0.065937f
C9291 a_33249_48695.n186 VSS 0.197755f
C9292 a_33249_48695.t21 VSS 0.065937f
C9293 a_33249_48695.t43 VSS 0.065937f
C9294 a_33249_48695.n187 VSS 0.153269f
C9295 a_33249_48695.n188 VSS 0.455172f
C9296 a_33249_48695.n189 VSS 0.395085f
C9297 a_33249_48695.t74 VSS 0.065937f
C9298 a_33249_48695.t97 VSS 0.065937f
C9299 a_33249_48695.n190 VSS 0.197755f
C9300 a_33249_48695.t72 VSS 0.065937f
C9301 a_33249_48695.t96 VSS 0.065937f
C9302 a_33249_48695.n191 VSS 0.153269f
C9303 a_33249_48695.n192 VSS 0.455172f
C9304 a_33249_48695.n193 VSS 0.710233f
C9305 a_33249_48695.t66 VSS 0.065937f
C9306 a_33249_48695.t104 VSS 0.065937f
C9307 a_33249_48695.n194 VSS 0.197755f
C9308 a_33249_48695.t64 VSS 0.065937f
C9309 a_33249_48695.t103 VSS 0.065937f
C9310 a_33249_48695.n195 VSS 0.153269f
C9311 a_33249_48695.n196 VSS 0.455172f
C9312 a_33249_48695.n197 VSS 0.710251f
C9313 a_33249_48695.t34 VSS 0.065937f
C9314 a_33249_48695.t61 VSS 0.065937f
C9315 a_33249_48695.n198 VSS 0.197755f
C9316 a_33249_48695.t33 VSS 0.065937f
C9317 a_33249_48695.t59 VSS 0.065937f
C9318 a_33249_48695.n199 VSS 0.153269f
C9319 a_33249_48695.n200 VSS 0.455172f
C9320 a_33249_48695.n201 VSS 0.700454f
C9321 a_33249_48695.t39 VSS 0.065937f
C9322 a_33249_48695.t53 VSS 0.065937f
C9323 a_33249_48695.n202 VSS 0.197755f
C9324 a_33249_48695.t37 VSS 0.065937f
C9325 a_33249_48695.t51 VSS 0.065937f
C9326 a_33249_48695.n203 VSS 0.153269f
C9327 a_33249_48695.n204 VSS 0.63464f
C9328 a_33249_48695.t38 VSS 0.065937f
C9329 a_33249_48695.t93 VSS 0.065937f
C9330 a_33249_48695.n205 VSS 0.197755f
C9331 a_33249_48695.t36 VSS 0.065937f
C9332 a_33249_48695.t92 VSS 0.065937f
C9333 a_33249_48695.n206 VSS 0.153269f
C9334 a_33249_48695.n207 VSS 0.455172f
C9335 a_33249_48695.n208 VSS 0.917033f
C9336 a_33249_48695.t44 VSS 0.065937f
C9337 a_33249_48695.t73 VSS 0.065937f
C9338 a_33249_48695.n209 VSS 0.197755f
C9339 a_33249_48695.t42 VSS 0.065937f
C9340 a_33249_48695.t70 VSS 0.065937f
C9341 a_33249_48695.n210 VSS 0.153269f
C9342 a_33249_48695.n211 VSS 0.455172f
C9343 a_33249_48695.n212 VSS 0.710233f
C9344 a_33249_48695.t77 VSS 0.065937f
C9345 a_33249_48695.t100 VSS 0.065937f
C9346 a_33249_48695.n213 VSS 0.197755f
C9347 a_33249_48695.t76 VSS 0.065937f
C9348 a_33249_48695.t99 VSS 0.065937f
C9349 a_33249_48695.n214 VSS 0.153269f
C9350 a_33249_48695.n215 VSS 0.455172f
C9351 a_33249_48695.n216 VSS 0.188713f
C9352 a_33249_48695.n217 VSS 0.554553f
C9353 a_33249_48695.n218 VSS 3.8908f
C9354 a_33249_48695.t81 VSS 0.065937f
C9355 a_33249_48695.t20 VSS 0.065937f
C9356 a_33249_48695.n219 VSS 0.263576f
C9357 a_33249_48695.n220 VSS 0.96226f
C9358 a_33249_48695.t71 VSS 0.261154f
C9359 a_33249_48695.n221 VSS 1.24524f
C9360 a_33249_48695.t48 VSS 0.506358f
C9361 a_33249_48695.t75 VSS 0.065937f
C9362 a_33249_48695.t101 VSS 0.065937f
C9363 a_33249_48695.n222 VSS 0.263576f
C9364 a_33249_48695.n223 VSS 1.78417f
C9365 a_33249_48695.n224 VSS 1.25132f
C9366 a_33249_48695.n225 VSS 2.79169f
C9367 a_33249_48695.n226 VSS 2.50126f
C9368 a_33249_48695.n227 VSS 1.25252f
C9369 a_33249_48695.n228 VSS 2.77274f
C9370 a_33249_48695.t31 VSS 0.065937f
C9371 a_33249_48695.t49 VSS 0.065937f
C9372 a_33249_48695.n229 VSS 0.197755f
C9373 a_33249_48695.t26 VSS 0.065937f
C9374 a_33249_48695.t47 VSS 0.065937f
C9375 a_33249_48695.n230 VSS 0.153269f
C9376 a_33249_48695.n231 VSS 0.63464f
C9377 a_33249_48695.t30 VSS 0.065937f
C9378 a_33249_48695.t88 VSS 0.065937f
C9379 a_33249_48695.n232 VSS 0.197755f
C9380 a_33249_48695.t25 VSS 0.065937f
C9381 a_33249_48695.t84 VSS 0.065937f
C9382 a_33249_48695.n233 VSS 0.153269f
C9383 a_33249_48695.n234 VSS 0.455172f
C9384 a_33249_48695.n235 VSS 0.917033f
C9385 a_33249_48695.t40 VSS 0.065937f
C9386 a_33249_48695.t65 VSS 0.065937f
C9387 a_33249_48695.n236 VSS 0.197755f
C9388 a_33249_48695.t29 VSS 0.065937f
C9389 a_33249_48695.t56 VSS 0.065937f
C9390 a_33249_48695.n237 VSS 0.153269f
C9391 a_33249_48695.n238 VSS 0.455172f
C9392 a_33249_48695.n239 VSS 0.710233f
C9393 a_33249_48695.t69 VSS 0.065937f
C9394 a_33249_48695.t94 VSS 0.065937f
C9395 a_33249_48695.n240 VSS 0.197755f
C9396 a_33249_48695.t60 VSS 0.065937f
C9397 a_33249_48695.t87 VSS 0.065937f
C9398 a_33249_48695.n241 VSS 0.153269f
C9399 a_33249_48695.n242 VSS 0.455172f
C9400 a_33249_48695.n243 VSS 0.188713f
C9401 a_33249_48695.n244 VSS 0.554553f
C9402 a_33249_48695.t28 VSS 0.065937f
C9403 a_33249_48695.t55 VSS 0.065937f
C9404 a_33249_48695.n245 VSS 0.197755f
C9405 a_33249_48695.t23 VSS 0.065937f
C9406 a_33249_48695.t50 VSS 0.065937f
C9407 a_33249_48695.n246 VSS 0.153269f
C9408 a_33249_48695.n247 VSS 0.455172f
C9409 a_33249_48695.n248 VSS 0.700454f
C9410 a_33249_48695.t58 VSS 0.065937f
C9411 a_33249_48695.t98 VSS 0.065937f
C9412 a_33249_48695.n249 VSS 0.197755f
C9413 a_33249_48695.t54 VSS 0.065937f
C9414 a_33249_48695.t89 VSS 0.065937f
C9415 a_33249_48695.n250 VSS 0.153269f
C9416 a_33249_48695.n251 VSS 0.455172f
C9417 a_33249_48695.n252 VSS 0.710251f
C9418 a_33249_48695.t67 VSS 0.065937f
C9419 a_33249_48695.t90 VSS 0.065937f
C9420 a_33249_48695.n253 VSS 0.197755f
C9421 a_33249_48695.t57 VSS 0.065937f
C9422 a_33249_48695.t86 VSS 0.065937f
C9423 a_33249_48695.n254 VSS 0.153269f
C9424 a_33249_48695.n255 VSS 0.455172f
C9425 a_33249_48695.n256 VSS 0.710233f
C9426 a_33249_48695.t19 VSS 0.065937f
C9427 a_33249_48695.t41 VSS 0.065937f
C9428 a_33249_48695.n257 VSS 0.197755f
C9429 a_33249_48695.t102 VSS 0.065937f
C9430 a_33249_48695.t32 VSS 0.065937f
C9431 a_33249_48695.n258 VSS 0.153269f
C9432 a_33249_48695.n259 VSS 0.455172f
C9433 a_33249_48695.n260 VSS 0.395085f
C9434 a_33249_48695.n261 VSS 2.54509f
C9435 a_33249_48695.n262 VSS 3.86208f
C9436 a_33249_48695.t78 VSS 0.065937f
C9437 a_33249_48695.t105 VSS 0.065937f
C9438 a_33249_48695.n263 VSS 0.263576f
C9439 a_33249_48695.n264 VSS 0.96226f
C9440 a_33249_48695.t63 VSS 0.261154f
C9441 a_33249_48695.n265 VSS 1.24524f
C9442 a_33249_48695.t46 VSS 0.506358f
C9443 a_33249_48695.t68 VSS 0.065937f
C9444 a_33249_48695.t95 VSS 0.065937f
C9445 a_33249_48695.n266 VSS 0.263576f
C9446 a_33249_48695.n267 VSS 1.78417f
C9447 a_33249_48695.n268 VSS 1.25132f
C9448 a_33249_48695.n269 VSS 3.1335f
C9449 a_33249_48695.n270 VSS 2.00968f
C9450 a_33249_48695.n271 VSS 2.08409f
C9451 a_33249_48695.n272 VSS 2.79169f
C9452 a_33249_48695.t337 VSS 0.065937f
C9453 a_33249_48695.t107 VSS 0.065937f
C9454 a_33249_48695.n273 VSS 0.361324f
C9455 a_33249_48695.t13 VSS 0.065937f
C9456 a_33249_48695.t148 VSS 0.065937f
C9457 a_33249_48695.n274 VSS 0.241202f
C9458 a_33249_48695.t9 VSS 0.065937f
C9459 a_33249_48695.t152 VSS 0.065937f
C9460 a_33249_48695.n275 VSS 0.241202f
C9461 a_33249_48695.t113 VSS 0.065937f
C9462 a_33249_48695.t5 VSS 0.065937f
C9463 a_33249_48695.n276 VSS 0.241202f
C9464 a_33249_48695.t124 VSS 0.065937f
C9465 a_33249_48695.t149 VSS 0.065937f
C9466 a_33249_48695.n277 VSS 0.241202f
C9467 a_33249_48695.t106 VSS 0.065937f
C9468 a_33249_48695.t12 VSS 0.065937f
C9469 a_33249_48695.n278 VSS 0.241202f
C9470 a_33249_48695.t118 VSS 0.065937f
C9471 a_33249_48695.t146 VSS 0.065937f
C9472 a_33249_48695.n279 VSS 0.241202f
C9473 a_33249_48695.t119 VSS 0.065937f
C9474 a_33249_48695.t346 VSS 0.065937f
C9475 a_33249_48695.n280 VSS 0.241202f
C9476 a_33249_48695.t140 VSS 0.065937f
C9477 a_33249_48695.t0 VSS 0.065937f
C9478 a_33249_48695.n281 VSS 0.181906f
C9479 a_33249_48695.t139 VSS 0.065937f
C9480 a_33249_48695.t334 VSS 0.065937f
C9481 a_33249_48695.n282 VSS 0.166113f
C9482 a_33249_48695.n283 VSS 1.02196f
C9483 a_33249_48695.t130 VSS 0.186098f
C9484 a_33249_48695.t128 VSS 0.172688f
C9485 a_33249_48695.n284 VSS 0.59185f
C9486 a_33249_48695.n285 VSS 1.17271f
C9487 a_33249_48695.t122 VSS 0.065937f
C9488 a_33249_48695.t343 VSS 0.065937f
C9489 a_33249_48695.n286 VSS 0.361324f
C9490 a_33249_48695.t132 VSS 0.065937f
C9491 a_33249_48695.t156 VSS 0.065937f
C9492 a_33249_48695.n287 VSS 0.241202f
C9493 a_33249_48695.t126 VSS 0.065937f
C9494 a_33249_48695.t338 VSS 0.065937f
C9495 a_33249_48695.n288 VSS 0.241202f
C9496 a_33249_48695.t108 VSS 0.065937f
C9497 a_33249_48695.t123 VSS 0.065937f
C9498 a_33249_48695.n289 VSS 0.241202f
C9499 a_33249_48695.t135 VSS 0.065937f
C9500 a_33249_48695.t340 VSS 0.065937f
C9501 a_33249_48695.n290 VSS 0.241202f
C9502 a_33249_48695.t341 VSS 0.065937f
C9503 a_33249_48695.t129 VSS 0.065937f
C9504 a_33249_48695.n291 VSS 0.241202f
C9505 a_33249_48695.t109 VSS 0.065937f
C9506 a_33249_48695.t153 VSS 0.065937f
C9507 a_33249_48695.n292 VSS 0.241202f
C9508 a_33249_48695.t15 VSS 0.065937f
C9509 a_33249_48695.t6 VSS 0.065937f
C9510 a_33249_48695.n293 VSS 0.241202f
C9511 a_33249_48695.n294 VSS 1.13487f
C9512 a_33249_48695.n295 VSS 3.83834f
C9513 a_33249_48695.n296 VSS 1.25143f
C9514 a_33249_48695.t134 VSS 0.065937f
C9515 a_33249_48695.t336 VSS 0.065937f
C9516 a_33249_48695.n297 VSS 0.181906f
C9517 a_33249_48695.t133 VSS 0.065937f
C9518 a_33249_48695.t335 VSS 0.065937f
C9519 a_33249_48695.n298 VSS 0.166113f
C9520 a_33249_48695.n299 VSS 0.458182f
C9521 a_33249_48695.n300 VSS 1.08733f
C9522 a_33249_48695.t350 VSS 0.186098f
C9523 a_33249_48695.t349 VSS 0.172688f
C9524 a_33249_48695.n301 VSS 0.59185f
C9525 a_33249_48695.n302 VSS 0.708323f
C9526 a_33249_48695.n303 VSS 4.22418f
C9527 a_33249_48695.t154 VSS 0.065937f
C9528 a_33249_48695.t117 VSS 0.065937f
C9529 a_33249_48695.n304 VSS 0.362253f
C9530 a_33249_48695.t8 VSS 0.065937f
C9531 a_33249_48695.t143 VSS 0.065937f
C9532 a_33249_48695.n305 VSS 0.241904f
C9533 a_33249_48695.n306 VSS 1.18974f
C9534 a_33249_48695.t2 VSS 0.065937f
C9535 a_33249_48695.t147 VSS 0.065937f
C9536 a_33249_48695.n307 VSS 0.241904f
C9537 a_33249_48695.n308 VSS 0.843784f
C9538 a_33249_48695.t333 VSS 0.065937f
C9539 a_33249_48695.t348 VSS 0.065937f
C9540 a_33249_48695.n309 VSS 0.241904f
C9541 a_33249_48695.n310 VSS 0.338896f
C9542 a_33249_48695.n311 VSS 0.549879f
C9543 a_33249_48695.t10 VSS 0.065937f
C9544 a_33249_48695.t145 VSS 0.065937f
C9545 a_33249_48695.n312 VSS 0.241904f
C9546 a_33249_48695.n313 VSS 0.822009f
C9547 a_33249_48695.t114 VSS 0.065937f
C9548 a_33249_48695.t7 VSS 0.065937f
C9549 a_33249_48695.n314 VSS 0.241904f
C9550 a_33249_48695.n315 VSS 0.843766f
C9551 a_33249_48695.t1 VSS 0.065937f
C9552 a_33249_48695.t141 VSS 0.065937f
C9553 a_33249_48695.n316 VSS 0.241904f
C9554 a_33249_48695.n317 VSS 0.843784f
C9555 a_33249_48695.t120 VSS 0.065937f
C9556 a_33249_48695.t342 VSS 0.065937f
C9557 a_33249_48695.n318 VSS 0.241904f
C9558 a_33249_48695.n319 VSS 0.518838f
C9559 a_33249_48695.n320 VSS 2.81996f
C9560 a_33249_48695.n321 VSS 2.71764f
C9561 a_33249_48695.n322 VSS 0.549826f
C9562 a_33249_48695.n323 VSS 2.6883f
C9563 a_33249_48695.t136 VSS 0.065937f
C9564 a_33249_48695.t116 VSS 0.065937f
C9565 a_33249_48695.n324 VSS 0.181906f
C9566 a_33249_48695.t131 VSS 0.065937f
C9567 a_33249_48695.t339 VSS 0.065937f
C9568 a_33249_48695.n325 VSS 0.166113f
C9569 a_33249_48695.n326 VSS 1.02196f
C9570 a_33249_48695.t125 VSS 0.186098f
C9571 a_33249_48695.t11 VSS 0.172688f
C9572 a_33249_48695.n327 VSS 0.59185f
C9573 a_33249_48695.n328 VSS 1.17271f
C9574 a_33249_48695.t345 VSS 0.186098f
C9575 a_33249_48695.t17 VSS 0.172688f
C9576 a_33249_48695.n329 VSS 0.59185f
C9577 a_33249_48695.n330 VSS 0.708323f
C9578 a_33249_48695.t127 VSS 0.065937f
C9579 a_33249_48695.t155 VSS 0.065937f
C9580 a_33249_48695.n331 VSS 0.181906f
C9581 a_33249_48695.t14 VSS 0.065937f
C9582 a_33249_48695.t150 VSS 0.065937f
C9583 a_33249_48695.n332 VSS 0.166113f
C9584 a_33249_48695.n333 VSS 0.458182f
C9585 a_33249_48695.n334 VSS 1.08733f
C9586 a_33249_48695.n335 VSS 1.25143f
C9587 a_33249_48695.n336 VSS 2.33745f
C9588 a_33249_48695.n337 VSS 3.07641f
C9589 a_33249_48695.n338 VSS 0.549879f
C9590 a_33249_48695.t4 VSS 0.065937f
C9591 a_33249_48695.t142 VSS 0.065937f
C9592 a_33249_48695.n339 VSS 0.241904f
C9593 a_33249_48695.n340 VSS 0.822009f
C9594 a_33249_48695.t121 VSS 0.065937f
C9595 a_33249_48695.t351 VSS 0.065937f
C9596 a_33249_48695.n341 VSS 0.241904f
C9597 a_33249_48695.n342 VSS 0.843766f
C9598 a_33249_48695.t110 VSS 0.065937f
C9599 a_33249_48695.t137 VSS 0.065937f
C9600 a_33249_48695.n343 VSS 0.241904f
C9601 a_33249_48695.n344 VSS 0.843784f
C9602 a_33249_48695.t111 VSS 0.065937f
C9603 a_33249_48695.t16 VSS 0.065937f
C9604 a_33249_48695.n345 VSS 0.241904f
C9605 a_33249_48695.n346 VSS 0.518838f
C9606 a_33249_48695.n347 VSS 3.43055f
C9607 a_33249_48695.n348 VSS 2.84218f
C9608 a_33249_48695.n349 VSS 3.04283f
C9609 a_33249_48695.n350 VSS 0.1838f
C9610 a_33249_48695.n351 VSS 0.1838f
C9611 a_33249_48695.n352 VSS 3.0578f
C9612 a_33249_48695.t171 VSS 0.162517f
C9613 a_33249_48695.t263 VSS 0.198291f
C9614 a_33249_48695.n353 VSS 1.06267f
C9615 a_33249_48695.t288 VSS 0.065937f
C9616 a_33249_48695.t190 VSS 0.065937f
C9617 a_33249_48695.n354 VSS 0.154318f
C9618 a_33249_48695.t208 VSS 0.065937f
C9619 a_33249_48695.t285 VSS 0.065937f
C9620 a_33249_48695.n355 VSS 0.196324f
C9621 a_33249_48695.n356 VSS 0.446847f
C9622 a_33249_48695.n357 VSS 0.976786f
C9623 a_33249_48695.t305 VSS 0.065937f
C9624 a_33249_48695.t230 VSS 0.065937f
C9625 a_33249_48695.n358 VSS 0.154318f
C9626 a_33249_48695.t223 VSS 0.065937f
C9627 a_33249_48695.t327 VSS 0.065937f
C9628 a_33249_48695.n359 VSS 0.196324f
C9629 a_33249_48695.n360 VSS 0.446847f
C9630 a_33249_48695.n361 VSS 0.776654f
C9631 a_33249_48695.t185 VSS 0.162517f
C9632 a_33249_48695.t280 VSS 0.198291f
C9633 a_33249_48695.n362 VSS 0.581116f
C9634 a_33249_48695.n363 VSS 1.18777f
C9635 a_33249_48695.n364 VSS 1.2517f
C9636 a_33249_48695.n365 VSS 2.70921f
C9637 a_33249_48695.n366 VSS 2.41819f
C9638 a_33249_48695.n367 VSS 0.183807f
C9639 a_33249_48695.t329 VSS 0.065937f
C9640 a_33249_48695.t291 VSS 0.065937f
C9641 a_33249_48695.n368 VSS 0.285449f
C9642 a_33249_48695.n369 VSS 0.428366f
C9643 a_33249_48695.t235 VSS 0.279755f
C9644 a_33249_48695.n370 VSS 0.806849f
C9645 a_33249_48695.t212 VSS 0.277438f
C9646 a_33249_48695.n371 VSS 0.80029f
C9647 a_33249_48695.t162 VSS 0.065937f
C9648 a_33249_48695.t277 VSS 0.065937f
C9649 a_33249_48695.n372 VSS 0.285449f
C9650 a_33249_48695.n373 VSS 0.542569f
C9651 a_33249_48695.t222 VSS 0.279833f
C9652 a_33249_48695.n374 VSS 0.795271f
C9653 a_33249_48695.t287 VSS 0.277438f
C9654 a_33249_48695.n375 VSS 0.720574f
C9655 a_33249_48695.t251 VSS 0.374369f
C9656 a_33249_48695.t169 VSS 0.065937f
C9657 a_33249_48695.t286 VSS 0.065937f
C9658 a_33249_48695.n376 VSS 0.285449f
C9659 a_33249_48695.n377 VSS 0.837958f
C9660 a_33249_48695.n378 VSS 0.183807f
C9661 a_33249_48695.n379 VSS 2.41819f
C9662 a_33249_48695.t255 VSS 0.372643f
C9663 a_33249_48695.t215 VSS 0.065937f
C9664 a_33249_48695.t159 VSS 0.065937f
C9665 a_33249_48695.n380 VSS 0.284868f
C9666 a_33249_48695.t279 VSS 0.279265f
C9667 a_33249_48695.t168 VSS 0.278903f
C9668 a_33249_48695.n381 VSS 0.1838f
C9669 a_33249_48695.t266 VSS 0.065937f
C9670 a_33249_48695.t233 VSS 0.065937f
C9671 a_33249_48695.n382 VSS 0.284868f
C9672 a_33249_48695.t173 VSS 0.279265f
C9673 a_33249_48695.t331 VSS 0.279265f
C9674 a_33249_48695.t276 VSS 0.065937f
C9675 a_33249_48695.t218 VSS 0.065937f
C9676 a_33249_48695.n383 VSS 0.284868f
C9677 a_33249_48695.t160 VSS 0.279265f
C9678 a_33249_48695.t228 VSS 0.278903f
C9679 a_33249_48695.t284 VSS 0.065937f
C9680 a_33249_48695.t226 VSS 0.065937f
C9681 a_33249_48695.n384 VSS 0.284868f
C9682 a_33249_48695.t188 VSS 0.373143f
C9683 a_33249_48695.n385 VSS 0.1838f
C9684 a_33249_48695.n386 VSS 2.69004f
C9685 a_33249_48695.n387 VSS 4.1989f
C9686 a_33249_48695.t232 VSS 0.065937f
C9687 a_33249_48695.t157 VSS 0.065937f
C9688 a_33249_48695.n388 VSS 0.154318f
C9689 a_33249_48695.t273 VSS 0.065937f
C9690 a_33249_48695.t198 VSS 0.065937f
C9691 a_33249_48695.n389 VSS 0.196324f
C9692 a_33249_48695.n390 VSS 0.446847f
C9693 a_33249_48695.n391 VSS 0.776654f
C9694 a_33249_48695.t290 VSS 0.162517f
C9695 a_33249_48695.t158 VSS 0.198291f
C9696 a_33249_48695.n392 VSS 0.581116f
C9697 a_33249_48695.n393 VSS 1.18777f
C9698 a_33249_48695.n394 VSS 1.2517f
C9699 a_33249_48695.n395 VSS 3.7876f
C9700 a_33249_48695.n396 VSS 0.642382f
C9701 a_33249_48695.n397 VSS 0.720563f
C9702 a_33249_48695.t332 VSS 0.277438f
C9703 a_106809_n17715.t1 VSS 0.995519f
C9704 a_106809_n17715.t0 VSS 1.00448f
C9705 a_71342_n30339.n0 VSS 10.6245f
C9706 a_71342_n30339.t2 VSS 0.843931f
C9707 a_71342_n30339.t3 VSS 0.685986f
C9708 a_71342_n30339.t1 VSS 0.632984f
C9709 a_71342_n30339.t0 VSS 0.812605f
C9710 a_65486_n36322.n0 VSS 11.550099f
C9711 a_65486_n36322.n1 VSS 0.727597f
C9712 a_65486_n36322.n2 VSS 11.477901f
C9713 a_65486_n36322.t14 VSS 0.458717f
C9714 a_65486_n36322.t20 VSS 0.45876f
C9715 a_65486_n36322.t2 VSS 0.278471f
C9716 a_65486_n36322.t23 VSS 0.452124f
C9717 a_65486_n36322.t8 VSS 0.452124f
C9718 a_65486_n36322.t19 VSS 0.450255f
C9719 a_65486_n36322.t11 VSS 0.450255f
C9720 a_65486_n36322.t22 VSS 0.45876f
C9721 a_65486_n36322.t9 VSS 0.450255f
C9722 a_65486_n36322.t16 VSS 0.450255f
C9723 a_65486_n36322.t17 VSS 0.452124f
C9724 a_65486_n36322.t10 VSS 0.450255f
C9725 a_65486_n36322.t15 VSS 0.452124f
C9726 a_65486_n36322.t18 VSS 0.450255f
C9727 a_65486_n36322.t13 VSS 0.458717f
C9728 a_65486_n36322.t21 VSS 0.450255f
C9729 a_65486_n36322.t12 VSS 0.450255f
C9730 a_65486_n36322.t5 VSS 0.410822f
C9731 a_65486_n36322.t6 VSS 0.242341f
C9732 a_65486_n36322.t7 VSS 0.273797f
C9733 a_65486_n36322.t4 VSS 0.423358f
C9734 a_65486_n36322.t1 VSS 0.39953f
C9735 a_65486_n36322.t3 VSS 0.50972f
C9736 a_65486_n36322.t0 VSS 0.260911f
C9737 a_50751_n19729.n0 VSS 0.022671f
C9738 a_50751_n19729.n1 VSS 0.027893f
C9739 a_50751_n19729.n2 VSS 0.037978f
C9740 a_50751_n19729.n3 VSS 0.022671f
C9741 a_50751_n19729.n4 VSS 0.027893f
C9742 a_50751_n19729.n5 VSS 0.022671f
C9743 a_50751_n19729.n6 VSS 0.249456f
C9744 a_50751_n19729.n7 VSS 0.027893f
C9745 a_50751_n19729.n8 VSS 0.022671f
C9746 a_50751_n19729.n9 VSS 0.027893f
C9747 a_50751_n19729.n10 VSS 0.022671f
C9748 a_50751_n19729.n11 VSS 0.027893f
C9749 a_50751_n19729.n12 VSS 0.02267f
C9750 a_50751_n19729.n13 VSS 0.027893f
C9751 a_50751_n19729.n14 VSS 0.022671f
C9752 a_50751_n19729.n15 VSS 0.027893f
C9753 a_50751_n19729.n16 VSS 0.022671f
C9754 a_50751_n19729.n17 VSS 0.027893f
C9755 a_50751_n19729.n18 VSS 0.022671f
C9756 a_50751_n19729.n19 VSS 0.110201f
C9757 a_50751_n19729.n20 VSS 0.027893f
C9758 a_50751_n19729.n21 VSS 0.022671f
C9759 a_50751_n19729.n22 VSS 0.154502f
C9760 a_50751_n19729.n23 VSS 0.027893f
C9761 a_50751_n19729.n24 VSS 0.022671f
C9762 a_50751_n19729.n25 VSS 0.027893f
C9763 a_50751_n19729.n26 VSS 0.022671f
C9764 a_50751_n19729.n27 VSS 0.173273f
C9765 a_50751_n19729.n28 VSS 0.027893f
C9766 a_50751_n19729.n29 VSS 0.02267f
C9767 a_50751_n19729.n30 VSS 0.027893f
C9768 a_50751_n19729.n31 VSS 0.022671f
C9769 a_50751_n19729.n32 VSS 0.027893f
C9770 a_50751_n19729.n33 VSS 0.022671f
C9771 a_50751_n19729.n34 VSS 0.027893f
C9772 a_50751_n19729.n35 VSS 0.022671f
C9773 a_50751_n19729.n36 VSS 0.055116f
C9774 a_50751_n19729.n37 VSS 0.027893f
C9775 a_50751_n19729.n38 VSS 0.022671f
C9776 a_50751_n19729.n39 VSS 0.027893f
C9777 a_50751_n19729.n40 VSS 0.02267f
C9778 a_50751_n19729.n41 VSS 0.027893f
C9779 a_50751_n19729.n42 VSS 0.022671f
C9780 a_50751_n19729.n43 VSS 0.027893f
C9781 a_50751_n19729.n44 VSS 0.022671f
C9782 a_50751_n19729.n45 VSS 0.027893f
C9783 a_50751_n19729.n46 VSS 0.022671f
C9784 a_50751_n19729.n47 VSS 0.110201f
C9785 a_50751_n19729.n48 VSS 0.027893f
C9786 a_50751_n19729.n49 VSS 0.022671f
C9787 a_50751_n19729.n50 VSS 0.200348f
C9788 a_50751_n19729.n51 VSS 0.027893f
C9789 a_50751_n19729.n52 VSS 0.022671f
C9790 a_50751_n19729.n53 VSS 0.027893f
C9791 a_50751_n19729.n54 VSS 0.02267f
C9792 a_50751_n19729.n55 VSS 0.027893f
C9793 a_50751_n19729.n56 VSS 0.022671f
C9794 a_50751_n19729.n57 VSS 0.027893f
C9795 a_50751_n19729.n58 VSS 0.022671f
C9796 a_50751_n19729.n59 VSS 0.027893f
C9797 a_50751_n19729.n60 VSS 0.022671f
C9798 a_50751_n19729.n61 VSS 0.027893f
C9799 a_50751_n19729.n62 VSS 0.022671f
C9800 a_50751_n19729.n63 VSS 0.027893f
C9801 a_50751_n19729.n64 VSS 0.037978f
C9802 a_50751_n19729.n65 VSS 0.022671f
C9803 a_50751_n19729.n66 VSS 0.027893f
C9804 a_50751_n19729.n67 VSS 0.022671f
C9805 a_50751_n19729.n68 VSS 0.249456f
C9806 a_50751_n19729.n69 VSS 0.027893f
C9807 a_50751_n19729.n70 VSS 0.022671f
C9808 a_50751_n19729.n71 VSS 0.027893f
C9809 a_50751_n19729.n72 VSS 0.022671f
C9810 a_50751_n19729.n73 VSS 0.027893f
C9811 a_50751_n19729.n74 VSS 0.02267f
C9812 a_50751_n19729.n75 VSS 0.110201f
C9813 a_50751_n19729.n76 VSS 0.027893f
C9814 a_50751_n19729.n77 VSS 0.022671f
C9815 a_50751_n19729.n78 VSS 0.027893f
C9816 a_50751_n19729.n79 VSS 0.022671f
C9817 a_50751_n19729.n80 VSS 0.055085f
C9818 a_50751_n19729.n81 VSS 0.027893f
C9819 a_50751_n19729.n82 VSS 0.022671f
C9820 a_50751_n19729.n83 VSS 0.027893f
C9821 a_50751_n19729.n84 VSS 0.022671f
C9822 a_50751_n19729.n85 VSS 0.027893f
C9823 a_50751_n19729.n86 VSS 0.022671f
C9824 a_50751_n19729.n87 VSS 0.154502f
C9825 a_50751_n19729.n88 VSS 0.027893f
C9826 a_50751_n19729.n89 VSS 0.022671f
C9827 a_50751_n19729.n90 VSS 0.173273f
C9828 a_50751_n19729.n91 VSS 0.027893f
C9829 a_50751_n19729.n92 VSS 0.02267f
C9830 a_50751_n19729.n93 VSS 0.027893f
C9831 a_50751_n19729.n94 VSS 0.022671f
C9832 a_50751_n19729.n95 VSS 0.027893f
C9833 a_50751_n19729.n96 VSS 0.022671f
C9834 a_50751_n19729.n97 VSS 0.027893f
C9835 a_50751_n19729.n98 VSS 0.022671f
C9836 a_50751_n19729.n99 VSS 0.055116f
C9837 a_50751_n19729.n100 VSS 0.027893f
C9838 a_50751_n19729.n101 VSS 0.022671f
C9839 a_50751_n19729.n102 VSS 0.027893f
C9840 a_50751_n19729.n103 VSS 0.02267f
C9841 a_50751_n19729.n104 VSS 0.027893f
C9842 a_50751_n19729.n105 VSS 0.022671f
C9843 a_50751_n19729.n106 VSS 0.027893f
C9844 a_50751_n19729.n107 VSS 0.022671f
C9845 a_50751_n19729.n108 VSS 0.027893f
C9846 a_50751_n19729.n109 VSS 0.022671f
C9847 a_50751_n19729.n110 VSS 0.110201f
C9848 a_50751_n19729.n111 VSS 0.027893f
C9849 a_50751_n19729.n112 VSS 0.022671f
C9850 a_50751_n19729.n113 VSS 0.200348f
C9851 a_50751_n19729.n114 VSS 0.027893f
C9852 a_50751_n19729.n115 VSS 0.022671f
C9853 a_50751_n19729.n116 VSS 0.027893f
C9854 a_50751_n19729.n117 VSS 0.02267f
C9855 a_50751_n19729.n118 VSS 0.027893f
C9856 a_50751_n19729.n119 VSS 0.022671f
C9857 a_50751_n19729.n120 VSS 0.027893f
C9858 a_50751_n19729.n121 VSS 0.022671f
C9859 a_50751_n19729.n122 VSS 0.027893f
C9860 a_50751_n19729.n123 VSS 0.022671f
C9861 a_50751_n19729.n124 VSS 0.027893f
C9862 a_50751_n19729.n125 VSS 0.02267f
C9863 a_50751_n19729.n126 VSS 0.027893f
C9864 a_50751_n19729.n127 VSS 0.022671f
C9865 a_50751_n19729.n128 VSS 0.027893f
C9866 a_50751_n19729.n129 VSS 0.022671f
C9867 a_50751_n19729.n130 VSS 0.027893f
C9868 a_50751_n19729.n131 VSS 0.022671f
C9869 a_50751_n19729.n132 VSS 0.027893f
C9870 a_50751_n19729.n133 VSS 0.022671f
C9871 a_50751_n19729.n134 VSS 0.027893f
C9872 a_50751_n19729.n135 VSS 0.037978f
C9873 a_50751_n19729.n136 VSS 0.022671f
C9874 a_50751_n19729.n137 VSS 0.027893f
C9875 a_50751_n19729.n138 VSS 0.022671f
C9876 a_50751_n19729.n139 VSS 0.249456f
C9877 a_50751_n19729.n140 VSS 0.027893f
C9878 a_50751_n19729.n141 VSS 0.022671f
C9879 a_50751_n19729.n142 VSS 0.027893f
C9880 a_50751_n19729.n143 VSS 0.022671f
C9881 a_50751_n19729.n144 VSS 0.027893f
C9882 a_50751_n19729.n145 VSS 0.02267f
C9883 a_50751_n19729.n146 VSS 0.110201f
C9884 a_50751_n19729.n147 VSS 0.027893f
C9885 a_50751_n19729.n148 VSS 0.022671f
C9886 a_50751_n19729.n149 VSS 0.027893f
C9887 a_50751_n19729.n150 VSS 0.022671f
C9888 a_50751_n19729.n151 VSS 0.055085f
C9889 a_50751_n19729.n152 VSS 0.027893f
C9890 a_50751_n19729.n153 VSS 0.022671f
C9891 a_50751_n19729.n154 VSS 0.027893f
C9892 a_50751_n19729.n155 VSS 0.022671f
C9893 a_50751_n19729.n156 VSS 0.027893f
C9894 a_50751_n19729.n157 VSS 0.022671f
C9895 a_50751_n19729.n158 VSS 0.154502f
C9896 a_50751_n19729.n159 VSS 0.027893f
C9897 a_50751_n19729.n160 VSS 0.022671f
C9898 a_50751_n19729.n161 VSS 0.173273f
C9899 a_50751_n19729.n162 VSS 0.027893f
C9900 a_50751_n19729.n163 VSS 0.02267f
C9901 a_50751_n19729.n164 VSS 0.027893f
C9902 a_50751_n19729.n165 VSS 0.022671f
C9903 a_50751_n19729.n166 VSS 0.027893f
C9904 a_50751_n19729.n167 VSS 0.022671f
C9905 a_50751_n19729.n168 VSS 0.027893f
C9906 a_50751_n19729.n169 VSS 0.022671f
C9907 a_50751_n19729.n170 VSS 0.055116f
C9908 a_50751_n19729.n171 VSS 0.027893f
C9909 a_50751_n19729.n172 VSS 0.022671f
C9910 a_50751_n19729.n173 VSS 0.027893f
C9911 a_50751_n19729.n174 VSS 0.02267f
C9912 a_50751_n19729.n175 VSS 0.027893f
C9913 a_50751_n19729.n176 VSS 0.022671f
C9914 a_50751_n19729.n177 VSS 0.027893f
C9915 a_50751_n19729.n178 VSS 0.022671f
C9916 a_50751_n19729.n179 VSS 0.027893f
C9917 a_50751_n19729.n180 VSS 0.022671f
C9918 a_50751_n19729.n181 VSS 0.110201f
C9919 a_50751_n19729.n182 VSS 0.027893f
C9920 a_50751_n19729.n183 VSS 0.022671f
C9921 a_50751_n19729.n184 VSS 0.200348f
C9922 a_50751_n19729.n185 VSS 0.027893f
C9923 a_50751_n19729.n186 VSS 0.022671f
C9924 a_50751_n19729.n187 VSS 0.027893f
C9925 a_50751_n19729.n188 VSS 0.02267f
C9926 a_50751_n19729.n189 VSS 0.027893f
C9927 a_50751_n19729.n190 VSS 0.022671f
C9928 a_50751_n19729.n191 VSS 0.027893f
C9929 a_50751_n19729.n192 VSS 0.022671f
C9930 a_50751_n19729.n193 VSS 0.027893f
C9931 a_50751_n19729.n194 VSS 0.022671f
C9932 a_50751_n19729.n195 VSS 0.027893f
C9933 a_50751_n19729.n196 VSS 0.02267f
C9934 a_50751_n19729.n197 VSS 0.027893f
C9935 a_50751_n19729.n198 VSS 0.022671f
C9936 a_50751_n19729.n199 VSS 0.027893f
C9937 a_50751_n19729.n200 VSS 0.022671f
C9938 a_50751_n19729.n201 VSS 0.027893f
C9939 a_50751_n19729.n202 VSS 0.022671f
C9940 a_50751_n19729.n203 VSS 0.027893f
C9941 a_50751_n19729.n204 VSS 0.02267f
C9942 a_50751_n19729.n205 VSS 0.027893f
C9943 a_50751_n19729.n206 VSS 0.022671f
C9944 a_50751_n19729.n207 VSS 0.027893f
C9945 a_50751_n19729.n208 VSS 0.022671f
C9946 a_50751_n19729.n209 VSS 0.027893f
C9947 a_50751_n19729.n210 VSS 0.022671f
C9948 a_50751_n19729.n211 VSS 0.027893f
C9949 a_50751_n19729.n212 VSS 0.023132f
C9950 a_50751_n19729.n213 VSS 0.028615f
C9951 a_50751_n19729.n214 VSS 0.023132f
C9952 a_50751_n19729.n215 VSS 0.032477f
C9953 a_50751_n19729.n216 VSS 0.023132f
C9954 a_50751_n19729.n217 VSS 0.028615f
C9955 a_50751_n19729.n218 VSS 0.023132f
C9956 a_50751_n19729.n219 VSS 0.032477f
C9957 a_50751_n19729.n220 VSS 0.023132f
C9958 a_50751_n19729.n221 VSS 0.028615f
C9959 a_50751_n19729.n222 VSS 0.023132f
C9960 a_50751_n19729.n223 VSS 0.032477f
C9961 a_50751_n19729.n224 VSS 0.055085f
C9962 a_50751_n19729.n225 VSS 0.024116f
C9963 a_50751_n19729.t41 VSS 0.007577f
C9964 a_50751_n19729.n226 VSS 0.021816f
C9965 a_50751_n19729.t31 VSS 0.007577f
C9966 a_50751_n19729.n227 VSS 0.016705f
C9967 a_50751_n19729.t9 VSS 0.007577f
C9968 a_50751_n19729.n228 VSS 0.021871f
C9969 a_50751_n19729.t358 VSS 0.039522f
C9970 a_50751_n19729.t237 VSS 0.039472f
C9971 a_50751_n19729.n229 VSS 0.02267f
C9972 a_50751_n19729.n230 VSS 0.045097f
C9973 a_50751_n19729.t229 VSS 0.042148f
C9974 a_50751_n19729.n231 VSS 0.045377f
C9975 a_50751_n19729.n232 VSS 0.045401f
C9976 a_50751_n19729.t357 VSS 0.042151f
C9977 a_50751_n19729.t152 VSS 0.039522f
C9978 a_50751_n19729.n233 VSS 0.045401f
C9979 a_50751_n19729.t227 VSS 0.039522f
C9980 a_50751_n19729.n234 VSS 0.045401f
C9981 a_50751_n19729.t137 VSS 0.042151f
C9982 a_50751_n19729.t224 VSS 0.039522f
C9983 a_50751_n19729.n235 VSS 0.045401f
C9984 a_50751_n19729.t138 VSS 0.039522f
C9985 a_50751_n19729.t315 VSS 0.039522f
C9986 a_50751_n19729.n236 VSS 0.045377f
C9987 a_50751_n19729.t308 VSS 0.042148f
C9988 a_50751_n19729.n237 VSS 0.045377f
C9989 a_50751_n19729.t307 VSS 0.039522f
C9990 a_50751_n19729.n238 VSS 0.045401f
C9991 a_50751_n19729.t122 VSS 0.042151f
C9992 a_50751_n19729.t216 VSS 0.039522f
C9993 a_50751_n19729.n239 VSS 0.045401f
C9994 a_50751_n19729.t123 VSS 0.039522f
C9995 a_50751_n19729.t303 VSS 0.039522f
C9996 a_50751_n19729.n240 VSS 0.045377f
C9997 a_50751_n19729.t296 VSS 0.042148f
C9998 a_50751_n19729.n241 VSS 0.045377f
C9999 a_50751_n19729.t294 VSS 0.039522f
C10000 a_50751_n19729.n242 VSS 0.045401f
C10001 a_50751_n19729.t194 VSS 0.042151f
C10002 a_50751_n19729.t290 VSS 0.039522f
C10003 a_50751_n19729.n243 VSS 0.045401f
C10004 a_50751_n19729.t40 VSS 0.039522f
C10005 a_50751_n19729.t88 VSS 0.039477f
C10006 a_50751_n19729.n244 VSS 0.045123f
C10007 a_50751_n19729.t81 VSS 0.042148f
C10008 a_50751_n19729.n245 VSS 0.045377f
C10009 a_50751_n19729.t70 VSS 0.039522f
C10010 a_50751_n19729.n246 VSS 0.045401f
C10011 a_50751_n19729.t274 VSS 0.042151f
C10012 a_50751_n19729.t76 VSS 0.039522f
C10013 a_50751_n19729.n247 VSS 0.045401f
C10014 a_50751_n19729.t30 VSS 0.039522f
C10015 a_50751_n19729.t155 VSS 0.039475f
C10016 a_50751_n19729.n248 VSS 0.045377f
C10017 a_50751_n19729.t149 VSS 0.042148f
C10018 a_50751_n19729.n249 VSS 0.04511f
C10019 a_50751_n19729.t48 VSS 0.039522f
C10020 a_50751_n19729.n250 VSS 0.045401f
C10021 a_50751_n19729.t346 VSS 0.042151f
C10022 a_50751_n19729.t145 VSS 0.039522f
C10023 a_50751_n19729.n251 VSS 0.045401f
C10024 a_50751_n19729.t8 VSS 0.039522f
C10025 a_50751_n19729.t228 VSS 0.039522f
C10026 a_50751_n19729.n252 VSS 0.045377f
C10027 a_50751_n19729.t222 VSS 0.042148f
C10028 a_50751_n19729.n253 VSS 0.045377f
C10029 a_50751_n19729.t36 VSS 0.039522f
C10030 a_50751_n19729.t57 VSS 0.007577f
C10031 a_50751_n19729.n254 VSS 0.021816f
C10032 a_50751_n19729.t65 VSS 0.007577f
C10033 a_50751_n19729.n255 VSS 0.016705f
C10034 a_50751_n19729.t47 VSS 0.007577f
C10035 a_50751_n19729.n256 VSS 0.021871f
C10036 a_50751_n19729.n257 VSS 0.045401f
C10037 a_50751_n19729.t250 VSS 0.042151f
C10038 a_50751_n19729.t146 VSS 0.039522f
C10039 a_50751_n19729.n258 VSS 0.045401f
C10040 a_50751_n19729.t56 VSS 0.039522f
C10041 a_50751_n19729.t263 VSS 0.039477f
C10042 a_50751_n19729.n259 VSS 0.045123f
C10043 a_50751_n19729.t188 VSS 0.042148f
C10044 a_50751_n19729.n260 VSS 0.045377f
C10045 a_50751_n19729.t14 VSS 0.039522f
C10046 a_50751_n19729.n261 VSS 0.045401f
C10047 a_50751_n19729.t231 VSS 0.042151f
C10048 a_50751_n19729.t134 VSS 0.039522f
C10049 a_50751_n19729.n262 VSS 0.045401f
C10050 a_50751_n19729.t64 VSS 0.039522f
C10051 a_50751_n19729.t251 VSS 0.039475f
C10052 a_50751_n19729.n263 VSS 0.045377f
C10053 a_50751_n19729.t177 VSS 0.042148f
C10054 a_50751_n19729.n264 VSS 0.04511f
C10055 a_50751_n19729.t18 VSS 0.039522f
C10056 a_50751_n19729.n265 VSS 0.045401f
C10057 a_50751_n19729.t297 VSS 0.042151f
C10058 a_50751_n19729.t185 VSS 0.039522f
C10059 a_50751_n19729.n266 VSS 0.045401f
C10060 a_50751_n19729.t46 VSS 0.039522f
C10061 a_50751_n19729.t311 VSS 0.039522f
C10062 a_50751_n19729.n267 VSS 0.045377f
C10063 a_50751_n19729.t242 VSS 0.042148f
C10064 a_50751_n19729.n268 VSS 0.045377f
C10065 a_50751_n19729.t66 VSS 0.039522f
C10066 a_50751_n19729.n269 VSS 0.046427f
C10067 a_50751_n19729.t204 VSS 0.04212f
C10068 a_50751_n19729.t105 VSS 0.039526f
C10069 a_50751_n19729.n270 VSS 0.0454f
C10070 a_50751_n19729.t75 VSS 0.039526f
C10071 a_50751_n19729.t223 VSS 0.039526f
C10072 a_50751_n19729.n271 VSS 0.046401f
C10073 a_50751_n19729.t154 VSS 0.042116f
C10074 a_50751_n19729.n272 VSS 0.045377f
C10075 a_50751_n19729.n273 VSS 0.025282f
C10076 a_50751_n19729.n274 VSS 0.025095f
C10077 a_50751_n19729.t298 VSS 0.039493f
C10078 a_50751_n19729.n275 VSS 0.045401f
C10079 a_50751_n19729.t132 VSS 0.042151f
C10080 a_50751_n19729.t326 VSS 0.039522f
C10081 a_50751_n19729.n276 VSS 0.045401f
C10082 a_50751_n19729.t288 VSS 0.039522f
C10083 a_50751_n19729.t150 VSS 0.039522f
C10084 a_50751_n19729.n277 VSS 0.045377f
C10085 a_50751_n19729.t86 VSS 0.042148f
C10086 a_50751_n19729.n278 VSS 0.045377f
C10087 a_50751_n19729.t219 VSS 0.039522f
C10088 a_50751_n19729.n279 VSS 0.045401f
C10089 a_50751_n19729.t83 VSS 0.042151f
C10090 a_50751_n19729.t268 VSS 0.039522f
C10091 a_50751_n19729.n280 VSS 0.045401f
C10092 a_50751_n19729.t225 VSS 0.039522f
C10093 a_50751_n19729.t96 VSS 0.039522f
C10094 a_50751_n19729.n281 VSS 0.045377f
C10095 a_50751_n19729.t321 VSS 0.042148f
C10096 a_50751_n19729.n282 VSS 0.045377f
C10097 a_50751_n19729.t161 VSS 0.039522f
C10098 a_50751_n19729.n283 VSS 0.02429f
C10099 a_50751_n19729.t67 VSS 0.007577f
C10100 a_50751_n19729.n284 VSS 0.021461f
C10101 a_50751_n19729.t19 VSS 0.007577f
C10102 a_50751_n19729.n285 VSS 0.016705f
C10103 a_50751_n19729.t15 VSS 0.007577f
C10104 a_50751_n19729.n286 VSS 0.021443f
C10105 a_50751_n19729.n287 VSS 0.024116f
C10106 a_50751_n19729.n288 VSS 0.045401f
C10107 a_50751_n19729.t167 VSS 0.042151f
C10108 a_50751_n19729.t78 VSS 0.039522f
C10109 a_50751_n19729.n289 VSS 0.045401f
C10110 a_50751_n19729.t327 VSS 0.039522f
C10111 a_50751_n19729.t182 VSS 0.039522f
C10112 a_50751_n19729.n290 VSS 0.045377f
C10113 a_50751_n19729.t118 VSS 0.042148f
C10114 a_50751_n19729.n291 VSS 0.045377f
C10115 a_50751_n19729.t260 VSS 0.039522f
C10116 a_50751_n19729.n292 VSS 0.045401f
C10117 a_50751_n19729.t100 VSS 0.042151f
C10118 a_50751_n19729.t292 VSS 0.039522f
C10119 a_50751_n19729.n293 VSS 0.045401f
C10120 a_50751_n19729.t253 VSS 0.039522f
C10121 a_50751_n19729.t109 VSS 0.039522f
C10122 a_50751_n19729.n294 VSS 0.045377f
C10123 a_50751_n19729.t337 VSS 0.042148f
C10124 a_50751_n19729.n295 VSS 0.045377f
C10125 a_50751_n19729.t180 VSS 0.039522f
C10126 a_50751_n19729.n296 VSS 0.045401f
C10127 a_50751_n19729.t106 VSS 0.042151f
C10128 a_50751_n19729.t305 VSS 0.039522f
C10129 a_50751_n19729.n297 VSS 0.045401f
C10130 a_50751_n19729.t266 VSS 0.039522f
C10131 a_50751_n19729.t124 VSS 0.039472f
C10132 a_50751_n19729.n298 VSS 0.045097f
C10133 a_50751_n19729.t351 VSS 0.042148f
C10134 a_50751_n19729.n299 VSS 0.045377f
C10135 a_50751_n19729.t192 VSS 0.039522f
C10136 a_50751_n19729.t73 VSS 0.077435f
C10137 a_50751_n19729.t72 VSS 0.063772f
C10138 a_50751_n19729.n300 VSS 0.723314f
C10139 a_50751_n19729.t55 VSS 0.007577f
C10140 a_50751_n19729.n301 VSS 0.021871f
C10141 a_50751_n19729.t3 VSS 0.007577f
C10142 a_50751_n19729.n302 VSS 0.016705f
C10143 a_50751_n19729.t29 VSS 0.007577f
C10144 a_50751_n19729.n303 VSS 0.021816f
C10145 a_50751_n19729.t141 VSS 0.039522f
C10146 a_50751_n19729.t241 VSS 0.039472f
C10147 a_50751_n19729.n304 VSS 0.02267f
C10148 a_50751_n19729.n305 VSS 0.045097f
C10149 a_50751_n19729.t80 VSS 0.042148f
C10150 a_50751_n19729.n306 VSS 0.045377f
C10151 a_50751_n19729.n307 VSS 0.045401f
C10152 a_50751_n19729.t140 VSS 0.042151f
C10153 a_50751_n19729.t265 VSS 0.039522f
C10154 a_50751_n19729.n308 VSS 0.045401f
C10155 a_50751_n19729.t147 VSS 0.039522f
C10156 a_50751_n19729.n309 VSS 0.045401f
C10157 a_50751_n19729.t212 VSS 0.042151f
C10158 a_50751_n19729.t336 VSS 0.039522f
C10159 a_50751_n19729.n310 VSS 0.045401f
C10160 a_50751_n19729.t214 VSS 0.039522f
C10161 a_50751_n19729.t320 VSS 0.039522f
C10162 a_50751_n19729.n311 VSS 0.045377f
C10163 a_50751_n19729.t148 VSS 0.042148f
C10164 a_50751_n19729.n312 VSS 0.045377f
C10165 a_50751_n19729.t220 VSS 0.039522f
C10166 a_50751_n19729.n313 VSS 0.045401f
C10167 a_50751_n19729.t196 VSS 0.042151f
C10168 a_50751_n19729.t325 VSS 0.039522f
C10169 a_50751_n19729.n314 VSS 0.045401f
C10170 a_50751_n19729.t199 VSS 0.039522f
C10171 a_50751_n19729.t306 VSS 0.039522f
C10172 a_50751_n19729.n315 VSS 0.045377f
C10173 a_50751_n19729.t136 VSS 0.042148f
C10174 a_50751_n19729.n316 VSS 0.045377f
C10175 a_50751_n19729.t207 VSS 0.039522f
C10176 a_50751_n19729.n317 VSS 0.045401f
C10177 a_50751_n19729.t129 VSS 0.042151f
C10178 a_50751_n19729.t259 VSS 0.039522f
C10179 a_50751_n19729.n318 VSS 0.045401f
C10180 a_50751_n19729.t54 VSS 0.039522f
C10181 a_50751_n19729.t232 VSS 0.039522f
C10182 a_50751_n19729.n319 VSS 0.045377f
C10183 a_50751_n19729.t361 VSS 0.042148f
C10184 a_50751_n19729.n320 VSS 0.045377f
C10185 a_50751_n19729.t52 VSS 0.039522f
C10186 a_50751_n19729.n321 VSS 0.045401f
C10187 a_50751_n19729.t348 VSS 0.042151f
C10188 a_50751_n19729.t176 VSS 0.039522f
C10189 a_50751_n19729.n322 VSS 0.045401f
C10190 a_50751_n19729.t2 VSS 0.039522f
C10191 a_50751_n19729.t158 VSS 0.039475f
C10192 a_50751_n19729.n323 VSS 0.04511f
C10193 a_50751_n19729.t285 VSS 0.042148f
C10194 a_50751_n19729.n324 VSS 0.045377f
C10195 a_50751_n19729.t0 VSS 0.039522f
C10196 a_50751_n19729.n325 VSS 0.045401f
C10197 a_50751_n19729.t276 VSS 0.042151f
C10198 a_50751_n19729.t104 VSS 0.039522f
C10199 a_50751_n19729.n326 VSS 0.045401f
C10200 a_50751_n19729.t28 VSS 0.039522f
C10201 a_50751_n19729.t93 VSS 0.039477f
C10202 a_50751_n19729.n327 VSS 0.045377f
C10203 a_50751_n19729.t209 VSS 0.042148f
C10204 a_50751_n19729.n328 VSS 0.045123f
C10205 a_50751_n19729.t24 VSS 0.039522f
C10206 a_50751_n19729.n329 VSS 0.024116f
C10207 a_50751_n19729.t25 VSS 0.007577f
C10208 a_50751_n19729.n330 VSS 0.021443f
C10209 a_50751_n19729.t1 VSS 0.007577f
C10210 a_50751_n19729.n331 VSS 0.016705f
C10211 a_50751_n19729.t53 VSS 0.007577f
C10212 a_50751_n19729.n332 VSS 0.021461f
C10213 a_50751_n19729.n333 VSS 0.02429f
C10214 a_50751_n19729.n334 VSS 0.045401f
C10215 a_50751_n19729.t115 VSS 0.042151f
C10216 a_50751_n19729.t247 VSS 0.039522f
C10217 a_50751_n19729.n335 VSS 0.045401f
C10218 a_50751_n19729.t116 VSS 0.039522f
C10219 a_50751_n19729.t221 VSS 0.039522f
C10220 a_50751_n19729.n336 VSS 0.045377f
C10221 a_50751_n19729.t344 VSS 0.042148f
C10222 a_50751_n19729.n337 VSS 0.045377f
C10223 a_50751_n19729.t125 VSS 0.039522f
C10224 a_50751_n19729.n338 VSS 0.045401f
C10225 a_50751_n19729.t184 VSS 0.042151f
C10226 a_50751_n19729.t323 VSS 0.039522f
C10227 a_50751_n19729.n339 VSS 0.045401f
C10228 a_50751_n19729.t186 VSS 0.039522f
C10229 a_50751_n19729.t300 VSS 0.039522f
C10230 a_50751_n19729.n340 VSS 0.045377f
C10231 a_50751_n19729.t126 VSS 0.042148f
C10232 a_50751_n19729.n341 VSS 0.045377f
C10233 a_50751_n19729.t198 VSS 0.039522f
C10234 a_50751_n19729.n342 VSS 0.046427f
C10235 a_50751_n19729.t254 VSS 0.04212f
C10236 a_50751_n19729.t92 VSS 0.039526f
C10237 a_50751_n19729.n343 VSS 0.0454f
C10238 a_50751_n19729.t256 VSS 0.039526f
C10239 a_50751_n19729.t359 VSS 0.039526f
C10240 a_50751_n19729.n344 VSS 0.046401f
C10241 a_50751_n19729.t181 VSS 0.042116f
C10242 a_50751_n19729.n345 VSS 0.045377f
C10243 a_50751_n19729.n346 VSS 0.025282f
C10244 a_50751_n19729.n347 VSS 0.025095f
C10245 a_50751_n19729.t262 VSS 0.039493f
C10246 a_50751_n19729.t27 VSS 0.007577f
C10247 a_50751_n19729.n348 VSS 0.021816f
C10248 a_50751_n19729.t33 VSS 0.007577f
C10249 a_50751_n19729.n349 VSS 0.016705f
C10250 a_50751_n19729.t17 VSS 0.007577f
C10251 a_50751_n19729.n350 VSS 0.021871f
C10252 a_50751_n19729.n351 VSS 0.045401f
C10253 a_50751_n19729.t127 VSS 0.042151f
C10254 a_50751_n19729.t189 VSS 0.039522f
C10255 a_50751_n19729.n352 VSS 0.045401f
C10256 a_50751_n19729.t26 VSS 0.039522f
C10257 a_50751_n19729.t244 VSS 0.039477f
C10258 a_50751_n19729.n353 VSS 0.045123f
C10259 a_50751_n19729.t312 VSS 0.042148f
C10260 a_50751_n19729.n354 VSS 0.045377f
C10261 a_50751_n19729.t6 VSS 0.039522f
C10262 a_50751_n19729.n355 VSS 0.045401f
C10263 a_50751_n19729.t110 VSS 0.042151f
C10264 a_50751_n19729.t178 VSS 0.039522f
C10265 a_50751_n19729.n356 VSS 0.045401f
C10266 a_50751_n19729.t32 VSS 0.039522f
C10267 a_50751_n19729.t226 VSS 0.039475f
C10268 a_50751_n19729.n357 VSS 0.045377f
C10269 a_50751_n19729.t301 VSS 0.042148f
C10270 a_50751_n19729.n358 VSS 0.04511f
C10271 a_50751_n19729.t12 VSS 0.039522f
C10272 a_50751_n19729.n359 VSS 0.045401f
C10273 a_50751_n19729.t169 VSS 0.042151f
C10274 a_50751_n19729.t243 VSS 0.039522f
C10275 a_50751_n19729.n360 VSS 0.045401f
C10276 a_50751_n19729.t16 VSS 0.039522f
C10277 a_50751_n19729.t291 VSS 0.039522f
C10278 a_50751_n19729.n361 VSS 0.045377f
C10279 a_50751_n19729.t360 VSS 0.042148f
C10280 a_50751_n19729.n362 VSS 0.045377f
C10281 a_50751_n19729.t60 VSS 0.039522f
C10282 a_50751_n19729.n363 VSS 0.046427f
C10283 a_50751_n19729.t94 VSS 0.04212f
C10284 a_50751_n19729.t156 VSS 0.039526f
C10285 a_50751_n19729.n364 VSS 0.0454f
C10286 a_50751_n19729.t246 VSS 0.039526f
C10287 a_50751_n19729.t201 VSS 0.039526f
C10288 a_50751_n19729.n365 VSS 0.046401f
C10289 a_50751_n19729.t271 VSS 0.042116f
C10290 a_50751_n19729.n366 VSS 0.045377f
C10291 a_50751_n19729.n367 VSS 0.025282f
C10292 a_50751_n19729.n368 VSS 0.025095f
C10293 a_50751_n19729.t313 VSS 0.039493f
C10294 a_50751_n19729.n369 VSS 0.045401f
C10295 a_50751_n19729.t309 VSS 0.042151f
C10296 a_50751_n19729.t87 VSS 0.039522f
C10297 a_50751_n19729.n370 VSS 0.045401f
C10298 a_50751_n19729.t165 VSS 0.039522f
C10299 a_50751_n19729.t128 VSS 0.039522f
C10300 a_50751_n19729.n371 VSS 0.045377f
C10301 a_50751_n19729.t190 VSS 0.042148f
C10302 a_50751_n19729.n372 VSS 0.045377f
C10303 a_50751_n19729.t235 VSS 0.039522f
C10304 a_50751_n19729.n373 VSS 0.045401f
C10305 a_50751_n19729.t252 VSS 0.042151f
C10306 a_50751_n19729.t322 VSS 0.039522f
C10307 a_50751_n19729.n374 VSS 0.045401f
C10308 a_50751_n19729.t107 VSS 0.039522f
C10309 a_50751_n19729.t77 VSS 0.039522f
C10310 a_50751_n19729.n375 VSS 0.045377f
C10311 a_50751_n19729.t139 VSS 0.042148f
C10312 a_50751_n19729.n376 VSS 0.045377f
C10313 a_50751_n19729.t172 VSS 0.039522f
C10314 a_50751_n19729.n377 VSS 0.02429f
C10315 a_50751_n19729.t61 VSS 0.007577f
C10316 a_50751_n19729.n378 VSS 0.021461f
C10317 a_50751_n19729.t13 VSS 0.007577f
C10318 a_50751_n19729.n379 VSS 0.016705f
C10319 a_50751_n19729.t7 VSS 0.007577f
C10320 a_50751_n19729.n380 VSS 0.021443f
C10321 a_50751_n19729.n381 VSS 0.024116f
C10322 a_50751_n19729.n382 VSS 0.045401f
C10323 a_50751_n19729.t345 VSS 0.042151f
C10324 a_50751_n19729.t119 VSS 0.039522f
C10325 a_50751_n19729.n383 VSS 0.045401f
C10326 a_50751_n19729.t203 VSS 0.039522f
C10327 a_50751_n19729.t164 VSS 0.039522f
C10328 a_50751_n19729.n384 VSS 0.045377f
C10329 a_50751_n19729.t234 VSS 0.042148f
C10330 a_50751_n19729.n385 VSS 0.045377f
C10331 a_50751_n19729.t275 VSS 0.039522f
C10332 a_50751_n19729.n386 VSS 0.045401f
C10333 a_50751_n19729.t272 VSS 0.042151f
C10334 a_50751_n19729.t338 VSS 0.039522f
C10335 a_50751_n19729.n387 VSS 0.045401f
C10336 a_50751_n19729.t131 VSS 0.039522f
C10337 a_50751_n19729.t97 VSS 0.039522f
C10338 a_50751_n19729.n388 VSS 0.045377f
C10339 a_50751_n19729.t160 VSS 0.042148f
C10340 a_50751_n19729.n389 VSS 0.045377f
C10341 a_50751_n19729.t195 VSS 0.039522f
C10342 a_50751_n19729.n390 VSS 0.045401f
C10343 a_50751_n19729.t286 VSS 0.042151f
C10344 a_50751_n19729.t352 VSS 0.039522f
C10345 a_50751_n19729.n391 VSS 0.045401f
C10346 a_50751_n19729.t144 VSS 0.039522f
C10347 a_50751_n19729.t102 VSS 0.039472f
C10348 a_50751_n19729.n392 VSS 0.045097f
C10349 a_50751_n19729.t168 VSS 0.042148f
C10350 a_50751_n19729.n393 VSS 0.045377f
C10351 a_50751_n19729.t211 VSS 0.039522f
C10352 a_50751_n19729.n394 VSS 0.107128f
C10353 a_50751_n19729.n395 VSS 0.440026f
C10354 a_50751_n19729.t43 VSS 0.007577f
C10355 a_50751_n19729.n396 VSS 0.021871f
C10356 a_50751_n19729.t63 VSS 0.007577f
C10357 a_50751_n19729.n397 VSS 0.016705f
C10358 a_50751_n19729.t21 VSS 0.007577f
C10359 a_50751_n19729.n398 VSS 0.021816f
C10360 a_50751_n19729.t175 VSS 0.039522f
C10361 a_50751_n19729.t293 VSS 0.039472f
C10362 a_50751_n19729.n399 VSS 0.02267f
C10363 a_50751_n19729.n400 VSS 0.045097f
C10364 a_50751_n19729.t215 VSS 0.042148f
C10365 a_50751_n19729.n401 VSS 0.045377f
C10366 a_50751_n19729.n402 VSS 0.045401f
C10367 a_50751_n19729.t257 VSS 0.042151f
C10368 a_50751_n19729.t282 VSS 0.039522f
C10369 a_50751_n19729.n403 VSS 0.045401f
C10370 a_50751_n19729.t95 VSS 0.039522f
C10371 a_50751_n19729.n404 VSS 0.045401f
C10372 a_50751_n19729.t328 VSS 0.042151f
C10373 a_50751_n19729.t356 VSS 0.039522f
C10374 a_50751_n19729.n405 VSS 0.045401f
C10375 a_50751_n19729.t258 VSS 0.039522f
C10376 a_50751_n19729.t79 VSS 0.039522f
C10377 a_50751_n19729.n406 VSS 0.045377f
C10378 a_50751_n19729.t289 VSS 0.042148f
C10379 a_50751_n19729.n407 VSS 0.045377f
C10380 a_50751_n19729.t162 VSS 0.039522f
C10381 a_50751_n19729.n408 VSS 0.045401f
C10382 a_50751_n19729.t319 VSS 0.042151f
C10383 a_50751_n19729.t340 VSS 0.039522f
C10384 a_50751_n19729.n409 VSS 0.045401f
C10385 a_50751_n19729.t245 VSS 0.039522f
C10386 a_50751_n19729.t354 VSS 0.039522f
C10387 a_50751_n19729.n410 VSS 0.045377f
C10388 a_50751_n19729.t280 VSS 0.042148f
C10389 a_50751_n19729.n411 VSS 0.045377f
C10390 a_50751_n19729.t151 VSS 0.039522f
C10391 a_50751_n19729.n412 VSS 0.045401f
C10392 a_50751_n19729.t249 VSS 0.042151f
C10393 a_50751_n19729.t273 VSS 0.039522f
C10394 a_50751_n19729.n413 VSS 0.045401f
C10395 a_50751_n19729.t42 VSS 0.039522f
C10396 a_50751_n19729.t283 VSS 0.039522f
C10397 a_50751_n19729.n414 VSS 0.045377f
C10398 a_50751_n19729.t202 VSS 0.042148f
C10399 a_50751_n19729.n415 VSS 0.045377f
C10400 a_50751_n19729.t68 VSS 0.039522f
C10401 a_50751_n19729.n416 VSS 0.045401f
C10402 a_50751_n19729.t166 VSS 0.042151f
C10403 a_50751_n19729.t193 VSS 0.039522f
C10404 a_50751_n19729.n417 VSS 0.045401f
C10405 a_50751_n19729.t62 VSS 0.039522f
C10406 a_50751_n19729.t206 VSS 0.039475f
C10407 a_50751_n19729.n418 VSS 0.04511f
C10408 a_50751_n19729.t130 VSS 0.042148f
C10409 a_50751_n19729.n419 VSS 0.045377f
C10410 a_50751_n19729.t22 VSS 0.039522f
C10411 a_50751_n19729.n420 VSS 0.045401f
C10412 a_50751_n19729.t99 VSS 0.042151f
C10413 a_50751_n19729.t121 VSS 0.039522f
C10414 a_50751_n19729.n421 VSS 0.045401f
C10415 a_50751_n19729.t20 VSS 0.039522f
C10416 a_50751_n19729.t135 VSS 0.039477f
C10417 a_50751_n19729.n422 VSS 0.045377f
C10418 a_50751_n19729.t350 VSS 0.042148f
C10419 a_50751_n19729.n423 VSS 0.045123f
C10420 a_50751_n19729.t34 VSS 0.039522f
C10421 a_50751_n19729.n424 VSS 0.024116f
C10422 a_50751_n19729.t35 VSS 0.007577f
C10423 a_50751_n19729.n425 VSS 0.021443f
C10424 a_50751_n19729.t23 VSS 0.007577f
C10425 a_50751_n19729.n426 VSS 0.016705f
C10426 a_50751_n19729.t69 VSS 0.007577f
C10427 a_50751_n19729.n427 VSS 0.021461f
C10428 a_50751_n19729.n428 VSS 0.02429f
C10429 a_50751_n19729.n429 VSS 0.045401f
C10430 a_50751_n19729.t230 VSS 0.042151f
C10431 a_50751_n19729.t261 VSS 0.039522f
C10432 a_50751_n19729.n430 VSS 0.045401f
C10433 a_50751_n19729.t159 VSS 0.039522f
C10434 a_50751_n19729.t270 VSS 0.039522f
C10435 a_50751_n19729.n431 VSS 0.045377f
C10436 a_50751_n19729.t187 VSS 0.042148f
C10437 a_50751_n19729.n432 VSS 0.045377f
C10438 a_50751_n19729.t74 VSS 0.039522f
C10439 a_50751_n19729.n433 VSS 0.045401f
C10440 a_50751_n19729.t310 VSS 0.042151f
C10441 a_50751_n19729.t330 VSS 0.039522f
C10442 a_50751_n19729.n434 VSS 0.045401f
C10443 a_50751_n19729.t233 VSS 0.039522f
C10444 a_50751_n19729.t343 VSS 0.039522f
C10445 a_50751_n19729.n435 VSS 0.045377f
C10446 a_50751_n19729.t269 VSS 0.042148f
C10447 a_50751_n19729.n436 VSS 0.045377f
C10448 a_50751_n19729.t142 VSS 0.039522f
C10449 a_50751_n19729.n437 VSS 0.046427f
C10450 a_50751_n19729.t82 VSS 0.04212f
C10451 a_50751_n19729.t101 VSS 0.039526f
C10452 a_50751_n19729.n438 VSS 0.0454f
C10453 a_50751_n19729.t299 VSS 0.039526f
C10454 a_50751_n19729.t108 VSS 0.039526f
C10455 a_50751_n19729.n439 VSS 0.046401f
C10456 a_50751_n19729.t329 VSS 0.042116f
C10457 a_50751_n19729.n440 VSS 0.045377f
C10458 a_50751_n19729.n441 VSS 0.025282f
C10459 a_50751_n19729.n442 VSS 0.025095f
C10460 a_50751_n19729.t200 VSS 0.039493f
C10461 a_50751_n19729.t5 VSS 0.007577f
C10462 a_50751_n19729.n443 VSS 0.021816f
C10463 a_50751_n19729.t11 VSS 0.007577f
C10464 a_50751_n19729.n444 VSS 0.016705f
C10465 a_50751_n19729.t59 VSS 0.007577f
C10466 a_50751_n19729.n445 VSS 0.021871f
C10467 a_50751_n19729.n446 VSS 0.045401f
C10468 a_50751_n19729.t98 VSS 0.042151f
C10469 a_50751_n19729.t191 VSS 0.039522f
C10470 a_50751_n19729.n447 VSS 0.045401f
C10471 a_50751_n19729.t4 VSS 0.039522f
C10472 a_50751_n19729.t117 VSS 0.039477f
C10473 a_50751_n19729.n448 VSS 0.045123f
C10474 a_50751_n19729.t183 VSS 0.042148f
C10475 a_50751_n19729.n449 VSS 0.045377f
C10476 a_50751_n19729.t44 VSS 0.039522f
C10477 a_50751_n19729.n450 VSS 0.045401f
C10478 a_50751_n19729.t91 VSS 0.042151f
C10479 a_50751_n19729.t179 VSS 0.039522f
C10480 a_50751_n19729.n451 VSS 0.045401f
C10481 a_50751_n19729.t10 VSS 0.039522f
C10482 a_50751_n19729.t103 VSS 0.039475f
C10483 a_50751_n19729.n452 VSS 0.045377f
C10484 a_50751_n19729.t174 VSS 0.042148f
C10485 a_50751_n19729.n453 VSS 0.04511f
C10486 a_50751_n19729.t50 VSS 0.039522f
C10487 a_50751_n19729.n454 VSS 0.045401f
C10488 a_50751_n19729.t143 VSS 0.042151f
C10489 a_50751_n19729.t248 VSS 0.039522f
C10490 a_50751_n19729.n455 VSS 0.045401f
C10491 a_50751_n19729.t58 VSS 0.039522f
C10492 a_50751_n19729.t163 VSS 0.039522f
C10493 a_50751_n19729.n456 VSS 0.045377f
C10494 a_50751_n19729.t238 VSS 0.042148f
C10495 a_50751_n19729.n457 VSS 0.045377f
C10496 a_50751_n19729.t38 VSS 0.039522f
C10497 a_50751_n19729.n458 VSS 0.046427f
C10498 a_50751_n19729.t349 VSS 0.04212f
C10499 a_50751_n19729.t157 VSS 0.039526f
C10500 a_50751_n19729.n459 VSS 0.0454f
C10501 a_50751_n19729.t314 VSS 0.039526f
C10502 a_50751_n19729.t85 VSS 0.039526f
C10503 a_50751_n19729.n460 VSS 0.046401f
C10504 a_50751_n19729.t153 VSS 0.042116f
C10505 a_50751_n19729.n461 VSS 0.045377f
C10506 a_50751_n19729.n462 VSS 0.025282f
C10507 a_50751_n19729.n463 VSS 0.025095f
C10508 a_50751_n19729.t113 VSS 0.039493f
C10509 a_50751_n19729.n464 VSS 0.045401f
C10510 a_50751_n19729.t279 VSS 0.042151f
C10511 a_50751_n19729.t90 VSS 0.039522f
C10512 a_50751_n19729.n465 VSS 0.045401f
C10513 a_50751_n19729.t236 VSS 0.039522f
C10514 a_50751_n19729.t302 VSS 0.039522f
C10515 a_50751_n19729.n466 VSS 0.045377f
C10516 a_50751_n19729.t84 VSS 0.042148f
C10517 a_50751_n19729.n467 VSS 0.045377f
C10518 a_50751_n19729.t333 VSS 0.039522f
C10519 a_50751_n19729.n468 VSS 0.045401f
C10520 a_50751_n19729.t218 VSS 0.042151f
C10521 a_50751_n19729.t324 VSS 0.039522f
C10522 a_50751_n19729.n469 VSS 0.045401f
C10523 a_50751_n19729.t173 VSS 0.039522f
C10524 a_50751_n19729.t240 VSS 0.039522f
C10525 a_50751_n19729.n470 VSS 0.045377f
C10526 a_50751_n19729.t317 VSS 0.042148f
C10527 a_50751_n19729.n471 VSS 0.045377f
C10528 a_50751_n19729.t281 VSS 0.039522f
C10529 a_50751_n19729.n472 VSS 0.02429f
C10530 a_50751_n19729.t39 VSS 0.007577f
C10531 a_50751_n19729.n473 VSS 0.021461f
C10532 a_50751_n19729.t51 VSS 0.007577f
C10533 a_50751_n19729.n474 VSS 0.016705f
C10534 a_50751_n19729.t45 VSS 0.007577f
C10535 a_50751_n19729.n475 VSS 0.021443f
C10536 a_50751_n19729.n476 VSS 0.024116f
C10537 a_50751_n19729.n477 VSS 0.045401f
C10538 a_50751_n19729.t318 VSS 0.042151f
C10539 a_50751_n19729.t120 VSS 0.039522f
C10540 a_50751_n19729.n478 VSS 0.045401f
C10541 a_50751_n19729.t277 VSS 0.039522f
C10542 a_50751_n19729.t335 VSS 0.039522f
C10543 a_50751_n19729.n479 VSS 0.045377f
C10544 a_50751_n19729.t114 VSS 0.042148f
C10545 a_50751_n19729.n480 VSS 0.045377f
C10546 a_50751_n19729.t89 VSS 0.039522f
C10547 a_50751_n19729.n481 VSS 0.045401f
C10548 a_50751_n19729.t239 VSS 0.042151f
C10549 a_50751_n19729.t339 VSS 0.039522f
C10550 a_50751_n19729.n482 VSS 0.045401f
C10551 a_50751_n19729.t197 VSS 0.039522f
C10552 a_50751_n19729.t264 VSS 0.039522f
C10553 a_50751_n19729.n483 VSS 0.045377f
C10554 a_50751_n19729.t334 VSS 0.042148f
C10555 a_50751_n19729.n484 VSS 0.045377f
C10556 a_50751_n19729.t304 VSS 0.039522f
C10557 a_50751_n19729.n485 VSS 0.045401f
C10558 a_50751_n19729.t255 VSS 0.042151f
C10559 a_50751_n19729.t355 VSS 0.039522f
C10560 a_50751_n19729.n486 VSS 0.045401f
C10561 a_50751_n19729.t213 VSS 0.039522f
C10562 a_50751_n19729.t278 VSS 0.039472f
C10563 a_50751_n19729.n487 VSS 0.045097f
C10564 a_50751_n19729.t347 VSS 0.042148f
C10565 a_50751_n19729.n488 VSS 0.045377f
C10566 a_50751_n19729.t316 VSS 0.039522f
C10567 a_50751_n19729.n489 VSS 0.107128f
C10568 a_50751_n19729.n490 VSS 0.256981f
C10569 a_50751_n19729.n491 VSS 0.208715f
C10570 a_50751_n19729.n492 VSS 0.046427f
C10571 a_50751_n19729.t170 VSS 0.04212f
C10572 a_50751_n19729.t267 VSS 0.039526f
C10573 a_50751_n19729.n493 VSS 0.0454f
C10574 a_50751_n19729.t171 VSS 0.039526f
C10575 a_50751_n19729.t353 VSS 0.039526f
C10576 a_50751_n19729.n494 VSS 0.046401f
C10577 a_50751_n19729.t342 VSS 0.042116f
C10578 a_50751_n19729.n495 VSS 0.045377f
C10579 a_50751_n19729.n496 VSS 0.025282f
C10580 a_50751_n19729.n497 VSS 0.025095f
C10581 a_50751_n19729.t341 VSS 0.039493f
C10582 a_50751_n19729.n498 VSS 0.045401f
C10583 a_50751_n19729.t111 VSS 0.042151f
C10584 a_50751_n19729.t205 VSS 0.039522f
C10585 a_50751_n19729.n499 VSS 0.045401f
C10586 a_50751_n19729.t112 VSS 0.039522f
C10587 a_50751_n19729.t295 VSS 0.039522f
C10588 a_50751_n19729.n500 VSS 0.045377f
C10589 a_50751_n19729.t287 VSS 0.042148f
C10590 a_50751_n19729.n501 VSS 0.045377f
C10591 a_50751_n19729.t284 VSS 0.039522f
C10592 a_50751_n19729.n502 VSS 0.045401f
C10593 a_50751_n19729.t331 VSS 0.042151f
C10594 a_50751_n19729.t133 VSS 0.039522f
C10595 a_50751_n19729.n503 VSS 0.045401f
C10596 a_50751_n19729.t332 VSS 0.039522f
C10597 a_50751_n19729.t217 VSS 0.039522f
C10598 a_50751_n19729.n504 VSS 0.045377f
C10599 a_50751_n19729.t210 VSS 0.042148f
C10600 a_50751_n19729.n505 VSS 0.045377f
C10601 a_50751_n19729.t208 VSS 0.039522f
C10602 a_50751_n19729.n506 VSS 0.02429f
C10603 a_50751_n19729.t37 VSS 0.007577f
C10604 a_50751_n19729.n507 VSS 0.021461f
C10605 a_50751_n19729.t49 VSS 0.007577f
C10606 a_50751_n19729.n508 VSS 0.016705f
C10607 a_50751_n19729.n509 VSS 0.021443f
C10608 a_50751_n19729.t71 VSS 0.007577f
C10609 a_52635_48695.n0 VSS 0.756922f
C10610 a_52635_48695.n1 VSS 1.21873f
C10611 a_52635_48695.n2 VSS 1.21872f
C10612 a_52635_48695.n3 VSS 1.18681f
C10613 a_52635_48695.n4 VSS 0.489342f
C10614 a_52635_48695.n5 VSS 1.21873f
C10615 a_52635_48695.n6 VSS 1.71719f
C10616 a_52635_48695.n7 VSS 1.52681f
C10617 a_52635_48695.n8 VSS 1.21873f
C10618 a_52635_48695.n9 VSS 1.21872f
C10619 a_52635_48695.n10 VSS 1.18681f
C10620 a_52635_48695.n11 VSS 0.489342f
C10621 a_52635_48695.n12 VSS 1.21873f
C10622 a_52635_48695.n13 VSS 1.71719f
C10623 a_52635_48695.n14 VSS 1.2057f
C10624 a_52635_48695.n15 VSS 1.0473f
C10625 a_52635_48695.n16 VSS 1.14869f
C10626 a_52635_48695.n17 VSS 0.784705f
C10627 a_52635_48695.n18 VSS 1.16549f
C10628 a_52635_48695.n19 VSS 1.16549f
C10629 a_52635_48695.n20 VSS 0.618892f
C10630 a_52635_48695.n21 VSS 1.0473f
C10631 a_52635_48695.n22 VSS 1.14869f
C10632 a_52635_48695.n23 VSS 1.36844f
C10633 a_52635_48695.n24 VSS 1.2057f
C10634 a_52635_48695.n25 VSS 1.0473f
C10635 a_52635_48695.n26 VSS 1.14869f
C10636 a_52635_48695.n27 VSS 0.784705f
C10637 a_52635_48695.n28 VSS 1.16549f
C10638 a_52635_48695.n29 VSS 1.16549f
C10639 a_52635_48695.n30 VSS 0.618892f
C10640 a_52635_48695.n31 VSS 1.0473f
C10641 a_52635_48695.n32 VSS 1.14869f
C10642 a_52635_48695.n33 VSS 1.36844f
C10643 a_52635_48695.t35 VSS 0.095327f
C10644 a_52635_48695.t13 VSS 0.095327f
C10645 a_52635_48695.t17 VSS 0.095327f
C10646 a_52635_48695.n34 VSS 0.349727f
C10647 a_52635_48695.n35 VSS 1.21985f
C10648 a_52635_48695.t2 VSS 0.095327f
C10649 a_52635_48695.t28 VSS 0.095327f
C10650 a_52635_48695.n36 VSS 0.523718f
C10651 a_52635_48695.t1 VSS 0.095327f
C10652 a_52635_48695.t58 VSS 0.095327f
C10653 a_52635_48695.n37 VSS 0.349727f
C10654 a_52635_48695.n38 VSS 1.72003f
C10655 a_52635_48695.t9 VSS 0.095327f
C10656 a_52635_48695.t45 VSS 0.095327f
C10657 a_52635_48695.n39 VSS 0.349727f
C10658 a_52635_48695.n40 VSS 1.21988f
C10659 a_52635_48695.t20 VSS 0.095327f
C10660 a_52635_48695.t12 VSS 0.095327f
C10661 a_52635_48695.n41 VSS 0.349727f
C10662 a_52635_48695.n42 VSS 0.489952f
C10663 a_52635_48695.n43 VSS 6.43054f
C10664 a_52635_48695.n44 VSS 3.88654f
C10665 a_52635_48695.t43 VSS 0.095327f
C10666 a_52635_48695.t34 VSS 0.095327f
C10667 a_52635_48695.n45 VSS 0.262987f
C10668 a_52635_48695.t48 VSS 0.095327f
C10669 a_52635_48695.t42 VSS 0.095327f
C10670 a_52635_48695.n46 VSS 0.240154f
C10671 a_52635_48695.n47 VSS 1.47747f
C10672 a_52635_48695.t66 VSS 0.269047f
C10673 a_52635_48695.t75 VSS 0.249659f
C10674 a_52635_48695.n48 VSS 0.855653f
C10675 a_52635_48695.n49 VSS 1.69542f
C10676 a_52635_48695.n50 VSS 4.5114f
C10677 a_52635_48695.t102 VSS 0.53874f
C10678 a_52635_48695.t134 VSS 0.095327f
C10679 a_52635_48695.t101 VSS 0.095327f
C10680 a_52635_48695.n51 VSS 0.411842f
C10681 a_52635_48695.t88 VSS 0.403741f
C10682 a_52635_48695.t108 VSS 0.403217f
C10683 a_52635_48695.n52 VSS 3.88906f
C10684 a_52635_48695.t161 VSS 0.533719f
C10685 a_52635_48695.t97 VSS 0.095327f
C10686 a_52635_48695.t160 VSS 0.095327f
C10687 a_52635_48695.n53 VSS 0.412681f
C10688 a_52635_48695.n54 VSS 1.35842f
C10689 a_52635_48695.t144 VSS 0.404562f
C10690 a_52635_48695.n55 VSS 1.14974f
C10691 a_52635_48695.t165 VSS 0.4011f
C10692 a_52635_48695.n56 VSS 1.04175f
C10693 a_52635_48695.t92 VSS 0.541236f
C10694 a_52635_48695.t137 VSS 0.095327f
C10695 a_52635_48695.t118 VSS 0.095327f
C10696 a_52635_48695.n57 VSS 0.412681f
C10697 a_52635_48695.n58 VSS 1.21146f
C10698 a_52635_48695.t142 VSS 0.541236f
C10699 a_52635_48695.t94 VSS 0.095327f
C10700 a_52635_48695.t172 VSS 0.095327f
C10701 a_52635_48695.n59 VSS 0.412681f
C10702 a_52635_48695.n60 VSS 1.21146f
C10703 a_52635_48695.n61 VSS 0.928757f
C10704 a_52635_48695.t166 VSS 0.234955f
C10705 a_52635_48695.t95 VSS 0.286675f
C10706 a_52635_48695.n62 VSS 1.53633f
C10707 a_52635_48695.t158 VSS 0.095327f
C10708 a_52635_48695.t109 VSS 0.095327f
C10709 a_52635_48695.n63 VSS 0.223101f
C10710 a_52635_48695.t93 VSS 0.095327f
C10711 a_52635_48695.t133 VSS 0.095327f
C10712 a_52635_48695.n64 VSS 0.283831f
C10713 a_52635_48695.n65 VSS 0.646018f
C10714 a_52635_48695.n66 VSS 1.41217f
C10715 a_52635_48695.t125 VSS 0.533719f
C10716 a_52635_48695.t154 VSS 0.095327f
C10717 a_52635_48695.t124 VSS 0.095327f
C10718 a_52635_48695.n67 VSS 0.412681f
C10719 a_52635_48695.n68 VSS 1.35842f
C10720 a_52635_48695.t99 VSS 0.404562f
C10721 a_52635_48695.n69 VSS 1.14974f
C10722 a_52635_48695.t127 VSS 0.4011f
C10723 a_52635_48695.n70 VSS 1.04175f
C10724 a_52635_48695.t138 VSS 0.4011f
C10725 a_52635_48695.n71 VSS 1.04175f
C10726 a_52635_48695.t135 VSS 0.404562f
C10727 a_52635_48695.n72 VSS 1.14974f
C10728 a_52635_48695.t162 VSS 0.095327f
C10729 a_52635_48695.t132 VSS 0.095327f
C10730 a_52635_48695.n73 VSS 0.412681f
C10731 a_52635_48695.n74 VSS 0.784406f
C10732 a_52635_48695.t123 VSS 0.4011f
C10733 a_52635_48695.n75 VSS 1.157f
C10734 a_52635_48695.t131 VSS 0.404449f
C10735 a_52635_48695.n76 VSS 1.16648f
C10736 a_52635_48695.t169 VSS 0.095327f
C10737 a_52635_48695.t141 VSS 0.095327f
C10738 a_52635_48695.n77 VSS 0.412681f
C10739 a_52635_48695.n78 VSS 0.6193f
C10740 a_52635_48695.n79 VSS 0.928757f
C10741 a_52635_48695.n80 VSS 5.47584f
C10742 a_52635_48695.n81 VSS 1.80962f
C10743 a_52635_48695.t106 VSS 0.234955f
C10744 a_52635_48695.t128 VSS 0.286675f
C10745 a_52635_48695.n82 VSS 0.840134f
C10746 a_52635_48695.n83 VSS 1.71719f
C10747 a_52635_48695.t167 VSS 0.095327f
C10748 a_52635_48695.t120 VSS 0.095327f
C10749 a_52635_48695.n84 VSS 0.223101f
C10750 a_52635_48695.t96 VSS 0.095327f
C10751 a_52635_48695.t143 VSS 0.095327f
C10752 a_52635_48695.n85 VSS 0.283831f
C10753 a_52635_48695.n86 VSS 0.646018f
C10754 a_52635_48695.n87 VSS 1.12283f
C10755 a_52635_48695.n88 VSS 6.07046f
C10756 a_52635_48695.t130 VSS 0.53874f
C10757 a_52635_48695.t159 VSS 0.095327f
C10758 a_52635_48695.t129 VSS 0.095327f
C10759 a_52635_48695.n89 VSS 0.411842f
C10760 a_52635_48695.t110 VSS 0.403741f
C10761 a_52635_48695.t136 VSS 0.403217f
C10762 a_52635_48695.n90 VSS 0.265724f
C10763 a_52635_48695.t89 VSS 0.095327f
C10764 a_52635_48695.t149 VSS 0.095327f
C10765 a_52635_48695.n91 VSS 0.411842f
C10766 a_52635_48695.t139 VSS 0.403741f
C10767 a_52635_48695.t126 VSS 0.403741f
C10768 a_52635_48695.t168 VSS 0.095327f
C10769 a_52635_48695.t140 VSS 0.095327f
C10770 a_52635_48695.n92 VSS 0.411842f
C10771 a_52635_48695.t145 VSS 0.403741f
C10772 a_52635_48695.t147 VSS 0.403217f
C10773 a_52635_48695.t103 VSS 0.095327f
C10774 a_52635_48695.t91 VSS 0.095327f
C10775 a_52635_48695.n93 VSS 0.411842f
C10776 a_52635_48695.t150 VSS 0.539462f
C10777 a_52635_48695.n94 VSS 0.265724f
C10778 a_52635_48695.n95 VSS 3.88906f
C10779 a_52635_48695.n96 VSS 3.49604f
C10780 a_52635_48695.n97 VSS 0.265735f
C10781 a_52635_48695.t175 VSS 0.4011f
C10782 a_52635_48695.n98 VSS 1.04175f
C10783 a_52635_48695.t174 VSS 0.404562f
C10784 a_52635_48695.n99 VSS 1.14974f
C10785 a_52635_48695.t107 VSS 0.095327f
C10786 a_52635_48695.t171 VSS 0.095327f
C10787 a_52635_48695.n100 VSS 0.412681f
C10788 a_52635_48695.n101 VSS 0.784406f
C10789 a_52635_48695.t157 VSS 0.4011f
C10790 a_52635_48695.n102 VSS 1.157f
C10791 a_52635_48695.t170 VSS 0.404449f
C10792 a_52635_48695.n103 VSS 1.16648f
C10793 a_52635_48695.t117 VSS 0.095327f
C10794 a_52635_48695.t90 VSS 0.095327f
C10795 a_52635_48695.n104 VSS 0.412681f
C10796 a_52635_48695.n105 VSS 0.6193f
C10797 a_52635_48695.n106 VSS 0.265735f
C10798 a_52635_48695.n107 VSS 3.49604f
C10799 a_52635_48695.t114 VSS 0.234955f
C10800 a_52635_48695.t163 VSS 0.286675f
C10801 a_52635_48695.n108 VSS 1.53633f
C10802 a_52635_48695.t105 VSS 0.095327f
C10803 a_52635_48695.t151 VSS 0.095327f
C10804 a_52635_48695.n109 VSS 0.223101f
C10805 a_52635_48695.t156 VSS 0.095327f
C10806 a_52635_48695.t104 VSS 0.095327f
C10807 a_52635_48695.n110 VSS 0.283831f
C10808 a_52635_48695.n111 VSS 0.646018f
C10809 a_52635_48695.n112 VSS 1.41217f
C10810 a_52635_48695.t115 VSS 0.095327f
C10811 a_52635_48695.t155 VSS 0.095327f
C10812 a_52635_48695.n113 VSS 0.223101f
C10813 a_52635_48695.t164 VSS 0.095327f
C10814 a_52635_48695.t113 VSS 0.095327f
C10815 a_52635_48695.n114 VSS 0.283831f
C10816 a_52635_48695.n115 VSS 0.646018f
C10817 a_52635_48695.n116 VSS 1.12283f
C10818 a_52635_48695.t148 VSS 0.234955f
C10819 a_52635_48695.t100 VSS 0.286675f
C10820 a_52635_48695.n117 VSS 0.840134f
C10821 a_52635_48695.n118 VSS 1.71719f
C10822 a_52635_48695.n119 VSS 1.80962f
C10823 a_52635_48695.n120 VSS 3.91678f
C10824 a_52635_48695.n121 VSS 4.55814f
C10825 a_52635_48695.n122 VSS 0.265724f
C10826 a_52635_48695.t152 VSS 0.095327f
C10827 a_52635_48695.t121 VSS 0.095327f
C10828 a_52635_48695.n123 VSS 0.411842f
C10829 a_52635_48695.t111 VSS 0.403741f
C10830 a_52635_48695.t98 VSS 0.403741f
C10831 a_52635_48695.t146 VSS 0.095327f
C10832 a_52635_48695.t112 VSS 0.095327f
C10833 a_52635_48695.n124 VSS 0.411842f
C10834 a_52635_48695.t116 VSS 0.403741f
C10835 a_52635_48695.t119 VSS 0.403217f
C10836 a_52635_48695.t173 VSS 0.095327f
C10837 a_52635_48695.t153 VSS 0.095327f
C10838 a_52635_48695.n125 VSS 0.411842f
C10839 a_52635_48695.t122 VSS 0.539462f
C10840 a_52635_48695.n126 VSS 0.265724f
C10841 a_52635_48695.n127 VSS 4.10938f
C10842 a_52635_48695.n128 VSS 6.28374f
C10843 a_52635_48695.t19 VSS 0.095327f
C10844 a_52635_48695.t54 VSS 0.095327f
C10845 a_52635_48695.n129 VSS 0.349727f
C10846 a_52635_48695.n130 VSS 1.21988f
C10847 a_52635_48695.t46 VSS 0.095327f
C10848 a_52635_48695.t21 VSS 0.095327f
C10849 a_52635_48695.n131 VSS 0.349727f
C10850 a_52635_48695.n132 VSS 0.750098f
C10851 a_52635_48695.n133 VSS 5.24514f
C10852 a_52635_48695.n134 VSS 6.10701f
C10853 a_52635_48695.t82 VSS 0.095327f
C10854 a_52635_48695.t24 VSS 0.095327f
C10855 a_52635_48695.n135 VSS 0.523718f
C10856 a_52635_48695.t81 VSS 0.095327f
C10857 a_52635_48695.t55 VSS 0.095327f
C10858 a_52635_48695.n136 VSS 0.349727f
C10859 a_52635_48695.n137 VSS 1.72003f
C10860 a_52635_48695.t3 VSS 0.095327f
C10861 a_52635_48695.t39 VSS 0.095327f
C10862 a_52635_48695.n138 VSS 0.349727f
C10863 a_52635_48695.n139 VSS 1.21988f
C10864 a_52635_48695.t15 VSS 0.095327f
C10865 a_52635_48695.t6 VSS 0.095327f
C10866 a_52635_48695.n140 VSS 0.349727f
C10867 a_52635_48695.n141 VSS 0.489952f
C10868 a_52635_48695.t61 VSS 0.095327f
C10869 a_52635_48695.t16 VSS 0.095327f
C10870 a_52635_48695.n142 VSS 0.522376f
C10871 a_52635_48695.t60 VSS 0.095327f
C10872 a_52635_48695.t50 VSS 0.095327f
C10873 a_52635_48695.n143 VSS 0.348711f
C10874 a_52635_48695.t65 VSS 0.095327f
C10875 a_52635_48695.t25 VSS 0.095327f
C10876 a_52635_48695.n144 VSS 0.348711f
C10877 a_52635_48695.t83 VSS 0.095327f
C10878 a_52635_48695.t68 VSS 0.095327f
C10879 a_52635_48695.n145 VSS 0.348711f
C10880 a_52635_48695.t56 VSS 0.095327f
C10881 a_52635_48695.t22 VSS 0.095327f
C10882 a_52635_48695.n146 VSS 0.348711f
C10883 a_52635_48695.t69 VSS 0.095327f
C10884 a_52635_48695.t76 VSS 0.095327f
C10885 a_52635_48695.n147 VSS 0.348711f
C10886 a_52635_48695.t78 VSS 0.095327f
C10887 a_52635_48695.t47 VSS 0.095327f
C10888 a_52635_48695.n148 VSS 0.348711f
C10889 a_52635_48695.t26 VSS 0.095327f
C10890 a_52635_48695.t84 VSS 0.095327f
C10891 a_52635_48695.n149 VSS 0.348711f
C10892 a_52635_48695.n150 VSS 1.64071f
C10893 a_52635_48695.t36 VSS 0.095327f
C10894 a_52635_48695.t29 VSS 0.095327f
C10895 a_52635_48695.n151 VSS 0.262987f
C10896 a_52635_48695.t38 VSS 0.095327f
C10897 a_52635_48695.t30 VSS 0.095327f
C10898 a_52635_48695.n152 VSS 0.240154f
C10899 a_52635_48695.n153 VSS 1.47747f
C10900 a_52635_48695.t62 VSS 0.269047f
C10901 a_52635_48695.t63 VSS 0.249659f
C10902 a_52635_48695.n154 VSS 0.855653f
C10903 a_52635_48695.n155 VSS 1.69542f
C10904 a_52635_48695.t71 VSS 0.269047f
C10905 a_52635_48695.t74 VSS 0.249659f
C10906 a_52635_48695.n156 VSS 0.855653f
C10907 a_52635_48695.n157 VSS 1.02404f
C10908 a_52635_48695.t57 VSS 0.095327f
C10909 a_52635_48695.t37 VSS 0.095327f
C10910 a_52635_48695.n158 VSS 0.262987f
C10911 a_52635_48695.t59 VSS 0.095327f
C10912 a_52635_48695.t40 VSS 0.095327f
C10913 a_52635_48695.n159 VSS 0.240154f
C10914 a_52635_48695.n160 VSS 0.662406f
C10915 a_52635_48695.n161 VSS 1.57198f
C10916 a_52635_48695.n162 VSS 1.80922f
C10917 a_52635_48695.n163 VSS 5.54919f
C10918 a_52635_48695.n164 VSS 4.03603f
C10919 a_52635_48695.n165 VSS 0.794975f
C10920 a_52635_48695.t77 VSS 0.095327f
C10921 a_52635_48695.t31 VSS 0.095327f
C10922 a_52635_48695.n166 VSS 0.349727f
C10923 a_52635_48695.n167 VSS 1.1884f
C10924 a_52635_48695.t7 VSS 0.095327f
C10925 a_52635_48695.t11 VSS 0.095327f
C10926 a_52635_48695.n168 VSS 0.349727f
C10927 a_52635_48695.n169 VSS 1.21985f
C10928 a_52635_48695.t14 VSS 0.095327f
C10929 a_52635_48695.t53 VSS 0.095327f
C10930 a_52635_48695.n170 VSS 0.349727f
C10931 a_52635_48695.n171 VSS 1.21988f
C10932 a_52635_48695.t41 VSS 0.095327f
C10933 a_52635_48695.t18 VSS 0.095327f
C10934 a_52635_48695.n172 VSS 0.349727f
C10935 a_52635_48695.n173 VSS 0.750098f
C10936 a_52635_48695.n174 VSS 4.07689f
C10937 a_52635_48695.t73 VSS 0.095327f
C10938 a_52635_48695.t23 VSS 0.095327f
C10939 a_52635_48695.n175 VSS 0.522376f
C10940 a_52635_48695.t72 VSS 0.095327f
C10941 a_52635_48695.t52 VSS 0.095327f
C10942 a_52635_48695.n176 VSS 0.348711f
C10943 a_52635_48695.t80 VSS 0.095327f
C10944 a_52635_48695.t32 VSS 0.095327f
C10945 a_52635_48695.n177 VSS 0.348711f
C10946 a_52635_48695.t8 VSS 0.095327f
C10947 a_52635_48695.t85 VSS 0.095327f
C10948 a_52635_48695.n178 VSS 0.348711f
C10949 a_52635_48695.n179 VSS 0.794898f
C10950 a_52635_48695.t67 VSS 0.095327f
C10951 a_52635_48695.t27 VSS 0.095327f
C10952 a_52635_48695.n180 VSS 0.348711f
C10953 a_52635_48695.t86 VSS 0.095327f
C10954 a_52635_48695.t4 VSS 0.095327f
C10955 a_52635_48695.n181 VSS 0.348711f
C10956 a_52635_48695.t5 VSS 0.095327f
C10957 a_52635_48695.t51 VSS 0.095327f
C10958 a_52635_48695.n182 VSS 0.348711f
C10959 a_52635_48695.t33 VSS 0.095327f
C10960 a_52635_48695.t10 VSS 0.095327f
C10961 a_52635_48695.n183 VSS 0.348711f
C10962 a_52635_48695.n184 VSS 3.92896f
C10963 a_52635_48695.n185 VSS 3.8188f
C10964 a_52635_48695.t79 VSS 0.269047f
C10965 a_52635_48695.t0 VSS 0.249659f
C10966 a_52635_48695.n186 VSS 0.855653f
C10967 a_52635_48695.n187 VSS 1.02404f
C10968 a_52635_48695.t64 VSS 0.095327f
C10969 a_52635_48695.t44 VSS 0.095327f
C10970 a_52635_48695.n188 VSS 0.262987f
C10971 a_52635_48695.t70 VSS 0.095327f
C10972 a_52635_48695.t49 VSS 0.095327f
C10973 a_52635_48695.n189 VSS 0.240154f
C10974 a_52635_48695.n190 VSS 0.662406f
C10975 a_52635_48695.n191 VSS 1.57198f
C10976 a_52635_48695.n192 VSS 1.80922f
C10977 a_52635_48695.n193 VSS 3.37931f
C10978 a_52635_48695.n194 VSS 4.6906f
C10979 a_52635_48695.n195 VSS 0.794975f
C10980 a_52635_48695.n196 VSS 1.1884f
C10981 a_52635_48695.n197 VSS 0.349727f
C10982 a_52635_48695.t87 VSS 0.095327f
C10983 a_35922_19591.n0 VSS 4.07049f
C10984 a_35922_19591.n1 VSS 0.727355f
C10985 a_35922_19591.n2 VSS 0.275511f
C10986 a_35922_19591.n3 VSS 0.95902f
C10987 a_35922_19591.t139 VSS 0.352198f
C10988 a_35922_19591.n4 VSS 0.743998f
C10989 a_35922_19591.n5 VSS 0.682821f
C10990 a_35922_19591.n6 VSS 0.367906f
C10991 a_35922_19591.n7 VSS 0.682821f
C10992 a_35922_19591.n8 VSS 0.743998f
C10993 a_35922_19591.n9 VSS 0.278311f
C10994 a_35922_19591.n10 VSS 0.952664f
C10995 a_35922_19591.n11 VSS 0.70044f
C10996 a_35922_19591.n12 VSS 0.952664f
C10997 a_35922_19591.n13 VSS 0.70044f
C10998 a_35922_19591.n14 VSS 0.424549f
C10999 a_35922_19591.n15 VSS 0.507406f
C11000 a_35922_19591.n16 VSS 0.531489f
C11001 a_35922_19591.n17 VSS 0.424549f
C11002 a_35922_19591.n18 VSS 0.507406f
C11003 a_35922_19591.n19 VSS 0.278537f
C11004 a_35922_19591.n20 VSS 0.531489f
C11005 a_35922_19591.n21 VSS 0.209745f
C11006 a_35922_19591.n22 VSS 0.209881f
C11007 a_35922_19591.n23 VSS 0.531489f
C11008 a_35922_19591.n24 VSS 0.271806f
C11009 a_35922_19591.n25 VSS 0.278537f
C11010 a_35922_19591.n26 VSS 0.209745f
C11011 a_35922_19591.n27 VSS 0.278537f
C11012 a_35922_19591.n28 VSS 0.209881f
C11013 a_35922_19591.n29 VSS 0.531489f
C11014 a_35922_19591.n30 VSS 0.271806f
C11015 a_35922_19591.n31 VSS 1.84527f
C11016 a_35922_19591.n32 VSS 0.670274f
C11017 a_35922_19591.n33 VSS 0.605009f
C11018 a_35922_19591.n34 VSS 1.84527f
C11019 a_35922_19591.n35 VSS 0.687543f
C11020 a_35922_19591.n36 VSS 0.749141f
C11021 a_35922_19591.n37 VSS 0.434127f
C11022 a_35922_19591.n38 VSS 0.605009f
C11023 a_35922_19591.n39 VSS 1.84527f
C11024 a_35922_19591.n40 VSS 0.670274f
C11025 a_35922_19591.n41 VSS 0.473019f
C11026 a_35922_19591.n42 VSS 0.749141f
C11027 a_35922_19591.n43 VSS 1.84527f
C11028 a_35922_19591.n44 VSS 0.687543f
C11029 a_35922_19591.n45 VSS 0.9613f
C11030 a_35922_19591.n46 VSS 0.742498f
C11031 a_35922_19591.n47 VSS 0.622834f
C11032 a_35922_19591.n48 VSS 1.8766f
C11033 a_35922_19591.n49 VSS 0.654383f
C11034 a_35922_19591.n50 VSS 1.88001f
C11035 a_35922_19591.n51 VSS 0.69152f
C11036 a_35922_19591.n52 VSS 0.441628f
C11037 a_35922_19591.n53 VSS 0.622828f
C11038 a_35922_19591.n54 VSS 1.8766f
C11039 a_35922_19591.n55 VSS 0.654382f
C11040 a_35922_19591.n56 VSS 1.88001f
C11041 a_35922_19591.n57 VSS 0.691539f
C11042 a_35922_19591.n58 VSS 0.742519f
C11043 a_35922_19591.n59 VSS 0.226402f
C11044 a_35922_19591.n60 VSS 0.110721f
C11045 a_35922_19591.n61 VSS 0.226784f
C11046 a_35922_19591.n62 VSS 0.226784f
C11047 a_35922_19591.n63 VSS 4.32896f
C11048 a_35922_19591.n64 VSS 1.31313f
C11049 a_35922_19591.n65 VSS 0.458534f
C11050 a_35922_19591.n66 VSS 1.31313f
C11051 a_35922_19591.n67 VSS 0.459143f
C11052 a_35922_19591.n68 VSS 1.31313f
C11053 a_35922_19591.n69 VSS 0.458534f
C11054 a_35922_19591.n70 VSS 1.31313f
C11055 a_35922_19591.n71 VSS 0.459143f
C11056 a_35922_19591.n72 VSS 1.78373f
C11057 a_35922_19591.n73 VSS 0.965859f
C11058 a_35922_19591.n74 VSS 1.78373f
C11059 a_35922_19591.n75 VSS 0.965859f
C11060 a_35922_19591.n76 VSS 1.37036f
C11061 a_35922_19591.n77 VSS 0.486448f
C11062 a_35922_19591.n78 VSS 1.37036f
C11063 a_35922_19591.n79 VSS 0.452424f
C11064 a_35922_19591.n80 VSS 1.37036f
C11065 a_35922_19591.n81 VSS 0.486508f
C11066 a_35922_19591.n82 VSS 1.37036f
C11067 a_35922_19591.n83 VSS 0.452437f
C11068 a_35922_19591.n84 VSS 1.80279f
C11069 a_35922_19591.n85 VSS 0.982133f
C11070 a_35922_19591.n86 VSS 1.80279f
C11071 a_35922_19591.n87 VSS 0.982133f
C11072 a_35922_19591.n88 VSS 0.473019f
C11073 a_35922_19591.n89 VSS 0.785866f
C11074 a_35922_19591.n90 VSS 1.78304f
C11075 a_35922_19591.n91 VSS 1.78304f
C11076 a_35922_19591.n92 VSS 0.785866f
C11077 a_35922_19591.n93 VSS 1.01659f
C11078 a_35922_19591.n94 VSS 1.79407f
C11079 a_35922_19591.n95 VSS 0.787626f
C11080 a_35922_19591.n96 VSS 0.46348f
C11081 a_35922_19591.n97 VSS 0.983076f
C11082 a_35922_19591.n98 VSS 0.787638f
C11083 a_35922_19591.n99 VSS 1.79407f
C11084 a_35922_19591.t188 VSS 0.377115f
C11085 a_35922_19591.n100 VSS 0.349439f
C11086 a_35922_19591.n101 VSS 0.349439f
C11087 a_35922_19591.t18 VSS 0.377115f
C11088 a_35922_19591.n102 VSS 0.041059f
C11089 a_35922_19591.n103 VSS 0.145445f
C11090 a_35922_19591.n104 VSS 0.041059f
C11091 a_35922_19591.n105 VSS 0.145445f
C11092 a_35922_19591.n106 VSS 0.145445f
C11093 a_35922_19591.n107 VSS 0.145445f
C11094 a_35922_19591.n108 VSS 0.179036f
C11095 a_35922_19591.n109 VSS 0.254443f
C11096 a_35922_19591.n110 VSS 0.145445f
C11097 a_35922_19591.n111 VSS 0.145445f
C11098 a_35922_19591.n112 VSS 0.145445f
C11099 a_35922_19591.n113 VSS 0.024141f
C11100 a_35922_19591.n114 VSS 0.040689f
C11101 a_35922_19591.n115 VSS 0.145445f
C11102 a_35922_19591.n116 VSS 0.041059f
C11103 a_35922_19591.n117 VSS 0.040689f
C11104 a_35922_19591.n118 VSS 0.145445f
C11105 a_35922_19591.n119 VSS 0.145445f
C11106 a_35922_19591.n120 VSS 0.163374f
C11107 a_35922_19591.n121 VSS 0.285649f
C11108 a_35922_19591.n122 VSS 0.024141f
C11109 a_35922_19591.n123 VSS 0.041059f
C11110 a_35922_19591.n124 VSS 0.145445f
C11111 a_35922_19591.n125 VSS 0.041059f
C11112 a_35922_19591.n126 VSS 0.145445f
C11113 a_35922_19591.t2 VSS 0.240828f
C11114 a_35922_19591.n127 VSS 2.45557f
C11115 a_35922_19591.n128 VSS 2.42356f
C11116 a_35922_19591.t69 VSS 0.341209f
C11117 a_35922_19591.t140 VSS 0.341209f
C11118 a_35922_19591.t54 VSS 0.341209f
C11119 a_35922_19591.t88 VSS 0.341209f
C11120 a_35922_19591.n129 VSS 0.04322f
C11121 a_35922_19591.t65 VSS 0.341209f
C11122 a_35922_19591.n130 VSS 0.04322f
C11123 a_35922_19591.t157 VSS 0.341209f
C11124 a_35922_19591.n131 VSS 0.177876f
C11125 a_35922_19591.t64 VSS 0.348542f
C11126 a_35922_19591.n132 VSS 0.25446f
C11127 a_35922_19591.n133 VSS 0.156818f
C11128 a_35922_19591.n134 VSS 0.040689f
C11129 a_35922_19591.n135 VSS 0.024141f
C11130 a_35922_19591.n136 VSS 0.04322f
C11131 a_35922_19591.n137 VSS 0.040689f
C11132 a_35922_19591.n138 VSS 0.024141f
C11133 a_35922_19591.n139 VSS 1.02835f
C11134 a_35922_19591.n140 VSS 0.199552f
C11135 a_35922_19591.n141 VSS 0.040689f
C11136 a_35922_19591.t145 VSS 0.341209f
C11137 a_35922_19591.n142 VSS 0.177876f
C11138 a_35922_19591.t38 VSS 0.348542f
C11139 a_35922_19591.n143 VSS 0.25446f
C11140 a_35922_19591.n144 VSS 0.156818f
C11141 a_35922_19591.n145 VSS 0.04322f
C11142 a_35922_19591.t39 VSS 0.341209f
C11143 a_35922_19591.n146 VSS 0.040689f
C11144 a_35922_19591.n147 VSS 0.04322f
C11145 a_35922_19591.n148 VSS 0.04322f
C11146 a_35922_19591.n149 VSS 0.024141f
C11147 a_35922_19591.t79 VSS 0.341209f
C11148 a_35922_19591.n150 VSS 0.114377f
C11149 a_35922_19591.t91 VSS 0.341209f
C11150 a_35922_19591.n151 VSS 0.276312f
C11151 a_35922_19591.t106 VSS 0.341209f
C11152 a_35922_19591.n152 VSS 0.227193f
C11153 a_35922_19591.t35 VSS 0.341209f
C11154 a_35922_19591.n153 VSS 0.275511f
C11155 a_35922_19591.n154 VSS 0.04322f
C11156 a_35922_19591.n155 VSS 0.051142f
C11157 a_35922_19591.t172 VSS 0.341209f
C11158 a_35922_19591.t10 VSS 0.341209f
C11159 a_35922_19591.n156 VSS 0.051139f
C11160 a_35922_19591.n157 VSS 0.04322f
C11161 a_35922_19591.t136 VSS 0.341209f
C11162 a_35922_19591.t7 VSS 0.341209f
C11163 a_35922_19591.n158 VSS 0.04322f
C11164 a_35922_19591.t184 VSS 0.341209f
C11165 a_35922_19591.t171 VSS 0.341209f
C11166 a_35922_19591.t67 VSS 0.341209f
C11167 a_35922_19591.t135 VSS 0.341209f
C11168 a_35922_19591.t189 VSS 0.341209f
C11169 a_35922_19591.t100 VSS 0.341209f
C11170 a_35922_19591.n159 VSS 0.278311f
C11171 a_35922_19591.t118 VSS 0.341209f
C11172 a_35922_19591.n160 VSS 0.227193f
C11173 a_35922_19591.t53 VSS 0.341209f
C11174 a_35922_19591.t96 VSS 0.341209f
C11175 a_35922_19591.t151 VSS 0.341209f
C11176 a_35922_19591.t164 VSS 0.341209f
C11177 a_35922_19591.t6 VSS 0.341209f
C11178 a_35922_19591.t115 VSS 0.341209f
C11179 a_35922_19591.t162 VSS 0.341209f
C11180 a_35922_19591.t156 VSS 0.341209f
C11181 a_35922_19591.t56 VSS 0.341209f
C11182 a_35922_19591.n161 VSS 0.278311f
C11183 a_35922_19591.t97 VSS 0.341209f
C11184 a_35922_19591.n162 VSS 0.227193f
C11185 a_35922_19591.t23 VSS 0.341209f
C11186 a_35922_19591.t73 VSS 0.341209f
C11187 a_35922_19591.t95 VSS 0.341209f
C11188 a_35922_19591.t150 VSS 0.350512f
C11189 a_35922_19591.t153 VSS 0.341209f
C11190 a_35922_19591.n163 VSS 3.64752f
C11191 a_35922_19591.n164 VSS 0.249586f
C11192 a_35922_19591.n165 VSS 0.04322f
C11193 a_35922_19591.t179 VSS 0.341209f
C11194 a_35922_19591.t83 VSS 0.341209f
C11195 a_35922_19591.n166 VSS 0.159294f
C11196 a_35922_19591.t120 VSS 0.341209f
C11197 a_35922_19591.t168 VSS 0.348659f
C11198 a_35922_19591.n167 VSS 0.041059f
C11199 a_35922_19591.n168 VSS 0.040689f
C11200 a_35922_19591.n169 VSS 0.04322f
C11201 a_35922_19591.n170 VSS 0.024141f
C11202 a_35922_19591.n171 VSS 0.041059f
C11203 a_35922_19591.n172 VSS 0.040689f
C11204 a_35922_19591.n173 VSS 0.04322f
C11205 a_35922_19591.n174 VSS 0.024141f
C11206 a_35922_19591.n175 VSS 0.074175f
C11207 a_35922_19591.n176 VSS 0.114068f
C11208 a_35922_19591.t192 VSS 0.341209f
C11209 a_35922_19591.n177 VSS 0.275511f
C11210 a_35922_19591.t90 VSS 0.341209f
C11211 a_35922_19591.n178 VSS 0.227193f
C11212 a_35922_19591.t41 VSS 0.341209f
C11213 a_35922_19591.n179 VSS 0.276312f
C11214 a_35922_19591.n180 VSS 0.114377f
C11215 a_35922_19591.n181 VSS 0.199552f
C11216 a_35922_19591.n182 VSS 0.024141f
C11217 a_35922_19591.n183 VSS 0.041059f
C11218 a_35922_19591.n184 VSS 0.040689f
C11219 a_35922_19591.n185 VSS 0.04322f
C11220 a_35922_19591.n186 VSS 0.024141f
C11221 a_35922_19591.n187 VSS 0.041059f
C11222 a_35922_19591.n188 VSS 0.040689f
C11223 a_35922_19591.n189 VSS 0.04322f
C11224 a_35922_19591.n190 VSS 0.024141f
C11225 a_35922_19591.n191 VSS 0.04322f
C11226 a_35922_19591.n192 VSS 0.041059f
C11227 a_35922_19591.n193 VSS 0.040689f
C11228 a_35922_19591.t48 VSS 0.341209f
C11229 a_35922_19591.n194 VSS 0.164008f
C11230 a_35922_19591.n195 VSS 0.285749f
C11231 a_35922_19591.n196 VSS 0.041059f
C11232 a_35922_19591.n197 VSS 0.040689f
C11233 a_35922_19591.n198 VSS 0.04322f
C11234 a_35922_19591.n199 VSS 0.024141f
C11235 a_35922_19591.n200 VSS 0.04322f
C11236 a_35922_19591.n201 VSS 0.041059f
C11237 a_35922_19591.t121 VSS 0.341209f
C11238 a_35922_19591.n202 VSS 0.024141f
C11239 a_35922_19591.n203 VSS 0.04322f
C11240 a_35922_19591.n204 VSS 0.04322f
C11241 a_35922_19591.t22 VSS 0.341209f
C11242 a_35922_19591.n205 VSS 0.114068f
C11243 a_35922_19591.n206 VSS 0.074175f
C11244 a_35922_19591.n207 VSS 0.249586f
C11245 a_35922_19591.n208 VSS 3.64752f
C11246 a_35922_19591.t142 VSS 0.341209f
C11247 a_35922_19591.t20 VSS 0.341209f
C11248 a_35922_19591.t72 VSS 0.341209f
C11249 a_35922_19591.t114 VSS 0.341209f
C11250 a_35922_19591.n209 VSS 0.278311f
C11251 a_35922_19591.t133 VSS 0.341209f
C11252 a_35922_19591.n210 VSS 0.227193f
C11253 a_35922_19591.t63 VSS 0.341209f
C11254 a_35922_19591.t110 VSS 0.341209f
C11255 a_35922_19591.t159 VSS 0.341209f
C11256 a_35922_19591.t126 VSS 0.341209f
C11257 a_35922_19591.t175 VSS 0.341209f
C11258 a_35922_19591.n211 VSS 0.356155f
C11259 a_35922_19591.t166 VSS 0.341209f
C11260 a_35922_19591.t161 VSS 0.341209f
C11261 a_35922_19591.t78 VSS 0.341209f
C11262 a_35922_19591.t107 VSS 0.341209f
C11263 a_35922_19591.t155 VSS 0.350512f
C11264 a_35922_19591.t40 VSS 0.341209f
C11265 a_35922_19591.n212 VSS 0.278537f
C11266 a_35922_19591.t112 VSS 0.341209f
C11267 a_35922_19591.n213 VSS 0.227193f
C11268 a_35922_19591.t68 VSS 0.341209f
C11269 a_35922_19591.t27 VSS 0.341209f
C11270 a_35922_19591.t177 VSS 0.341209f
C11271 a_35922_19591.t186 VSS 0.341209f
C11272 a_35922_19591.n214 VSS 2.42356f
C11273 a_35922_19591.n215 VSS 2.42356f
C11274 a_35922_19591.t131 VSS 0.341209f
C11275 a_35922_19591.t45 VSS 0.341209f
C11276 a_35922_19591.t147 VSS 0.341209f
C11277 a_35922_19591.t44 VSS 0.341209f
C11278 a_35922_19591.t80 VSS 0.341209f
C11279 a_35922_19591.t143 VSS 0.341209f
C11280 a_35922_19591.t74 VSS 0.341209f
C11281 a_35922_19591.t125 VSS 0.341209f
C11282 a_35922_19591.t174 VSS 0.341209f
C11283 a_35922_19591.t15 VSS 0.341209f
C11284 a_35922_19591.t13 VSS 0.341209f
C11285 a_35922_19591.t62 VSS 0.341209f
C11286 a_35922_19591.t167 VSS 0.341209f
C11287 a_35922_19591.t119 VSS 0.341209f
C11288 a_35922_19591.t154 VSS 0.341209f
C11289 a_35922_19591.t103 VSS 0.341209f
C11290 a_35922_19591.t89 VSS 0.341209f
C11291 a_35922_19591.t30 VSS 0.341209f
C11292 a_35922_19591.t144 VSS 0.341209f
C11293 a_35922_19591.t31 VSS 0.341209f
C11294 a_35922_19591.t77 VSS 0.341209f
C11295 a_35922_19591.t98 VSS 0.341209f
C11296 a_35922_19591.t25 VSS 0.341209f
C11297 a_35922_19591.t12 VSS 0.341209f
C11298 a_35922_19591.t117 VSS 0.341209f
C11299 a_35922_19591.t165 VSS 0.341209f
C11300 a_35922_19591.t190 VSS 0.341209f
C11301 a_35922_19591.t87 VSS 0.341209f
C11302 a_35922_19591.t182 VSS 0.341209f
C11303 a_35922_19591.t170 VSS 0.341209f
C11304 a_35922_19591.t82 VSS 0.341209f
C11305 a_35922_19591.t116 VSS 0.341209f
C11306 a_35922_19591.t163 VSS 0.341209f
C11307 a_35922_19591.t33 VSS 0.341209f
C11308 a_35922_19591.t178 VSS 0.341209f
C11309 a_35922_19591.t187 VSS 0.341209f
C11310 a_35922_19591.t134 VSS 0.341209f
C11311 a_35922_19591.t37 VSS 0.341209f
C11312 a_35922_19591.n216 VSS 3.78794f
C11313 a_35922_19591.t108 VSS 0.341209f
C11314 a_35922_19591.t70 VSS 0.341209f
C11315 a_35922_19591.t9 VSS 0.341209f
C11316 a_35922_19591.t137 VSS 0.341209f
C11317 a_35922_19591.t8 VSS 0.341209f
C11318 a_35922_19591.t123 VSS 0.341209f
C11319 a_35922_19591.t57 VSS 0.341209f
C11320 a_35922_19591.t181 VSS 0.341209f
C11321 a_35922_19591.t169 VSS 0.341209f
C11322 a_35922_19591.t19 VSS 0.341209f
C11323 a_35922_19591.t160 VSS 0.341209f
C11324 a_35922_19591.t105 VSS 0.341209f
C11325 a_35922_19591.t34 VSS 0.341209f
C11326 a_35922_19591.t75 VSS 0.341209f
C11327 a_35922_19591.t101 VSS 0.341209f
C11328 a_35922_19591.t152 VSS 0.341209f
C11329 a_35922_19591.t158 VSS 0.341209f
C11330 a_35922_19591.n217 VSS 3.78794f
C11331 a_35922_19591.t50 VSS 0.341209f
C11332 a_35922_19591.t21 VSS 0.341209f
C11333 a_35922_19591.t130 VSS 0.341209f
C11334 a_35922_19591.t28 VSS 0.341209f
C11335 a_35922_19591.t81 VSS 0.341209f
C11336 a_35922_19591.t148 VSS 0.341209f
C11337 a_35922_19591.t47 VSS 0.341209f
C11338 a_35922_19591.t49 VSS 0.341209f
C11339 a_35922_19591.t113 VSS 0.341209f
C11340 a_35922_19591.t42 VSS 0.341209f
C11341 a_35922_19591.t93 VSS 0.341209f
C11342 a_35922_19591.t180 VSS 0.341209f
C11343 a_35922_19591.t55 VSS 0.341209f
C11344 a_35922_19591.t141 VSS 0.341209f
C11345 a_35922_19591.t17 VSS 0.341209f
C11346 a_35922_19591.t193 VSS 0.341209f
C11347 a_35922_19591.t92 VSS 0.341209f
C11348 a_35922_19591.t11 VSS 0.341209f
C11349 a_35922_19591.t185 VSS 0.341209f
C11350 a_35922_19591.t85 VSS 0.341209f
C11351 a_35922_19591.t127 VSS 0.341209f
C11352 a_35922_19591.t176 VSS 0.341209f
C11353 a_35922_19591.n218 VSS 2.42356f
C11354 a_35922_19591.n219 VSS 2.03211f
C11355 a_35922_19591.n220 VSS 0.434127f
C11356 a_35922_19591.t191 VSS 0.341209f
C11357 a_35922_19591.t128 VSS 0.341209f
C11358 a_35922_19591.t59 VSS 0.341209f
C11359 a_35922_19591.t183 VSS 0.341209f
C11360 a_35922_19591.t84 VSS 0.341209f
C11361 a_35922_19591.t122 VSS 0.341209f
C11362 a_35922_19591.t173 VSS 0.341209f
C11363 a_35922_19591.t76 VSS 0.341209f
C11364 a_35922_19591.t138 VSS 0.341209f
C11365 a_35922_19591.t52 VSS 0.341209f
C11366 a_35922_19591.t26 VSS 0.341209f
C11367 a_35922_19591.n221 VSS 2.26597f
C11368 a_35922_19591.n222 VSS 2.92955f
C11369 a_35922_19591.n223 VSS 2.13722f
C11370 a_35922_19591.n224 VSS 0.367115f
C11371 a_35922_19591.n225 VSS 0.199552f
C11372 a_35922_19591.n226 VSS 0.114377f
C11373 a_35922_19591.t111 VSS 0.341209f
C11374 a_35922_19591.n227 VSS 0.276312f
C11375 a_35922_19591.t129 VSS 0.341209f
C11376 a_35922_19591.n228 VSS 0.227193f
C11377 a_35922_19591.t60 VSS 0.341209f
C11378 a_35922_19591.t16 VSS 0.341209f
C11379 a_35922_19591.t46 VSS 0.341209f
C11380 a_35922_19591.t146 VSS 0.341209f
C11381 a_35922_19591.t43 VSS 0.341209f
C11382 a_35922_19591.t32 VSS 0.341209f
C11383 a_35922_19591.t66 VSS 0.341209f
C11384 a_35922_19591.t109 VSS 0.341209f
C11385 a_35922_19591.t36 VSS 0.341209f
C11386 a_35922_19591.t14 VSS 0.348659f
C11387 a_35922_19591.t94 VSS 0.341209f
C11388 a_35922_19591.t24 VSS 0.341209f
C11389 a_35922_19591.n229 VSS 2.13722f
C11390 a_35922_19591.n230 VSS 8.488879f
C11391 a_35922_19591.t1 VSS 0.058657f
C11392 a_35922_19591.t0 VSS 0.222881f
C11393 a_35922_19591.n231 VSS 0.288911f
C11394 a_35922_19591.t124 VSS 0.248352f
C11395 a_35922_19591.n232 VSS 0.280777f
C11396 a_35922_19591.t99 VSS 0.264051f
C11397 a_35922_19591.t58 VSS 0.248352f
C11398 a_35922_19591.n233 VSS 0.417235f
C11399 a_35922_19591.t132 VSS 0.251241f
C11400 a_35922_19591.t104 VSS 0.264023f
C11401 a_35922_19591.t61 VSS 0.248352f
C11402 a_35922_19591.n234 VSS 0.416873f
C11403 a_35922_19591.t71 VSS 0.251248f
C11404 a_35922_19591.t51 VSS 0.264262f
C11405 a_35922_19591.t149 VSS 0.248352f
C11406 a_35922_19591.n235 VSS 0.419944f
C11407 a_35922_19591.t102 VSS 0.251248f
C11408 a_35922_19591.t86 VSS 0.264234f
C11409 a_35922_19591.t29 VSS 0.248352f
C11410 a_35922_19591.n236 VSS 0.419583f
C11411 a_35922_19591.n237 VSS 10.4498f
C11412 a_35922_19591.t3 VSS 0.208804f
C11413 a_35922_19591.t4 VSS 0.235371f
C11414 a_35922_19591.n238 VSS 0.734704f
C11415 a_35922_19591.n239 VSS 3.23651f
C11416 a_35922_19591.n240 VSS 0.873591f
C11417 a_35922_19591.t5 VSS 0.182449f
C11418 a_71281_n8397.n0 VSS 1.83357f
C11419 a_71281_n8397.n1 VSS 5.784431f
C11420 a_71281_n8397.t41 VSS 0.033548f
C11421 a_71281_n8397.t45 VSS 0.159066f
C11422 a_71281_n8397.n2 VSS 0.051472f
C11423 a_71281_n8397.n3 VSS 0.047376f
C11424 a_71281_n8397.n4 VSS 0.43613f
C11425 a_71281_n8397.t269 VSS 0.418638f
C11426 a_71281_n8397.n5 VSS 0.419773f
C11427 a_71281_n8397.t234 VSS 0.382252f
C11428 a_71281_n8397.n6 VSS 0.43064f
C11429 a_71281_n8397.n7 VSS 0.047376f
C11430 a_71281_n8397.t81 VSS 0.421756f
C11431 a_71281_n8397.t144 VSS 0.382162f
C11432 a_71281_n8397.n8 VSS 0.43613f
C11433 a_71281_n8397.n9 VSS 0.042199f
C11434 a_71281_n8397.n10 VSS 0.14932f
C11435 a_71281_n8397.t311 VSS 0.33632f
C11436 a_71281_n8397.n11 VSS 0.14932f
C11437 a_71281_n8397.n12 VSS 0.042199f
C11438 a_71281_n8397.n13 VSS 0.01957f
C11439 a_71281_n8397.n14 VSS 0.533769f
C11440 a_71281_n8397.n15 VSS 0.267172f
C11441 a_71281_n8397.n16 VSS 0.047376f
C11442 a_71281_n8397.n17 VSS 0.43613f
C11443 a_71281_n8397.t335 VSS 0.421781f
C11444 a_71281_n8397.n18 VSS 0.43064f
C11445 a_71281_n8397.t300 VSS 0.382252f
C11446 a_71281_n8397.n19 VSS 0.43064f
C11447 a_71281_n8397.n20 VSS 0.047376f
C11448 a_71281_n8397.t154 VSS 0.421756f
C11449 a_71281_n8397.t216 VSS 0.382162f
C11450 a_71281_n8397.n21 VSS 0.43613f
C11451 a_71281_n8397.n22 VSS 0.01957f
C11452 a_71281_n8397.n23 VSS 0.042199f
C11453 a_71281_n8397.n24 VSS 0.14932f
C11454 a_71281_n8397.t127 VSS 0.33632f
C11455 a_71281_n8397.n25 VSS 0.14932f
C11456 a_71281_n8397.n26 VSS 0.042199f
C11457 a_71281_n8397.n27 VSS 0.01957f
C11458 a_71281_n8397.n28 VSS 0.267172f
C11459 a_71281_n8397.n29 VSS 0.267467f
C11460 a_71281_n8397.n30 VSS 0.047376f
C11461 a_71281_n8397.n31 VSS 0.43613f
C11462 a_71281_n8397.t328 VSS 0.421781f
C11463 a_71281_n8397.n32 VSS 0.43064f
C11464 a_71281_n8397.t292 VSS 0.382252f
C11465 a_71281_n8397.n33 VSS 0.43064f
C11466 a_71281_n8397.n34 VSS 0.047376f
C11467 a_71281_n8397.t151 VSS 0.421756f
C11468 a_71281_n8397.t212 VSS 0.382162f
C11469 a_71281_n8397.n35 VSS 0.43613f
C11470 a_71281_n8397.n36 VSS 0.01957f
C11471 a_71281_n8397.n37 VSS 0.042199f
C11472 a_71281_n8397.n38 VSS 0.14932f
C11473 a_71281_n8397.t119 VSS 0.33632f
C11474 a_71281_n8397.n39 VSS 0.14932f
C11475 a_71281_n8397.n40 VSS 0.042199f
C11476 a_71281_n8397.n41 VSS 0.01957f
C11477 a_71281_n8397.n42 VSS 0.267467f
C11478 a_71281_n8397.n43 VSS 0.268058f
C11479 a_71281_n8397.n44 VSS 0.047376f
C11480 a_71281_n8397.n45 VSS 0.43613f
C11481 a_71281_n8397.t141 VSS 0.421781f
C11482 a_71281_n8397.n46 VSS 0.43064f
C11483 a_71281_n8397.t109 VSS 0.382252f
C11484 a_71281_n8397.n47 VSS 0.43064f
C11485 a_71281_n8397.n48 VSS 0.047376f
C11486 a_71281_n8397.t222 VSS 0.421756f
C11487 a_71281_n8397.t278 VSS 0.382162f
C11488 a_71281_n8397.n49 VSS 0.43613f
C11489 a_71281_n8397.n50 VSS 0.01957f
C11490 a_71281_n8397.n51 VSS 0.042199f
C11491 a_71281_n8397.n52 VSS 0.14932f
C11492 a_71281_n8397.t193 VSS 0.33632f
C11493 a_71281_n8397.n53 VSS 0.14932f
C11494 a_71281_n8397.n54 VSS 0.042199f
C11495 a_71281_n8397.n55 VSS 0.01957f
C11496 a_71281_n8397.n56 VSS 0.221362f
C11497 a_71281_n8397.t67 VSS 0.159066f
C11498 a_71281_n8397.t43 VSS 0.033548f
C11499 a_71281_n8397.t11 VSS 0.033548f
C11500 a_71281_n8397.n57 VSS 0.136945f
C11501 a_71281_n8397.n58 VSS 0.382877f
C11502 a_71281_n8397.n59 VSS 0.092801f
C11503 a_71281_n8397.n60 VSS 0.221362f
C11504 a_71281_n8397.n61 VSS 0.047376f
C11505 a_71281_n8397.n62 VSS 0.43613f
C11506 a_71281_n8397.t134 VSS 0.421781f
C11507 a_71281_n8397.n63 VSS 0.43064f
C11508 a_71281_n8397.t66 VSS 0.382252f
C11509 a_71281_n8397.n64 VSS 0.43064f
C11510 a_71281_n8397.n65 VSS 0.047376f
C11511 a_71281_n8397.t214 VSS 0.421756f
C11512 a_71281_n8397.t10 VSS 0.382162f
C11513 a_71281_n8397.n66 VSS 0.43613f
C11514 a_71281_n8397.n67 VSS 0.01957f
C11515 a_71281_n8397.n68 VSS 0.042199f
C11516 a_71281_n8397.n69 VSS 0.14932f
C11517 a_71281_n8397.t42 VSS 0.33632f
C11518 a_71281_n8397.n70 VSS 0.14932f
C11519 a_71281_n8397.n71 VSS 0.042199f
C11520 a_71281_n8397.n72 VSS 0.01957f
C11521 a_71281_n8397.n73 VSS 0.267467f
C11522 a_71281_n8397.n74 VSS 0.267467f
C11523 a_71281_n8397.n75 VSS 0.047376f
C11524 a_71281_n8397.n76 VSS 0.43613f
C11525 a_71281_n8397.t210 VSS 0.421781f
C11526 a_71281_n8397.n77 VSS 0.43064f
C11527 a_71281_n8397.t46 VSS 0.382252f
C11528 a_71281_n8397.n78 VSS 0.43064f
C11529 a_71281_n8397.n79 VSS 0.047376f
C11530 a_71281_n8397.t281 VSS 0.421756f
C11531 a_71281_n8397.t2 VSS 0.382162f
C11532 a_71281_n8397.n80 VSS 0.43613f
C11533 a_71281_n8397.n81 VSS 0.01957f
C11534 a_71281_n8397.n82 VSS 0.042199f
C11535 a_71281_n8397.n83 VSS 0.14932f
C11536 a_71281_n8397.t20 VSS 0.33632f
C11537 a_71281_n8397.n84 VSS 0.14932f
C11538 a_71281_n8397.n85 VSS 0.042199f
C11539 a_71281_n8397.n86 VSS 0.01957f
C11540 a_71281_n8397.n87 VSS 0.221067f
C11541 a_71281_n8397.t47 VSS 0.033548f
C11542 a_71281_n8397.t21 VSS 0.033548f
C11543 a_71281_n8397.n88 VSS 0.136714f
C11544 a_71281_n8397.t3 VSS 0.159292f
C11545 a_71281_n8397.n89 VSS 0.384352f
C11546 a_71281_n8397.n90 VSS 0.092801f
C11547 a_71281_n8397.n91 VSS 0.220771f
C11548 a_71281_n8397.n92 VSS 0.047376f
C11549 a_71281_n8397.n93 VSS 0.43613f
C11550 a_71281_n8397.t184 VSS 0.421781f
C11551 a_71281_n8397.n94 VSS 0.43064f
C11552 a_71281_n8397.t152 VSS 0.382252f
C11553 a_71281_n8397.n95 VSS 0.43064f
C11554 a_71281_n8397.n96 VSS 0.047376f
C11555 a_71281_n8397.t261 VSS 0.421756f
C11556 a_71281_n8397.t310 VSS 0.382162f
C11557 a_71281_n8397.n97 VSS 0.43613f
C11558 a_71281_n8397.n98 VSS 0.01957f
C11559 a_71281_n8397.n99 VSS 0.042199f
C11560 a_71281_n8397.n100 VSS 0.14932f
C11561 a_71281_n8397.t227 VSS 0.33632f
C11562 a_71281_n8397.n101 VSS 0.14932f
C11563 a_71281_n8397.n102 VSS 0.042199f
C11564 a_71281_n8397.n103 VSS 0.01957f
C11565 a_71281_n8397.n104 VSS 0.267172f
C11566 a_71281_n8397.n105 VSS 0.267467f
C11567 a_71281_n8397.n106 VSS 0.047376f
C11568 a_71281_n8397.n107 VSS 0.43613f
C11569 a_71281_n8397.t252 VSS 0.421781f
C11570 a_71281_n8397.n108 VSS 0.43064f
C11571 a_71281_n8397.t224 VSS 0.382252f
C11572 a_71281_n8397.n109 VSS 0.43064f
C11573 a_71281_n8397.n110 VSS 0.047376f
C11574 a_71281_n8397.t326 VSS 0.421756f
C11575 a_71281_n8397.t125 VSS 0.382162f
C11576 a_71281_n8397.n111 VSS 0.43613f
C11577 a_71281_n8397.n112 VSS 0.01957f
C11578 a_71281_n8397.n113 VSS 0.042199f
C11579 a_71281_n8397.n114 VSS 0.14932f
C11580 a_71281_n8397.t295 VSS 0.33632f
C11581 a_71281_n8397.n115 VSS 0.14932f
C11582 a_71281_n8397.n116 VSS 0.042199f
C11583 a_71281_n8397.n117 VSS 0.01957f
C11584 a_71281_n8397.n118 VSS 0.267467f
C11585 a_71281_n8397.n119 VSS 0.268058f
C11586 a_71281_n8397.n120 VSS 0.047376f
C11587 a_71281_n8397.n121 VSS 0.43613f
C11588 a_71281_n8397.t242 VSS 0.421781f
C11589 a_71281_n8397.n122 VSS 0.43064f
C11590 a_71281_n8397.t217 VSS 0.382252f
C11591 a_71281_n8397.n123 VSS 0.43064f
C11592 a_71281_n8397.n124 VSS 0.047376f
C11593 a_71281_n8397.n125 VSS 0.01957f
C11594 a_71281_n8397.t318 VSS 0.421756f
C11595 a_71281_n8397.t118 VSS 0.382162f
C11596 a_71281_n8397.n126 VSS 0.43613f
C11597 a_71281_n8397.n127 VSS 0.042199f
C11598 a_71281_n8397.n128 VSS 0.14932f
C11599 a_71281_n8397.t286 VSS 0.33632f
C11600 a_71281_n8397.n129 VSS 0.14932f
C11601 a_71281_n8397.n130 VSS 0.042199f
C11602 a_71281_n8397.n131 VSS 0.01957f
C11603 a_71281_n8397.n132 VSS 0.268058f
C11604 a_71281_n8397.n133 VSS 0.267467f
C11605 a_71281_n8397.n134 VSS 0.047376f
C11606 a_71281_n8397.n135 VSS 0.43613f
C11607 a_71281_n8397.t309 VSS 0.421781f
C11608 a_71281_n8397.n136 VSS 0.43064f
C11609 a_71281_n8397.t282 VSS 0.382252f
C11610 a_71281_n8397.n137 VSS 0.43064f
C11611 a_71281_n8397.n138 VSS 0.047376f
C11612 a_71281_n8397.n139 VSS 0.01957f
C11613 a_71281_n8397.t131 VSS 0.421756f
C11614 a_71281_n8397.t191 VSS 0.382162f
C11615 a_71281_n8397.n140 VSS 0.43613f
C11616 a_71281_n8397.n141 VSS 0.042199f
C11617 a_71281_n8397.n142 VSS 0.14932f
C11618 a_71281_n8397.t98 VSS 0.33632f
C11619 a_71281_n8397.n143 VSS 0.14932f
C11620 a_71281_n8397.n144 VSS 0.042199f
C11621 a_71281_n8397.n145 VSS 0.01957f
C11622 a_71281_n8397.n146 VSS 0.605274f
C11623 a_71281_n8397.n147 VSS 0.052547f
C11624 a_71281_n8397.n148 VSS 0.047376f
C11625 a_71281_n8397.n149 VSS 0.43613f
C11626 a_71281_n8397.t178 VSS 0.421781f
C11627 a_71281_n8397.n150 VSS 0.43064f
C11628 a_71281_n8397.t113 VSS 0.382252f
C11629 a_71281_n8397.n151 VSS 0.43064f
C11630 a_71281_n8397.n152 VSS 0.047376f
C11631 a_71281_n8397.t264 VSS 0.421756f
C11632 a_71281_n8397.t255 VSS 0.382162f
C11633 a_71281_n8397.n153 VSS 0.43613f
C11634 a_71281_n8397.n154 VSS 0.042199f
C11635 a_71281_n8397.n155 VSS 0.14932f
C11636 a_71281_n8397.t268 VSS 0.33632f
C11637 a_71281_n8397.n156 VSS 0.14932f
C11638 a_71281_n8397.n157 VSS 0.042199f
C11639 a_71281_n8397.n158 VSS 0.01957f
C11640 a_71281_n8397.n159 VSS 0.542742f
C11641 a_71281_n8397.n160 VSS 0.268058f
C11642 a_71281_n8397.n161 VSS 0.047376f
C11643 a_71281_n8397.n162 VSS 0.43613f
C11644 a_71281_n8397.t111 VSS 0.421781f
C11645 a_71281_n8397.n163 VSS 0.43064f
C11646 a_71281_n8397.t298 VSS 0.382252f
C11647 a_71281_n8397.n164 VSS 0.43064f
C11648 a_71281_n8397.n165 VSS 0.047376f
C11649 a_71281_n8397.t200 VSS 0.421756f
C11650 a_71281_n8397.t187 VSS 0.382162f
C11651 a_71281_n8397.n166 VSS 0.43613f
C11652 a_71281_n8397.n167 VSS 0.01957f
C11653 a_71281_n8397.n168 VSS 0.042199f
C11654 a_71281_n8397.n169 VSS 0.14932f
C11655 a_71281_n8397.t205 VSS 0.33632f
C11656 a_71281_n8397.n170 VSS 0.14932f
C11657 a_71281_n8397.n171 VSS 0.042199f
C11658 a_71281_n8397.n172 VSS 0.01957f
C11659 a_71281_n8397.n173 VSS 0.268058f
C11660 a_71281_n8397.n174 VSS 0.267467f
C11661 a_71281_n8397.n175 VSS 0.047376f
C11662 a_71281_n8397.n176 VSS 0.43613f
C11663 a_71281_n8397.t236 VSS 0.421781f
C11664 a_71281_n8397.n177 VSS 0.43064f
C11665 a_71281_n8397.t169 VSS 0.382252f
C11666 a_71281_n8397.n178 VSS 0.43064f
C11667 a_71281_n8397.n179 VSS 0.047376f
C11668 a_71281_n8397.n180 VSS 0.01957f
C11669 a_71281_n8397.t319 VSS 0.421756f
C11670 a_71281_n8397.t307 VSS 0.382162f
C11671 a_71281_n8397.n181 VSS 0.43613f
C11672 a_71281_n8397.n182 VSS 0.042199f
C11673 a_71281_n8397.n183 VSS 0.14932f
C11674 a_71281_n8397.t324 VSS 0.33632f
C11675 a_71281_n8397.n184 VSS 0.14932f
C11676 a_71281_n8397.n185 VSS 0.042199f
C11677 a_71281_n8397.n186 VSS 0.01957f
C11678 a_71281_n8397.n187 VSS 0.267467f
C11679 a_71281_n8397.n188 VSS 0.267172f
C11680 a_71281_n8397.n189 VSS 0.047376f
C11681 a_71281_n8397.n190 VSS 0.43613f
C11682 a_71281_n8397.t164 VSS 0.421781f
C11683 a_71281_n8397.n191 VSS 0.43064f
C11684 a_71281_n8397.t96 VSS 0.382252f
C11685 a_71281_n8397.n192 VSS 0.43064f
C11686 a_71281_n8397.n193 VSS 0.047376f
C11687 a_71281_n8397.n194 VSS 0.01957f
C11688 a_71281_n8397.t253 VSS 0.421756f
C11689 a_71281_n8397.t240 VSS 0.382162f
C11690 a_71281_n8397.n195 VSS 0.43613f
C11691 a_71281_n8397.n196 VSS 0.042199f
C11692 a_71281_n8397.n197 VSS 0.14932f
C11693 a_71281_n8397.t259 VSS 0.33632f
C11694 a_71281_n8397.n198 VSS 0.14932f
C11695 a_71281_n8397.n199 VSS 0.042199f
C11696 a_71281_n8397.n200 VSS 0.01957f
C11697 a_71281_n8397.n201 VSS 0.220771f
C11698 a_71281_n8397.t65 VSS 0.033548f
C11699 a_71281_n8397.t13 VSS 0.033548f
C11700 a_71281_n8397.n202 VSS 0.136714f
C11701 a_71281_n8397.t17 VSS 0.159292f
C11702 a_71281_n8397.n203 VSS 0.384352f
C11703 a_71281_n8397.n204 VSS 0.092801f
C11704 a_71281_n8397.n205 VSS 0.221067f
C11705 a_71281_n8397.n206 VSS 0.047376f
C11706 a_71281_n8397.n207 VSS 0.43613f
C11707 a_71281_n8397.t177 VSS 0.421781f
C11708 a_71281_n8397.n208 VSS 0.43064f
C11709 a_71281_n8397.t64 VSS 0.382252f
C11710 a_71281_n8397.n209 VSS 0.43064f
C11711 a_71281_n8397.n210 VSS 0.047376f
C11712 a_71281_n8397.n211 VSS 0.01957f
C11713 a_71281_n8397.t262 VSS 0.421756f
C11714 a_71281_n8397.t16 VSS 0.382162f
C11715 a_71281_n8397.n212 VSS 0.43613f
C11716 a_71281_n8397.n213 VSS 0.042199f
C11717 a_71281_n8397.n214 VSS 0.14932f
C11718 a_71281_n8397.t12 VSS 0.33632f
C11719 a_71281_n8397.n215 VSS 0.14932f
C11720 a_71281_n8397.n216 VSS 0.042199f
C11721 a_71281_n8397.n217 VSS 0.01957f
C11722 a_71281_n8397.n218 VSS 0.267467f
C11723 a_71281_n8397.n219 VSS 0.267467f
C11724 a_71281_n8397.n220 VSS 0.047376f
C11725 a_71281_n8397.n221 VSS 0.43613f
C11726 a_71281_n8397.t103 VSS 0.421781f
C11727 a_71281_n8397.n222 VSS 0.43064f
C11728 a_71281_n8397.t6 VSS 0.382252f
C11729 a_71281_n8397.n223 VSS 0.43064f
C11730 a_71281_n8397.n224 VSS 0.047376f
C11731 a_71281_n8397.n225 VSS 0.01957f
C11732 a_71281_n8397.t197 VSS 0.421756f
C11733 a_71281_n8397.t38 VSS 0.382162f
C11734 a_71281_n8397.n226 VSS 0.43613f
C11735 a_71281_n8397.n227 VSS 0.042199f
C11736 a_71281_n8397.n228 VSS 0.14932f
C11737 a_71281_n8397.t30 VSS 0.33632f
C11738 a_71281_n8397.n229 VSS 0.14932f
C11739 a_71281_n8397.n230 VSS 0.042199f
C11740 a_71281_n8397.n231 VSS 0.01957f
C11741 a_71281_n8397.n232 VSS 0.221362f
C11742 a_71281_n8397.t7 VSS 0.159066f
C11743 a_71281_n8397.t31 VSS 0.033548f
C11744 a_71281_n8397.t39 VSS 0.033548f
C11745 a_71281_n8397.n233 VSS 0.136945f
C11746 a_71281_n8397.n234 VSS 0.382877f
C11747 a_71281_n8397.n235 VSS 0.092801f
C11748 a_71281_n8397.n236 VSS 0.221362f
C11749 a_71281_n8397.n237 VSS 0.047376f
C11750 a_71281_n8397.n238 VSS 0.43613f
C11751 a_71281_n8397.t116 VSS 0.421781f
C11752 a_71281_n8397.n239 VSS 0.43064f
C11753 a_71281_n8397.t301 VSS 0.382252f
C11754 a_71281_n8397.n240 VSS 0.43064f
C11755 a_71281_n8397.n241 VSS 0.047376f
C11756 a_71281_n8397.n242 VSS 0.01957f
C11757 a_71281_n8397.t204 VSS 0.421756f
C11758 a_71281_n8397.t196 VSS 0.382162f
C11759 a_71281_n8397.n243 VSS 0.43613f
C11760 a_71281_n8397.n244 VSS 0.042199f
C11761 a_71281_n8397.n245 VSS 0.14932f
C11762 a_71281_n8397.t211 VSS 0.33632f
C11763 a_71281_n8397.n246 VSS 0.14932f
C11764 a_71281_n8397.n247 VSS 0.042199f
C11765 a_71281_n8397.n248 VSS 0.01957f
C11766 a_71281_n8397.n249 VSS 0.268058f
C11767 a_71281_n8397.n250 VSS 0.267467f
C11768 a_71281_n8397.n251 VSS 0.047376f
C11769 a_71281_n8397.n252 VSS 0.43613f
C11770 a_71281_n8397.t105 VSS 0.421781f
C11771 a_71281_n8397.n253 VSS 0.43064f
C11772 a_71281_n8397.t294 VSS 0.382252f
C11773 a_71281_n8397.n254 VSS 0.43064f
C11774 a_71281_n8397.n255 VSS 0.047376f
C11775 a_71281_n8397.n256 VSS 0.01957f
C11776 a_71281_n8397.t198 VSS 0.421756f
C11777 a_71281_n8397.t183 VSS 0.382162f
C11778 a_71281_n8397.n257 VSS 0.43613f
C11779 a_71281_n8397.n258 VSS 0.042199f
C11780 a_71281_n8397.n259 VSS 0.14932f
C11781 a_71281_n8397.t202 VSS 0.33632f
C11782 a_71281_n8397.n260 VSS 0.14932f
C11783 a_71281_n8397.n261 VSS 0.042199f
C11784 a_71281_n8397.n262 VSS 0.01957f
C11785 a_71281_n8397.n263 VSS 0.267467f
C11786 a_71281_n8397.n264 VSS 0.267172f
C11787 a_71281_n8397.n265 VSS 0.047376f
C11788 a_71281_n8397.n266 VSS 0.43613f
C11789 a_71281_n8397.t129 VSS 0.421781f
C11790 a_71281_n8397.n267 VSS 0.43064f
C11791 a_71281_n8397.t317 VSS 0.382252f
C11792 a_71281_n8397.n268 VSS 0.43064f
C11793 a_71281_n8397.n269 VSS 0.047376f
C11794 a_71281_n8397.n270 VSS 0.01957f
C11795 a_71281_n8397.t215 VSS 0.421756f
C11796 a_71281_n8397.t209 VSS 0.382162f
C11797 a_71281_n8397.n271 VSS 0.43613f
C11798 a_71281_n8397.n272 VSS 0.042199f
C11799 a_71281_n8397.n273 VSS 0.14932f
C11800 a_71281_n8397.t219 VSS 0.33632f
C11801 a_71281_n8397.n274 VSS 0.14932f
C11802 a_71281_n8397.n275 VSS 0.042199f
C11803 a_71281_n8397.n276 VSS 0.01957f
C11804 a_71281_n8397.n277 VSS 0.267172f
C11805 a_71281_n8397.n278 VSS 0.267467f
C11806 a_71281_n8397.n279 VSS 0.047376f
C11807 a_71281_n8397.n280 VSS 0.43613f
C11808 a_71281_n8397.t312 VSS 0.418638f
C11809 a_71281_n8397.n281 VSS 0.43064f
C11810 a_71281_n8397.t249 VSS 0.382252f
C11811 a_71281_n8397.n282 VSS 0.419773f
C11812 a_71281_n8397.n283 VSS 0.047376f
C11813 a_71281_n8397.n284 VSS 0.01957f
C11814 a_71281_n8397.t143 VSS 0.421756f
C11815 a_71281_n8397.t133 VSS 0.382162f
C11816 a_71281_n8397.n285 VSS 0.43613f
C11817 a_71281_n8397.n286 VSS 0.042199f
C11818 a_71281_n8397.n287 VSS 0.14932f
C11819 a_71281_n8397.t148 VSS 0.33632f
C11820 a_71281_n8397.n288 VSS 0.14932f
C11821 a_71281_n8397.n289 VSS 0.042199f
C11822 a_71281_n8397.n290 VSS 0.01957f
C11823 a_71281_n8397.n291 VSS 0.607638f
C11824 a_71281_n8397.n292 VSS 2.23771f
C11825 a_71281_n8397.n293 VSS 0.051472f
C11826 a_71281_n8397.n294 VSS 0.047376f
C11827 a_71281_n8397.n295 VSS 0.43613f
C11828 a_71281_n8397.t226 VSS 0.418638f
C11829 a_71281_n8397.n296 VSS 0.419773f
C11830 a_71281_n8397.t190 VSS 0.382252f
C11831 a_71281_n8397.n297 VSS 0.43064f
C11832 a_71281_n8397.n298 VSS 0.047376f
C11833 a_71281_n8397.t126 VSS 0.421756f
C11834 a_71281_n8397.t91 VSS 0.382162f
C11835 a_71281_n8397.n299 VSS 0.43613f
C11836 a_71281_n8397.n300 VSS 0.042199f
C11837 a_71281_n8397.n301 VSS 0.14932f
C11838 a_71281_n8397.t277 VSS 0.33632f
C11839 a_71281_n8397.n302 VSS 0.14932f
C11840 a_71281_n8397.n303 VSS 0.042199f
C11841 a_71281_n8397.n304 VSS 0.01957f
C11842 a_71281_n8397.n305 VSS 0.533769f
C11843 a_71281_n8397.n306 VSS 0.267172f
C11844 a_71281_n8397.n307 VSS 0.047376f
C11845 a_71281_n8397.n308 VSS 0.43613f
C11846 a_71281_n8397.t289 VSS 0.421781f
C11847 a_71281_n8397.n309 VSS 0.43064f
C11848 a_71281_n8397.t258 VSS 0.382252f
C11849 a_71281_n8397.n310 VSS 0.43064f
C11850 a_71281_n8397.n311 VSS 0.047376f
C11851 a_71281_n8397.t201 VSS 0.421756f
C11852 a_71281_n8397.t166 VSS 0.382162f
C11853 a_71281_n8397.n312 VSS 0.43613f
C11854 a_71281_n8397.n313 VSS 0.01957f
C11855 a_71281_n8397.n314 VSS 0.042199f
C11856 a_71281_n8397.n315 VSS 0.14932f
C11857 a_71281_n8397.t76 VSS 0.33632f
C11858 a_71281_n8397.n316 VSS 0.14932f
C11859 a_71281_n8397.n317 VSS 0.042199f
C11860 a_71281_n8397.n318 VSS 0.01957f
C11861 a_71281_n8397.n319 VSS 0.267172f
C11862 a_71281_n8397.n320 VSS 0.267467f
C11863 a_71281_n8397.n321 VSS 0.047376f
C11864 a_71281_n8397.n322 VSS 0.43613f
C11865 a_71281_n8397.t283 VSS 0.421781f
C11866 a_71281_n8397.n323 VSS 0.43064f
C11867 a_71281_n8397.t247 VSS 0.382252f
C11868 a_71281_n8397.n324 VSS 0.43064f
C11869 a_71281_n8397.n325 VSS 0.047376f
C11870 a_71281_n8397.t192 VSS 0.421756f
C11871 a_71281_n8397.t160 VSS 0.382162f
C11872 a_71281_n8397.n326 VSS 0.43613f
C11873 a_71281_n8397.n327 VSS 0.01957f
C11874 a_71281_n8397.n328 VSS 0.042199f
C11875 a_71281_n8397.n329 VSS 0.14932f
C11876 a_71281_n8397.t332 VSS 0.33632f
C11877 a_71281_n8397.n330 VSS 0.14932f
C11878 a_71281_n8397.n331 VSS 0.042199f
C11879 a_71281_n8397.n332 VSS 0.01957f
C11880 a_71281_n8397.n333 VSS 0.267467f
C11881 a_71281_n8397.n334 VSS 0.268058f
C11882 a_71281_n8397.n335 VSS 0.047376f
C11883 a_71281_n8397.n336 VSS 0.43613f
C11884 a_71281_n8397.t90 VSS 0.421781f
C11885 a_71281_n8397.n337 VSS 0.43064f
C11886 a_71281_n8397.t315 VSS 0.382252f
C11887 a_71281_n8397.n338 VSS 0.43064f
C11888 a_71281_n8397.n339 VSS 0.047376f
C11889 a_71281_n8397.t260 VSS 0.421756f
C11890 a_71281_n8397.t230 VSS 0.382162f
C11891 a_71281_n8397.n340 VSS 0.43613f
C11892 a_71281_n8397.n341 VSS 0.01957f
C11893 a_71281_n8397.n342 VSS 0.042199f
C11894 a_71281_n8397.n343 VSS 0.14932f
C11895 a_71281_n8397.t146 VSS 0.33632f
C11896 a_71281_n8397.n344 VSS 0.14932f
C11897 a_71281_n8397.n345 VSS 0.042199f
C11898 a_71281_n8397.n346 VSS 0.01957f
C11899 a_71281_n8397.n347 VSS 0.221362f
C11900 a_71281_n8397.t5 VSS 0.159066f
C11901 a_71281_n8397.t55 VSS 0.033548f
C11902 a_71281_n8397.t25 VSS 0.033548f
C11903 a_71281_n8397.n348 VSS 0.136945f
C11904 a_71281_n8397.n349 VSS 0.382877f
C11905 a_71281_n8397.n350 VSS 0.092801f
C11906 a_71281_n8397.n351 VSS 0.221362f
C11907 a_71281_n8397.n352 VSS 0.047376f
C11908 a_71281_n8397.n353 VSS 0.43613f
C11909 a_71281_n8397.t85 VSS 0.421781f
C11910 a_71281_n8397.n354 VSS 0.43064f
C11911 a_71281_n8397.t4 VSS 0.382252f
C11912 a_71281_n8397.n355 VSS 0.43064f
C11913 a_71281_n8397.n356 VSS 0.047376f
C11914 a_71281_n8397.t248 VSS 0.421756f
C11915 a_71281_n8397.t24 VSS 0.382162f
C11916 a_71281_n8397.n357 VSS 0.43613f
C11917 a_71281_n8397.n358 VSS 0.01957f
C11918 a_71281_n8397.n359 VSS 0.042199f
C11919 a_71281_n8397.n360 VSS 0.14932f
C11920 a_71281_n8397.t54 VSS 0.33632f
C11921 a_71281_n8397.n361 VSS 0.14932f
C11922 a_71281_n8397.n362 VSS 0.042199f
C11923 a_71281_n8397.n363 VSS 0.01957f
C11924 a_71281_n8397.n364 VSS 0.267467f
C11925 a_71281_n8397.n365 VSS 0.267467f
C11926 a_71281_n8397.n366 VSS 0.047376f
C11927 a_71281_n8397.n367 VSS 0.43613f
C11928 a_71281_n8397.t158 VSS 0.421781f
C11929 a_71281_n8397.n368 VSS 0.43064f
C11930 a_71281_n8397.t58 VSS 0.382252f
C11931 a_71281_n8397.n369 VSS 0.43064f
C11932 a_71281_n8397.n370 VSS 0.047376f
C11933 a_71281_n8397.t316 VSS 0.421756f
C11934 a_71281_n8397.t8 VSS 0.382162f
C11935 a_71281_n8397.n371 VSS 0.43613f
C11936 a_71281_n8397.n372 VSS 0.01957f
C11937 a_71281_n8397.n373 VSS 0.042199f
C11938 a_71281_n8397.n374 VSS 0.14932f
C11939 a_71281_n8397.t26 VSS 0.33632f
C11940 a_71281_n8397.n375 VSS 0.14932f
C11941 a_71281_n8397.n376 VSS 0.042199f
C11942 a_71281_n8397.n377 VSS 0.01957f
C11943 a_71281_n8397.n378 VSS 0.221067f
C11944 a_71281_n8397.t59 VSS 0.033548f
C11945 a_71281_n8397.t27 VSS 0.033548f
C11946 a_71281_n8397.n379 VSS 0.136714f
C11947 a_71281_n8397.t9 VSS 0.159292f
C11948 a_71281_n8397.n380 VSS 0.384352f
C11949 a_71281_n8397.n381 VSS 0.092801f
C11950 a_71281_n8397.n382 VSS 0.220771f
C11951 a_71281_n8397.n383 VSS 0.047376f
C11952 a_71281_n8397.n384 VSS 0.43613f
C11953 a_71281_n8397.t139 VSS 0.421781f
C11954 a_71281_n8397.n385 VSS 0.43064f
C11955 a_71281_n8397.t93 VSS 0.382252f
C11956 a_71281_n8397.n386 VSS 0.43064f
C11957 a_71281_n8397.n387 VSS 0.047376f
C11958 a_71281_n8397.t293 VSS 0.421756f
C11959 a_71281_n8397.t275 VSS 0.382162f
C11960 a_71281_n8397.n388 VSS 0.43613f
C11961 a_71281_n8397.n389 VSS 0.01957f
C11962 a_71281_n8397.n390 VSS 0.042199f
C11963 a_71281_n8397.n391 VSS 0.14932f
C11964 a_71281_n8397.t189 VSS 0.33632f
C11965 a_71281_n8397.n392 VSS 0.14932f
C11966 a_71281_n8397.n393 VSS 0.042199f
C11967 a_71281_n8397.n394 VSS 0.01957f
C11968 a_71281_n8397.n395 VSS 0.267172f
C11969 a_71281_n8397.n396 VSS 0.267467f
C11970 a_71281_n8397.n397 VSS 0.047376f
C11971 a_71281_n8397.n398 VSS 0.43613f
C11972 a_71281_n8397.t213 VSS 0.421781f
C11973 a_71281_n8397.n399 VSS 0.43064f
C11974 a_71281_n8397.t167 VSS 0.382252f
C11975 a_71281_n8397.n400 VSS 0.43064f
C11976 a_71281_n8397.n401 VSS 0.047376f
C11977 a_71281_n8397.t110 VSS 0.421756f
C11978 a_71281_n8397.t74 VSS 0.382162f
C11979 a_71281_n8397.n402 VSS 0.43613f
C11980 a_71281_n8397.n403 VSS 0.01957f
C11981 a_71281_n8397.n404 VSS 0.042199f
C11982 a_71281_n8397.n405 VSS 0.14932f
C11983 a_71281_n8397.t257 VSS 0.33632f
C11984 a_71281_n8397.n406 VSS 0.14932f
C11985 a_71281_n8397.n407 VSS 0.042199f
C11986 a_71281_n8397.n408 VSS 0.01957f
C11987 a_71281_n8397.n409 VSS 0.267467f
C11988 a_71281_n8397.n410 VSS 0.268058f
C11989 a_71281_n8397.n411 VSS 0.047376f
C11990 a_71281_n8397.n412 VSS 0.43613f
C11991 a_71281_n8397.t207 VSS 0.421781f
C11992 a_71281_n8397.n413 VSS 0.43064f
C11993 a_71281_n8397.t161 VSS 0.382252f
C11994 a_71281_n8397.n414 VSS 0.43064f
C11995 a_71281_n8397.n415 VSS 0.047376f
C11996 a_71281_n8397.n416 VSS 0.01957f
C11997 a_71281_n8397.t97 VSS 0.421756f
C11998 a_71281_n8397.t331 VSS 0.382162f
C11999 a_71281_n8397.n417 VSS 0.43613f
C12000 a_71281_n8397.n418 VSS 0.042199f
C12001 a_71281_n8397.n419 VSS 0.14932f
C12002 a_71281_n8397.t246 VSS 0.33632f
C12003 a_71281_n8397.n420 VSS 0.14932f
C12004 a_71281_n8397.n421 VSS 0.042199f
C12005 a_71281_n8397.n422 VSS 0.01957f
C12006 a_71281_n8397.n423 VSS 0.268058f
C12007 a_71281_n8397.n424 VSS 0.267467f
C12008 a_71281_n8397.n425 VSS 0.047376f
C12009 a_71281_n8397.n426 VSS 0.43613f
C12010 a_71281_n8397.t274 VSS 0.421781f
C12011 a_71281_n8397.n427 VSS 0.43064f
C12012 a_71281_n8397.t231 VSS 0.382252f
C12013 a_71281_n8397.n428 VSS 0.43064f
C12014 a_71281_n8397.n429 VSS 0.047376f
C12015 a_71281_n8397.n430 VSS 0.01957f
C12016 a_71281_n8397.t170 VSS 0.421756f
C12017 a_71281_n8397.t145 VSS 0.382162f
C12018 a_71281_n8397.n431 VSS 0.43613f
C12019 a_71281_n8397.n432 VSS 0.042199f
C12020 a_71281_n8397.n433 VSS 0.14932f
C12021 a_71281_n8397.t314 VSS 0.33632f
C12022 a_71281_n8397.n434 VSS 0.14932f
C12023 a_71281_n8397.n435 VSS 0.042199f
C12024 a_71281_n8397.n436 VSS 0.01957f
C12025 a_71281_n8397.n437 VSS 0.605274f
C12026 a_71281_n8397.n438 VSS 0.052547f
C12027 a_71281_n8397.n439 VSS 0.047376f
C12028 a_71281_n8397.n440 VSS 0.43613f
C12029 a_71281_n8397.t75 VSS 0.421781f
C12030 a_71281_n8397.n441 VSS 0.43064f
C12031 a_71281_n8397.t188 VSS 0.382252f
C12032 a_71281_n8397.n442 VSS 0.43064f
C12033 a_71281_n8397.n443 VSS 0.047376f
C12034 a_71281_n8397.t173 VSS 0.421756f
C12035 a_71281_n8397.t157 VSS 0.382162f
C12036 a_71281_n8397.n444 VSS 0.43613f
C12037 a_71281_n8397.n445 VSS 0.042199f
C12038 a_71281_n8397.n446 VSS 0.14932f
C12039 a_71281_n8397.t172 VSS 0.33632f
C12040 a_71281_n8397.n447 VSS 0.14932f
C12041 a_71281_n8397.n448 VSS 0.042199f
C12042 a_71281_n8397.n449 VSS 0.01957f
C12043 a_71281_n8397.n450 VSS 0.542742f
C12044 a_71281_n8397.n451 VSS 0.268058f
C12045 a_71281_n8397.n452 VSS 0.047376f
C12046 a_71281_n8397.n453 VSS 0.43613f
C12047 a_71281_n8397.t276 VSS 0.421781f
C12048 a_71281_n8397.n454 VSS 0.43064f
C12049 a_71281_n8397.t117 VSS 0.382252f
C12050 a_71281_n8397.n455 VSS 0.43064f
C12051 a_71281_n8397.n456 VSS 0.047376f
C12052 a_71281_n8397.t101 VSS 0.421756f
C12053 a_71281_n8397.t84 VSS 0.382162f
C12054 a_71281_n8397.n457 VSS 0.43613f
C12055 a_71281_n8397.n458 VSS 0.01957f
C12056 a_71281_n8397.n459 VSS 0.042199f
C12057 a_71281_n8397.n460 VSS 0.14932f
C12058 a_71281_n8397.t99 VSS 0.33632f
C12059 a_71281_n8397.n461 VSS 0.14932f
C12060 a_71281_n8397.n462 VSS 0.042199f
C12061 a_71281_n8397.n463 VSS 0.01957f
C12062 a_71281_n8397.n464 VSS 0.268058f
C12063 a_71281_n8397.n465 VSS 0.267467f
C12064 a_71281_n8397.n466 VSS 0.047376f
C12065 a_71281_n8397.n467 VSS 0.43613f
C12066 a_71281_n8397.t142 VSS 0.421781f
C12067 a_71281_n8397.n468 VSS 0.43064f
C12068 a_71281_n8397.t244 VSS 0.382252f
C12069 a_71281_n8397.n469 VSS 0.43064f
C12070 a_71281_n8397.n470 VSS 0.047376f
C12071 a_71281_n8397.n471 VSS 0.01957f
C12072 a_71281_n8397.t232 VSS 0.421756f
C12073 a_71281_n8397.t221 VSS 0.382162f
C12074 a_71281_n8397.n472 VSS 0.43613f
C12075 a_71281_n8397.n473 VSS 0.042199f
C12076 a_71281_n8397.n474 VSS 0.14932f
C12077 a_71281_n8397.t229 VSS 0.33632f
C12078 a_71281_n8397.n475 VSS 0.14932f
C12079 a_71281_n8397.n476 VSS 0.042199f
C12080 a_71281_n8397.n477 VSS 0.01957f
C12081 a_71281_n8397.n478 VSS 0.267467f
C12082 a_71281_n8397.n479 VSS 0.267172f
C12083 a_71281_n8397.n480 VSS 0.047376f
C12084 a_71281_n8397.n481 VSS 0.43613f
C12085 a_71281_n8397.t330 VSS 0.421781f
C12086 a_71281_n8397.n482 VSS 0.43064f
C12087 a_71281_n8397.t175 VSS 0.382252f
C12088 a_71281_n8397.n483 VSS 0.43064f
C12089 a_71281_n8397.n484 VSS 0.047376f
C12090 a_71281_n8397.n485 VSS 0.01957f
C12091 a_71281_n8397.t162 VSS 0.421756f
C12092 a_71281_n8397.t150 VSS 0.382162f
C12093 a_71281_n8397.n486 VSS 0.43613f
C12094 a_71281_n8397.n487 VSS 0.042199f
C12095 a_71281_n8397.n488 VSS 0.14932f
C12096 a_71281_n8397.t159 VSS 0.33632f
C12097 a_71281_n8397.n489 VSS 0.14932f
C12098 a_71281_n8397.n490 VSS 0.042199f
C12099 a_71281_n8397.n491 VSS 0.01957f
C12100 a_71281_n8397.n492 VSS 0.220771f
C12101 a_71281_n8397.t37 VSS 0.033548f
C12102 a_71281_n8397.t49 VSS 0.033548f
C12103 a_71281_n8397.n493 VSS 0.136714f
C12104 a_71281_n8397.t51 VSS 0.159292f
C12105 a_71281_n8397.n494 VSS 0.384352f
C12106 a_71281_n8397.n495 VSS 0.092801f
C12107 a_71281_n8397.n496 VSS 0.221067f
C12108 a_71281_n8397.n497 VSS 0.047376f
C12109 a_71281_n8397.n498 VSS 0.43613f
C12110 a_71281_n8397.t336 VSS 0.421781f
C12111 a_71281_n8397.n499 VSS 0.43064f
C12112 a_71281_n8397.t36 VSS 0.382252f
C12113 a_71281_n8397.n500 VSS 0.43064f
C12114 a_71281_n8397.n501 VSS 0.047376f
C12115 a_71281_n8397.n502 VSS 0.01957f
C12116 a_71281_n8397.t168 VSS 0.421756f
C12117 a_71281_n8397.t50 VSS 0.382162f
C12118 a_71281_n8397.n503 VSS 0.43613f
C12119 a_71281_n8397.n504 VSS 0.042199f
C12120 a_71281_n8397.n505 VSS 0.14932f
C12121 a_71281_n8397.t48 VSS 0.33632f
C12122 a_71281_n8397.n506 VSS 0.14932f
C12123 a_71281_n8397.n507 VSS 0.042199f
C12124 a_71281_n8397.n508 VSS 0.01957f
C12125 a_71281_n8397.n509 VSS 0.267467f
C12126 a_71281_n8397.n510 VSS 0.267467f
C12127 a_71281_n8397.n511 VSS 0.047376f
C12128 a_71281_n8397.n512 VSS 0.43613f
C12129 a_71281_n8397.t271 VSS 0.421781f
C12130 a_71281_n8397.n513 VSS 0.43064f
C12131 a_71281_n8397.t62 VSS 0.382252f
C12132 a_71281_n8397.n514 VSS 0.43064f
C12133 a_71281_n8397.n515 VSS 0.047376f
C12134 a_71281_n8397.n516 VSS 0.01957f
C12135 a_71281_n8397.t94 VSS 0.421756f
C12136 a_71281_n8397.t70 VSS 0.382162f
C12137 a_71281_n8397.n517 VSS 0.43613f
C12138 a_71281_n8397.n518 VSS 0.042199f
C12139 a_71281_n8397.n519 VSS 0.14932f
C12140 a_71281_n8397.t68 VSS 0.33632f
C12141 a_71281_n8397.n520 VSS 0.14932f
C12142 a_71281_n8397.n521 VSS 0.042199f
C12143 a_71281_n8397.n522 VSS 0.01957f
C12144 a_71281_n8397.n523 VSS 0.221362f
C12145 a_71281_n8397.t63 VSS 0.159066f
C12146 a_71281_n8397.t69 VSS 0.033548f
C12147 a_71281_n8397.t71 VSS 0.033548f
C12148 a_71281_n8397.n524 VSS 0.136945f
C12149 a_71281_n8397.n525 VSS 0.382877f
C12150 a_71281_n8397.n526 VSS 0.092801f
C12151 a_71281_n8397.n527 VSS 0.221362f
C12152 a_71281_n8397.n528 VSS 0.047376f
C12153 a_71281_n8397.n529 VSS 0.43613f
C12154 a_71281_n8397.t280 VSS 0.421781f
C12155 a_71281_n8397.n530 VSS 0.43064f
C12156 a_71281_n8397.t122 VSS 0.382252f
C12157 a_71281_n8397.n531 VSS 0.43064f
C12158 a_71281_n8397.n532 VSS 0.047376f
C12159 a_71281_n8397.n533 VSS 0.01957f
C12160 a_71281_n8397.t108 VSS 0.421756f
C12161 a_71281_n8397.t88 VSS 0.382162f
C12162 a_71281_n8397.n534 VSS 0.43613f
C12163 a_71281_n8397.n535 VSS 0.042199f
C12164 a_71281_n8397.n536 VSS 0.14932f
C12165 a_71281_n8397.t107 VSS 0.33632f
C12166 a_71281_n8397.n537 VSS 0.14932f
C12167 a_71281_n8397.n538 VSS 0.042199f
C12168 a_71281_n8397.n539 VSS 0.01957f
C12169 a_71281_n8397.n540 VSS 0.268058f
C12170 a_71281_n8397.n541 VSS 0.267467f
C12171 a_71281_n8397.n542 VSS 0.047376f
C12172 a_71281_n8397.n543 VSS 0.43613f
C12173 a_71281_n8397.t272 VSS 0.421781f
C12174 a_71281_n8397.n544 VSS 0.43064f
C12175 a_71281_n8397.t114 VSS 0.382252f
C12176 a_71281_n8397.n545 VSS 0.43064f
C12177 a_71281_n8397.n546 VSS 0.047376f
C12178 a_71281_n8397.n547 VSS 0.01957f
C12179 a_71281_n8397.t95 VSS 0.421756f
C12180 a_71281_n8397.t80 VSS 0.382162f
C12181 a_71281_n8397.n548 VSS 0.43613f
C12182 a_71281_n8397.n549 VSS 0.042199f
C12183 a_71281_n8397.n550 VSS 0.14932f
C12184 a_71281_n8397.t92 VSS 0.33632f
C12185 a_71281_n8397.n551 VSS 0.14932f
C12186 a_71281_n8397.n552 VSS 0.042199f
C12187 a_71281_n8397.n553 VSS 0.01957f
C12188 a_71281_n8397.n554 VSS 0.267467f
C12189 a_71281_n8397.n555 VSS 0.267172f
C12190 a_71281_n8397.n556 VSS 0.047376f
C12191 a_71281_n8397.n557 VSS 0.43613f
C12192 a_71281_n8397.t285 VSS 0.421781f
C12193 a_71281_n8397.n558 VSS 0.43064f
C12194 a_71281_n8397.t135 VSS 0.382252f
C12195 a_71281_n8397.n559 VSS 0.43064f
C12196 a_71281_n8397.n560 VSS 0.047376f
C12197 a_71281_n8397.n561 VSS 0.01957f
C12198 a_71281_n8397.t123 VSS 0.421756f
C12199 a_71281_n8397.t106 VSS 0.382162f
C12200 a_71281_n8397.n562 VSS 0.43613f
C12201 a_71281_n8397.n563 VSS 0.042199f
C12202 a_71281_n8397.n564 VSS 0.14932f
C12203 a_71281_n8397.t121 VSS 0.33632f
C12204 a_71281_n8397.n565 VSS 0.14932f
C12205 a_71281_n8397.n566 VSS 0.042199f
C12206 a_71281_n8397.n567 VSS 0.01957f
C12207 a_71281_n8397.n568 VSS 0.267172f
C12208 a_71281_n8397.n569 VSS 0.267467f
C12209 a_71281_n8397.n570 VSS 0.047376f
C12210 a_71281_n8397.n571 VSS 0.43613f
C12211 a_71281_n8397.t225 VSS 0.418638f
C12212 a_71281_n8397.n572 VSS 0.43064f
C12213 a_71281_n8397.t320 VSS 0.382252f
C12214 a_71281_n8397.n573 VSS 0.419773f
C12215 a_71281_n8397.n574 VSS 0.047376f
C12216 a_71281_n8397.n575 VSS 0.01957f
C12217 a_71281_n8397.t304 VSS 0.421756f
C12218 a_71281_n8397.t291 VSS 0.382162f
C12219 a_71281_n8397.n576 VSS 0.43613f
C12220 a_71281_n8397.n577 VSS 0.042199f
C12221 a_71281_n8397.n578 VSS 0.14932f
C12222 a_71281_n8397.t303 VSS 0.33632f
C12223 a_71281_n8397.n579 VSS 0.14932f
C12224 a_71281_n8397.n580 VSS 0.042199f
C12225 a_71281_n8397.n581 VSS 0.01957f
C12226 a_71281_n8397.n582 VSS 0.607638f
C12227 a_71281_n8397.n583 VSS 0.863579f
C12228 a_71281_n8397.n584 VSS 2.75402f
C12229 a_71281_n8397.t0 VSS 0.413362f
C12230 a_71281_n8397.t1 VSS 0.96901f
C12231 a_71281_n8397.n585 VSS 8.049689f
C12232 a_71281_n8397.n586 VSS 0.051472f
C12233 a_71281_n8397.n587 VSS 0.047376f
C12234 a_71281_n8397.n588 VSS 0.43613f
C12235 a_71281_n8397.t206 VSS 0.418638f
C12236 a_71281_n8397.n589 VSS 0.419773f
C12237 a_71281_n8397.t256 VSS 0.382252f
C12238 a_71281_n8397.n590 VSS 0.43064f
C12239 a_71281_n8397.n591 VSS 0.047376f
C12240 a_71281_n8397.t120 VSS 0.421756f
C12241 a_71281_n8397.t321 VSS 0.382162f
C12242 a_71281_n8397.n592 VSS 0.43613f
C12243 a_71281_n8397.n593 VSS 0.042199f
C12244 a_71281_n8397.n594 VSS 0.14932f
C12245 a_71281_n8397.t265 VSS 0.33632f
C12246 a_71281_n8397.n595 VSS 0.14932f
C12247 a_71281_n8397.n596 VSS 0.042199f
C12248 a_71281_n8397.n597 VSS 0.01957f
C12249 a_71281_n8397.n598 VSS 0.533769f
C12250 a_71281_n8397.n599 VSS 0.267172f
C12251 a_71281_n8397.n600 VSS 0.047376f
C12252 a_71281_n8397.n601 VSS 0.43613f
C12253 a_71281_n8397.t270 VSS 0.421781f
C12254 a_71281_n8397.n602 VSS 0.43064f
C12255 a_71281_n8397.t323 VSS 0.382252f
C12256 a_71281_n8397.n603 VSS 0.43064f
C12257 a_71281_n8397.n604 VSS 0.047376f
C12258 a_71281_n8397.t195 VSS 0.421756f
C12259 a_71281_n8397.t136 VSS 0.382162f
C12260 a_71281_n8397.n605 VSS 0.43613f
C12261 a_71281_n8397.n606 VSS 0.01957f
C12262 a_71281_n8397.n607 VSS 0.042199f
C12263 a_71281_n8397.n608 VSS 0.14932f
C12264 a_71281_n8397.t333 VSS 0.33632f
C12265 a_71281_n8397.n609 VSS 0.14932f
C12266 a_71281_n8397.n610 VSS 0.042199f
C12267 a_71281_n8397.n611 VSS 0.01957f
C12268 a_71281_n8397.n612 VSS 0.267172f
C12269 a_71281_n8397.n613 VSS 0.267467f
C12270 a_71281_n8397.n614 VSS 0.047376f
C12271 a_71281_n8397.n615 VSS 0.43613f
C12272 a_71281_n8397.t263 VSS 0.421781f
C12273 a_71281_n8397.n616 VSS 0.43064f
C12274 a_71281_n8397.t313 VSS 0.382252f
C12275 a_71281_n8397.n617 VSS 0.43064f
C12276 a_71281_n8397.n618 VSS 0.047376f
C12277 a_71281_n8397.t182 VSS 0.421756f
C12278 a_71281_n8397.t128 VSS 0.382162f
C12279 a_71281_n8397.n619 VSS 0.43613f
C12280 a_71281_n8397.n620 VSS 0.01957f
C12281 a_71281_n8397.n621 VSS 0.042199f
C12282 a_71281_n8397.n622 VSS 0.14932f
C12283 a_71281_n8397.t325 VSS 0.33632f
C12284 a_71281_n8397.n623 VSS 0.14932f
C12285 a_71281_n8397.n624 VSS 0.042199f
C12286 a_71281_n8397.n625 VSS 0.01957f
C12287 a_71281_n8397.n626 VSS 0.267467f
C12288 a_71281_n8397.n627 VSS 0.268058f
C12289 a_71281_n8397.n628 VSS 0.047376f
C12290 a_71281_n8397.n629 VSS 0.43613f
C12291 a_71281_n8397.t329 VSS 0.421781f
C12292 a_71281_n8397.n630 VSS 0.43064f
C12293 a_71281_n8397.t130 VSS 0.382252f
C12294 a_71281_n8397.n631 VSS 0.43064f
C12295 a_71281_n8397.n632 VSS 0.047376f
C12296 a_71281_n8397.t251 VSS 0.421756f
C12297 a_71281_n8397.t203 VSS 0.382162f
C12298 a_71281_n8397.n633 VSS 0.43613f
C12299 a_71281_n8397.n634 VSS 0.01957f
C12300 a_71281_n8397.n635 VSS 0.042199f
C12301 a_71281_n8397.n636 VSS 0.14932f
C12302 a_71281_n8397.t138 VSS 0.33632f
C12303 a_71281_n8397.n637 VSS 0.14932f
C12304 a_71281_n8397.n638 VSS 0.042199f
C12305 a_71281_n8397.n639 VSS 0.01957f
C12306 a_71281_n8397.n640 VSS 0.221362f
C12307 a_71281_n8397.t61 VSS 0.159066f
C12308 a_71281_n8397.t57 VSS 0.033548f
C12309 a_71281_n8397.t35 VSS 0.033548f
C12310 a_71281_n8397.n641 VSS 0.136945f
C12311 a_71281_n8397.n642 VSS 0.382877f
C12312 a_71281_n8397.n643 VSS 0.092801f
C12313 a_71281_n8397.n644 VSS 0.221362f
C12314 a_71281_n8397.n645 VSS 0.047376f
C12315 a_71281_n8397.n646 VSS 0.43613f
C12316 a_71281_n8397.t322 VSS 0.421781f
C12317 a_71281_n8397.n647 VSS 0.43064f
C12318 a_71281_n8397.t60 VSS 0.382252f
C12319 a_71281_n8397.n648 VSS 0.43064f
C12320 a_71281_n8397.n649 VSS 0.047376f
C12321 a_71281_n8397.t241 VSS 0.421756f
C12322 a_71281_n8397.t34 VSS 0.382162f
C12323 a_71281_n8397.n650 VSS 0.43613f
C12324 a_71281_n8397.n651 VSS 0.01957f
C12325 a_71281_n8397.n652 VSS 0.042199f
C12326 a_71281_n8397.n653 VSS 0.14932f
C12327 a_71281_n8397.t56 VSS 0.33632f
C12328 a_71281_n8397.n654 VSS 0.14932f
C12329 a_71281_n8397.n655 VSS 0.042199f
C12330 a_71281_n8397.n656 VSS 0.01957f
C12331 a_71281_n8397.n657 VSS 0.267467f
C12332 a_71281_n8397.n658 VSS 0.267467f
C12333 a_71281_n8397.n659 VSS 0.047376f
C12334 a_71281_n8397.n660 VSS 0.43613f
C12335 a_71281_n8397.t137 VSS 0.421781f
C12336 a_71281_n8397.n661 VSS 0.43064f
C12337 a_71281_n8397.t32 VSS 0.382252f
C12338 a_71281_n8397.n662 VSS 0.43064f
C12339 a_71281_n8397.n663 VSS 0.047376f
C12340 a_71281_n8397.t308 VSS 0.421756f
C12341 a_71281_n8397.t14 VSS 0.382162f
C12342 a_71281_n8397.n664 VSS 0.43613f
C12343 a_71281_n8397.n665 VSS 0.01957f
C12344 a_71281_n8397.n666 VSS 0.042199f
C12345 a_71281_n8397.n667 VSS 0.14932f
C12346 a_71281_n8397.t28 VSS 0.33632f
C12347 a_71281_n8397.n668 VSS 0.14932f
C12348 a_71281_n8397.n669 VSS 0.042199f
C12349 a_71281_n8397.n670 VSS 0.01957f
C12350 a_71281_n8397.n671 VSS 0.221067f
C12351 a_71281_n8397.t33 VSS 0.033548f
C12352 a_71281_n8397.t29 VSS 0.033548f
C12353 a_71281_n8397.n672 VSS 0.136714f
C12354 a_71281_n8397.t15 VSS 0.159292f
C12355 a_71281_n8397.n673 VSS 0.384352f
C12356 a_71281_n8397.n674 VSS 0.092801f
C12357 a_71281_n8397.n675 VSS 0.220771f
C12358 a_71281_n8397.n676 VSS 0.047376f
C12359 a_71281_n8397.n677 VSS 0.43613f
C12360 a_71281_n8397.t115 VSS 0.421781f
C12361 a_71281_n8397.n678 VSS 0.43064f
C12362 a_71281_n8397.t165 VSS 0.382252f
C12363 a_71281_n8397.n679 VSS 0.43064f
C12364 a_71281_n8397.n680 VSS 0.047376f
C12365 a_71281_n8397.t287 VSS 0.421756f
C12366 a_71281_n8397.t235 VSS 0.382162f
C12367 a_71281_n8397.n681 VSS 0.43613f
C12368 a_71281_n8397.n682 VSS 0.01957f
C12369 a_71281_n8397.n683 VSS 0.042199f
C12370 a_71281_n8397.n684 VSS 0.14932f
C12371 a_71281_n8397.t180 VSS 0.33632f
C12372 a_71281_n8397.n685 VSS 0.14932f
C12373 a_71281_n8397.n686 VSS 0.042199f
C12374 a_71281_n8397.n687 VSS 0.01957f
C12375 a_71281_n8397.n688 VSS 0.267172f
C12376 a_71281_n8397.n689 VSS 0.267467f
C12377 a_71281_n8397.n690 VSS 0.047376f
C12378 a_71281_n8397.n691 VSS 0.43613f
C12379 a_71281_n8397.t185 VSS 0.421781f
C12380 a_71281_n8397.n692 VSS 0.43064f
C12381 a_71281_n8397.t237 VSS 0.382252f
C12382 a_71281_n8397.n693 VSS 0.43064f
C12383 a_71281_n8397.n694 VSS 0.047376f
C12384 a_71281_n8397.t100 VSS 0.421756f
C12385 a_71281_n8397.t302 VSS 0.382162f
C12386 a_71281_n8397.n695 VSS 0.43613f
C12387 a_71281_n8397.n696 VSS 0.01957f
C12388 a_71281_n8397.n697 VSS 0.042199f
C12389 a_71281_n8397.n698 VSS 0.14932f
C12390 a_71281_n8397.t250 VSS 0.33632f
C12391 a_71281_n8397.n699 VSS 0.14932f
C12392 a_71281_n8397.n700 VSS 0.042199f
C12393 a_71281_n8397.n701 VSS 0.01957f
C12394 a_71281_n8397.n702 VSS 0.267467f
C12395 a_71281_n8397.n703 VSS 0.268058f
C12396 a_71281_n8397.n704 VSS 0.047376f
C12397 a_71281_n8397.n705 VSS 0.43613f
C12398 a_71281_n8397.t176 VSS 0.421781f
C12399 a_71281_n8397.n706 VSS 0.43064f
C12400 a_71281_n8397.t228 VSS 0.382252f
C12401 a_71281_n8397.n707 VSS 0.43064f
C12402 a_71281_n8397.n708 VSS 0.047376f
C12403 a_71281_n8397.n709 VSS 0.01957f
C12404 a_71281_n8397.t89 VSS 0.421756f
C12405 a_71281_n8397.t296 VSS 0.382162f
C12406 a_71281_n8397.n710 VSS 0.43613f
C12407 a_71281_n8397.n711 VSS 0.042199f
C12408 a_71281_n8397.n712 VSS 0.14932f
C12409 a_71281_n8397.t238 VSS 0.33632f
C12410 a_71281_n8397.n713 VSS 0.14932f
C12411 a_71281_n8397.n714 VSS 0.042199f
C12412 a_71281_n8397.n715 VSS 0.01957f
C12413 a_71281_n8397.n716 VSS 0.268058f
C12414 a_71281_n8397.n717 VSS 0.267467f
C12415 a_71281_n8397.n718 VSS 0.047376f
C12416 a_71281_n8397.n719 VSS 0.43613f
C12417 a_71281_n8397.t245 VSS 0.421781f
C12418 a_71281_n8397.n720 VSS 0.43064f
C12419 a_71281_n8397.t297 VSS 0.382252f
C12420 a_71281_n8397.n721 VSS 0.43064f
C12421 a_71281_n8397.n722 VSS 0.047376f
C12422 a_71281_n8397.n723 VSS 0.01957f
C12423 a_71281_n8397.t163 VSS 0.421756f
C12424 a_71281_n8397.t112 VSS 0.382162f
C12425 a_71281_n8397.n724 VSS 0.43613f
C12426 a_71281_n8397.n725 VSS 0.042199f
C12427 a_71281_n8397.n726 VSS 0.14932f
C12428 a_71281_n8397.t305 VSS 0.33632f
C12429 a_71281_n8397.n727 VSS 0.14932f
C12430 a_71281_n8397.n728 VSS 0.042199f
C12431 a_71281_n8397.n729 VSS 0.01957f
C12432 a_71281_n8397.n730 VSS 0.58961f
C12433 a_71281_n8397.n731 VSS 0.605438f
C12434 a_71281_n8397.n732 VSS 0.047376f
C12435 a_71281_n8397.n733 VSS 0.43613f
C12436 a_71281_n8397.t223 VSS 0.418638f
C12437 a_71281_n8397.n734 VSS 0.419773f
C12438 a_71281_n8397.t124 VSS 0.382252f
C12439 a_71281_n8397.n735 VSS 0.43064f
C12440 a_71281_n8397.n736 VSS 0.047376f
C12441 a_71281_n8397.t290 VSS 0.421756f
C12442 a_71281_n8397.t132 VSS 0.382162f
C12443 a_71281_n8397.n737 VSS 0.43613f
C12444 a_71281_n8397.n738 VSS 0.01957f
C12445 a_71281_n8397.n739 VSS 0.042199f
C12446 a_71281_n8397.n740 VSS 0.14932f
C12447 a_71281_n8397.t288 VSS 0.33632f
C12448 a_71281_n8397.n741 VSS 0.14932f
C12449 a_71281_n8397.n742 VSS 0.042199f
C12450 a_71281_n8397.n743 VSS 0.01957f
C12451 a_71281_n8397.n744 VSS 0.267467f
C12452 a_71281_n8397.n745 VSS 0.267172f
C12453 a_71281_n8397.n746 VSS 0.047376f
C12454 a_71281_n8397.n747 VSS 0.43613f
C12455 a_71281_n8397.t284 VSS 0.421781f
C12456 a_71281_n8397.n748 VSS 0.43064f
C12457 a_71281_n8397.t199 VSS 0.382252f
C12458 a_71281_n8397.n749 VSS 0.43064f
C12459 a_71281_n8397.n750 VSS 0.047376f
C12460 a_71281_n8397.t104 VSS 0.421756f
C12461 a_71281_n8397.t208 VSS 0.382162f
C12462 a_71281_n8397.n751 VSS 0.43613f
C12463 a_71281_n8397.n752 VSS 0.01957f
C12464 a_71281_n8397.n753 VSS 0.042199f
C12465 a_71281_n8397.n754 VSS 0.14932f
C12466 a_71281_n8397.t102 VSS 0.33632f
C12467 a_71281_n8397.n755 VSS 0.14932f
C12468 a_71281_n8397.n756 VSS 0.042199f
C12469 a_71281_n8397.n757 VSS 0.01957f
C12470 a_71281_n8397.n758 VSS 0.267172f
C12471 a_71281_n8397.n759 VSS 0.267467f
C12472 a_71281_n8397.n760 VSS 0.047376f
C12473 a_71281_n8397.n761 VSS 0.43613f
C12474 a_71281_n8397.t267 VSS 0.421781f
C12475 a_71281_n8397.n762 VSS 0.43064f
C12476 a_71281_n8397.t171 VSS 0.382252f
C12477 a_71281_n8397.n763 VSS 0.43064f
C12478 a_71281_n8397.n764 VSS 0.047376f
C12479 a_71281_n8397.t79 VSS 0.421756f
C12480 a_71281_n8397.t181 VSS 0.382162f
C12481 a_71281_n8397.n765 VSS 0.43613f
C12482 a_71281_n8397.n766 VSS 0.01957f
C12483 a_71281_n8397.n767 VSS 0.042199f
C12484 a_71281_n8397.n768 VSS 0.14932f
C12485 a_71281_n8397.t77 VSS 0.33632f
C12486 a_71281_n8397.n769 VSS 0.14932f
C12487 a_71281_n8397.n770 VSS 0.042199f
C12488 a_71281_n8397.n771 VSS 0.01957f
C12489 a_71281_n8397.n772 VSS 0.267467f
C12490 a_71281_n8397.n773 VSS 0.268058f
C12491 a_71281_n8397.n774 VSS 0.047376f
C12492 a_71281_n8397.n775 VSS 0.43613f
C12493 a_71281_n8397.t279 VSS 0.421781f
C12494 a_71281_n8397.n776 VSS 0.43064f
C12495 a_71281_n8397.t179 VSS 0.382252f
C12496 a_71281_n8397.n777 VSS 0.43064f
C12497 a_71281_n8397.n778 VSS 0.047376f
C12498 a_71281_n8397.t87 VSS 0.421756f
C12499 a_71281_n8397.t194 VSS 0.382162f
C12500 a_71281_n8397.n779 VSS 0.43613f
C12501 a_71281_n8397.n780 VSS 0.01957f
C12502 a_71281_n8397.n781 VSS 0.042199f
C12503 a_71281_n8397.n782 VSS 0.14932f
C12504 a_71281_n8397.t86 VSS 0.33632f
C12505 a_71281_n8397.n783 VSS 0.14932f
C12506 a_71281_n8397.n784 VSS 0.042199f
C12507 a_71281_n8397.n785 VSS 0.01957f
C12508 a_71281_n8397.n786 VSS 0.221362f
C12509 a_71281_n8397.n787 VSS 0.052547f
C12510 a_71281_n8397.n788 VSS 0.047376f
C12511 a_71281_n8397.n789 VSS 0.43613f
C12512 a_71281_n8397.t337 VSS 0.421781f
C12513 a_71281_n8397.n790 VSS 0.43064f
C12514 a_71281_n8397.t243 VSS 0.382252f
C12515 a_71281_n8397.n791 VSS 0.43064f
C12516 a_71281_n8397.n792 VSS 0.047376f
C12517 a_71281_n8397.t156 VSS 0.421756f
C12518 a_71281_n8397.t254 VSS 0.382162f
C12519 a_71281_n8397.n793 VSS 0.43613f
C12520 a_71281_n8397.n794 VSS 0.042199f
C12521 a_71281_n8397.n795 VSS 0.14932f
C12522 a_71281_n8397.t155 VSS 0.33632f
C12523 a_71281_n8397.n796 VSS 0.14932f
C12524 a_71281_n8397.n797 VSS 0.042199f
C12525 a_71281_n8397.n798 VSS 0.01957f
C12526 a_71281_n8397.n799 VSS 0.542742f
C12527 a_71281_n8397.n800 VSS 0.268058f
C12528 a_71281_n8397.n801 VSS 0.047376f
C12529 a_71281_n8397.n802 VSS 0.43613f
C12530 a_71281_n8397.t273 VSS 0.421781f
C12531 a_71281_n8397.n803 VSS 0.43064f
C12532 a_71281_n8397.t174 VSS 0.382252f
C12533 a_71281_n8397.n804 VSS 0.43064f
C12534 a_71281_n8397.n805 VSS 0.047376f
C12535 a_71281_n8397.t83 VSS 0.421756f
C12536 a_71281_n8397.t186 VSS 0.382162f
C12537 a_71281_n8397.n806 VSS 0.43613f
C12538 a_71281_n8397.n807 VSS 0.01957f
C12539 a_71281_n8397.n808 VSS 0.042199f
C12540 a_71281_n8397.n809 VSS 0.14932f
C12541 a_71281_n8397.t82 VSS 0.33632f
C12542 a_71281_n8397.n810 VSS 0.14932f
C12543 a_71281_n8397.n811 VSS 0.042199f
C12544 a_71281_n8397.n812 VSS 0.01957f
C12545 a_71281_n8397.n813 VSS 0.268058f
C12546 a_71281_n8397.n814 VSS 0.267467f
C12547 a_71281_n8397.n815 VSS 0.047376f
C12548 a_71281_n8397.n816 VSS 0.43613f
C12549 a_71281_n8397.t140 VSS 0.421781f
C12550 a_71281_n8397.n817 VSS 0.43064f
C12551 a_71281_n8397.t299 VSS 0.382252f
C12552 a_71281_n8397.n818 VSS 0.43064f
C12553 a_71281_n8397.n819 VSS 0.047376f
C12554 a_71281_n8397.n820 VSS 0.01957f
C12555 a_71281_n8397.t220 VSS 0.421756f
C12556 a_71281_n8397.t306 VSS 0.382162f
C12557 a_71281_n8397.n821 VSS 0.43613f
C12558 a_71281_n8397.n822 VSS 0.042199f
C12559 a_71281_n8397.n823 VSS 0.14932f
C12560 a_71281_n8397.t218 VSS 0.33632f
C12561 a_71281_n8397.n824 VSS 0.14932f
C12562 a_71281_n8397.n825 VSS 0.042199f
C12563 a_71281_n8397.n826 VSS 0.01957f
C12564 a_71281_n8397.n827 VSS 0.267467f
C12565 a_71281_n8397.n828 VSS 0.267172f
C12566 a_71281_n8397.n829 VSS 0.047376f
C12567 a_71281_n8397.n830 VSS 0.43613f
C12568 a_71281_n8397.t327 VSS 0.421781f
C12569 a_71281_n8397.n831 VSS 0.43064f
C12570 a_71281_n8397.t233 VSS 0.382252f
C12571 a_71281_n8397.n832 VSS 0.43064f
C12572 a_71281_n8397.n833 VSS 0.047376f
C12573 a_71281_n8397.n834 VSS 0.01957f
C12574 a_71281_n8397.t149 VSS 0.421756f
C12575 a_71281_n8397.t239 VSS 0.382162f
C12576 a_71281_n8397.n835 VSS 0.43613f
C12577 a_71281_n8397.n836 VSS 0.042199f
C12578 a_71281_n8397.n837 VSS 0.14932f
C12579 a_71281_n8397.t147 VSS 0.33632f
C12580 a_71281_n8397.n838 VSS 0.14932f
C12581 a_71281_n8397.n839 VSS 0.042199f
C12582 a_71281_n8397.n840 VSS 0.01957f
C12583 a_71281_n8397.n841 VSS 0.220771f
C12584 a_71281_n8397.t23 VSS 0.033548f
C12585 a_71281_n8397.t53 VSS 0.033548f
C12586 a_71281_n8397.n842 VSS 0.136714f
C12587 a_71281_n8397.t19 VSS 0.159292f
C12588 a_71281_n8397.n843 VSS 0.384352f
C12589 a_71281_n8397.n844 VSS 0.092801f
C12590 a_71281_n8397.n845 VSS 0.221067f
C12591 a_71281_n8397.n846 VSS 0.047376f
C12592 a_71281_n8397.n847 VSS 0.43613f
C12593 a_71281_n8397.t334 VSS 0.421781f
C12594 a_71281_n8397.n848 VSS 0.43064f
C12595 a_71281_n8397.t22 VSS 0.382252f
C12596 a_71281_n8397.n849 VSS 0.43064f
C12597 a_71281_n8397.n850 VSS 0.047376f
C12598 a_71281_n8397.n851 VSS 0.01957f
C12599 a_71281_n8397.t153 VSS 0.421756f
C12600 a_71281_n8397.t18 VSS 0.382162f
C12601 a_71281_n8397.n852 VSS 0.43613f
C12602 a_71281_n8397.n853 VSS 0.042199f
C12603 a_71281_n8397.n854 VSS 0.14932f
C12604 a_71281_n8397.t52 VSS 0.33632f
C12605 a_71281_n8397.n855 VSS 0.14932f
C12606 a_71281_n8397.n856 VSS 0.042199f
C12607 a_71281_n8397.n857 VSS 0.01957f
C12608 a_71281_n8397.n858 VSS 0.267467f
C12609 a_71281_n8397.n859 VSS 0.267467f
C12610 a_71281_n8397.n860 VSS 0.047376f
C12611 a_71281_n8397.n861 VSS 0.43613f
C12612 a_71281_n8397.t266 VSS 0.421781f
C12613 a_71281_n8397.n862 VSS 0.43064f
C12614 a_71281_n8397.t44 VSS 0.382252f
C12615 a_71281_n8397.n863 VSS 0.43064f
C12616 a_71281_n8397.n864 VSS 0.047376f
C12617 a_71281_n8397.n865 VSS 0.01957f
C12618 a_71281_n8397.t78 VSS 0.421756f
C12619 a_71281_n8397.t40 VSS 0.382162f
C12620 a_71281_n8397.n866 VSS 0.43613f
C12621 a_71281_n8397.n867 VSS 0.042199f
C12622 a_71281_n8397.n868 VSS 0.14932f
C12623 a_71281_n8397.t72 VSS 0.33632f
C12624 a_71281_n8397.n869 VSS 0.14932f
C12625 a_71281_n8397.n870 VSS 0.042199f
C12626 a_71281_n8397.n871 VSS 0.01957f
C12627 a_71281_n8397.n872 VSS 0.221362f
C12628 a_71281_n8397.n873 VSS 0.092801f
C12629 a_71281_n8397.n874 VSS 0.382877f
C12630 a_71281_n8397.n875 VSS 0.136945f
C12631 a_71281_n8397.t73 VSS 0.033548f
C12632 a_41891_4481.t8 VSS 3.64456f
C12633 a_41891_4481.n0 VSS 0.449404f
C12634 a_41891_4481.n1 VSS 7.74464f
C12635 a_41891_4481.t10 VSS 0.182047f
C12636 a_41891_4481.t5 VSS 0.177333f
C12637 a_41891_4481.t3 VSS 0.152849f
C12638 a_41891_4481.t4 VSS 0.296925f
C12639 a_41891_4481.t13 VSS 0.284336f
C12640 a_41891_4481.t15 VSS 0.293711f
C12641 a_41891_4481.t22 VSS 0.296925f
C12642 a_41891_4481.t11 VSS 0.284336f
C12643 a_41891_4481.t16 VSS 0.296925f
C12644 a_41891_4481.t17 VSS 0.284336f
C12645 a_41891_4481.t0 VSS 0.294005f
C12646 a_41891_4481.t18 VSS 0.284359f
C12647 a_41891_4481.t7 VSS 0.177256f
C12648 a_41891_4481.t1 VSS 0.152918f
C12649 a_41891_4481.t6 VSS 0.296925f
C12650 a_41891_4481.t19 VSS 0.284336f
C12651 a_41891_4481.t21 VSS 0.293956f
C12652 a_41891_4481.t20 VSS 0.284359f
C12653 a_41891_4481.t12 VSS 0.284359f
C12654 a_41891_4481.t2 VSS 0.293809f
C12655 a_41891_4481.t14 VSS 0.284359f
C12656 a_41891_4481.t9 VSS 0.181041f
C12657 a_35502_24538.n0 VSS 0.201745f
C12658 a_35502_24538.n1 VSS 0.078965f
C12659 a_35502_24538.n2 VSS 0.096477f
C12660 a_35502_24538.n3 VSS 0.632723f
C12661 a_35502_24538.n4 VSS 0.137716f
C12662 a_35502_24538.n5 VSS 0.193543f
C12663 a_35502_24538.n6 VSS 0.104977f
C12664 a_35502_24538.n7 VSS 0.600521f
C12665 a_35502_24538.n8 VSS 0.113978f
C12666 a_35502_24538.n9 VSS 0.109075f
C12667 a_35502_24538.n10 VSS 0.096479f
C12668 a_35502_24538.n11 VSS 0.629354f
C12669 a_35502_24538.n12 VSS 0.136805f
C12670 a_35502_24538.n13 VSS 0.635197f
C12671 a_35502_24538.n14 VSS 0.137729f
C12672 a_35502_24538.n15 VSS 0.190479f
C12673 a_35502_24538.n16 VSS 0.073508f
C12674 a_35502_24538.n17 VSS 0.619589f
C12675 a_35502_24538.n18 VSS 0.114969f
C12676 a_35502_24538.n19 VSS 0.109124f
C12677 a_35502_24538.n20 VSS 0.090985f
C12678 a_35502_24538.n21 VSS 0.602671f
C12679 a_35502_24538.n22 VSS 0.136797f
C12680 a_35502_24538.n23 VSS 0.141765f
C12681 a_35502_24538.n24 VSS 0.142077f
C12682 a_35502_24538.n25 VSS 0.570993f
C12683 a_35502_24538.n26 VSS 0.222694f
C12684 a_35502_24538.n27 VSS 0.085585f
C12685 a_35502_24538.n28 VSS 0.124773f
C12686 a_35502_24538.n29 VSS 0.028484f
C12687 a_35502_24538.n30 VSS 0.128481f
C12688 a_35502_24538.n31 VSS 0.079331f
C12689 a_35502_24538.n32 VSS 0.139369f
C12690 a_35502_24538.n33 VSS 0.059376f
C12691 a_35502_24538.n34 VSS 0.36666f
C12692 a_35502_24538.n35 VSS 0.218793f
C12693 a_35502_24538.n36 VSS 0.121372f
C12694 a_35502_24538.n37 VSS 0.083195f
C12695 a_35502_24538.n38 VSS 0.103461f
C12696 a_35502_24538.n39 VSS 0.071225f
C12697 a_35502_24538.n40 VSS 0.011258f
C12698 a_35502_24538.n41 VSS 0.117227f
C12699 a_35502_24538.n42 VSS 0.083694f
C12700 a_35502_24538.t15 VSS 0.139537f
C12701 a_35502_24538.t17 VSS 0.138296f
C12702 a_35502_24538.n43 VSS 0.224747f
C12703 a_35502_24538.n44 VSS 0.028183f
C12704 a_35502_24538.t12 VSS 0.069849f
C12705 a_35502_24538.t9 VSS 0.070288f
C12706 a_35502_24538.t7 VSS 0.143318f
C12707 a_35502_24538.t22 VSS 0.027467f
C12708 a_35502_24538.t16 VSS 0.027467f
C12709 a_35502_24538.n45 VSS 0.106345f
C12710 a_35502_24538.n46 VSS 0.365826f
C12711 a_35502_24538.t6 VSS 0.105876f
C12712 a_35502_24538.n47 VSS 0.222541f
C12713 a_35502_24538.t2 VSS 0.027467f
C12714 a_35502_24538.t20 VSS 0.027467f
C12715 a_35502_24538.n48 VSS 0.106848f
C12716 a_35502_24538.n49 VSS 0.188808f
C12717 a_35502_24538.n50 VSS 0.011258f
C12718 a_35502_24538.n51 VSS 0.117541f
C12719 a_35502_24538.n52 VSS 0.077316f
C12720 a_35502_24538.t10 VSS 0.027467f
C12721 a_35502_24538.t19 VSS 0.027467f
C12722 a_35502_24538.n53 VSS 0.066763f
C12723 a_35502_24538.n54 VSS 0.10193f
C12724 a_35502_24538.n55 VSS 0.066459f
C12725 a_35502_24538.n56 VSS 0.718125f
C12726 a_35502_24538.t34 VSS 0.169702f
C12727 a_35502_24538.t36 VSS 0.170464f
C12728 a_35502_24538.n57 VSS 0.293172f
C12729 a_35502_24538.t56 VSS 0.169697f
C12730 a_35502_24538.t59 VSS 0.170495f
C12731 a_35502_24538.n58 VSS 0.282922f
C12732 a_35502_24538.n59 VSS 0.460003f
C12733 a_35502_24538.t41 VSS 0.169697f
C12734 a_35502_24538.t1 VSS 0.039575f
C12735 a_35502_24538.t0 VSS 0.148476f
C12736 a_35502_24538.n60 VSS 0.165749f
C12737 a_35502_24538.n61 VSS 0.199677f
C12738 a_35502_24538.n62 VSS 0.354733f
C12739 a_35502_24538.t26 VSS 0.228116f
C12740 a_35502_24538.n63 VSS 0.190127f
C12741 a_35502_24538.n64 VSS 0.13653f
C12742 a_35502_24538.t24 VSS 0.228116f
C12743 a_35502_24538.n65 VSS 0.137964f
C12744 a_35502_24538.t53 VSS 0.228116f
C12745 a_35502_24538.t42 VSS 0.228116f
C12746 a_35502_24538.n66 VSS 0.081574f
C12747 a_35502_24538.n67 VSS 0.066113f
C12748 a_35502_24538.t55 VSS 0.228116f
C12749 a_35502_24538.t40 VSS 0.228116f
C12750 a_35502_24538.t48 VSS 0.228116f
C12751 a_35502_24538.t50 VSS 0.228116f
C12752 a_35502_24538.t38 VSS 0.228116f
C12753 a_35502_24538.n68 VSS 0.028483f
C12754 a_35502_24538.n69 VSS 0.076493f
C12755 a_35502_24538.n70 VSS 0.146275f
C12756 a_35502_24538.t46 VSS 0.228116f
C12757 a_35502_24538.n71 VSS 0.183849f
C12758 a_35502_24538.n72 VSS 0.137994f
C12759 a_35502_24538.t37 VSS 0.228116f
C12760 a_35502_24538.t49 VSS 0.228116f
C12761 a_35502_24538.n73 VSS 0.138006f
C12762 a_35502_24538.t64 VSS 0.228116f
C12763 a_35502_24538.n74 VSS 0.081616f
C12764 a_35502_24538.n75 VSS 0.066093f
C12765 a_35502_24538.t32 VSS 0.228116f
C12766 a_35502_24538.t60 VSS 0.228116f
C12767 a_35502_24538.t33 VSS 0.228116f
C12768 a_35502_24538.n76 VSS 0.141777f
C12769 a_35502_24538.t62 VSS 0.228116f
C12770 a_35502_24538.n77 VSS 0.126233f
C12771 a_35502_24538.n78 VSS 0.080239f
C12772 a_35502_24538.t31 VSS 0.228116f
C12773 a_35502_24538.n79 VSS 2.41886f
C12774 a_35502_24538.n80 VSS 0.135374f
C12775 a_35502_24538.n81 VSS 0.023547f
C12776 a_35502_24538.n82 VSS 0.122525f
C12777 a_35502_24538.t47 VSS 0.231588f
C12778 a_35502_24538.n83 VSS 0.176835f
C12779 a_35502_24538.t35 VSS 0.228116f
C12780 a_35502_24538.n84 VSS 0.112114f
C12781 a_35502_24538.n85 VSS 0.009506f
C12782 a_35502_24538.n86 VSS 0.023547f
C12783 a_35502_24538.n87 VSS 0.024786f
C12784 a_35502_24538.n88 VSS 0.024786f
C12785 a_35502_24538.n89 VSS 0.016219f
C12786 a_35502_24538.n90 VSS 0.009443f
C12787 a_35502_24538.t63 VSS 0.228116f
C12788 a_35502_24538.n91 VSS 0.088267f
C12789 a_35502_24538.n92 VSS 0.077816f
C12790 a_35502_24538.t45 VSS 0.228116f
C12791 a_35502_24538.n93 VSS 0.18615f
C12792 a_35502_24538.t30 VSS 0.228116f
C12793 a_35502_24538.n94 VSS 0.150147f
C12794 a_35502_24538.t57 VSS 0.228116f
C12795 a_35502_24538.n95 VSS 0.184907f
C12796 a_35502_24538.n96 VSS 0.026715f
C12797 a_35502_24538.t61 VSS 0.233364f
C12798 a_35502_24538.t29 VSS 0.228116f
C12799 a_35502_24538.n97 VSS 0.116813f
C12800 a_35502_24538.n98 VSS 0.195195f
C12801 a_35502_24538.n99 VSS 0.147461f
C12802 a_35502_24538.t28 VSS 0.228116f
C12803 a_35502_24538.n100 VSS 0.62344f
C12804 a_35502_24538.n101 VSS 0.134066f
C12805 a_35502_24538.n102 VSS 0.016219f
C12806 a_35502_24538.n103 VSS 0.027585f
C12807 a_35502_24538.t25 VSS 0.233246f
C12808 a_35502_24538.n104 VSS 0.190643f
C12809 a_35502_24538.t54 VSS 0.228116f
C12810 a_35502_24538.n105 VSS 0.116626f
C12811 a_35502_24538.n106 VSS 0.026591f
C12812 a_35502_24538.n107 VSS 0.133837f
C12813 a_35502_24538.n108 VSS 0.029037f
C12814 a_35502_24538.n109 VSS 0.016219f
C12815 a_35502_24538.n110 VSS 0.008201f
C12816 a_35502_24538.t43 VSS 0.228116f
C12817 a_35502_24538.n111 VSS 0.088267f
C12818 a_35502_24538.n112 VSS 0.077738f
C12819 a_35502_24538.t27 VSS 0.228116f
C12820 a_35502_24538.n113 VSS 0.185901f
C12821 a_35502_24538.t58 VSS 0.228116f
C12822 a_35502_24538.n114 VSS 0.151062f
C12823 a_35502_24538.t44 VSS 0.228116f
C12824 a_35502_24538.n115 VSS 0.183966f
C12825 a_35502_24538.n116 VSS 0.027585f
C12826 a_35502_24538.t39 VSS 0.231588f
C12827 a_35502_24538.n117 VSS 0.182036f
C12828 a_35502_24538.t52 VSS 0.228116f
C12829 a_35502_24538.n118 VSS 0.111126f
C12830 a_35502_24538.n119 VSS 0.008698f
C12831 a_35502_24538.n120 VSS 0.126334f
C12832 a_35502_24538.n121 VSS 0.029037f
C12833 a_35502_24538.n122 VSS 0.029037f
C12834 a_35502_24538.n123 VSS 0.026094f
C12835 a_35502_24538.t51 VSS 0.228116f
C12836 a_35502_24538.n124 VSS 0.088267f
C12837 a_35502_24538.n125 VSS 0.009195f
C12838 a_35502_24538.n126 VSS 0.076193f
C12839 a_35502_24538.n127 VSS 0.049833f
C12840 a_35502_24538.n128 VSS 0.167681f
C12841 a_35502_24538.n129 VSS 2.23998f
C12842 a_35502_24538.n130 VSS 4.67369f
C12843 a_35502_24538.n131 VSS 4.46256f
C12844 a_35502_24538.n132 VSS 2.59861f
C12845 a_35502_24538.n133 VSS 0.015737f
C12846 a_35502_24538.n134 VSS 0.22611f
C12847 a_35502_24538.t8 VSS 0.027467f
C12848 a_35502_24538.t18 VSS 0.027467f
C12849 a_35502_24538.n135 VSS 0.067342f
C12850 a_35502_24538.t11 VSS 0.106676f
C12851 a_35502_24538.t14 VSS 0.027467f
C12852 a_35502_24538.t5 VSS 0.027467f
C12853 a_35502_24538.n136 VSS 0.106232f
C12854 a_35502_24538.n137 VSS 0.187325f
C12855 a_35502_24538.t21 VSS 0.027467f
C12856 a_35502_24538.t13 VSS 0.027467f
C12857 a_35502_24538.n138 VSS 0.10729f
C12858 a_35502_24538.t4 VSS 0.144332f
C12859 a_35502_24538.t3 VSS 0.070259f
C12860 a_35502_24538.n139 VSS 0.027073f
C12861 a_35502_24538.n140 VSS 0.081594f
C12862 a_35502_24538.n141 VSS 0.117852f
C12863 a_35502_24538.t23 VSS 0.069878f
C12864 a_31699_20742.n0 VSS 0.33657f
C12865 a_31699_20742.n1 VSS 0.252378f
C12866 a_31699_20742.n2 VSS 0.119729f
C12867 a_31699_20742.n3 VSS 0.252378f
C12868 a_31699_20742.n4 VSS 0.119608f
C12869 a_31699_20742.n5 VSS 0.252378f
C12870 a_31699_20742.n6 VSS 0.227077f
C12871 a_31699_20742.n7 VSS 0.33657f
C12872 a_31699_20742.n8 VSS 0.252378f
C12873 a_31699_20742.n9 VSS 0.119729f
C12874 a_31699_20742.n10 VSS 0.229433f
C12875 a_31699_20742.n11 VSS 0.252378f
C12876 a_31699_20742.n12 VSS 0.119608f
C12877 a_31699_20742.n13 VSS 0.33657f
C12878 a_31699_20742.n14 VSS 0.252378f
C12879 a_31699_20742.n15 VSS 0.227077f
C12880 a_31699_20742.n16 VSS 0.25941f
C12881 a_31699_20742.n17 VSS 0.230515f
C12882 a_31699_20742.n18 VSS 0.25941f
C12883 a_31699_20742.n19 VSS 0.127036f
C12884 a_31699_20742.n20 VSS 0.25941f
C12885 a_31699_20742.n21 VSS 0.127153f
C12886 a_31699_20742.n22 VSS 0.25941f
C12887 a_31699_20742.n23 VSS 0.230515f
C12888 a_31699_20742.n24 VSS 0.25941f
C12889 a_31699_20742.n25 VSS 0.127036f
C12890 a_31699_20742.n26 VSS 0.25941f
C12891 a_31699_20742.n27 VSS 0.127153f
C12892 a_31699_20742.n28 VSS 0.343765f
C12893 a_31699_20742.n29 VSS 0.149348f
C12894 a_31699_20742.n30 VSS 0.343765f
C12895 a_31699_20742.n31 VSS 0.149348f
C12896 a_31699_20742.n32 VSS 0.343765f
C12897 a_31699_20742.n33 VSS 0.149348f
C12898 a_31699_20742.n34 VSS 0.343765f
C12899 a_31699_20742.n35 VSS 0.149348f
C12900 a_31699_20742.n36 VSS 0.283994f
C12901 a_31699_20742.n37 VSS 0.33657f
C12902 a_31699_20742.n38 VSS 0.283994f
C12903 a_31699_20742.n39 VSS 0.283994f
C12904 a_31699_20742.n40 VSS 0.283994f
C12905 a_31699_20742.n41 VSS 0.340692f
C12906 a_31699_20742.n42 VSS 0.145738f
C12907 a_31699_20742.n43 VSS 0.257836f
C12908 a_31699_20742.n44 VSS 0.232767f
C12909 a_31699_20742.n45 VSS 0.257836f
C12910 a_31699_20742.n46 VSS 0.109525f
C12911 a_31699_20742.n47 VSS 0.257836f
C12912 a_31699_20742.n48 VSS 0.125496f
C12913 a_31699_20742.n49 VSS 0.341462f
C12914 a_31699_20742.n50 VSS 0.288981f
C12915 a_31699_20742.n51 VSS 0.145738f
C12916 a_31699_20742.n52 VSS 0.340692f
C12917 a_31699_20742.n53 VSS 0.257836f
C12918 a_31699_20742.n54 VSS 0.125496f
C12919 a_31699_20742.n55 VSS 0.257836f
C12920 a_31699_20742.n56 VSS 0.125352f
C12921 a_31699_20742.n57 VSS 0.257836f
C12922 a_31699_20742.n58 VSS 0.109525f
C12923 a_31699_20742.n59 VSS 0.341462f
C12924 a_31699_20742.n60 VSS 0.288981f
C12925 a_31699_20742.n61 VSS 0.340692f
C12926 a_31699_20742.n62 VSS 0.145738f
C12927 a_31699_20742.n63 VSS 0.257836f
C12928 a_31699_20742.n64 VSS 0.232767f
C12929 a_31699_20742.n65 VSS 0.257836f
C12930 a_31699_20742.n66 VSS 0.109525f
C12931 a_31699_20742.n67 VSS 0.257836f
C12932 a_31699_20742.n68 VSS 0.125496f
C12933 a_31699_20742.n69 VSS 0.341462f
C12934 a_31699_20742.n70 VSS 0.288981f
C12935 a_31699_20742.n71 VSS 0.340692f
C12936 a_31699_20742.n72 VSS 0.145738f
C12937 a_31699_20742.n73 VSS 0.257836f
C12938 a_31699_20742.n74 VSS 0.125496f
C12939 a_31699_20742.n75 VSS 0.257836f
C12940 a_31699_20742.n76 VSS 0.125352f
C12941 a_31699_20742.n77 VSS 0.257836f
C12942 a_31699_20742.n78 VSS 0.109525f
C12943 a_31699_20742.n79 VSS 0.341462f
C12944 a_31699_20742.n80 VSS 0.288981f
C12945 a_31699_20742.n81 VSS 0.257731f
C12946 a_31699_20742.n82 VSS 0.109266f
C12947 a_31699_20742.n83 VSS 1.05167f
C12948 a_31699_20742.n84 VSS 0.247803f
C12949 a_31699_20742.n85 VSS 0.245079f
C12950 a_31699_20742.n86 VSS 1.07804f
C12951 a_31699_20742.n87 VSS 1.05555f
C12952 a_31699_20742.n88 VSS 0.507149f
C12953 a_31699_20742.n89 VSS 0.507183f
C12954 a_31699_20742.n90 VSS 2.03605f
C12955 a_31699_20742.n91 VSS 0.828639f
C12956 a_31699_20742.n92 VSS 1.07804f
C12957 a_31699_20742.n93 VSS 1.05167f
C12958 a_31699_20742.n94 VSS 0.247811f
C12959 a_31699_20742.n95 VSS 0.245088f
C12960 a_31699_20742.n96 VSS 1.07804f
C12961 a_31699_20742.n97 VSS 1.05555f
C12962 a_31699_20742.n98 VSS 0.507129f
C12963 a_31699_20742.n99 VSS 0.507162f
C12964 a_31699_20742.n100 VSS 2.03605f
C12965 a_31699_20742.n101 VSS 0.828643f
C12966 a_31699_20742.n102 VSS 1.07386f
C12967 a_31699_20742.n103 VSS 1.0203f
C12968 a_31699_20742.n104 VSS 0.507172f
C12969 a_31699_20742.n105 VSS 0.507172f
C12970 a_31699_20742.n106 VSS 1.07386f
C12971 a_31699_20742.n107 VSS 1.0203f
C12972 a_31699_20742.n108 VSS 0.24561f
C12973 a_31699_20742.n109 VSS 0.245082f
C12974 a_31699_20742.n110 VSS 1.0203f
C12975 a_31699_20742.n111 VSS 0.507172f
C12976 a_31699_20742.n112 VSS 0.507172f
C12977 a_31699_20742.n113 VSS 1.0203f
C12978 a_31699_20742.n114 VSS 0.24561f
C12979 a_31699_20742.n115 VSS 0.245082f
C12980 a_31699_20742.n116 VSS 0.281749f
C12981 a_31699_20742.n117 VSS 0.37602f
C12982 a_31699_20742.n118 VSS 0.506958f
C12983 a_31699_20742.n119 VSS 0.506958f
C12984 a_31699_20742.n120 VSS 0.950455f
C12985 a_31699_20742.n121 VSS 1.07386f
C12986 a_31699_20742.n122 VSS 0.378143f
C12987 a_31699_20742.n123 VSS 0.460311f
C12988 a_31699_20742.n124 VSS 1.07386f
C12989 a_31699_20742.n125 VSS 0.281749f
C12990 a_31699_20742.n126 VSS 0.37602f
C12991 a_31699_20742.n127 VSS 1.07386f
C12992 a_31699_20742.n128 VSS 0.506958f
C12993 a_31699_20742.n129 VSS 0.506958f
C12994 a_31699_20742.n130 VSS 0.950455f
C12995 a_31699_20742.n131 VSS 1.07386f
C12996 a_31699_20742.n132 VSS 0.378143f
C12997 a_31699_20742.n133 VSS 0.460311f
C12998 a_31699_20742.n134 VSS 1.00324f
C12999 a_31699_20742.n135 VSS 0.374031f
C13000 a_31699_20742.n136 VSS 1.00324f
C13001 a_31699_20742.n137 VSS 0.374031f
C13002 a_31699_20742.n138 VSS 0.255397f
C13003 a_31699_20742.n139 VSS 0.358947f
C13004 a_31699_20742.n140 VSS 0.358947f
C13005 a_31699_20742.n141 VSS 0.255397f
C13006 a_31699_20742.n142 VSS 0.232798f
C13007 a_31699_20742.n143 VSS 0.38794f
C13008 a_31699_20742.n144 VSS 0.232798f
C13009 a_31699_20742.n145 VSS 0.38794f
C13010 a_31699_20742.n146 VSS 0.380618f
C13011 a_31699_20742.n147 VSS 0.229433f
C13012 a_31699_20742.n148 VSS 0.380618f
C13013 a_31699_20742.n149 VSS 0.281749f
C13014 a_31699_20742.n150 VSS 0.375336f
C13015 a_31699_20742.n151 VSS 0.506964f
C13016 a_31699_20742.n152 VSS 0.507147f
C13017 a_31699_20742.n153 VSS 1.07804f
C13018 a_31699_20742.n154 VSS 0.379124f
C13019 a_31699_20742.n155 VSS 0.460319f
C13020 a_31699_20742.n156 VSS 0.281745f
C13021 a_31699_20742.n157 VSS 0.375333f
C13022 a_31699_20742.n158 VSS 0.967909f
C13023 a_31699_20742.n159 VSS 1.07804f
C13024 a_31699_20742.n160 VSS 0.379124f
C13025 a_31699_20742.n161 VSS 0.460319f
C13026 a_31699_20742.n162 VSS 1.07804f
C13027 a_31699_20742.n163 VSS 0.506972f
C13028 a_31699_20742.n164 VSS 0.507155f
C13029 a_31699_20742.n165 VSS 1.0203f
C13030 a_31699_20742.n166 VSS 0.32944f
C13031 a_31699_20742.n167 VSS 0.330046f
C13032 a_31699_20742.n168 VSS 1.0203f
C13033 a_31699_20742.n169 VSS 0.32944f
C13034 a_31699_20742.n170 VSS 0.330046f
C13035 a_31699_20742.n171 VSS 0.390877f
C13036 a_31699_20742.n172 VSS 0.390877f
C13037 a_31699_20742.n173 VSS 1.02306f
C13038 a_31699_20742.n174 VSS 0.248142f
C13039 a_31699_20742.n175 VSS 0.467178f
C13040 a_31699_20742.n176 VSS 1.02306f
C13041 a_31699_20742.n177 VSS 0.248142f
C13042 a_31699_20742.n178 VSS 0.467178f
C13043 a_31699_20742.n179 VSS 1.02306f
C13044 a_31699_20742.n180 VSS 0.248142f
C13045 a_31699_20742.n181 VSS 0.467178f
C13046 a_31699_20742.n182 VSS 1.02306f
C13047 a_31699_20742.n183 VSS 0.248142f
C13048 a_31699_20742.n184 VSS 0.237296f
C13049 a_31699_20742.n185 VSS 0.15405f
C13050 a_31699_20742.n186 VSS 0.232006f
C13051 a_31699_20742.n187 VSS 0.375474f
C13052 a_31699_20742.n188 VSS 0.359299f
C13053 a_31699_20742.n189 VSS 0.249781f
C13054 a_31699_20742.n190 VSS 0.232006f
C13055 a_31699_20742.n191 VSS 0.375474f
C13056 a_31699_20742.n192 VSS 0.249781f
C13057 a_31699_20742.n193 VSS 0.359299f
C13058 a_31699_20742.n194 VSS 0.31207f
C13059 a_31699_20742.n195 VSS 0.31207f
C13060 a_31699_20742.n196 VSS 0.317556f
C13061 a_31699_20742.n197 VSS 1.06707f
C13062 a_31699_20742.n198 VSS 1.06813f
C13063 a_31699_20742.n199 VSS 0.248121f
C13064 a_31699_20742.n200 VSS 0.487063f
C13065 a_31699_20742.n201 VSS 1.06813f
C13066 a_31699_20742.n202 VSS 0.248121f
C13067 a_31699_20742.n203 VSS 0.487063f
C13068 a_31699_20742.n204 VSS 1.06813f
C13069 a_31699_20742.n205 VSS 0.248121f
C13070 a_31699_20742.n206 VSS 1.06813f
C13071 a_31699_20742.n207 VSS 0.248121f
C13072 a_31699_20742.n208 VSS 1.04026f
C13073 a_31699_20742.n209 VSS 2.17076f
C13074 a_31699_20742.n210 VSS 0.238189f
C13075 a_31699_20742.n211 VSS 0.35906f
C13076 a_31699_20742.n212 VSS 0.238189f
C13077 a_31699_20742.n213 VSS 0.35906f
C13078 a_31699_20742.n214 VSS 0.967909f
C13079 a_31699_20742.n215 VSS 0.411198f
C13080 a_31699_20742.n216 VSS 0.411198f
C13081 a_31699_20742.n217 VSS 0.712129f
C13082 a_31699_20742.n218 VSS 0.497515f
C13083 a_31699_20742.n219 VSS 0.467178f
C13084 a_31699_20742.n220 VSS 0.22427f
C13085 a_31699_20742.n221 VSS 0.22427f
C13086 a_31699_20742.n222 VSS 0.22427f
C13087 a_31699_20742.n223 VSS 0.22427f
C13088 a_31699_20742.n224 VSS 0.376149f
C13089 a_31699_20742.n225 VSS 0.376149f
C13090 a_31699_20742.n226 VSS 0.487063f
C13091 a_31699_20742.n227 VSS 0.224273f
C13092 a_31699_20742.n228 VSS 0.338926f
C13093 a_31699_20742.n229 VSS 0.22429f
C13094 a_31699_20742.n230 VSS 0.487063f
C13095 a_31699_20742.n231 VSS 0.338925f
C13096 a_31699_20742.n232 VSS 0.537276f
C13097 a_31699_20742.n233 VSS 0.529413f
C13098 a_31699_20742.n234 VSS 0.14727f
C13099 a_31699_20742.n235 VSS 0.49195f
C13100 a_31699_20742.n236 VSS 0.964513f
C13101 a_31699_20742.n237 VSS 1.07595f
C13102 a_31699_20742.n238 VSS 0.37478f
C13103 a_31699_20742.n239 VSS 0.94551f
C13104 a_31699_20742.n240 VSS 0.363125f
C13105 a_31699_20742.n241 VSS 0.627318f
C13106 a_31699_20742.t20 VSS 0.046398f
C13107 a_31699_20742.t12 VSS 0.246181f
C13108 a_31699_20742.t6 VSS 0.182618f
C13109 a_31699_20742.t32 VSS 0.182353f
C13110 a_31699_20742.t22 VSS 0.046398f
C13111 a_31699_20742.t10 VSS 0.046398f
C13112 a_31699_20742.n242 VSS 0.184107f
C13113 a_31699_20742.t2 VSS 0.249568f
C13114 a_31699_20742.t34 VSS 0.046398f
C13115 a_31699_20742.t8 VSS 0.046398f
C13116 a_31699_20742.n243 VSS 0.18758f
C13117 a_31699_20742.n244 VSS 0.635542f
C13118 a_31699_20742.t38 VSS 0.185553f
C13119 a_31699_20742.n245 VSS 0.541928f
C13120 a_31699_20742.t26 VSS 0.185553f
C13121 a_31699_20742.n246 VSS 0.534748f
C13122 a_31699_20742.t28 VSS 0.249791f
C13123 a_31699_20742.t16 VSS 0.046398f
C13124 a_31699_20742.t42 VSS 0.046398f
C13125 a_31699_20742.n247 VSS 0.18758f
C13126 a_31699_20742.t24 VSS 0.046398f
C13127 a_31699_20742.t14 VSS 0.046398f
C13128 a_31699_20742.n248 VSS 0.117306f
C13129 a_31699_20742.t18 VSS 0.046398f
C13130 a_31699_20742.t40 VSS 0.046398f
C13131 a_31699_20742.n249 VSS 0.107477f
C13132 a_31699_20742.n250 VSS 0.662865f
C13133 a_31699_20742.t4 VSS 0.121773f
C13134 a_31699_20742.t30 VSS 0.113301f
C13135 a_31699_20742.n251 VSS 3.58253f
C13136 a_31699_20742.n252 VSS 2.7071f
C13137 a_31699_20742.n253 VSS 2.75045f
C13138 a_31699_20742.t146 VSS 0.38723f
C13139 a_31699_20742.t90 VSS 0.38723f
C13140 a_31699_20742.t238 VSS 0.38723f
C13141 a_31699_20742.t187 VSS 0.38723f
C13142 a_31699_20742.t156 VSS 0.38723f
C13143 a_31699_20742.t221 VSS 0.38723f
C13144 a_31699_20742.t124 VSS 0.38723f
C13145 a_31699_20742.t166 VSS 0.38723f
C13146 a_31699_20742.t217 VSS 0.38723f
C13147 a_31699_20742.t70 VSS 0.38723f
C13148 a_31699_20742.t237 VSS 0.38723f
C13149 a_31699_20742.t63 VSS 0.38723f
C13150 a_31699_20742.t168 VSS 0.38723f
C13151 a_31699_20742.t97 VSS 0.38723f
C13152 a_31699_20742.t152 VSS 0.38723f
C13153 a_31699_20742.t106 VSS 0.38723f
C13154 a_31699_20742.t100 VSS 0.38723f
C13155 a_31699_20742.t181 VSS 0.38723f
C13156 a_31699_20742.t230 VSS 0.38723f
C13157 a_31699_20742.t77 VSS 0.38723f
C13158 a_31699_20742.t145 VSS 0.38723f
C13159 a_31699_20742.t174 VSS 0.38723f
C13160 a_31699_20742.t74 VSS 0.38723f
C13161 a_31699_20742.t66 VSS 0.38723f
C13162 a_31699_20742.t161 VSS 0.38723f
C13163 a_31699_20742.t209 VSS 0.38723f
C13164 a_31699_20742.t59 VSS 0.38723f
C13165 a_31699_20742.t154 VSS 0.38723f
C13166 a_31699_20742.t247 VSS 0.38723f
C13167 a_31699_20742.t214 VSS 0.38723f
C13168 a_31699_20742.t139 VSS 0.38723f
C13169 a_31699_20742.t216 VSS 0.38723f
C13170 a_31699_20742.t258 VSS 0.38723f
C13171 a_31699_20742.t78 VSS 0.38723f
C13172 a_31699_20742.t76 VSS 0.38723f
C13173 a_31699_20742.t227 VSS 0.38723f
C13174 a_31699_20742.t151 VSS 0.38723f
C13175 a_31699_20742.t84 VSS 0.38723f
C13176 a_31699_20742.n254 VSS 4.29884f
C13177 a_31699_20742.n255 VSS 0.376149f
C13178 a_31699_20742.t83 VSS 0.38723f
C13179 a_31699_20742.t93 VSS 0.38723f
C13180 a_31699_20742.t245 VSS 0.38723f
C13181 a_31699_20742.t170 VSS 0.38723f
C13182 a_31699_20742.t125 VSS 0.38723f
C13183 a_31699_20742.t157 VSS 0.38723f
C13184 a_31699_20742.t56 VSS 0.38723f
C13185 a_31699_20742.t236 VSS 0.38723f
C13186 a_31699_20742.t229 VSS 0.38723f
C13187 a_31699_20742.t249 VSS 0.38723f
C13188 a_31699_20742.t243 VSS 0.38723f
C13189 a_31699_20742.t136 VSS 0.38723f
C13190 a_31699_20742.t233 VSS 0.38723f
C13191 a_31699_20742.t86 VSS 0.38723f
C13192 a_31699_20742.t159 VSS 0.38723f
C13193 a_31699_20742.t205 VSS 0.38723f
C13194 a_31699_20742.t158 VSS 0.38723f
C13195 a_31699_20742.n256 VSS 4.29884f
C13196 a_31699_20742.t211 VSS 0.38723f
C13197 a_31699_20742.t193 VSS 0.38723f
C13198 a_31699_20742.t68 VSS 0.38723f
C13199 a_31699_20742.t200 VSS 0.38723f
C13200 a_31699_20742.t54 VSS 0.38723f
C13201 a_31699_20742.t135 VSS 0.38723f
C13202 a_31699_20742.t88 VSS 0.38723f
C13203 a_31699_20742.t210 VSS 0.38723f
C13204 a_31699_20742.t80 VSS 0.38723f
C13205 a_31699_20742.t203 VSS 0.38723f
C13206 a_31699_20742.t232 VSS 0.38723f
C13207 a_31699_20742.n257 VSS 0.486196f
C13208 a_31699_20742.t117 VSS 0.38723f
C13209 a_31699_20742.t215 VSS 0.38723f
C13210 a_31699_20742.t57 VSS 0.38723f
C13211 a_31699_20742.t133 VSS 0.38723f
C13212 a_31699_20742.t206 VSS 0.38723f
C13213 a_31699_20742.t61 VSS 0.38723f
C13214 a_31699_20742.t155 VSS 0.38723f
C13215 a_31699_20742.t122 VSS 0.38723f
C13216 a_31699_20742.t49 VSS 0.38723f
C13217 a_31699_20742.t123 VSS 0.38723f
C13218 a_31699_20742.t167 VSS 0.38723f
C13219 a_31699_20742.n258 VSS 2.75045f
C13220 a_31699_20742.n259 VSS 2.75045f
C13221 a_31699_20742.t113 VSS 0.38723f
C13222 a_31699_20742.n260 VSS 0.186129f
C13223 a_31699_20742.t188 VSS 0.38723f
C13224 a_31699_20742.t96 VSS 0.38723f
C13225 a_31699_20742.t176 VSS 0.38723f
C13226 a_31699_20742.t109 VSS 0.38723f
C13227 a_31699_20742.t253 VSS 0.38723f
C13228 a_31699_20742.n261 VSS 0.201867f
C13229 a_31699_20742.t207 VSS 0.395552f
C13230 a_31699_20742.n262 VSS 0.28878f
C13231 a_31699_20742.n263 VSS 0.193918f
C13232 a_31699_20742.n264 VSS 0.046177f
C13233 a_31699_20742.n265 VSS 1.06707f
C13234 a_31699_20742.n266 VSS 0.046177f
C13235 a_31699_20742.t194 VSS 0.38723f
C13236 a_31699_20742.n267 VSS 0.201867f
C13237 a_31699_20742.t142 VSS 0.395552f
C13238 a_31699_20742.n268 VSS 0.28878f
C13239 a_31699_20742.n269 VSS 0.193918f
C13240 a_31699_20742.t262 VSS 0.38723f
C13241 a_31699_20742.t112 VSS 0.38723f
C13242 a_31699_20742.t64 VSS 0.38723f
C13243 a_31699_20742.n270 VSS 0.31358f
C13244 a_31699_20742.t137 VSS 0.38723f
C13245 a_31699_20742.n271 VSS 0.257836f
C13246 a_31699_20742.t257 VSS 0.38723f
C13247 a_31699_20742.n272 VSS 0.312671f
C13248 a_31699_20742.t171 VSS 0.38723f
C13249 a_31699_20742.t246 VSS 0.38723f
C13250 a_31699_20742.n273 VSS 0.073985f
C13251 a_31699_20742.t115 VSS 0.38723f
C13252 a_31699_20742.t190 VSS 0.38723f
C13253 a_31699_20742.t261 VSS 0.38723f
C13254 a_31699_20742.t47 VSS 0.38723f
C13255 a_31699_20742.t129 VSS 0.38723f
C13256 a_31699_20742.t208 VSS 0.38723f
C13257 a_31699_20742.t160 VSS 0.398966f
C13258 a_31699_20742.t58 VSS 0.38723f
C13259 a_31699_20742.t120 VSS 0.38723f
C13260 a_31699_20742.n274 VSS 0.315849f
C13261 a_31699_20742.t195 VSS 0.38723f
C13262 a_31699_20742.n275 VSS 0.257836f
C13263 a_31699_20742.t95 VSS 0.38723f
C13264 a_31699_20742.n276 VSS 0.316105f
C13265 a_31699_20742.t140 VSS 0.38723f
C13266 a_31699_20742.t189 VSS 0.38723f
C13267 a_31699_20742.t260 VSS 0.38723f
C13268 a_31699_20742.t65 VSS 0.38723f
C13269 a_31699_20742.t132 VSS 0.38723f
C13270 a_31699_20742.t204 VSS 0.38723f
C13271 a_31699_20742.t55 VSS 0.38723f
C13272 a_31699_20742.t99 VSS 0.38723f
C13273 a_31699_20742.n277 VSS 0.315849f
C13274 a_31699_20742.t173 VSS 0.38723f
C13275 a_31699_20742.n278 VSS 0.257836f
C13276 a_31699_20742.t264 VSS 0.38723f
C13277 a_31699_20742.n279 VSS 0.316105f
C13278 a_31699_20742.t121 VSS 0.38723f
C13279 a_31699_20742.t198 VSS 0.38723f
C13280 a_31699_20742.t242 VSS 0.397787f
C13281 a_31699_20742.t196 VSS 0.38723f
C13282 a_31699_20742.n280 VSS 4.13948f
C13283 a_31699_20742.n281 VSS 0.31207f
C13284 a_31699_20742.t177 VSS 0.38723f
C13285 a_31699_20742.t105 VSS 0.38723f
C13286 a_31699_20742.t179 VSS 0.38723f
C13287 a_31699_20742.t228 VSS 0.398677f
C13288 a_31699_20742.t212 VSS 0.38723f
C13289 a_31699_20742.n282 VSS 0.312671f
C13290 a_31699_20742.t119 VSS 0.38723f
C13291 a_31699_20742.n283 VSS 0.257836f
C13292 a_31699_20742.t263 VSS 0.38723f
C13293 a_31699_20742.n284 VSS 0.31358f
C13294 a_31699_20742.n285 VSS 0.046177f
C13295 a_31699_20742.t48 VSS 0.38723f
C13296 a_31699_20742.n286 VSS 0.186129f
C13297 a_31699_20742.n287 VSS 0.331197f
C13298 a_31699_20742.t126 VSS 0.38723f
C13299 a_31699_20742.t251 VSS 0.38723f
C13300 a_31699_20742.n288 VSS 4.13948f
C13301 a_31699_20742.t67 VSS 0.398966f
C13302 a_31699_20742.t116 VSS 0.38723f
C13303 a_31699_20742.t191 VSS 0.38723f
C13304 a_31699_20742.t254 VSS 0.38723f
C13305 a_31699_20742.t248 VSS 0.38723f
C13306 a_31699_20742.n289 VSS 0.315849f
C13307 a_31699_20742.t101 VSS 0.38723f
C13308 a_31699_20742.n290 VSS 0.257836f
C13309 a_31699_20742.t225 VSS 0.38723f
C13310 a_31699_20742.n291 VSS 0.316105f
C13311 a_31699_20742.t50 VSS 0.38723f
C13312 a_31699_20742.t98 VSS 0.38723f
C13313 a_31699_20742.t259 VSS 0.38723f
C13314 a_31699_20742.t114 VSS 0.38723f
C13315 a_31699_20742.n292 VSS 0.317556f
C13316 a_31699_20742.t186 VSS 0.38723f
C13317 a_31699_20742.t102 VSS 0.38723f
C13318 a_31699_20742.t250 VSS 0.38723f
C13319 a_31699_20742.t103 VSS 0.38723f
C13320 a_31699_20742.t148 VSS 0.397787f
C13321 a_31699_20742.t175 VSS 0.38723f
C13322 a_31699_20742.n293 VSS 0.316105f
C13323 a_31699_20742.t79 VSS 0.38723f
C13324 a_31699_20742.n294 VSS 0.257836f
C13325 a_31699_20742.t231 VSS 0.38723f
C13326 a_31699_20742.n295 VSS 0.315849f
C13327 a_31699_20742.t197 VSS 0.38723f
C13328 a_31699_20742.t169 VSS 0.38723f
C13329 a_31699_20742.t178 VSS 0.38723f
C13330 a_31699_20742.n296 VSS 2.75045f
C13331 a_31699_20742.n297 VSS 2.49429f
C13332 a_31699_20742.n298 VSS 0.31207f
C13333 a_31699_20742.t130 VSS 0.38723f
C13334 a_31699_20742.n299 VSS 0.31358f
C13335 a_31699_20742.t202 VSS 0.38723f
C13336 a_31699_20742.n300 VSS 0.257836f
C13337 a_31699_20742.t104 VSS 0.38723f
C13338 a_31699_20742.n301 VSS 0.312671f
C13339 a_31699_20742.t239 VSS 0.38723f
C13340 a_31699_20742.t91 VSS 0.38723f
C13341 a_31699_20742.n302 VSS 0.331197f
C13342 a_31699_20742.n303 VSS 0.073985f
C13343 a_31699_20742.n304 VSS 0.046177f
C13344 a_31699_20742.t182 VSS 0.38723f
C13345 a_31699_20742.t252 VSS 0.38723f
C13346 a_31699_20742.t107 VSS 0.38723f
C13347 a_31699_20742.t110 VSS 0.38723f
C13348 a_31699_20742.n305 VSS 0.31358f
C13349 a_31699_20742.t183 VSS 0.38723f
C13350 a_31699_20742.n306 VSS 0.257836f
C13351 a_31699_20742.t53 VSS 0.38723f
C13352 a_31699_20742.n307 VSS 0.312671f
C13353 a_31699_20742.t69 VSS 0.398677f
C13354 a_31699_20742.t241 VSS 0.38723f
C13355 a_31699_20742.t165 VSS 0.38723f
C13356 a_31699_20742.t240 VSS 0.38723f
C13357 a_31699_20742.n308 VSS 2.74435f
C13358 a_31699_20742.n309 VSS 3.41548f
C13359 a_31699_20742.n310 VSS 2.37271f
C13360 a_31699_20742.n311 VSS 0.376149f
C13361 a_31699_20742.t87 VSS 0.38723f
C13362 a_31699_20742.t201 VSS 0.38723f
C13363 a_31699_20742.t73 VSS 0.38723f
C13364 a_31699_20742.t222 VSS 0.38723f
C13365 a_31699_20742.t147 VSS 0.38723f
C13366 a_31699_20742.t223 VSS 0.38723f
C13367 a_31699_20742.t51 VSS 0.38723f
C13368 a_31699_20742.t128 VSS 0.38723f
C13369 a_31699_20742.t162 VSS 0.38723f
C13370 a_31699_20742.t94 VSS 0.38723f
C13371 a_31699_20742.t75 VSS 0.38723f
C13372 a_31699_20742.n312 VSS 2.37271f
C13373 a_31699_20742.n313 VSS 16.538599f
C13374 a_31699_20742.t1 VSS 0.436569f
C13375 a_31699_20742.t33 VSS 0.41901f
C13376 a_31699_20742.n314 VSS 0.567026f
C13377 a_31699_20742.t7 VSS 0.419016f
C13378 a_31699_20742.n315 VSS 0.301485f
C13379 a_31699_20742.t37 VSS 0.419016f
C13380 a_31699_20742.n316 VSS 0.329307f
C13381 a_31699_20742.t185 VSS 0.419124f
C13382 a_31699_20742.n317 VSS 0.331307f
C13383 a_31699_20742.t256 VSS 0.419016f
C13384 a_31699_20742.n318 VSS 0.303598f
C13385 a_31699_20742.t89 VSS 0.419022f
C13386 a_31699_20742.n319 VSS 0.258958f
C13387 a_31699_20742.t27 VSS 0.436777f
C13388 a_31699_20742.t41 VSS 0.418993f
C13389 a_31699_20742.n320 VSS 0.570836f
C13390 a_31699_20742.t15 VSS 0.418993f
C13391 a_31699_20742.n321 VSS 0.301614f
C13392 a_31699_20742.t25 VSS 0.418993f
C13393 a_31699_20742.n322 VSS 0.305037f
C13394 a_31699_20742.n323 VSS 0.177663f
C13395 a_31699_20742.t131 VSS 0.436569f
C13396 a_31699_20742.t180 VSS 0.41901f
C13397 a_31699_20742.n324 VSS 0.567026f
C13398 a_31699_20742.t108 VSS 0.419016f
C13399 a_31699_20742.n325 VSS 0.301485f
C13400 a_31699_20742.t153 VSS 0.419016f
C13401 a_31699_20742.n326 VSS 0.329307f
C13402 a_31699_20742.t52 VSS 0.419124f
C13403 a_31699_20742.n327 VSS 0.331307f
C13404 a_31699_20742.t127 VSS 0.419016f
C13405 a_31699_20742.n328 VSS 0.303598f
C13406 a_31699_20742.t172 VSS 0.419022f
C13407 a_31699_20742.n329 VSS 0.258958f
C13408 a_31699_20742.t213 VSS 0.436777f
C13409 a_31699_20742.t138 VSS 0.418993f
C13410 a_31699_20742.n330 VSS 0.570836f
C13411 a_31699_20742.t72 VSS 0.418993f
C13412 a_31699_20742.n331 VSS 0.301614f
C13413 a_31699_20742.t218 VSS 0.418993f
C13414 a_31699_20742.n332 VSS 0.305037f
C13415 a_31699_20742.n333 VSS 0.099804f
C13416 a_31699_20742.n334 VSS 1.54854f
C13417 a_31699_20742.t220 VSS 0.439404f
C13418 a_31699_20742.t46 VSS 0.41901f
C13419 a_31699_20742.n335 VSS 0.609926f
C13420 a_31699_20742.t199 VSS 0.419016f
C13421 a_31699_20742.n336 VSS 0.301485f
C13422 a_31699_20742.t244 VSS 0.419016f
C13423 a_31699_20742.n337 VSS 0.329307f
C13424 a_31699_20742.t23 VSS 0.419124f
C13425 a_31699_20742.n338 VSS 0.331307f
C13426 a_31699_20742.t13 VSS 0.419016f
C13427 a_31699_20742.n339 VSS 0.303598f
C13428 a_31699_20742.t3 VSS 0.419022f
C13429 a_31699_20742.n340 VSS 0.258958f
C13430 a_31699_20742.t81 VSS 0.437037f
C13431 a_31699_20742.t234 VSS 0.418993f
C13432 a_31699_20742.n341 VSS 0.574774f
C13433 a_31699_20742.t163 VSS 0.418993f
C13434 a_31699_20742.n342 VSS 0.301614f
C13435 a_31699_20742.t92 VSS 0.418993f
C13436 a_31699_20742.n343 VSS 0.305037f
C13437 a_31699_20742.n344 VSS 0.099804f
C13438 a_31699_20742.n345 VSS 1.03208f
C13439 a_31699_20742.t60 VSS 0.436774f
C13440 a_31699_20742.t111 VSS 0.41901f
C13441 a_31699_20742.n346 VSS 0.570135f
C13442 a_31699_20742.t255 VSS 0.419016f
C13443 a_31699_20742.n347 VSS 0.301485f
C13444 a_31699_20742.t85 VSS 0.419016f
C13445 a_31699_20742.n348 VSS 0.329307f
C13446 a_31699_20742.t17 VSS 0.419124f
C13447 a_31699_20742.n349 VSS 0.331307f
C13448 a_31699_20742.t39 VSS 0.419016f
C13449 a_31699_20742.n350 VSS 0.303598f
C13450 a_31699_20742.t29 VSS 0.419022f
C13451 a_31699_20742.n351 VSS 0.258958f
C13452 a_31699_20742.t143 VSS 0.436572f
C13453 a_31699_20742.t71 VSS 0.418993f
C13454 a_31699_20742.n352 VSS 0.567727f
C13455 a_31699_20742.t226 VSS 0.418993f
C13456 a_31699_20742.n353 VSS 0.301614f
C13457 a_31699_20742.t150 VSS 0.418993f
C13458 a_31699_20742.n354 VSS 0.305037f
C13459 a_31699_20742.n355 VSS 0.099804f
C13460 a_31699_20742.t141 VSS 0.436569f
C13461 a_31699_20742.t192 VSS 0.41901f
C13462 a_31699_20742.n356 VSS 0.567026f
C13463 a_31699_20742.t118 VSS 0.419016f
C13464 a_31699_20742.n357 VSS 0.301485f
C13465 a_31699_20742.t164 VSS 0.419016f
C13466 a_31699_20742.n358 VSS 0.329307f
C13467 a_31699_20742.t62 VSS 0.419124f
C13468 a_31699_20742.n359 VSS 0.331307f
C13469 a_31699_20742.t134 VSS 0.419016f
C13470 a_31699_20742.n360 VSS 0.303598f
C13471 a_31699_20742.t184 VSS 0.419022f
C13472 a_31699_20742.n361 VSS 0.258958f
C13473 a_31699_20742.t224 VSS 0.436777f
C13474 a_31699_20742.t149 VSS 0.418993f
C13475 a_31699_20742.n362 VSS 0.570836f
C13476 a_31699_20742.t82 VSS 0.418993f
C13477 a_31699_20742.n363 VSS 0.301614f
C13478 a_31699_20742.t235 VSS 0.418993f
C13479 a_31699_20742.n364 VSS 0.305037f
C13480 a_31699_20742.n365 VSS 0.099804f
C13481 a_31699_20742.t43 VSS 0.38723f
C13482 a_31699_20742.n366 VSS 0.202043f
C13483 a_31699_20742.t11 VSS 0.395572f
C13484 a_31699_20742.n367 VSS 0.288798f
C13485 a_31699_20742.n368 VSS 0.193926f
C13486 a_31699_20742.n369 VSS 0.046177f
C13487 a_31699_20742.t19 VSS 0.38723f
C13488 a_31699_20742.t5 VSS 0.38723f
C13489 a_31699_20742.t144 VSS 0.419124f
C13490 a_31699_20742.n370 VSS 0.331512f
C13491 a_31699_20742.t219 VSS 0.419016f
C13492 a_31699_20742.n371 VSS 0.303598f
C13493 a_31699_20742.t45 VSS 0.419022f
C13494 a_31699_20742.n372 VSS 0.258958f
C13495 a_31699_20742.t31 VSS 0.38723f
C13496 a_31699_20742.n373 VSS 0.186798f
C13497 a_31699_20742.n374 VSS 0.049049f
C13498 a_31699_20742.t21 VSS 0.38723f
C13499 a_31699_20742.n375 VSS 0.046597f
C13500 a_31699_20742.t35 VSS 0.395626f
C13501 a_31699_20742.n376 VSS 0.289107f
C13502 a_31699_20742.t9 VSS 0.38723f
C13503 a_31699_20742.n377 VSS 0.20248f
C13504 a_31699_20742.n378 VSS 0.046597f
C13505 a_31699_20742.n379 VSS 0.180313f
C13506 a_31699_20742.n380 VSS 0.049049f
C13507 a_31699_20742.n381 VSS 0.027397f
C13508 a_31699_20742.n382 VSS 0.164642f
C13509 a_31699_20742.n383 VSS 0.046597f
C13510 a_31699_20742.n384 VSS 0.046597f
C13511 a_31699_20742.n385 VSS 0.058036f
C13512 a_31699_20742.n386 VSS 0.079208f
C13513 a_31699_20742.n387 VSS 0.092177f
C13514 a_31699_20742.n388 VSS 13.563499f
C13515 a_31699_20742.t0 VSS 1.11866f
C13516 a_31699_20742.n389 VSS 3.50557f
C13517 a_31699_20742.n390 VSS 2.18128f
C13518 a_31699_20742.t36 VSS 0.247033f
C13519 a_31699_20742.n391 VSS 0.184107f
C13520 a_31699_20742.t44 VSS 0.046398f
C13521 a_31953_n19727.n0 VSS 0.022916f
C13522 a_31953_n19727.n1 VSS 0.028194f
C13523 a_31953_n19727.n2 VSS 0.022916f
C13524 a_31953_n19727.n3 VSS 0.202509f
C13525 a_31953_n19727.n4 VSS 0.028194f
C13526 a_31953_n19727.n5 VSS 0.022916f
C13527 a_31953_n19727.n6 VSS 0.028194f
C13528 a_31953_n19727.n7 VSS 0.022916f
C13529 a_31953_n19727.n8 VSS 0.028194f
C13530 a_31953_n19727.n9 VSS 0.022916f
C13531 a_31953_n19727.n10 VSS 0.111389f
C13532 a_31953_n19727.n11 VSS 0.028194f
C13533 a_31953_n19727.n12 VSS 0.022916f
C13534 a_31953_n19727.n13 VSS 0.028194f
C13535 a_31953_n19727.n14 VSS 0.022914f
C13536 a_31953_n19727.n15 VSS 0.028194f
C13537 a_31953_n19727.n16 VSS 0.022916f
C13538 a_31953_n19727.n17 VSS 0.028194f
C13539 a_31953_n19727.n18 VSS 0.022916f
C13540 a_31953_n19727.n19 VSS 0.05571f
C13541 a_31953_n19727.n20 VSS 0.028194f
C13542 a_31953_n19727.n21 VSS 0.022914f
C13543 a_31953_n19727.n22 VSS 0.028194f
C13544 a_31953_n19727.n23 VSS 0.022916f
C13545 a_31953_n19727.n24 VSS 0.028194f
C13546 a_31953_n19727.n25 VSS 0.022916f
C13547 a_31953_n19727.n26 VSS 0.028194f
C13548 a_31953_n19727.n27 VSS 0.022916f
C13549 a_31953_n19727.n28 VSS 0.028194f
C13550 a_31953_n19727.n29 VSS 0.022916f
C13551 a_31953_n19727.n30 VSS 0.175142f
C13552 a_31953_n19727.n31 VSS 0.028194f
C13553 a_31953_n19727.n32 VSS 0.022914f
C13554 a_31953_n19727.n33 VSS 0.028194f
C13555 a_31953_n19727.n34 VSS 0.022916f
C13556 a_31953_n19727.n35 VSS 0.028194f
C13557 a_31953_n19727.n36 VSS 0.022916f
C13558 a_31953_n19727.n37 VSS 0.028194f
C13559 a_31953_n19727.n38 VSS 0.022916f
C13560 a_31953_n19727.n39 VSS 0.156168f
C13561 a_31953_n19727.n40 VSS 0.028194f
C13562 a_31953_n19727.n41 VSS 0.022916f
C13563 a_31953_n19727.n42 VSS 0.028194f
C13564 a_31953_n19727.n43 VSS 0.022916f
C13565 a_31953_n19727.n44 VSS 0.028194f
C13566 a_31953_n19727.n45 VSS 0.022916f
C13567 a_31953_n19727.n46 VSS 0.028194f
C13568 a_31953_n19727.n47 VSS 0.022916f
C13569 a_31953_n19727.n48 VSS 0.055679f
C13570 a_31953_n19727.n49 VSS 0.028194f
C13571 a_31953_n19727.n50 VSS 0.022914f
C13572 a_31953_n19727.n51 VSS 0.028194f
C13573 a_31953_n19727.n52 VSS 0.022916f
C13574 a_31953_n19727.n53 VSS 0.111389f
C13575 a_31953_n19727.n54 VSS 0.028194f
C13576 a_31953_n19727.n55 VSS 0.022916f
C13577 a_31953_n19727.n56 VSS 0.028194f
C13578 a_31953_n19727.n57 VSS 0.022914f
C13579 a_31953_n19727.n58 VSS 0.028194f
C13580 a_31953_n19727.n59 VSS 0.022916f
C13581 a_31953_n19727.n60 VSS 0.252146f
C13582 a_31953_n19727.n61 VSS 0.028194f
C13583 a_31953_n19727.n62 VSS 0.022916f
C13584 a_31953_n19727.n63 VSS 0.028194f
C13585 a_31953_n19727.n64 VSS 0.022916f
C13586 a_31953_n19727.n65 VSS 0.028194f
C13587 a_31953_n19727.n66 VSS 0.022916f
C13588 a_31953_n19727.n67 VSS 0.028194f
C13589 a_31953_n19727.n68 VSS 0.038388f
C13590 a_31953_n19727.n69 VSS 0.022916f
C13591 a_31953_n19727.n70 VSS 0.028194f
C13592 a_31953_n19727.n71 VSS 0.022916f
C13593 a_31953_n19727.n72 VSS 0.028194f
C13594 a_31953_n19727.n73 VSS 0.022916f
C13595 a_31953_n19727.n74 VSS 0.202509f
C13596 a_31953_n19727.n75 VSS 0.028194f
C13597 a_31953_n19727.n76 VSS 0.022916f
C13598 a_31953_n19727.n77 VSS 0.028194f
C13599 a_31953_n19727.n78 VSS 0.022916f
C13600 a_31953_n19727.n79 VSS 0.028194f
C13601 a_31953_n19727.n80 VSS 0.022916f
C13602 a_31953_n19727.n81 VSS 0.111389f
C13603 a_31953_n19727.n82 VSS 0.028194f
C13604 a_31953_n19727.n83 VSS 0.022916f
C13605 a_31953_n19727.n84 VSS 0.028194f
C13606 a_31953_n19727.n85 VSS 0.022914f
C13607 a_31953_n19727.n86 VSS 0.028194f
C13608 a_31953_n19727.n87 VSS 0.022916f
C13609 a_31953_n19727.n88 VSS 0.028194f
C13610 a_31953_n19727.n89 VSS 0.022916f
C13611 a_31953_n19727.n90 VSS 0.05571f
C13612 a_31953_n19727.n91 VSS 0.028194f
C13613 a_31953_n19727.n92 VSS 0.022914f
C13614 a_31953_n19727.n93 VSS 0.028194f
C13615 a_31953_n19727.n94 VSS 0.022916f
C13616 a_31953_n19727.n95 VSS 0.028194f
C13617 a_31953_n19727.n96 VSS 0.022916f
C13618 a_31953_n19727.n97 VSS 0.028194f
C13619 a_31953_n19727.n98 VSS 0.022916f
C13620 a_31953_n19727.n99 VSS 0.028194f
C13621 a_31953_n19727.n100 VSS 0.022916f
C13622 a_31953_n19727.n101 VSS 0.174613f
C13623 a_31953_n19727.n102 VSS 0.028194f
C13624 a_31953_n19727.n103 VSS 0.022914f
C13625 a_31953_n19727.n104 VSS 0.028194f
C13626 a_31953_n19727.n105 VSS 0.022916f
C13627 a_31953_n19727.n106 VSS 0.028194f
C13628 a_31953_n19727.n107 VSS 0.022916f
C13629 a_31953_n19727.n108 VSS 0.154833f
C13630 a_31953_n19727.n109 VSS 0.028194f
C13631 a_31953_n19727.n110 VSS 0.022916f
C13632 a_31953_n19727.n111 VSS 0.028194f
C13633 a_31953_n19727.n112 VSS 0.022916f
C13634 a_31953_n19727.n113 VSS 0.055679f
C13635 a_31953_n19727.n114 VSS 0.028194f
C13636 a_31953_n19727.n115 VSS 0.022916f
C13637 a_31953_n19727.n116 VSS 0.028194f
C13638 a_31953_n19727.n117 VSS 0.022916f
C13639 a_31953_n19727.n118 VSS 0.028194f
C13640 a_31953_n19727.n119 VSS 0.022916f
C13641 a_31953_n19727.n120 VSS 0.028194f
C13642 a_31953_n19727.n121 VSS 0.022914f
C13643 a_31953_n19727.n122 VSS 0.028194f
C13644 a_31953_n19727.n123 VSS 0.022916f
C13645 a_31953_n19727.n124 VSS 0.111389f
C13646 a_31953_n19727.n125 VSS 0.028194f
C13647 a_31953_n19727.n126 VSS 0.022916f
C13648 a_31953_n19727.n127 VSS 0.028194f
C13649 a_31953_n19727.n128 VSS 0.022914f
C13650 a_31953_n19727.n129 VSS 0.028194f
C13651 a_31953_n19727.n130 VSS 0.022916f
C13652 a_31953_n19727.n131 VSS 0.252146f
C13653 a_31953_n19727.n132 VSS 0.028194f
C13654 a_31953_n19727.n133 VSS 0.022916f
C13655 a_31953_n19727.n134 VSS 0.028194f
C13656 a_31953_n19727.n135 VSS 0.022916f
C13657 a_31953_n19727.n136 VSS 0.028194f
C13658 a_31953_n19727.n137 VSS 0.022916f
C13659 a_31953_n19727.n138 VSS 0.028194f
C13660 a_31953_n19727.n139 VSS 0.038388f
C13661 a_31953_n19727.n140 VSS 0.022916f
C13662 a_31953_n19727.n141 VSS 0.028194f
C13663 a_31953_n19727.n142 VSS 0.022916f
C13664 a_31953_n19727.n143 VSS 0.028194f
C13665 a_31953_n19727.n144 VSS 0.022916f
C13666 a_31953_n19727.n145 VSS 0.202509f
C13667 a_31953_n19727.n146 VSS 0.028194f
C13668 a_31953_n19727.n147 VSS 0.022916f
C13669 a_31953_n19727.n148 VSS 0.028194f
C13670 a_31953_n19727.n149 VSS 0.022916f
C13671 a_31953_n19727.n150 VSS 0.028194f
C13672 a_31953_n19727.n151 VSS 0.022916f
C13673 a_31953_n19727.n152 VSS 0.111389f
C13674 a_31953_n19727.n153 VSS 0.028194f
C13675 a_31953_n19727.n154 VSS 0.022916f
C13676 a_31953_n19727.n155 VSS 0.028194f
C13677 a_31953_n19727.n156 VSS 0.022914f
C13678 a_31953_n19727.n157 VSS 0.028194f
C13679 a_31953_n19727.n158 VSS 0.022916f
C13680 a_31953_n19727.n159 VSS 0.028194f
C13681 a_31953_n19727.n160 VSS 0.022916f
C13682 a_31953_n19727.n161 VSS 0.05571f
C13683 a_31953_n19727.n162 VSS 0.028194f
C13684 a_31953_n19727.n163 VSS 0.022914f
C13685 a_31953_n19727.n164 VSS 0.028194f
C13686 a_31953_n19727.n165 VSS 0.022916f
C13687 a_31953_n19727.n166 VSS 0.028194f
C13688 a_31953_n19727.n167 VSS 0.022916f
C13689 a_31953_n19727.n168 VSS 0.028194f
C13690 a_31953_n19727.n169 VSS 0.022916f
C13691 a_31953_n19727.n170 VSS 0.028194f
C13692 a_31953_n19727.n171 VSS 0.022916f
C13693 a_31953_n19727.n172 VSS 0.175142f
C13694 a_31953_n19727.n173 VSS 0.028194f
C13695 a_31953_n19727.n174 VSS 0.022914f
C13696 a_31953_n19727.n175 VSS 0.028194f
C13697 a_31953_n19727.n176 VSS 0.022916f
C13698 a_31953_n19727.n177 VSS 0.028194f
C13699 a_31953_n19727.n178 VSS 0.022916f
C13700 a_31953_n19727.n179 VSS 0.156168f
C13701 a_31953_n19727.n180 VSS 0.028194f
C13702 a_31953_n19727.n181 VSS 0.022916f
C13703 a_31953_n19727.n182 VSS 0.028194f
C13704 a_31953_n19727.n183 VSS 0.022916f
C13705 a_31953_n19727.n184 VSS 0.055679f
C13706 a_31953_n19727.n185 VSS 0.028194f
C13707 a_31953_n19727.n186 VSS 0.022916f
C13708 a_31953_n19727.n187 VSS 0.028194f
C13709 a_31953_n19727.n188 VSS 0.022916f
C13710 a_31953_n19727.n189 VSS 0.028194f
C13711 a_31953_n19727.n190 VSS 0.022916f
C13712 a_31953_n19727.n191 VSS 0.028194f
C13713 a_31953_n19727.n192 VSS 0.022914f
C13714 a_31953_n19727.n193 VSS 0.028194f
C13715 a_31953_n19727.n194 VSS 0.022916f
C13716 a_31953_n19727.n195 VSS 0.111389f
C13717 a_31953_n19727.n196 VSS 0.028194f
C13718 a_31953_n19727.n197 VSS 0.022916f
C13719 a_31953_n19727.n198 VSS 0.028194f
C13720 a_31953_n19727.n199 VSS 0.022914f
C13721 a_31953_n19727.n200 VSS 0.028194f
C13722 a_31953_n19727.n201 VSS 0.022916f
C13723 a_31953_n19727.n202 VSS 0.252146f
C13724 a_31953_n19727.n203 VSS 0.028194f
C13725 a_31953_n19727.n204 VSS 0.022916f
C13726 a_31953_n19727.n205 VSS 0.028194f
C13727 a_31953_n19727.n206 VSS 0.022916f
C13728 a_31953_n19727.n207 VSS 0.028194f
C13729 a_31953_n19727.n208 VSS 0.022916f
C13730 a_31953_n19727.n209 VSS 0.028194f
C13731 a_31953_n19727.n210 VSS 0.038388f
C13732 a_31953_n19727.n211 VSS 0.022916f
C13733 a_31953_n19727.n212 VSS 0.028194f
C13734 a_31953_n19727.n213 VSS 0.023381f
C13735 a_31953_n19727.n214 VSS 0.032827f
C13736 a_31953_n19727.n215 VSS 0.023381f
C13737 a_31953_n19727.n216 VSS 0.028924f
C13738 a_31953_n19727.n217 VSS 0.023381f
C13739 a_31953_n19727.n218 VSS 0.032827f
C13740 a_31953_n19727.n219 VSS 0.023381f
C13741 a_31953_n19727.n220 VSS 0.028924f
C13742 a_31953_n19727.n221 VSS 0.023381f
C13743 a_31953_n19727.n222 VSS 0.032827f
C13744 a_31953_n19727.n223 VSS 0.023381f
C13745 a_31953_n19727.n224 VSS 0.028924f
C13746 a_31953_n19727.n225 VSS 0.17012f
C13747 a_31953_n19727.n226 VSS 0.710578f
C13748 a_31953_n19727.t13 VSS 0.007658f
C13749 a_31953_n19727.n227 VSS 0.016885f
C13750 a_31953_n19727.t19 VSS 0.007658f
C13751 a_31953_n19727.n228 VSS 0.021674f
C13752 a_31953_n19727.t21 VSS 0.007658f
C13753 a_31953_n19727.n229 VSS 0.022051f
C13754 a_31953_n19727.t17 VSS 0.007658f
C13755 a_31953_n19727.n230 VSS 0.016885f
C13756 a_31953_n19727.t39 VSS 0.007658f
C13757 a_31953_n19727.n231 VSS 0.022107f
C13758 a_31953_n19727.n232 VSS 0.046928f
C13759 a_31953_n19727.t99 VSS 0.042575f
C13760 a_31953_n19727.t195 VSS 0.039952f
C13761 a_31953_n19727.n233 VSS 0.04589f
C13762 a_31953_n19727.t100 VSS 0.039952f
C13763 a_31953_n19727.t208 VSS 0.039952f
C13764 a_31953_n19727.n234 VSS 0.046902f
C13765 a_31953_n19727.t197 VSS 0.042571f
C13766 a_31953_n19727.n235 VSS 0.045866f
C13767 a_31953_n19727.n236 VSS 0.025554f
C13768 a_31953_n19727.n237 VSS 0.025366f
C13769 a_31953_n19727.t273 VSS 0.039919f
C13770 a_31953_n19727.n238 VSS 0.045891f
C13771 a_31953_n19727.t174 VSS 0.042606f
C13772 a_31953_n19727.t271 VSS 0.039948f
C13773 a_31953_n19727.n239 VSS 0.045891f
C13774 a_31953_n19727.t175 VSS 0.039948f
C13775 a_31953_n19727.t281 VSS 0.039948f
C13776 a_31953_n19727.n240 VSS 0.045866f
C13777 a_31953_n19727.t276 VSS 0.042602f
C13778 a_31953_n19727.n241 VSS 0.045866f
C13779 a_31953_n19727.t345 VSS 0.039948f
C13780 a_31953_n19727.n242 VSS 0.045891f
C13781 a_31953_n19727.t159 VSS 0.042606f
C13782 a_31953_n19727.t259 VSS 0.039948f
C13783 a_31953_n19727.n243 VSS 0.045891f
C13784 a_31953_n19727.t160 VSS 0.039948f
C13785 a_31953_n19727.t270 VSS 0.039948f
C13786 a_31953_n19727.n244 VSS 0.045866f
C13787 a_31953_n19727.t262 VSS 0.042602f
C13788 a_31953_n19727.n245 VSS 0.045866f
C13789 a_31953_n19727.t329 VSS 0.039948f
C13790 a_31953_n19727.n246 VSS 0.045891f
C13791 a_31953_n19727.t299 VSS 0.042606f
C13792 a_31953_n19727.t95 VSS 0.039948f
C13793 a_31953_n19727.n247 VSS 0.045891f
C13794 a_31953_n19727.t20 VSS 0.039948f
C13795 a_31953_n19727.t111 VSS 0.039903f
C13796 a_31953_n19727.n248 VSS 0.04561f
C13797 a_31953_n19727.t102 VSS 0.042602f
C13798 a_31953_n19727.n249 VSS 0.045866f
C13799 a_31953_n19727.t52 VSS 0.039948f
C13800 a_31953_n19727.n250 VSS 0.045891f
C13801 a_31953_n19727.t311 VSS 0.042606f
C13802 a_31953_n19727.t112 VSS 0.039948f
C13803 a_31953_n19727.n251 VSS 0.045891f
C13804 a_31953_n19727.t16 VSS 0.039948f
C13805 a_31953_n19727.t121 VSS 0.039901f
C13806 a_31953_n19727.n252 VSS 0.045866f
C13807 a_31953_n19727.t117 VSS 0.042602f
C13808 a_31953_n19727.n253 VSS 0.045597f
C13809 a_31953_n19727.t48 VSS 0.039948f
C13810 a_31953_n19727.n254 VSS 0.045891f
C13811 a_31953_n19727.t238 VSS 0.042606f
C13812 a_31953_n19727.t327 VSS 0.039948f
C13813 a_31953_n19727.n255 VSS 0.045891f
C13814 a_31953_n19727.t38 VSS 0.039948f
C13815 a_31953_n19727.t342 VSS 0.039948f
C13816 a_31953_n19727.n256 VSS 0.045866f
C13817 a_31953_n19727.t333 VSS 0.042602f
C13818 a_31953_n19727.n257 VSS 0.045866f
C13819 a_31953_n19727.t60 VSS 0.039948f
C13820 a_31953_n19727.n258 VSS 0.024552f
C13821 a_31953_n19727.t61 VSS 0.007658f
C13822 a_31953_n19727.n259 VSS 0.021693f
C13823 a_31953_n19727.t49 VSS 0.007658f
C13824 a_31953_n19727.n260 VSS 0.016885f
C13825 a_31953_n19727.t53 VSS 0.007658f
C13826 a_31953_n19727.n261 VSS 0.021674f
C13827 a_31953_n19727.n262 VSS 0.024376f
C13828 a_31953_n19727.n263 VSS 0.045891f
C13829 a_31953_n19727.t78 VSS 0.042606f
C13830 a_31953_n19727.t170 VSS 0.039948f
C13831 a_31953_n19727.n264 VSS 0.045891f
C13832 a_31953_n19727.t79 VSS 0.039948f
C13833 a_31953_n19727.t186 VSS 0.039948f
C13834 a_31953_n19727.n265 VSS 0.045866f
C13835 a_31953_n19727.t177 VSS 0.042602f
C13836 a_31953_n19727.n266 VSS 0.045866f
C13837 a_31953_n19727.t250 VSS 0.039948f
C13838 a_31953_n19727.n267 VSS 0.045891f
C13839 a_31953_n19727.t146 VSS 0.042606f
C13840 a_31953_n19727.t248 VSS 0.039948f
C13841 a_31953_n19727.n268 VSS 0.045891f
C13842 a_31953_n19727.t149 VSS 0.039948f
C13843 a_31953_n19727.t261 VSS 0.039948f
C13844 a_31953_n19727.n269 VSS 0.045866f
C13845 a_31953_n19727.t253 VSS 0.042602f
C13846 a_31953_n19727.n270 VSS 0.045866f
C13847 a_31953_n19727.t319 VSS 0.039948f
C13848 a_31953_n19727.n271 VSS 0.045891f
C13849 a_31953_n19727.t128 VSS 0.042606f
C13850 a_31953_n19727.t221 VSS 0.039948f
C13851 a_31953_n19727.n272 VSS 0.045891f
C13852 a_31953_n19727.t129 VSS 0.039948f
C13853 a_31953_n19727.t229 VSS 0.039898f
C13854 a_31953_n19727.n273 VSS 0.045583f
C13855 a_31953_n19727.t224 VSS 0.042602f
C13856 a_31953_n19727.n274 VSS 0.045866f
C13857 a_31953_n19727.t295 VSS 0.039948f
C13858 a_31953_n19727.t69 VSS 0.007658f
C13859 a_31953_n19727.n275 VSS 0.022051f
C13860 a_31953_n19727.t65 VSS 0.007658f
C13861 a_31953_n19727.n276 VSS 0.016885f
C13862 a_31953_n19727.t15 VSS 0.007658f
C13863 a_31953_n19727.n277 VSS 0.022107f
C13864 a_31953_n19727.n278 VSS 0.046928f
C13865 a_31953_n19727.t180 VSS 0.042575f
C13866 a_31953_n19727.t275 VSS 0.039952f
C13867 a_31953_n19727.n279 VSS 0.04589f
C13868 a_31953_n19727.t181 VSS 0.039952f
C13869 a_31953_n19727.t286 VSS 0.039952f
C13870 a_31953_n19727.n280 VSS 0.046902f
C13871 a_31953_n19727.t114 VSS 0.042571f
C13872 a_31953_n19727.n281 VSS 0.045866f
C13873 a_31953_n19727.n282 VSS 0.025554f
C13874 a_31953_n19727.n283 VSS 0.025366f
C13875 a_31953_n19727.t187 VSS 0.039919f
C13876 a_31953_n19727.n284 VSS 0.045891f
C13877 a_31953_n19727.t255 VSS 0.042606f
C13878 a_31953_n19727.t347 VSS 0.039948f
C13879 a_31953_n19727.n285 VSS 0.045891f
C13880 a_31953_n19727.t256 VSS 0.039948f
C13881 a_31953_n19727.t357 VSS 0.039948f
C13882 a_31953_n19727.n286 VSS 0.045866f
C13883 a_31953_n19727.t189 VSS 0.042602f
C13884 a_31953_n19727.n287 VSS 0.045866f
C13885 a_31953_n19727.t264 VSS 0.039948f
C13886 a_31953_n19727.n288 VSS 0.045891f
C13887 a_31953_n19727.t240 VSS 0.042606f
C13888 a_31953_n19727.t331 VSS 0.039948f
C13889 a_31953_n19727.n289 VSS 0.045891f
C13890 a_31953_n19727.t242 VSS 0.039948f
C13891 a_31953_n19727.t343 VSS 0.039948f
C13892 a_31953_n19727.n290 VSS 0.045866f
C13893 a_31953_n19727.t172 VSS 0.042602f
C13894 a_31953_n19727.n291 VSS 0.045866f
C13895 a_31953_n19727.t249 VSS 0.039948f
C13896 a_31953_n19727.n292 VSS 0.045891f
C13897 a_31953_n19727.t81 VSS 0.042606f
C13898 a_31953_n19727.t173 VSS 0.039948f
C13899 a_31953_n19727.n293 VSS 0.045891f
C13900 a_31953_n19727.t68 VSS 0.039948f
C13901 a_31953_n19727.t188 VSS 0.039903f
C13902 a_31953_n19727.n294 VSS 0.04561f
C13903 a_31953_n19727.t310 VSS 0.042602f
C13904 a_31953_n19727.n295 VSS 0.045866f
C13905 a_31953_n19727.t66 VSS 0.039948f
C13906 a_31953_n19727.n296 VSS 0.045891f
C13907 a_31953_n19727.t91 VSS 0.042606f
C13908 a_31953_n19727.t191 VSS 0.039948f
C13909 a_31953_n19727.n297 VSS 0.045891f
C13910 a_31953_n19727.t64 VSS 0.039948f
C13911 a_31953_n19727.t201 VSS 0.039901f
C13912 a_31953_n19727.n298 VSS 0.045866f
C13913 a_31953_n19727.t320 VSS 0.042602f
C13914 a_31953_n19727.n299 VSS 0.045597f
C13915 a_31953_n19727.t62 VSS 0.039948f
C13916 a_31953_n19727.n300 VSS 0.045891f
C13917 a_31953_n19727.t312 VSS 0.042606f
C13918 a_31953_n19727.t116 VSS 0.039948f
C13919 a_31953_n19727.n301 VSS 0.045891f
C13920 a_31953_n19727.t14 VSS 0.039948f
C13921 a_31953_n19727.t124 VSS 0.039948f
C13922 a_31953_n19727.n302 VSS 0.045866f
C13923 a_31953_n19727.t251 VSS 0.042602f
C13924 a_31953_n19727.n303 VSS 0.045866f
C13925 a_31953_n19727.t10 VSS 0.039948f
C13926 a_31953_n19727.n304 VSS 0.024552f
C13927 a_31953_n19727.t11 VSS 0.007658f
C13928 a_31953_n19727.n305 VSS 0.021693f
C13929 a_31953_n19727.t63 VSS 0.007658f
C13930 a_31953_n19727.n306 VSS 0.016885f
C13931 a_31953_n19727.t67 VSS 0.007658f
C13932 a_31953_n19727.n307 VSS 0.021674f
C13933 a_31953_n19727.n308 VSS 0.024376f
C13934 a_31953_n19727.n309 VSS 0.045891f
C13935 a_31953_n19727.t151 VSS 0.042606f
C13936 a_31953_n19727.t252 VSS 0.039948f
C13937 a_31953_n19727.n310 VSS 0.045891f
C13938 a_31953_n19727.t153 VSS 0.039948f
C13939 a_31953_n19727.t265 VSS 0.039948f
C13940 a_31953_n19727.n311 VSS 0.045866f
C13941 a_31953_n19727.t89 VSS 0.042602f
C13942 a_31953_n19727.n312 VSS 0.045866f
C13943 a_31953_n19727.t163 VSS 0.039948f
C13944 a_31953_n19727.n313 VSS 0.045891f
C13945 a_31953_n19727.t231 VSS 0.042606f
C13946 a_31953_n19727.t321 VSS 0.039948f
C13947 a_31953_n19727.n314 VSS 0.045891f
C13948 a_31953_n19727.t232 VSS 0.039948f
C13949 a_31953_n19727.t335 VSS 0.039948f
C13950 a_31953_n19727.n315 VSS 0.045866f
C13951 a_31953_n19727.t164 VSS 0.042602f
C13952 a_31953_n19727.n316 VSS 0.045866f
C13953 a_31953_n19727.t241 VSS 0.039948f
C13954 a_31953_n19727.n317 VSS 0.045891f
C13955 a_31953_n19727.t210 VSS 0.042606f
C13956 a_31953_n19727.t297 VSS 0.039948f
C13957 a_31953_n19727.n318 VSS 0.045891f
C13958 a_31953_n19727.t211 VSS 0.039948f
C13959 a_31953_n19727.t306 VSS 0.039898f
C13960 a_31953_n19727.n319 VSS 0.045583f
C13961 a_31953_n19727.t139 VSS 0.042602f
C13962 a_31953_n19727.n320 VSS 0.045866f
C13963 a_31953_n19727.t216 VSS 0.039948f
C13964 a_31953_n19727.t72 VSS 0.073404f
C13965 a_31953_n19727.t73 VSS 0.061873f
C13966 a_31953_n19727.n321 VSS 1.21075f
C13967 a_31953_n19727.t59 VSS 0.007658f
C13968 a_31953_n19727.n322 VSS 0.022107f
C13969 a_31953_n19727.t43 VSS 0.007658f
C13970 a_31953_n19727.n323 VSS 0.016885f
C13971 a_31953_n19727.t31 VSS 0.007658f
C13972 a_31953_n19727.n324 VSS 0.022051f
C13973 a_31953_n19727.n325 VSS 0.045891f
C13974 a_31953_n19727.t266 VSS 0.042606f
C13975 a_31953_n19727.t156 VSS 0.039948f
C13976 a_31953_n19727.n326 VSS 0.045891f
C13977 a_31953_n19727.t58 VSS 0.039948f
C13978 a_31953_n19727.t82 VSS 0.039948f
C13979 a_31953_n19727.n327 VSS 0.045866f
C13980 a_31953_n19727.t145 VSS 0.042602f
C13981 a_31953_n19727.n328 VSS 0.045866f
C13982 a_31953_n19727.t44 VSS 0.039948f
C13983 a_31953_n19727.n329 VSS 0.045891f
C13984 a_31953_n19727.t336 VSS 0.042606f
C13985 a_31953_n19727.t236 VSS 0.039948f
C13986 a_31953_n19727.n330 VSS 0.045891f
C13987 a_31953_n19727.t42 VSS 0.039948f
C13988 a_31953_n19727.t154 VSS 0.039901f
C13989 a_31953_n19727.n331 VSS 0.045597f
C13990 a_31953_n19727.t226 VSS 0.042602f
C13991 a_31953_n19727.n332 VSS 0.045866f
C13992 a_31953_n19727.t24 VSS 0.039948f
C13993 a_31953_n19727.n333 VSS 0.045891f
C13994 a_31953_n19727.t103 VSS 0.042606f
C13995 a_31953_n19727.t294 VSS 0.039948f
C13996 a_31953_n19727.n334 VSS 0.045891f
C13997 a_31953_n19727.t30 VSS 0.039948f
C13998 a_31953_n19727.t219 VSS 0.039903f
C13999 a_31953_n19727.n335 VSS 0.045866f
C14000 a_31953_n19727.t288 VSS 0.042602f
C14001 a_31953_n19727.n336 VSS 0.04561f
C14002 a_31953_n19727.t8 VSS 0.039948f
C14003 a_31953_n19727.t167 VSS 0.039948f
C14004 a_31953_n19727.t133 VSS 0.039898f
C14005 a_31953_n19727.n337 VSS 0.022914f
C14006 a_31953_n19727.n338 VSS 0.045583f
C14007 a_31953_n19727.t202 VSS 0.042602f
C14008 a_31953_n19727.n339 VSS 0.045866f
C14009 a_31953_n19727.n340 VSS 0.045891f
C14010 a_31953_n19727.t309 VSS 0.042606f
C14011 a_31953_n19727.t213 VSS 0.039948f
C14012 a_31953_n19727.n341 VSS 0.045891f
C14013 a_31953_n19727.t239 VSS 0.039948f
C14014 a_31953_n19727.n342 VSS 0.045891f
C14015 a_31953_n19727.t235 VSS 0.042606f
C14016 a_31953_n19727.t134 VSS 0.039948f
C14017 a_31953_n19727.n343 VSS 0.045891f
C14018 a_31953_n19727.t93 VSS 0.039948f
C14019 a_31953_n19727.t352 VSS 0.039948f
C14020 a_31953_n19727.n344 VSS 0.045866f
C14021 a_31953_n19727.t125 VSS 0.042602f
C14022 a_31953_n19727.n345 VSS 0.045866f
C14023 a_31953_n19727.t162 VSS 0.039948f
C14024 a_31953_n19727.n346 VSS 0.045891f
C14025 a_31953_n19727.t179 VSS 0.042606f
C14026 a_31953_n19727.t75 VSS 0.039948f
C14027 a_31953_n19727.n347 VSS 0.045891f
C14028 a_31953_n19727.t332 VSS 0.039948f
C14029 a_31953_n19727.t291 VSS 0.039948f
C14030 a_31953_n19727.n348 VSS 0.045866f
C14031 a_31953_n19727.t359 VSS 0.042602f
C14032 a_31953_n19727.n349 VSS 0.045866f
C14033 a_31953_n19727.t105 VSS 0.039948f
C14034 a_31953_n19727.n350 VSS 0.024376f
C14035 a_31953_n19727.t9 VSS 0.007658f
C14036 a_31953_n19727.n351 VSS 0.021674f
C14037 a_31953_n19727.t25 VSS 0.007658f
C14038 a_31953_n19727.n352 VSS 0.016885f
C14039 a_31953_n19727.t45 VSS 0.007658f
C14040 a_31953_n19727.n353 VSS 0.021693f
C14041 a_31953_n19727.n354 VSS 0.024552f
C14042 a_31953_n19727.n355 VSS 0.045891f
C14043 a_31953_n19727.t279 VSS 0.042606f
C14044 a_31953_n19727.t171 VSS 0.039948f
C14045 a_31953_n19727.n356 VSS 0.045891f
C14046 a_31953_n19727.t136 VSS 0.039948f
C14047 a_31953_n19727.t92 VSS 0.039948f
C14048 a_31953_n19727.n357 VSS 0.045866f
C14049 a_31953_n19727.t161 VSS 0.042602f
C14050 a_31953_n19727.n358 VSS 0.045866f
C14051 a_31953_n19727.t206 VSS 0.039948f
C14052 a_31953_n19727.n359 VSS 0.045891f
C14053 a_31953_n19727.t203 VSS 0.042606f
C14054 a_31953_n19727.t96 VSS 0.039948f
C14055 a_31953_n19727.n360 VSS 0.045891f
C14056 a_31953_n19727.t353 VSS 0.039948f
C14057 a_31953_n19727.t313 VSS 0.039948f
C14058 a_31953_n19727.n361 VSS 0.045866f
C14059 a_31953_n19727.t87 VSS 0.042602f
C14060 a_31953_n19727.n362 VSS 0.045866f
C14061 a_31953_n19727.t131 VSS 0.039948f
C14062 a_31953_n19727.n363 VSS 0.046928f
C14063 a_31953_n19727.t126 VSS 0.042575f
C14064 a_31953_n19727.t315 VSS 0.039952f
C14065 a_31953_n19727.n364 VSS 0.04589f
C14066 a_31953_n19727.t283 VSS 0.039952f
C14067 a_31953_n19727.t243 VSS 0.039952f
C14068 a_31953_n19727.n365 VSS 0.046902f
C14069 a_31953_n19727.t305 VSS 0.042571f
C14070 a_31953_n19727.n366 VSS 0.045866f
C14071 a_31953_n19727.n367 VSS 0.025554f
C14072 a_31953_n19727.n368 VSS 0.025366f
C14073 a_31953_n19727.t350 VSS 0.039919f
C14074 a_31953_n19727.t33 VSS 0.007658f
C14075 a_31953_n19727.n369 VSS 0.022051f
C14076 a_31953_n19727.t29 VSS 0.007658f
C14077 a_31953_n19727.n370 VSS 0.016885f
C14078 a_31953_n19727.t47 VSS 0.007658f
C14079 a_31953_n19727.n371 VSS 0.022107f
C14080 a_31953_n19727.n372 VSS 0.046928f
C14081 a_31953_n19727.t293 VSS 0.042575f
C14082 a_31953_n19727.t316 VSS 0.039952f
C14083 a_31953_n19727.n373 VSS 0.04589f
C14084 a_31953_n19727.t348 VSS 0.039952f
C14085 a_31953_n19727.t132 VSS 0.039952f
C14086 a_31953_n19727.n374 VSS 0.046902f
C14087 a_31953_n19727.t258 VSS 0.042571f
C14088 a_31953_n19727.n375 VSS 0.045866f
C14089 a_31953_n19727.n376 VSS 0.025554f
C14090 a_31953_n19727.n377 VSS 0.025366f
C14091 a_31953_n19727.t130 VSS 0.039919f
C14092 a_31953_n19727.n378 VSS 0.045891f
C14093 a_31953_n19727.t74 VSS 0.042606f
C14094 a_31953_n19727.t97 VSS 0.039948f
C14095 a_31953_n19727.n379 VSS 0.045891f
C14096 a_31953_n19727.t127 VSS 0.039948f
C14097 a_31953_n19727.t207 VSS 0.039948f
C14098 a_31953_n19727.n380 VSS 0.045866f
C14099 a_31953_n19727.t326 VSS 0.042602f
C14100 a_31953_n19727.n381 VSS 0.045866f
C14101 a_31953_n19727.t205 VSS 0.039948f
C14102 a_31953_n19727.n382 VSS 0.045891f
C14103 a_31953_n19727.t356 VSS 0.042606f
C14104 a_31953_n19727.t85 VSS 0.039948f
C14105 a_31953_n19727.n383 VSS 0.045891f
C14106 a_31953_n19727.t118 VSS 0.039948f
C14107 a_31953_n19727.t194 VSS 0.039948f
C14108 a_31953_n19727.n384 VSS 0.045866f
C14109 a_31953_n19727.t314 VSS 0.042602f
C14110 a_31953_n19727.n385 VSS 0.045866f
C14111 a_31953_n19727.t192 VSS 0.039948f
C14112 a_31953_n19727.n386 VSS 0.045891f
C14113 a_31953_n19727.t200 VSS 0.042606f
C14114 a_31953_n19727.t225 VSS 0.039948f
C14115 a_31953_n19727.n387 VSS 0.045891f
C14116 a_31953_n19727.t32 VSS 0.039948f
C14117 a_31953_n19727.t324 VSS 0.039903f
C14118 a_31953_n19727.n388 VSS 0.04561f
C14119 a_31953_n19727.t155 VSS 0.042602f
C14120 a_31953_n19727.n389 VSS 0.045866f
C14121 a_31953_n19727.t6 VSS 0.039948f
C14122 a_31953_n19727.n390 VSS 0.045891f
C14123 a_31953_n19727.t215 VSS 0.042606f
C14124 a_31953_n19727.t237 VSS 0.039948f
C14125 a_31953_n19727.n391 VSS 0.045891f
C14126 a_31953_n19727.t28 VSS 0.039948f
C14127 a_31953_n19727.t341 VSS 0.039901f
C14128 a_31953_n19727.n392 VSS 0.045866f
C14129 a_31953_n19727.t168 VSS 0.042602f
C14130 a_31953_n19727.n393 VSS 0.045597f
C14131 a_31953_n19727.t4 VSS 0.039948f
C14132 a_31953_n19727.n394 VSS 0.045891f
C14133 a_31953_n19727.t138 VSS 0.042606f
C14134 a_31953_n19727.t157 VSS 0.039948f
C14135 a_31953_n19727.n395 VSS 0.045891f
C14136 a_31953_n19727.t46 VSS 0.039948f
C14137 a_31953_n19727.t269 VSS 0.039948f
C14138 a_31953_n19727.n396 VSS 0.045866f
C14139 a_31953_n19727.t94 VSS 0.042602f
C14140 a_31953_n19727.n397 VSS 0.045866f
C14141 a_31953_n19727.t26 VSS 0.039948f
C14142 a_31953_n19727.n398 VSS 0.024552f
C14143 a_31953_n19727.t27 VSS 0.007658f
C14144 a_31953_n19727.n399 VSS 0.021693f
C14145 a_31953_n19727.t5 VSS 0.007658f
C14146 a_31953_n19727.n400 VSS 0.016885f
C14147 a_31953_n19727.t7 VSS 0.007658f
C14148 a_31953_n19727.n401 VSS 0.021674f
C14149 a_31953_n19727.n402 VSS 0.024376f
C14150 a_31953_n19727.n403 VSS 0.045891f
C14151 a_31953_n19727.t278 VSS 0.042606f
C14152 a_31953_n19727.t298 VSS 0.039948f
C14153 a_31953_n19727.n404 VSS 0.045891f
C14154 a_31953_n19727.t322 VSS 0.039948f
C14155 a_31953_n19727.t109 VSS 0.039948f
C14156 a_31953_n19727.n405 VSS 0.045866f
C14157 a_31953_n19727.t234 VSS 0.042602f
C14158 a_31953_n19727.n406 VSS 0.045866f
C14159 a_31953_n19727.t107 VSS 0.039948f
C14160 a_31953_n19727.n407 VSS 0.045891f
C14161 a_31953_n19727.t351 VSS 0.042606f
C14162 a_31953_n19727.t77 VSS 0.039948f
C14163 a_31953_n19727.n408 VSS 0.045891f
C14164 a_31953_n19727.t106 VSS 0.039948f
C14165 a_31953_n19727.t185 VSS 0.039948f
C14166 a_31953_n19727.n409 VSS 0.045866f
C14167 a_31953_n19727.t308 VSS 0.042602f
C14168 a_31953_n19727.n410 VSS 0.045866f
C14169 a_31953_n19727.t183 VSS 0.039948f
C14170 a_31953_n19727.n411 VSS 0.045891f
C14171 a_31953_n19727.t318 VSS 0.042606f
C14172 a_31953_n19727.t349 VSS 0.039948f
C14173 a_31953_n19727.n412 VSS 0.045891f
C14174 a_31953_n19727.t76 VSS 0.039948f
C14175 a_31953_n19727.t150 VSS 0.039898f
C14176 a_31953_n19727.n413 VSS 0.045583f
C14177 a_31953_n19727.t285 VSS 0.042602f
C14178 a_31953_n19727.n414 VSS 0.045866f
C14179 a_31953_n19727.t147 VSS 0.039948f
C14180 a_31953_n19727.t3 VSS 0.007658f
C14181 a_31953_n19727.n415 VSS 0.022107f
C14182 a_31953_n19727.t55 VSS 0.007658f
C14183 a_31953_n19727.n416 VSS 0.016885f
C14184 a_31953_n19727.t41 VSS 0.007658f
C14185 a_31953_n19727.n417 VSS 0.022051f
C14186 a_31953_n19727.n418 VSS 0.045891f
C14187 a_31953_n19727.t230 VSS 0.042606f
C14188 a_31953_n19727.t328 VSS 0.039948f
C14189 a_31953_n19727.n419 VSS 0.045891f
C14190 a_31953_n19727.t2 VSS 0.039948f
C14191 a_31953_n19727.t263 VSS 0.039948f
C14192 a_31953_n19727.n420 VSS 0.045866f
C14193 a_31953_n19727.t323 VSS 0.042602f
C14194 a_31953_n19727.n421 VSS 0.045866f
C14195 a_31953_n19727.t22 VSS 0.039948f
C14196 a_31953_n19727.n422 VSS 0.045891f
C14197 a_31953_n19727.t304 VSS 0.042606f
C14198 a_31953_n19727.t113 VSS 0.039948f
C14199 a_31953_n19727.n423 VSS 0.045891f
C14200 a_31953_n19727.t54 VSS 0.039948f
C14201 a_31953_n19727.t334 VSS 0.039901f
C14202 a_31953_n19727.n424 VSS 0.045597f
C14203 a_31953_n19727.t108 VSS 0.042602f
C14204 a_31953_n19727.n425 VSS 0.045866f
C14205 a_31953_n19727.t0 VSS 0.039948f
C14206 a_31953_n19727.n426 VSS 0.045891f
C14207 a_31953_n19727.t360 VSS 0.042606f
C14208 a_31953_n19727.t169 VSS 0.039948f
C14209 a_31953_n19727.n427 VSS 0.045891f
C14210 a_31953_n19727.t40 VSS 0.039948f
C14211 a_31953_n19727.t101 VSS 0.039903f
C14212 a_31953_n19727.n428 VSS 0.045866f
C14213 a_31953_n19727.t165 VSS 0.042602f
C14214 a_31953_n19727.n429 VSS 0.04561f
C14215 a_31953_n19727.t56 VSS 0.039948f
C14216 a_31953_n19727.t120 VSS 0.039948f
C14217 a_31953_n19727.t307 VSS 0.039898f
C14218 a_31953_n19727.n430 VSS 0.022914f
C14219 a_31953_n19727.n431 VSS 0.045583f
C14220 a_31953_n19727.t80 VSS 0.042602f
C14221 a_31953_n19727.n432 VSS 0.045866f
C14222 a_31953_n19727.n433 VSS 0.045891f
C14223 a_31953_n19727.t282 VSS 0.042606f
C14224 a_31953_n19727.t84 VSS 0.039948f
C14225 a_31953_n19727.n434 VSS 0.045891f
C14226 a_31953_n19727.t339 VSS 0.039948f
C14227 a_31953_n19727.n435 VSS 0.045891f
C14228 a_31953_n19727.t209 VSS 0.042606f
C14229 a_31953_n19727.t303 VSS 0.039948f
C14230 a_31953_n19727.n436 VSS 0.045891f
C14231 a_31953_n19727.t338 VSS 0.039948f
C14232 a_31953_n19727.t233 VSS 0.039948f
C14233 a_31953_n19727.n437 VSS 0.045866f
C14234 a_31953_n19727.t300 VSS 0.042602f
C14235 a_31953_n19727.n438 VSS 0.045866f
C14236 a_31953_n19727.t267 VSS 0.039948f
C14237 a_31953_n19727.n439 VSS 0.045891f
C14238 a_31953_n19727.t142 VSS 0.042606f
C14239 a_31953_n19727.t247 VSS 0.039948f
C14240 a_31953_n19727.n440 VSS 0.045891f
C14241 a_31953_n19727.t287 VSS 0.039948f
C14242 a_31953_n19727.t176 VSS 0.039948f
C14243 a_31953_n19727.n441 VSS 0.045866f
C14244 a_31953_n19727.t244 VSS 0.042602f
C14245 a_31953_n19727.n442 VSS 0.045866f
C14246 a_31953_n19727.t212 VSS 0.039948f
C14247 a_31953_n19727.n443 VSS 0.024376f
C14248 a_31953_n19727.t57 VSS 0.007658f
C14249 a_31953_n19727.n444 VSS 0.021674f
C14250 a_31953_n19727.t1 VSS 0.007658f
C14251 a_31953_n19727.n445 VSS 0.016885f
C14252 a_31953_n19727.t23 VSS 0.007658f
C14253 a_31953_n19727.n446 VSS 0.021693f
C14254 a_31953_n19727.n447 VSS 0.024552f
C14255 a_31953_n19727.n448 VSS 0.045891f
C14256 a_31953_n19727.t245 VSS 0.042606f
C14257 a_31953_n19727.t344 VSS 0.039948f
C14258 a_31953_n19727.n449 VSS 0.045891f
C14259 a_31953_n19727.t83 VSS 0.039948f
C14260 a_31953_n19727.t277 VSS 0.039948f
C14261 a_31953_n19727.n450 VSS 0.045866f
C14262 a_31953_n19727.t340 VSS 0.042602f
C14263 a_31953_n19727.n451 VSS 0.045866f
C14264 a_31953_n19727.t302 VSS 0.039948f
C14265 a_31953_n19727.n452 VSS 0.045891f
C14266 a_31953_n19727.t166 VSS 0.042606f
C14267 a_31953_n19727.t272 VSS 0.039948f
C14268 a_31953_n19727.n453 VSS 0.045891f
C14269 a_31953_n19727.t301 VSS 0.039948f
C14270 a_31953_n19727.t199 VSS 0.039948f
C14271 a_31953_n19727.n454 VSS 0.045866f
C14272 a_31953_n19727.t268 VSS 0.042602f
C14273 a_31953_n19727.n455 VSS 0.045866f
C14274 a_31953_n19727.t228 VSS 0.039948f
C14275 a_31953_n19727.n456 VSS 0.046928f
C14276 a_31953_n19727.t90 VSS 0.042575f
C14277 a_31953_n19727.t196 VSS 0.039952f
C14278 a_31953_n19727.n457 VSS 0.04589f
C14279 a_31953_n19727.t227 VSS 0.039952f
C14280 a_31953_n19727.t123 VSS 0.039952f
C14281 a_31953_n19727.n458 VSS 0.046902f
C14282 a_31953_n19727.t193 VSS 0.042571f
C14283 a_31953_n19727.n459 VSS 0.045866f
C14284 a_31953_n19727.n460 VSS 0.025554f
C14285 a_31953_n19727.n461 VSS 0.025366f
C14286 a_31953_n19727.t148 VSS 0.039919f
C14287 a_31953_n19727.n462 VSS 0.108284f
C14288 a_31953_n19727.n463 VSS 0.28434f
C14289 a_31953_n19727.n464 VSS 0.210966f
C14290 a_31953_n19727.n465 VSS 0.046928f
C14291 a_31953_n19727.t246 VSS 0.042575f
C14292 a_31953_n19727.t141 VSS 0.039952f
C14293 a_31953_n19727.n466 VSS 0.04589f
C14294 a_31953_n19727.t104 VSS 0.039952f
C14295 a_31953_n19727.t358 VSS 0.039952f
C14296 a_31953_n19727.n467 VSS 0.046902f
C14297 a_31953_n19727.t290 VSS 0.042571f
C14298 a_31953_n19727.n468 VSS 0.045866f
C14299 a_31953_n19727.n469 VSS 0.025554f
C14300 a_31953_n19727.n470 VSS 0.025366f
C14301 a_31953_n19727.t330 VSS 0.039919f
C14302 a_31953_n19727.n471 VSS 0.045891f
C14303 a_31953_n19727.t317 VSS 0.042606f
C14304 a_31953_n19727.t220 VSS 0.039948f
C14305 a_31953_n19727.n472 VSS 0.045891f
C14306 a_31953_n19727.t182 VSS 0.039948f
C14307 a_31953_n19727.t140 VSS 0.039948f
C14308 a_31953_n19727.n473 VSS 0.045866f
C14309 a_31953_n19727.t361 VSS 0.042602f
C14310 a_31953_n19727.n474 VSS 0.045866f
C14311 a_31953_n19727.t115 VSS 0.039948f
C14312 a_31953_n19727.n475 VSS 0.045891f
C14313 a_31953_n19727.t98 VSS 0.042606f
C14314 a_31953_n19727.t292 VSS 0.039948f
C14315 a_31953_n19727.n476 VSS 0.045891f
C14316 a_31953_n19727.t260 VSS 0.039948f
C14317 a_31953_n19727.t217 VSS 0.039948f
C14318 a_31953_n19727.n477 VSS 0.045866f
C14319 a_31953_n19727.t143 VSS 0.042602f
C14320 a_31953_n19727.n478 VSS 0.045866f
C14321 a_31953_n19727.t190 VSS 0.039948f
C14322 a_31953_n19727.t37 VSS 0.007658f
C14323 a_31953_n19727.n479 VSS 0.022107f
C14324 a_31953_n19727.t35 VSS 0.007658f
C14325 a_31953_n19727.n480 VSS 0.016885f
C14326 a_31953_n19727.t51 VSS 0.007658f
C14327 a_31953_n19727.n481 VSS 0.021693f
C14328 a_31953_n19727.n482 VSS 0.024552f
C14329 a_31953_n19727.n483 VSS 0.045891f
C14330 a_31953_n19727.t86 VSS 0.042606f
C14331 a_31953_n19727.t284 VSS 0.039948f
C14332 a_31953_n19727.n484 VSS 0.045891f
C14333 a_31953_n19727.t36 VSS 0.039948f
C14334 a_31953_n19727.t204 VSS 0.039948f
C14335 a_31953_n19727.n485 VSS 0.045866f
C14336 a_31953_n19727.t135 VSS 0.042602f
C14337 a_31953_n19727.n486 VSS 0.045866f
C14338 a_31953_n19727.t50 VSS 0.039948f
C14339 a_31953_n19727.n487 VSS 0.045891f
C14340 a_31953_n19727.t158 VSS 0.042606f
C14341 a_31953_n19727.t355 VSS 0.039948f
C14342 a_31953_n19727.n488 VSS 0.045891f
C14343 a_31953_n19727.t12 VSS 0.039948f
C14344 a_31953_n19727.t280 VSS 0.039901f
C14345 a_31953_n19727.n489 VSS 0.045597f
C14346 a_31953_n19727.t214 VSS 0.042602f
C14347 a_31953_n19727.n490 VSS 0.045866f
C14348 a_31953_n19727.t34 VSS 0.039948f
C14349 a_31953_n19727.n491 VSS 0.045891f
C14350 a_31953_n19727.t222 VSS 0.042606f
C14351 a_31953_n19727.t122 VSS 0.039948f
C14352 a_31953_n19727.n492 VSS 0.045891f
C14353 a_31953_n19727.t70 VSS 0.039948f
C14354 a_31953_n19727.t337 VSS 0.039903f
C14355 a_31953_n19727.n493 VSS 0.045866f
C14356 a_31953_n19727.t274 VSS 0.042602f
C14357 a_31953_n19727.n494 VSS 0.04561f
C14358 a_31953_n19727.t18 VSS 0.039948f
C14359 a_31953_n19727.t289 VSS 0.039948f
C14360 a_31953_n19727.t254 VSS 0.039898f
C14361 a_31953_n19727.n495 VSS 0.022914f
C14362 a_31953_n19727.n496 VSS 0.045583f
C14363 a_31953_n19727.t184 VSS 0.042602f
C14364 a_31953_n19727.n497 VSS 0.045866f
C14365 a_31953_n19727.n498 VSS 0.045891f
C14366 a_31953_n19727.t137 VSS 0.042606f
C14367 a_31953_n19727.t325 VSS 0.039948f
C14368 a_31953_n19727.n499 VSS 0.045891f
C14369 a_31953_n19727.t223 VSS 0.039948f
C14370 a_31953_n19727.n500 VSS 0.045891f
C14371 a_31953_n19727.t354 VSS 0.042606f
C14372 a_31953_n19727.t257 VSS 0.039948f
C14373 a_31953_n19727.n501 VSS 0.045891f
C14374 a_31953_n19727.t218 VSS 0.039948f
C14375 a_31953_n19727.t178 VSS 0.039948f
C14376 a_31953_n19727.n502 VSS 0.045866f
C14377 a_31953_n19727.t110 VSS 0.042602f
C14378 a_31953_n19727.n503 VSS 0.045866f
C14379 a_31953_n19727.t144 VSS 0.039948f
C14380 a_31953_n19727.n504 VSS 0.045891f
C14381 a_31953_n19727.t296 VSS 0.042606f
C14382 a_31953_n19727.t198 VSS 0.039948f
C14383 a_31953_n19727.n505 VSS 0.045891f
C14384 a_31953_n19727.t152 VSS 0.039948f
C14385 a_31953_n19727.t119 VSS 0.039948f
C14386 a_31953_n19727.n506 VSS 0.045866f
C14387 a_31953_n19727.t346 VSS 0.042602f
C14388 a_31953_n19727.n507 VSS 0.045866f
C14389 a_31953_n19727.t88 VSS 0.039948f
C14390 a_31953_n19727.n508 VSS 0.024376f
C14391 a_31953_n19727.n509 VSS 0.022051f
C14392 a_31953_n19727.t71 VSS 0.007658f
C14393 a_33249_35053.n0 VSS 1.83524f
C14394 a_33249_35053.n1 VSS 1.4665f
C14395 a_33249_35053.n2 VSS 1.57152f
C14396 a_33249_35053.n3 VSS 1.92894f
C14397 a_33249_35053.n4 VSS 1.68723f
C14398 a_33249_35053.n5 VSS 1.08952f
C14399 a_33249_35053.n6 VSS 1.92894f
C14400 a_33249_35053.n7 VSS 1.68723f
C14401 a_33249_35053.n8 VSS 1.08952f
C14402 a_33249_35053.n9 VSS 2.09988f
C14403 a_33249_35053.n10 VSS 4.85677f
C14404 a_33249_35053.t109 VSS 0.07106f
C14405 a_33249_35053.t122 VSS 0.07106f
C14406 a_33249_35053.n11 VSS 0.177102f
C14407 a_33249_35053.t107 VSS 0.07106f
C14408 a_33249_35053.t119 VSS 0.07106f
C14409 a_33249_35053.n12 VSS 0.190759f
C14410 a_33249_35053.n13 VSS 0.637527f
C14411 a_33249_35053.n14 VSS 7.50995f
C14412 a_33249_35053.n15 VSS 3.02979f
C14413 a_33249_35053.t5 VSS 0.196574f
C14414 a_33249_35053.t4 VSS 0.20931f
C14415 a_33249_35053.n16 VSS 0.794625f
C14416 a_33249_35053.t28 VSS 0.074613f
C14417 a_33249_35053.t57 VSS 0.074613f
C14418 a_33249_35053.n17 VSS 0.189335f
C14419 a_33249_35053.t26 VSS 0.074613f
C14420 a_33249_35053.t55 VSS 0.074613f
C14421 a_33249_35053.n18 VSS 0.204335f
C14422 a_33249_35053.n19 VSS 0.518601f
C14423 a_33249_35053.n20 VSS 0.432177f
C14424 a_33249_35053.t36 VSS 0.196574f
C14425 a_33249_35053.t34 VSS 0.20931f
C14426 a_33249_35053.n21 VSS 0.79384f
C14427 a_33249_35053.t76 VSS 0.074613f
C14428 a_33249_35053.t22 VSS 0.074613f
C14429 a_33249_35053.n22 VSS 0.189335f
C14430 a_33249_35053.t75 VSS 0.074613f
C14431 a_33249_35053.t20 VSS 0.074613f
C14432 a_33249_35053.n23 VSS 0.204335f
C14433 a_33249_35053.n24 VSS 0.518601f
C14434 a_33249_35053.n25 VSS 0.547885f
C14435 a_33249_35053.t21 VSS 0.196574f
C14436 a_33249_35053.t19 VSS 0.20931f
C14437 a_33249_35053.n26 VSS 0.659973f
C14438 a_33249_35053.n27 VSS 0.604093f
C14439 a_33249_35053.t56 VSS 0.196574f
C14440 a_33249_35053.t53 VSS 0.20931f
C14441 a_33249_35053.n28 VSS 0.662721f
C14442 a_33249_35053.n29 VSS 0.510661f
C14443 a_33249_35053.n30 VSS 4.45672f
C14444 a_33249_35053.t78 VSS 0.074613f
C14445 a_33249_35053.t29 VSS 0.074613f
C14446 a_33249_35053.n31 VSS 0.717178f
C14447 a_33249_35053.t51 VSS 0.335476f
C14448 a_33249_35053.n32 VSS 1.92412f
C14449 a_33249_35053.n33 VSS 1.99746f
C14450 a_33249_35053.t88 VSS 0.074613f
C14451 a_33249_35053.t46 VSS 0.074613f
C14452 a_33249_35053.n34 VSS 0.344546f
C14453 a_33249_35053.n35 VSS 1.69025f
C14454 a_33249_35053.t61 VSS 0.335476f
C14455 a_33249_35053.n36 VSS 1.57565f
C14456 a_33249_35053.t2 VSS 0.196574f
C14457 a_33249_35053.t85 VSS 0.20931f
C14458 a_33249_35053.n37 VSS 0.794625f
C14459 a_33249_35053.t24 VSS 0.074613f
C14460 a_33249_35053.t50 VSS 0.074613f
C14461 a_33249_35053.n38 VSS 0.189335f
C14462 a_33249_35053.t15 VSS 0.074613f
C14463 a_33249_35053.t40 VSS 0.074613f
C14464 a_33249_35053.n39 VSS 0.204335f
C14465 a_33249_35053.n40 VSS 0.518601f
C14466 a_33249_35053.n41 VSS 0.432177f
C14467 a_33249_35053.t32 VSS 0.196574f
C14468 a_33249_35053.t30 VSS 0.20931f
C14469 a_33249_35053.n42 VSS 0.79384f
C14470 a_33249_35053.t71 VSS 0.074613f
C14471 a_33249_35053.t14 VSS 0.074613f
C14472 a_33249_35053.n43 VSS 0.189335f
C14473 a_33249_35053.t67 VSS 0.074613f
C14474 a_33249_35053.t9 VSS 0.074613f
C14475 a_33249_35053.n44 VSS 0.204335f
C14476 a_33249_35053.n45 VSS 0.518601f
C14477 a_33249_35053.n46 VSS 0.547885f
C14478 a_33249_35053.t13 VSS 0.196574f
C14479 a_33249_35053.t8 VSS 0.20931f
C14480 a_33249_35053.n47 VSS 0.659973f
C14481 a_33249_35053.n48 VSS 0.604093f
C14482 a_33249_35053.t48 VSS 0.196574f
C14483 a_33249_35053.t39 VSS 0.20931f
C14484 a_33249_35053.n49 VSS 0.662721f
C14485 a_33249_35053.n50 VSS 0.510661f
C14486 a_33249_35053.n51 VSS 0.205287f
C14487 a_33249_35053.t77 VSS 0.074613f
C14488 a_33249_35053.t23 VSS 0.074613f
C14489 a_33249_35053.n52 VSS 0.189335f
C14490 a_33249_35053.t70 VSS 0.074613f
C14491 a_33249_35053.t12 VSS 0.074613f
C14492 a_33249_35053.n53 VSS 0.204335f
C14493 a_33249_35053.n54 VSS 0.518601f
C14494 a_33249_35053.n55 VSS 0.288394f
C14495 a_33249_35053.t52 VSS 0.196574f
C14496 a_33249_35053.t43 VSS 0.20931f
C14497 a_33249_35053.n56 VSS 0.669825f
C14498 a_33249_35053.n57 VSS 0.61504f
C14499 a_33249_35053.t38 VSS 0.196574f
C14500 a_33249_35053.t33 VSS 0.20931f
C14501 a_33249_35053.n58 VSS 0.669825f
C14502 a_33249_35053.n59 VSS 0.615019f
C14503 a_33249_35053.t81 VSS 0.074613f
C14504 a_33249_35053.t11 VSS 0.074613f
C14505 a_33249_35053.n60 VSS 0.189335f
C14506 a_33249_35053.t72 VSS 0.074613f
C14507 a_33249_35053.t6 VSS 0.074613f
C14508 a_33249_35053.n61 VSS 0.204335f
C14509 a_33249_35053.n62 VSS 0.518601f
C14510 a_33249_35053.n63 VSS 0.405037f
C14511 a_33249_35053.t41 VSS 0.196574f
C14512 a_33249_35053.t37 VSS 0.20931f
C14513 a_33249_35053.n64 VSS 0.659973f
C14514 a_33249_35053.n65 VSS 0.604093f
C14515 a_33249_35053.t73 VSS 0.196574f
C14516 a_33249_35053.t69 VSS 0.20931f
C14517 a_33249_35053.n66 VSS 0.662721f
C14518 a_33249_35053.n67 VSS 0.510661f
C14519 a_33249_35053.n68 VSS 0.205287f
C14520 a_33249_35053.n69 VSS 4.86153f
C14521 a_33249_35053.n70 VSS 3.25477f
C14522 a_33249_35053.t66 VSS 0.074613f
C14523 a_33249_35053.t7 VSS 0.074613f
C14524 a_33249_35053.n71 VSS 0.347301f
C14525 a_33249_35053.t62 VSS 0.337446f
C14526 a_33249_35053.t63 VSS 0.074613f
C14527 a_33249_35053.t1 VSS 0.074613f
C14528 a_33249_35053.n72 VSS 0.347301f
C14529 a_33249_35053.t35 VSS 0.611504f
C14530 a_33249_35053.n73 VSS 1.41648f
C14531 a_33249_35053.n74 VSS 2.82773f
C14532 a_33249_35053.t64 VSS 0.335476f
C14533 a_33249_35053.n75 VSS 1.11142f
C14534 a_33249_35053.t3 VSS 0.074613f
C14535 a_33249_35053.t54 VSS 0.074613f
C14536 a_33249_35053.n76 VSS 0.344546f
C14537 a_33249_35053.n77 VSS 1.69025f
C14538 a_33249_35053.t84 VSS 0.074613f
C14539 a_33249_35053.t31 VSS 0.074613f
C14540 a_33249_35053.n78 VSS 0.717178f
C14541 a_33249_35053.t58 VSS 0.335476f
C14542 a_33249_35053.n79 VSS 1.92412f
C14543 a_33249_35053.n80 VSS 1.41725f
C14544 a_33249_35053.n81 VSS 2.74097f
C14545 a_33249_35053.n82 VSS 3.27733f
C14546 a_33249_35053.n83 VSS 0.205287f
C14547 a_33249_35053.t83 VSS 0.074613f
C14548 a_33249_35053.t27 VSS 0.074613f
C14549 a_33249_35053.n84 VSS 0.189335f
C14550 a_33249_35053.t82 VSS 0.074613f
C14551 a_33249_35053.t25 VSS 0.074613f
C14552 a_33249_35053.n85 VSS 0.204335f
C14553 a_33249_35053.n86 VSS 0.518601f
C14554 a_33249_35053.n87 VSS 0.288394f
C14555 a_33249_35053.t60 VSS 0.196574f
C14556 a_33249_35053.t59 VSS 0.20931f
C14557 a_33249_35053.n88 VSS 0.669825f
C14558 a_33249_35053.n89 VSS 0.61504f
C14559 a_33249_35053.t44 VSS 0.196574f
C14560 a_33249_35053.t42 VSS 0.20931f
C14561 a_33249_35053.n90 VSS 0.669825f
C14562 a_33249_35053.n91 VSS 0.615019f
C14563 a_33249_35053.t87 VSS 0.074613f
C14564 a_33249_35053.t17 VSS 0.074613f
C14565 a_33249_35053.n92 VSS 0.189335f
C14566 a_33249_35053.t86 VSS 0.074613f
C14567 a_33249_35053.t16 VSS 0.074613f
C14568 a_33249_35053.n93 VSS 0.204335f
C14569 a_33249_35053.n94 VSS 0.518601f
C14570 a_33249_35053.n95 VSS 0.405037f
C14571 a_33249_35053.t49 VSS 0.196574f
C14572 a_33249_35053.t47 VSS 0.20931f
C14573 a_33249_35053.n96 VSS 0.659973f
C14574 a_33249_35053.n97 VSS 0.604093f
C14575 a_33249_35053.t80 VSS 0.196574f
C14576 a_33249_35053.t79 VSS 0.20931f
C14577 a_33249_35053.n98 VSS 0.662721f
C14578 a_33249_35053.n99 VSS 0.510661f
C14579 a_33249_35053.n100 VSS 0.205287f
C14580 a_33249_35053.n101 VSS 3.27733f
C14581 a_33249_35053.t74 VSS 0.074613f
C14582 a_33249_35053.t18 VSS 0.074613f
C14583 a_33249_35053.n102 VSS 0.347301f
C14584 a_33249_35053.t65 VSS 0.337446f
C14585 a_33249_35053.t68 VSS 0.074613f
C14586 a_33249_35053.t10 VSS 0.074613f
C14587 a_33249_35053.n103 VSS 0.347301f
C14588 a_33249_35053.t45 VSS 0.611504f
C14589 a_33249_35053.n104 VSS 1.41648f
C14590 a_33249_35053.n105 VSS 4.42321f
C14591 a_33249_35053.n106 VSS 12.737201f
C14592 a_33249_35053.t92 VSS 0.528339f
C14593 a_33249_35053.t89 VSS 0.07106f
C14594 a_33249_35053.t95 VSS 0.07106f
C14595 a_33249_35053.n107 VSS 0.278463f
C14596 a_33249_35053.n108 VSS 2.09739f
C14597 a_33249_35053.n109 VSS 9.46617f
C14598 a_33249_35053.t91 VSS 0.22239f
C14599 a_33249_35053.t105 VSS 0.182969f
C14600 a_33249_35053.n110 VSS 0.795201f
C14601 a_33249_35053.t100 VSS 0.07106f
C14602 a_33249_35053.t97 VSS 0.07106f
C14603 a_33249_35053.n111 VSS 0.20821f
C14604 a_33249_35053.t98 VSS 0.07106f
C14605 a_33249_35053.t93 VSS 0.07106f
C14606 a_33249_35053.n112 VSS 0.163168f
C14607 a_33249_35053.n113 VSS 0.528707f
C14608 a_33249_35053.n114 VSS 0.979027f
C14609 a_33249_35053.t101 VSS 0.07106f
C14610 a_33249_35053.t104 VSS 0.07106f
C14611 a_33249_35053.n115 VSS 0.20821f
C14612 a_33249_35053.t90 VSS 0.07106f
C14613 a_33249_35053.t94 VSS 0.07106f
C14614 a_33249_35053.n116 VSS 0.163168f
C14615 a_33249_35053.n117 VSS 0.528707f
C14616 a_33249_35053.n118 VSS 0.802261f
C14617 a_33249_35053.t0 VSS 0.22239f
C14618 a_33249_35053.t96 VSS 0.182969f
C14619 a_33249_35053.n119 VSS 0.643953f
C14620 a_33249_35053.n120 VSS 0.300334f
C14621 a_33249_35053.n121 VSS 2.86645f
C14622 a_33249_35053.t103 VSS 0.287637f
C14623 a_33249_35053.t99 VSS 0.07106f
C14624 a_33249_35053.t102 VSS 0.07106f
C14625 a_33249_35053.n122 VSS 0.602285f
C14626 a_33249_35053.n123 VSS 3.53981f
C14627 a_33249_35053.n124 VSS 5.24967f
C14628 a_33249_35053.t128 VSS 0.07106f
C14629 a_33249_35053.t141 VSS 0.07106f
C14630 a_33249_35053.n125 VSS 0.638798f
C14631 a_33249_35053.t130 VSS 0.326634f
C14632 a_33249_35053.n126 VSS 1.84327f
C14633 a_33249_35053.n127 VSS 1.20691f
C14634 a_33249_35053.t114 VSS 0.07106f
C14635 a_33249_35053.t129 VSS 0.07106f
C14636 a_33249_35053.n128 VSS 0.322136f
C14637 a_33249_35053.n129 VSS 1.48873f
C14638 a_33249_35053.t117 VSS 0.326634f
C14639 a_33249_35053.n130 VSS 1.06366f
C14640 a_33249_35053.n131 VSS 4.2966f
C14641 a_33249_35053.t113 VSS 0.07106f
C14642 a_33249_35053.t111 VSS 0.07106f
C14643 a_33249_35053.n132 VSS 0.324656f
C14644 a_33249_35053.t126 VSS 0.328556f
C14645 a_33249_35053.n133 VSS 5.31934f
C14646 a_33249_35053.n134 VSS 0.4889f
C14647 a_33249_35053.t120 VSS 0.195319f
C14648 a_33249_35053.t115 VSS 0.207237f
C14649 a_33249_35053.n135 VSS 0.639651f
C14650 a_33249_35053.n136 VSS 0.514924f
C14651 a_33249_35053.t124 VSS 0.195319f
C14652 a_33249_35053.t123 VSS 0.207237f
C14653 a_33249_35053.n137 VSS 0.636903f
C14654 a_33249_35053.n138 VSS 0.605515f
C14655 a_33249_35053.t138 VSS 0.07106f
C14656 a_33249_35053.t110 VSS 0.07106f
C14657 a_33249_35053.n139 VSS 0.177102f
C14658 a_33249_35053.t135 VSS 0.07106f
C14659 a_33249_35053.t108 VSS 0.07106f
C14660 a_33249_35053.n140 VSS 0.190759f
C14661 a_33249_35053.n141 VSS 0.532224f
C14662 a_33249_35053.n142 VSS 0.804026f
C14663 a_33249_35053.t121 VSS 0.07106f
C14664 a_33249_35053.t133 VSS 0.07106f
C14665 a_33249_35053.n143 VSS 0.177102f
C14666 a_33249_35053.t116 VSS 0.07106f
C14667 a_33249_35053.t131 VSS 0.07106f
C14668 a_33249_35053.n144 VSS 0.190759f
C14669 a_33249_35053.n145 VSS 0.532224f
C14670 a_33249_35053.n146 VSS 0.687283f
C14671 a_33249_35053.t118 VSS 0.07106f
C14672 a_33249_35053.t136 VSS 0.07106f
C14673 a_33249_35053.n147 VSS 0.177102f
C14674 a_33249_35053.t112 VSS 0.07106f
C14675 a_33249_35053.t132 VSS 0.07106f
C14676 a_33249_35053.n148 VSS 0.190759f
C14677 a_33249_35053.n149 VSS 0.775507f
C14678 a_33249_35053.t106 VSS 0.195319f
C14679 a_33249_35053.t139 VSS 0.207237f
C14680 a_33249_35053.n150 VSS 0.636903f
C14681 a_33249_35053.n151 VSS 0.889874f
C14682 a_33249_35053.t137 VSS 0.195319f
C14683 a_33249_35053.t134 VSS 0.207237f
C14684 a_33249_35053.n152 VSS 0.639651f
C14685 a_33249_35053.n153 VSS 0.514924f
C14686 a_33249_35053.n154 VSS 0.202572f
C14687 a_33249_35053.n155 VSS 4.69303f
C14688 a_33249_35053.n156 VSS 1.94054f
C14689 a_33249_35053.t127 VSS 0.07106f
C14690 a_33249_35053.t125 VSS 0.07106f
C14691 a_33249_35053.n157 VSS 0.324656f
C14692 a_33249_35053.t140 VSS 0.567904f
C14693 a_35502_25545.n0 VSS 0.054238f
C14694 a_35502_25545.n1 VSS 0.201858f
C14695 a_35502_25545.n2 VSS 0.169544f
C14696 a_35502_25545.n3 VSS 0.02883f
C14697 a_35502_25545.n4 VSS 0.028228f
C14698 a_35502_25545.n5 VSS 0.163138f
C14699 a_35502_25545.n6 VSS 0.195374f
C14700 a_35502_25545.n7 VSS 0.057098f
C14701 a_35502_25545.n8 VSS 0.163138f
C14702 a_35502_25545.n9 VSS 0.195374f
C14703 a_35502_25545.n10 VSS 0.057098f
C14704 a_35502_25545.n11 VSS 0.068083f
C14705 a_35502_25545.n12 VSS 0.031561f
C14706 a_35502_25545.n13 VSS 0.068083f
C14707 a_35502_25545.n14 VSS 0.031561f
C14708 a_35502_25545.n15 VSS 0.129052f
C14709 a_35502_25545.n16 VSS 0.074307f
C14710 a_35502_25545.n17 VSS 0.131171f
C14711 a_35502_25545.n18 VSS 0.129052f
C14712 a_35502_25545.n19 VSS 0.072194f
C14713 a_35502_25545.n20 VSS 0.169544f
C14714 a_35502_25545.n21 VSS 0.024914f
C14715 a_35502_25545.n22 VSS 0.072194f
C14716 a_35502_25545.n23 VSS 0.169544f
C14717 a_35502_25545.n24 VSS 0.024914f
C14718 a_35502_25545.n25 VSS 0.025009f
C14719 a_35502_25545.n26 VSS 0.072519f
C14720 a_35502_25545.n27 VSS 0.074307f
C14721 a_35502_25545.n28 VSS 0.16987f
C14722 a_35502_25545.n29 VSS 0.025009f
C14723 a_35502_25545.n30 VSS 0.074307f
C14724 a_35502_25545.n31 VSS 0.16987f
C14725 a_35502_25545.n32 VSS 0.025009f
C14726 a_35502_25545.n33 VSS 0.10095f
C14727 a_35502_25545.n34 VSS 0.1331f
C14728 a_35502_25545.n35 VSS 0.043969f
C14729 a_35502_25545.n36 VSS 0.04169f
C14730 a_35502_25545.n37 VSS 0.124713f
C14731 a_35502_25545.n38 VSS 0.024358f
C14732 a_35502_25545.n39 VSS 0.043969f
C14733 a_35502_25545.n40 VSS 0.1331f
C14734 a_35502_25545.n41 VSS 0.04169f
C14735 a_35502_25545.n42 VSS 0.061624f
C14736 a_35502_25545.n43 VSS 0.130169f
C14737 a_35502_25545.n44 VSS 0.04169f
C14738 a_35502_25545.n45 VSS 0.044881f
C14739 a_35502_25545.n46 VSS 0.392837f
C14740 a_35502_25545.n47 VSS 0.02135f
C14741 a_35502_25545.n48 VSS 0.044881f
C14742 a_35502_25545.n49 VSS 0.061624f
C14743 a_35502_25545.n50 VSS 0.130169f
C14744 a_35502_25545.n51 VSS 0.04169f
C14745 a_35502_25545.n52 VSS 0.025532f
C14746 a_35502_25545.n53 VSS 0.074307f
C14747 a_35502_25545.n54 VSS 0.061624f
C14748 a_35502_25545.n55 VSS 0.171655f
C14749 a_35502_25545.n56 VSS 0.025532f
C14750 a_35502_25545.n57 VSS 0.171655f
C14751 a_35502_25545.n58 VSS 0.025532f
C14752 a_35502_25545.n59 VSS 0.025532f
C14753 a_35502_25545.n60 VSS 0.072194f
C14754 a_35502_25545.n61 VSS 0.135361f
C14755 a_35502_25545.n62 VSS 0.095594f
C14756 a_35502_25545.n63 VSS 0.04215f
C14757 a_35502_25545.n64 VSS 0.072194f
C14758 a_35502_25545.n65 VSS 0.135361f
C14759 a_35502_25545.n66 VSS 0.095594f
C14760 a_35502_25545.n67 VSS 0.04215f
C14761 a_35502_25545.n68 VSS 0.163138f
C14762 a_35502_25545.n69 VSS 0.08974f
C14763 a_35502_25545.n70 VSS 0.072194f
C14764 a_35502_25545.n71 VSS 0.16987f
C14765 a_35502_25545.n72 VSS 0.024914f
C14766 a_35502_25545.n73 VSS 0.025009f
C14767 a_35502_25545.n74 VSS 0.072194f
C14768 a_35502_25545.n75 VSS 0.16987f
C14769 a_35502_25545.n76 VSS 0.024914f
C14770 a_35502_25545.n77 VSS 0.025009f
C14771 a_35502_25545.n78 VSS 0.171655f
C14772 a_35502_25545.n79 VSS 0.025532f
C14773 a_35502_25545.n80 VSS 0.025532f
C14774 a_35502_25545.n81 VSS 0.06894f
C14775 a_35502_25545.n82 VSS 0.171654f
C14776 a_35502_25545.n83 VSS 0.086209f
C14777 a_35502_25545.n84 VSS 0.08875f
C14778 a_35502_25545.n85 VSS 0.041717f
C14779 a_35502_25545.n86 VSS 0.171654f
C14780 a_35502_25545.n87 VSS 0.024914f
C14781 a_35502_25545.n88 VSS 0.025532f
C14782 a_35502_25545.n89 VSS 0.06894f
C14783 a_35502_25545.n90 VSS 0.171654f
C14784 a_35502_25545.n91 VSS 0.028228f
C14785 a_35502_25545.n92 VSS 0.02883f
C14786 a_35502_25545.n93 VSS 0.162625f
C14787 a_35502_25545.n94 VSS 0.089858f
C14788 a_35502_25545.n95 VSS 0.084816f
C14789 a_35502_25545.n96 VSS 0.138411f
C14790 a_35502_25545.n97 VSS 0.068636f
C14791 a_35502_25545.n98 VSS 0.019526f
C14792 a_35502_25545.n99 VSS 0.018822f
C14793 a_35502_25545.n100 VSS 0.068636f
C14794 a_35502_25545.n101 VSS 0.068636f
C14795 a_35502_25545.n102 VSS 0.02135f
C14796 a_35502_25545.n103 VSS 0.02436f
C14797 a_35502_25545.n104 VSS 0.088546f
C14798 a_35502_25545.n105 VSS 0.028259f
C14799 a_35502_25545.n106 VSS 0.027763f
C14800 a_35502_25545.n107 VSS 0.027763f
C14801 a_35502_25545.n108 VSS 0.068284f
C14802 a_35502_25545.n109 VSS 0.079891f
C14803 a_35502_25545.n110 VSS 0.132962f
C14804 a_35502_25545.n111 VSS 0.019526f
C14805 a_35502_25545.n112 VSS 0.068284f
C14806 a_35502_25545.n113 VSS 0.132284f
C14807 a_35502_25545.n114 VSS 0.020097f
C14808 a_35502_25545.n115 VSS 0.077331f
C14809 a_35502_25545.n116 VSS 0.01148f
C14810 a_35502_25545.n117 VSS 0.019614f
C14811 a_35502_25545.n118 VSS 0.068196f
C14812 a_35502_25545.n119 VSS 0.068196f
C14813 a_35502_25545.n120 VSS 0.064876f
C14814 a_35502_25545.n121 VSS 0.064876f
C14815 a_35502_25545.n122 VSS 0.098651f
C14816 a_35502_25545.n123 VSS 0.042029f
C14817 a_35502_25545.n124 VSS 0.072194f
C14818 a_35502_25545.n125 VSS 0.13155f
C14819 a_35502_25545.n126 VSS 0.042363f
C14820 a_35502_25545.n127 VSS 0.072194f
C14821 a_35502_25545.n128 VSS 0.13155f
C14822 a_35502_25545.n129 VSS 0.042363f
C14823 a_35502_25545.n130 VSS 0.01148f
C14824 a_35502_25545.n131 VSS 0.072519f
C14825 a_35502_25545.n132 VSS 0.098326f
C14826 a_35502_25545.n133 VSS 0.098326f
C14827 a_35502_25545.n134 VSS 0.285733f
C14828 a_35502_25545.n135 VSS 0.157254f
C14829 a_35502_25545.n136 VSS 0.083613f
C14830 a_35502_25545.n137 VSS 0.058769f
C14831 a_35502_25545.n138 VSS 0.281135f
C14832 a_35502_25545.n139 VSS 0.019866f
C14833 a_35502_25545.n140 VSS 0.058867f
C14834 a_35502_25545.n141 VSS 0.00797f
C14835 a_35502_25545.n142 VSS 0.086736f
C14836 a_35502_25545.t21 VSS 0.092644f
C14837 a_35502_25545.n143 VSS 1.05169f
C14838 a_35502_25545.n144 VSS 0.460139f
C14839 a_35502_25545.n145 VSS 0.095824f
C14840 a_35502_25545.n146 VSS 0.016667f
C14841 a_35502_25545.n147 VSS 0.01148f
C14842 a_35502_25545.n148 VSS 0.024921f
C14843 a_35502_25545.n149 VSS 0.020646f
C14844 a_35502_25545.t87 VSS 0.16147f
C14845 a_35502_25545.n150 VSS 0.392837f
C14846 a_35502_25545.n151 VSS 0.02436f
C14847 a_35502_25545.t79 VSS 0.16147f
C14848 a_35502_25545.n152 VSS 0.134579f
C14849 a_35502_25545.t96 VSS 0.16147f
C14850 a_35502_25545.t73 VSS 0.16147f
C14851 a_35502_25545.n153 VSS 0.02135f
C14852 a_35502_25545.n154 VSS 0.02135f
C14853 a_35502_25545.t76 VSS 0.16147f
C14854 a_35502_25545.n155 VSS 0.04212f
C14855 a_35502_25545.n156 VSS 0.024349f
C14856 a_35502_25545.n157 VSS 0.068292f
C14857 a_35502_25545.t82 VSS 0.16147f
C14858 a_35502_25545.n158 VSS 0.027662f
C14859 a_35502_25545.t53 VSS 0.16147f
C14860 a_35502_25545.t68 VSS 0.16147f
C14861 a_35502_25545.t40 VSS 0.16147f
C14862 a_35502_25545.n159 VSS 0.128168f
C14863 a_35502_25545.t95 VSS 0.16147f
C14864 a_35502_25545.t75 VSS 0.16147f
C14865 a_35502_25545.t49 VSS 0.16147f
C14866 a_35502_25545.n160 VSS 0.02135f
C14867 a_35502_25545.n161 VSS 0.04212f
C14868 a_35502_25545.t41 VSS 0.16147f
C14869 a_35502_25545.n162 VSS 0.02436f
C14870 a_35502_25545.t52 VSS 0.16147f
C14871 a_35502_25545.n163 VSS 0.134579f
C14872 a_35502_25545.n164 VSS 0.024349f
C14873 a_35502_25545.n165 VSS 0.068292f
C14874 a_35502_25545.t54 VSS 0.16147f
C14875 a_35502_25545.n166 VSS 0.027662f
C14876 a_35502_25545.t28 VSS 0.16147f
C14877 a_35502_25545.t103 VSS 0.16147f
C14878 a_35502_25545.t78 VSS 0.16147f
C14879 a_35502_25545.t44 VSS 0.16147f
C14880 a_35502_25545.n167 VSS 0.090742f
C14881 a_35502_25545.n168 VSS 0.02767f
C14882 a_35502_25545.n169 VSS 0.02436f
C14883 a_35502_25545.t56 VSS 0.16147f
C14884 a_35502_25545.n170 VSS 0.130136f
C14885 a_35502_25545.n171 VSS 0.028259f
C14886 a_35502_25545.t51 VSS 0.16147f
C14887 a_35502_25545.t80 VSS 0.16147f
C14888 a_35502_25545.n172 VSS 0.028259f
C14889 a_35502_25545.t45 VSS 0.16147f
C14890 a_35502_25545.n173 VSS 0.023957f
C14891 a_35502_25545.n174 VSS 0.02436f
C14892 a_35502_25545.t83 VSS 0.16147f
C14893 a_35502_25545.n175 VSS 0.130136f
C14894 a_35502_25545.t81 VSS 0.16147f
C14895 a_35502_25545.n176 VSS 0.02135f
C14896 a_35502_25545.t77 VSS 0.16147f
C14897 a_35502_25545.n177 VSS 0.080622f
C14898 a_35502_25545.t102 VSS 0.16147f
C14899 a_35502_25545.n178 VSS 0.080614f
C14900 a_35502_25545.n179 VSS 0.02135f
C14901 a_35502_25545.n180 VSS 0.02135f
C14902 a_35502_25545.n181 VSS 0.02135f
C14903 a_35502_25545.n182 VSS 0.042119f
C14904 a_35502_25545.n183 VSS 0.024348f
C14905 a_35502_25545.n184 VSS 0.064403f
C14906 a_35502_25545.t86 VSS 0.16147f
C14907 a_35502_25545.t57 VSS 0.16147f
C14908 a_35502_25545.t72 VSS 0.16147f
C14909 a_35502_25545.n185 VSS 0.01148f
C14910 a_35502_25545.n186 VSS 0.092213f
C14911 a_35502_25545.n187 VSS 0.032845f
C14912 a_35502_25545.n188 VSS 0.040756f
C14913 a_35502_25545.n189 VSS 0.01148f
C14914 a_35502_25545.n190 VSS 0.023957f
C14915 a_35502_25545.n191 VSS 0.028259f
C14916 a_35502_25545.t100 VSS 0.16147f
C14917 a_35502_25545.n192 VSS 0.131013f
C14918 a_35502_25545.n193 VSS 0.03317f
C14919 a_35502_25545.n194 VSS 0.131013f
C14920 a_35502_25545.n195 VSS 0.028259f
C14921 a_35502_25545.n196 VSS 0.02135f
C14922 a_35502_25545.n197 VSS 0.02135f
C14923 a_35502_25545.n198 VSS 0.061624f
C14924 a_35502_25545.n199 VSS 0.02135f
C14925 a_35502_25545.t47 VSS 0.16147f
C14926 a_35502_25545.n200 VSS 0.042119f
C14927 a_35502_25545.n201 VSS 0.024348f
C14928 a_35502_25545.n202 VSS 0.064403f
C14929 a_35502_25545.t59 VSS 0.16147f
C14930 a_35502_25545.t29 VSS 0.16147f
C14931 a_35502_25545.n203 VSS 0.040756f
C14932 a_35502_25545.n204 VSS 0.01148f
C14933 a_35502_25545.n205 VSS 0.023957f
C14934 a_35502_25545.t85 VSS 0.16147f
C14935 a_35502_25545.n206 VSS 0.087831f
C14936 a_35502_25545.t50 VSS 0.161797f
C14937 a_35502_25545.n207 VSS 0.023957f
C14938 a_35502_25545.t30 VSS 0.16147f
C14939 a_35502_25545.n208 VSS 0.032845f
C14940 a_35502_25545.n209 VSS 0.092213f
C14941 a_35502_25545.n210 VSS 1.68497f
C14942 a_35502_25545.n211 VSS 0.124713f
C14943 a_35502_25545.n212 VSS 0.024358f
C14944 a_35502_25545.n213 VSS 0.02436f
C14945 a_35502_25545.n214 VSS 0.128099f
C14946 a_35502_25545.n215 VSS 0.040603f
C14947 a_35502_25545.n216 VSS 0.128747f
C14948 a_35502_25545.n217 VSS 0.128701f
C14949 a_35502_25545.n218 VSS 0.027673f
C14950 a_35502_25545.n219 VSS 0.02767f
C14951 a_35502_25545.n220 VSS 1.79682f
C14952 a_35502_25545.n221 VSS 1.28081f
C14953 a_35502_25545.n222 VSS 0.094898f
C14954 a_35502_25545.n223 VSS 0.01148f
C14955 a_35502_25545.t39 VSS 0.165101f
C14956 a_35502_25545.n224 VSS 0.134945f
C14957 a_35502_25545.t94 VSS 0.16147f
C14958 a_35502_25545.n225 VSS 0.082553f
C14959 a_35502_25545.n226 VSS 0.018822f
C14960 a_35502_25545.n227 VSS 0.094735f
C14961 a_35502_25545.n228 VSS 0.020553f
C14962 a_35502_25545.n229 VSS 0.01148f
C14963 a_35502_25545.t98 VSS 0.16147f
C14964 a_35502_25545.n230 VSS 0.055026f
C14965 a_35502_25545.t63 VSS 0.16147f
C14966 a_35502_25545.n231 VSS 0.131588f
C14967 a_35502_25545.t67 VSS 0.16147f
C14968 a_35502_25545.n232 VSS 0.106928f
C14969 a_35502_25545.t38 VSS 0.16147f
C14970 a_35502_25545.n233 VSS 0.130219f
C14971 a_35502_25545.n234 VSS 0.020553f
C14972 a_35502_25545.n235 VSS 0.024319f
C14973 a_35502_25545.n236 VSS 0.020553f
C14974 a_35502_25545.t74 VSS 0.16147f
C14975 a_35502_25545.t66 VSS 0.16147f
C14976 a_35502_25545.n237 VSS 0.006509f
C14977 a_35502_25545.n238 VSS 0.098925f
C14978 a_35502_25545.t46 VSS 0.16147f
C14979 a_35502_25545.n239 VSS 0.062479f
C14980 a_35502_25545.t101 VSS 0.16147f
C14981 a_35502_25545.t69 VSS 0.165422f
C14982 a_35502_25545.n240 VSS 0.019526f
C14983 a_35502_25545.n241 VSS 0.01847f
C14984 a_35502_25545.n242 VSS 0.020553f
C14985 a_35502_25545.n243 VSS 0.01148f
C14986 a_35502_25545.n244 VSS 0.035274f
C14987 a_35502_25545.n245 VSS 0.053933f
C14988 a_35502_25545.t88 VSS 0.16147f
C14989 a_35502_25545.n246 VSS 0.130219f
C14990 a_35502_25545.t42 VSS 0.16147f
C14991 a_35502_25545.n247 VSS 0.106928f
C14992 a_35502_25545.t36 VSS 0.16147f
C14993 a_35502_25545.n248 VSS 0.131588f
C14994 a_35502_25545.n249 VSS 0.055026f
C14995 a_35502_25545.n250 VSS 0.094898f
C14996 a_35502_25545.n251 VSS 0.01148f
C14997 a_35502_25545.n252 VSS 0.019526f
C14998 a_35502_25545.n253 VSS 0.018822f
C14999 a_35502_25545.n254 VSS 0.020553f
C15000 a_35502_25545.n255 VSS 0.01148f
C15001 a_35502_25545.n256 VSS 0.020553f
C15002 a_35502_25545.n257 VSS 0.019526f
C15003 a_35502_25545.n258 VSS 0.01847f
C15004 a_35502_25545.t97 VSS 0.16147f
C15005 a_35502_25545.n259 VSS 0.077654f
C15006 a_35502_25545.n260 VSS 0.133088f
C15007 a_35502_25545.t37 VSS 0.16147f
C15008 a_35502_25545.n261 VSS 0.024322f
C15009 a_35502_25545.n262 VSS 0.019526f
C15010 a_35502_25545.t65 VSS 0.16147f
C15011 a_35502_25545.n263 VSS 0.01148f
C15012 a_35502_25545.n264 VSS 0.020553f
C15013 a_35502_25545.n265 VSS 0.020553f
C15014 a_35502_25545.n266 VSS 0.01847f
C15015 a_35502_25545.t89 VSS 0.16147f
C15016 a_35502_25545.n267 VSS 0.062479f
C15017 a_35502_25545.n268 VSS 0.006509f
C15018 a_35502_25545.n269 VSS 0.053933f
C15019 a_35502_25545.n270 VSS 0.035274f
C15020 a_35502_25545.n271 VSS 0.460139f
C15021 a_35502_25545.n272 VSS 1.66281f
C15022 a_35502_25545.n273 VSS 0.121006f
C15023 a_35502_25545.t93 VSS 0.16147f
C15024 a_35502_25545.n274 VSS 0.062479f
C15025 a_35502_25545.n275 VSS 0.017545f
C15026 a_35502_25545.n276 VSS 0.006728f
C15027 a_35502_25545.t90 VSS 0.16147f
C15028 a_35502_25545.n277 VSS 0.079359f
C15029 a_35502_25545.t35 VSS 0.163927f
C15030 a_35502_25545.n278 VSS 0.125171f
C15031 a_35502_25545.n279 VSS 0.086728f
C15032 a_35502_25545.n280 VSS 0.017545f
C15033 a_35502_25545.n281 VSS 0.016667f
C15034 a_35502_25545.n282 VSS 0.016667f
C15035 a_35502_25545.n283 VSS 0.006685f
C15036 a_35502_25545.n284 VSS 0.01148f
C15037 a_35502_25545.n285 VSS 0.095824f
C15038 a_35502_25545.n286 VSS 0.055082f
C15039 a_35502_25545.t55 VSS 0.16147f
C15040 a_35502_25545.n287 VSS 0.131764f
C15041 a_35502_25545.t58 VSS 0.16147f
C15042 a_35502_25545.n288 VSS 0.10628f
C15043 a_35502_25545.t32 VSS 0.16147f
C15044 a_35502_25545.n289 VSS 0.130885f
C15045 a_35502_25545.n290 VSS 0.054994f
C15046 a_35502_25545.n291 VSS 0.036663f
C15047 a_35502_25545.n292 VSS 0.01148f
C15048 a_35502_25545.n293 VSS 0.019614f
C15049 a_35502_25545.t60 VSS 0.16147f
C15050 a_35502_25545.n294 VSS 0.01891f
C15051 a_35502_25545.n295 VSS 0.020646f
C15052 a_35502_25545.n296 VSS 0.01148f
C15053 a_35502_25545.n297 VSS 0.021155f
C15054 a_35502_25545.n298 VSS 0.020097f
C15055 a_35502_25545.n299 VSS 0.01847f
C15056 a_35502_25545.t34 VSS 0.16147f
C15057 a_35502_25545.n300 VSS 0.078447f
C15058 a_35502_25545.n301 VSS 0.132614f
C15059 a_35502_25545.t92 VSS 0.16147f
C15060 a_35502_25545.n302 VSS 0.024924f
C15061 a_35502_25545.n303 VSS 0.021155f
C15062 a_35502_25545.n304 VSS 0.018822f
C15063 a_35502_25545.t70 VSS 0.16147f
C15064 a_35502_25545.n305 VSS 0.062479f
C15065 a_35502_25545.n306 VSS 0.006728f
C15066 a_35502_25545.n307 VSS 0.016667f
C15067 a_35502_25545.n308 VSS 0.017545f
C15068 a_35502_25545.n309 VSS 0.017545f
C15069 a_35502_25545.n310 VSS 0.01148f
C15070 a_35502_25545.n311 VSS 0.006685f
C15071 a_35502_25545.t61 VSS 0.16147f
C15072 a_35502_25545.n312 VSS 0.062479f
C15073 a_35502_25545.n313 VSS 0.055082f
C15074 a_35502_25545.t31 VSS 0.16147f
C15075 a_35502_25545.n314 VSS 0.131764f
C15076 a_35502_25545.t33 VSS 0.16147f
C15077 a_35502_25545.n315 VSS 0.10628f
C15078 a_35502_25545.t84 VSS 0.16147f
C15079 a_35502_25545.n316 VSS 0.130885f
C15080 a_35502_25545.n317 VSS 0.01891f
C15081 a_35502_25545.t64 VSS 0.165184f
C15082 a_35502_25545.t99 VSS 0.16147f
C15083 a_35502_25545.n318 VSS 0.082685f
C15084 a_35502_25545.n319 VSS 0.138167f
C15085 a_35502_25545.n320 VSS 0.0977f
C15086 a_35502_25545.n321 VSS 0.020646f
C15087 a_35502_25545.t43 VSS 0.16147f
C15088 a_35502_25545.n322 VSS 0.054994f
C15089 a_35502_25545.n323 VSS 0.036663f
C15090 a_35502_25545.n324 VSS 0.121006f
C15091 a_35502_25545.n325 VSS 1.66281f
C15092 a_35502_25545.n326 VSS 2.38102f
C15093 a_35502_25545.t17 VSS 0.100583f
C15094 a_35502_25545.t0 VSS 0.093958f
C15095 a_35502_25545.t16 VSS 0.019442f
C15096 a_35502_25545.n327 VSS 0.256639f
C15097 a_35502_25545.t19 VSS 0.074305f
C15098 a_35502_25545.n328 VSS 0.130254f
C15099 a_35502_25545.t14 VSS 0.050299f
C15100 a_35502_25545.t7 VSS 0.048952f
C15101 a_35502_25545.n329 VSS 0.082342f
C15102 a_35502_25545.t5 VSS 0.100915f
C15103 a_35502_25545.t13 VSS 0.093958f
C15104 a_35502_25545.t18 VSS 0.019442f
C15105 a_35502_25545.n330 VSS 0.255029f
C15106 a_35502_25545.n331 VSS 0.057799f
C15107 a_35502_25545.t1 VSS 0.095983f
C15108 a_35502_25545.t9 VSS 0.019442f
C15109 a_35502_25545.n332 VSS 0.119925f
C15110 a_35502_25545.n333 VSS 0.350036f
C15111 a_35502_25545.n334 VSS 0.007407f
C15112 a_35502_25545.t12 VSS 0.074674f
C15113 a_35502_25545.t4 VSS 0.087321f
C15114 a_35502_25545.t11 VSS 0.10138f
C15115 a_35502_25545.t10 VSS 0.09656f
C15116 a_35502_25545.t15 VSS 0.019442f
C15117 a_35502_25545.n335 VSS 0.132071f
C15118 a_35502_25545.t2 VSS 0.100992f
C15119 a_35502_25545.t8 VSS 0.087321f
C15120 a_35502_25545.t6 VSS 0.049237f
C15121 a_35502_25545.n336 VSS 0.016089f
C15122 a_35502_25545.n337 VSS 0.007969f
C15123 a_35502_25545.t3 VSS 0.050405f
C15124 a_35502_25545.n338 VSS 0.087006f
C15125 a_35502_25545.n339 VSS 0.051468f
C15126 a_35502_25545.n340 VSS 0.00574f
C15127 a_35502_25545.n341 VSS 2.05391f
C15128 a_35502_25545.n342 VSS 3.03378f
C15129 a_35502_25545.t23 VSS 0.103728f
C15130 a_35502_25545.t25 VSS 0.080762f
C15131 a_35502_25545.n343 VSS 0.305516f
C15132 a_35502_25545.n344 VSS 0.810129f
C15133 a_35502_25545.t22 VSS 0.199995f
C15134 a_35502_25545.t24 VSS 0.192538f
C15135 a_35502_25545.n345 VSS 0.261445f
C15136 a_35502_25545.t48 VSS 0.192541f
C15137 a_35502_25545.n346 VSS 0.127292f
C15138 a_35502_25545.t91 VSS 0.195808f
C15139 a_35502_25545.n347 VSS 0.13645f
C15140 a_35502_25545.n348 VSS 0.178301f
C15141 a_35502_25545.t71 VSS 0.199995f
C15142 a_35502_25545.t62 VSS 0.192538f
C15143 a_35502_25545.n349 VSS 0.261445f
C15144 a_35502_25545.t26 VSS 0.192541f
C15145 a_35502_25545.n350 VSS 0.127292f
C15146 a_35502_25545.t20 VSS 0.195808f
C15147 a_35502_25545.n351 VSS 0.13645f
C15148 a_35502_25545.n352 VSS 0.342272f
C15149 a_35502_25545.n353 VSS 0.364067f
C15150 a_35502_25545.t27 VSS 0.102707f
C15151 a_36032_n36322.t3 VSS 0.792603f
C15152 a_36032_n36322.t2 VSS 0.676033f
C15153 a_36032_n36322.n0 VSS 8.260099f
C15154 a_36032_n36322.t1 VSS 0.752866f
C15155 a_36032_n36322.n1 VSS 8.13687f
C15156 a_36032_n36322.t0 VSS 0.781529f
C15157 a_53829_n36382.n0 VSS 2.53786f
C15158 a_53829_n36382.n1 VSS 9.92737f
C15159 a_53829_n36382.n2 VSS 0.941684f
C15160 a_53829_n36382.n3 VSS 1.60401f
C15161 a_53829_n36382.n4 VSS 5.88446f
C15162 a_53829_n36382.n5 VSS 7.95021f
C15163 a_53829_n36382.n6 VSS 0.911784f
C15164 a_53829_n36382.t12 VSS 0.572572f
C15165 a_53829_n36382.t13 VSS 0.605718f
C15166 a_53829_n36382.t22 VSS 0.572368f
C15167 a_53829_n36382.t6 VSS 0.347085f
C15168 a_53829_n36382.t0 VSS 0.599022f
C15169 a_53829_n36382.t2 VSS 0.321538f
C15170 a_53829_n36382.t3 VSS 0.32663f
C15171 a_53829_n36382.t1 VSS 0.49853f
C15172 a_53829_n36382.t5 VSS 0.52604f
C15173 a_53829_n36382.t21 VSS 0.563936f
C15174 a_53829_n36382.t10 VSS 0.563895f
C15175 a_53829_n36382.t16 VSS 0.561709f
C15176 a_53829_n36382.t11 VSS 0.561709f
C15177 a_53829_n36382.t17 VSS 0.561709f
C15178 a_53829_n36382.t20 VSS 0.561709f
C15179 a_53829_n36382.t23 VSS 0.563801f
C15180 a_53829_n36382.t9 VSS 0.563957f
C15181 a_53829_n36382.t15 VSS 0.561709f
C15182 a_53829_n36382.t14 VSS 0.561709f
C15183 a_53829_n36382.t18 VSS 0.561709f
C15184 a_53829_n36382.t8 VSS 0.571948f
C15185 a_53829_n36382.t19 VSS 0.561709f
C15186 a_53829_n36382.t7 VSS 0.523325f
C15187 a_53829_n36382.n7 VSS 0.912676f
C15188 a_53829_n36382.t4 VSS 0.315883f
C15189 a_100820_10448.t0 VSS 20.5853f
C15190 a_100820_10448.t3 VSS 1.77451f
C15191 a_100820_10448.t9 VSS 0.34777f
C15192 a_100820_10448.t2 VSS 0.330207f
C15193 a_100820_10448.t1 VSS 0.329925f
C15194 a_100820_10448.t14 VSS 0.568066f
C15195 a_100820_10448.t17 VSS 0.544019f
C15196 a_100820_10448.t23 VSS 0.544019f
C15197 a_100820_10448.t4 VSS 0.562597f
C15198 a_100820_10448.t18 VSS 0.568066f
C15199 a_100820_10448.t12 VSS 0.544019f
C15200 a_100820_10448.t10 VSS 0.568066f
C15201 a_100820_10448.t15 VSS 0.544019f
C15202 a_100820_10448.t19 VSS 0.544019f
C15203 a_100820_10448.t21 VSS 0.562597f
C15204 a_100820_10448.t11 VSS 0.34777f
C15205 a_100820_10448.t7 VSS 0.30485f
C15206 a_100820_10448.t6 VSS 0.562597f
C15207 a_100820_10448.t13 VSS 0.544019f
C15208 a_100820_10448.t8 VSS 0.568066f
C15209 a_100820_10448.t16 VSS 0.544019f
C15210 a_100820_10448.t22 VSS 0.562597f
C15211 a_100820_10448.t20 VSS 0.544019f
C15212 a_100820_10448.t5 VSS 0.30485f
C15213 a_31284_4481.t1 VSS 5.04925f
C15214 a_31284_4481.t2 VSS 40.732197f
C15215 a_31284_4481.t0 VSS 37.7185f
C15216 a_30324_4421.t0 VSS 25.4694f
C15217 a_30324_4421.t1 VSS 13.3715f
C15218 a_30324_4421.t2 VSS 1.15913f
C15219 a_100820_11614.n0 VSS 0.727613f
C15220 a_100820_11614.n1 VSS 11.477901f
C15221 a_100820_11614.n2 VSS 11.550099f
C15222 a_100820_11614.t20 VSS 0.458761f
C15223 a_100820_11614.t12 VSS 0.458717f
C15224 a_100820_11614.t1 VSS 0.509737f
C15225 a_100820_11614.t3 VSS 0.260912f
C15226 a_100820_11614.t2 VSS 0.278471f
C15227 a_100820_11614.t10 VSS 0.452124f
C15228 a_100820_11614.t14 VSS 0.452124f
C15229 a_100820_11614.t15 VSS 0.450255f
C15230 a_100820_11614.t11 VSS 0.450255f
C15231 a_100820_11614.t18 VSS 0.450255f
C15232 a_100820_11614.t16 VSS 0.458761f
C15233 a_100820_11614.t21 VSS 0.450255f
C15234 a_100820_11614.t17 VSS 0.452124f
C15235 a_100820_11614.t8 VSS 0.452124f
C15236 a_100820_11614.t9 VSS 0.450255f
C15237 a_100820_11614.t19 VSS 0.450255f
C15238 a_100820_11614.t23 VSS 0.450255f
C15239 a_100820_11614.t22 VSS 0.458717f
C15240 a_100820_11614.t13 VSS 0.450255f
C15241 a_100820_11614.t6 VSS 0.410823f
C15242 a_100820_11614.t5 VSS 0.242329f
C15243 a_100820_11614.t4 VSS 0.273794f
C15244 a_100820_11614.t7 VSS 0.423369f
C15245 a_100820_11614.t0 VSS 0.399525f
C15246 a_57977_n12421.t0 VSS 59.2863f
C15247 a_57977_n12421.t2 VSS 2.43373f
C15248 a_57977_n12421.t1 VSS 31.18f
C15249 a_52635_49681.n0 VSS 2.5012f
C15250 a_52635_49681.n1 VSS 2.18773f
C15251 a_52635_49681.n2 VSS 2.5012f
C15252 a_52635_49681.n3 VSS 2.18779f
C15253 a_52635_49681.n4 VSS 1.41275f
C15254 a_52635_49681.n5 VSS 2.60963f
C15255 a_52635_49681.n6 VSS 1.8458f
C15256 a_52635_49681.n7 VSS 1.76011f
C15257 a_52635_49681.n8 VSS 2.60963f
C15258 a_52635_49681.n9 VSS 1.8458f
C15259 a_52635_49681.n10 VSS 1.34268f
C15260 a_52635_49681.n11 VSS 1.41272f
C15261 a_52635_49681.t92 VSS 0.096749f
C15262 a_52635_49681.t126 VSS 0.437557f
C15263 a_52635_49681.t121 VSS 0.096749f
C15264 a_52635_49681.t93 VSS 0.096749f
C15265 a_52635_49681.n12 VSS 0.450336f
C15266 a_52635_49681.t136 VSS 0.79292f
C15267 a_52635_49681.n13 VSS 5.77891f
C15268 a_52635_49681.n14 VSS 4.24962f
C15269 a_52635_49681.t88 VSS 0.096749f
C15270 a_52635_49681.t128 VSS 0.096749f
C15271 a_52635_49681.n15 VSS 0.929945f
C15272 a_52635_49681.t111 VSS 0.435002f
C15273 a_52635_49681.n16 VSS 2.49496f
C15274 a_52635_49681.n17 VSS 2.59005f
C15275 a_52635_49681.t170 VSS 0.096749f
C15276 a_52635_49681.t115 VSS 0.096749f
C15277 a_52635_49681.n18 VSS 0.446763f
C15278 a_52635_49681.n19 VSS 2.1917f
C15279 a_52635_49681.t175 VSS 0.435002f
C15280 a_52635_49681.n20 VSS 2.0431f
C15281 a_52635_49681.t113 VSS 0.254893f
C15282 a_52635_49681.t140 VSS 0.271406f
C15283 a_52635_49681.n21 VSS 1.03037f
C15284 a_52635_49681.t143 VSS 0.096749f
C15285 a_52635_49681.t112 VSS 0.096749f
C15286 a_52635_49681.n22 VSS 0.245505f
C15287 a_52635_49681.t171 VSS 0.096749f
C15288 a_52635_49681.t139 VSS 0.096749f
C15289 a_52635_49681.n23 VSS 0.264956f
C15290 a_52635_49681.n24 VSS 0.672455f
C15291 a_52635_49681.n25 VSS 0.560391f
C15292 a_52635_49681.t135 VSS 0.254893f
C15293 a_52635_49681.t156 VSS 0.271406f
C15294 a_52635_49681.n26 VSS 1.02935f
C15295 a_52635_49681.t91 VSS 0.096749f
C15296 a_52635_49681.t166 VSS 0.096749f
C15297 a_52635_49681.n27 VSS 0.245505f
C15298 a_52635_49681.t108 VSS 0.096749f
C15299 a_52635_49681.t97 VSS 0.096749f
C15300 a_52635_49681.n28 VSS 0.264956f
C15301 a_52635_49681.n29 VSS 0.672455f
C15302 a_52635_49681.n30 VSS 0.710427f
C15303 a_52635_49681.t133 VSS 0.254893f
C15304 a_52635_49681.t150 VSS 0.271406f
C15305 a_52635_49681.n31 VSS 0.855769f
C15306 a_52635_49681.n32 VSS 0.783311f
C15307 a_52635_49681.t129 VSS 0.254893f
C15308 a_52635_49681.t147 VSS 0.271406f
C15309 a_52635_49681.n33 VSS 0.859332f
C15310 a_52635_49681.n34 VSS 0.662159f
C15311 a_52635_49681.n35 VSS 0.266191f
C15312 a_52635_49681.t155 VSS 0.096749f
C15313 a_52635_49681.t125 VSS 0.096749f
C15314 a_52635_49681.n36 VSS 0.245505f
C15315 a_52635_49681.t89 VSS 0.096749f
C15316 a_52635_49681.t145 VSS 0.096749f
C15317 a_52635_49681.n37 VSS 0.264956f
C15318 a_52635_49681.n38 VSS 0.672455f
C15319 a_52635_49681.n39 VSS 0.373952f
C15320 a_52635_49681.t109 VSS 0.254893f
C15321 a_52635_49681.t138 VSS 0.271406f
C15322 a_52635_49681.n40 VSS 0.868543f
C15323 a_52635_49681.n41 VSS 0.797505f
C15324 a_52635_49681.t124 VSS 0.254893f
C15325 a_52635_49681.t144 VSS 0.271406f
C15326 a_52635_49681.n42 VSS 0.868543f
C15327 a_52635_49681.n43 VSS 0.797478f
C15328 a_52635_49681.t163 VSS 0.096749f
C15329 a_52635_49681.t134 VSS 0.096749f
C15330 a_52635_49681.n44 VSS 0.245505f
C15331 a_52635_49681.t96 VSS 0.096749f
C15332 a_52635_49681.t153 VSS 0.096749f
C15333 a_52635_49681.n45 VSS 0.264956f
C15334 a_52635_49681.n46 VSS 0.672455f
C15335 a_52635_49681.n47 VSS 0.525201f
C15336 a_52635_49681.t119 VSS 0.254893f
C15337 a_52635_49681.t142 VSS 0.271406f
C15338 a_52635_49681.n48 VSS 0.855769f
C15339 a_52635_49681.n49 VSS 0.783311f
C15340 a_52635_49681.t98 VSS 0.254893f
C15341 a_52635_49681.t116 VSS 0.271406f
C15342 a_52635_49681.n50 VSS 0.859332f
C15343 a_52635_49681.n51 VSS 0.662159f
C15344 a_52635_49681.n52 VSS 0.266191f
C15345 a_52635_49681.n53 VSS 6.30381f
C15346 a_52635_49681.n54 VSS 4.22046f
C15347 a_52635_49681.n55 VSS 6.23036f
C15348 a_52635_49681.t158 VSS 0.096749f
C15349 a_52635_49681.t146 VSS 0.096749f
C15350 a_52635_49681.n56 VSS 0.450336f
C15351 a_52635_49681.t100 VSS 0.437557f
C15352 a_52635_49681.t99 VSS 0.096749f
C15353 a_52635_49681.t159 VSS 0.096749f
C15354 a_52635_49681.n57 VSS 0.450336f
C15355 a_52635_49681.t102 VSS 0.79292f
C15356 a_52635_49681.n58 VSS 3.70414f
C15357 a_52635_49681.n59 VSS 4.69402f
C15358 a_52635_49681.t46 VSS 0.38248f
C15359 a_52635_49681.t52 VSS 0.096749f
C15360 a_52635_49681.t25 VSS 0.096749f
C15361 a_52635_49681.n60 VSS 0.385894f
C15362 a_52635_49681.t27 VSS 0.38248f
C15363 a_52635_49681.t45 VSS 0.096749f
C15364 a_52635_49681.t15 VSS 0.096749f
C15365 a_52635_49681.n61 VSS 0.885379f
C15366 a_52635_49681.t31 VSS 0.38248f
C15367 a_52635_49681.t55 VSS 0.096749f
C15368 a_52635_49681.t26 VSS 0.096749f
C15369 a_52635_49681.n62 VSS 0.885379f
C15370 a_52635_49681.n63 VSS 2.61926f
C15371 a_52635_49681.t57 VSS 0.38248f
C15372 a_52635_49681.t62 VSS 0.096749f
C15373 a_52635_49681.t29 VSS 0.096749f
C15374 a_52635_49681.n64 VSS 0.385894f
C15375 a_52635_49681.n65 VSS 6.50148f
C15376 a_52635_49681.t20 VSS 0.096749f
C15377 a_52635_49681.t65 VSS 0.096749f
C15378 a_52635_49681.n66 VSS 0.290163f
C15379 a_52635_49681.t18 VSS 0.096749f
C15380 a_52635_49681.t64 VSS 0.096749f
C15381 a_52635_49681.n67 VSS 0.224889f
C15382 a_52635_49681.n68 VSS 0.667866f
C15383 a_52635_49681.n69 VSS 0.579701f
C15384 a_52635_49681.t21 VSS 0.096749f
C15385 a_52635_49681.t34 VSS 0.096749f
C15386 a_52635_49681.n70 VSS 0.290163f
C15387 a_52635_49681.t19 VSS 0.096749f
C15388 a_52635_49681.t33 VSS 0.096749f
C15389 a_52635_49681.n71 VSS 0.224889f
C15390 a_52635_49681.n72 VSS 0.667866f
C15391 a_52635_49681.n73 VSS 1.04211f
C15392 a_52635_49681.t11 VSS 0.096749f
C15393 a_52635_49681.t56 VSS 0.096749f
C15394 a_52635_49681.n74 VSS 0.290163f
C15395 a_52635_49681.t10 VSS 0.096749f
C15396 a_52635_49681.t53 VSS 0.096749f
C15397 a_52635_49681.n75 VSS 0.224889f
C15398 a_52635_49681.n76 VSS 0.667866f
C15399 a_52635_49681.n77 VSS 1.04214f
C15400 a_52635_49681.t79 VSS 0.096749f
C15401 a_52635_49681.t8 VSS 0.096749f
C15402 a_52635_49681.n78 VSS 0.290163f
C15403 a_52635_49681.t76 VSS 0.096749f
C15404 a_52635_49681.t5 VSS 0.096749f
C15405 a_52635_49681.n79 VSS 0.224889f
C15406 a_52635_49681.n80 VSS 0.667866f
C15407 a_52635_49681.n81 VSS 1.02776f
C15408 a_52635_49681.t54 VSS 0.096749f
C15409 a_52635_49681.t77 VSS 0.096749f
C15410 a_52635_49681.n82 VSS 0.290163f
C15411 a_52635_49681.t51 VSS 0.096749f
C15412 a_52635_49681.t75 VSS 0.096749f
C15413 a_52635_49681.n83 VSS 0.224889f
C15414 a_52635_49681.n84 VSS 0.931197f
C15415 a_52635_49681.t83 VSS 0.096749f
C15416 a_52635_49681.t37 VSS 0.096749f
C15417 a_52635_49681.n85 VSS 0.290163f
C15418 a_52635_49681.t82 VSS 0.096749f
C15419 a_52635_49681.t36 VSS 0.096749f
C15420 a_52635_49681.n86 VSS 0.224889f
C15421 a_52635_49681.n87 VSS 0.667866f
C15422 a_52635_49681.n88 VSS 1.34555f
C15423 a_52635_49681.t6 VSS 0.096749f
C15424 a_52635_49681.t87 VSS 0.096749f
C15425 a_52635_49681.n89 VSS 0.290163f
C15426 a_52635_49681.t4 VSS 0.096749f
C15427 a_52635_49681.t86 VSS 0.096749f
C15428 a_52635_49681.n90 VSS 0.224889f
C15429 a_52635_49681.n91 VSS 0.667866f
C15430 a_52635_49681.n92 VSS 1.04211f
C15431 a_52635_49681.t24 VSS 0.096749f
C15432 a_52635_49681.t61 VSS 0.096749f
C15433 a_52635_49681.n93 VSS 0.290163f
C15434 a_52635_49681.t23 VSS 0.096749f
C15435 a_52635_49681.t60 VSS 0.096749f
C15436 a_52635_49681.n94 VSS 0.224889f
C15437 a_52635_49681.n95 VSS 0.667866f
C15438 a_52635_49681.n96 VSS 0.276895f
C15439 a_52635_49681.n97 VSS 0.813686f
C15440 a_52635_49681.n98 VSS 5.7089f
C15441 a_52635_49681.t41 VSS 0.096749f
C15442 a_52635_49681.t47 VSS 0.096749f
C15443 a_52635_49681.n99 VSS 0.38674f
C15444 a_52635_49681.n100 VSS 1.41191f
C15445 a_52635_49681.t17 VSS 0.383187f
C15446 a_52635_49681.n101 VSS 1.82711f
C15447 a_52635_49681.t2 VSS 0.742971f
C15448 a_52635_49681.t22 VSS 0.096749f
C15449 a_52635_49681.t40 VSS 0.096749f
C15450 a_52635_49681.n102 VSS 0.38674f
C15451 a_52635_49681.n103 VSS 2.61788f
C15452 a_52635_49681.n104 VSS 1.83604f
C15453 a_52635_49681.n105 VSS 4.09621f
C15454 a_52635_49681.n106 VSS 3.67005f
C15455 a_52635_49681.n107 VSS 1.83781f
C15456 a_52635_49681.n108 VSS 4.06839f
C15457 a_52635_49681.t48 VSS 0.096749f
C15458 a_52635_49681.t70 VSS 0.096749f
C15459 a_52635_49681.n109 VSS 0.290163f
C15460 a_52635_49681.t43 VSS 0.096749f
C15461 a_52635_49681.t66 VSS 0.096749f
C15462 a_52635_49681.n110 VSS 0.224889f
C15463 a_52635_49681.n111 VSS 0.931197f
C15464 a_52635_49681.t74 VSS 0.096749f
C15465 a_52635_49681.t35 VSS 0.096749f
C15466 a_52635_49681.n112 VSS 0.290163f
C15467 a_52635_49681.t68 VSS 0.096749f
C15468 a_52635_49681.t30 VSS 0.096749f
C15469 a_52635_49681.n113 VSS 0.224889f
C15470 a_52635_49681.n114 VSS 0.667866f
C15471 a_52635_49681.n115 VSS 1.34555f
C15472 a_52635_49681.t84 VSS 0.096749f
C15473 a_52635_49681.t78 VSS 0.096749f
C15474 a_52635_49681.n116 VSS 0.290163f
C15475 a_52635_49681.t72 VSS 0.096749f
C15476 a_52635_49681.t69 VSS 0.096749f
C15477 a_52635_49681.n117 VSS 0.224889f
C15478 a_52635_49681.n118 VSS 0.667866f
C15479 a_52635_49681.n119 VSS 1.04211f
C15480 a_52635_49681.t16 VSS 0.096749f
C15481 a_52635_49681.t58 VSS 0.096749f
C15482 a_52635_49681.n120 VSS 0.290163f
C15483 a_52635_49681.t7 VSS 0.096749f
C15484 a_52635_49681.t50 VSS 0.096749f
C15485 a_52635_49681.n121 VSS 0.224889f
C15486 a_52635_49681.n122 VSS 0.667866f
C15487 a_52635_49681.n123 VSS 0.276895f
C15488 a_52635_49681.n124 VSS 0.813686f
C15489 a_52635_49681.t71 VSS 0.096749f
C15490 a_52635_49681.t85 VSS 0.096749f
C15491 a_52635_49681.n125 VSS 0.290163f
C15492 a_52635_49681.t67 VSS 0.096749f
C15493 a_52635_49681.t73 VSS 0.096749f
C15494 a_52635_49681.n126 VSS 0.224889f
C15495 a_52635_49681.n127 VSS 0.667866f
C15496 a_52635_49681.n128 VSS 1.02776f
C15497 a_52635_49681.t3 VSS 0.096749f
C15498 a_52635_49681.t49 VSS 0.096749f
C15499 a_52635_49681.n129 VSS 0.290163f
C15500 a_52635_49681.t80 VSS 0.096749f
C15501 a_52635_49681.t44 VSS 0.096749f
C15502 a_52635_49681.n130 VSS 0.224889f
C15503 a_52635_49681.n131 VSS 0.667866f
C15504 a_52635_49681.n132 VSS 1.04214f
C15505 a_52635_49681.t13 VSS 0.096749f
C15506 a_52635_49681.t32 VSS 0.096749f
C15507 a_52635_49681.n133 VSS 0.290163f
C15508 a_52635_49681.t1 VSS 0.096749f
C15509 a_52635_49681.t28 VSS 0.096749f
C15510 a_52635_49681.n134 VSS 0.224889f
C15511 a_52635_49681.n135 VSS 0.667866f
C15512 a_52635_49681.n136 VSS 1.04211f
C15513 a_52635_49681.t12 VSS 0.096749f
C15514 a_52635_49681.t63 VSS 0.096749f
C15515 a_52635_49681.n137 VSS 0.290163f
C15516 a_52635_49681.t0 VSS 0.096749f
C15517 a_52635_49681.t59 VSS 0.096749f
C15518 a_52635_49681.n138 VSS 0.224889f
C15519 a_52635_49681.n139 VSS 0.667866f
C15520 a_52635_49681.n140 VSS 0.579701f
C15521 a_52635_49681.n141 VSS 3.73436f
C15522 a_52635_49681.n142 VSS 5.4662f
C15523 a_52635_49681.t39 VSS 0.096749f
C15524 a_52635_49681.t42 VSS 0.096749f
C15525 a_52635_49681.n143 VSS 0.38674f
C15526 a_52635_49681.n144 VSS 1.41191f
C15527 a_52635_49681.t9 VSS 0.383187f
C15528 a_52635_49681.n145 VSS 1.82711f
C15529 a_52635_49681.t81 VSS 0.742971f
C15530 a_52635_49681.t14 VSS 0.096749f
C15531 a_52635_49681.t38 VSS 0.096749f
C15532 a_52635_49681.n146 VSS 0.38674f
C15533 a_52635_49681.n147 VSS 2.61788f
C15534 a_52635_49681.n148 VSS 1.83604f
C15535 a_52635_49681.n149 VSS 4.41262f
C15536 a_52635_49681.n150 VSS 6.29237f
C15537 a_52635_49681.n151 VSS 4.92683f
C15538 a_52635_49681.n152 VSS 1.8367f
C15539 a_52635_49681.n153 VSS 5.00434f
C15540 a_52635_49681.t154 VSS 0.254893f
C15541 a_52635_49681.t107 VSS 0.271406f
C15542 a_52635_49681.n154 VSS 1.03037f
C15543 a_52635_49681.t95 VSS 0.096749f
C15544 a_52635_49681.t152 VSS 0.096749f
C15545 a_52635_49681.n155 VSS 0.245505f
C15546 a_52635_49681.t141 VSS 0.096749f
C15547 a_52635_49681.t106 VSS 0.096749f
C15548 a_52635_49681.n156 VSS 0.264956f
C15549 a_52635_49681.n157 VSS 0.672455f
C15550 a_52635_49681.n158 VSS 0.560391f
C15551 a_52635_49681.t173 VSS 0.254893f
C15552 a_52635_49681.t131 VSS 0.271406f
C15553 a_52635_49681.n159 VSS 1.02935f
C15554 a_52635_49681.t132 VSS 0.096749f
C15555 a_52635_49681.t104 VSS 0.096749f
C15556 a_52635_49681.n160 VSS 0.245505f
C15557 a_52635_49681.t90 VSS 0.096749f
C15558 a_52635_49681.t161 VSS 0.096749f
C15559 a_52635_49681.n161 VSS 0.264956f
C15560 a_52635_49681.n162 VSS 0.672455f
C15561 a_52635_49681.n163 VSS 0.710427f
C15562 a_52635_49681.t169 VSS 0.254893f
C15563 a_52635_49681.t127 VSS 0.271406f
C15564 a_52635_49681.n164 VSS 0.855769f
C15565 a_52635_49681.n165 VSS 0.783311f
C15566 a_52635_49681.t168 VSS 0.254893f
C15567 a_52635_49681.t123 VSS 0.271406f
C15568 a_52635_49681.n166 VSS 0.859332f
C15569 a_52635_49681.n167 VSS 0.662159f
C15570 a_52635_49681.n168 VSS 0.266191f
C15571 a_52635_49681.t101 VSS 0.096749f
C15572 a_52635_49681.t165 VSS 0.096749f
C15573 a_52635_49681.n169 VSS 0.245505f
C15574 a_52635_49681.t148 VSS 0.096749f
C15575 a_52635_49681.t118 VSS 0.096749f
C15576 a_52635_49681.n170 VSS 0.264956f
C15577 a_52635_49681.n171 VSS 0.672455f
C15578 a_52635_49681.n172 VSS 0.373952f
C15579 a_52635_49681.t149 VSS 0.254893f
C15580 a_52635_49681.t105 VSS 0.271406f
C15581 a_52635_49681.n173 VSS 0.868543f
C15582 a_52635_49681.n174 VSS 0.797505f
C15583 a_52635_49681.t164 VSS 0.254893f
C15584 a_52635_49681.t117 VSS 0.271406f
C15585 a_52635_49681.n175 VSS 0.868543f
C15586 a_52635_49681.n176 VSS 0.797478f
C15587 a_52635_49681.t103 VSS 0.096749f
C15588 a_52635_49681.t172 VSS 0.096749f
C15589 a_52635_49681.n177 VSS 0.245505f
C15590 a_52635_49681.t160 VSS 0.096749f
C15591 a_52635_49681.t130 VSS 0.096749f
C15592 a_52635_49681.n178 VSS 0.264956f
C15593 a_52635_49681.n179 VSS 0.672455f
C15594 a_52635_49681.n180 VSS 0.525201f
C15595 a_52635_49681.t162 VSS 0.254893f
C15596 a_52635_49681.t114 VSS 0.271406f
C15597 a_52635_49681.n181 VSS 0.855769f
C15598 a_52635_49681.n182 VSS 0.783311f
C15599 a_52635_49681.t137 VSS 0.254893f
C15600 a_52635_49681.t94 VSS 0.271406f
C15601 a_52635_49681.n183 VSS 0.859332f
C15602 a_52635_49681.n184 VSS 0.662159f
C15603 a_52635_49681.n185 VSS 0.266191f
C15604 a_52635_49681.n186 VSS 4.24962f
C15605 a_52635_49681.n187 VSS 3.92865f
C15606 a_52635_49681.t120 VSS 0.435002f
C15607 a_52635_49681.n188 VSS 1.44115f
C15608 a_52635_49681.t110 VSS 0.096749f
C15609 a_52635_49681.t157 VSS 0.096749f
C15610 a_52635_49681.n189 VSS 0.446763f
C15611 a_52635_49681.n190 VSS 2.1917f
C15612 a_52635_49681.t122 VSS 0.096749f
C15613 a_52635_49681.t167 VSS 0.096749f
C15614 a_52635_49681.n191 VSS 0.929945f
C15615 a_52635_49681.t151 VSS 0.435002f
C15616 a_52635_49681.n192 VSS 2.49496f
C15617 a_52635_49681.n193 VSS 1.8377f
C15618 a_52635_49681.n194 VSS 3.55414f
C15619 a_52635_49681.n195 VSS 3.66664f
C15620 a_52635_49681.n196 VSS 1.8367f
C15621 a_52635_49681.n197 VSS 0.450336f
C15622 a_52635_49681.t174 VSS 0.096749f
C15623 VDD.n0 VSS 0.250507f
C15624 VDD.n1 VSS 0.309686f
C15625 VDD.n3 VSS 0.018249f
C15626 VDD.n5 VSS 0.01487f
C15627 VDD.n6 VSS 2.53555f
C15628 VDD.n7 VSS 1.05204f
C15629 VDD.n8 VSS 0.009688f
C15630 VDD.n9 VSS 0.101314f
C15631 VDD.t2665 VSS 0.066856f
C15632 VDD.n11 VSS 0.14405f
C15633 VDD.t1468 VSS 0.025104f
C15634 VDD.n12 VSS 0.087217f
C15635 VDD.n13 VSS 1.05032f
C15636 VDD.n14 VSS 0.207221f
C15637 VDD.t836 VSS 1.45905f
C15638 VDD.t1484 VSS 1.96535f
C15639 VDD.t331 VSS 1.96535f
C15640 VDD.t329 VSS 1.36988f
C15641 VDD.n15 VSS 0.645798f
C15642 VDD.t1221 VSS 1.45794f
C15643 VDD.n16 VSS 0.208771f
C15644 VDD.n17 VSS 0.206947f
C15645 VDD.t4045 VSS 0.028519f
C15646 VDD.t2654 VSS 0.028519f
C15647 VDD.n18 VSS 0.009191f
C15648 VDD.t3873 VSS 0.028519f
C15649 VDD.t2865 VSS 0.028519f
C15650 VDD.n19 VSS 0.009191f
C15651 VDD.n20 VSS 0.471397f
C15652 VDD.t3449 VSS 0.028519f
C15653 VDD.t1968 VSS 0.028519f
C15654 VDD.n21 VSS 0.009191f
C15655 VDD.t3448 VSS 0.066856f
C15656 VDD.t3308 VSS 0.066856f
C15657 VDD.t3806 VSS 0.066856f
C15658 VDD.t3638 VSS 0.066856f
C15659 VDD.t3807 VSS 0.028519f
C15660 VDD.t2417 VSS 0.028519f
C15661 VDD.n22 VSS 0.009191f
C15662 VDD.t1220 VSS 0.066856f
C15663 VDD.t1088 VSS 0.066856f
C15664 VDD.t1222 VSS 0.028519f
C15665 VDD.t3945 VSS 0.028519f
C15666 VDD.n23 VSS 0.009191f
C15667 VDD.t1292 VSS 0.066856f
C15668 VDD.n24 VSS 0.125227f
C15669 VDD.t3917 VSS 0.025104f
C15670 VDD.t847 VSS 0.066856f
C15671 VDD.n25 VSS 0.125227f
C15672 VDD.t4267 VSS 0.025104f
C15673 VDD.n26 VSS 0.099723f
C15674 VDD.t4135 VSS 0.028519f
C15675 VDD.t4329 VSS 0.028519f
C15676 VDD.n27 VSS 0.009191f
C15677 VDD.t3975 VSS 0.028519f
C15678 VDD.t2961 VSS 0.028519f
C15679 VDD.n28 VSS 0.009191f
C15680 VDD.n29 VSS 0.471397f
C15681 VDD.n30 VSS 0.207221f
C15682 VDD.n31 VSS 0.208771f
C15683 VDD.n32 VSS 0.206947f
C15684 VDD.t1572 VSS 1.96535f
C15685 VDD.t1293 VSS 1.96535f
C15686 VDD.t1542 VSS 1.36988f
C15687 VDD.n33 VSS 0.645798f
C15688 VDD.n34 VSS 0.595476f
C15689 VDD.t848 VSS 1.31955f
C15690 VDD.t1906 VSS 1.96535f
C15691 VDD.t1158 VSS 1.96535f
C15692 VDD.t1886 VSS 1.45794f
C15693 VDD.n35 VSS 0.865258f
C15694 VDD.n36 VSS 0.902999f
C15695 VDD.t640 VSS 0.028519f
C15696 VDD.t894 VSS 0.028519f
C15697 VDD.n37 VSS 0.009191f
C15698 VDD.t4401 VSS 0.028519f
C15699 VDD.t1651 VSS 0.028519f
C15700 VDD.n38 VSS 0.009191f
C15701 VDD.n39 VSS 0.475536f
C15702 VDD.t4231 VSS 0.028519f
C15703 VDD.t4405 VSS 0.028519f
C15704 VDD.n40 VSS 0.009191f
C15705 VDD.t3821 VSS 0.028519f
C15706 VDD.t1078 VSS 0.028519f
C15707 VDD.n41 VSS 0.009191f
C15708 VDD.n42 VSS 0.528101f
C15709 VDD.n43 VSS 0.208771f
C15710 VDD.n44 VSS 0.207221f
C15711 VDD.t2242 VSS 0.066856f
C15712 VDD.n45 VSS 0.125227f
C15713 VDD.t1999 VSS 0.025104f
C15714 VDD.n46 VSS 0.035132f
C15715 VDD.t3129 VSS 0.025104f
C15716 VDD.t1494 VSS 0.066856f
C15717 VDD.n47 VSS 0.125227f
C15718 VDD.t3153 VSS 0.025104f
C15719 VDD.t3152 VSS 0.066856f
C15720 VDD.n48 VSS 0.125227f
C15721 VDD.n49 VSS 0.101294f
C15722 VDD.n50 VSS 0.016021f
C15723 VDD.t1495 VSS 0.025104f
C15724 VDD.n51 VSS 0.081176f
C15725 VDD.n52 VSS 0.048151f
C15726 VDD.n53 VSS 0.083673f
C15727 VDD.t3128 VSS 0.066856f
C15728 VDD.n54 VSS 0.125227f
C15729 VDD.n55 VSS 0.006598f
C15730 VDD.n56 VSS 0.010188f
C15731 VDD.t531 VSS 0.020387f
C15732 VDD.t534 VSS 0.022137f
C15733 VDD.n57 VSS 0.069721f
C15734 VDD.n58 VSS 0.040089f
C15735 VDD.t539 VSS 0.022115f
C15736 VDD.t536 VSS 0.020371f
C15737 VDD.n59 VSS 0.027128f
C15738 VDD.n60 VSS 0.036577f
C15739 VDD.n61 VSS 0.044801f
C15740 VDD.n62 VSS 0.278297f
C15741 VDD.n63 VSS 0.040089f
C15742 VDD.t532 VSS 0.020387f
C15743 VDD.n64 VSS 0.049653f
C15744 VDD.t533 VSS 0.017093f
C15745 VDD.n65 VSS 0.042104f
C15746 VDD.n66 VSS 0.069461f
C15747 VDD.t538 VSS 0.017093f
C15748 VDD.n67 VSS 0.035483f
C15749 VDD.t537 VSS 0.020371f
C15750 VDD.n68 VSS 0.027128f
C15751 VDD.n69 VSS 0.016538f
C15752 VDD.n70 VSS 0.027213f
C15753 VDD.n71 VSS 0.204333f
C15754 VDD.n72 VSS 0.030906f
C15755 VDD.t1854 VSS 0.066856f
C15756 VDD.n73 VSS 0.045867f
C15757 VDD.n74 VSS 0.015693f
C15758 VDD.n75 VSS 0.010881f
C15759 VDD.n76 VSS 0.044227f
C15760 VDD.n77 VSS 0.094696f
C15761 VDD.n78 VSS 0.016021f
C15762 VDD.t1855 VSS 0.025104f
C15763 VDD.n79 VSS 0.08403f
C15764 VDD.t4230 VSS 0.066856f
C15765 VDD.t3820 VSS 0.066856f
C15766 VDD.t1077 VSS 0.066856f
C15767 VDD.t4404 VSS 0.066856f
C15768 VDD.n80 VSS 0.696076f
C15769 VDD.t4550 VSS 0.066856f
C15770 VDD.t4220 VSS 0.066856f
C15771 VDD.t1417 VSS 0.066856f
C15772 VDD.t628 VSS 0.066856f
C15773 VDD.n81 VSS 0.696076f
C15774 VDD.t4551 VSS 0.028519f
C15775 VDD.t630 VSS 0.028519f
C15776 VDD.n82 VSS 0.009191f
C15777 VDD.t4221 VSS 0.028519f
C15778 VDD.t1418 VSS 0.028519f
C15779 VDD.n83 VSS 0.009191f
C15780 VDD.n84 VSS 0.650522f
C15781 VDD.t2033 VSS 0.066856f
C15782 VDD.t1612 VSS 0.066856f
C15783 VDD.t3104 VSS 0.066856f
C15784 VDD.t2266 VSS 0.066856f
C15785 VDD.n85 VSS 0.715442f
C15786 VDD.t2034 VSS 0.028519f
C15787 VDD.t2267 VSS 0.028519f
C15788 VDD.n86 VSS 0.009191f
C15789 VDD.t1614 VSS 0.028519f
C15790 VDD.t3105 VSS 0.028519f
C15791 VDD.n87 VSS 0.009191f
C15792 VDD.n88 VSS 0.263202f
C15793 VDD.n89 VSS 0.62638f
C15794 VDD.n90 VSS 0.099723f
C15795 VDD.t1997 VSS 0.066856f
C15796 VDD.n91 VSS 0.125227f
C15797 VDD.n92 VSS 0.101294f
C15798 VDD.n93 VSS 0.016021f
C15799 VDD.t2244 VSS 0.025104f
C15800 VDD.n94 VSS 0.081176f
C15801 VDD.n95 VSS 0.048151f
C15802 VDD.t639 VSS 1.45794f
C15803 VDD.t629 VSS 1.96535f
C15804 VDD.t1998 VSS 1.96535f
C15805 VDD.t2243 VSS 1.36988f
C15806 VDD.t1427 VSS 1.45794f
C15807 VDD.n96 VSS 0.208771f
C15808 VDD.n97 VSS 0.206947f
C15809 VDD.t2513 VSS 0.028519f
C15810 VDD.t2725 VSS 0.028519f
C15811 VDD.n98 VSS 0.009191f
C15812 VDD.t987 VSS 0.028519f
C15813 VDD.t1156 VSS 0.028519f
C15814 VDD.n99 VSS 0.009191f
C15815 VDD.n100 VSS 0.471397f
C15816 VDD.t1792 VSS 0.028519f
C15817 VDD.t2057 VSS 0.028519f
C15818 VDD.n101 VSS 0.009191f
C15819 VDD.t1791 VSS 0.066856f
C15820 VDD.t4490 VSS 0.066856f
C15821 VDD.t2223 VSS 0.066856f
C15822 VDD.t750 VSS 0.066856f
C15823 VDD.t2224 VSS 0.028519f
C15824 VDD.t2503 VSS 0.028519f
C15825 VDD.n102 VSS 0.009191f
C15826 VDD.t3794 VSS 0.066856f
C15827 VDD.t2410 VSS 0.066856f
C15828 VDD.t3795 VSS 0.028519f
C15829 VDD.t4017 VSS 0.028519f
C15830 VDD.n103 VSS 0.009191f
C15831 VDD.t3772 VSS 0.066856f
C15832 VDD.n104 VSS 0.125227f
C15833 VDD.t3997 VSS 0.025104f
C15834 VDD.t2524 VSS 0.066856f
C15835 VDD.n105 VSS 0.125227f
C15836 VDD.t906 VSS 0.025104f
C15837 VDD.n106 VSS 0.099723f
C15838 VDD.t2600 VSS 0.028519f
C15839 VDD.t971 VSS 0.028519f
C15840 VDD.n107 VSS 0.009191f
C15841 VDD.t1050 VSS 0.028519f
C15842 VDD.t1236 VSS 0.028519f
C15843 VDD.n108 VSS 0.009191f
C15844 VDD.n109 VSS 0.471397f
C15845 VDD.n110 VSS 0.207221f
C15846 VDD.n111 VSS 0.208771f
C15847 VDD.n112 VSS 0.206947f
C15848 VDD.t1655 VSS 1.96535f
C15849 VDD.t551 VSS 1.96535f
C15850 VDD.t550 VSS 1.36988f
C15851 VDD.n113 VSS 0.645798f
C15852 VDD.n114 VSS 0.595476f
C15853 VDD.t548 VSS 1.31955f
C15854 VDD.t549 VSS 1.96535f
C15855 VDD.t831 VSS 1.96535f
C15856 VDD.t623 VSS 1.45794f
C15857 VDD.n115 VSS 0.865258f
C15858 VDD.n116 VSS 0.902999f
C15859 VDD.t2015 VSS 0.028519f
C15860 VDD.t4587 VSS 0.028519f
C15861 VDD.n117 VSS 0.009191f
C15862 VDD.t2893 VSS 0.028519f
C15863 VDD.t3097 VSS 0.028519f
C15864 VDD.n118 VSS 0.009191f
C15865 VDD.n119 VSS 0.475536f
C15866 VDD.t1396 VSS 0.028519f
C15867 VDD.t4031 VSS 0.028519f
C15868 VDD.n120 VSS 0.009191f
C15869 VDD.t2239 VSS 0.028519f
C15870 VDD.t2517 VSS 0.028519f
C15871 VDD.n121 VSS 0.009191f
C15872 VDD.n122 VSS 0.528101f
C15873 VDD.n123 VSS 0.208771f
C15874 VDD.n124 VSS 0.207221f
C15875 VDD.t4630 VSS 0.066856f
C15876 VDD.n125 VSS 0.125227f
C15877 VDD.t4407 VSS 0.025104f
C15878 VDD.t1395 VSS 0.066856f
C15879 VDD.t2238 VSS 0.066856f
C15880 VDD.t2516 VSS 0.066856f
C15881 VDD.t4030 VSS 0.066856f
C15882 VDD.n126 VSS 0.696076f
C15883 VDD.t1765 VSS 0.066856f
C15884 VDD.t2673 VSS 0.066856f
C15885 VDD.t2880 VSS 0.066856f
C15886 VDD.t4376 VSS 0.066856f
C15887 VDD.n127 VSS 0.696076f
C15888 VDD.t1766 VSS 0.028519f
C15889 VDD.t4377 VSS 0.028519f
C15890 VDD.n128 VSS 0.009191f
C15891 VDD.t2674 VSS 0.028519f
C15892 VDD.t2881 VSS 0.028519f
C15893 VDD.n129 VSS 0.009191f
C15894 VDD.n130 VSS 0.650522f
C15895 VDD.t3393 VSS 0.066856f
C15896 VDD.t4196 VSS 0.066856f
C15897 VDD.t4382 VSS 0.066856f
C15898 VDD.t1788 VSS 0.066856f
C15899 VDD.n131 VSS 0.715442f
C15900 VDD.t3394 VSS 0.028519f
C15901 VDD.t1790 VSS 0.028519f
C15902 VDD.n132 VSS 0.009191f
C15903 VDD.t4197 VSS 0.028519f
C15904 VDD.t4383 VSS 0.028519f
C15905 VDD.n133 VSS 0.009191f
C15906 VDD.n134 VSS 0.263202f
C15907 VDD.n135 VSS 0.035132f
C15908 VDD.t4229 VSS 0.025104f
C15909 VDD.t4078 VSS 0.066856f
C15910 VDD.n136 VSS 0.125227f
C15911 VDD.t3859 VSS 0.025104f
C15912 VDD.t3858 VSS 0.066856f
C15913 VDD.n137 VSS 0.125227f
C15914 VDD.n138 VSS 0.101294f
C15915 VDD.n139 VSS 0.016021f
C15916 VDD.t4079 VSS 0.025104f
C15917 VDD.n140 VSS 0.081176f
C15918 VDD.n141 VSS 0.048151f
C15919 VDD.n142 VSS 0.083673f
C15920 VDD.t4228 VSS 0.066856f
C15921 VDD.n143 VSS 0.125227f
C15922 VDD.n144 VSS 0.006598f
C15923 VDD.n145 VSS 0.010188f
C15924 VDD.t4759 VSS 0.020387f
C15925 VDD.t4765 VSS 0.022137f
C15926 VDD.n146 VSS 0.069721f
C15927 VDD.n147 VSS 0.040089f
C15928 VDD.t4763 VSS 0.022115f
C15929 VDD.t4758 VSS 0.020371f
C15930 VDD.n148 VSS 0.027128f
C15931 VDD.n149 VSS 0.036577f
C15932 VDD.n150 VSS 0.044801f
C15933 VDD.n151 VSS 0.278297f
C15934 VDD.n152 VSS 0.040089f
C15935 VDD.t4761 VSS 0.020387f
C15936 VDD.n153 VSS 0.049653f
C15937 VDD.t4764 VSS 0.017093f
C15938 VDD.n154 VSS 0.042104f
C15939 VDD.n155 VSS 0.069461f
C15940 VDD.t4762 VSS 0.017093f
C15941 VDD.n156 VSS 0.035483f
C15942 VDD.t4760 VSS 0.020371f
C15943 VDD.n157 VSS 0.027128f
C15944 VDD.n158 VSS 0.016538f
C15945 VDD.n159 VSS 0.027213f
C15946 VDD.n160 VSS 0.204333f
C15947 VDD.n161 VSS 0.030906f
C15948 VDD.t2730 VSS 0.066856f
C15949 VDD.n162 VSS 0.045867f
C15950 VDD.n163 VSS 0.015693f
C15951 VDD.n164 VSS 0.010881f
C15952 VDD.n165 VSS 0.044227f
C15953 VDD.n166 VSS 0.094696f
C15954 VDD.n167 VSS 0.016021f
C15955 VDD.t2732 VSS 0.025104f
C15956 VDD.n168 VSS 0.08403f
C15957 VDD.n169 VSS 0.62638f
C15958 VDD.n170 VSS 0.099723f
C15959 VDD.t4406 VSS 0.066856f
C15960 VDD.n171 VSS 0.125227f
C15961 VDD.n172 VSS 0.101294f
C15962 VDD.n173 VSS 0.016021f
C15963 VDD.t4631 VSS 0.025104f
C15964 VDD.n174 VSS 0.081176f
C15965 VDD.n175 VSS 0.048151f
C15966 VDD.t1055 VSS 1.45794f
C15967 VDD.t1789 VSS 1.96535f
C15968 VDD.t2100 VSS 1.96535f
C15969 VDD.t2385 VSS 1.36988f
C15970 VDD.t1130 VSS 1.45794f
C15971 VDD.n176 VSS 0.208771f
C15972 VDD.n177 VSS 0.206947f
C15973 VDD.t2110 VSS 0.028519f
C15974 VDD.t1023 VSS 0.028519f
C15975 VDD.n178 VSS 0.009191f
C15976 VDD.t615 VSS 0.028519f
C15977 VDD.t3602 VSS 0.028519f
C15978 VDD.n179 VSS 0.009191f
C15979 VDD.n180 VSS 0.471397f
C15980 VDD.t1478 VSS 0.028519f
C15981 VDD.t4533 VSS 0.028519f
C15982 VDD.n181 VSS 0.009191f
C15983 VDD.t1477 VSS 0.066856f
C15984 VDD.t4216 VSS 0.066856f
C15985 VDD.t1860 VSS 0.066856f
C15986 VDD.t4534 VSS 0.066856f
C15987 VDD.t1861 VSS 0.028519f
C15988 VDD.t796 VSS 0.028519f
C15989 VDD.n182 VSS 0.009191f
C15990 VDD.t3486 VSS 0.066856f
C15991 VDD.t2004 VSS 0.066856f
C15992 VDD.t3487 VSS 0.028519f
C15993 VDD.t2457 VSS 0.028519f
C15994 VDD.n183 VSS 0.009191f
C15995 VDD.n184 VSS 0.099723f
C15996 VDD.t4604 VSS 0.066856f
C15997 VDD.n185 VSS 0.125227f
C15998 VDD.t2047 VSS 0.025104f
C15999 VDD.n186 VSS 0.083673f
C16000 VDD.t2045 VSS 0.066856f
C16001 VDD.n187 VSS 0.125227f
C16002 VDD.n188 VSS 0.101294f
C16003 VDD.n189 VSS 0.016021f
C16004 VDD.t4605 VSS 0.025104f
C16005 VDD.n190 VSS 0.099723f
C16006 VDD.n191 VSS 0.012131f
C16007 VDD.n192 VSS 0.012131f
C16008 VDD.n193 VSS 0.012131f
C16009 VDD.n194 VSS 0.012131f
C16010 VDD.n195 VSS 0.027719f
C16011 VDD.n196 VSS 0.012131f
C16012 VDD.n197 VSS 0.012131f
C16013 VDD.n198 VSS 0.012131f
C16014 VDD.n199 VSS 0.012131f
C16015 VDD.n200 VSS 0.012131f
C16016 VDD.n201 VSS 0.012131f
C16017 VDD.n202 VSS 0.012131f
C16018 VDD.n203 VSS 0.012131f
C16019 VDD.n204 VSS 0.012131f
C16020 VDD.n205 VSS 0.012131f
C16021 VDD.n206 VSS 0.012131f
C16022 VDD.n207 VSS 0.012131f
C16023 VDD.n208 VSS 0.012131f
C16024 VDD.n209 VSS 0.012131f
C16025 VDD.n210 VSS 0.012131f
C16026 VDD.n211 VSS 0.012131f
C16027 VDD.n212 VSS 0.012131f
C16028 VDD.n213 VSS 0.012131f
C16029 VDD.n214 VSS 0.012131f
C16030 VDD.n215 VSS 0.012131f
C16031 VDD.n216 VSS 0.012131f
C16032 VDD.n217 VSS 0.012131f
C16033 VDD.n218 VSS 0.012131f
C16034 VDD.n219 VSS 0.012131f
C16035 VDD.n220 VSS 0.012131f
C16036 VDD.n221 VSS 0.012131f
C16037 VDD.n222 VSS 0.012131f
C16038 VDD.n223 VSS 0.012131f
C16039 VDD.n224 VSS 0.012131f
C16040 VDD.n225 VSS 0.012131f
C16041 VDD.n226 VSS 0.012131f
C16042 VDD.n227 VSS 0.012131f
C16043 VDD.n228 VSS 0.012131f
C16044 VDD.n229 VSS 0.012131f
C16045 VDD.n230 VSS 0.012131f
C16046 VDD.n231 VSS 0.012131f
C16047 VDD.n232 VSS 0.012131f
C16048 VDD.n233 VSS 0.012131f
C16049 VDD.n234 VSS 0.012131f
C16050 VDD.n235 VSS 0.012131f
C16051 VDD.n236 VSS 0.012131f
C16052 VDD.n237 VSS 0.012131f
C16053 VDD.n238 VSS 0.012131f
C16054 VDD.n239 VSS 0.012131f
C16055 VDD.n240 VSS 0.012131f
C16056 VDD.n241 VSS 0.012131f
C16057 VDD.n242 VSS 0.012131f
C16058 VDD.n243 VSS 0.012131f
C16059 VDD.n244 VSS 0.012131f
C16060 VDD.n245 VSS 0.012131f
C16061 VDD.n246 VSS 0.012131f
C16062 VDD.n247 VSS 0.012131f
C16063 VDD.n248 VSS 0.012131f
C16064 VDD.n249 VSS 0.012131f
C16065 VDD.n250 VSS 0.012131f
C16066 VDD.n251 VSS 0.012131f
C16067 VDD.n252 VSS 0.012131f
C16068 VDD.n253 VSS 0.012131f
C16069 VDD.n254 VSS 0.012131f
C16070 VDD.n255 VSS 0.012131f
C16071 VDD.n256 VSS 0.012131f
C16072 VDD.n257 VSS 0.012131f
C16073 VDD.n258 VSS 0.012131f
C16074 VDD.n259 VSS 0.012131f
C16075 VDD.n260 VSS 0.012131f
C16076 VDD.n261 VSS 0.012131f
C16077 VDD.n262 VSS 0.012131f
C16078 VDD.n263 VSS 0.012131f
C16079 VDD.n264 VSS 0.012131f
C16080 VDD.n265 VSS 0.012131f
C16081 VDD.n266 VSS 0.012131f
C16082 VDD.n267 VSS 0.012131f
C16083 VDD.n268 VSS 0.012131f
C16084 VDD.n269 VSS 0.012131f
C16085 VDD.n270 VSS 0.012131f
C16086 VDD.n271 VSS 0.012131f
C16087 VDD.n272 VSS 0.012131f
C16088 VDD.n273 VSS 0.012131f
C16089 VDD.n274 VSS 0.012131f
C16090 VDD.n275 VSS 0.012131f
C16091 VDD.n276 VSS 0.012131f
C16092 VDD.n277 VSS 0.012131f
C16093 VDD.n278 VSS 0.012131f
C16094 VDD.n279 VSS 0.012131f
C16095 VDD.n280 VSS 0.012131f
C16096 VDD.n281 VSS 0.012131f
C16097 VDD.n282 VSS 0.012131f
C16098 VDD.n283 VSS 0.012131f
C16099 VDD.n284 VSS 0.012131f
C16100 VDD.n285 VSS 0.012131f
C16101 VDD.n286 VSS 0.012131f
C16102 VDD.n287 VSS 0.012131f
C16103 VDD.n288 VSS 0.012131f
C16104 VDD.n289 VSS 0.012131f
C16105 VDD.n290 VSS 0.012131f
C16106 VDD.n291 VSS 0.012131f
C16107 VDD.n292 VSS 0.012131f
C16108 VDD.n293 VSS 0.012131f
C16109 VDD.n294 VSS 0.012131f
C16110 VDD.n295 VSS 0.012131f
C16111 VDD.n296 VSS 0.012131f
C16112 VDD.n297 VSS 0.012131f
C16113 VDD.n298 VSS 0.012131f
C16114 VDD.n299 VSS 0.012131f
C16115 VDD.n300 VSS 0.012131f
C16116 VDD.n301 VSS 0.012131f
C16117 VDD.n302 VSS 0.012131f
C16118 VDD.n303 VSS 0.012131f
C16119 VDD.n304 VSS 0.012131f
C16120 VDD.n305 VSS 0.012131f
C16121 VDD.n306 VSS 0.012131f
C16122 VDD.n307 VSS 0.012131f
C16123 VDD.n308 VSS 0.012131f
C16124 VDD.n309 VSS 0.012131f
C16125 VDD.n310 VSS 0.012131f
C16126 VDD.n311 VSS 0.012131f
C16127 VDD.n312 VSS 0.012131f
C16128 VDD.n313 VSS 0.012131f
C16129 VDD.n314 VSS 0.012131f
C16130 VDD.n315 VSS 0.012131f
C16131 VDD.n316 VSS 0.012131f
C16132 VDD.n317 VSS 0.012131f
C16133 VDD.n318 VSS 0.012131f
C16134 VDD.n319 VSS 0.012131f
C16135 VDD.n320 VSS 0.012131f
C16136 VDD.n321 VSS 0.012131f
C16137 VDD.n322 VSS 0.012131f
C16138 VDD.n323 VSS 0.012131f
C16139 VDD.n324 VSS 0.012131f
C16140 VDD.n325 VSS 0.012131f
C16141 VDD.n326 VSS 0.012131f
C16142 VDD.n327 VSS 0.012131f
C16143 VDD.n328 VSS 0.012131f
C16144 VDD.n329 VSS 0.012131f
C16145 VDD.n330 VSS 0.012131f
C16146 VDD.n331 VSS 0.012131f
C16147 VDD.n332 VSS 0.012131f
C16148 VDD.n333 VSS 0.012131f
C16149 VDD.n334 VSS 0.012131f
C16150 VDD.n335 VSS 0.012131f
C16151 VDD.n336 VSS 0.012131f
C16152 VDD.n337 VSS 0.012131f
C16153 VDD.n338 VSS 0.012131f
C16154 VDD.n339 VSS 0.012131f
C16155 VDD.n340 VSS 0.012131f
C16156 VDD.n341 VSS 0.012131f
C16157 VDD.n342 VSS 0.012131f
C16158 VDD.n343 VSS 0.012131f
C16159 VDD.n344 VSS 0.012131f
C16160 VDD.n345 VSS 0.012131f
C16161 VDD.n346 VSS 0.012131f
C16162 VDD.n347 VSS 0.012131f
C16163 VDD.n348 VSS 0.012131f
C16164 VDD.n349 VSS 0.012131f
C16165 VDD.n350 VSS 0.012131f
C16166 VDD.n351 VSS 0.012131f
C16167 VDD.n352 VSS 0.012131f
C16168 VDD.n353 VSS 0.012131f
C16169 VDD.n354 VSS 0.012131f
C16170 VDD.n355 VSS 0.012131f
C16171 VDD.n356 VSS 0.012131f
C16172 VDD.n357 VSS 0.012131f
C16173 VDD.n358 VSS 0.012131f
C16174 VDD.n359 VSS 0.012131f
C16175 VDD.n360 VSS 0.012131f
C16176 VDD.n361 VSS 0.012131f
C16177 VDD.n362 VSS 0.012131f
C16178 VDD.n363 VSS 0.012131f
C16179 VDD.n364 VSS 0.012131f
C16180 VDD.n365 VSS 0.012131f
C16181 VDD.n366 VSS 0.012131f
C16182 VDD.n367 VSS 0.012131f
C16183 VDD.n368 VSS 0.012131f
C16184 VDD.n369 VSS 0.012131f
C16185 VDD.n370 VSS 0.012131f
C16186 VDD.n371 VSS 0.012131f
C16187 VDD.n372 VSS 0.012131f
C16188 VDD.n373 VSS 0.012131f
C16189 VDD.n374 VSS 0.012131f
C16190 VDD.n375 VSS 0.012131f
C16191 VDD.n376 VSS 0.012131f
C16192 VDD.n377 VSS 0.012131f
C16193 VDD.n378 VSS 0.012131f
C16194 VDD.n379 VSS 0.012131f
C16195 VDD.n380 VSS 0.012131f
C16196 VDD.n381 VSS 0.012131f
C16197 VDD.n382 VSS 0.012131f
C16198 VDD.n383 VSS 0.012131f
C16199 VDD.n384 VSS 0.007954f
C16200 VDD.n385 VSS 0.012131f
C16201 VDD.n386 VSS 0.012131f
C16202 VDD.n387 VSS 0.012131f
C16203 VDD.n388 VSS 0.012131f
C16204 VDD.n389 VSS 0.012131f
C16205 VDD.n390 VSS 0.012131f
C16206 VDD.n391 VSS 0.012131f
C16207 VDD.n392 VSS 0.012131f
C16208 VDD.n393 VSS 0.012131f
C16209 VDD.n394 VSS 0.012131f
C16210 VDD.n395 VSS 0.012131f
C16211 VDD.n396 VSS 0.012131f
C16212 VDD.n397 VSS 0.012131f
C16213 VDD.n398 VSS 0.012131f
C16214 VDD.n399 VSS 0.012131f
C16215 VDD.n400 VSS 0.012131f
C16216 VDD.n401 VSS 0.012131f
C16217 VDD.n402 VSS 0.012131f
C16218 VDD.n403 VSS 0.012131f
C16219 VDD.n404 VSS 0.012131f
C16220 VDD.n405 VSS 0.032438f
C16221 VDD.n406 VSS 0.012131f
C16222 VDD.n407 VSS 0.012131f
C16223 VDD.n408 VSS 0.012131f
C16224 VDD.n409 VSS 0.012131f
C16225 VDD.n410 VSS 0.012131f
C16226 VDD.n411 VSS 0.012131f
C16227 VDD.n412 VSS 0.012131f
C16228 VDD.n413 VSS 0.012131f
C16229 VDD.n414 VSS 0.012131f
C16230 VDD.n415 VSS 0.012131f
C16231 VDD.n416 VSS 0.012131f
C16232 VDD.n417 VSS 0.012131f
C16233 VDD.n418 VSS 0.012131f
C16234 VDD.n419 VSS 0.012131f
C16235 VDD.n420 VSS 0.012131f
C16236 VDD.n421 VSS 0.012131f
C16237 VDD.n422 VSS 0.012131f
C16238 VDD.n423 VSS 0.012131f
C16239 VDD.n424 VSS 0.012131f
C16240 VDD.n425 VSS 0.012131f
C16241 VDD.n426 VSS 0.012131f
C16242 VDD.n427 VSS 0.012131f
C16243 VDD.n428 VSS 0.012131f
C16244 VDD.n429 VSS 0.012131f
C16245 VDD.n430 VSS 0.012131f
C16246 VDD.n431 VSS 0.012131f
C16247 VDD.n432 VSS 0.012131f
C16248 VDD.n433 VSS 0.012131f
C16249 VDD.n434 VSS 0.012131f
C16250 VDD.n435 VSS 0.012131f
C16251 VDD.n436 VSS 0.012131f
C16252 VDD.n437 VSS 0.012131f
C16253 VDD.n438 VSS 0.012131f
C16254 VDD.n439 VSS 0.012131f
C16255 VDD.n440 VSS 0.012131f
C16256 VDD.n441 VSS 0.012131f
C16257 VDD.n442 VSS 0.012131f
C16258 VDD.n443 VSS 0.012131f
C16259 VDD.n444 VSS 0.012131f
C16260 VDD.n445 VSS 0.012131f
C16261 VDD.n446 VSS 0.012131f
C16262 VDD.n447 VSS 0.012131f
C16263 VDD.n448 VSS 0.012131f
C16264 VDD.n449 VSS 0.012131f
C16265 VDD.n450 VSS 0.012131f
C16266 VDD.n451 VSS 0.012131f
C16267 VDD.n452 VSS 0.012131f
C16268 VDD.n453 VSS 0.012131f
C16269 VDD.n454 VSS 0.012131f
C16270 VDD.n455 VSS 0.012131f
C16271 VDD.n456 VSS 0.012131f
C16272 VDD.n457 VSS 0.012131f
C16273 VDD.n458 VSS 0.012131f
C16274 VDD.n459 VSS 0.012131f
C16275 VDD.n460 VSS 0.012131f
C16276 VDD.n461 VSS 0.012131f
C16277 VDD.n462 VSS 0.012131f
C16278 VDD.n463 VSS 0.012131f
C16279 VDD.n464 VSS 0.012131f
C16280 VDD.n465 VSS 0.012131f
C16281 VDD.n466 VSS 0.012131f
C16282 VDD.n467 VSS 0.012131f
C16283 VDD.n468 VSS 0.012131f
C16284 VDD.n469 VSS 0.012131f
C16285 VDD.n470 VSS 0.012131f
C16286 VDD.n471 VSS 0.012131f
C16287 VDD.n472 VSS 0.012131f
C16288 VDD.n473 VSS 0.012131f
C16289 VDD.n474 VSS 0.012131f
C16290 VDD.n475 VSS 0.012131f
C16291 VDD.n476 VSS 0.012131f
C16292 VDD.n477 VSS 0.012131f
C16293 VDD.n478 VSS 0.012131f
C16294 VDD.n479 VSS 0.012131f
C16295 VDD.n480 VSS 0.012131f
C16296 VDD.n481 VSS 0.012131f
C16297 VDD.n482 VSS 0.012131f
C16298 VDD.n483 VSS 0.012131f
C16299 VDD.n484 VSS 0.012131f
C16300 VDD.n485 VSS 0.012131f
C16301 VDD.n486 VSS 0.012131f
C16302 VDD.n487 VSS 0.012131f
C16303 VDD.n488 VSS 0.012131f
C16304 VDD.n489 VSS 0.012131f
C16305 VDD.n490 VSS 0.012131f
C16306 VDD.n491 VSS 0.012131f
C16307 VDD.n492 VSS 0.012131f
C16308 VDD.n493 VSS 0.012131f
C16309 VDD.n494 VSS 0.012131f
C16310 VDD.n495 VSS 0.012131f
C16311 VDD.n496 VSS 0.012131f
C16312 VDD.n497 VSS 0.012131f
C16313 VDD.n498 VSS 0.012131f
C16314 VDD.n499 VSS 0.012131f
C16315 VDD.n500 VSS 0.012131f
C16316 VDD.n501 VSS 0.012131f
C16317 VDD.n502 VSS 0.012131f
C16318 VDD.n503 VSS 0.012131f
C16319 VDD.n504 VSS 0.012131f
C16320 VDD.n505 VSS 0.012131f
C16321 VDD.n506 VSS 0.012131f
C16322 VDD.n507 VSS 0.012131f
C16323 VDD.n508 VSS 0.012131f
C16324 VDD.n509 VSS 0.012131f
C16325 VDD.n510 VSS 0.012131f
C16326 VDD.n511 VSS 0.012131f
C16327 VDD.n512 VSS 0.012131f
C16328 VDD.n513 VSS 0.012131f
C16329 VDD.n514 VSS 0.012131f
C16330 VDD.n515 VSS 0.012131f
C16331 VDD.n516 VSS 0.012131f
C16332 VDD.n517 VSS 0.012131f
C16333 VDD.n518 VSS 0.012131f
C16334 VDD.n519 VSS 0.012131f
C16335 VDD.n520 VSS 0.012131f
C16336 VDD.n521 VSS 0.012131f
C16337 VDD.n522 VSS 0.012131f
C16338 VDD.n523 VSS 0.012131f
C16339 VDD.n524 VSS 0.012131f
C16340 VDD.n525 VSS 0.012131f
C16341 VDD.n526 VSS 0.012131f
C16342 VDD.n527 VSS 0.012131f
C16343 VDD.n528 VSS 0.012131f
C16344 VDD.n529 VSS 0.012131f
C16345 VDD.n530 VSS 0.012131f
C16346 VDD.n531 VSS 0.012131f
C16347 VDD.n532 VSS 0.012131f
C16348 VDD.n533 VSS 0.012131f
C16349 VDD.n534 VSS 0.012131f
C16350 VDD.n535 VSS 0.012131f
C16351 VDD.n536 VSS 0.012131f
C16352 VDD.n537 VSS 0.012131f
C16353 VDD.n538 VSS 0.012131f
C16354 VDD.n539 VSS 0.012131f
C16355 VDD.n540 VSS 0.012131f
C16356 VDD.n541 VSS 0.012131f
C16357 VDD.n542 VSS 0.012131f
C16358 VDD.n543 VSS 0.012131f
C16359 VDD.n544 VSS 0.012131f
C16360 VDD.n545 VSS 0.012131f
C16361 VDD.n546 VSS 0.012131f
C16362 VDD.n547 VSS 0.012131f
C16363 VDD.n548 VSS 0.012131f
C16364 VDD.n549 VSS 0.012131f
C16365 VDD.n550 VSS 0.012131f
C16366 VDD.n551 VSS 0.012131f
C16367 VDD.n552 VSS 0.012131f
C16368 VDD.n553 VSS 0.012131f
C16369 VDD.n554 VSS 0.012131f
C16370 VDD.n555 VSS 0.012131f
C16371 VDD.n556 VSS 0.012131f
C16372 VDD.n557 VSS 0.012131f
C16373 VDD.n558 VSS 0.012131f
C16374 VDD.n559 VSS 0.012131f
C16375 VDD.n560 VSS 0.012131f
C16376 VDD.n561 VSS 0.012131f
C16377 VDD.n562 VSS 0.012131f
C16378 VDD.n563 VSS 0.012131f
C16379 VDD.n564 VSS 0.012131f
C16380 VDD.n565 VSS 0.012131f
C16381 VDD.n566 VSS 0.012131f
C16382 VDD.n567 VSS 0.012131f
C16383 VDD.n568 VSS 0.012131f
C16384 VDD.n569 VSS 0.012131f
C16385 VDD.n570 VSS 0.012131f
C16386 VDD.n571 VSS 0.012131f
C16387 VDD.n572 VSS 0.012131f
C16388 VDD.n573 VSS 0.012131f
C16389 VDD.n574 VSS 0.012131f
C16390 VDD.n575 VSS 0.012131f
C16391 VDD.n576 VSS 0.012131f
C16392 VDD.n577 VSS 0.012131f
C16393 VDD.n578 VSS 0.012131f
C16394 VDD.n579 VSS 0.012131f
C16395 VDD.n580 VSS 0.012131f
C16396 VDD.n581 VSS 0.012131f
C16397 VDD.n582 VSS 0.012131f
C16398 VDD.n583 VSS 0.012131f
C16399 VDD.n584 VSS 0.012131f
C16400 VDD.n585 VSS 0.012131f
C16401 VDD.n586 VSS 0.012131f
C16402 VDD.n587 VSS 0.012131f
C16403 VDD.n588 VSS 0.012131f
C16404 VDD.n589 VSS 0.012131f
C16405 VDD.n590 VSS 0.012131f
C16406 VDD.n591 VSS 0.012131f
C16407 VDD.n592 VSS 0.012131f
C16408 VDD.n593 VSS 0.012131f
C16409 VDD.n594 VSS 0.012131f
C16410 VDD.n595 VSS 0.012131f
C16411 VDD.n596 VSS 0.012131f
C16412 VDD.n597 VSS 0.012131f
C16413 VDD.n598 VSS 0.012131f
C16414 VDD.n599 VSS 0.012131f
C16415 VDD.n600 VSS 0.012131f
C16416 VDD.n601 VSS 0.012131f
C16417 VDD.n602 VSS 0.012131f
C16418 VDD.n603 VSS 0.012131f
C16419 VDD.n604 VSS 0.012131f
C16420 VDD.n605 VSS 0.012131f
C16421 VDD.n606 VSS 0.012131f
C16422 VDD.n607 VSS 0.012131f
C16423 VDD.n608 VSS 0.012131f
C16424 VDD.n609 VSS 0.012131f
C16425 VDD.n610 VSS 0.012131f
C16426 VDD.n611 VSS 0.012131f
C16427 VDD.n612 VSS 0.012131f
C16428 VDD.n613 VSS 0.012131f
C16429 VDD.n614 VSS 0.012131f
C16430 VDD.n615 VSS 0.012131f
C16431 VDD.n616 VSS 0.012131f
C16432 VDD.n617 VSS 0.012131f
C16433 VDD.n618 VSS 0.012131f
C16434 VDD.n619 VSS 0.012131f
C16435 VDD.n620 VSS 0.012131f
C16436 VDD.n621 VSS 0.012131f
C16437 VDD.n622 VSS 0.012131f
C16438 VDD.n623 VSS 0.012131f
C16439 VDD.n624 VSS 0.012131f
C16440 VDD.n625 VSS 0.012131f
C16441 VDD.n626 VSS 0.012131f
C16442 VDD.n627 VSS 0.012131f
C16443 VDD.n628 VSS 0.012131f
C16444 VDD.n629 VSS 0.012131f
C16445 VDD.n630 VSS 0.012131f
C16446 VDD.n631 VSS 0.269046f
C16447 VDD.n632 VSS 0.012131f
C16448 VDD.n633 VSS 0.031727f
C16449 VDD.n634 VSS 0.009688f
C16450 VDD.n635 VSS 0.01502f
C16451 VDD.n636 VSS 0.01487f
C16452 VDD.n637 VSS 0.018625f
C16453 VDD.n638 VSS 0.009312f
C16454 VDD.n640 VSS 0.134523f
C16455 VDD.t3943 VSS 0.028519f
C16456 VDD.t2044 VSS 0.028519f
C16457 VDD.n641 VSS 0.009191f
C16458 VDD.n642 VSS 0.147389f
C16459 VDD.n644 VSS 0.183585f
C16460 VDD.n645 VSS 0.012131f
C16461 VDD.n646 VSS 0.269046f
C16462 VDD.n647 VSS 0.012131f
C16463 VDD.t969 VSS 0.028519f
C16464 VDD.t2394 VSS 0.028519f
C16465 VDD.n648 VSS 0.009191f
C16466 VDD.n649 VSS 0.149927f
C16467 VDD.n650 VSS 0.012131f
C16468 VDD.t967 VSS 0.066856f
C16469 VDD.t2393 VSS 0.066856f
C16470 VDD.n651 VSS 0.182387f
C16471 VDD.n652 VSS 0.012131f
C16472 VDD.n653 VSS 0.269046f
C16473 VDD.n654 VSS 0.012131f
C16474 VDD.n655 VSS 0.227166f
C16475 VDD.n656 VSS 0.012131f
C16476 VDD.n657 VSS 0.134523f
C16477 VDD.n658 VSS 0.012131f
C16478 VDD.n659 VSS 0.257624f
C16479 VDD.n660 VSS 0.012131f
C16480 VDD.t3882 VSS 0.066856f
C16481 VDD.t1101 VSS 0.066856f
C16482 VDD.n661 VSS 0.182387f
C16483 VDD.n662 VSS 0.012131f
C16484 VDD.n663 VSS 0.269046f
C16485 VDD.n664 VSS 0.012131f
C16486 VDD.n665 VSS 0.257624f
C16487 VDD.n666 VSS 0.012131f
C16488 VDD.n667 VSS 0.269046f
C16489 VDD.n668 VSS 0.012131f
C16490 VDD.t1671 VSS 0.066856f
C16491 VDD.t3126 VSS 0.066856f
C16492 VDD.n669 VSS 0.115126f
C16493 VDD.n673 VSS 0.139599f
C16494 VDD.n674 VSS 0.018249f
C16495 VDD.n675 VSS 0.018625f
C16496 VDD.n676 VSS 0.131985f
C16497 VDD.n677 VSS 0.009688f
C16498 VDD.n678 VSS 0.104438f
C16499 VDD.t1172 VSS 0.034186f
C16500 VDD.n679 VSS 0.095183f
C16501 VDD.n680 VSS 0.089932f
C16502 VDD.n682 VSS 0.549746f
C16503 VDD.t3050 VSS 0.080309f
C16504 VDD.n683 VSS 0.17245f
C16505 VDD.t740 VSS 0.080309f
C16506 VDD.n684 VSS 0.17245f
C16507 VDD.t4641 VSS 0.016021f
C16508 VDD.n685 VSS 0.121516f
C16509 VDD.n686 VSS 0.304439f
C16510 VDD.n687 VSS 0.303418f
C16511 VDD.t431 VSS 3.20156f
C16512 VDD.n688 VSS 0.304763f
C16513 VDD.n689 VSS 0.304763f
C16514 VDD.t422 VSS 7.65735f
C16515 VDD.t426 VSS 7.734359f
C16516 VDD.t471 VSS 9.533179f
C16517 VDD.t686 VSS 7.54183f
C16518 VDD.n690 VSS 3.54262f
C16519 VDD.n691 VSS 0.304439f
C16520 VDD.n692 VSS 0.303418f
C16521 VDD.t1106 VSS 0.080309f
C16522 VDD.t1290 VSS 0.080309f
C16523 VDD.n693 VSS 0.24784f
C16524 VDD.n694 VSS 0.016021f
C16525 VDD.t1288 VSS 0.080309f
C16526 VDD.t1505 VSS 0.080309f
C16527 VDD.n695 VSS 0.385661f
C16528 VDD.t1291 VSS 0.016021f
C16529 VDD.t1289 VSS 0.025104f
C16530 VDD.t1154 VSS 0.034186f
C16531 VDD.t486 VSS 0.092978f
C16532 VDD.n696 VSS 0.255649f
C16533 VDD.t1153 VSS 0.080309f
C16534 VDD.t1370 VSS 0.080309f
C16535 VDD.n697 VSS 0.342138f
C16536 VDD.t1575 VSS 0.034186f
C16537 VDD.t1574 VSS 0.080309f
C16538 VDD.t1784 VSS 0.080309f
C16539 VDD.n698 VSS 0.385661f
C16540 VDD.n699 VSS 0.332862f
C16541 VDD.n700 VSS 0.29513f
C16542 VDD.t3537 VSS 0.034186f
C16543 VDD.t3245 VSS 0.034186f
C16544 VDD.n701 VSS 0.278056f
C16545 VDD.t3244 VSS 0.080308f
C16546 VDD.t4637 VSS 0.034186f
C16547 VDD.t4295 VSS 0.034186f
C16548 VDD.n702 VSS 0.278056f
C16549 VDD.t4294 VSS 0.080308f
C16550 VDD.t4503 VSS 0.034186f
C16551 VDD.t4193 VSS 0.034186f
C16552 VDD.n703 VSS 0.278056f
C16553 VDD.t4192 VSS 0.080308f
C16554 VDD.t1460 VSS 0.034186f
C16555 VDD.t1133 VSS 0.034186f
C16556 VDD.n704 VSS 0.278056f
C16557 VDD.t1132 VSS 0.080308f
C16558 VDD.t1143 VSS 0.034186f
C16559 VDD.t819 VSS 0.034186f
C16560 VDD.n705 VSS 0.278056f
C16561 VDD.t818 VSS 0.080308f
C16562 VDD.n706 VSS 0.096875f
C16563 VDD.n707 VSS 0.304944f
C16564 VDD.n708 VSS 0.304763f
C16565 VDD.t469 VSS 9.533179f
C16566 VDD.t745 VSS 7.54183f
C16567 VDD.n709 VSS 3.4106f
C16568 VDD.n710 VSS 0.304439f
C16569 VDD.n711 VSS 0.304763f
C16570 VDD.t428 VSS 7.65735f
C16571 VDD.n712 VSS 0.303418f
C16572 VDD.t2720 VSS 0.080309f
C16573 VDD.t2944 VSS 0.080309f
C16574 VDD.n713 VSS 0.24784f
C16575 VDD.n714 VSS 0.016021f
C16576 VDD.t2940 VSS 0.080309f
C16577 VDD.t3136 VSS 0.080309f
C16578 VDD.n715 VSS 0.385661f
C16579 VDD.t2723 VSS 0.025104f
C16580 VDD.t2508 VSS 0.080309f
C16581 VDD.t2722 VSS 0.080309f
C16582 VDD.n716 VSS 0.385661f
C16583 VDD.t4068 VSS 0.080309f
C16584 VDD.t4286 VSS 0.080309f
C16585 VDD.n717 VSS 0.385661f
C16586 VDD.t4069 VSS 0.034186f
C16587 VDD.t2251 VSS 0.080309f
C16588 VDD.t2536 VSS 0.080309f
C16589 VDD.n718 VSS 0.385661f
C16590 VDD.t2252 VSS 0.034186f
C16591 VDD.t2537 VSS 0.034186f
C16592 VDD.n719 VSS 0.327288f
C16593 VDD.n720 VSS 0.327288f
C16594 VDD.t4287 VSS 0.034186f
C16595 VDD.n721 VSS 0.298193f
C16596 VDD.n722 VSS 0.298193f
C16597 VDD.t2509 VSS 0.025104f
C16598 VDD.t2721 VSS 0.016021f
C16599 VDD.n723 VSS 0.016021f
C16600 VDD.n724 VSS 0.289935f
C16601 VDD.n725 VSS 0.016021f
C16602 VDD.t2945 VSS 0.016021f
C16603 VDD.t2941 VSS 0.025104f
C16604 VDD.t2701 VSS 0.034186f
C16605 VDD.t2700 VSS 0.080309f
C16606 VDD.t2912 VSS 0.080309f
C16607 VDD.n726 VSS 0.385661f
C16608 VDD.t3107 VSS 0.034186f
C16609 VDD.t3106 VSS 0.080309f
C16610 VDD.t3296 VSS 0.080309f
C16611 VDD.n727 VSS 0.385661f
C16612 VDD.n728 VSS 0.332862f
C16613 VDD.n729 VSS 0.29513f
C16614 VDD.t1475 VSS 0.080308f
C16615 VDD.t481 VSS 0.017997f
C16616 VDD.t2149 VSS 0.034186f
C16617 VDD.t1476 VSS 0.034186f
C16618 VDD.n730 VSS 0.328513f
C16619 VDD.t4514 VSS 0.080308f
C16620 VDD.t474 VSS 0.017997f
C16621 VDD.t1029 VSS 0.034186f
C16622 VDD.t4515 VSS 0.034186f
C16623 VDD.n731 VSS 0.328513f
C16624 VDD.t712 VSS 0.080308f
C16625 VDD.t1323 VSS 0.034186f
C16626 VDD.t713 VSS 0.034186f
C16627 VDD.n732 VSS 0.278056f
C16628 VDD.t4736 VSS 0.080308f
C16629 VDD.t1215 VSS 0.034186f
C16630 VDD.t4737 VSS 0.034186f
C16631 VDD.n733 VSS 0.278056f
C16632 VDD.t714 VSS 0.080308f
C16633 VDD.t1328 VSS 0.034186f
C16634 VDD.t715 VSS 0.034186f
C16635 VDD.n734 VSS 0.278056f
C16636 VDD.t465 VSS 0.030249f
C16637 VDD.n735 VSS 0.077873f
C16638 VDD.n736 VSS 0.064716f
C16639 VDD.t456 VSS 0.008011f
C16640 VDD.t436 VSS 0.008011f
C16641 VDD.n737 VSS 0.030367f
C16642 VDD.n738 VSS 0.063471f
C16643 VDD.n739 VSS 0.063471f
C16644 VDD.t353 VSS 0.008011f
C16645 VDD.t346 VSS 0.008011f
C16646 VDD.n740 VSS 0.030367f
C16647 VDD.n741 VSS 0.064716f
C16648 VDD.n742 VSS 0.234959f
C16649 VDD.t336 VSS 0.008011f
C16650 VDD.t341 VSS 0.008011f
C16651 VDD.n743 VSS 0.030367f
C16652 VDD.n744 VSS 0.064716f
C16653 VDD.n745 VSS 0.234959f
C16654 VDD.t342 VSS 0.008011f
C16655 VDD.t356 VSS 0.008011f
C16656 VDD.n746 VSS 0.030367f
C16657 VDD.n747 VSS 0.031651f
C16658 VDD.t4621 VSS 0.034186f
C16659 VDD.n748 VSS 0.136328f
C16660 VDD.t4745 VSS 0.034186f
C16661 VDD.n749 VSS 0.136328f
C16662 VDD.t3633 VSS 0.034186f
C16663 VDD.n750 VSS 0.136328f
C16664 VDD.t386 VSS 0.019806f
C16665 VDD.t1522 VSS 0.035116f
C16666 VDD.n751 VSS 0.087326f
C16667 VDD.n752 VSS 0.15353f
C16668 VDD.t4553 VSS 0.034186f
C16669 VDD.n753 VSS 0.136328f
C16670 VDD.t3118 VSS 0.080309f
C16671 VDD.n754 VSS 0.132968f
C16672 VDD.t2710 VSS 0.080309f
C16673 VDD.n755 VSS 0.17245f
C16674 VDD.t1091 VSS 0.080309f
C16675 VDD.n756 VSS 0.17245f
C16676 VDD.t2746 VSS 0.016021f
C16677 VDD.t2745 VSS 0.080309f
C16678 VDD.n757 VSS 0.113227f
C16679 VDD.n758 VSS 0.304439f
C16680 VDD.n759 VSS 0.303418f
C16681 VDD.t314 VSS 3.20156f
C16682 VDD.n760 VSS 0.304944f
C16683 VDD.t321 VSS 7.65735f
C16684 VDD.n761 VSS 0.304763f
C16685 VDD.n762 VSS 0.304439f
C16686 VDD.t306 VSS 9.533179f
C16687 VDD.t578 VSS 7.54183f
C16688 VDD.n763 VSS 3.58663f
C16689 VDD.n764 VSS 0.303418f
C16690 VDD.t3542 VSS 0.080309f
C16691 VDD.n765 VSS 0.113227f
C16692 VDD.t3342 VSS 0.080309f
C16693 VDD.n766 VSS 0.17245f
C16694 VDD.t3543 VSS 0.016021f
C16695 VDD.t2139 VSS 0.080309f
C16696 VDD.n767 VSS 0.17245f
C16697 VDD.t2936 VSS 0.080309f
C16698 VDD.n768 VSS 0.132968f
C16699 VDD.t3410 VSS 0.034186f
C16700 VDD.n769 VSS 0.371358f
C16701 VDD.n770 VSS 0.32759f
C16702 VDD.n771 VSS 0.238069f
C16703 VDD.t4523 VSS 0.034186f
C16704 VDD.t4522 VSS 0.231787f
C16705 VDD.n772 VSS 0.32759f
C16706 VDD.t2326 VSS 0.034186f
C16707 VDD.n773 VSS 0.393929f
C16708 VDD.n774 VSS 0.275158f
C16709 VDD.t4589 VSS 0.034186f
C16710 VDD.n775 VSS 0.26663f
C16711 VDD.t2484 VSS 0.034186f
C16712 VDD.n776 VSS 0.26663f
C16713 VDD.n777 VSS 0.242279f
C16714 VDD.t1259 VSS 0.034186f
C16715 VDD.n778 VSS 0.26663f
C16716 VDD.n779 VSS 0.275158f
C16717 VDD.t924 VSS 0.034186f
C16718 VDD.n780 VSS 0.26663f
C16719 VDD.t1390 VSS 0.034186f
C16720 VDD.n781 VSS 0.26663f
C16721 VDD.n782 VSS 0.20535f
C16722 VDD.n783 VSS 0.064716f
C16723 VDD.t350 VSS 0.030249f
C16724 VDD.n784 VSS 0.077873f
C16725 VDD.t4476 VSS 0.080308f
C16726 VDD.t1698 VSS 0.034186f
C16727 VDD.t4477 VSS 0.034186f
C16728 VDD.n785 VSS 0.278056f
C16729 VDD.t656 VSS 0.080308f
C16730 VDD.t2073 VSS 0.034186f
C16731 VDD.t658 VSS 0.034186f
C16732 VDD.n786 VSS 0.278056f
C16733 VDD.t3699 VSS 0.080308f
C16734 VDD.t961 VSS 0.034186f
C16735 VDD.t3700 VSS 0.034186f
C16736 VDD.n787 VSS 0.278056f
C16737 VDD.t3836 VSS 0.081403f
C16738 VDD.t4716 VSS 0.080308f
C16739 VDD.t3969 VSS 0.034186f
C16740 VDD.t4717 VSS 0.034186f
C16741 VDD.n788 VSS 0.278056f
C16742 VDD.t3618 VSS 0.080308f
C16743 VDD.t2917 VSS 0.034186f
C16744 VDD.t3619 VSS 0.034186f
C16745 VDD.n789 VSS 0.278056f
C16746 VDD.t3952 VSS 0.080308f
C16747 VDD.t3227 VSS 0.034186f
C16748 VDD.t3953 VSS 0.034186f
C16749 VDD.n790 VSS 0.278056f
C16750 VDD.t3822 VSS 0.080308f
C16751 VDD.t3117 VSS 0.034186f
C16752 VDD.t3823 VSS 0.034186f
C16753 VDD.n791 VSS 0.278056f
C16754 VDD.t3960 VSS 0.080308f
C16755 VDD.t3233 VSS 0.034186f
C16756 VDD.t3961 VSS 0.034186f
C16757 VDD.n792 VSS 0.278056f
C16758 VDD.n793 VSS 0.234544f
C16759 VDD.t3232 VSS 0.080308f
C16760 VDD.n794 VSS 0.299675f
C16761 VDD.n795 VSS 0.299675f
C16762 VDD.t3116 VSS 0.080308f
C16763 VDD.n796 VSS 0.299675f
C16764 VDD.n797 VSS 0.299675f
C16765 VDD.t3226 VSS 0.080308f
C16766 VDD.n798 VSS 0.299675f
C16767 VDD.n799 VSS 0.299675f
C16768 VDD.t2916 VSS 0.080308f
C16769 VDD.n800 VSS 0.299675f
C16770 VDD.n801 VSS 0.299675f
C16771 VDD.t3968 VSS 0.080308f
C16772 VDD.n802 VSS 0.332862f
C16773 VDD.t2802 VSS 0.042371f
C16774 VDD.t1070 VSS 0.042371f
C16775 VDD.t385 VSS 0.020844f
C16776 VDD.t3837 VSS 0.034186f
C16777 VDD.n803 VSS 0.129126f
C16778 VDD.t382 VSS 0.020844f
C16779 VDD.t4125 VSS 0.034186f
C16780 VDD.n804 VSS 0.129126f
C16781 VDD.t2113 VSS 0.080309f
C16782 VDD.t2408 VSS 0.080309f
C16783 VDD.n805 VSS 0.385661f
C16784 VDD.t2114 VSS 0.034186f
C16785 VDD.t4408 VSS 0.080309f
C16786 VDD.t4638 VSS 0.080309f
C16787 VDD.n806 VSS 0.385661f
C16788 VDD.t4409 VSS 0.034186f
C16789 VDD.t4654 VSS 0.080309f
C16790 VDD.t738 VSS 0.080309f
C16791 VDD.n807 VSS 0.385661f
C16792 VDD.t4655 VSS 0.025104f
C16793 VDD.t1909 VSS 0.016021f
C16794 VDD.n808 VSS 0.144967f
C16795 VDD.t1472 VSS 0.025104f
C16796 VDD.t1471 VSS 0.080309f
C16797 VDD.t1683 VSS 0.080309f
C16798 VDD.n809 VSS 0.385661f
C16799 VDD.t1681 VSS 0.080309f
C16800 VDD.t1908 VSS 0.080309f
C16801 VDD.n810 VSS 0.24784f
C16802 VDD.t1695 VSS 0.080309f
C16803 VDD.t1929 VSS 0.080309f
C16804 VDD.n811 VSS 0.385661f
C16805 VDD.t1696 VSS 0.034186f
C16806 VDD.t1546 VSS 0.080309f
C16807 VDD.t1771 VSS 0.080309f
C16808 VDD.n812 VSS 0.385661f
C16809 VDD.t1547 VSS 0.034186f
C16810 VDD.n813 VSS 0.241596f
C16811 VDD.t310 VSS 0.020844f
C16812 VDD.t2766 VSS 0.034186f
C16813 VDD.n814 VSS 0.129126f
C16814 VDD.t4071 VSS 0.042371f
C16815 VDD.t1532 VSS 0.042371f
C16816 VDD.t2422 VSS 0.080309f
C16817 VDD.t2659 VSS 0.080309f
C16818 VDD.n815 VSS 0.385661f
C16819 VDD.t2423 VSS 0.034186f
C16820 VDD.t4660 VSS 0.080309f
C16821 VDD.t742 VSS 0.080309f
C16822 VDD.n816 VSS 0.385661f
C16823 VDD.t4661 VSS 0.034186f
C16824 VDD.t4510 VSS 0.080309f
C16825 VDD.t4738 VSS 0.080309f
C16826 VDD.n817 VSS 0.385661f
C16827 VDD.t4511 VSS 0.025104f
C16828 VDD.t4513 VSS 0.016021f
C16829 VDD.n818 VSS 0.144967f
C16830 VDD.t1700 VSS 0.025104f
C16831 VDD.t1699 VSS 0.080309f
C16832 VDD.t1933 VSS 0.080309f
C16833 VDD.n819 VSS 0.385661f
C16834 VDD.t4314 VSS 0.080309f
C16835 VDD.t4512 VSS 0.080309f
C16836 VDD.n820 VSS 0.24784f
C16837 VDD.n821 VSS 0.0787f
C16838 VDD.t3932 VSS 0.080309f
C16839 VDD.t4156 VSS 0.080309f
C16840 VDD.n822 VSS 0.385661f
C16841 VDD.t3933 VSS 0.034186f
C16842 VDD.t2747 VSS 0.082281f
C16843 VDD.n824 VSS 0.29513f
C16844 VDD.t1722 VSS 0.080308f
C16845 VDD.t2476 VSS 0.034186f
C16846 VDD.t1723 VSS 0.034186f
C16847 VDD.n825 VSS 0.278056f
C16848 VDD.t609 VSS 0.080308f
C16849 VDD.t472 VSS 0.017997f
C16850 VDD.t1250 VSS 0.034186f
C16851 VDD.t610 VSS 0.034186f
C16852 VDD.n826 VSS 0.328513f
C16853 VDD.t990 VSS 0.080308f
C16854 VDD.t1585 VSS 0.034186f
C16855 VDD.t991 VSS 0.034186f
C16856 VDD.n827 VSS 0.278056f
C16857 VDD.t873 VSS 0.080308f
C16858 VDD.t1456 VSS 0.034186f
C16859 VDD.t874 VSS 0.034186f
C16860 VDD.n828 VSS 0.278056f
C16861 VDD.t999 VSS 0.080308f
C16862 VDD.t1589 VSS 0.034186f
C16863 VDD.t1000 VSS 0.034186f
C16864 VDD.n829 VSS 0.278056f
C16865 VDD.n830 VSS 0.234544f
C16866 VDD.t1588 VSS 0.080308f
C16867 VDD.n831 VSS 0.299675f
C16868 VDD.n832 VSS 0.299675f
C16869 VDD.t1455 VSS 0.080308f
C16870 VDD.n833 VSS 0.299675f
C16871 VDD.n834 VSS 0.299675f
C16872 VDD.t1584 VSS 0.080308f
C16873 VDD.n835 VSS 0.299675f
C16874 VDD.n836 VSS 0.299675f
C16875 VDD.t1249 VSS 0.080308f
C16876 VDD.n837 VSS 0.299675f
C16877 VDD.n838 VSS 0.299675f
C16878 VDD.t2475 VSS 0.080308f
C16879 VDD.n839 VSS 0.332862f
C16880 VDD.t4137 VSS 0.034186f
C16881 VDD.t3775 VSS 0.034186f
C16882 VDD.n840 VSS 0.278056f
C16883 VDD.t3774 VSS 0.080308f
C16884 VDD.t4011 VSS 0.034186f
C16885 VDD.t3635 VSS 0.034186f
C16886 VDD.n841 VSS 0.278056f
C16887 VDD.t3634 VSS 0.080308f
C16888 VDD.t985 VSS 0.034186f
C16889 VDD.t562 VSS 0.034186f
C16890 VDD.n842 VSS 0.278056f
C16891 VDD.t560 VSS 0.080308f
C16892 VDD.t595 VSS 0.034186f
C16893 VDD.t4415 VSS 0.034186f
C16894 VDD.n843 VSS 0.278056f
C16895 VDD.t4414 VSS 0.080308f
C16896 VDD.n844 VSS 0.017494f
C16897 VDD.n845 VSS 0.304944f
C16898 VDD.n846 VSS 0.304763f
C16899 VDD.t561 VSS 7.54183f
C16900 VDD.n847 VSS 0.303418f
C16901 VDD.n848 VSS 0.304439f
C16902 VDD.t567 VSS 7.54183f
C16903 VDD.n849 VSS 0.304763f
C16904 VDD.n850 VSS 0.304944f
C16905 VDD.n851 VSS 0.234544f
C16906 VDD.n852 VSS 0.234959f
C16907 VDD.t459 VSS 0.030289f
C16908 VDD.n853 VSS 0.077802f
C16909 VDD.t425 VSS 0.008011f
C16910 VDD.t457 VSS 0.008011f
C16911 VDD.n854 VSS 0.030319f
C16912 VDD.n855 VSS 0.039264f
C16913 VDD.t442 VSS 0.008011f
C16914 VDD.t429 VSS 0.008011f
C16915 VDD.n856 VSS 0.030367f
C16916 VDD.n857 VSS 0.039375f
C16917 VDD.t440 VSS 0.030249f
C16918 VDD.n858 VSS 0.077873f
C16919 VDD.n859 VSS 0.303418f
C16920 VDD.t4338 VSS 0.080308f
C16921 VDD.t4681 VSS 0.034186f
C16922 VDD.t4339 VSS 0.034186f
C16923 VDD.n860 VSS 0.278056f
C16924 VDD.t4658 VSS 0.080308f
C16925 VDD.t882 VSS 0.034186f
C16926 VDD.t4659 VSS 0.034186f
C16927 VDD.n861 VSS 0.278056f
C16928 VDD.t3554 VSS 0.080308f
C16929 VDD.t3905 VSS 0.034186f
C16930 VDD.t3555 VSS 0.034186f
C16931 VDD.n862 VSS 0.278056f
C16932 VDD.t3666 VSS 0.080308f
C16933 VDD.t4039 VSS 0.034186f
C16934 VDD.t3667 VSS 0.034186f
C16935 VDD.n863 VSS 0.278056f
C16936 VDD.t2647 VSS 0.080308f
C16937 VDD.t2999 VSS 0.034186f
C16938 VDD.t2648 VSS 0.034186f
C16939 VDD.n864 VSS 0.278056f
C16940 VDD.t2998 VSS 0.080308f
C16941 VDD.n865 VSS 0.299675f
C16942 VDD.n866 VSS 0.299675f
C16943 VDD.t4038 VSS 0.080308f
C16944 VDD.n867 VSS 0.299675f
C16945 VDD.n868 VSS 0.299675f
C16946 VDD.t3904 VSS 0.080308f
C16947 VDD.n869 VSS 0.299675f
C16948 VDD.n870 VSS 0.299675f
C16949 VDD.t880 VSS 0.080308f
C16950 VDD.n871 VSS 0.299675f
C16951 VDD.n872 VSS 0.299675f
C16952 VDD.t4680 VSS 0.080308f
C16953 VDD.n873 VSS 0.234544f
C16954 VDD.t470 VSS 9.533179f
C16955 VDD.t660 VSS 7.54183f
C16956 VDD.n874 VSS 3.4106f
C16957 VDD.n875 VSS 0.304439f
C16958 VDD.t2027 VSS 0.080309f
C16959 VDD.n876 VSS 0.113227f
C16960 VDD.t4592 VSS 0.080309f
C16961 VDD.n877 VSS 0.17245f
C16962 VDD.t583 VSS 0.025104f
C16963 VDD.t3286 VSS 0.080309f
C16964 VDD.n878 VSS 0.17245f
C16965 VDD.t2891 VSS 0.034186f
C16966 VDD.t2198 VSS 0.034186f
C16967 VDD.n879 VSS 0.205873f
C16968 VDD.t2197 VSS 0.080308f
C16969 VDD.t4347 VSS 0.034186f
C16970 VDD.t3706 VSS 0.034186f
C16971 VDD.n880 VSS 0.278056f
C16972 VDD.t3705 VSS 0.080308f
C16973 VDD.t1283 VSS 0.034186f
C16974 VDD.t661 VSS 0.034186f
C16975 VDD.n881 VSS 0.278056f
C16976 VDD.t659 VSS 0.080308f
C16977 VDD.t3422 VSS 0.034186f
C16978 VDD.t2853 VSS 0.034186f
C16979 VDD.n882 VSS 0.278056f
C16980 VDD.t2852 VSS 0.080308f
C16981 VDD.t4499 VSS 0.034186f
C16982 VDD.t3887 VSS 0.034186f
C16983 VDD.n883 VSS 0.278056f
C16984 VDD.t3886 VSS 0.080308f
C16985 VDD.t4381 VSS 0.034186f
C16986 VDD.t3767 VSS 0.034186f
C16987 VDD.n884 VSS 0.278056f
C16988 VDD.t3766 VSS 0.080308f
C16989 VDD.n885 VSS 0.234544f
C16990 VDD.t4380 VSS 0.080308f
C16991 VDD.n886 VSS 0.299675f
C16992 VDD.n887 VSS 0.299675f
C16993 VDD.t4498 VSS 0.080308f
C16994 VDD.n888 VSS 0.299675f
C16995 VDD.n889 VSS 0.299675f
C16996 VDD.t3421 VSS 0.080308f
C16997 VDD.n890 VSS 0.299675f
C16998 VDD.n891 VSS 0.299675f
C16999 VDD.t1282 VSS 0.080308f
C17000 VDD.n892 VSS 0.299675f
C17001 VDD.n893 VSS 0.299675f
C17002 VDD.t4346 VSS 0.080308f
C17003 VDD.n894 VSS 0.348626f
C17004 VDD.n895 VSS 0.348626f
C17005 VDD.t2890 VSS 0.080308f
C17006 VDD.n896 VSS 0.357338f
C17007 VDD.t1724 VSS 0.080309f
C17008 VDD.n897 VSS 0.17245f
C17009 VDD.t1985 VSS 0.080309f
C17010 VDD.n898 VSS 0.17245f
C17011 VDD.t1747 VSS 0.016021f
C17012 VDD.t1527 VSS 0.080309f
C17013 VDD.n899 VSS 0.17245f
C17014 VDD.t3258 VSS 0.080309f
C17015 VDD.n900 VSS 0.17245f
C17016 VDD.t4462 VSS 0.080309f
C17017 VDD.n901 VSS 0.17245f
C17018 VDD.t4582 VSS 0.080309f
C17019 VDD.n902 VSS 0.17245f
C17020 VDD.t4379 VSS 0.016021f
C17021 VDD.t2826 VSS 0.080309f
C17022 VDD.n903 VSS 0.17245f
C17023 VDD.t1648 VSS 0.080309f
C17024 VDD.n904 VSS 0.17245f
C17025 VDD.n905 VSS 0.133386f
C17026 VDD.t1649 VSS 0.034186f
C17027 VDD.n906 VSS 0.129218f
C17028 VDD.n907 VSS 0.129218f
C17029 VDD.t2827 VSS 0.025104f
C17030 VDD.n908 VSS 0.016021f
C17031 VDD.n909 VSS 0.124587f
C17032 VDD.t4378 VSS 0.080309f
C17033 VDD.n910 VSS 0.113227f
C17034 VDD.n911 VSS 0.062293f
C17035 VDD.n912 VSS 0.121516f
C17036 VDD.n913 VSS 0.016021f
C17037 VDD.t4583 VSS 0.025104f
C17038 VDD.n914 VSS 0.129218f
C17039 VDD.n915 VSS 0.129218f
C17040 VDD.t4463 VSS 0.034186f
C17041 VDD.n916 VSS 0.133386f
C17042 VDD.t1348 VSS 0.034186f
C17043 VDD.t746 VSS 0.034186f
C17044 VDD.n917 VSS 0.205873f
C17045 VDD.t744 VSS 0.080308f
C17046 VDD.t2995 VSS 0.034186f
C17047 VDD.t2318 VSS 0.034186f
C17048 VDD.n918 VSS 0.278056f
C17049 VDD.t2317 VSS 0.080308f
C17050 VDD.t4037 VSS 0.034186f
C17051 VDD.t3398 VSS 0.034186f
C17052 VDD.n919 VSS 0.278056f
C17053 VDD.t3397 VSS 0.080308f
C17054 VDD.t1964 VSS 0.034186f
C17055 VDD.t1300 VSS 0.034186f
C17056 VDD.n920 VSS 0.278056f
C17057 VDD.t1299 VSS 0.080308f
C17058 VDD.t3145 VSS 0.034186f
C17059 VDD.t2527 VSS 0.034186f
C17060 VDD.n921 VSS 0.278056f
C17061 VDD.t2526 VSS 0.080308f
C17062 VDD.t3035 VSS 0.034186f
C17063 VDD.t2400 VSS 0.034186f
C17064 VDD.n922 VSS 0.278056f
C17065 VDD.t2399 VSS 0.080308f
C17066 VDD.t4081 VSS 0.034186f
C17067 VDD.t3457 VSS 0.034186f
C17068 VDD.n923 VSS 0.278056f
C17069 VDD.t3456 VSS 0.080308f
C17070 VDD.t3963 VSS 0.034186f
C17071 VDD.t3329 VSS 0.034186f
C17072 VDD.n924 VSS 0.278056f
C17073 VDD.t3328 VSS 0.080308f
C17074 VDD.t4073 VSS 0.034186f
C17075 VDD.t3453 VSS 0.034186f
C17076 VDD.n925 VSS 0.278056f
C17077 VDD.t3452 VSS 0.080308f
C17078 VDD.t480 VSS 0.017997f
C17079 VDD.t3740 VSS 0.034186f
C17080 VDD.t3161 VSS 0.034186f
C17081 VDD.n926 VSS 0.328513f
C17082 VDD.t3160 VSS 0.080308f
C17083 VDD.t482 VSS 0.017997f
C17084 VDD.t693 VSS 0.034186f
C17085 VDD.t4233 VSS 0.034186f
C17086 VDD.n927 VSS 0.328513f
C17087 VDD.t4232 VSS 0.080308f
C17088 VDD.t691 VSS 0.080308f
C17089 VDD.n928 VSS 0.299675f
C17090 VDD.n929 VSS 0.299675f
C17091 VDD.t3739 VSS 0.080308f
C17092 VDD.n930 VSS 0.299675f
C17093 VDD.n931 VSS 0.299675f
C17094 VDD.t4072 VSS 0.080308f
C17095 VDD.n932 VSS 0.299675f
C17096 VDD.n933 VSS 0.299675f
C17097 VDD.t3962 VSS 0.080308f
C17098 VDD.n934 VSS 0.299675f
C17099 VDD.n935 VSS 0.299675f
C17100 VDD.t4080 VSS 0.080308f
C17101 VDD.n936 VSS 0.234959f
C17102 VDD.t2630 VSS 0.034186f
C17103 VDD.n937 VSS 0.44766f
C17104 VDD.t2501 VSS 0.034186f
C17105 VDD.n938 VSS 0.44766f
C17106 VDD.t2624 VSS 0.034186f
C17107 VDD.n939 VSS 0.44766f
C17108 VDD.t2228 VSS 0.034186f
C17109 VDD.n940 VSS 0.44766f
C17110 VDD.t485 VSS 0.017997f
C17111 VDD.t3331 VSS 0.034186f
C17112 VDD.n941 VSS 0.498117f
C17113 VDD.t687 VSS 0.034186f
C17114 VDD.n942 VSS 0.44766f
C17115 VDD.t2622 VSS 0.034186f
C17116 VDD.t2621 VSS 0.080309f
C17117 VDD.t2830 VSS 0.080309f
C17118 VDD.n943 VSS 0.385661f
C17119 VDD.t3600 VSS 0.025104f
C17120 VDD.t3599 VSS 0.080309f
C17121 VDD.t3816 VSS 0.080309f
C17122 VDD.n944 VSS 0.385661f
C17123 VDD.t1107 VSS 0.016021f
C17124 VDD.n945 VSS 0.016021f
C17125 VDD.n946 VSS 0.289935f
C17126 VDD.n947 VSS 0.016021f
C17127 VDD.t3817 VSS 0.025104f
C17128 VDD.n948 VSS 0.223912f
C17129 VDD.t475 VSS 0.242099f
C17130 VDD.n949 VSS 0.469073f
C17131 VDD.n950 VSS 0.280724f
C17132 VDD.t2831 VSS 0.034186f
C17133 VDD.n951 VSS 0.307891f
C17134 VDD.n952 VSS 0.227298f
C17135 VDD.n953 VSS 0.018249f
C17136 VDD.n954 VSS 0.01487f
C17137 VDD.n956 VSS 0.12547f
C17138 VDD.n957 VSS 0.018625f
C17139 VDD.t941 VSS 0.034186f
C17140 VDD.n958 VSS 0.44766f
C17141 VDD.t2933 VSS 0.034186f
C17142 VDD.n959 VSS 0.44766f
C17143 VDD.t3979 VSS 0.034186f
C17144 VDD.n960 VSS 0.44766f
C17145 VDD.t3847 VSS 0.034186f
C17146 VDD.n961 VSS 0.44766f
C17147 VDD.t809 VSS 0.034186f
C17148 VDD.n962 VSS 0.44766f
C17149 VDD.t4611 VSS 0.034186f
C17150 VDD.n963 VSS 0.44766f
C17151 VDD.t1562 VSS 0.034186f
C17152 VDD.n964 VSS 0.44766f
C17153 VDD.t1434 VSS 0.034186f
C17154 VDD.n965 VSS 0.44766f
C17155 VDD.t2670 VSS 0.034186f
C17156 VDD.n966 VSS 0.44766f
C17157 VDD.t2547 VSS 0.034186f
C17158 VDD.n967 VSS 0.44766f
C17159 VDD.t484 VSS 0.017997f
C17160 VDD.t3582 VSS 0.034186f
C17161 VDD.n968 VSS 0.498117f
C17162 VDD.t3581 VSS 0.080308f
C17163 VDD.n969 VSS 0.464166f
C17164 VDD.n970 VSS 0.464166f
C17165 VDD.t2546 VSS 0.080308f
C17166 VDD.n971 VSS 0.464166f
C17167 VDD.n972 VSS 0.464166f
C17168 VDD.t2669 VSS 0.080308f
C17169 VDD.n973 VSS 0.464166f
C17170 VDD.n974 VSS 0.464166f
C17171 VDD.t1433 VSS 0.080308f
C17172 VDD.n975 VSS 0.464166f
C17173 VDD.n976 VSS 0.464166f
C17174 VDD.t1561 VSS 0.080308f
C17175 VDD.n977 VSS 0.351025f
C17176 VDD.t437 VSS 0.008011f
C17177 VDD.t423 VSS 0.008011f
C17178 VDD.n978 VSS 0.030367f
C17179 VDD.t430 VSS 0.030249f
C17180 VDD.n979 VSS 0.077873f
C17181 VDD.n980 VSS 0.039375f
C17182 VDD.t463 VSS 0.008011f
C17183 VDD.t451 VSS 0.008011f
C17184 VDD.n981 VSS 0.030319f
C17185 VDD.n982 VSS 0.039264f
C17186 VDD.t453 VSS 0.030289f
C17187 VDD.n983 VSS 0.077802f
C17188 VDD.n984 VSS 0.1297f
C17189 VDD.n985 VSS 0.113141f
C17190 VDD.n986 VSS 0.3503f
C17191 VDD.t4610 VSS 0.080308f
C17192 VDD.n987 VSS 0.464166f
C17193 VDD.n988 VSS 0.464166f
C17194 VDD.t808 VSS 0.080308f
C17195 VDD.n989 VSS 0.464166f
C17196 VDD.n990 VSS 0.464166f
C17197 VDD.t3846 VSS 0.080308f
C17198 VDD.n991 VSS 0.464166f
C17199 VDD.n992 VSS 0.464166f
C17200 VDD.t3978 VSS 0.080308f
C17201 VDD.n993 VSS 0.464166f
C17202 VDD.n994 VSS 0.464166f
C17203 VDD.t2932 VSS 0.080308f
C17204 VDD.n995 VSS 0.549746f
C17205 VDD.n996 VSS 0.549746f
C17206 VDD.t940 VSS 0.080308f
C17207 VDD.n997 VSS 0.431529f
C17208 VDD.n1000 VSS 0.009312f
C17209 VDD.n1001 VSS 0.009688f
C17210 VDD.n1002 VSS 0.271248f
C17211 VDD.n1003 VSS 0.01502f
C17212 VDD.n1004 VSS 0.316214f
C17213 VDD.n1005 VSS 0.522186f
C17214 VDD.t685 VSS 0.080308f
C17215 VDD.n1006 VSS 0.549746f
C17216 VDD.n1007 VSS 0.549746f
C17217 VDD.t3330 VSS 0.080308f
C17218 VDD.n1008 VSS 0.464166f
C17219 VDD.n1009 VSS 0.464166f
C17220 VDD.t2227 VSS 0.080308f
C17221 VDD.n1010 VSS 0.464166f
C17222 VDD.n1011 VSS 0.464166f
C17223 VDD.t2623 VSS 0.080308f
C17224 VDD.n1012 VSS 0.464166f
C17225 VDD.n1013 VSS 0.464166f
C17226 VDD.t2500 VSS 0.080308f
C17227 VDD.n1014 VSS 0.464166f
C17228 VDD.n1015 VSS 0.464166f
C17229 VDD.t2629 VSS 0.080308f
C17230 VDD.n1016 VSS 0.351025f
C17231 VDD.t1400 VSS 0.034186f
C17232 VDD.n1017 VSS 0.44766f
C17233 VDD.t1513 VSS 0.034186f
C17234 VDD.n1018 VSS 0.44766f
C17235 VDD.t4545 VSS 0.034186f
C17236 VDD.n1019 VSS 0.44766f
C17237 VDD.t2568 VSS 0.034186f
C17238 VDD.n1020 VSS 0.44766f
C17239 VDD.t1344 VSS 0.034186f
C17240 VDD.n1021 VSS 0.44766f
C17241 VDD.n1022 VSS 0.508406f
C17242 VDD.t1343 VSS 0.080308f
C17243 VDD.n1023 VSS 0.464166f
C17244 VDD.n1024 VSS 0.464166f
C17245 VDD.t2567 VSS 0.080308f
C17246 VDD.n1025 VSS 0.464166f
C17247 VDD.n1026 VSS 0.464166f
C17248 VDD.t4544 VSS 0.080308f
C17249 VDD.n1027 VSS 0.464166f
C17250 VDD.n1028 VSS 0.464166f
C17251 VDD.t1512 VSS 0.080308f
C17252 VDD.n1029 VSS 0.464166f
C17253 VDD.n1030 VSS 0.464166f
C17254 VDD.t1399 VSS 0.080308f
C17255 VDD.n1031 VSS 0.3503f
C17256 VDD.n1032 VSS 0.113141f
C17257 VDD.n1033 VSS 0.1297f
C17258 VDD.t462 VSS 0.030289f
C17259 VDD.n1034 VSS 0.077802f
C17260 VDD.t427 VSS 0.008011f
C17261 VDD.t445 VSS 0.008011f
C17262 VDD.n1035 VSS 0.030319f
C17263 VDD.n1036 VSS 0.039264f
C17264 VDD.t432 VSS 0.008011f
C17265 VDD.t435 VSS 0.008011f
C17266 VDD.n1037 VSS 0.030367f
C17267 VDD.n1038 VSS 0.039375f
C17268 VDD.t449 VSS 0.030249f
C17269 VDD.n1039 VSS 0.077873f
C17270 VDD.t454 VSS 0.008011f
C17271 VDD.t455 VSS 0.008011f
C17272 VDD.n1040 VSS 0.030367f
C17273 VDD.n1041 VSS 0.039375f
C17274 VDD.t461 VSS 0.008011f
C17275 VDD.t464 VSS 0.008011f
C17276 VDD.n1042 VSS 0.030319f
C17277 VDD.n1043 VSS 0.039264f
C17278 VDD.t448 VSS 0.030289f
C17279 VDD.n1044 VSS 0.077802f
C17280 VDD.n1045 VSS 0.096875f
C17281 VDD.n1046 VSS 0.064716f
C17282 VDD.n1047 VSS 0.234544f
C17283 VDD.t3034 VSS 0.080308f
C17284 VDD.n1048 VSS 0.299675f
C17285 VDD.n1049 VSS 0.299675f
C17286 VDD.t3144 VSS 0.080308f
C17287 VDD.n1050 VSS 0.299675f
C17288 VDD.n1051 VSS 0.299675f
C17289 VDD.t1963 VSS 0.080308f
C17290 VDD.n1052 VSS 0.299675f
C17291 VDD.n1053 VSS 0.299675f
C17292 VDD.t4036 VSS 0.080308f
C17293 VDD.n1054 VSS 0.299675f
C17294 VDD.n1055 VSS 0.299675f
C17295 VDD.t2994 VSS 0.080308f
C17296 VDD.n1056 VSS 0.348626f
C17297 VDD.n1057 VSS 0.348626f
C17298 VDD.t1347 VSS 0.080308f
C17299 VDD.n1058 VSS 0.357338f
C17300 VDD.n1059 VSS 0.250403f
C17301 VDD.n1060 VSS 0.133386f
C17302 VDD.t3259 VSS 0.034186f
C17303 VDD.n1061 VSS 0.129218f
C17304 VDD.n1062 VSS 0.129218f
C17305 VDD.t1528 VSS 0.025104f
C17306 VDD.n1063 VSS 0.016021f
C17307 VDD.n1064 VSS 0.124587f
C17308 VDD.t1746 VSS 0.080309f
C17309 VDD.n1065 VSS 0.113227f
C17310 VDD.n1066 VSS 0.062293f
C17311 VDD.n1067 VSS 0.121516f
C17312 VDD.n1068 VSS 0.016021f
C17313 VDD.t1986 VSS 0.025104f
C17314 VDD.n1069 VSS 0.129218f
C17315 VDD.n1070 VSS 0.129218f
C17316 VDD.t1725 VSS 0.034186f
C17317 VDD.n1071 VSS 0.133386f
C17318 VDD.n1072 VSS 0.250403f
C17319 VDD.n1073 VSS 0.133386f
C17320 VDD.t3287 VSS 0.034186f
C17321 VDD.n1074 VSS 0.129218f
C17322 VDD.n1075 VSS 0.129218f
C17323 VDD.t582 VSS 0.080309f
C17324 VDD.n1076 VSS 0.17245f
C17325 VDD.n1077 VSS 0.124587f
C17326 VDD.n1078 VSS 0.016021f
C17327 VDD.t2028 VSS 0.016021f
C17328 VDD.t1995 VSS 0.080309f
C17329 VDD.n1079 VSS 0.17245f
C17330 VDD.t3498 VSS 0.080309f
C17331 VDD.n1080 VSS 0.17245f
C17332 VDD.t891 VSS 0.080309f
C17333 VDD.n1081 VSS 0.17245f
C17334 VDD.t3479 VSS 0.016021f
C17335 VDD.n1082 VSS 0.121516f
C17336 VDD.n1083 VSS 0.303418f
C17337 VDD.t317 VSS 9.533179f
C17338 VDD.t315 VSS 7.734359f
C17339 VDD.t319 VSS 3.20156f
C17340 VDD.n1084 VSS 3.4106f
C17341 VDD.n1085 VSS 0.234544f
C17342 VDD.t371 VSS 0.030289f
C17343 VDD.n1086 VSS 0.077802f
C17344 VDD.t347 VSS 0.008011f
C17345 VDD.t357 VSS 0.008011f
C17346 VDD.n1087 VSS 0.030319f
C17347 VDD.n1088 VSS 0.039264f
C17348 VDD.t340 VSS 0.008011f
C17349 VDD.t358 VSS 0.008011f
C17350 VDD.n1089 VSS 0.030367f
C17351 VDD.n1090 VSS 0.039375f
C17352 VDD.t487 VSS 0.030249f
C17353 VDD.n1091 VSS 0.077873f
C17354 VDD.t3344 VSS 0.080308f
C17355 VDD.t4719 VSS 0.034186f
C17356 VDD.t3345 VSS 0.034186f
C17357 VDD.n1092 VSS 0.278056f
C17358 VDD.t3656 VSS 0.080308f
C17359 VDD.t926 VSS 0.034186f
C17360 VDD.t3657 VSS 0.034186f
C17361 VDD.n1093 VSS 0.278056f
C17362 VDD.t2639 VSS 0.080308f
C17363 VDD.t3957 VSS 0.034186f
C17364 VDD.t2640 VSS 0.034186f
C17365 VDD.n1094 VSS 0.278056f
C17366 VDD.n1095 VSS 0.299675f
C17367 VDD.t3956 VSS 0.080308f
C17368 VDD.n1096 VSS 0.299675f
C17369 VDD.n1097 VSS 0.299675f
C17370 VDD.t925 VSS 0.080308f
C17371 VDD.n1098 VSS 0.299675f
C17372 VDD.n1099 VSS 0.299675f
C17373 VDD.t4718 VSS 0.080308f
C17374 VDD.n1100 VSS 0.234959f
C17375 VDD.t362 VSS 0.008011f
C17376 VDD.t372 VSS 0.008011f
C17377 VDD.n1101 VSS 0.030367f
C17378 VDD.n1102 VSS 0.039375f
C17379 VDD.t370 VSS 0.008011f
C17380 VDD.t335 VSS 0.008011f
C17381 VDD.n1103 VSS 0.030319f
C17382 VDD.n1104 VSS 0.039264f
C17383 VDD.t352 VSS 0.030289f
C17384 VDD.n1105 VSS 0.077802f
C17385 VDD.n1106 VSS 0.096875f
C17386 VDD.t1705 VSS 0.080309f
C17387 VDD.n1107 VSS 0.113227f
C17388 VDD.t1845 VSS 0.080309f
C17389 VDD.n1108 VSS 0.17245f
C17390 VDD.t4675 VSS 0.025104f
C17391 VDD.t3194 VSS 0.080309f
C17392 VDD.n1109 VSS 0.17245f
C17393 VDD.t2479 VSS 0.080309f
C17394 VDD.n1110 VSS 0.17245f
C17395 VDD.t4670 VSS 0.080309f
C17396 VDD.n1111 VSS 0.17245f
C17397 VDD.t3485 VSS 0.016021f
C17398 VDD.t3658 VSS 0.080309f
C17399 VDD.n1112 VSS 0.17245f
C17400 VDD.t720 VSS 0.080309f
C17401 VDD.n1113 VSS 0.17245f
C17402 VDD.t4730 VSS 0.080309f
C17403 VDD.n1114 VSS 0.17245f
C17404 VDD.t1761 VSS 0.080309f
C17405 VDD.n1115 VSS 0.17245f
C17406 VDD.t1990 VSS 0.016021f
C17407 VDD.t4566 VSS 0.080309f
C17408 VDD.n1116 VSS 0.17245f
C17409 VDD.t1629 VSS 0.080309f
C17410 VDD.n1117 VSS 0.17245f
C17411 VDD.n1118 VSS 0.357338f
C17412 VDD.t954 VSS 0.034186f
C17413 VDD.t2248 VSS 0.034186f
C17414 VDD.t2247 VSS 0.080308f
C17415 VDD.t3318 VSS 0.080308f
C17416 VDD.t479 VSS 0.017997f
C17417 VDD.t3627 VSS 0.034186f
C17418 VDD.t3319 VSS 0.034186f
C17419 VDD.n1119 VSS 0.328513f
C17420 VDD.t2190 VSS 0.080308f
C17421 VDD.t478 VSS 0.017997f
C17422 VDD.t2608 VSS 0.034186f
C17423 VDD.t2191 VSS 0.034186f
C17424 VDD.n1120 VSS 0.328513f
C17425 VDD.t2368 VSS 0.080308f
C17426 VDD.t2727 VSS 0.034186f
C17427 VDD.t2369 VSS 0.034186f
C17428 VDD.n1121 VSS 0.278056f
C17429 VDD.t1162 VSS 0.080308f
C17430 VDD.t1500 VSS 0.034186f
C17431 VDD.t1163 VSS 0.034186f
C17432 VDD.n1122 VSS 0.278056f
C17433 VDD.t1276 VSS 0.080308f
C17434 VDD.t1632 VSS 0.034186f
C17435 VDD.t1277 VSS 0.034186f
C17436 VDD.n1123 VSS 0.278056f
C17437 VDD.t1631 VSS 0.080308f
C17438 VDD.n1124 VSS 0.299675f
C17439 VDD.n1125 VSS 0.299675f
C17440 VDD.t1499 VSS 0.080308f
C17441 VDD.n1126 VSS 0.299675f
C17442 VDD.n1127 VSS 0.299675f
C17443 VDD.t2726 VSS 0.080308f
C17444 VDD.n1128 VSS 0.299675f
C17445 VDD.n1129 VSS 0.299675f
C17446 VDD.t2607 VSS 0.080308f
C17447 VDD.n1130 VSS 0.299675f
C17448 VDD.n1131 VSS 0.299675f
C17449 VDD.t3626 VSS 0.080308f
C17450 VDD.n1132 VSS 0.348626f
C17451 VDD.t953 VSS 0.080308f
C17452 VDD.n1133 VSS 0.348626f
C17453 VDD.n1134 VSS 0.205873f
C17454 VDD.t1479 VSS 0.080309f
C17455 VDD.n1135 VSS 0.17245f
C17456 VDD.t4140 VSS 0.080309f
C17457 VDD.n1136 VSS 0.17245f
C17458 VDD.t3005 VSS 0.016021f
C17459 VDD.t1685 VSS 0.080309f
C17460 VDD.n1137 VSS 0.17245f
C17461 VDD.t1218 VSS 0.080309f
C17462 VDD.n1138 VSS 0.17245f
C17463 VDD.n1139 VSS 0.357338f
C17464 VDD.t3608 VSS 0.034186f
C17465 VDD.t754 VSS 0.034186f
C17466 VDD.t753 VSS 0.080308f
C17467 VDD.t3914 VSS 0.080308f
C17468 VDD.t483 VSS 0.017997f
C17469 VDD.t4265 VSS 0.034186f
C17470 VDD.t3915 VSS 0.034186f
C17471 VDD.n1140 VSS 0.328513f
C17472 VDD.t2876 VSS 0.080308f
C17473 VDD.t476 VSS 0.017997f
C17474 VDD.t3197 VSS 0.034186f
C17475 VDD.t2877 VSS 0.034186f
C17476 VDD.n1141 VSS 0.328513f
C17477 VDD.t3006 VSS 0.080308f
C17478 VDD.t3303 VSS 0.034186f
C17479 VDD.t3007 VSS 0.034186f
C17480 VDD.n1142 VSS 0.278056f
C17481 VDD.t1773 VSS 0.080308f
C17482 VDD.t2162 VSS 0.034186f
C17483 VDD.t1774 VSS 0.034186f
C17484 VDD.n1143 VSS 0.278056f
C17485 VDD.t1914 VSS 0.080308f
C17486 VDD.t2324 VSS 0.034186f
C17487 VDD.t1915 VSS 0.034186f
C17488 VDD.n1144 VSS 0.278056f
C17489 VDD.n1145 VSS 0.234959f
C17490 VDD.t2323 VSS 0.080308f
C17491 VDD.n1146 VSS 0.299675f
C17492 VDD.n1147 VSS 0.299675f
C17493 VDD.t2161 VSS 0.080308f
C17494 VDD.n1148 VSS 0.299675f
C17495 VDD.n1149 VSS 0.299675f
C17496 VDD.t3302 VSS 0.080308f
C17497 VDD.n1150 VSS 0.299675f
C17498 VDD.n1151 VSS 0.299675f
C17499 VDD.t3196 VSS 0.080308f
C17500 VDD.n1152 VSS 0.299675f
C17501 VDD.n1153 VSS 0.299675f
C17502 VDD.t4264 VSS 0.080308f
C17503 VDD.n1154 VSS 0.348626f
C17504 VDD.t3607 VSS 0.080308f
C17505 VDD.n1155 VSS 0.348626f
C17506 VDD.n1156 VSS 0.205873f
C17507 VDD.t4198 VSS 0.080309f
C17508 VDD.n1157 VSS 0.17245f
C17509 VDD.t1679 VSS 0.080309f
C17510 VDD.n1158 VSS 0.17245f
C17511 VDD.n1159 VSS 0.016021f
C17512 VDD.t1680 VSS 0.025104f
C17513 VDD.n1160 VSS 0.129218f
C17514 VDD.n1161 VSS 0.129218f
C17515 VDD.t4199 VSS 0.034186f
C17516 VDD.n1162 VSS 0.133386f
C17517 VDD.n1163 VSS 0.250403f
C17518 VDD.n1164 VSS 0.133386f
C17519 VDD.t1219 VSS 0.034186f
C17520 VDD.n1165 VSS 0.129218f
C17521 VDD.n1166 VSS 0.129218f
C17522 VDD.t1686 VSS 0.025104f
C17523 VDD.n1167 VSS 0.016021f
C17524 VDD.n1168 VSS 0.124587f
C17525 VDD.t3004 VSS 0.080309f
C17526 VDD.n1169 VSS 0.113227f
C17527 VDD.n1170 VSS 0.062293f
C17528 VDD.n1171 VSS 0.121516f
C17529 VDD.n1172 VSS 0.016021f
C17530 VDD.t4141 VSS 0.025104f
C17531 VDD.n1173 VSS 0.129218f
C17532 VDD.n1174 VSS 0.129218f
C17533 VDD.t1480 VSS 0.034186f
C17534 VDD.n1175 VSS 0.133386f
C17535 VDD.n1176 VSS 0.250403f
C17536 VDD.n1177 VSS 0.133386f
C17537 VDD.t1630 VSS 0.034186f
C17538 VDD.n1178 VSS 0.129218f
C17539 VDD.n1179 VSS 0.129218f
C17540 VDD.t4567 VSS 0.025104f
C17541 VDD.n1180 VSS 0.016021f
C17542 VDD.n1181 VSS 0.124587f
C17543 VDD.t1989 VSS 0.080309f
C17544 VDD.n1182 VSS 0.113227f
C17545 VDD.n1183 VSS 0.062293f
C17546 VDD.n1184 VSS 0.121516f
C17547 VDD.n1185 VSS 0.016021f
C17548 VDD.t1762 VSS 0.025104f
C17549 VDD.n1186 VSS 0.129218f
C17550 VDD.n1187 VSS 0.129218f
C17551 VDD.t4731 VSS 0.034186f
C17552 VDD.n1188 VSS 0.133386f
C17553 VDD.n1189 VSS 0.357338f
C17554 VDD.t4181 VSS 0.034186f
C17555 VDD.t1273 VSS 0.034186f
C17556 VDD.t1272 VSS 0.080308f
C17557 VDD.t3387 VSS 0.080308f
C17558 VDD.t3724 VSS 0.034186f
C17559 VDD.t3388 VSS 0.034186f
C17560 VDD.n1190 VSS 0.278056f
C17561 VDD.t2313 VSS 0.080308f
C17562 VDD.t477 VSS 0.017997f
C17563 VDD.t2699 VSS 0.034186f
C17564 VDD.t2314 VSS 0.034186f
C17565 VDD.n1191 VSS 0.328513f
C17566 VDD.t2477 VSS 0.080308f
C17567 VDD.t2821 VSS 0.034186f
C17568 VDD.t2478 VSS 0.034186f
C17569 VDD.n1192 VSS 0.278056f
C17570 VDD.t1256 VSS 0.080308f
C17571 VDD.t1601 VSS 0.034186f
C17572 VDD.t1257 VSS 0.034186f
C17573 VDD.n1193 VSS 0.278056f
C17574 VDD.t1378 VSS 0.080308f
C17575 VDD.t1719 VSS 0.034186f
C17576 VDD.t1379 VSS 0.034186f
C17577 VDD.n1194 VSS 0.278056f
C17578 VDD.t1718 VSS 0.080308f
C17579 VDD.n1195 VSS 0.299675f
C17580 VDD.n1196 VSS 0.299675f
C17581 VDD.t1600 VSS 0.080308f
C17582 VDD.n1197 VSS 0.299675f
C17583 VDD.n1198 VSS 0.299675f
C17584 VDD.t2820 VSS 0.080308f
C17585 VDD.n1199 VSS 0.299675f
C17586 VDD.n1200 VSS 0.299675f
C17587 VDD.t2698 VSS 0.080308f
C17588 VDD.n1201 VSS 0.299675f
C17589 VDD.n1202 VSS 0.299675f
C17590 VDD.t3723 VSS 0.080308f
C17591 VDD.n1203 VSS 0.348626f
C17592 VDD.t4180 VSS 0.080308f
C17593 VDD.n1204 VSS 0.348626f
C17594 VDD.n1205 VSS 0.205873f
C17595 VDD.n1206 VSS 0.250403f
C17596 VDD.n1207 VSS 0.133386f
C17597 VDD.t721 VSS 0.034186f
C17598 VDD.n1208 VSS 0.129218f
C17599 VDD.n1209 VSS 0.129218f
C17600 VDD.t3659 VSS 0.025104f
C17601 VDD.n1210 VSS 0.016021f
C17602 VDD.n1211 VSS 0.124587f
C17603 VDD.t3484 VSS 0.080309f
C17604 VDD.n1212 VSS 0.113227f
C17605 VDD.n1213 VSS 0.062293f
C17606 VDD.n1214 VSS 0.121516f
C17607 VDD.n1215 VSS 0.016021f
C17608 VDD.t4671 VSS 0.025104f
C17609 VDD.n1216 VSS 0.129218f
C17610 VDD.n1217 VSS 0.129218f
C17611 VDD.t2480 VSS 0.034186f
C17612 VDD.n1218 VSS 0.133386f
C17613 VDD.n1219 VSS 0.357338f
C17614 VDD.t1787 VSS 0.034186f
C17615 VDD.t4205 VSS 0.034186f
C17616 VDD.t4204 VSS 0.080308f
C17617 VDD.t2360 VSS 0.080308f
C17618 VDD.t3671 VSS 0.034186f
C17619 VDD.t2361 VSS 0.034186f
C17620 VDD.n1220 VSS 0.278056f
C17621 VDD.t1151 VSS 0.080308f
C17622 VDD.t2650 VSS 0.034186f
C17623 VDD.t1152 VSS 0.034186f
C17624 VDD.n1221 VSS 0.278056f
C17625 VDD.t1270 VSS 0.080308f
C17626 VDD.t2784 VSS 0.034186f
C17627 VDD.t1271 VSS 0.034186f
C17628 VDD.n1222 VSS 0.278056f
C17629 VDD.t4334 VSS 0.080308f
C17630 VDD.t1536 VSS 0.034186f
C17631 VDD.t4335 VSS 0.034186f
C17632 VDD.n1223 VSS 0.278056f
C17633 VDD.t4446 VSS 0.080308f
C17634 VDD.t1670 VSS 0.034186f
C17635 VDD.t4447 VSS 0.034186f
C17636 VDD.n1224 VSS 0.278056f
C17637 VDD.t1669 VSS 0.080308f
C17638 VDD.n1225 VSS 0.299675f
C17639 VDD.n1226 VSS 0.299675f
C17640 VDD.t1535 VSS 0.080308f
C17641 VDD.n1227 VSS 0.299675f
C17642 VDD.n1228 VSS 0.299675f
C17643 VDD.t2783 VSS 0.080308f
C17644 VDD.n1229 VSS 0.299675f
C17645 VDD.n1230 VSS 0.299675f
C17646 VDD.t2649 VSS 0.080308f
C17647 VDD.n1231 VSS 0.299675f
C17648 VDD.n1232 VSS 0.299675f
C17649 VDD.t3670 VSS 0.080308f
C17650 VDD.n1233 VSS 0.348626f
C17651 VDD.t1786 VSS 0.080308f
C17652 VDD.n1234 VSS 0.348626f
C17653 VDD.n1235 VSS 0.205873f
C17654 VDD.n1236 VSS 0.250403f
C17655 VDD.n1237 VSS 0.133386f
C17656 VDD.t3195 VSS 0.034186f
C17657 VDD.n1238 VSS 0.129218f
C17658 VDD.n1239 VSS 0.129218f
C17659 VDD.t4674 VSS 0.080309f
C17660 VDD.n1240 VSS 0.17245f
C17661 VDD.n1241 VSS 0.124587f
C17662 VDD.n1242 VSS 0.016021f
C17663 VDD.t1706 VSS 0.016021f
C17664 VDD.t3419 VSS 0.080309f
C17665 VDD.n1243 VSS 0.17245f
C17666 VDD.t4598 VSS 0.080309f
C17667 VDD.n1244 VSS 0.17245f
C17668 VDD.t3434 VSS 0.080309f
C17669 VDD.n1245 VSS 0.17245f
C17670 VDD.n1246 VSS 0.124587f
C17671 VDD.n1247 VSS 0.016021f
C17672 VDD.t3435 VSS 0.025104f
C17673 VDD.n1248 VSS 0.129218f
C17674 VDD.n1249 VSS 0.129218f
C17675 VDD.t4599 VSS 0.034186f
C17676 VDD.n1250 VSS 0.133386f
C17677 VDD.n1251 VSS 0.357338f
C17678 VDD.t2907 VSS 0.034186f
C17679 VDD.t1043 VSS 0.034186f
C17680 VDD.t1042 VSS 0.080308f
C17681 VDD.t3466 VSS 0.080308f
C17682 VDD.t666 VSS 0.034186f
C17683 VDD.t3467 VSS 0.034186f
C17684 VDD.n1252 VSS 0.278056f
C17685 VDD.t2406 VSS 0.080308f
C17686 VDD.t3716 VSS 0.034186f
C17687 VDD.t2407 VSS 0.034186f
C17688 VDD.n1253 VSS 0.278056f
C17689 VDD.t2532 VSS 0.080308f
C17690 VDD.t3839 VSS 0.034186f
C17691 VDD.t2533 VSS 0.034186f
C17692 VDD.n1254 VSS 0.278056f
C17693 VDD.t1304 VSS 0.080308f
C17694 VDD.t2812 VSS 0.034186f
C17695 VDD.t1305 VSS 0.034186f
C17696 VDD.n1255 VSS 0.278056f
C17697 VDD.t1429 VSS 0.080308f
C17698 VDD.t2919 VSS 0.034186f
C17699 VDD.t1430 VSS 0.034186f
C17700 VDD.n1256 VSS 0.278056f
C17701 VDD.n1257 VSS 0.234544f
C17702 VDD.t2918 VSS 0.080308f
C17703 VDD.n1258 VSS 0.299675f
C17704 VDD.n1259 VSS 0.299675f
C17705 VDD.t2811 VSS 0.080308f
C17706 VDD.n1260 VSS 0.299675f
C17707 VDD.n1261 VSS 0.299675f
C17708 VDD.t3838 VSS 0.080308f
C17709 VDD.n1262 VSS 0.299675f
C17710 VDD.n1263 VSS 0.299675f
C17711 VDD.t3715 VSS 0.080308f
C17712 VDD.n1264 VSS 0.299675f
C17713 VDD.n1265 VSS 0.299675f
C17714 VDD.t664 VSS 0.080308f
C17715 VDD.n1266 VSS 0.348626f
C17716 VDD.t2906 VSS 0.080308f
C17717 VDD.n1267 VSS 0.348626f
C17718 VDD.n1268 VSS 0.205873f
C17719 VDD.n1269 VSS 0.250403f
C17720 VDD.n1270 VSS 0.133386f
C17721 VDD.t3420 VSS 0.034186f
C17722 VDD.n1271 VSS 0.129218f
C17723 VDD.n1272 VSS 0.129218f
C17724 VDD.t1846 VSS 0.025104f
C17725 VDD.n1273 VSS 0.016021f
C17726 VDD.n1274 VSS 0.121516f
C17727 VDD.n1275 VSS 0.062293f
C17728 VDD.n1276 VSS 0.304763f
C17729 VDD.n1277 VSS 0.303418f
C17730 VDD.t703 VSS 7.54183f
C17731 VDD.t316 VSS 9.533179f
C17732 VDD.t332 VSS 7.734359f
C17733 VDD.t320 VSS 3.18057f
C17734 VDD.t866 VSS 0.080309f
C17735 VDD.n1278 VSS 0.113227f
C17736 VDD.t3798 VSS 0.080309f
C17737 VDD.n1279 VSS 0.17245f
C17738 VDD.t593 VSS 0.025104f
C17739 VDD.t883 VSS 0.080309f
C17740 VDD.n1280 VSS 0.17245f
C17741 VDD.t3812 VSS 0.080309f
C17742 VDD.n1281 VSS 0.17245f
C17743 VDD.t3668 VSS 0.080309f
C17744 VDD.n1282 VSS 0.17245f
C17745 VDD.n1283 VSS 0.016021f
C17746 VDD.t3669 VSS 0.025104f
C17747 VDD.n1284 VSS 0.129218f
C17748 VDD.n1285 VSS 0.129218f
C17749 VDD.t3813 VSS 0.034186f
C17750 VDD.n1286 VSS 0.133386f
C17751 VDD.t704 VSS 0.034186f
C17752 VDD.t1458 VSS 0.034186f
C17753 VDD.n1287 VSS 0.205873f
C17754 VDD.t1457 VSS 0.080308f
C17755 VDD.t380 VSS 0.017997f
C17756 VDD.t2279 VSS 0.034186f
C17757 VDD.t3089 VSS 0.034186f
C17758 VDD.n1288 VSS 0.328513f
C17759 VDD.t3088 VSS 0.080308f
C17760 VDD.t381 VSS 0.017997f
C17761 VDD.t3364 VSS 0.034186f
C17762 VDD.t4155 VSS 0.034186f
C17763 VDD.n1289 VSS 0.328513f
C17764 VDD.t4154 VSS 0.080308f
C17765 VDD.t1281 VSS 0.034186f
C17766 VDD.t2094 VSS 0.034186f
C17767 VDD.n1290 VSS 0.278056f
C17768 VDD.t2093 VSS 0.080308f
C17769 VDD.t2511 VSS 0.034186f
C17770 VDD.t3253 VSS 0.034186f
C17771 VDD.n1291 VSS 0.278056f
C17772 VDD.t3252 VSS 0.080308f
C17773 VDD.t2371 VSS 0.034186f
C17774 VDD.t3139 VSS 0.034186f
C17775 VDD.n1292 VSS 0.278056f
C17776 VDD.t3138 VSS 0.080308f
C17777 VDD.t2370 VSS 0.080308f
C17778 VDD.n1293 VSS 0.299675f
C17779 VDD.n1294 VSS 0.299675f
C17780 VDD.t2510 VSS 0.080308f
C17781 VDD.n1295 VSS 0.299675f
C17782 VDD.n1296 VSS 0.299675f
C17783 VDD.t1280 VSS 0.080308f
C17784 VDD.n1297 VSS 0.299675f
C17785 VDD.n1298 VSS 0.299675f
C17786 VDD.t3363 VSS 0.080308f
C17787 VDD.n1299 VSS 0.299675f
C17788 VDD.n1300 VSS 0.299675f
C17789 VDD.t2278 VSS 0.080308f
C17790 VDD.n1301 VSS 0.348626f
C17791 VDD.n1302 VSS 0.348626f
C17792 VDD.t702 VSS 0.080308f
C17793 VDD.n1303 VSS 0.357338f
C17794 VDD.n1304 VSS 0.250403f
C17795 VDD.n1305 VSS 0.133386f
C17796 VDD.t884 VSS 0.034186f
C17797 VDD.n1306 VSS 0.129218f
C17798 VDD.n1307 VSS 0.129218f
C17799 VDD.t592 VSS 0.080309f
C17800 VDD.n1308 VSS 0.17245f
C17801 VDD.n1309 VSS 0.124587f
C17802 VDD.n1310 VSS 0.016021f
C17803 VDD.t867 VSS 0.016021f
C17804 VDD.t3573 VSS 0.080309f
C17805 VDD.n1311 VSS 0.17245f
C17806 VDD.t2378 VSS 0.080309f
C17807 VDD.n1312 VSS 0.17245f
C17808 VDD.t3848 VSS 0.080309f
C17809 VDD.n1313 VSS 0.17245f
C17810 VDD.n1314 VSS 0.124587f
C17811 VDD.n1315 VSS 0.016021f
C17812 VDD.t3849 VSS 0.025104f
C17813 VDD.n1316 VSS 0.129218f
C17814 VDD.n1317 VSS 0.129218f
C17815 VDD.t2379 VSS 0.034186f
C17816 VDD.n1318 VSS 0.133386f
C17817 VDD.t4609 VSS 0.034186f
C17818 VDD.t1224 VSS 0.034186f
C17819 VDD.n1319 VSS 0.205873f
C17820 VDD.t1223 VSS 0.080308f
C17821 VDD.t378 VSS 0.017997f
C17822 VDD.t2003 VSS 0.034186f
C17823 VDD.t2859 VSS 0.034186f
C17824 VDD.n1320 VSS 0.328513f
C17825 VDD.t2858 VSS 0.080308f
C17826 VDD.t384 VSS 0.017997f
C17827 VDD.t3181 VSS 0.034186f
C17828 VDD.t3895 VSS 0.034186f
C17829 VDD.n1321 VSS 0.328513f
C17830 VDD.t3894 VSS 0.080308f
C17831 VDD.t1072 VSS 0.034186f
C17832 VDD.t1814 VSS 0.034186f
C17833 VDD.n1322 VSS 0.278056f
C17834 VDD.t1813 VSS 0.080308f
C17835 VDD.t2202 VSS 0.034186f
C17836 VDD.t3033 VSS 0.034186f
C17837 VDD.n1323 VSS 0.278056f
C17838 VDD.t3032 VSS 0.080308f
C17839 VDD.t2075 VSS 0.034186f
C17840 VDD.t2911 VSS 0.034186f
C17841 VDD.n1324 VSS 0.278056f
C17842 VDD.t2910 VSS 0.080308f
C17843 VDD.t2074 VSS 0.080308f
C17844 VDD.n1325 VSS 0.299675f
C17845 VDD.n1326 VSS 0.299675f
C17846 VDD.t2201 VSS 0.080308f
C17847 VDD.n1327 VSS 0.299675f
C17848 VDD.n1328 VSS 0.299675f
C17849 VDD.t1071 VSS 0.080308f
C17850 VDD.n1329 VSS 0.299675f
C17851 VDD.n1330 VSS 0.299675f
C17852 VDD.t3180 VSS 0.080308f
C17853 VDD.n1331 VSS 0.299675f
C17854 VDD.n1332 VSS 0.299675f
C17855 VDD.t2002 VSS 0.080308f
C17856 VDD.n1333 VSS 0.348626f
C17857 VDD.n1334 VSS 0.348626f
C17858 VDD.t4608 VSS 0.080308f
C17859 VDD.n1335 VSS 0.357338f
C17860 VDD.n1336 VSS 0.250403f
C17861 VDD.n1337 VSS 0.133386f
C17862 VDD.t3574 VSS 0.034186f
C17863 VDD.n1338 VSS 0.129218f
C17864 VDD.n1339 VSS 0.129218f
C17865 VDD.t3799 VSS 0.025104f
C17866 VDD.n1340 VSS 0.016021f
C17867 VDD.n1341 VSS 0.121516f
C17868 VDD.n1342 VSS 0.062293f
C17869 VDD.n1343 VSS 0.304944f
C17870 VDD.t313 VSS 7.65735f
C17871 VDD.n1344 VSS 0.304439f
C17872 VDD.t308 VSS 9.533179f
C17873 VDD.t657 VSS 7.54183f
C17874 VDD.t311 VSS 7.734359f
C17875 VDD.t312 VSS 9.533179f
C17876 VDD.t665 VSS 7.54183f
C17877 VDD.n1345 VSS 3.4106f
C17878 VDD.n1346 VSS 3.4106f
C17879 VDD.n1347 VSS 0.303418f
C17880 VDD.n1348 VSS 0.304763f
C17881 VDD.n1349 VSS 3.12105f
C17882 VDD.n1350 VSS 0.304944f
C17883 VDD.n1351 VSS 0.304439f
C17884 VDD.n1352 VSS 0.064716f
C17885 VDD.n1353 VSS 0.303418f
C17886 VDD.n1354 VSS 3.4106f
C17887 VDD.t821 VSS 7.54183f
C17888 VDD.t309 VSS 9.533179f
C17889 VDD.t318 VSS 7.65735f
C17890 VDD.n1355 VSS 0.304763f
C17891 VDD.n1356 VSS 3.12455f
C17892 VDD.n1357 VSS 0.304944f
C17893 VDD.n1358 VSS 0.062293f
C17894 VDD.t3478 VSS 0.080309f
C17895 VDD.n1359 VSS 0.113227f
C17896 VDD.n1360 VSS 0.124587f
C17897 VDD.n1361 VSS 0.016021f
C17898 VDD.t892 VSS 0.025104f
C17899 VDD.n1362 VSS 0.129218f
C17900 VDD.n1363 VSS 0.129218f
C17901 VDD.t3499 VSS 0.034186f
C17902 VDD.n1364 VSS 0.133386f
C17903 VDD.t3121 VSS 0.034186f
C17904 VDD.t2515 VSS 0.034186f
C17905 VDD.n1365 VSS 0.205873f
C17906 VDD.t2514 VSS 0.080308f
C17907 VDD.t388 VSS 0.017997f
C17908 VDD.t4565 VSS 0.034186f
C17909 VDD.t3973 VSS 0.034186f
C17910 VDD.n1366 VSS 0.328513f
C17911 VDD.t3972 VSS 0.080308f
C17912 VDD.t1526 VSS 0.034186f
C17913 VDD.t943 VSS 0.034186f
C17914 VDD.n1367 VSS 0.278056f
C17915 VDD.t942 VSS 0.080308f
C17916 VDD.t3637 VSS 0.034186f
C17917 VDD.t3087 VSS 0.034186f
C17918 VDD.n1368 VSS 0.278056f
C17919 VDD.t3086 VSS 0.080308f
C17920 VDD.t568 VSS 0.034186f
C17921 VDD.t4147 VSS 0.034186f
C17922 VDD.n1369 VSS 0.278056f
C17923 VDD.t4146 VSS 0.080308f
C17924 VDD.t4633 VSS 0.034186f
C17925 VDD.t4023 VSS 0.034186f
C17926 VDD.n1370 VSS 0.278056f
C17927 VDD.t4022 VSS 0.080308f
C17928 VDD.n1371 VSS 0.234544f
C17929 VDD.t4632 VSS 0.080308f
C17930 VDD.n1372 VSS 0.299675f
C17931 VDD.n1373 VSS 0.299675f
C17932 VDD.t566 VSS 0.080308f
C17933 VDD.n1374 VSS 0.299675f
C17934 VDD.n1375 VSS 0.299675f
C17935 VDD.t3636 VSS 0.080308f
C17936 VDD.n1376 VSS 0.299675f
C17937 VDD.n1377 VSS 0.299675f
C17938 VDD.t1525 VSS 0.080308f
C17939 VDD.n1378 VSS 0.299675f
C17940 VDD.n1379 VSS 0.299675f
C17941 VDD.t4564 VSS 0.080308f
C17942 VDD.n1380 VSS 0.348626f
C17943 VDD.n1381 VSS 0.348626f
C17944 VDD.t3120 VSS 0.080308f
C17945 VDD.n1382 VSS 0.357338f
C17946 VDD.n1383 VSS 0.250403f
C17947 VDD.n1384 VSS 0.133386f
C17948 VDD.t1996 VSS 0.034186f
C17949 VDD.n1385 VSS 0.129218f
C17950 VDD.n1386 VSS 0.129218f
C17951 VDD.t4593 VSS 0.025104f
C17952 VDD.n1387 VSS 0.016021f
C17953 VDD.n1388 VSS 0.121516f
C17954 VDD.n1389 VSS 0.062293f
C17955 VDD.n1390 VSS 0.304763f
C17956 VDD.t468 VSS 9.533179f
C17957 VDD.t433 VSS 7.65735f
C17958 VDD.t2968 VSS 0.080309f
C17959 VDD.t3158 VSS 0.080309f
C17960 VDD.n1391 VSS 0.24784f
C17961 VDD.n1392 VSS 0.016021f
C17962 VDD.t1297 VSS 0.080309f
C17963 VDD.t1510 VSS 0.080309f
C17964 VDD.n1393 VSS 0.385661f
C17965 VDD.t1676 VSS 0.025104f
C17966 VDD.t1449 VSS 0.080309f
C17967 VDD.t1675 VSS 0.080309f
C17968 VDD.n1394 VSS 0.385661f
C17969 VDD.t4116 VSS 0.080309f
C17970 VDD.t4312 VSS 0.080309f
C17971 VDD.n1395 VSS 0.385661f
C17972 VDD.t4117 VSS 0.034186f
C17973 VDD.t3662 VSS 0.080309f
C17974 VDD.t3890 VSS 0.080309f
C17975 VDD.n1396 VSS 0.385661f
C17976 VDD.t3663 VSS 0.034186f
C17977 VDD.t3891 VSS 0.034186f
C17978 VDD.n1397 VSS 0.327288f
C17979 VDD.n1398 VSS 0.327288f
C17980 VDD.t4313 VSS 0.034186f
C17981 VDD.n1399 VSS 0.298193f
C17982 VDD.n1400 VSS 0.298193f
C17983 VDD.t1450 VSS 0.025104f
C17984 VDD.t2969 VSS 0.016021f
C17985 VDD.n1401 VSS 0.016021f
C17986 VDD.n1402 VSS 0.289935f
C17987 VDD.n1403 VSS 0.016021f
C17988 VDD.t3159 VSS 0.016021f
C17989 VDD.t1298 VSS 0.025104f
C17990 VDD.t2955 VSS 0.034186f
C17991 VDD.t2954 VSS 0.080309f
C17992 VDD.t3146 VSS 0.080309f
C17993 VDD.n1404 VSS 0.385661f
C17994 VDD.t3313 VSS 0.034186f
C17995 VDD.t3312 VSS 0.080309f
C17996 VDD.t3510 VSS 0.080309f
C17997 VDD.n1405 VSS 0.385661f
C17998 VDD.t3511 VSS 0.034186f
C17999 VDD.n1406 VSS 0.327288f
C18000 VDD.n1407 VSS 0.327288f
C18001 VDD.t3147 VSS 0.034186f
C18002 VDD.n1408 VSS 0.298193f
C18003 VDD.n1409 VSS 0.298193f
C18004 VDD.t1511 VSS 0.025104f
C18005 VDD.n1410 VSS 0.016021f
C18006 VDD.n1411 VSS 0.282788f
C18007 VDD.n1412 VSS 0.144967f
C18008 VDD.n1413 VSS 0.304944f
C18009 VDD.n1414 VSS 3.12455f
C18010 VDD.t443 VSS 3.20156f
C18011 VDD.t438 VSS 7.734359f
C18012 VDD.t473 VSS 9.533179f
C18013 VDD.t881 VSS 7.54183f
C18014 VDD.n1415 VSS 3.4106f
C18015 VDD.n1416 VSS 0.304439f
C18016 VDD.n1417 VSS 0.064716f
C18017 VDD.n1418 VSS 0.096875f
C18018 VDD.t446 VSS 0.030289f
C18019 VDD.n1419 VSS 0.077802f
C18020 VDD.t460 VSS 0.008011f
C18021 VDD.t458 VSS 0.008011f
C18022 VDD.n1420 VSS 0.030319f
C18023 VDD.n1421 VSS 0.039264f
C18024 VDD.t444 VSS 0.008011f
C18025 VDD.t434 VSS 0.008011f
C18026 VDD.n1422 VSS 0.030367f
C18027 VDD.n1423 VSS 0.039375f
C18028 VDD.t447 VSS 0.030249f
C18029 VDD.n1424 VSS 0.077877f
C18030 VDD.n1425 VSS 0.017566f
C18031 VDD.n1426 VSS 0.063471f
C18032 VDD.n1427 VSS 0.304439f
C18033 VDD.n1428 VSS 3.4106f
C18034 VDD.n1429 VSS 3.4106f
C18035 VDD.n1430 VSS 0.303418f
C18036 VDD.n1431 VSS 0.063471f
C18037 VDD.n1432 VSS 0.234544f
C18038 VDD.t594 VSS 0.080308f
C18039 VDD.n1433 VSS 0.299675f
C18040 VDD.n1434 VSS 0.299675f
C18041 VDD.t984 VSS 0.080308f
C18042 VDD.n1435 VSS 0.299675f
C18043 VDD.n1436 VSS 0.299675f
C18044 VDD.t4010 VSS 0.080308f
C18045 VDD.n1437 VSS 0.299675f
C18046 VDD.n1438 VSS 0.299675f
C18047 VDD.t4136 VSS 0.080308f
C18048 VDD.n1439 VSS 0.299675f
C18049 VDD.n1440 VSS 0.241596f
C18050 VDD.t3074 VSS 0.082281f
C18051 VDD.t2748 VSS 0.042371f
C18052 VDD.t383 VSS 0.020844f
C18053 VDD.t3075 VSS 0.034186f
C18054 VDD.n1441 VSS 0.129126f
C18055 VDD.n1442 VSS 1.16761f
C18056 VDD.n1443 VSS 0.29513f
C18057 VDD.t4157 VSS 0.034186f
C18058 VDD.n1444 VSS 0.327288f
C18059 VDD.t4345 VSS 0.034186f
C18060 VDD.t4529 VSS 0.034186f
C18061 VDD.n1445 VSS 0.327288f
C18062 VDD.t4344 VSS 0.080309f
C18063 VDD.t4528 VSS 0.080309f
C18064 VDD.n1446 VSS 0.359117f
C18065 VDD.n1447 VSS 0.145214f
C18066 VDD.t387 VSS 0.19852f
C18067 VDD.n1448 VSS 0.440195f
C18068 VDD.n1449 VSS 0.137821f
C18069 VDD.n1450 VSS 0.261441f
C18070 VDD.t1934 VSS 0.025104f
C18071 VDD.n1451 VSS 0.016021f
C18072 VDD.n1452 VSS 0.289935f
C18073 VDD.n1453 VSS 0.016021f
C18074 VDD.t4315 VSS 0.016021f
C18075 VDD.n1454 VSS 0.016021f
C18076 VDD.n1455 VSS 0.282788f
C18077 VDD.n1456 VSS 0.016021f
C18078 VDD.t4739 VSS 0.025104f
C18079 VDD.n1457 VSS 0.298193f
C18080 VDD.n1458 VSS 0.298193f
C18081 VDD.t743 VSS 0.034186f
C18082 VDD.n1459 VSS 0.327288f
C18083 VDD.n1460 VSS 0.327288f
C18084 VDD.t2660 VSS 0.034186f
C18085 VDD.n1461 VSS 0.29513f
C18086 VDD.t820 VSS 0.080308f
C18087 VDD.t4215 VSS 0.034186f
C18088 VDD.t822 VSS 0.034186f
C18089 VDD.n1462 VSS 0.278056f
C18090 VDD.t3856 VSS 0.080308f
C18091 VDD.t3149 VSS 0.034186f
C18092 VDD.t3857 VSS 0.034186f
C18093 VDD.n1463 VSS 0.278056f
C18094 VDD.t4200 VSS 0.080308f
C18095 VDD.t3429 VSS 0.034186f
C18096 VDD.t4201 VSS 0.034186f
C18097 VDD.n1464 VSS 0.278056f
C18098 VDD.t4066 VSS 0.080308f
C18099 VDD.t3325 VSS 0.034186f
C18100 VDD.t4067 VSS 0.034186f
C18101 VDD.n1465 VSS 0.278056f
C18102 VDD.t4208 VSS 0.080308f
C18103 VDD.t3437 VSS 0.034186f
C18104 VDD.t4209 VSS 0.034186f
C18105 VDD.n1466 VSS 0.278056f
C18106 VDD.n1467 VSS 0.234544f
C18107 VDD.t3436 VSS 0.080308f
C18108 VDD.n1468 VSS 0.299675f
C18109 VDD.n1469 VSS 0.299675f
C18110 VDD.t3324 VSS 0.080308f
C18111 VDD.n1470 VSS 0.299675f
C18112 VDD.n1471 VSS 0.299675f
C18113 VDD.t3428 VSS 0.080308f
C18114 VDD.n1472 VSS 0.299675f
C18115 VDD.n1473 VSS 0.299675f
C18116 VDD.t3148 VSS 0.080308f
C18117 VDD.n1474 VSS 0.299675f
C18118 VDD.n1475 VSS 0.299675f
C18119 VDD.t4214 VSS 0.080308f
C18120 VDD.n1476 VSS 0.332862f
C18121 VDD.t4070 VSS 0.081403f
C18122 VDD.t3030 VSS 0.082281f
C18123 VDD.n1477 VSS 0.224389f
C18124 VDD.t2765 VSS 0.081403f
C18125 VDD.t1531 VSS 0.082281f
C18126 VDD.n1478 VSS 0.224389f
C18127 VDD.t379 VSS 0.020844f
C18128 VDD.t3031 VSS 0.034186f
C18129 VDD.n1479 VSS 0.129126f
C18130 VDD.n1480 VSS 1.50435f
C18131 VDD.n1481 VSS 0.29513f
C18132 VDD.t1772 VSS 0.034186f
C18133 VDD.n1482 VSS 0.327288f
C18134 VDD.n1483 VSS 0.327288f
C18135 VDD.t1930 VSS 0.034186f
C18136 VDD.n1484 VSS 0.298193f
C18137 VDD.n1485 VSS 0.298193f
C18138 VDD.t1684 VSS 0.025104f
C18139 VDD.n1486 VSS 0.016021f
C18140 VDD.n1487 VSS 0.289935f
C18141 VDD.n1488 VSS 0.016021f
C18142 VDD.t1682 VSS 0.016021f
C18143 VDD.n1489 VSS 0.016021f
C18144 VDD.n1490 VSS 0.282788f
C18145 VDD.n1491 VSS 0.016021f
C18146 VDD.t739 VSS 0.025104f
C18147 VDD.n1492 VSS 0.298193f
C18148 VDD.n1493 VSS 0.298193f
C18149 VDD.t4639 VSS 0.034186f
C18150 VDD.n1494 VSS 0.327288f
C18151 VDD.n1495 VSS 0.327288f
C18152 VDD.t2409 VSS 0.034186f
C18153 VDD.n1496 VSS 0.29513f
C18154 VDD.t1311 VSS 0.034186f
C18155 VDD.t1310 VSS 0.080309f
C18156 VDD.t1523 VSS 0.080309f
C18157 VDD.n1497 VSS 0.385661f
C18158 VDD.t3221 VSS 0.034186f
C18159 VDD.t3220 VSS 0.080309f
C18160 VDD.t3395 VSS 0.080309f
C18161 VDD.n1498 VSS 0.385661f
C18162 VDD.t4697 VSS 0.025104f
C18163 VDD.t4696 VSS 0.080309f
C18164 VDD.t785 VSS 0.080309f
C18165 VDD.n1499 VSS 0.385661f
C18166 VDD.t3728 VSS 0.016021f
C18167 VDD.n1500 VSS 0.016021f
C18168 VDD.t3523 VSS 0.016021f
C18169 VDD.n1501 VSS 0.016021f
C18170 VDD.t1942 VSS 0.080309f
C18171 VDD.t2188 VSS 0.080309f
C18172 VDD.n1502 VSS 0.385661f
C18173 VDD.t1943 VSS 0.025104f
C18174 VDD.t3507 VSS 0.034186f
C18175 VDD.t3506 VSS 0.080309f
C18176 VDD.t3707 VSS 0.080309f
C18177 VDD.n1503 VSS 0.385661f
C18178 VDD.t3925 VSS 0.034186f
C18179 VDD.t3924 VSS 0.080309f
C18180 VDD.t4150 VSS 0.080309f
C18181 VDD.n1504 VSS 0.29378f
C18182 VDD.t2756 VSS 0.034186f
C18183 VDD.n1505 VSS 0.136328f
C18184 VDD.t307 VSS 0.019806f
C18185 VDD.t3785 VSS 0.035116f
C18186 VDD.n1506 VSS 0.087326f
C18187 VDD.n1507 VSS 0.15353f
C18188 VDD.t3643 VSS 0.034186f
C18189 VDD.n1508 VSS 0.136328f
C18190 VDD.t579 VSS 0.034186f
C18191 VDD.n1509 VSS 0.136328f
C18192 VDD.t3874 VSS 0.231787f
C18193 VDD.n1510 VSS 0.227269f
C18194 VDD.t3875 VSS 0.034186f
C18195 VDD.t4429 VSS 0.034186f
C18196 VDD.t1666 VSS 0.231805f
C18197 VDD.n1511 VSS 0.451142f
C18198 VDD.t4207 VSS 0.025104f
C18199 VDD.n1512 VSS 0.02945f
C18200 VDD.t694 VSS 0.231805f
C18201 VDD.n1513 VSS 0.451142f
C18202 VDD.t2432 VSS 0.025104f
C18203 VDD.t2431 VSS 0.231805f
C18204 VDD.n1514 VSS 0.451142f
C18205 VDD.n1515 VSS 0.29843f
C18206 VDD.n1516 VSS 0.016021f
C18207 VDD.t696 VSS 0.025104f
C18208 VDD.n1517 VSS 0.186367f
C18209 VDD.n1518 VSS 0.185495f
C18210 VDD.t1080 VSS 0.034186f
C18211 VDD.n1519 VSS 0.23881f
C18212 VDD.n1520 VSS 0.060699f
C18213 VDD.n1521 VSS 1.52188f
C18214 VDD.t3061 VSS 0.034186f
C18215 VDD.n1522 VSS 0.249436f
C18216 VDD.t3017 VSS 0.034186f
C18217 VDD.n1523 VSS 0.179934f
C18218 VDD.t1625 VSS 0.231805f
C18219 VDD.n1524 VSS 0.451142f
C18220 VDD.t1872 VSS 0.025104f
C18221 VDD.t1871 VSS 0.231805f
C18222 VDD.n1525 VSS 0.451142f
C18223 VDD.n1526 VSS 0.29843f
C18224 VDD.n1527 VSS 0.016021f
C18225 VDD.t1626 VSS 0.025104f
C18226 VDD.n1528 VSS 0.238069f
C18227 VDD.n1529 VSS 0.563325f
C18228 VDD.t3016 VSS 0.233178f
C18229 VDD.n1530 VSS 0.381077f
C18230 VDD.n1531 VSS 0.381077f
C18231 VDD.t3060 VSS 0.231787f
C18232 VDD.n1532 VSS 0.33592f
C18233 VDD.n1533 VSS 0.320606f
C18234 VDD.t3604 VSS 0.034186f
C18235 VDD.t3445 VSS 0.034186f
C18236 VDD.n1534 VSS 0.249436f
C18237 VDD.t2303 VSS 0.034186f
C18238 VDD.n1535 VSS 0.180326f
C18239 VDD.t996 VSS 0.231805f
C18240 VDD.n1536 VSS 0.451142f
C18241 VDD.t1192 VSS 0.025104f
C18242 VDD.n1537 VSS 0.185495f
C18243 VDD.t1190 VSS 0.231805f
C18244 VDD.n1538 VSS 0.451142f
C18245 VDD.n1539 VSS 0.29843f
C18246 VDD.n1540 VSS 0.016021f
C18247 VDD.t998 VSS 0.025104f
C18248 VDD.n1541 VSS 0.238069f
C18249 VDD.n1542 VSS 0.562943f
C18250 VDD.t2301 VSS 0.233168f
C18251 VDD.n1543 VSS 0.381077f
C18252 VDD.n1544 VSS 0.381077f
C18253 VDD.t3444 VSS 0.231787f
C18254 VDD.n1545 VSS 0.33592f
C18255 VDD.t3603 VSS 0.231787f
C18256 VDD.n1546 VSS 0.33592f
C18257 VDD.n1547 VSS 0.147735f
C18258 VDD.n1548 VSS 0.117015f
C18259 VDD.n1549 VSS 1.52159f
C18260 VDD.t923 VSS 3.32223f
C18261 VDD.t1667 VSS 3.93704f
C18262 VDD.t695 VSS 2.74191f
C18263 VDD.n1550 VSS 0.269232f
C18264 VDD.t2302 VSS 3.32223f
C18265 VDD.t997 VSS 3.93704f
C18266 VDD.t1191 VSS 2.7319f
C18267 VDD.n1551 VSS 2.04987f
C18268 VDD.n1552 VSS 0.266386f
C18269 VDD.n1553 VSS 0.02945f
C18270 VDD.n1554 VSS 0.091202f
C18271 VDD.t4776 VSS 0.017093f
C18272 VDD.t4779 VSS 0.017093f
C18273 VDD.n1555 VSS 0.155393f
C18274 VDD.t4778 VSS 0.017093f
C18275 VDD.t4781 VSS 0.017093f
C18276 VDD.n1556 VSS 0.173624f
C18277 VDD.t4777 VSS 0.017093f
C18278 VDD.t4780 VSS 0.017093f
C18279 VDD.n1557 VSS 0.155393f
C18280 VDD.n1558 VSS 0.091202f
C18281 VDD.n1559 VSS 0.186367f
C18282 VDD.t4206 VSS 0.231805f
C18283 VDD.n1560 VSS 0.451142f
C18284 VDD.n1561 VSS 0.29843f
C18285 VDD.n1562 VSS 0.016021f
C18286 VDD.t1668 VSS 0.025104f
C18287 VDD.n1563 VSS 0.238069f
C18288 VDD.n1564 VSS 0.329848f
C18289 VDD.n1565 VSS 0.118255f
C18290 VDD.n1566 VSS 0.26663f
C18291 VDD.n1567 VSS 0.275158f
C18292 VDD.t4428 VSS 0.080308f
C18293 VDD.n1568 VSS 0.337025f
C18294 VDD.n1569 VSS 0.255139f
C18295 VDD.t577 VSS 0.080308f
C18296 VDD.n1570 VSS 0.147087f
C18297 VDD.n1571 VSS 0.147087f
C18298 VDD.t3642 VSS 0.080308f
C18299 VDD.n1572 VSS 0.147087f
C18300 VDD.n1573 VSS 0.118683f
C18301 VDD.t3784 VSS 0.080308f
C18302 VDD.n1574 VSS 0.118683f
C18303 VDD.n1575 VSS 0.147087f
C18304 VDD.t2755 VSS 0.080308f
C18305 VDD.n1576 VSS 0.163319f
C18306 VDD.t2465 VSS 0.034186f
C18307 VDD.n1577 VSS 0.136328f
C18308 VDD.t1240 VSS 0.034186f
C18309 VDD.n1578 VSS 0.136328f
C18310 VDD.t1570 VSS 0.034186f
C18311 VDD.n1579 VSS 0.136328f
C18312 VDD.t1448 VSS 0.034186f
C18313 VDD.n1580 VSS 0.136328f
C18314 VDD.t1581 VSS 0.034186f
C18315 VDD.n1581 VSS 0.136328f
C18316 VDD.n1582 VSS 0.115234f
C18317 VDD.t1580 VSS 0.080308f
C18318 VDD.n1583 VSS 0.147087f
C18319 VDD.n1584 VSS 0.147087f
C18320 VDD.t1447 VSS 0.080308f
C18321 VDD.n1585 VSS 0.147087f
C18322 VDD.n1586 VSS 0.147087f
C18323 VDD.t1569 VSS 0.080308f
C18324 VDD.n1587 VSS 0.147087f
C18325 VDD.n1588 VSS 0.147087f
C18326 VDD.t1239 VSS 0.080308f
C18327 VDD.n1589 VSS 0.147087f
C18328 VDD.n1590 VSS 0.147087f
C18329 VDD.t2464 VSS 0.080308f
C18330 VDD.n1591 VSS 0.163319f
C18331 VDD.n1592 VSS 0.302817f
C18332 VDD.n1593 VSS 0.357405f
C18333 VDD.t4151 VSS 0.034186f
C18334 VDD.n1594 VSS 0.327288f
C18335 VDD.n1595 VSS 0.327288f
C18336 VDD.t3708 VSS 0.034186f
C18337 VDD.n1596 VSS 0.298193f
C18338 VDD.n1597 VSS 0.298193f
C18339 VDD.t2189 VSS 0.025104f
C18340 VDD.n1598 VSS 0.016021f
C18341 VDD.n1599 VSS 0.282788f
C18342 VDD.n1600 VSS 0.144967f
C18343 VDD.t3522 VSS 0.080309f
C18344 VDD.t3727 VSS 0.080309f
C18345 VDD.n1601 VSS 0.24784f
C18346 VDD.n1602 VSS 0.289935f
C18347 VDD.n1603 VSS 0.016021f
C18348 VDD.t786 VSS 0.025104f
C18349 VDD.n1604 VSS 0.298193f
C18350 VDD.n1605 VSS 0.298193f
C18351 VDD.t3396 VSS 0.034186f
C18352 VDD.n1606 VSS 0.327288f
C18353 VDD.n1607 VSS 0.327288f
C18354 VDD.t1524 VSS 0.034186f
C18355 VDD.n1608 VSS 0.29513f
C18356 VDD.t2801 VSS 0.082281f
C18357 VDD.n1609 VSS 0.224389f
C18358 VDD.n1610 VSS 1.50435f
C18359 VDD.t4124 VSS 0.082281f
C18360 VDD.n1611 VSS 0.224389f
C18361 VDD.t1069 VSS 0.081403f
C18362 VDD.n1612 VSS 0.241596f
C18363 VDD.n1613 VSS 0.299675f
C18364 VDD.t960 VSS 0.080308f
C18365 VDD.n1614 VSS 0.299675f
C18366 VDD.n1615 VSS 0.299675f
C18367 VDD.t2072 VSS 0.080308f
C18368 VDD.n1616 VSS 0.299675f
C18369 VDD.n1617 VSS 0.299675f
C18370 VDD.t1697 VSS 0.080308f
C18371 VDD.n1618 VSS 0.234959f
C18372 VDD.n1619 VSS 0.096875f
C18373 VDD.t360 VSS 0.030289f
C18374 VDD.n1620 VSS 0.077802f
C18375 VDD.t337 VSS 0.008011f
C18376 VDD.t338 VSS 0.008011f
C18377 VDD.n1621 VSS 0.030319f
C18378 VDD.n1622 VSS 0.039264f
C18379 VDD.t354 VSS 0.008011f
C18380 VDD.t349 VSS 0.008011f
C18381 VDD.n1623 VSS 0.030367f
C18382 VDD.n1624 VSS 0.039375f
C18383 VDD.t327 VSS 0.030249f
C18384 VDD.n1625 VSS 0.077873f
C18385 VDD.n1626 VSS 0.145738f
C18386 VDD.n1627 VSS 0.131514f
C18387 VDD.t1389 VSS 0.080308f
C18388 VDD.n1628 VSS 0.297077f
C18389 VDD.n1629 VSS 0.32759f
C18390 VDD.t922 VSS 0.231787f
C18391 VDD.n1630 VSS 0.336864f
C18392 VDD.t1258 VSS 0.080308f
C18393 VDD.n1631 VSS 0.329955f
C18394 VDD.n1632 VSS 0.32759f
C18395 VDD.t1079 VSS 0.231787f
C18396 VDD.n1633 VSS 0.336864f
C18397 VDD.t2483 VSS 0.080308f
C18398 VDD.n1634 VSS 0.329955f
C18399 VDD.n1635 VSS 0.32759f
C18400 VDD.t4588 VSS 0.231787f
C18401 VDD.n1636 VSS 0.336864f
C18402 VDD.n1637 VSS 0.299606f
C18403 VDD.t2325 VSS 0.080308f
C18404 VDD.n1638 VSS 0.275158f
C18405 VDD.n1639 VSS 0.244711f
C18406 VDD.n1640 VSS 0.214352f
C18407 VDD.n1641 VSS 0.17315f
C18408 VDD.t3409 VSS 0.080308f
C18409 VDD.n1642 VSS 0.158502f
C18410 VDD.n1643 VSS 0.295034f
C18411 VDD.t2937 VSS 0.035031f
C18412 VDD.n1644 VSS 0.141721f
C18413 VDD.n1645 VSS 0.141721f
C18414 VDD.t2140 VSS 0.034186f
C18415 VDD.n1646 VSS 0.129218f
C18416 VDD.n1647 VSS 0.129218f
C18417 VDD.t3343 VSS 0.025104f
C18418 VDD.n1648 VSS 0.016021f
C18419 VDD.n1649 VSS 0.121516f
C18420 VDD.n1650 VSS 0.062293f
C18421 VDD.n1651 VSS 0.304763f
C18422 VDD.n1652 VSS 3.12455f
C18423 VDD.n1653 VSS 0.304944f
C18424 VDD.n1654 VSS 0.062293f
C18425 VDD.n1655 VSS 0.121516f
C18426 VDD.n1656 VSS 0.016021f
C18427 VDD.t1092 VSS 0.025104f
C18428 VDD.n1657 VSS 0.129218f
C18429 VDD.n1658 VSS 0.129218f
C18430 VDD.t2711 VSS 0.034186f
C18431 VDD.n1659 VSS 0.141721f
C18432 VDD.n1660 VSS 0.141721f
C18433 VDD.t3119 VSS 0.035031f
C18434 VDD.n1661 VSS 0.295034f
C18435 VDD.n1662 VSS 0.163319f
C18436 VDD.t4552 VSS 0.080308f
C18437 VDD.n1663 VSS 0.147087f
C18438 VDD.n1664 VSS 0.118683f
C18439 VDD.t1521 VSS 0.080308f
C18440 VDD.n1665 VSS 0.118683f
C18441 VDD.n1666 VSS 0.147087f
C18442 VDD.t3632 VSS 0.080308f
C18443 VDD.n1667 VSS 0.147087f
C18444 VDD.n1668 VSS 0.147087f
C18445 VDD.t4744 VSS 0.080308f
C18446 VDD.n1669 VSS 0.147087f
C18447 VDD.n1670 VSS 0.147087f
C18448 VDD.t4620 VSS 0.080308f
C18449 VDD.n1671 VSS 0.115436f
C18450 VDD.n1672 VSS 0.047764f
C18451 VDD.t348 VSS 0.030249f
C18452 VDD.n1673 VSS 0.077873f
C18453 VDD.n1674 VSS 0.039375f
C18454 VDD.t345 VSS 0.008011f
C18455 VDD.t361 VSS 0.008011f
C18456 VDD.n1675 VSS 0.030319f
C18457 VDD.n1676 VSS 0.039264f
C18458 VDD.t343 VSS 0.030289f
C18459 VDD.n1677 VSS 0.077802f
C18460 VDD.n1678 VSS 0.096875f
C18461 VDD.t364 VSS 0.030249f
C18462 VDD.n1679 VSS 0.077873f
C18463 VDD.n1680 VSS 0.039375f
C18464 VDD.t344 VSS 0.008011f
C18465 VDD.t377 VSS 0.008011f
C18466 VDD.n1681 VSS 0.030319f
C18467 VDD.n1682 VSS 0.039264f
C18468 VDD.t333 VSS 0.030289f
C18469 VDD.n1683 VSS 0.077802f
C18470 VDD.n1684 VSS 0.096875f
C18471 VDD.t359 VSS 0.030249f
C18472 VDD.n1685 VSS 0.077873f
C18473 VDD.n1686 VSS 0.039375f
C18474 VDD.t355 VSS 0.008011f
C18475 VDD.t4984 VSS 0.008011f
C18476 VDD.n1687 VSS 0.030319f
C18477 VDD.n1688 VSS 0.039264f
C18478 VDD.t363 VSS 0.030289f
C18479 VDD.n1689 VSS 0.077802f
C18480 VDD.n1690 VSS 0.017494f
C18481 VDD.n1691 VSS 0.017569f
C18482 VDD.t450 VSS 0.030249f
C18483 VDD.n1692 VSS 0.077873f
C18484 VDD.n1693 VSS 0.039375f
C18485 VDD.t452 VSS 0.008011f
C18486 VDD.t466 VSS 0.008011f
C18487 VDD.n1694 VSS 0.030319f
C18488 VDD.n1695 VSS 0.039264f
C18489 VDD.t439 VSS 0.030289f
C18490 VDD.n1696 VSS 0.077802f
C18491 VDD.n1697 VSS 0.096875f
C18492 VDD.n1698 VSS 0.234959f
C18493 VDD.t1327 VSS 0.080308f
C18494 VDD.n1699 VSS 0.299675f
C18495 VDD.n1700 VSS 0.299675f
C18496 VDD.t1214 VSS 0.080308f
C18497 VDD.n1701 VSS 0.299675f
C18498 VDD.n1702 VSS 0.299675f
C18499 VDD.t1322 VSS 0.080308f
C18500 VDD.n1703 VSS 0.299675f
C18501 VDD.n1704 VSS 0.299675f
C18502 VDD.t1028 VSS 0.080308f
C18503 VDD.n1705 VSS 0.299675f
C18504 VDD.n1706 VSS 0.299675f
C18505 VDD.t2148 VSS 0.080308f
C18506 VDD.n1707 VSS 0.332862f
C18507 VDD.n1708 VSS 0.592265f
C18508 VDD.n1709 VSS 0.29513f
C18509 VDD.t3297 VSS 0.034186f
C18510 VDD.n1710 VSS 0.327288f
C18511 VDD.n1711 VSS 0.327288f
C18512 VDD.t2913 VSS 0.034186f
C18513 VDD.n1712 VSS 0.298193f
C18514 VDD.n1713 VSS 0.298193f
C18515 VDD.t3137 VSS 0.025104f
C18516 VDD.n1714 VSS 0.016021f
C18517 VDD.n1715 VSS 0.282788f
C18518 VDD.n1716 VSS 0.144967f
C18519 VDD.n1717 VSS 0.304944f
C18520 VDD.n1718 VSS 3.12105f
C18521 VDD.t441 VSS 3.18057f
C18522 VDD.t424 VSS 7.734359f
C18523 VDD.t467 VSS 9.533179f
C18524 VDD.t692 VSS 7.54183f
C18525 VDD.n1719 VSS 3.4106f
C18526 VDD.n1720 VSS 0.304439f
C18527 VDD.n1721 VSS 0.064716f
C18528 VDD.n1722 VSS 0.234544f
C18529 VDD.t1142 VSS 0.080308f
C18530 VDD.n1723 VSS 0.299675f
C18531 VDD.n1724 VSS 0.299675f
C18532 VDD.t1459 VSS 0.080308f
C18533 VDD.n1725 VSS 0.299675f
C18534 VDD.n1726 VSS 0.299675f
C18535 VDD.t4502 VSS 0.080308f
C18536 VDD.n1727 VSS 0.299675f
C18537 VDD.n1728 VSS 0.299675f
C18538 VDD.t4636 VSS 0.080308f
C18539 VDD.n1729 VSS 0.299675f
C18540 VDD.n1730 VSS 0.299675f
C18541 VDD.t3536 VSS 0.080308f
C18542 VDD.n1731 VSS 0.332862f
C18543 VDD.n1732 VSS 0.592265f
C18544 VDD.n1733 VSS 0.29513f
C18545 VDD.t1785 VSS 0.034186f
C18546 VDD.n1734 VSS 0.327288f
C18547 VDD.n1735 VSS 0.327288f
C18548 VDD.t1371 VSS 0.034186f
C18549 VDD.n1736 VSS 0.234091f
C18550 VDD.n1737 VSS 0.298193f
C18551 VDD.t1506 VSS 0.025104f
C18552 VDD.n1738 VSS 0.016021f
C18553 VDD.n1739 VSS 0.282788f
C18554 VDD.n1740 VSS 0.144967f
C18555 VDD.n1741 VSS 0.304944f
C18556 VDD.n1742 VSS 3.12455f
C18557 VDD.n1743 VSS 0.304944f
C18558 VDD.n1744 VSS 0.062293f
C18559 VDD.t4640 VSS 0.080309f
C18560 VDD.n1745 VSS 0.113227f
C18561 VDD.n1746 VSS 0.124587f
C18562 VDD.n1747 VSS 0.016021f
C18563 VDD.t741 VSS 0.025104f
C18564 VDD.n1748 VSS 0.129218f
C18565 VDD.n1749 VSS 0.129218f
C18566 VDD.t3051 VSS 0.034186f
C18567 VDD.n1750 VSS 0.133386f
C18568 VDD.n1751 VSS 0.789016f
C18569 VDD.t1171 VSS 0.080666f
C18570 VDD.n1752 VSS 0.445309f
C18571 VDD.n1754 VSS 0.018625f
C18572 VDD.n1755 VSS 0.01502f
C18573 VDD.n1756 VSS 0.191469f
C18574 VDD.n1757 VSS 0.01487f
C18575 VDD.n1759 VSS 0.018249f
C18576 VDD.n1760 VSS 0.009312f
C18577 VDD.n1761 VSS 2.45645f
C18578 VDD.n1762 VSS 1.92254f
C18579 VDD.n1763 VSS 0.43261f
C18580 VDD.n1764 VSS 0.009688f
C18581 VDD.t1672 VSS 0.028519f
C18582 VDD.t3127 VSS 0.028519f
C18583 VDD.n1765 VSS 0.009191f
C18584 VDD.n1766 VSS 0.113124f
C18585 VDD.n1767 VSS 0.012131f
C18586 VDD.n1768 VSS 0.269046f
C18587 VDD.t3591 VSS 0.066856f
C18588 VDD.n1769 VSS 0.125227f
C18589 VDD.t1244 VSS 0.025104f
C18590 VDD.n1770 VSS 0.083673f
C18591 VDD.n1771 VSS 1.05032f
C18592 VDD.n1772 VSS 0.207221f
C18593 VDD.t968 VSS 1.45905f
C18594 VDD.t1102 VSS 1.96535f
C18595 VDD.t376 VSS 1.96535f
C18596 VDD.t373 VSS 1.36988f
C18597 VDD.t374 VSS 1.31955f
C18598 VDD.t584 VSS 0.066856f
C18599 VDD.n1773 VSS 0.14405f
C18600 VDD.t3947 VSS 0.025104f
C18601 VDD.n1774 VSS 0.116823f
C18602 VDD.t3946 VSS 0.066856f
C18603 VDD.n1775 VSS 0.14405f
C18604 VDD.n1776 VSS 0.120118f
C18605 VDD.n1777 VSS 0.016021f
C18606 VDD.t585 VSS 0.025104f
C18607 VDD.n1778 VSS 0.105404f
C18608 VDD.t2615 VSS 0.066856f
C18609 VDD.n1779 VSS 0.14405f
C18610 VDD.t3694 VSS 0.025104f
C18611 VDD.n1780 VSS 0.04911f
C18612 VDD.t4307 VSS 0.028519f
C18613 VDD.t4703 VSS 0.028519f
C18614 VDD.n1781 VSS 0.009191f
C18615 VDD.t2837 VSS 0.028519f
C18616 VDD.t4561 VSS 0.028519f
C18617 VDD.n1782 VSS 0.009191f
C18618 VDD.n1783 VSS 0.523473f
C18619 VDD.n1784 VSS 0.206947f
C18620 VDD.n1785 VSS 0.208771f
C18621 VDD.t375 VSS 1.96535f
C18622 VDD.t1422 VSS 1.96535f
C18623 VDD.t1644 VSS 1.45794f
C18624 VDD.n1786 VSS 0.865258f
C18625 VDD.n1787 VSS 0.865258f
C18626 VDD.t3779 VSS 0.028519f
C18627 VDD.t2489 VSS 0.028519f
C18628 VDD.n1788 VSS 0.009191f
C18629 VDD.t2237 VSS 0.028519f
C18630 VDD.t4057 VSS 0.028519f
C18631 VDD.n1789 VSS 0.009191f
C18632 VDD.n1790 VSS 0.523473f
C18633 VDD.t1194 VSS 0.028519f
C18634 VDD.t4003 VSS 0.028519f
C18635 VDD.n1791 VSS 0.009191f
C18636 VDD.t3811 VSS 0.028519f
C18637 VDD.t1474 VSS 0.028519f
C18638 VDD.n1792 VSS 0.009191f
C18639 VDD.n1793 VSS 0.471397f
C18640 VDD.n1794 VSS 0.206947f
C18641 VDD.n1795 VSS 0.207221f
C18642 VDD.t2692 VSS 0.066856f
C18643 VDD.n1796 VSS 0.14405f
C18644 VDD.t2889 VSS 0.025104f
C18645 VDD.t1193 VSS 0.066856f
C18646 VDD.t3810 VSS 0.066856f
C18647 VDD.t1473 VSS 0.066856f
C18648 VDD.t4002 VSS 0.066856f
C18649 VDD.n1797 VSS 0.690489f
C18650 VDD.t854 VSS 0.066856f
C18651 VDD.t3450 VSS 0.066856f
C18652 VDD.t1114 VSS 0.066856f
C18653 VDD.t3620 VSS 0.066856f
C18654 VDD.n1798 VSS 0.690489f
C18655 VDD.t856 VSS 0.028519f
C18656 VDD.t3621 VSS 0.028519f
C18657 VDD.n1799 VSS 0.009191f
C18658 VDD.t3451 VSS 0.028519f
C18659 VDD.t1116 VSS 0.028519f
C18660 VDD.n1800 VSS 0.009191f
C18661 VDD.n1801 VSS 0.644755f
C18662 VDD.t2886 VSS 0.066856f
C18663 VDD.t2233 VSS 0.066856f
C18664 VDD.t3114 VSS 0.066856f
C18665 VDD.t4034 VSS 0.066856f
C18666 VDD.n1802 VSS 0.709674f
C18667 VDD.t2887 VSS 0.028519f
C18668 VDD.t4035 VSS 0.028519f
C18669 VDD.n1803 VSS 0.009191f
C18670 VDD.t2235 VSS 0.028519f
C18671 VDD.t3115 VSS 0.028519f
C18672 VDD.n1804 VSS 0.009191f
C18673 VDD.n1805 VSS 0.309003f
C18674 VDD.t4452 VSS 0.066856f
C18675 VDD.n1806 VSS 0.14405f
C18676 VDD.t3317 VSS 0.025104f
C18677 VDD.t1359 VSS 0.066856f
C18678 VDD.n1807 VSS 0.14405f
C18679 VDD.t1556 VSS 0.025104f
C18680 VDD.n1808 VSS 0.033925f
C18681 VDD.t417 VSS 0.019767f
C18682 VDD.t295 VSS 0.018805f
C18683 VDD.n1809 VSS 0.054793f
C18684 VDD.t294 VSS 0.018792f
C18685 VDD.t416 VSS 0.019781f
C18686 VDD.n1810 VSS 0.077486f
C18687 VDD.n1811 VSS 0.252514f
C18688 VDD.n1812 VSS 0.199549f
C18689 VDD.n1813 VSS 0.060108f
C18690 VDD.t1555 VSS 0.066856f
C18691 VDD.n1814 VSS 0.131361f
C18692 VDD.n1815 VSS 0.120118f
C18693 VDD.n1816 VSS 0.016021f
C18694 VDD.t1360 VSS 0.025104f
C18695 VDD.n1817 VSS 0.105404f
C18696 VDD.n1818 VSS 0.057098f
C18697 VDD.n1819 VSS 0.087217f
C18698 VDD.t3316 VSS 0.066856f
C18699 VDD.n1820 VSS 0.14405f
C18700 VDD.n1821 VSS 0.120118f
C18701 VDD.n1822 VSS 0.016021f
C18702 VDD.t4453 VSS 0.025104f
C18703 VDD.n1823 VSS 0.116823f
C18704 VDD.n1824 VSS 0.77922f
C18705 VDD.n1825 VSS 0.116823f
C18706 VDD.t2888 VSS 0.066856f
C18707 VDD.n1826 VSS 0.14405f
C18708 VDD.n1827 VSS 0.120118f
C18709 VDD.n1828 VSS 0.016021f
C18710 VDD.t2693 VSS 0.025104f
C18711 VDD.n1829 VSS 0.105404f
C18712 VDD.n1830 VSS 0.057098f
C18713 VDD.t855 VSS 1.45794f
C18714 VDD.t2488 VSS 1.96535f
C18715 VDD.t324 VSS 1.96535f
C18716 VDD.t325 VSS 1.36988f
C18717 VDD.n1831 VSS 0.645798f
C18718 VDD.t792 VSS 1.45794f
C18719 VDD.n1832 VSS 0.206947f
C18720 VDD.n1833 VSS 0.208771f
C18721 VDD.t3353 VSS 0.028519f
C18722 VDD.t1970 VSS 0.028519f
C18723 VDD.n1834 VSS 0.009191f
C18724 VDD.t3169 VSS 0.028519f
C18725 VDD.t3013 VSS 0.028519f
C18726 VDD.n1835 VSS 0.009191f
C18727 VDD.n1836 VSS 0.528101f
C18728 VDD.t793 VSS 0.028519f
C18729 VDD.t3567 VSS 0.028519f
C18730 VDD.n1837 VSS 0.009191f
C18731 VDD.t791 VSS 0.066856f
C18732 VDD.t4698 VSS 0.066856f
C18733 VDD.t4530 VSS 0.066856f
C18734 VDD.t4326 VSS 0.066856f
C18735 VDD.t4531 VSS 0.028519f
C18736 VDD.t3247 VSS 0.028519f
C18737 VDD.n1838 VSS 0.009191f
C18738 VDD.t3844 VSS 0.066856f
C18739 VDD.t3140 VSS 0.066856f
C18740 VDD.t3845 VSS 0.028519f
C18741 VDD.t921 VSS 0.028519f
C18742 VDD.n1839 VSS 0.009191f
C18743 VDD.t2520 VSS 0.066856f
C18744 VDD.n1840 VSS 0.14405f
C18745 VDD.t3629 VSS 0.025104f
C18746 VDD.t1331 VSS 0.066856f
C18747 VDD.n1841 VSS 0.14405f
C18748 VDD.t1139 VSS 0.025104f
C18749 VDD.n1842 VSS 0.04911f
C18750 VDD.t1033 VSS 0.028519f
C18751 VDD.t3805 VSS 0.028519f
C18752 VDD.n1843 VSS 0.009191f
C18753 VDD.t2780 VSS 0.028519f
C18754 VDD.t1285 VSS 0.028519f
C18755 VDD.n1844 VSS 0.009191f
C18756 VDD.n1845 VSS 0.523473f
C18757 VDD.n1846 VSS 0.207221f
C18758 VDD.n1847 VSS 0.206947f
C18759 VDD.n1848 VSS 0.208771f
C18760 VDD.t920 VSS 1.96535f
C18761 VDD.t503 VSS 1.96535f
C18762 VDD.t502 VSS 1.36988f
C18763 VDD.n1849 VSS 0.645798f
C18764 VDD.n1850 VSS 0.595476f
C18765 VDD.t501 VSS 1.31955f
C18766 VDD.t500 VSS 1.96535f
C18767 VDD.t2779 VSS 1.96535f
C18768 VDD.t1145 VSS 1.45794f
C18769 VDD.n1851 VSS 0.865258f
C18770 VDD.n1852 VSS 0.865258f
C18771 VDD.t4629 VSS 0.028519f
C18772 VDD.t3738 VSS 0.028519f
C18773 VDD.n1853 VSS 0.009191f
C18774 VDD.t2157 VSS 0.028519f
C18775 VDD.t784 VSS 0.028519f
C18776 VDD.n1854 VSS 0.009191f
C18777 VDD.n1855 VSS 0.523473f
C18778 VDD.t2096 VSS 0.028519f
C18779 VDD.t1161 VSS 0.028519f
C18780 VDD.n1856 VSS 0.009191f
C18781 VDD.t3744 VSS 0.028519f
C18782 VDD.t2446 VSS 0.028519f
C18783 VDD.n1857 VSS 0.009191f
C18784 VDD.n1858 VSS 0.471397f
C18785 VDD.n1859 VSS 0.206947f
C18786 VDD.n1860 VSS 0.207221f
C18787 VDD.t1444 VSS 0.066856f
C18788 VDD.n1861 VSS 0.14405f
C18789 VDD.t4403 VSS 0.025104f
C18790 VDD.t1901 VSS 0.066856f
C18791 VDD.n1862 VSS 0.14405f
C18792 VDD.t2120 VSS 0.025104f
C18793 VDD.t705 VSS 0.066856f
C18794 VDD.n1863 VSS 0.14405f
C18795 VDD.t3655 VSS 0.025104f
C18796 VDD.n1864 VSS 0.033925f
C18797 VDD.t4770 VSS 0.019767f
C18798 VDD.t4768 VSS 0.018805f
C18799 VDD.n1865 VSS 0.054793f
C18800 VDD.t4771 VSS 0.018792f
C18801 VDD.t4769 VSS 0.019781f
C18802 VDD.n1866 VSS 0.077486f
C18803 VDD.n1867 VSS 0.252514f
C18804 VDD.n1868 VSS 0.199549f
C18805 VDD.n1869 VSS 0.060108f
C18806 VDD.t3654 VSS 0.066856f
C18807 VDD.n1870 VSS 0.131361f
C18808 VDD.n1871 VSS 0.120118f
C18809 VDD.n1872 VSS 0.016021f
C18810 VDD.t706 VSS 0.025104f
C18811 VDD.n1873 VSS 0.105404f
C18812 VDD.n1874 VSS 0.057098f
C18813 VDD.n1875 VSS 0.087217f
C18814 VDD.t2119 VSS 0.066856f
C18815 VDD.n1876 VSS 0.14405f
C18816 VDD.n1877 VSS 0.120118f
C18817 VDD.n1878 VSS 0.016021f
C18818 VDD.t1902 VSS 0.025104f
C18819 VDD.n1879 VSS 0.116823f
C18820 VDD.t2095 VSS 0.066856f
C18821 VDD.t3743 VSS 0.066856f
C18822 VDD.t2445 VSS 0.066856f
C18823 VDD.t1160 VSS 0.066856f
C18824 VDD.n1880 VSS 0.690489f
C18825 VDD.t1687 VSS 0.066856f
C18826 VDD.t3375 VSS 0.066856f
C18827 VDD.t1983 VSS 0.066856f
C18828 VDD.t803 VSS 0.066856f
C18829 VDD.n1881 VSS 0.690489f
C18830 VDD.t1688 VSS 0.028519f
C18831 VDD.t805 VSS 0.028519f
C18832 VDD.n1882 VSS 0.009191f
C18833 VDD.t3376 VSS 0.028519f
C18834 VDD.t1984 VSS 0.028519f
C18835 VDD.n1883 VSS 0.009191f
C18836 VDD.n1884 VSS 0.644755f
C18837 VDD.t1659 VSS 0.066856f
C18838 VDD.t699 VSS 0.066856f
C18839 VDD.t1903 VSS 0.066856f
C18840 VDD.t1439 VSS 0.066856f
C18841 VDD.n1885 VSS 0.709674f
C18842 VDD.t1661 VSS 0.028519f
C18843 VDD.t1440 VSS 0.028519f
C18844 VDD.n1886 VSS 0.009191f
C18845 VDD.t701 VSS 0.028519f
C18846 VDD.t1904 VSS 0.028519f
C18847 VDD.n1887 VSS 0.009191f
C18848 VDD.n1888 VSS 0.309003f
C18849 VDD.n1889 VSS 0.77922f
C18850 VDD.n1890 VSS 0.116823f
C18851 VDD.t4402 VSS 0.066856f
C18852 VDD.n1891 VSS 0.14405f
C18853 VDD.n1892 VSS 0.120118f
C18854 VDD.n1893 VSS 0.016021f
C18855 VDD.t1446 VSS 0.025104f
C18856 VDD.n1894 VSS 0.105404f
C18857 VDD.n1895 VSS 0.057098f
C18858 VDD.t1660 VSS 1.45794f
C18859 VDD.t804 VSS 1.96535f
C18860 VDD.t647 VSS 1.96535f
C18861 VDD.t1445 VSS 1.36988f
C18862 VDD.n1896 VSS 0.645798f
C18863 VDD.t858 VSS 1.45794f
C18864 VDD.n1897 VSS 0.206947f
C18865 VDD.n1898 VSS 0.208771f
C18866 VDD.t3095 VSS 0.028519f
C18867 VDD.t2123 VSS 0.028519f
C18868 VDD.n1899 VSS 0.009191f
C18869 VDD.t3993 VSS 0.028519f
C18870 VDD.t2683 VSS 0.028519f
C18871 VDD.n1900 VSS 0.009191f
C18872 VDD.n1901 VSS 0.528101f
C18873 VDD.t4603 VSS 0.028519f
C18874 VDD.t3718 VSS 0.028519f
C18875 VDD.n1902 VSS 0.009191f
C18876 VDD.t4602 VSS 0.066856f
C18877 VDD.t1401 VSS 0.066856f
C18878 VDD.t4254 VSS 0.066856f
C18879 VDD.t1051 VSS 0.066856f
C18880 VDD.t4255 VSS 0.028519f
C18881 VDD.t3341 VSS 0.028519f
C18882 VDD.n1903 VSS 0.009191f
C18883 VDD.t2443 VSS 0.066856f
C18884 VDD.t1925 VSS 0.066856f
C18885 VDD.t2444 VSS 0.028519f
C18886 VDD.t2179 VSS 0.028519f
C18887 VDD.n1904 VSS 0.009191f
C18888 VDD.t3568 VSS 0.066856f
C18889 VDD.n1905 VSS 0.14405f
C18890 VDD.t576 VSS 0.025104f
C18891 VDD.t3570 VSS 0.066856f
C18892 VDD.n1906 VSS 0.14405f
C18893 VDD.t3370 VSS 0.025104f
C18894 VDD.n1907 VSS 0.04911f
C18895 VDD.t2573 VSS 0.028519f
C18896 VDD.t4321 VSS 0.028519f
C18897 VDD.n1908 VSS 0.009191f
C18898 VDD.t4161 VSS 0.028519f
C18899 VDD.t3815 VSS 0.028519f
C18900 VDD.n1909 VSS 0.009191f
C18901 VDD.n1910 VSS 0.523473f
C18902 VDD.n1911 VSS 0.207221f
C18903 VDD.n1912 VSS 0.206947f
C18904 VDD.n1913 VSS 0.208771f
C18905 VDD.t2122 VSS 1.96535f
C18906 VDD.t1843 VSS 1.96535f
C18907 VDD.t575 VSS 1.36988f
C18908 VDD.n1914 VSS 0.645798f
C18909 VDD.n1915 VSS 0.595476f
C18910 VDD.t3571 VSS 1.31955f
C18911 VDD.t2926 VSS 1.96535f
C18912 VDD.t1186 VSS 1.96535f
C18913 VDD.t908 VSS 1.45794f
C18914 VDD.n1916 VSS 0.865258f
C18915 VDD.n1917 VSS 0.865258f
C18916 VDD.n1918 VSS 0.092503f
C18917 VDD.n1919 VSS 0.236396f
C18918 VDD.n1920 VSS 0.206947f
C18919 VDD.n1921 VSS 0.207221f
C18920 VDD.n1922 VSS 0.057098f
C18921 VDD.t1938 VSS 1.45794f
C18922 VDD.t878 VSS 1.96535f
C18923 VDD.t1381 VSS 1.96535f
C18924 VDD.t869 VSS 1.36988f
C18925 VDD.n1923 VSS 0.645798f
C18926 VDD.t801 VSS 1.45794f
C18927 VDD.n1924 VSS 0.206947f
C18928 VDD.n1925 VSS 0.208771f
C18929 VDD.t802 VSS 0.028519f
C18930 VDD.t3275 VSS 0.028519f
C18931 VDD.n1926 VSS 0.009191f
C18932 VDD.t1266 VSS 0.028519f
C18933 VDD.t4187 VSS 0.028519f
C18934 VDD.n1927 VSS 0.009191f
C18935 VDD.n1928 VSS 0.528101f
C18936 VDD.t2486 VSS 0.028519f
C18937 VDD.t643 VSS 0.028519f
C18938 VDD.n1929 VSS 0.009191f
C18939 VDD.t2485 VSS 0.066856f
C18940 VDD.t2966 VSS 0.066856f
C18941 VDD.t2025 VSS 0.066856f
C18942 VDD.t2597 VSS 0.066856f
C18943 VDD.t2026 VSS 0.028519f
C18944 VDD.t4413 VSS 0.028519f
C18945 VDD.n1930 VSS 0.009191f
C18946 VDD.t3216 VSS 0.066856f
C18947 VDD.t4168 VSS 0.066856f
C18948 VDD.t3217 VSS 0.028519f
C18949 VDD.t4333 VSS 0.028519f
C18950 VDD.n1931 VSS 0.009191f
C18951 VDD.t2097 VSS 0.066856f
C18952 VDD.n1932 VSS 0.14405f
C18953 VDD.t3015 VSS 0.025104f
C18954 VDD.t667 VSS 0.066856f
C18955 VDD.n1933 VSS 0.14405f
C18956 VDD.t2545 VSS 0.025104f
C18957 VDD.n1934 VSS 0.04911f
C18958 VDD.t3081 VSS 0.028519f
C18959 VDD.t2760 VSS 0.028519f
C18960 VDD.n1935 VSS 0.009191f
C18961 VDD.t2576 VSS 0.028519f
C18962 VDD.t4325 VSS 0.028519f
C18963 VDD.n1936 VSS 0.009191f
C18964 VDD.n1937 VSS 0.523473f
C18965 VDD.n1938 VSS 0.207221f
C18966 VDD.n1939 VSS 0.206947f
C18967 VDD.n1940 VSS 0.208771f
C18968 VDD.t642 VSS 1.96535f
C18969 VDD.t493 VSS 1.96535f
C18970 VDD.t495 VSS 1.36988f
C18971 VDD.n1941 VSS 0.645798f
C18972 VDD.n1942 VSS 0.595476f
C18973 VDD.t494 VSS 1.31955f
C18974 VDD.t492 VSS 1.96535f
C18975 VDD.t2575 VSS 1.96535f
C18976 VDD.t1376 VSS 1.45794f
C18977 VDD.n1943 VSS 0.865258f
C18978 VDD.n1944 VSS 0.865258f
C18979 VDD.t678 VSS 0.028519f
C18980 VDD.t4489 VSS 0.028519f
C18981 VDD.n1945 VSS 0.009191f
C18982 VDD.t4323 VSS 0.028519f
C18983 VDD.t2013 VSS 0.028519f
C18984 VDD.n1946 VSS 0.009191f
C18985 VDD.n1947 VSS 0.523473f
C18986 VDD.t2357 VSS 0.028519f
C18987 VDD.t1945 VSS 0.028519f
C18988 VDD.n1948 VSS 0.009191f
C18989 VDD.t1743 VSS 0.028519f
C18990 VDD.t3610 VSS 0.028519f
C18991 VDD.n1949 VSS 0.009191f
C18992 VDD.n1950 VSS 0.471397f
C18993 VDD.n1951 VSS 0.206947f
C18994 VDD.n1952 VSS 0.207221f
C18995 VDD.t4432 VSS 0.066856f
C18996 VDD.n1953 VSS 0.14405f
C18997 VDD.t4635 VSS 0.025104f
C18998 VDD.t3678 VSS 0.066856f
C18999 VDD.n1954 VSS 0.14405f
C19000 VDD.t1409 VSS 0.025104f
C19001 VDD.t3676 VSS 0.066856f
C19002 VDD.n1955 VSS 0.14405f
C19003 VDD.t3889 VSS 0.025104f
C19004 VDD.n1956 VSS 0.033925f
C19005 VDD.t508 VSS 0.019767f
C19006 VDD.t511 VSS 0.018805f
C19007 VDD.n1957 VSS 0.054793f
C19008 VDD.t509 VSS 0.018792f
C19009 VDD.t510 VSS 0.019781f
C19010 VDD.n1958 VSS 0.077486f
C19011 VDD.n1959 VSS 0.252514f
C19012 VDD.n1960 VSS 0.199549f
C19013 VDD.n1961 VSS 0.060108f
C19014 VDD.t3888 VSS 0.066856f
C19015 VDD.n1962 VSS 0.131361f
C19016 VDD.n1963 VSS 0.120118f
C19017 VDD.n1964 VSS 0.016021f
C19018 VDD.t3677 VSS 0.025104f
C19019 VDD.n1965 VSS 0.105404f
C19020 VDD.n1966 VSS 0.057098f
C19021 VDD.n1967 VSS 0.087217f
C19022 VDD.t1407 VSS 0.066856f
C19023 VDD.n1968 VSS 0.14405f
C19024 VDD.n1969 VSS 0.120118f
C19025 VDD.n1970 VSS 0.016021f
C19026 VDD.t3680 VSS 0.025104f
C19027 VDD.n1971 VSS 0.116823f
C19028 VDD.t2356 VSS 0.066856f
C19029 VDD.t1742 VSS 0.066856f
C19030 VDD.t3609 VSS 0.066856f
C19031 VDD.t1944 VSS 0.066856f
C19032 VDD.n1972 VSS 0.690489f
C19033 VDD.t1897 VSS 0.066856f
C19034 VDD.t1372 VSS 0.066856f
C19035 VDD.t3284 VSS 0.066856f
C19036 VDD.t1550 VSS 0.066856f
C19037 VDD.n1973 VSS 0.690489f
C19038 VDD.t1898 VSS 0.028519f
C19039 VDD.t1552 VSS 0.028519f
C19040 VDD.n1974 VSS 0.009191f
C19041 VDD.t1374 VSS 0.028519f
C19042 VDD.t3285 VSS 0.028519f
C19043 VDD.n1975 VSS 0.009191f
C19044 VDD.n1976 VSS 0.644755f
C19045 VDD.t2052 VSS 0.066856f
C19046 VDD.t4494 VSS 0.066856f
C19047 VDD.t1182 VSS 0.066856f
C19048 VDD.t2182 VSS 0.066856f
C19049 VDD.n1977 VSS 0.709674f
C19050 VDD.t2053 VSS 0.028519f
C19051 VDD.t2183 VSS 0.028519f
C19052 VDD.n1978 VSS 0.009191f
C19053 VDD.t4495 VSS 0.028519f
C19054 VDD.t1184 VSS 0.028519f
C19055 VDD.n1979 VSS 0.009191f
C19056 VDD.n1980 VSS 0.309003f
C19057 VDD.n1981 VSS 0.77922f
C19058 VDD.n1982 VSS 0.116823f
C19059 VDD.t4634 VSS 0.066856f
C19060 VDD.n1983 VSS 0.14405f
C19061 VDD.n1984 VSS 0.120118f
C19062 VDD.n1985 VSS 0.016021f
C19063 VDD.t4433 VSS 0.025104f
C19064 VDD.n1986 VSS 0.105404f
C19065 VDD.n1987 VSS 0.057098f
C19066 VDD.t677 VSS 1.45794f
C19067 VDD.t1551 VSS 1.96535f
C19068 VDD.t496 VSS 1.96535f
C19069 VDD.t498 VSS 1.36988f
C19070 VDD.n1988 VSS 0.645798f
C19071 VDD.t1167 VSS 1.45794f
C19072 VDD.n1989 VSS 0.206947f
C19073 VDD.n1990 VSS 0.208771f
C19074 VDD.t1878 VSS 0.028519f
C19075 VDD.t4667 VSS 0.028519f
C19076 VDD.n1991 VSS 0.009191f
C19077 VDD.t2935 VSS 0.028519f
C19078 VDD.t1443 VSS 0.028519f
C19079 VDD.n1992 VSS 0.009191f
C19080 VDD.n1993 VSS 0.528101f
C19081 VDD.t3505 VSS 0.028519f
C19082 VDD.t2118 VSS 0.028519f
C19083 VDD.n1994 VSS 0.009191f
C19084 VDD.t3504 VSS 0.066856f
C19085 VDD.t4430 VSS 0.066856f
C19086 VDD.t3174 VSS 0.066856f
C19087 VDD.t4074 VSS 0.066856f
C19088 VDD.t3175 VSS 0.028519f
C19089 VDD.t1717 VSS 0.028519f
C19090 VDD.n1995 VSS 0.009191f
C19091 VDD.t1166 VSS 0.066856f
C19092 VDD.t772 VSS 0.066856f
C19093 VDD.n1996 VSS 0.018249f
C19094 VDD.n1997 VSS 0.018625f
C19095 VDD.t1168 VSS 0.028519f
C19096 VDD.t2472 VSS 0.028519f
C19097 VDD.n1998 VSS 0.009191f
C19098 VDD.t773 VSS 0.028519f
C19099 VDD.t1957 VSS 0.028519f
C19100 VDD.n1999 VSS 0.009191f
C19101 VDD.n2000 VSS 0.10689f
C19102 VDD.n2001 VSS 0.01502f
C19103 VDD.n2002 VSS 0.009688f
C19104 VDD.n2004 VSS 0.074698f
C19105 VDD.t3938 VSS 0.066856f
C19106 VDD.n2005 VSS 0.14405f
C19107 VDD.t1004 VSS 0.025104f
C19108 VDD.t2938 VSS 0.066856f
C19109 VDD.n2006 VSS 0.14405f
C19110 VDD.t2742 VSS 0.025104f
C19111 VDD.n2007 VSS 0.04911f
C19112 VDD.t1326 VSS 0.028519f
C19113 VDD.t4153 VSS 0.028519f
C19114 VDD.n2008 VSS 0.009191f
C19115 VDD.t1210 VSS 0.028519f
C19116 VDD.t4029 VSS 0.028519f
C19117 VDD.n2009 VSS 0.009191f
C19118 VDD.n2010 VSS 0.523473f
C19119 VDD.n2011 VSS 0.207221f
C19120 VDD.n2012 VSS 0.206947f
C19121 VDD.n2013 VSS 0.208771f
C19122 VDD.t1716 VSS 1.96535f
C19123 VDD.t290 VSS 1.96535f
C19124 VDD.t293 VSS 1.36988f
C19125 VDD.n2014 VSS 0.645798f
C19126 VDD.n2015 VSS 0.595476f
C19127 VDD.t292 VSS 1.31955f
C19128 VDD.t291 VSS 1.96535f
C19129 VDD.t1209 VSS 1.96535f
C19130 VDD.t1084 VSS 1.45794f
C19131 VDD.n2016 VSS 0.865258f
C19132 VDD.n2017 VSS 0.865258f
C19133 VDD.t3251 VSS 0.028519f
C19134 VDD.t2353 VSS 0.028519f
C19135 VDD.n2018 VSS 0.009191f
C19136 VDD.t681 VSS 0.028519f
C19137 VDD.t3489 VSS 0.028519f
C19138 VDD.n2019 VSS 0.009191f
C19139 VDD.n2020 VSS 0.523473f
C19140 VDD.t603 VSS 0.028519f
C19141 VDD.t3881 VSS 0.028519f
C19142 VDD.n2021 VSS 0.009191f
C19143 VDD.t2363 VSS 0.028519f
C19144 VDD.t934 VSS 0.028519f
C19145 VDD.n2022 VSS 0.009191f
C19146 VDD.n2023 VSS 0.471397f
C19147 VDD.n2024 VSS 0.206947f
C19148 VDD.n2025 VSS 1.049f
C19149 VDD.t3040 VSS 0.066856f
C19150 VDD.n2026 VSS 0.14405f
C19151 VDD.t1733 VSS 0.025104f
C19152 VDD.t601 VSS 0.066856f
C19153 VDD.t2362 VSS 0.066856f
C19154 VDD.t932 VSS 0.066856f
C19155 VDD.t3880 VSS 0.066856f
C19156 VDD.n2027 VSS 0.690489f
C19157 VDD.t4394 VSS 0.066856f
C19158 VDD.t1899 VSS 0.066856f
C19159 VDD.t4684 VSS 0.066856f
C19160 VDD.t3512 VSS 0.066856f
C19161 VDD.n2028 VSS 0.690489f
C19162 VDD.t4395 VSS 0.028519f
C19163 VDD.t3513 VSS 0.028519f
C19164 VDD.n2029 VSS 0.009191f
C19165 VDD.t1900 VSS 0.028519f
C19166 VDD.t4685 VSS 0.028519f
C19167 VDD.n2030 VSS 0.009191f
C19168 VDD.n2031 VSS 0.644755f
C19169 VDD.t3222 VSS 0.066856f
C19170 VDD.t2229 VSS 0.066856f
C19171 VDD.t3426 VSS 0.066856f
C19172 VDD.t3038 VSS 0.066856f
C19173 VDD.n2032 VSS 0.709674f
C19174 VDD.t3223 VSS 0.028519f
C19175 VDD.t3039 VSS 0.028519f
C19176 VDD.n2033 VSS 0.009191f
C19177 VDD.t2230 VSS 0.028519f
C19178 VDD.t3427 VSS 0.028519f
C19179 VDD.n2034 VSS 0.009191f
C19180 VDD.n2035 VSS 0.309003f
C19181 VDD.t3423 VSS 0.066856f
C19182 VDD.n2036 VSS 0.14405f
C19183 VDD.t3615 VSS 0.025104f
C19184 VDD.t1712 VSS 0.066856f
C19185 VDD.n2037 VSS 0.14405f
C19186 VDD.t4683 VSS 0.025104f
C19187 VDD.n2038 VSS 0.033925f
C19188 VDD.t507 VSS 0.019767f
C19189 VDD.t506 VSS 0.018805f
C19190 VDD.n2039 VSS 0.054793f
C19191 VDD.t504 VSS 0.018792f
C19192 VDD.t505 VSS 0.019781f
C19193 VDD.n2040 VSS 0.077486f
C19194 VDD.n2041 VSS 0.252514f
C19195 VDD.n2042 VSS 0.199549f
C19196 VDD.n2043 VSS 0.060108f
C19197 VDD.t4682 VSS 0.066856f
C19198 VDD.n2044 VSS 0.131361f
C19199 VDD.n2045 VSS 0.120118f
C19200 VDD.n2046 VSS 0.016021f
C19201 VDD.t1714 VSS 0.025104f
C19202 VDD.n2047 VSS 0.105404f
C19203 VDD.n2048 VSS 0.057098f
C19204 VDD.n2049 VSS 0.087217f
C19205 VDD.t3613 VSS 0.066856f
C19206 VDD.n2050 VSS 0.14405f
C19207 VDD.n2051 VSS 0.120118f
C19208 VDD.n2052 VSS 0.016021f
C19209 VDD.t3425 VSS 0.025104f
C19210 VDD.n2053 VSS 0.116823f
C19211 VDD.n2054 VSS 0.77922f
C19212 VDD.n2055 VSS 0.116823f
C19213 VDD.t1732 VSS 0.066856f
C19214 VDD.n2056 VSS 0.14405f
C19215 VDD.n2057 VSS 0.120118f
C19216 VDD.n2058 VSS 0.016021f
C19217 VDD.t3041 VSS 0.025104f
C19218 VDD.n2059 VSS 0.105404f
C19219 VDD.t672 VSS 0.066856f
C19220 VDD.n2060 VSS 0.14405f
C19221 VDD.t4617 VSS 0.025104f
C19222 VDD.n2061 VSS 0.054485f
C19223 VDD.n2062 VSS 0.106951f
C19224 VDD.n2063 VSS 0.012131f
C19225 VDD.t3036 VSS 0.066856f
C19226 VDD.t4184 VSS 0.066856f
C19227 VDD.n2064 VSS 0.10134f
C19228 VDD.n2065 VSS 0.012131f
C19229 VDD.n2066 VSS 0.106951f
C19230 VDD.n2067 VSS 0.012131f
C19231 VDD.n2068 VSS 0.080214f
C19232 VDD.n2069 VSS 0.012131f
C19233 VDD.n2070 VSS 0.106951f
C19234 VDD.n2071 VSS 0.012131f
C19235 VDD.n2072 VSS 0.090303f
C19236 VDD.n2073 VSS 0.012131f
C19237 VDD.n2074 VSS 0.053476f
C19238 VDD.n2075 VSS 0.012131f
C19239 VDD.n2076 VSS 0.102411f
C19240 VDD.n2077 VSS 0.012131f
C19241 VDD.t4304 VSS 0.066856f
C19242 VDD.t3020 VSS 0.066856f
C19243 VDD.n2078 VSS 0.10134f
C19244 VDD.n2079 VSS 0.012131f
C19245 VDD.n2080 VSS 0.106951f
C19246 VDD.n2081 VSS 0.012131f
C19247 VDD.n2082 VSS 0.102411f
C19248 VDD.n2083 VSS 0.012131f
C19249 VDD.n2084 VSS 0.106951f
C19250 VDD.n2085 VSS 0.012131f
C19251 VDD.n2086 VSS 0.106951f
C19252 VDD.n2087 VSS 0.012131f
C19253 VDD.n2088 VSS 0.068106f
C19254 VDD.n2089 VSS 0.035132f
C19255 VDD.t2151 VSS 0.025104f
C19256 VDD.t1981 VSS 0.066856f
C19257 VDD.n2090 VSS 0.125227f
C19258 VDD.t3368 VSS 0.025104f
C19259 VDD.t3550 VSS 0.066856f
C19260 VDD.n2091 VSS 0.125227f
C19261 VDD.t4451 VSS 0.025104f
C19262 VDD.t4298 VSS 0.066856f
C19263 VDD.n2092 VSS 0.125227f
C19264 VDD.t1498 VSS 0.025104f
C19265 VDD.t3335 VSS 0.028519f
C19266 VDD.t1932 VSS 0.028519f
C19267 VDD.n2093 VSS 0.009191f
C19268 VDD.t3334 VSS 0.066856f
C19269 VDD.t3256 VSS 0.066856f
C19270 VDD.t3043 VSS 0.028519f
C19271 VDD.t1566 VSS 0.028519f
C19272 VDD.n2094 VSS 0.009191f
C19273 VDD.t3042 VSS 0.066856f
C19274 VDD.t2928 VSS 0.066856f
C19275 VDD.t1324 VSS 0.066856f
C19276 VDD.t1208 VSS 0.066856f
C19277 VDD.t4028 VSS 0.066856f
C19278 VDD.t4152 VSS 0.066856f
C19279 VDD.n2095 VSS 0.690489f
C19280 VDD.t1435 VSS 0.066856f
C19281 VDD.t1565 VSS 0.066856f
C19282 VDD.n2096 VSS 0.690489f
C19283 VDD.t2929 VSS 0.028519f
C19284 VDD.t1436 VSS 0.028519f
C19285 VDD.n2097 VSS 0.009191f
C19286 VDD.n2098 VSS 0.644755f
C19287 VDD.t1795 VSS 0.066856f
C19288 VDD.t1931 VSS 0.066856f
C19289 VDD.n2099 VSS 0.709674f
C19290 VDD.t3257 VSS 0.028519f
C19291 VDD.t1796 VSS 0.028519f
C19292 VDD.n2100 VSS 0.009191f
C19293 VDD.n2101 VSS 0.261039f
C19294 VDD.t4106 VSS 0.066856f
C19295 VDD.n2102 VSS 0.125227f
C19296 VDD.t865 VSS 0.025104f
C19297 VDD.t674 VSS 0.066856f
C19298 VDD.n2103 VSS 0.125227f
C19299 VDD.t2085 VSS 0.025104f
C19300 VDD.n2104 VSS 0.08403f
C19301 VDD.n2105 VSS 0.471009f
C19302 VDD.t3865 VSS 0.028519f
C19303 VDD.t2570 VSS 0.028519f
C19304 VDD.n2106 VSS 0.009191f
C19305 VDD.n2109 VSS 0.01487f
C19306 VDD.n2110 VSS 0.018625f
C19307 VDD.t3864 VSS 0.066856f
C19308 VDD.t651 VSS 0.066856f
C19309 VDD.t3517 VSS 0.028519f
C19310 VDD.t2138 VSS 0.028519f
C19311 VDD.n2111 VSS 0.009191f
C19312 VDD.t3516 VSS 0.066856f
C19313 VDD.t4456 VSS 0.066856f
C19314 VDD.t1877 VSS 0.066856f
C19315 VDD.t2934 VSS 0.066856f
C19316 VDD.t1441 VSS 0.066856f
C19317 VDD.t4666 VSS 0.066856f
C19318 VDD.n2112 VSS 0.696076f
C19319 VDD.t3154 VSS 0.066856f
C19320 VDD.t2137 VSS 0.066856f
C19321 VDD.n2113 VSS 0.696076f
C19322 VDD.t4457 VSS 0.028519f
C19323 VDD.t3155 VSS 0.028519f
C19324 VDD.n2114 VSS 0.009191f
C19325 VDD.n2115 VSS 0.650522f
C19326 VDD.t3464 VSS 0.066856f
C19327 VDD.t2569 VSS 0.066856f
C19328 VDD.n2116 VSS 0.635903f
C19329 VDD.n2118 VSS 0.018249f
C19330 VDD.n2119 VSS 0.020119f
C19331 VDD.n2120 VSS 0.058553f
C19332 VDD.t4687 VSS 0.019983f
C19333 VDD.n2121 VSS 0.336192f
C19334 VDD.t863 VSS 0.014798f
C19335 VDD.t862 VSS 0.043485f
C19336 VDD.n2122 VSS 0.095207f
C19337 VDD.n2123 VSS 1.83791f
C19338 VDD.n2124 VSS 0.154958f
C19339 VDD.t965 VSS 3.35166f
C19340 VDD.t389 VSS 4.24765f
C19341 VDD.t406 VSS 2.51852f
C19342 VDD.t401 VSS 2.42329f
C19343 VDD.t944 VSS 0.043485f
C19344 VDD.n2125 VSS 0.081263f
C19345 VDD.t2842 VSS 0.043485f
C19346 VDD.n2126 VSS 0.097632f
C19347 VDD.t2086 VSS 0.043485f
C19348 VDD.n2127 VSS 0.097632f
C19349 VDD.t1027 VSS 0.019983f
C19350 VDD.t2413 VSS 0.019983f
C19351 VDD.t2299 VSS 0.043485f
C19352 VDD.t3327 VSS 0.019983f
C19353 VDD.t2300 VSS 0.019983f
C19354 VDD.t775 VSS 0.019983f
C19355 VDD.t3871 VSS 0.019983f
C19356 VDD.t3870 VSS 0.043485f
C19357 VDD.t2846 VSS 0.043485f
C19358 VDD.t3803 VSS 0.019983f
C19359 VDD.t2847 VSS 0.019983f
C19360 VDD.t964 VSS 0.043485f
C19361 VDD.t413 VSS 0.011309f
C19362 VDD.n2128 VSS 0.076307f
C19363 VDD.t1992 VSS 0.019983f
C19364 VDD.t966 VSS 0.019983f
C19365 VDD.n2129 VSS 0.380982f
C19366 VDD.n2130 VSS 0.176495f
C19367 VDD.t1991 VSS 0.043485f
C19368 VDD.n2131 VSS 0.206328f
C19369 VDD.n2132 VSS 0.279289f
C19370 VDD.t3802 VSS 0.043485f
C19371 VDD.n2133 VSS 0.240634f
C19372 VDD.t774 VSS 0.043485f
C19373 VDD.n2134 VSS 0.240634f
C19374 VDD.n2135 VSS 0.231506f
C19375 VDD.n2136 VSS 0.239326f
C19376 VDD.n2137 VSS 0.224971f
C19377 VDD.t3326 VSS 0.043485f
C19378 VDD.n2138 VSS 0.200074f
C19379 VDD.t2412 VSS 0.043485f
C19380 VDD.n2139 VSS 0.116954f
C19381 VDD.n2140 VSS 0.139266f
C19382 VDD.t1026 VSS 0.043485f
C19383 VDD.n2141 VSS 0.14628f
C19384 VDD.n2142 VSS 0.211734f
C19385 VDD.n2143 VSS 0.098613f
C19386 VDD.t2087 VSS 0.019983f
C19387 VDD.n2144 VSS 0.083454f
C19388 VDD.n2145 VSS 0.083454f
C19389 VDD.t945 VSS 0.014798f
C19390 VDD.t1362 VSS 0.014798f
C19391 VDD.t1100 VSS 0.034186f
C19392 VDD.n2146 VSS 0.232449f
C19393 VDD.t573 VSS 0.019983f
C19394 VDD.t1913 VSS 0.019983f
C19395 VDD.n2147 VSS 0.124683f
C19396 VDD.t1119 VSS 0.066856f
C19397 VDD.n2148 VSS 0.154846f
C19398 VDD.t3781 VSS 0.034186f
C19399 VDD.t2200 VSS 0.034186f
C19400 VDD.t927 VSS 0.066856f
C19401 VDD.n2149 VSS 0.215845f
C19402 VDD.n2150 VSS 0.00473f
C19403 VDD.n2151 VSS 0.00473f
C19404 VDD.n2152 VSS 0.00473f
C19405 VDD.n2153 VSS 0.00473f
C19406 VDD.n2154 VSS 0.00473f
C19407 VDD.n2155 VSS 0.00473f
C19408 VDD.t1912 VSS 0.043485f
C19409 VDD.n2156 VSS 0.142069f
C19410 VDD.t3753 VSS 0.034186f
C19411 VDD.n2157 VSS 0.135294f
C19412 VDD.t1830 VSS 0.043485f
C19413 VDD.n2158 VSS 0.14041f
C19414 VDD.t3752 VSS 0.066856f
C19415 VDD.n2159 VSS 0.114368f
C19416 VDD.t1831 VSS 0.019983f
C19417 VDD.n2160 VSS 0.171561f
C19418 VDD.t2172 VSS 0.066856f
C19419 VDD.n2161 VSS 0.142163f
C19420 VDD.n2162 VSS 0.123623f
C19421 VDD.t2173 VSS 0.034186f
C19422 VDD.n2163 VSS 0.140273f
C19423 VDD.t3475 VSS 0.019983f
C19424 VDD.n2164 VSS 0.109749f
C19425 VDD.t3474 VSS 0.043485f
C19426 VDD.n2165 VSS 0.155344f
C19427 VDD.t2430 VSS 0.019983f
C19428 VDD.t914 VSS 0.034186f
C19429 VDD.t4276 VSS 0.066856f
C19430 VDD.n2166 VSS 0.126716f
C19431 VDD.t3378 VSS 0.016021f
C19432 VDD.t4728 VSS 0.066856f
C19433 VDD.n2167 VSS 0.126716f
C19434 VDD.t3835 VSS 0.025104f
C19435 VDD.t1586 VSS 0.066856f
C19436 VDD.n2168 VSS 0.126716f
C19437 VDD.t4375 VSS 0.016021f
C19438 VDD.t3494 VSS 0.066856f
C19439 VDD.n2169 VSS 0.126716f
C19440 VDD.t2671 VSS 0.066856f
C19441 VDD.n2170 VSS 0.126716f
C19442 VDD.t1189 VSS 0.016021f
C19443 VDD.t4108 VSS 0.066856f
C19444 VDD.n2171 VSS 0.126716f
C19445 VDD.t2804 VSS 0.025104f
C19446 VDD.t929 VSS 0.034186f
C19447 VDD.n2172 VSS 0.273827f
C19448 VDD.n2173 VSS 0.137101f
C19449 VDD.t2803 VSS 0.066856f
C19450 VDD.n2174 VSS 0.126716f
C19451 VDD.n2175 VSS 0.102784f
C19452 VDD.n2176 VSS 0.016021f
C19453 VDD.t4109 VSS 0.016021f
C19454 VDD.n2177 VSS 0.016021f
C19455 VDD.n2178 VSS 0.102784f
C19456 VDD.t1188 VSS 0.066856f
C19457 VDD.n2179 VSS 0.126716f
C19458 VDD.n2180 VSS 0.102784f
C19459 VDD.n2181 VSS 0.016021f
C19460 VDD.t2672 VSS 0.025104f
C19461 VDD.n2182 VSS 0.107953f
C19462 VDD.n2183 VSS 0.107953f
C19463 VDD.t3495 VSS 0.025104f
C19464 VDD.n2184 VSS 0.016021f
C19465 VDD.n2185 VSS 0.102784f
C19466 VDD.t4374 VSS 0.066856f
C19467 VDD.n2186 VSS 0.082381f
C19468 VDD.n2187 VSS 0.310374f
C19469 VDD.n2188 VSS 1.94948f
C19470 VDD.t30 VSS 3.42569f
C19471 VDD.t928 VSS 3.43836f
C19472 VDD.t37 VSS 3.66626f
C19473 VDD.t23 VSS 2.8468f
C19474 VDD.t28 VSS 2.8468f
C19475 VDD.t35 VSS 3.52342f
C19476 VDD.t17 VSS 3.52342f
C19477 VDD.t26 VSS 1.52113f
C19478 VDD.n2189 VSS 0.218448f
C19479 VDD.t2008 VSS 0.066856f
C19480 VDD.n2190 VSS 0.272089f
C19481 VDD.t2474 VSS 0.016021f
C19482 VDD.t3793 VSS 0.025104f
C19483 VDD.t1020 VSS 0.066856f
C19484 VDD.n2191 VSS 0.272089f
C19485 VDD.n2192 VSS 0.248157f
C19486 VDD.n2193 VSS 0.251491f
C19487 VDD.t3646 VSS 0.066856f
C19488 VDD.n2194 VSS 0.259856f
C19489 VDD.t2473 VSS 0.066856f
C19490 VDD.n2195 VSS 0.272089f
C19491 VDD.t3401 VSS 0.066856f
C19492 VDD.n2196 VSS 0.272089f
C19493 VDD.t1431 VSS 0.066856f
C19494 VDD.n2197 VSS 0.309663f
C19495 VDD.t2442 VSS 0.016021f
C19496 VDD.t3687 VSS 0.066856f
C19497 VDD.n2198 VSS 0.27209f
C19498 VDD.n2199 VSS 0.649726f
C19499 VDD.t1884 VSS 0.025104f
C19500 VDD.t3350 VSS 0.066856f
C19501 VDD.n2200 VSS 0.27209f
C19502 VDD.t1013 VSS 0.066856f
C19503 VDD.n2201 VSS 0.254614f
C19504 VDD.n2202 VSS 0.25586f
C19505 VDD.t1307 VSS 0.016021f
C19506 VDD.t2758 VSS 0.034186f
C19507 VDD.n2203 VSS 0.183335f
C19508 VDD.t1384 VSS 0.034186f
C19509 VDD.n2204 VSS 0.155079f
C19510 VDD.t2785 VSS 0.066856f
C19511 VDD.n2205 VSS 0.168108f
C19512 VDD.n2206 VSS 0.280079f
C19513 VDD.t1216 VSS 0.066856f
C19514 VDD.n2207 VSS 0.309663f
C19515 VDD.t1217 VSS 0.025104f
C19516 VDD.t4467 VSS 0.025104f
C19517 VDD.t1204 VSS 0.066856f
C19518 VDD.n2208 VSS 0.126927f
C19519 VDD.t2196 VSS 0.034186f
C19520 VDD.n2209 VSS 0.198913f
C19521 VDD.n2210 VSS 0.279865f
C19522 VDD.t3062 VSS 0.066856f
C19523 VDD.n2211 VSS 0.244128f
C19524 VDD.n2212 VSS 0.248157f
C19525 VDD.t3063 VSS 0.016021f
C19526 VDD.t4481 VSS 0.025104f
C19527 VDD.t1693 VSS 0.066856f
C19528 VDD.n2213 VSS 0.272089f
C19529 VDD.t4386 VSS 0.066856f
C19530 VDD.n2214 VSS 0.272089f
C19531 VDD.n2215 VSS 0.255859f
C19532 VDD.n2216 VSS 0.255859f
C19533 VDD.t4480 VSS 0.066856f
C19534 VDD.n2217 VSS 0.259856f
C19535 VDD.t3380 VSS 0.025104f
C19536 VDD.n2218 VSS 0.251491f
C19537 VDD.n2219 VSS 0.247995f
C19538 VDD.t4360 VSS 0.066856f
C19539 VDD.n2220 VSS 0.272089f
C19540 VDD.t3379 VSS 0.066856f
C19541 VDD.n2221 VSS 0.272089f
C19542 VDD.t4361 VSS 0.025104f
C19543 VDD.n2222 VSS 0.016021f
C19544 VDD.n2223 VSS 0.248157f
C19545 VDD.n2224 VSS 0.248157f
C19546 VDD.n2225 VSS 0.016021f
C19547 VDD.t1994 VSS 0.016021f
C19548 VDD.n2226 VSS 0.016021f
C19549 VDD.t4387 VSS 0.025104f
C19550 VDD.n2227 VSS 0.255859f
C19551 VDD.n2228 VSS 0.248157f
C19552 VDD.n2229 VSS 0.016021f
C19553 VDD.t1694 VSS 0.016021f
C19554 VDD.n2230 VSS 0.016021f
C19555 VDD.n2231 VSS 0.248157f
C19556 VDD.t1993 VSS 0.066856f
C19557 VDD.n2232 VSS 0.056262f
C19558 VDD.n2233 VSS 0.243788f
C19559 VDD.n2234 VSS 0.283109f
C19560 VDD.t597 VSS 9.19382f
C19561 VDD.n2235 VSS 0.283088f
C19562 VDD.n2236 VSS 0.283088f
C19563 VDD.n2237 VSS 0.279865f
C19564 VDD.n2238 VSS 0.283109f
C19565 VDD.t4121 VSS 0.034186f
C19566 VDD.n2239 VSS 0.198913f
C19567 VDD.t1012 VSS 0.034186f
C19568 VDD.t598 VSS 0.034186f
C19569 VDD.t4336 VSS 0.066856f
C19570 VDD.t2332 VSS 0.066856f
C19571 VDD.n2240 VSS 0.191511f
C19572 VDD.n2241 VSS 0.266053f
C19573 VDD.t2055 VSS 0.034186f
C19574 VDD.t1665 VSS 0.034186f
C19575 VDD.n2242 VSS 0.007954f
C19576 VDD.n2243 VSS 0.260606f
C19577 VDD.n2244 VSS 0.012131f
C19578 VDD.n2245 VSS 0.012131f
C19579 VDD.n2246 VSS 0.260606f
C19580 VDD.n2247 VSS 0.012131f
C19581 VDD.t3955 VSS 0.034186f
C19582 VDD.t3954 VSS 0.066856f
C19583 VDD.n2248 VSS 0.284538f
C19584 VDD.n2249 VSS 0.012131f
C19585 VDD.t3587 VSS 0.066856f
C19586 VDD.n2250 VSS 0.154235f
C19587 VDD.n2251 VSS 0.012131f
C19588 VDD.t3588 VSS 0.034186f
C19589 VDD.n2252 VSS 0.145708f
C19590 VDD.n2253 VSS 0.012131f
C19591 VDD.n2254 VSS 0.260606f
C19592 VDD.n2255 VSS 0.012131f
C19593 VDD.n2256 VSS 0.260606f
C19594 VDD.n2257 VSS 0.012131f
C19595 VDD.n2258 VSS 0.233562f
C19596 VDD.n2259 VSS 0.012131f
C19597 VDD.t1082 VSS 0.034186f
C19598 VDD.n2260 VSS 0.145708f
C19599 VDD.n2261 VSS 0.260606f
C19600 VDD.n2262 VSS 0.012131f
C19601 VDD.n2263 VSS 0.260606f
C19602 VDD.n2264 VSS 0.012131f
C19603 VDD.n2265 VSS 0.385214f
C19604 VDD.n2266 VSS 0.260606f
C19605 VDD.n2267 VSS 0.012131f
C19606 VDD.n2268 VSS 0.260606f
C19607 VDD.n2269 VSS 0.012131f
C19608 VDD.t1094 VSS 0.034186f
C19609 VDD.n2270 VSS 0.145708f
C19610 VDD.n2271 VSS 0.012131f
C19611 VDD.t1093 VSS 0.066856f
C19612 VDD.n2272 VSS 0.154235f
C19613 VDD.n2273 VSS 0.012131f
C19614 VDD.n2274 VSS 0.260606f
C19615 VDD.n2275 VSS 0.012131f
C19616 VDD.n2276 VSS 0.260606f
C19617 VDD.n2277 VSS 0.012131f
C19618 VDD.t2829 VSS 0.034186f
C19619 VDD.n2278 VSS 0.260606f
C19620 VDD.n2279 VSS 0.012131f
C19621 VDD.n2280 VSS 0.232332f
C19622 VDD.n2281 VSS 0.012131f
C19623 VDD.t2454 VSS 0.066856f
C19624 VDD.n2282 VSS 0.154235f
C19625 VDD.t2455 VSS 0.034186f
C19626 VDD.n2283 VSS 0.145708f
C19627 VDD.n2284 VSS 0.012131f
C19628 VDD.n2285 VSS 0.260606f
C19629 VDD.n2286 VSS 0.012131f
C19630 VDD.n2287 VSS 0.260606f
C19631 VDD.n2288 VSS 0.012131f
C19632 VDD.n2289 VSS 0.222498f
C19633 VDD.n2290 VSS 0.012131f
C19634 VDD.t2713 VSS 0.034186f
C19635 VDD.n2291 VSS 0.145708f
C19636 VDD.t2712 VSS 0.066856f
C19637 VDD.n2292 VSS 0.154235f
C19638 VDD.n2293 VSS 0.012131f
C19639 VDD.t2316 VSS 0.034186f
C19640 VDD.t2628 VSS 0.034186f
C19641 VDD.t2195 VSS 0.066856f
C19642 VDD.n2294 VSS 0.164998f
C19643 VDD.t2627 VSS 0.066856f
C19644 VDD.n2295 VSS 0.164998f
C19645 VDD.n2296 VSS 0.274982f
C19646 VDD.t915 VSS 0.066856f
C19647 VDD.t1977 VSS 0.066856f
C19648 VDD.n2297 VSS 0.191511f
C19649 VDD.t916 VSS 0.034186f
C19650 VDD.t1635 VSS 0.066856f
C19651 VDD.t2834 VSS 0.066856f
C19652 VDD.n2298 VSS 0.256005f
C19653 VDD.t1636 VSS 0.025104f
C19654 VDD.t3645 VSS 0.016021f
C19655 VDD.t2643 VSS 0.066856f
C19656 VDD.t3644 VSS 0.066856f
C19657 VDD.n2299 VSS 0.256005f
C19658 VDD.t3951 VSS 0.016021f
C19659 VDD.t3950 VSS 0.066856f
C19660 VDD.t910 VSS 0.066856f
C19661 VDD.n2300 VSS 0.256005f
C19662 VDD.t3653 VSS 0.025104f
C19663 VDD.t2655 VSS 0.066856f
C19664 VDD.t3652 VSS 0.066856f
C19665 VDD.n2301 VSS 0.256005f
C19666 VDD.t1548 VSS 0.066856f
C19667 VDD.t2761 VSS 0.066856f
C19668 VDD.n2302 VSS 0.256005f
C19669 VDD.t1549 VSS 0.025104f
C19670 VDD.t4399 VSS 0.016021f
C19671 VDD.t3332 VSS 0.066856f
C19672 VDD.t4398 VSS 0.066856f
C19673 VDD.n2303 VSS 0.163661f
C19674 VDD.t4689 VSS 0.025104f
C19675 VDD.t4688 VSS 0.066856f
C19676 VDD.t1621 VSS 0.066856f
C19677 VDD.n2304 VSS 0.256005f
C19678 VDD.n2305 VSS 0.10407f
C19679 VDD.t988 VSS 0.066856f
C19680 VDD.t2076 VSS 0.066856f
C19681 VDD.n2306 VSS 0.256005f
C19682 VDD.t989 VSS 0.025104f
C19683 VDD.t3455 VSS 0.016021f
C19684 VDD.t2414 VSS 0.066856f
C19685 VDD.t3454 VSS 0.066856f
C19686 VDD.n2307 VSS 0.256005f
C19687 VDD.t3714 VSS 0.016021f
C19688 VDD.t3713 VSS 0.066856f
C19689 VDD.t644 VSS 0.066856f
C19690 VDD.n2308 VSS 0.256005f
C19691 VDD.t1917 VSS 0.025104f
C19692 VDD.t850 VSS 0.066856f
C19693 VDD.t1916 VSS 0.066856f
C19694 VDD.n2309 VSS 0.256005f
C19695 VDD.n2310 VSS 0.225377f
C19696 VDD.t1953 VSS 0.034186f
C19697 VDD.t1597 VSS 0.034186f
C19698 VDD.n2311 VSS 0.33406f
C19699 VDD.t887 VSS 0.034186f
C19700 VDD.t4665 VSS 0.034186f
C19701 VDD.t4664 VSS 0.066856f
C19702 VDD.t2604 VSS 0.034186f
C19703 VDD.t2181 VSS 0.034186f
C19704 VDD.t2180 VSS 0.066856f
C19705 VDD.t1775 VSS 0.066856f
C19706 VDD.t2167 VSS 0.034186f
C19707 VDD.t1776 VSS 0.034186f
C19708 VDD.n2312 VSS 0.283088f
C19709 VDD.t2218 VSS 0.034186f
C19710 VDD.t1829 VSS 0.034186f
C19711 VDD.t1828 VSS 0.066856f
C19712 VDD.t1465 VSS 0.066856f
C19713 VDD.t1806 VSS 0.034186f
C19714 VDD.t1466 VSS 0.034186f
C19715 VDD.n2313 VSS 0.556001f
C19716 VDD.t1805 VSS 0.066856f
C19717 VDD.n2314 VSS 0.333277f
C19718 VDD.t2217 VSS 0.066856f
C19719 VDD.n2315 VSS 0.333277f
C19720 VDD.n2316 VSS 0.43943f
C19721 VDD.n2317 VSS 1.26071f
C19722 VDD.n2318 VSS 0.280759f
C19723 VDD.t886 VSS 9.19382f
C19724 VDD.n2319 VSS 0.280759f
C19725 VDD.t4093 VSS 0.034186f
C19726 VDD.t3734 VSS 0.034186f
C19727 VDD.n2320 VSS 0.402094f
C19728 VDD.n2321 VSS 0.283088f
C19729 VDD.t995 VSS 0.034186f
C19730 VDD.t588 VSS 0.034186f
C19731 VDD.t586 VSS 0.066856f
C19732 VDD.t4396 VSS 0.066856f
C19733 VDD.t4743 VSS 0.034186f
C19734 VDD.t4397 VSS 0.034186f
C19735 VDD.t1890 VSS 0.066856f
C19736 VDD.t2296 VSS 0.034186f
C19737 VDD.t1891 VSS 0.034186f
C19738 VDD.n2322 VSS 0.225377f
C19739 VDD.t4311 VSS 0.034186f
C19740 VDD.t3981 VSS 0.034186f
C19741 VDD.n2323 VSS 0.333645f
C19742 VDD.t4285 VSS 0.025104f
C19743 VDD.t4284 VSS 0.066856f
C19744 VDD.t2249 VSS 0.066856f
C19745 VDD.n2324 VSS 0.256005f
C19746 VDD.t975 VSS 0.016021f
C19747 VDD.n2325 VSS 0.016021f
C19748 VDD.t3082 VSS 0.066856f
C19749 VDD.t3083 VSS 0.016021f
C19750 VDD.n2326 VSS 0.016021f
C19751 VDD.t1615 VSS 0.066856f
C19752 VDD.t3725 VSS 0.066856f
C19753 VDD.n2327 VSS 0.256005f
C19754 VDD.t2428 VSS 0.025104f
C19755 VDD.t1616 VSS 0.016021f
C19756 VDD.n2328 VSS 0.016021f
C19757 VDD.t4392 VSS 0.066856f
C19758 VDD.t4393 VSS 0.025104f
C19759 VDD.t4005 VSS 0.025104f
C19760 VDD.t4004 VSS 0.066856f
C19761 VDD.t1921 VSS 0.066856f
C19762 VDD.n2329 VSS 0.256005f
C19763 VDD.t4701 VSS 0.016021f
C19764 VDD.n2330 VSS 0.016021f
C19765 VDD.t52 VSS 9.81076f
C19766 VDD.t69 VSS 7.61793f
C19767 VDD.t137 VSS 7.61793f
C19768 VDD.t65 VSS 9.428519f
C19769 VDD.t79 VSS 9.213929f
C19770 VDD.n2331 VSS 0.283109f
C19771 VDD.n2332 VSS 0.283109f
C19772 VDD.t58 VSS 9.81076f
C19773 VDD.t125 VSS 7.61793f
C19774 VDD.t54 VSS 7.61793f
C19775 VDD.t123 VSS 9.428519f
C19776 VDD.t61 VSS 9.428519f
C19777 VDD.t76 VSS 4.02355f
C19778 VDD.n2333 VSS 0.34593f
C19779 VDD.t3532 VSS 0.066856f
C19780 VDD.n2334 VSS 0.016021f
C19781 VDD.t1751 VSS 0.066856f
C19782 VDD.t1736 VSS 0.066856f
C19783 VDD.n2335 VSS 0.414447f
C19784 VDD.t1147 VSS 0.066856f
C19785 VDD.t1134 VSS 0.066856f
C19786 VDD.n2336 VSS 0.414447f
C19787 VDD.t1148 VSS 0.025104f
C19788 VDD.t2618 VSS 0.016021f
C19789 VDD.t2633 VSS 0.066856f
C19790 VDD.t2617 VSS 0.066856f
C19791 VDD.n2337 VSS 0.414447f
C19792 VDD.t3927 VSS 0.016021f
C19793 VDD.t3926 VSS 0.066856f
C19794 VDD.t3908 VSS 0.066856f
C19795 VDD.n2338 VSS 0.414447f
C19796 VDD.t1025 VSS 0.025104f
C19797 VDD.t1036 VSS 0.066856f
C19798 VDD.t1024 VSS 0.066856f
C19799 VDD.n2339 VSS 0.414447f
C19800 VDD.t1073 VSS 0.066856f
C19801 VDD.t1063 VSS 0.066856f
C19802 VDD.n2340 VSS 0.414447f
C19803 VDD.t1074 VSS 0.034186f
C19804 VDD.t2806 VSS 0.034186f
C19805 VDD.t2453 VSS 0.034186f
C19806 VDD.n2341 VSS 0.556001f
C19807 VDD.n2342 VSS 0.369079f
C19808 VDD.t3980 VSS 0.066856f
C19809 VDD.t4310 VSS 0.066856f
C19810 VDD.n2343 VSS 0.58882f
C19811 VDD.t2019 VSS 0.034186f
C19812 VDD.t1658 VSS 0.034186f
C19813 VDD.n2344 VSS 0.571765f
C19814 VDD.t1657 VSS 0.066856f
C19815 VDD.t2018 VSS 0.066856f
C19816 VDD.n2345 VSS 0.333277f
C19817 VDD.t1286 VSS 0.066856f
C19818 VDD.t1641 VSS 0.066856f
C19819 VDD.n2346 VSS 0.333277f
C19820 VDD.t1642 VSS 0.034186f
C19821 VDD.t1287 VSS 0.034186f
C19822 VDD.n2347 VSS 0.402094f
C19823 VDD.n2348 VSS 0.279865f
C19824 VDD.n2349 VSS 0.280759f
C19825 VDD.n2350 VSS 0.183291f
C19826 VDD.t81 VSS 9.213929f
C19827 VDD.n2351 VSS 0.283109f
C19828 VDD.n2352 VSS 0.283109f
C19829 VDD.n2353 VSS 0.283109f
C19830 VDD.t404 VSS 3.66626f
C19831 VDD.t572 VSS 3.43571f
C19832 VDD.n2354 VSS 1.55371f
C19833 VDD.n2355 VSS 1.55371f
C19834 VDD.t913 VSS 3.43571f
C19835 VDD.t15 VSS 3.66626f
C19836 VDD.t41 VSS 1.73916f
C19837 VDD.t19 VSS 3.52342f
C19838 VDD.t21 VSS 2.53105f
C19839 VDD.n2356 VSS 4.61542f
C19840 VDD.t587 VSS 8.89876f
C19841 VDD.t73 VSS 9.81076f
C19842 VDD.t118 VSS 7.61793f
C19843 VDD.t56 VSS 7.61793f
C19844 VDD.t50 VSS 9.428519f
C19845 VDD.t67 VSS 9.428519f
C19846 VDD.t99 VSS 4.02355f
C19847 VDD.n2357 VSS 0.279865f
C19848 VDD.t2452 VSS 0.066856f
C19849 VDD.t2805 VSS 0.066856f
C19850 VDD.n2358 VSS 0.333277f
C19851 VDD.t2006 VSS 0.066856f
C19852 VDD.t2435 VSS 0.066856f
C19853 VDD.n2359 VSS 0.333277f
C19854 VDD.t2436 VSS 0.034186f
C19855 VDD.t2007 VSS 0.034186f
C19856 VDD.n2360 VSS 0.402094f
C19857 VDD.t2689 VSS 0.034186f
C19858 VDD.t2310 VSS 0.034186f
C19859 VDD.t2309 VSS 0.066856f
C19860 VDD.t1881 VSS 0.066856f
C19861 VDD.t2275 VSS 0.034186f
C19862 VDD.t1882 VSS 0.034186f
C19863 VDD.t1596 VSS 0.066856f
C19864 VDD.t1952 VSS 0.066856f
C19865 VDD.n2361 VSS 0.58882f
C19866 VDD.n2362 VSS 0.571765f
C19867 VDD.t2274 VSS 0.066856f
C19868 VDD.n2363 VSS 0.333277f
C19869 VDD.t2688 VSS 0.066856f
C19870 VDD.n2364 VSS 0.333277f
C19871 VDD.n2365 VSS 0.43943f
C19872 VDD.n2366 VSS 0.532659f
C19873 VDD.n2367 VSS 0.283088f
C19874 VDD.n2368 VSS 0.279865f
C19875 VDD.n2369 VSS 0.280759f
C19876 VDD.n2370 VSS 0.096993f
C19877 VDD.t2651 VSS 0.066856f
C19878 VDD.n2371 VSS 0.126716f
C19879 VDD.t726 VSS 0.016021f
C19880 VDD.t3150 VSS 0.066856f
C19881 VDD.n2372 VSS 0.126716f
C19882 VDD.t1315 VSS 0.016021f
C19883 VDD.t4554 VSS 0.066856f
C19884 VDD.n2373 VSS 0.126716f
C19885 VDD.t3271 VSS 0.025104f
C19886 VDD.t3270 VSS 0.066856f
C19887 VDD.n2374 VSS 0.057673f
C19888 VDD.n2375 VSS 0.05157f
C19889 VDD.n2376 VSS 0.283978f
C19890 VDD.t185 VSS 0.008011f
C19891 VDD.t233 VSS 0.008011f
C19892 VDD.n2377 VSS 0.04401f
C19893 VDD.t72 VSS 0.008011f
C19894 VDD.t154 VSS 0.008011f
C19895 VDD.n2378 VSS 0.029389f
C19896 VDD.n2379 VSS 0.144542f
C19897 VDD.t51 VSS 0.008011f
C19898 VDD.t165 VSS 0.008011f
C19899 VDD.n2380 VSS 0.029389f
C19900 VDD.n2381 VSS 0.102512f
C19901 VDD.t214 VSS 0.008011f
C19902 VDD.t285 VSS 0.008011f
C19903 VDD.n2382 VSS 0.029389f
C19904 VDD.n2383 VSS 0.041173f
C19905 VDD.n2384 VSS 0.041824f
C19906 VDD.t3589 VSS 0.066856f
C19907 VDD.n2385 VSS 0.057673f
C19908 VDD.t2897 VSS 0.034186f
C19909 VDD.t4459 VSS 0.034186f
C19910 VDD.t4120 VSS 0.066856f
C19911 VDD.n2386 VSS 0.164998f
C19912 VDD.t4458 VSS 0.066856f
C19913 VDD.n2387 VSS 0.164998f
C19914 VDD.n2388 VSS 0.282774f
C19915 VDD.t2896 VSS 0.066856f
C19916 VDD.n2389 VSS 0.291301f
C19917 VDD.n2390 VSS 0.277083f
C19918 VDD.t4475 VSS 0.016021f
C19919 VDD.t1689 VSS 0.066856f
C19920 VDD.n2391 VSS 0.126716f
C19921 VDD.t4479 VSS 0.025104f
C19922 VDD.t3514 VSS 0.066856f
C19923 VDD.n2392 VSS 0.126716f
C19924 VDD.t1096 VSS 0.016021f
C19925 VDD.t2556 VSS 0.066856f
C19926 VDD.n2393 VSS 0.126716f
C19927 VDD.t2976 VSS 0.066856f
C19928 VDD.n2394 VSS 0.126716f
C19929 VDD.t4269 VSS 0.016021f
C19930 VDD.t1463 VSS 0.066856f
C19931 VDD.n2395 VSS 0.126716f
C19932 VDD.t2845 VSS 0.025104f
C19933 VDD.n2396 VSS 0.105419f
C19934 VDD.t2875 VSS 0.034186f
C19935 VDD.t2529 VSS 0.034186f
C19936 VDD.t2528 VSS 0.066856f
C19937 VDD.t4427 VSS 0.034186f
C19938 VDD.t4115 VSS 0.034186f
C19939 VDD.t4114 VSS 0.066856f
C19940 VDD.t3733 VSS 0.066856f
C19941 VDD.t4092 VSS 0.066856f
C19942 VDD.n2397 VSS 0.333277f
C19943 VDD.t4426 VSS 0.066856f
C19944 VDD.n2398 VSS 0.333277f
C19945 VDD.n2399 VSS 0.571765f
C19946 VDD.t2874 VSS 0.066856f
C19947 VDD.n2400 VSS 0.58882f
C19948 VDD.n2401 VSS 0.172271f
C19949 VDD.n2402 VSS 0.437712f
C19950 VDD.n2403 VSS 0.111391f
C19951 VDD.t2844 VSS 0.066856f
C19952 VDD.n2404 VSS 0.111632f
C19953 VDD.n2405 VSS 0.306702f
C19954 VDD.t1007 VSS 0.066856f
C19955 VDD.n2406 VSS 0.08105f
C19956 VDD.t4244 VSS 0.066856f
C19957 VDD.n2407 VSS 0.126716f
C19958 VDD.n2408 VSS 0.104062f
C19959 VDD.n2409 VSS 0.051804f
C19960 VDD.n2410 VSS 0.151757f
C19961 VDD.n2412 VSS 0.012131f
C19962 VDD.n2413 VSS 0.012131f
C19963 VDD.n2414 VSS 0.012131f
C19964 VDD.n2415 VSS 0.012131f
C19965 VDD.n2416 VSS 0.012131f
C19966 VDD.n2417 VSS 0.012131f
C19967 VDD.n2418 VSS 0.012131f
C19968 VDD.n2419 VSS 0.012131f
C19969 VDD.n2420 VSS 0.012131f
C19970 VDD.n2421 VSS 0.012131f
C19971 VDD.n2422 VSS 0.012131f
C19972 VDD.n2423 VSS 0.012131f
C19973 VDD.n2425 VSS 0.012131f
C19974 VDD.n2426 VSS 0.012131f
C19975 VDD.n2427 VSS 0.012131f
C19976 VDD.n2428 VSS 0.012131f
C19977 VDD.n2429 VSS 0.012131f
C19978 VDD.n2430 VSS 0.012131f
C19979 VDD.n2431 VSS 0.012131f
C19980 VDD.n2432 VSS 0.012131f
C19981 VDD.n2433 VSS 0.012131f
C19982 VDD.n2434 VSS 0.012131f
C19983 VDD.n2435 VSS 0.012131f
C19984 VDD.n2436 VSS 0.012131f
C19985 VDD.n2437 VSS 0.012131f
C19986 VDD.n2438 VSS 0.012131f
C19987 VDD.n2439 VSS 0.012131f
C19988 VDD.n2440 VSS 0.012131f
C19989 VDD.n2441 VSS 0.012131f
C19990 VDD.n2442 VSS 0.012131f
C19991 VDD.n2443 VSS 0.012131f
C19992 VDD.n2444 VSS 0.012131f
C19993 VDD.n2445 VSS 0.012131f
C19994 VDD.n2446 VSS 0.012131f
C19995 VDD.n2447 VSS 0.012131f
C19996 VDD.n2448 VSS 0.012131f
C19997 VDD.n2449 VSS 0.012131f
C19998 VDD.n2450 VSS 0.012131f
C19999 VDD.n2451 VSS 0.012131f
C20000 VDD.n2452 VSS 0.012131f
C20001 VDD.n2453 VSS 0.012131f
C20002 VDD.n2454 VSS 0.012131f
C20003 VDD.n2455 VSS 0.012131f
C20004 VDD.n2456 VSS 0.012131f
C20005 VDD.n2457 VSS 0.012131f
C20006 VDD.n2458 VSS 0.012131f
C20007 VDD.n2459 VSS 0.012131f
C20008 VDD.n2460 VSS 0.012131f
C20009 VDD.n2461 VSS 0.012131f
C20010 VDD.n2462 VSS 0.012131f
C20011 VDD.n2463 VSS 0.012131f
C20012 VDD.n2464 VSS 0.012131f
C20013 VDD.n2465 VSS 0.012131f
C20014 VDD.n2466 VSS 0.012131f
C20015 VDD.n2467 VSS 0.012131f
C20016 VDD.n2468 VSS 0.012131f
C20017 VDD.n2469 VSS 0.012131f
C20018 VDD.n2470 VSS 0.012131f
C20019 VDD.n2471 VSS 0.012131f
C20020 VDD.n2472 VSS 0.012131f
C20021 VDD.n2473 VSS 0.012131f
C20022 VDD.n2474 VSS 0.012131f
C20023 VDD.n2475 VSS 0.012131f
C20024 VDD.n2476 VSS 0.012131f
C20025 VDD.n2477 VSS 0.012131f
C20026 VDD.n2478 VSS 0.012131f
C20027 VDD.n2479 VSS 0.012131f
C20028 VDD.n2480 VSS 0.012131f
C20029 VDD.n2481 VSS 0.012131f
C20030 VDD.n2482 VSS 0.012131f
C20031 VDD.n2483 VSS 0.012131f
C20032 VDD.n2484 VSS 0.012131f
C20033 VDD.n2485 VSS 0.012131f
C20034 VDD.n2486 VSS 0.012131f
C20035 VDD.n2487 VSS 0.012131f
C20036 VDD.n2488 VSS 0.012131f
C20037 VDD.n2489 VSS 0.012131f
C20038 VDD.n2490 VSS 0.012131f
C20039 VDD.n2491 VSS 0.012131f
C20040 VDD.n2492 VSS 0.012131f
C20041 VDD.n2493 VSS 0.012131f
C20042 VDD.n2494 VSS 0.012131f
C20043 VDD.n2495 VSS 0.012131f
C20044 VDD.n2496 VSS 0.012131f
C20045 VDD.n2497 VSS 0.012131f
C20046 VDD.n2498 VSS 0.012131f
C20047 VDD.n2499 VSS 0.012131f
C20048 VDD.n2500 VSS 0.012131f
C20049 VDD.n2501 VSS 0.012131f
C20050 VDD.n2502 VSS 0.012131f
C20051 VDD.n2503 VSS 0.012131f
C20052 VDD.n2504 VSS 0.012131f
C20053 VDD.n2505 VSS 0.012131f
C20054 VDD.n2506 VSS 0.012131f
C20055 VDD.n2507 VSS 0.012131f
C20056 VDD.n2508 VSS 0.012131f
C20057 VDD.n2509 VSS 0.012131f
C20058 VDD.n2510 VSS 0.012131f
C20059 VDD.n2511 VSS 0.012131f
C20060 VDD.n2512 VSS 0.012131f
C20061 VDD.n2513 VSS 0.012131f
C20062 VDD.n2514 VSS 0.012131f
C20063 VDD.n2515 VSS 0.012131f
C20064 VDD.n2516 VSS 0.012131f
C20065 VDD.n2517 VSS 0.012131f
C20066 VDD.n2518 VSS 0.012131f
C20067 VDD.n2519 VSS 0.012131f
C20068 VDD.n2520 VSS 0.012131f
C20069 VDD.n2521 VSS 0.012131f
C20070 VDD.n2522 VSS 0.012131f
C20071 VDD.n2523 VSS 0.012131f
C20072 VDD.n2524 VSS 0.012131f
C20073 VDD.n2525 VSS 0.012131f
C20074 VDD.n2526 VSS 0.012131f
C20075 VDD.n2527 VSS 0.012131f
C20076 VDD.n2528 VSS 0.012131f
C20077 VDD.n2529 VSS 0.012131f
C20078 VDD.n2530 VSS 0.012131f
C20079 VDD.n2531 VSS 0.012131f
C20080 VDD.n2532 VSS 0.012131f
C20081 VDD.n2533 VSS 0.012131f
C20082 VDD.n2534 VSS 0.012131f
C20083 VDD.n2535 VSS 0.012131f
C20084 VDD.n2536 VSS 0.012131f
C20085 VDD.n2537 VSS 0.012131f
C20086 VDD.n2538 VSS 0.012131f
C20087 VDD.n2539 VSS 0.012131f
C20088 VDD.n2540 VSS 0.012131f
C20089 VDD.n2541 VSS 0.012131f
C20090 VDD.n2542 VSS 0.012131f
C20091 VDD.n2543 VSS 0.012131f
C20092 VDD.n2544 VSS 0.012131f
C20093 VDD.n2545 VSS 0.012131f
C20094 VDD.n2546 VSS 0.012131f
C20095 VDD.n2547 VSS 0.012131f
C20096 VDD.n2548 VSS 0.012131f
C20097 VDD.n2549 VSS 0.012131f
C20098 VDD.n2550 VSS 0.012131f
C20099 VDD.n2551 VSS 0.012131f
C20100 VDD.n2552 VSS 0.012131f
C20101 VDD.n2553 VSS 0.012131f
C20102 VDD.n2554 VSS 0.012131f
C20103 VDD.n2555 VSS 0.012131f
C20104 VDD.n2556 VSS 0.012131f
C20105 VDD.n2557 VSS 0.012131f
C20106 VDD.n2558 VSS 0.012131f
C20107 VDD.n2559 VSS 0.012131f
C20108 VDD.n2560 VSS 0.012131f
C20109 VDD.n2561 VSS 0.012131f
C20110 VDD.n2562 VSS 0.012131f
C20111 VDD.n2563 VSS 0.012131f
C20112 VDD.n2564 VSS 0.012131f
C20113 VDD.n2565 VSS 0.012131f
C20114 VDD.n2566 VSS 0.012131f
C20115 VDD.n2567 VSS 0.012131f
C20116 VDD.n2568 VSS 0.012131f
C20117 VDD.n2569 VSS 0.012131f
C20118 VDD.n2570 VSS 0.012131f
C20119 VDD.n2571 VSS 0.012131f
C20120 VDD.n2572 VSS 0.012131f
C20121 VDD.n2573 VSS 0.012131f
C20122 VDD.n2574 VSS 0.012131f
C20123 VDD.n2575 VSS 0.012131f
C20124 VDD.n2576 VSS 0.012131f
C20125 VDD.n2577 VSS 0.012131f
C20126 VDD.n2578 VSS 0.012131f
C20127 VDD.n2579 VSS 0.012131f
C20128 VDD.n2580 VSS 0.012131f
C20129 VDD.n2581 VSS 0.012131f
C20130 VDD.n2582 VSS 0.012131f
C20131 VDD.n2583 VSS 0.012131f
C20132 VDD.n2584 VSS 0.012131f
C20133 VDD.n2585 VSS 0.012131f
C20134 VDD.n2586 VSS 0.012131f
C20135 VDD.n2587 VSS 0.012131f
C20136 VDD.n2588 VSS 0.012131f
C20137 VDD.n2589 VSS 0.012131f
C20138 VDD.n2590 VSS 0.012131f
C20139 VDD.n2591 VSS 0.012131f
C20140 VDD.n2592 VSS 0.012131f
C20141 VDD.n2593 VSS 0.012131f
C20142 VDD.n2594 VSS 0.012131f
C20143 VDD.n2595 VSS 0.012131f
C20144 VDD.n2596 VSS 0.012131f
C20145 VDD.n2597 VSS 0.012131f
C20146 VDD.n2598 VSS 0.012131f
C20147 VDD.n2599 VSS 0.012131f
C20148 VDD.n2600 VSS 0.012131f
C20149 VDD.n2601 VSS 0.012131f
C20150 VDD.n2602 VSS 0.012131f
C20151 VDD.n2603 VSS 0.012131f
C20152 VDD.n2604 VSS 0.012131f
C20153 VDD.n2605 VSS 0.012131f
C20154 VDD.n2606 VSS 0.012131f
C20155 VDD.n2607 VSS 0.012131f
C20156 VDD.n2608 VSS 0.012131f
C20157 VDD.n2609 VSS 0.012131f
C20158 VDD.n2610 VSS 0.012131f
C20159 VDD.n2611 VSS 0.012131f
C20160 VDD.n2612 VSS 0.012131f
C20161 VDD.n2613 VSS 0.012131f
C20162 VDD.n2614 VSS 0.012131f
C20163 VDD.n2615 VSS 0.012131f
C20164 VDD.n2616 VSS 0.012131f
C20165 VDD.n2617 VSS 0.012131f
C20166 VDD.n2618 VSS 0.012131f
C20167 VDD.n2619 VSS 0.012131f
C20168 VDD.n2620 VSS 0.012131f
C20169 VDD.n2621 VSS 0.012131f
C20170 VDD.n2622 VSS 0.012131f
C20171 VDD.n2623 VSS 0.012131f
C20172 VDD.n2624 VSS 0.012131f
C20173 VDD.n2625 VSS 0.012131f
C20174 VDD.n2626 VSS 0.012131f
C20175 VDD.n2627 VSS 0.012131f
C20176 VDD.n2628 VSS 0.012131f
C20177 VDD.n2629 VSS 0.012131f
C20178 VDD.n2630 VSS 0.012131f
C20179 VDD.n2631 VSS 0.012131f
C20180 VDD.n2632 VSS 0.012131f
C20181 VDD.n2633 VSS 0.012131f
C20182 VDD.n2634 VSS 0.012131f
C20183 VDD.n2635 VSS 0.012131f
C20184 VDD.n2636 VSS 0.012131f
C20185 VDD.n2637 VSS 0.012131f
C20186 VDD.n2638 VSS 0.012131f
C20187 VDD.n2639 VSS 0.012131f
C20188 VDD.n2640 VSS 0.012131f
C20189 VDD.n2641 VSS 0.012131f
C20190 VDD.n2642 VSS 0.012131f
C20191 VDD.n2643 VSS 0.012131f
C20192 VDD.n2644 VSS 0.012131f
C20193 VDD.n2645 VSS 0.012131f
C20194 VDD.n2646 VSS 0.012131f
C20195 VDD.n2647 VSS 0.012131f
C20196 VDD.n2648 VSS 0.012131f
C20197 VDD.n2649 VSS 0.012131f
C20198 VDD.n2650 VSS 0.012131f
C20199 VDD.n2651 VSS 0.012131f
C20200 VDD.n2652 VSS 0.012131f
C20201 VDD.n2653 VSS 0.012131f
C20202 VDD.n2654 VSS 0.012131f
C20203 VDD.n2655 VSS 0.012131f
C20204 VDD.n2656 VSS 0.012131f
C20205 VDD.n2657 VSS 0.012131f
C20206 VDD.n2658 VSS 0.012131f
C20207 VDD.n2659 VSS 0.012131f
C20208 VDD.n2660 VSS 0.012131f
C20209 VDD.n2661 VSS 0.012131f
C20210 VDD.n2662 VSS 0.012131f
C20211 VDD.n2663 VSS 0.012131f
C20212 VDD.n2664 VSS 0.012131f
C20213 VDD.n2665 VSS 0.012131f
C20214 VDD.n2666 VSS 0.012131f
C20215 VDD.n2667 VSS 0.012131f
C20216 VDD.n2668 VSS 0.012131f
C20217 VDD.n2669 VSS 0.012131f
C20218 VDD.n2670 VSS 0.012131f
C20219 VDD.n2671 VSS 0.012131f
C20220 VDD.n2672 VSS 0.012131f
C20221 VDD.n2673 VSS 0.012131f
C20222 VDD.n2674 VSS 0.012131f
C20223 VDD.n2675 VSS 0.012131f
C20224 VDD.n2676 VSS 0.012131f
C20225 VDD.n2677 VSS 0.012131f
C20226 VDD.n2678 VSS 0.012131f
C20227 VDD.n2679 VSS 0.012131f
C20228 VDD.n2680 VSS 0.012131f
C20229 VDD.n2681 VSS 0.012131f
C20230 VDD.n2682 VSS 0.012131f
C20231 VDD.n2683 VSS 0.012131f
C20232 VDD.n2684 VSS 0.012131f
C20233 VDD.n2685 VSS 0.012131f
C20234 VDD.n2686 VSS 0.012131f
C20235 VDD.n2687 VSS 0.012131f
C20236 VDD.n2688 VSS 0.012131f
C20237 VDD.n2689 VSS 0.012131f
C20238 VDD.n2690 VSS 0.012131f
C20239 VDD.n2691 VSS 0.012131f
C20240 VDD.n2692 VSS 0.012131f
C20241 VDD.n2693 VSS 0.012131f
C20242 VDD.n2694 VSS 0.012131f
C20243 VDD.n2695 VSS 0.012131f
C20244 VDD.n2696 VSS 0.012131f
C20245 VDD.n2697 VSS 0.012131f
C20246 VDD.n2698 VSS 0.012131f
C20247 VDD.n2699 VSS 0.012131f
C20248 VDD.n2700 VSS 0.012131f
C20249 VDD.n2701 VSS 0.012131f
C20250 VDD.n2702 VSS 0.012131f
C20251 VDD.n2703 VSS 0.012131f
C20252 VDD.n2704 VSS 0.012131f
C20253 VDD.n2705 VSS 0.012131f
C20254 VDD.n2706 VSS 0.012131f
C20255 VDD.n2707 VSS 0.012131f
C20256 VDD.n2708 VSS 0.012131f
C20257 VDD.n2709 VSS 0.012131f
C20258 VDD.n2710 VSS 0.012131f
C20259 VDD.n2711 VSS 0.012131f
C20260 VDD.n2712 VSS 0.012131f
C20261 VDD.n2713 VSS 0.012131f
C20262 VDD.n2714 VSS 0.012131f
C20263 VDD.n2715 VSS 0.012131f
C20264 VDD.n2716 VSS 0.012131f
C20265 VDD.n2717 VSS 0.012131f
C20266 VDD.n2718 VSS 0.012131f
C20267 VDD.n2719 VSS 0.012131f
C20268 VDD.n2720 VSS 0.012131f
C20269 VDD.n2721 VSS 0.012131f
C20270 VDD.n2722 VSS 0.012131f
C20271 VDD.n2723 VSS 0.012131f
C20272 VDD.n2724 VSS 0.012131f
C20273 VDD.n2725 VSS 0.012131f
C20274 VDD.n2726 VSS 0.012131f
C20275 VDD.n2727 VSS 0.012131f
C20276 VDD.n2728 VSS 0.012131f
C20277 VDD.n2729 VSS 0.012131f
C20278 VDD.n2730 VSS 0.012131f
C20279 VDD.n2731 VSS 0.012131f
C20280 VDD.n2732 VSS 0.012131f
C20281 VDD.n2733 VSS 0.012131f
C20282 VDD.n2734 VSS 0.012131f
C20283 VDD.n2735 VSS 0.012131f
C20284 VDD.n2736 VSS 0.012131f
C20285 VDD.n2737 VSS 0.012131f
C20286 VDD.n2738 VSS 0.012131f
C20287 VDD.n2739 VSS 0.012131f
C20288 VDD.n2740 VSS 0.012131f
C20289 VDD.n2741 VSS 0.012131f
C20290 VDD.n2742 VSS 0.012131f
C20291 VDD.n2743 VSS 0.012131f
C20292 VDD.n2744 VSS 0.012131f
C20293 VDD.n2745 VSS 0.026818f
C20294 VDD.n2746 VSS 0.012131f
C20295 VDD.n2747 VSS 0.012131f
C20296 VDD.n2748 VSS 0.012131f
C20297 VDD.n2749 VSS 0.012131f
C20298 VDD.n2750 VSS 0.012131f
C20299 VDD.n2751 VSS 0.012131f
C20300 VDD.n2752 VSS 0.012131f
C20301 VDD.n2753 VSS 0.012131f
C20302 VDD.n2754 VSS 0.012131f
C20303 VDD.n2755 VSS 0.012131f
C20304 VDD.n2756 VSS 0.012131f
C20305 VDD.n2757 VSS 0.012131f
C20306 VDD.n2758 VSS 0.012131f
C20307 VDD.n2759 VSS 0.012131f
C20308 VDD.n2760 VSS 0.012131f
C20309 VDD.n2761 VSS 0.012131f
C20310 VDD.n2762 VSS 0.012131f
C20311 VDD.n2763 VSS 0.012131f
C20312 VDD.n2764 VSS 0.012131f
C20313 VDD.n2765 VSS 0.012131f
C20314 VDD.n2766 VSS 0.012131f
C20315 VDD.n2767 VSS 0.012131f
C20316 VDD.n2768 VSS 0.012131f
C20317 VDD.n2769 VSS 0.012131f
C20318 VDD.n2770 VSS 0.012131f
C20319 VDD.n2771 VSS 0.012131f
C20320 VDD.n2772 VSS 0.012131f
C20321 VDD.n2773 VSS 0.012131f
C20322 VDD.n2774 VSS 0.012131f
C20323 VDD.n2775 VSS 0.012131f
C20324 VDD.n2776 VSS 0.012131f
C20325 VDD.n2777 VSS 0.012131f
C20326 VDD.n2778 VSS 0.012131f
C20327 VDD.n2779 VSS 0.012131f
C20328 VDD.n2780 VSS 0.012131f
C20329 VDD.n2781 VSS 0.012131f
C20330 VDD.n2782 VSS 0.012131f
C20331 VDD.n2783 VSS 0.012131f
C20332 VDD.n2784 VSS 0.012131f
C20333 VDD.n2785 VSS 0.012131f
C20334 VDD.n2786 VSS 0.012131f
C20335 VDD.n2787 VSS 0.012131f
C20336 VDD.n2788 VSS 0.012131f
C20337 VDD.n2789 VSS 0.012131f
C20338 VDD.n2790 VSS 0.012131f
C20339 VDD.n2791 VSS 0.012131f
C20340 VDD.n2792 VSS 0.012131f
C20341 VDD.n2793 VSS 0.012131f
C20342 VDD.n2794 VSS 0.012131f
C20343 VDD.n2795 VSS 0.012131f
C20344 VDD.n2796 VSS 0.012131f
C20345 VDD.n2797 VSS 0.012131f
C20346 VDD.n2798 VSS 0.012131f
C20347 VDD.n2799 VSS 0.012131f
C20348 VDD.n2800 VSS 0.012131f
C20349 VDD.n2801 VSS 0.012131f
C20350 VDD.n2802 VSS 0.012131f
C20351 VDD.n2803 VSS 0.012131f
C20352 VDD.n2804 VSS 0.012131f
C20353 VDD.n2805 VSS 0.012131f
C20354 VDD.n2806 VSS 0.012131f
C20355 VDD.n2807 VSS 0.012131f
C20356 VDD.n2808 VSS 0.012131f
C20357 VDD.n2809 VSS 0.012131f
C20358 VDD.n2810 VSS 0.012131f
C20359 VDD.n2811 VSS 0.012131f
C20360 VDD.n2812 VSS 0.012131f
C20361 VDD.n2813 VSS 0.012131f
C20362 VDD.n2814 VSS 0.012131f
C20363 VDD.n2815 VSS 0.012131f
C20364 VDD.n2816 VSS 0.012131f
C20365 VDD.n2817 VSS 0.012131f
C20366 VDD.n2818 VSS 0.012131f
C20367 VDD.n2819 VSS 0.012131f
C20368 VDD.n2820 VSS 0.012131f
C20369 VDD.n2821 VSS 0.012131f
C20370 VDD.n2822 VSS 0.012131f
C20371 VDD.n2823 VSS 0.012131f
C20372 VDD.n2824 VSS 0.012131f
C20373 VDD.n2825 VSS 0.012131f
C20374 VDD.n2826 VSS 0.012131f
C20375 VDD.n2827 VSS 0.012131f
C20376 VDD.n2828 VSS 0.012131f
C20377 VDD.n2829 VSS 0.012131f
C20378 VDD.n2830 VSS 0.012131f
C20379 VDD.n2831 VSS 0.012131f
C20380 VDD.n2832 VSS 0.012131f
C20381 VDD.n2833 VSS 0.012131f
C20382 VDD.n2834 VSS 0.012131f
C20383 VDD.n2835 VSS 0.012131f
C20384 VDD.n2836 VSS 0.012131f
C20385 VDD.n2837 VSS 0.012131f
C20386 VDD.n2838 VSS 0.012131f
C20387 VDD.n2839 VSS 0.012131f
C20388 VDD.n2840 VSS 0.012131f
C20389 VDD.n2841 VSS 0.012131f
C20390 VDD.n2842 VSS 0.012131f
C20391 VDD.n2843 VSS 0.012131f
C20392 VDD.n2844 VSS 0.012131f
C20393 VDD.n2845 VSS 0.012131f
C20394 VDD.n2846 VSS 0.012131f
C20395 VDD.n2847 VSS 0.012131f
C20396 VDD.n2848 VSS 0.012131f
C20397 VDD.n2849 VSS 0.012131f
C20398 VDD.n2850 VSS 0.012131f
C20399 VDD.n2851 VSS 0.012131f
C20400 VDD.n2852 VSS 0.012131f
C20401 VDD.n2853 VSS 0.012131f
C20402 VDD.n2854 VSS 0.012131f
C20403 VDD.n2855 VSS 0.012131f
C20404 VDD.n2856 VSS 0.012131f
C20405 VDD.n2857 VSS 0.012131f
C20406 VDD.n2858 VSS 0.012131f
C20407 VDD.n2859 VSS 0.012131f
C20408 VDD.n2860 VSS 0.012131f
C20409 VDD.n2861 VSS 0.012131f
C20410 VDD.n2862 VSS 0.012131f
C20411 VDD.n2863 VSS 0.012131f
C20412 VDD.n2864 VSS 0.012131f
C20413 VDD.n2865 VSS 0.012131f
C20414 VDD.n2866 VSS 0.012131f
C20415 VDD.n2867 VSS 0.012131f
C20416 VDD.n2868 VSS 0.012131f
C20417 VDD.n2869 VSS 0.012131f
C20418 VDD.n2870 VSS 0.012131f
C20419 VDD.n2871 VSS 0.012131f
C20420 VDD.n2872 VSS 0.012131f
C20421 VDD.n2873 VSS 0.012131f
C20422 VDD.n2874 VSS 0.012131f
C20423 VDD.n2875 VSS 0.012131f
C20424 VDD.n2876 VSS 0.012131f
C20425 VDD.n2877 VSS 0.012131f
C20426 VDD.n2878 VSS 0.012131f
C20427 VDD.n2879 VSS 0.012131f
C20428 VDD.n2880 VSS 0.012131f
C20429 VDD.n2881 VSS 0.012131f
C20430 VDD.n2882 VSS 0.012131f
C20431 VDD.n2883 VSS 0.012131f
C20432 VDD.n2884 VSS 0.012131f
C20433 VDD.n2885 VSS 0.012131f
C20434 VDD.n2886 VSS 0.012131f
C20435 VDD.n2887 VSS 0.012131f
C20436 VDD.n2888 VSS 0.012131f
C20437 VDD.n2889 VSS 0.012131f
C20438 VDD.n2890 VSS 0.012131f
C20439 VDD.n2891 VSS 0.012131f
C20440 VDD.n2892 VSS 0.012131f
C20441 VDD.n2893 VSS 0.012131f
C20442 VDD.n2894 VSS 0.012131f
C20443 VDD.n2895 VSS 0.012131f
C20444 VDD.n2896 VSS 0.012131f
C20445 VDD.n2897 VSS 0.012131f
C20446 VDD.n2898 VSS 0.012131f
C20447 VDD.n2899 VSS 0.012131f
C20448 VDD.n2900 VSS 0.012131f
C20449 VDD.n2901 VSS 0.012131f
C20450 VDD.n2902 VSS 0.012131f
C20451 VDD.n2903 VSS 0.012131f
C20452 VDD.n2904 VSS 0.012131f
C20453 VDD.n2905 VSS 0.012131f
C20454 VDD.n2906 VSS 0.012131f
C20455 VDD.n2907 VSS 0.012131f
C20456 VDD.n2908 VSS 0.012131f
C20457 VDD.n2909 VSS 0.012131f
C20458 VDD.n2910 VSS 0.012131f
C20459 VDD.n2911 VSS 0.012131f
C20460 VDD.n2912 VSS 0.012131f
C20461 VDD.n2913 VSS 0.012131f
C20462 VDD.n2914 VSS 0.012131f
C20463 VDD.n2915 VSS 0.012131f
C20464 VDD.n2916 VSS 0.012131f
C20465 VDD.n2917 VSS 0.012131f
C20466 VDD.n2918 VSS 0.012131f
C20467 VDD.n2919 VSS 0.012131f
C20468 VDD.n2920 VSS 0.012131f
C20469 VDD.n2921 VSS 0.012131f
C20470 VDD.n2922 VSS 0.012131f
C20471 VDD.n2923 VSS 0.012131f
C20472 VDD.n2924 VSS 0.012131f
C20473 VDD.n2925 VSS 0.012131f
C20474 VDD.n2926 VSS 0.012131f
C20475 VDD.n2927 VSS 0.012131f
C20476 VDD.n2928 VSS 0.012131f
C20477 VDD.n2929 VSS 0.012131f
C20478 VDD.n2930 VSS 0.012131f
C20479 VDD.n2931 VSS 0.012131f
C20480 VDD.n2932 VSS 0.012131f
C20481 VDD.n2933 VSS 0.012131f
C20482 VDD.n2934 VSS 0.012131f
C20483 VDD.n2935 VSS 0.012131f
C20484 VDD.n2936 VSS 0.012131f
C20485 VDD.n2937 VSS 0.012131f
C20486 VDD.n2938 VSS 0.012131f
C20487 VDD.n2939 VSS 0.012131f
C20488 VDD.n2940 VSS 0.012131f
C20489 VDD.n2941 VSS 0.012131f
C20490 VDD.n2942 VSS 0.012131f
C20491 VDD.n2943 VSS 0.012131f
C20492 VDD.n2944 VSS 0.012131f
C20493 VDD.n2945 VSS 0.012131f
C20494 VDD.n2946 VSS 0.012131f
C20495 VDD.n2947 VSS 0.012131f
C20496 VDD.n2948 VSS 0.012131f
C20497 VDD.n2949 VSS 0.012131f
C20498 VDD.n2950 VSS 0.012131f
C20499 VDD.n2951 VSS 0.012131f
C20500 VDD.n2952 VSS 0.012131f
C20501 VDD.n2953 VSS 0.012131f
C20502 VDD.n2954 VSS 0.012131f
C20503 VDD.n2955 VSS 0.012131f
C20504 VDD.n2956 VSS 0.012131f
C20505 VDD.n2957 VSS 0.012131f
C20506 VDD.n2958 VSS 0.012131f
C20507 VDD.n2959 VSS 0.012131f
C20508 VDD.n2960 VSS 0.012131f
C20509 VDD.n2961 VSS 0.012131f
C20510 VDD.n2962 VSS 0.012131f
C20511 VDD.n2963 VSS 0.012131f
C20512 VDD.n2964 VSS 0.012131f
C20513 VDD.n2965 VSS 0.012131f
C20514 VDD.n2966 VSS 0.269046f
C20515 VDD.n2967 VSS 0.012131f
C20516 VDD.n2968 VSS 0.012131f
C20517 VDD.n2969 VSS 0.206985f
C20518 VDD.n2970 VSS 0.011174f
C20519 VDD.n2971 VSS 0.012131f
C20520 VDD.n2972 VSS 0.012131f
C20521 VDD.n2973 VSS 0.012131f
C20522 VDD.n2974 VSS 0.012131f
C20523 VDD.n2975 VSS 0.012131f
C20524 VDD.n2976 VSS 0.012131f
C20525 VDD.n2977 VSS 0.012131f
C20526 VDD.n2978 VSS 0.012131f
C20527 VDD.n2979 VSS 0.012131f
C20528 VDD.n2980 VSS 0.012131f
C20529 VDD.n2981 VSS 0.012131f
C20530 VDD.n2982 VSS 0.012131f
C20531 VDD.n2983 VSS 0.012131f
C20532 VDD.n2984 VSS 0.012131f
C20533 VDD.n2985 VSS 0.012131f
C20534 VDD.n2986 VSS 0.012131f
C20535 VDD.n2987 VSS 0.012131f
C20536 VDD.n2988 VSS 0.012131f
C20537 VDD.n2989 VSS 0.012131f
C20538 VDD.n2990 VSS 0.012131f
C20539 VDD.n2991 VSS 0.012131f
C20540 VDD.n2992 VSS 0.012131f
C20541 VDD.n2993 VSS 0.012131f
C20542 VDD.n2994 VSS 0.012131f
C20543 VDD.n2995 VSS 0.012131f
C20544 VDD.n2996 VSS 0.012131f
C20545 VDD.n2997 VSS 0.012131f
C20546 VDD.n2998 VSS 0.012131f
C20547 VDD.n2999 VSS 0.012131f
C20548 VDD.n3000 VSS 0.012131f
C20549 VDD.n3001 VSS 0.012131f
C20550 VDD.n3002 VSS 0.012131f
C20551 VDD.n3003 VSS 0.012131f
C20552 VDD.n3004 VSS 0.012131f
C20553 VDD.n3005 VSS 0.012131f
C20554 VDD.n3006 VSS 0.012131f
C20555 VDD.n3007 VSS 0.012131f
C20556 VDD.n3008 VSS 0.012131f
C20557 VDD.n3009 VSS 0.012131f
C20558 VDD.n3010 VSS 0.012131f
C20559 VDD.n3011 VSS 0.012131f
C20560 VDD.n3012 VSS 0.012131f
C20561 VDD.n3013 VSS 0.012131f
C20562 VDD.n3014 VSS 0.012131f
C20563 VDD.n3015 VSS 0.012131f
C20564 VDD.n3016 VSS 0.012131f
C20565 VDD.n3017 VSS 0.012131f
C20566 VDD.n3018 VSS 0.012131f
C20567 VDD.n3019 VSS 0.012131f
C20568 VDD.n3020 VSS 0.012131f
C20569 VDD.n3021 VSS 0.012131f
C20570 VDD.n3022 VSS 0.012131f
C20571 VDD.n3023 VSS 0.012131f
C20572 VDD.n3024 VSS 0.012131f
C20573 VDD.n3025 VSS 0.012131f
C20574 VDD.n3026 VSS 0.012131f
C20575 VDD.n3027 VSS 0.012131f
C20576 VDD.n3028 VSS 0.012131f
C20577 VDD.n3029 VSS 0.012131f
C20578 VDD.n3030 VSS 0.012131f
C20579 VDD.n3031 VSS 0.012131f
C20580 VDD.n3032 VSS 0.012131f
C20581 VDD.n3033 VSS 0.012131f
C20582 VDD.n3034 VSS 0.012131f
C20583 VDD.n3035 VSS 0.012131f
C20584 VDD.n3036 VSS 0.012131f
C20585 VDD.n3037 VSS 0.012131f
C20586 VDD.n3038 VSS 0.012131f
C20587 VDD.n3039 VSS 0.012131f
C20588 VDD.n3040 VSS 0.012131f
C20589 VDD.n3041 VSS 0.012131f
C20590 VDD.n3042 VSS 0.012131f
C20591 VDD.n3043 VSS 0.012131f
C20592 VDD.n3044 VSS 0.012131f
C20593 VDD.n3045 VSS 0.012131f
C20594 VDD.n3046 VSS 0.012131f
C20595 VDD.n3047 VSS 0.012131f
C20596 VDD.n3048 VSS 0.012131f
C20597 VDD.n3049 VSS 0.012131f
C20598 VDD.n3050 VSS 0.012131f
C20599 VDD.n3051 VSS 0.012131f
C20600 VDD.n3052 VSS 0.012131f
C20601 VDD.n3053 VSS 0.012131f
C20602 VDD.n3054 VSS 0.012131f
C20603 VDD.n3055 VSS 0.012131f
C20604 VDD.n3056 VSS 0.012131f
C20605 VDD.n3057 VSS 0.012131f
C20606 VDD.n3058 VSS 0.012131f
C20607 VDD.n3059 VSS 0.012131f
C20608 VDD.n3060 VSS 0.012131f
C20609 VDD.n3061 VSS 0.012131f
C20610 VDD.n3062 VSS 0.012131f
C20611 VDD.n3063 VSS 0.012131f
C20612 VDD.n3064 VSS 0.012131f
C20613 VDD.n3065 VSS 0.012131f
C20614 VDD.n3066 VSS 0.012131f
C20615 VDD.n3067 VSS 0.012131f
C20616 VDD.n3068 VSS 0.012131f
C20617 VDD.n3069 VSS 0.012131f
C20618 VDD.n3070 VSS 0.012131f
C20619 VDD.n3071 VSS 0.012131f
C20620 VDD.n3072 VSS 0.012131f
C20621 VDD.n3073 VSS 0.012131f
C20622 VDD.n3074 VSS 0.012131f
C20623 VDD.n3075 VSS 0.012131f
C20624 VDD.n3076 VSS 0.012131f
C20625 VDD.n3077 VSS 0.012131f
C20626 VDD.n3078 VSS 0.012131f
C20627 VDD.n3079 VSS 0.012131f
C20628 VDD.n3080 VSS 0.012131f
C20629 VDD.n3081 VSS 0.012131f
C20630 VDD.n3082 VSS 0.012131f
C20631 VDD.n3083 VSS 0.012131f
C20632 VDD.n3084 VSS 0.012131f
C20633 VDD.n3085 VSS 0.012131f
C20634 VDD.n3086 VSS 0.012131f
C20635 VDD.n3087 VSS 0.012131f
C20636 VDD.n3088 VSS 0.012131f
C20637 VDD.n3089 VSS 0.012131f
C20638 VDD.n3090 VSS 0.012131f
C20639 VDD.n3091 VSS 0.012131f
C20640 VDD.n3092 VSS 0.012131f
C20641 VDD.n3093 VSS 0.012131f
C20642 VDD.n3094 VSS 0.012131f
C20643 VDD.n3095 VSS 0.012131f
C20644 VDD.n3096 VSS 0.012131f
C20645 VDD.n3097 VSS 0.012131f
C20646 VDD.n3098 VSS 0.012131f
C20647 VDD.n3099 VSS 0.012131f
C20648 VDD.n3100 VSS 0.012131f
C20649 VDD.n3101 VSS 0.012131f
C20650 VDD.n3102 VSS 0.012131f
C20651 VDD.n3103 VSS 0.012131f
C20652 VDD.n3104 VSS 0.012131f
C20653 VDD.n3105 VSS 0.012131f
C20654 VDD.n3106 VSS 0.012131f
C20655 VDD.n3107 VSS 0.012131f
C20656 VDD.n3108 VSS 0.012131f
C20657 VDD.n3109 VSS 0.012131f
C20658 VDD.n3110 VSS 0.012131f
C20659 VDD.n3111 VSS 0.012131f
C20660 VDD.n3112 VSS 0.012131f
C20661 VDD.n3113 VSS 0.012131f
C20662 VDD.n3114 VSS 0.012131f
C20663 VDD.n3115 VSS 0.012131f
C20664 VDD.n3116 VSS 0.012131f
C20665 VDD.n3117 VSS 0.012131f
C20666 VDD.n3118 VSS 0.012131f
C20667 VDD.n3119 VSS 0.012131f
C20668 VDD.n3120 VSS 0.012131f
C20669 VDD.n3121 VSS 0.012131f
C20670 VDD.n3122 VSS 0.012131f
C20671 VDD.n3123 VSS 0.012131f
C20672 VDD.n3124 VSS 0.012131f
C20673 VDD.n3125 VSS 0.012131f
C20674 VDD.n3126 VSS 0.012131f
C20675 VDD.n3127 VSS 0.012131f
C20676 VDD.n3128 VSS 0.012131f
C20677 VDD.n3129 VSS 0.012131f
C20678 VDD.n3130 VSS 0.012131f
C20679 VDD.n3131 VSS 0.012131f
C20680 VDD.n3132 VSS 0.012131f
C20681 VDD.n3133 VSS 0.012131f
C20682 VDD.n3134 VSS 0.012131f
C20683 VDD.n3135 VSS 0.012131f
C20684 VDD.n3136 VSS 0.012131f
C20685 VDD.n3137 VSS 0.012131f
C20686 VDD.n3138 VSS 0.012131f
C20687 VDD.n3139 VSS 0.012131f
C20688 VDD.n3140 VSS 0.012131f
C20689 VDD.n3141 VSS 0.012131f
C20690 VDD.n3142 VSS 0.012131f
C20691 VDD.n3143 VSS 0.012131f
C20692 VDD.n3144 VSS 0.012131f
C20693 VDD.n3145 VSS 0.012131f
C20694 VDD.n3146 VSS 0.012131f
C20695 VDD.n3147 VSS 0.012131f
C20696 VDD.n3148 VSS 0.012131f
C20697 VDD.n3149 VSS 0.012131f
C20698 VDD.n3150 VSS 0.012131f
C20699 VDD.n3151 VSS 0.012131f
C20700 VDD.n3152 VSS 0.012131f
C20701 VDD.n3153 VSS 0.012131f
C20702 VDD.n3154 VSS 0.012131f
C20703 VDD.n3155 VSS 0.012131f
C20704 VDD.n3156 VSS 0.012131f
C20705 VDD.n3157 VSS 0.012131f
C20706 VDD.n3158 VSS 0.012131f
C20707 VDD.n3159 VSS 0.012131f
C20708 VDD.n3160 VSS 0.012131f
C20709 VDD.n3161 VSS 0.012131f
C20710 VDD.n3162 VSS 0.012131f
C20711 VDD.n3163 VSS 0.012131f
C20712 VDD.n3164 VSS 0.012131f
C20713 VDD.n3165 VSS 0.012131f
C20714 VDD.n3166 VSS 0.012131f
C20715 VDD.n3167 VSS 0.012131f
C20716 VDD.n3168 VSS 0.012131f
C20717 VDD.n3169 VSS 0.012131f
C20718 VDD.n3170 VSS 0.012131f
C20719 VDD.n3171 VSS 0.012131f
C20720 VDD.n3172 VSS 0.012131f
C20721 VDD.n3173 VSS 0.012131f
C20722 VDD.n3174 VSS 0.012131f
C20723 VDD.n3175 VSS 0.012131f
C20724 VDD.n3176 VSS 0.012131f
C20725 VDD.n3177 VSS 0.012131f
C20726 VDD.n3178 VSS 0.012131f
C20727 VDD.n3179 VSS 0.012131f
C20728 VDD.n3180 VSS 0.012131f
C20729 VDD.n3181 VSS 0.012131f
C20730 VDD.n3182 VSS 0.012131f
C20731 VDD.n3183 VSS 0.012131f
C20732 VDD.n3184 VSS 0.012131f
C20733 VDD.n3185 VSS 0.012131f
C20734 VDD.n3186 VSS 0.012131f
C20735 VDD.n3187 VSS 0.012131f
C20736 VDD.n3188 VSS 0.012131f
C20737 VDD.n3189 VSS 0.012131f
C20738 VDD.n3190 VSS 0.012131f
C20739 VDD.n3191 VSS 0.012131f
C20740 VDD.n3192 VSS 0.012131f
C20741 VDD.n3193 VSS 0.012131f
C20742 VDD.n3194 VSS 0.012131f
C20743 VDD.n3195 VSS 0.012131f
C20744 VDD.n3196 VSS 0.012131f
C20745 VDD.n3197 VSS 0.012131f
C20746 VDD.n3198 VSS 0.012131f
C20747 VDD.n3199 VSS 0.012131f
C20748 VDD.n3200 VSS 0.012131f
C20749 VDD.n3201 VSS 0.012131f
C20750 VDD.n3202 VSS 0.012131f
C20751 VDD.n3203 VSS 0.012131f
C20752 VDD.n3204 VSS 0.012131f
C20753 VDD.n3205 VSS 0.012131f
C20754 VDD.n3206 VSS 0.012131f
C20755 VDD.n3207 VSS 0.012131f
C20756 VDD.n3208 VSS 0.012131f
C20757 VDD.n3209 VSS 0.012131f
C20758 VDD.n3210 VSS 0.012131f
C20759 VDD.n3211 VSS 0.012131f
C20760 VDD.n3212 VSS 0.012131f
C20761 VDD.n3213 VSS 0.012131f
C20762 VDD.n3214 VSS 0.012131f
C20763 VDD.n3215 VSS 0.012131f
C20764 VDD.n3216 VSS 0.012131f
C20765 VDD.n3217 VSS 0.012131f
C20766 VDD.n3218 VSS 0.012131f
C20767 VDD.n3219 VSS 0.012131f
C20768 VDD.n3220 VSS 0.012131f
C20769 VDD.n3221 VSS 0.012131f
C20770 VDD.n3222 VSS 0.012131f
C20771 VDD.n3223 VSS 0.012131f
C20772 VDD.n3224 VSS 0.012131f
C20773 VDD.n3225 VSS 0.012131f
C20774 VDD.n3226 VSS 0.012131f
C20775 VDD.n3227 VSS 0.012131f
C20776 VDD.n3228 VSS 0.012131f
C20777 VDD.n3229 VSS 0.012131f
C20778 VDD.n3230 VSS 0.012131f
C20779 VDD.n3231 VSS 0.012131f
C20780 VDD.n3232 VSS 0.012131f
C20781 VDD.n3233 VSS 0.012131f
C20782 VDD.n3234 VSS 0.012131f
C20783 VDD.n3235 VSS 0.012131f
C20784 VDD.n3236 VSS 0.012131f
C20785 VDD.n3237 VSS 0.012131f
C20786 VDD.n3238 VSS 0.012131f
C20787 VDD.n3239 VSS 0.012131f
C20788 VDD.n3240 VSS 0.012131f
C20789 VDD.n3241 VSS 0.012131f
C20790 VDD.n3242 VSS 0.012131f
C20791 VDD.n3243 VSS 0.012131f
C20792 VDD.n3244 VSS 0.012131f
C20793 VDD.n3245 VSS 0.012131f
C20794 VDD.n3246 VSS 0.012131f
C20795 VDD.n3247 VSS 0.012131f
C20796 VDD.n3248 VSS 0.012131f
C20797 VDD.n3249 VSS 0.012131f
C20798 VDD.n3250 VSS 0.012131f
C20799 VDD.n3251 VSS 0.012131f
C20800 VDD.n3252 VSS 0.012131f
C20801 VDD.n3253 VSS 0.012131f
C20802 VDD.n3254 VSS 0.012131f
C20803 VDD.n3255 VSS 0.012131f
C20804 VDD.n3256 VSS 0.012131f
C20805 VDD.n3257 VSS 0.012131f
C20806 VDD.n3258 VSS 0.012131f
C20807 VDD.n3259 VSS 0.012131f
C20808 VDD.n3260 VSS 0.012131f
C20809 VDD.n3261 VSS 0.012131f
C20810 VDD.n3262 VSS 0.012131f
C20811 VDD.n3263 VSS 0.012131f
C20812 VDD.n3264 VSS 0.012131f
C20813 VDD.n3265 VSS 0.012131f
C20814 VDD.n3266 VSS 0.012131f
C20815 VDD.n3267 VSS 0.012131f
C20816 VDD.n3268 VSS 0.012131f
C20817 VDD.n3269 VSS 0.012131f
C20818 VDD.n3270 VSS 0.012131f
C20819 VDD.n3271 VSS 0.012131f
C20820 VDD.n3272 VSS 0.012131f
C20821 VDD.n3273 VSS 0.012131f
C20822 VDD.n3274 VSS 0.012131f
C20823 VDD.n3275 VSS 0.012131f
C20824 VDD.n3276 VSS 0.012131f
C20825 VDD.n3277 VSS 0.012131f
C20826 VDD.n3278 VSS 0.012131f
C20827 VDD.n3279 VSS 0.012131f
C20828 VDD.n3280 VSS 0.012131f
C20829 VDD.n3281 VSS 0.012131f
C20830 VDD.n3282 VSS 0.012131f
C20831 VDD.n3283 VSS 0.012131f
C20832 VDD.n3284 VSS 0.012131f
C20833 VDD.n3285 VSS 0.012131f
C20834 VDD.n3286 VSS 0.012131f
C20835 VDD.n3287 VSS 0.012131f
C20836 VDD.n3288 VSS 0.012131f
C20837 VDD.n3289 VSS 0.012131f
C20838 VDD.n3290 VSS 0.012131f
C20839 VDD.n3291 VSS 0.012131f
C20840 VDD.n3292 VSS 0.012131f
C20841 VDD.n3293 VSS 0.012131f
C20842 VDD.n3294 VSS 0.012131f
C20843 VDD.n3295 VSS 0.012131f
C20844 VDD.n3296 VSS 0.012131f
C20845 VDD.n3297 VSS 0.012131f
C20846 VDD.n3298 VSS 0.012131f
C20847 VDD.n3299 VSS 0.012131f
C20848 VDD.n3300 VSS 0.012131f
C20849 VDD.n3301 VSS 0.012131f
C20850 VDD.n3302 VSS 0.012131f
C20851 VDD.n3303 VSS 0.012131f
C20852 VDD.n3304 VSS 0.012131f
C20853 VDD.n3305 VSS 0.012131f
C20854 VDD.n3306 VSS 0.012131f
C20855 VDD.n3307 VSS 0.012131f
C20856 VDD.n3308 VSS 0.012131f
C20857 VDD.n3309 VSS 0.012131f
C20858 VDD.n3310 VSS 0.012131f
C20859 VDD.n3311 VSS 0.012131f
C20860 VDD.n3312 VSS 0.012131f
C20861 VDD.n3313 VSS 0.012131f
C20862 VDD.n3314 VSS 0.012131f
C20863 VDD.n3315 VSS 0.012131f
C20864 VDD.n3316 VSS 0.012131f
C20865 VDD.n3317 VSS 0.012131f
C20866 VDD.n3318 VSS 0.012131f
C20867 VDD.n3319 VSS 0.012131f
C20868 VDD.n3320 VSS 0.012131f
C20869 VDD.n3321 VSS 0.012131f
C20870 VDD.n3322 VSS 0.012131f
C20871 VDD.n3323 VSS 0.012131f
C20872 VDD.n3324 VSS 0.012131f
C20873 VDD.n3325 VSS 0.012131f
C20874 VDD.n3326 VSS 0.012131f
C20875 VDD.n3327 VSS 0.012131f
C20876 VDD.n3328 VSS 0.012131f
C20877 VDD.n3329 VSS 0.012131f
C20878 VDD.n3330 VSS 0.012131f
C20879 VDD.n3331 VSS 0.012131f
C20880 VDD.n3332 VSS 0.012131f
C20881 VDD.n3333 VSS 0.012131f
C20882 VDD.n3334 VSS 0.012131f
C20883 VDD.n3335 VSS 0.012131f
C20884 VDD.n3336 VSS 0.012131f
C20885 VDD.n3337 VSS 0.012131f
C20886 VDD.n3338 VSS 0.012131f
C20887 VDD.n3339 VSS 0.012131f
C20888 VDD.n3340 VSS 0.012131f
C20889 VDD.n3341 VSS 0.012131f
C20890 VDD.n3342 VSS 0.012131f
C20891 VDD.n3343 VSS 0.012131f
C20892 VDD.n3344 VSS 0.012131f
C20893 VDD.n3345 VSS 0.012131f
C20894 VDD.n3346 VSS 0.012131f
C20895 VDD.n3347 VSS 0.012131f
C20896 VDD.n3348 VSS 0.012131f
C20897 VDD.n3349 VSS 0.012131f
C20898 VDD.n3350 VSS 0.012131f
C20899 VDD.n3351 VSS 0.012131f
C20900 VDD.n3352 VSS 0.012131f
C20901 VDD.n3353 VSS 0.012131f
C20902 VDD.n3354 VSS 0.012131f
C20903 VDD.n3355 VSS 0.012131f
C20904 VDD.n3356 VSS 0.012131f
C20905 VDD.n3357 VSS 0.012131f
C20906 VDD.n3358 VSS 0.012131f
C20907 VDD.n3359 VSS 0.012131f
C20908 VDD.n3360 VSS 0.012131f
C20909 VDD.n3361 VSS 0.012131f
C20910 VDD.n3362 VSS 0.012131f
C20911 VDD.n3363 VSS 0.012131f
C20912 VDD.n3364 VSS 0.012131f
C20913 VDD.n3365 VSS 0.012131f
C20914 VDD.n3366 VSS 0.012131f
C20915 VDD.n3367 VSS 0.012131f
C20916 VDD.n3368 VSS 0.012131f
C20917 VDD.n3369 VSS 0.012131f
C20918 VDD.n3370 VSS 0.012131f
C20919 VDD.n3371 VSS 0.012131f
C20920 VDD.n3372 VSS 0.012131f
C20921 VDD.n3373 VSS 0.012131f
C20922 VDD.n3374 VSS 0.012131f
C20923 VDD.n3375 VSS 0.012131f
C20924 VDD.n3376 VSS 0.012131f
C20925 VDD.n3377 VSS 0.012131f
C20926 VDD.n3378 VSS 0.012131f
C20927 VDD.n3379 VSS 0.012131f
C20928 VDD.n3380 VSS 0.012131f
C20929 VDD.n3381 VSS 0.012131f
C20930 VDD.n3382 VSS 0.012131f
C20931 VDD.n3383 VSS 0.012131f
C20932 VDD.n3384 VSS 0.012131f
C20933 VDD.n3385 VSS 0.012131f
C20934 VDD.n3386 VSS 0.012131f
C20935 VDD.n3387 VSS 0.012131f
C20936 VDD.n3388 VSS 0.012131f
C20937 VDD.n3389 VSS 0.012131f
C20938 VDD.n3390 VSS 0.012131f
C20939 VDD.n3391 VSS 0.012131f
C20940 VDD.n3392 VSS 0.012131f
C20941 VDD.n3393 VSS 0.012131f
C20942 VDD.n3394 VSS 0.012131f
C20943 VDD.n3395 VSS 0.012131f
C20944 VDD.n3396 VSS 0.012131f
C20945 VDD.n3397 VSS 0.012131f
C20946 VDD.n3398 VSS 0.012131f
C20947 VDD.n3399 VSS 0.012131f
C20948 VDD.n3400 VSS 0.012131f
C20949 VDD.n3401 VSS 0.012131f
C20950 VDD.n3402 VSS 0.012131f
C20951 VDD.n3403 VSS 0.012131f
C20952 VDD.n3404 VSS 0.012131f
C20953 VDD.n3405 VSS 0.012131f
C20954 VDD.n3406 VSS 0.012131f
C20955 VDD.n3407 VSS 0.012131f
C20956 VDD.n3408 VSS 0.012131f
C20957 VDD.n3409 VSS 0.012131f
C20958 VDD.n3410 VSS 0.012131f
C20959 VDD.n3411 VSS 0.012131f
C20960 VDD.n3412 VSS 0.012131f
C20961 VDD.n3413 VSS 0.012131f
C20962 VDD.n3414 VSS 0.012131f
C20963 VDD.n3415 VSS 0.012131f
C20964 VDD.n3416 VSS 0.012131f
C20965 VDD.n3417 VSS 0.012131f
C20966 VDD.n3418 VSS 0.012131f
C20967 VDD.n3419 VSS 0.012131f
C20968 VDD.n3420 VSS 0.012131f
C20969 VDD.n3421 VSS 0.012131f
C20970 VDD.n3422 VSS 0.012131f
C20971 VDD.n3423 VSS 0.012131f
C20972 VDD.n3424 VSS 0.012131f
C20973 VDD.n3425 VSS 0.012131f
C20974 VDD.n3426 VSS 0.012131f
C20975 VDD.n3427 VSS 0.012131f
C20976 VDD.n3428 VSS 0.012131f
C20977 VDD.n3429 VSS 0.012131f
C20978 VDD.n3430 VSS 0.012131f
C20979 VDD.n3431 VSS 0.012131f
C20980 VDD.n3432 VSS 0.012131f
C20981 VDD.n3433 VSS 0.012131f
C20982 VDD.n3434 VSS 0.012131f
C20983 VDD.n3435 VSS 0.012131f
C20984 VDD.n3436 VSS 0.012131f
C20985 VDD.n3437 VSS 0.012131f
C20986 VDD.n3438 VSS 0.012131f
C20987 VDD.n3439 VSS 0.012131f
C20988 VDD.n3440 VSS 0.012131f
C20989 VDD.n3441 VSS 0.012131f
C20990 VDD.n3442 VSS 0.012131f
C20991 VDD.n3443 VSS 0.012131f
C20992 VDD.n3444 VSS 0.012131f
C20993 VDD.n3445 VSS 0.012131f
C20994 VDD.n3446 VSS 0.012131f
C20995 VDD.n3447 VSS 0.012131f
C20996 VDD.n3448 VSS 0.012131f
C20997 VDD.n3449 VSS 0.012131f
C20998 VDD.n3450 VSS 0.012131f
C20999 VDD.n3451 VSS 0.012131f
C21000 VDD.n3452 VSS 0.012131f
C21001 VDD.n3453 VSS 0.012131f
C21002 VDD.n3454 VSS 0.012131f
C21003 VDD.n3455 VSS 0.012131f
C21004 VDD.n3456 VSS 0.012131f
C21005 VDD.n3457 VSS 0.012131f
C21006 VDD.n3458 VSS 0.012131f
C21007 VDD.n3459 VSS 0.012131f
C21008 VDD.n3460 VSS 0.012131f
C21009 VDD.n3461 VSS 0.012131f
C21010 VDD.n3462 VSS 0.012131f
C21011 VDD.n3463 VSS 0.012131f
C21012 VDD.n3464 VSS 0.012131f
C21013 VDD.n3465 VSS 0.012131f
C21014 VDD.n3466 VSS 0.012131f
C21015 VDD.n3467 VSS 0.012131f
C21016 VDD.n3468 VSS 0.012131f
C21017 VDD.n3469 VSS 0.012131f
C21018 VDD.n3470 VSS 0.012131f
C21019 VDD.n3471 VSS 0.012131f
C21020 VDD.n3472 VSS 0.012131f
C21021 VDD.n3473 VSS 0.012131f
C21022 VDD.n3474 VSS 0.012131f
C21023 VDD.n3475 VSS 0.012131f
C21024 VDD.n3476 VSS 0.012131f
C21025 VDD.n3477 VSS 0.012131f
C21026 VDD.n3478 VSS 0.012131f
C21027 VDD.n3479 VSS 0.012131f
C21028 VDD.n3480 VSS 0.012131f
C21029 VDD.n3481 VSS 0.012131f
C21030 VDD.n3482 VSS 0.012131f
C21031 VDD.n3483 VSS 0.012131f
C21032 VDD.n3484 VSS 0.012131f
C21033 VDD.n3485 VSS 0.012131f
C21034 VDD.n3486 VSS 0.012131f
C21035 VDD.n3487 VSS 0.012131f
C21036 VDD.n3488 VSS 0.012131f
C21037 VDD.n3489 VSS 0.012131f
C21038 VDD.n3490 VSS 0.012131f
C21039 VDD.n3491 VSS 0.012131f
C21040 VDD.n3492 VSS 0.012131f
C21041 VDD.n3493 VSS 0.012131f
C21042 VDD.n3494 VSS 0.012131f
C21043 VDD.n3495 VSS 0.012131f
C21044 VDD.n3496 VSS 0.012131f
C21045 VDD.n3497 VSS 0.012131f
C21046 VDD.n3498 VSS 0.012131f
C21047 VDD.n3499 VSS 0.012131f
C21048 VDD.n3500 VSS 0.012131f
C21049 VDD.n3501 VSS 0.012131f
C21050 VDD.n3502 VSS 0.012131f
C21051 VDD.n3503 VSS 0.012131f
C21052 VDD.n3504 VSS 0.012131f
C21053 VDD.n3505 VSS 0.012131f
C21054 VDD.n3506 VSS 0.012131f
C21055 VDD.n3507 VSS 0.012131f
C21056 VDD.n3508 VSS 0.012131f
C21057 VDD.n3509 VSS 0.012131f
C21058 VDD.n3510 VSS 0.012131f
C21059 VDD.n3511 VSS 0.012131f
C21060 VDD.n3512 VSS 0.012131f
C21061 VDD.n3513 VSS 0.012131f
C21062 VDD.n3514 VSS 0.012131f
C21063 VDD.n3515 VSS 0.012131f
C21064 VDD.n3516 VSS 0.012131f
C21065 VDD.n3517 VSS 0.012131f
C21066 VDD.n3518 VSS 0.012131f
C21067 VDD.n3519 VSS 0.012131f
C21068 VDD.n3520 VSS 0.012131f
C21069 VDD.n3521 VSS 0.012131f
C21070 VDD.n3522 VSS 0.012131f
C21071 VDD.n3523 VSS 0.012131f
C21072 VDD.n3524 VSS 0.012131f
C21073 VDD.n3525 VSS 0.012131f
C21074 VDD.n3526 VSS 0.012131f
C21075 VDD.n3527 VSS 0.012131f
C21076 VDD.n3528 VSS 0.012131f
C21077 VDD.n3529 VSS 0.012131f
C21078 VDD.n3530 VSS 0.012131f
C21079 VDD.n3531 VSS 0.012131f
C21080 VDD.n3532 VSS 0.012131f
C21081 VDD.n3533 VSS 0.012131f
C21082 VDD.n3534 VSS 0.012131f
C21083 VDD.n3535 VSS 0.012131f
C21084 VDD.n3536 VSS 0.012131f
C21085 VDD.n3537 VSS 0.012131f
C21086 VDD.n3538 VSS 0.012131f
C21087 VDD.n3539 VSS 0.012131f
C21088 VDD.n3540 VSS 0.012131f
C21089 VDD.n3541 VSS 0.012131f
C21090 VDD.n3542 VSS 0.012131f
C21091 VDD.n3543 VSS 0.012131f
C21092 VDD.n3544 VSS 0.012131f
C21093 VDD.n3545 VSS 0.012131f
C21094 VDD.n3546 VSS 0.012131f
C21095 VDD.n3547 VSS 0.012131f
C21096 VDD.n3548 VSS 0.012131f
C21097 VDD.n3549 VSS 0.012131f
C21098 VDD.n3550 VSS 0.012131f
C21099 VDD.n3551 VSS 0.012131f
C21100 VDD.n3552 VSS 0.012131f
C21101 VDD.n3553 VSS 0.012131f
C21102 VDD.n3554 VSS 0.012131f
C21103 VDD.n3555 VSS 0.012131f
C21104 VDD.n3556 VSS 0.012131f
C21105 VDD.n3557 VSS 0.012131f
C21106 VDD.n3558 VSS 0.012131f
C21107 VDD.n3559 VSS 0.012131f
C21108 VDD.n3560 VSS 0.012131f
C21109 VDD.n3561 VSS 0.012131f
C21110 VDD.n3562 VSS 0.012131f
C21111 VDD.n3563 VSS 0.012131f
C21112 VDD.n3564 VSS 0.012131f
C21113 VDD.n3565 VSS 0.012131f
C21114 VDD.n3566 VSS 0.012131f
C21115 VDD.n3567 VSS 0.012131f
C21116 VDD.n3568 VSS 0.012131f
C21117 VDD.n3569 VSS 0.012131f
C21118 VDD.n3570 VSS 0.012131f
C21119 VDD.n3571 VSS 0.012131f
C21120 VDD.n3572 VSS 0.012131f
C21121 VDD.n3573 VSS 0.012131f
C21122 VDD.n3574 VSS 0.012131f
C21123 VDD.n3575 VSS 0.012131f
C21124 VDD.n3576 VSS 0.012131f
C21125 VDD.n3577 VSS 0.012131f
C21126 VDD.n3578 VSS 0.012131f
C21127 VDD.n3579 VSS 0.012131f
C21128 VDD.n3580 VSS 0.012131f
C21129 VDD.n3581 VSS 0.012131f
C21130 VDD.n3582 VSS 0.012131f
C21131 VDD.n3583 VSS 0.012131f
C21132 VDD.n3584 VSS 0.012131f
C21133 VDD.n3585 VSS 0.012131f
C21134 VDD.n3586 VSS 0.012131f
C21135 VDD.n3587 VSS 0.012131f
C21136 VDD.n3588 VSS 0.012131f
C21137 VDD.n3589 VSS 0.012131f
C21138 VDD.n3590 VSS 0.012131f
C21139 VDD.n3591 VSS 0.012131f
C21140 VDD.n3592 VSS 0.012131f
C21141 VDD.n3593 VSS 0.012131f
C21142 VDD.n3594 VSS 0.012131f
C21143 VDD.n3595 VSS 0.012131f
C21144 VDD.n3596 VSS 0.012131f
C21145 VDD.n3597 VSS 0.012131f
C21146 VDD.n3598 VSS 0.012131f
C21147 VDD.n3599 VSS 0.012131f
C21148 VDD.n3600 VSS 0.012131f
C21149 VDD.n3601 VSS 0.012131f
C21150 VDD.n3602 VSS 0.012131f
C21151 VDD.n3603 VSS 0.012131f
C21152 VDD.n3604 VSS 0.012131f
C21153 VDD.n3605 VSS 0.012131f
C21154 VDD.n3606 VSS 0.012131f
C21155 VDD.n3607 VSS 0.012131f
C21156 VDD.n3608 VSS 0.012131f
C21157 VDD.n3609 VSS 0.012131f
C21158 VDD.n3610 VSS 0.012131f
C21159 VDD.n3611 VSS 0.012131f
C21160 VDD.n3612 VSS 0.012131f
C21161 VDD.n3613 VSS 0.012131f
C21162 VDD.n3614 VSS 0.012131f
C21163 VDD.n3615 VSS 0.012131f
C21164 VDD.n3616 VSS 0.012131f
C21165 VDD.n3617 VSS 0.012131f
C21166 VDD.n3618 VSS 0.012131f
C21167 VDD.n3619 VSS 0.012131f
C21168 VDD.n3620 VSS 0.012131f
C21169 VDD.n3621 VSS 0.012131f
C21170 VDD.n3622 VSS 0.012131f
C21171 VDD.n3623 VSS 0.012131f
C21172 VDD.n3624 VSS 0.012131f
C21173 VDD.n3625 VSS 0.012131f
C21174 VDD.n3626 VSS 0.012131f
C21175 VDD.n3627 VSS 0.012131f
C21176 VDD.n3628 VSS 0.032462f
C21177 VDD.n3629 VSS 0.032462f
C21178 VDD.n3630 VSS 0.026818f
C21179 VDD.n3631 VSS 0.012131f
C21180 VDD.n3632 VSS 0.012131f
C21181 VDD.n3633 VSS 0.012131f
C21182 VDD.n3634 VSS 0.012131f
C21183 VDD.n3635 VSS 0.012131f
C21184 VDD.n3636 VSS 0.012131f
C21185 VDD.n3637 VSS 0.012131f
C21186 VDD.n3638 VSS 0.012131f
C21187 VDD.n3639 VSS 0.012131f
C21188 VDD.n3640 VSS 0.012131f
C21189 VDD.n3641 VSS 0.012131f
C21190 VDD.n3642 VSS 0.012131f
C21191 VDD.n3643 VSS 0.012131f
C21192 VDD.n3644 VSS 0.012131f
C21193 VDD.n3645 VSS 0.012131f
C21194 VDD.n3646 VSS 0.012131f
C21195 VDD.n3647 VSS 0.012131f
C21196 VDD.n3648 VSS 0.012131f
C21197 VDD.n3649 VSS 0.012131f
C21198 VDD.n3650 VSS 0.012131f
C21199 VDD.n3651 VSS 0.012131f
C21200 VDD.n3652 VSS 0.012131f
C21201 VDD.n3653 VSS 0.012131f
C21202 VDD.n3654 VSS 0.012131f
C21203 VDD.n3655 VSS 0.012131f
C21204 VDD.n3656 VSS 0.012131f
C21205 VDD.n3657 VSS 0.012131f
C21206 VDD.n3658 VSS 0.012131f
C21207 VDD.n3659 VSS 0.012131f
C21208 VDD.n3660 VSS 0.012131f
C21209 VDD.n3661 VSS 0.012131f
C21210 VDD.n3662 VSS 0.012131f
C21211 VDD.n3663 VSS 0.012131f
C21212 VDD.n3664 VSS 0.012131f
C21213 VDD.n3665 VSS 0.012131f
C21214 VDD.n3666 VSS 0.012131f
C21215 VDD.n3667 VSS 0.012131f
C21216 VDD.n3668 VSS 0.012131f
C21217 VDD.n3669 VSS 0.012131f
C21218 VDD.n3670 VSS 0.012131f
C21219 VDD.n3671 VSS 0.012131f
C21220 VDD.n3672 VSS 0.012131f
C21221 VDD.n3673 VSS 0.012131f
C21222 VDD.n3674 VSS 0.012131f
C21223 VDD.n3675 VSS 0.012131f
C21224 VDD.n3676 VSS 0.012131f
C21225 VDD.n3677 VSS 0.012131f
C21226 VDD.n3678 VSS 0.012131f
C21227 VDD.n3679 VSS 0.012131f
C21228 VDD.n3680 VSS 0.012131f
C21229 VDD.n3681 VSS 0.012131f
C21230 VDD.n3682 VSS 0.012131f
C21231 VDD.n3683 VSS 0.012131f
C21232 VDD.n3684 VSS 0.012131f
C21233 VDD.n3685 VSS 0.012131f
C21234 VDD.n3686 VSS 0.012131f
C21235 VDD.n3687 VSS 0.012131f
C21236 VDD.n3688 VSS 0.012131f
C21237 VDD.n3689 VSS 0.012131f
C21238 VDD.n3690 VSS 0.012131f
C21239 VDD.n3691 VSS 0.012131f
C21240 VDD.n3692 VSS 0.012131f
C21241 VDD.n3693 VSS 0.012131f
C21242 VDD.n3694 VSS 0.012131f
C21243 VDD.n3695 VSS 0.012131f
C21244 VDD.n3696 VSS 0.012131f
C21245 VDD.n3697 VSS 0.012131f
C21246 VDD.n3698 VSS 0.012131f
C21247 VDD.n3699 VSS 0.012131f
C21248 VDD.n3700 VSS 0.012131f
C21249 VDD.n3701 VSS 0.012131f
C21250 VDD.n3702 VSS 0.012131f
C21251 VDD.n3703 VSS 0.012131f
C21252 VDD.n3704 VSS 0.012131f
C21253 VDD.n3705 VSS 0.012131f
C21254 VDD.n3706 VSS 0.012131f
C21255 VDD.n3707 VSS 0.012131f
C21256 VDD.n3708 VSS 0.012131f
C21257 VDD.n3709 VSS 0.012131f
C21258 VDD.n3710 VSS 0.012131f
C21259 VDD.n3711 VSS 0.012131f
C21260 VDD.n3712 VSS 0.012131f
C21261 VDD.n3713 VSS 0.012131f
C21262 VDD.n3714 VSS 0.012131f
C21263 VDD.n3715 VSS 0.012131f
C21264 VDD.n3716 VSS 0.012131f
C21265 VDD.n3717 VSS 0.012131f
C21266 VDD.n3718 VSS 0.012131f
C21267 VDD.n3719 VSS 0.012131f
C21268 VDD.n3720 VSS 0.012131f
C21269 VDD.n3721 VSS 0.012131f
C21270 VDD.n3722 VSS 0.012131f
C21271 VDD.n3723 VSS 0.012131f
C21272 VDD.n3724 VSS 0.012131f
C21273 VDD.n3725 VSS 0.012131f
C21274 VDD.n3726 VSS 0.012131f
C21275 VDD.n3727 VSS 0.012131f
C21276 VDD.n3728 VSS 0.012131f
C21277 VDD.n3729 VSS 0.012131f
C21278 VDD.n3730 VSS 0.012131f
C21279 VDD.n3731 VSS 0.012131f
C21280 VDD.n3732 VSS 0.012131f
C21281 VDD.n3733 VSS 0.012131f
C21282 VDD.n3734 VSS 0.012131f
C21283 VDD.n3735 VSS 0.012131f
C21284 VDD.n3736 VSS 0.012131f
C21285 VDD.n3737 VSS 0.012131f
C21286 VDD.n3738 VSS 0.012131f
C21287 VDD.n3739 VSS 0.012131f
C21288 VDD.n3740 VSS 0.012131f
C21289 VDD.n3741 VSS 0.012131f
C21290 VDD.n3742 VSS 0.012131f
C21291 VDD.n3743 VSS 0.012131f
C21292 VDD.n3744 VSS 0.012131f
C21293 VDD.n3745 VSS 0.012131f
C21294 VDD.n3746 VSS 0.012131f
C21295 VDD.n3747 VSS 0.012131f
C21296 VDD.n3748 VSS 0.012131f
C21297 VDD.n3749 VSS 0.012131f
C21298 VDD.n3750 VSS 0.012131f
C21299 VDD.n3751 VSS 0.012131f
C21300 VDD.n3752 VSS 0.012131f
C21301 VDD.n3753 VSS 0.012131f
C21302 VDD.n3754 VSS 0.012131f
C21303 VDD.n3755 VSS 0.012131f
C21304 VDD.n3756 VSS 0.012131f
C21305 VDD.n3757 VSS 0.012131f
C21306 VDD.n3758 VSS 0.012131f
C21307 VDD.n3759 VSS 0.012131f
C21308 VDD.n3760 VSS 0.012131f
C21309 VDD.n3761 VSS 0.012131f
C21310 VDD.n3762 VSS 0.012131f
C21311 VDD.n3763 VSS 0.012131f
C21312 VDD.n3764 VSS 0.012131f
C21313 VDD.n3765 VSS 0.012131f
C21314 VDD.n3766 VSS 0.012131f
C21315 VDD.n3767 VSS 0.012131f
C21316 VDD.n3768 VSS 0.012131f
C21317 VDD.n3769 VSS 0.012131f
C21318 VDD.n3770 VSS 0.012131f
C21319 VDD.n3771 VSS 0.012131f
C21320 VDD.n3772 VSS 0.012131f
C21321 VDD.n3773 VSS 0.012131f
C21322 VDD.n3774 VSS 0.012131f
C21323 VDD.n3775 VSS 0.012131f
C21324 VDD.n3776 VSS 0.012131f
C21325 VDD.n3777 VSS 0.012131f
C21326 VDD.n3778 VSS 0.012131f
C21327 VDD.n3779 VSS 0.012131f
C21328 VDD.n3780 VSS 0.012131f
C21329 VDD.n3781 VSS 0.012131f
C21330 VDD.n3782 VSS 0.012131f
C21331 VDD.n3783 VSS 0.012131f
C21332 VDD.n3784 VSS 0.012131f
C21333 VDD.n3785 VSS 0.012131f
C21334 VDD.n3786 VSS 0.012131f
C21335 VDD.n3787 VSS 0.012131f
C21336 VDD.n3788 VSS 0.012131f
C21337 VDD.n3789 VSS 0.012131f
C21338 VDD.n3790 VSS 0.012131f
C21339 VDD.n3791 VSS 0.012131f
C21340 VDD.n3792 VSS 0.012131f
C21341 VDD.n3793 VSS 0.012131f
C21342 VDD.n3794 VSS 0.012131f
C21343 VDD.n3795 VSS 0.012131f
C21344 VDD.n3796 VSS 0.012131f
C21345 VDD.n3797 VSS 0.012131f
C21346 VDD.n3798 VSS 0.012131f
C21347 VDD.n3799 VSS 0.012131f
C21348 VDD.n3800 VSS 0.012131f
C21349 VDD.n3801 VSS 0.012131f
C21350 VDD.n3802 VSS 0.012131f
C21351 VDD.n3803 VSS 0.012131f
C21352 VDD.n3804 VSS 0.012131f
C21353 VDD.n3805 VSS 0.012131f
C21354 VDD.n3806 VSS 0.012131f
C21355 VDD.n3807 VSS 0.012131f
C21356 VDD.n3808 VSS 0.012131f
C21357 VDD.n3809 VSS 0.012131f
C21358 VDD.n3810 VSS 0.012131f
C21359 VDD.n3811 VSS 0.012131f
C21360 VDD.n3812 VSS 0.012131f
C21361 VDD.n3813 VSS 0.012131f
C21362 VDD.n3814 VSS 0.012131f
C21363 VDD.n3815 VSS 0.012131f
C21364 VDD.n3816 VSS 0.012131f
C21365 VDD.n3817 VSS 0.012131f
C21366 VDD.n3818 VSS 0.012131f
C21367 VDD.n3819 VSS 0.012131f
C21368 VDD.n3820 VSS 0.012131f
C21369 VDD.n3821 VSS 0.012131f
C21370 VDD.n3822 VSS 0.012131f
C21371 VDD.n3823 VSS 0.012131f
C21372 VDD.n3824 VSS 0.012131f
C21373 VDD.n3825 VSS 0.012131f
C21374 VDD.n3826 VSS 0.012131f
C21375 VDD.n3827 VSS 0.012131f
C21376 VDD.n3828 VSS 0.012131f
C21377 VDD.n3829 VSS 0.012131f
C21378 VDD.n3830 VSS 0.012131f
C21379 VDD.n3831 VSS 0.012131f
C21380 VDD.n3832 VSS 0.012131f
C21381 VDD.n3833 VSS 0.012131f
C21382 VDD.n3834 VSS 0.012131f
C21383 VDD.n3835 VSS 0.012131f
C21384 VDD.n3836 VSS 0.012131f
C21385 VDD.n3837 VSS 0.012131f
C21386 VDD.n3838 VSS 0.012131f
C21387 VDD.n3839 VSS 0.012131f
C21388 VDD.n3840 VSS 0.012131f
C21389 VDD.n3841 VSS 0.012131f
C21390 VDD.n3842 VSS 0.012131f
C21391 VDD.n3843 VSS 0.012131f
C21392 VDD.n3844 VSS 0.012131f
C21393 VDD.n3845 VSS 0.012131f
C21394 VDD.n3846 VSS 0.012131f
C21395 VDD.n3847 VSS 0.012131f
C21396 VDD.n3848 VSS 0.012131f
C21397 VDD.n3849 VSS 0.012131f
C21398 VDD.n3850 VSS 0.012131f
C21399 VDD.n3851 VSS 0.012131f
C21400 VDD.n3852 VSS 0.012131f
C21401 VDD.n3853 VSS 0.012131f
C21402 VDD.n3854 VSS 0.012131f
C21403 VDD.n3855 VSS 0.012131f
C21404 VDD.n3856 VSS 0.012131f
C21405 VDD.n3857 VSS 0.012131f
C21406 VDD.n3858 VSS 0.012131f
C21407 VDD.n3859 VSS 0.012131f
C21408 VDD.n3860 VSS 0.012131f
C21409 VDD.n3861 VSS 0.012131f
C21410 VDD.n3862 VSS 0.012131f
C21411 VDD.n3863 VSS 0.012131f
C21412 VDD.n3864 VSS 0.012131f
C21413 VDD.n3865 VSS 0.012131f
C21414 VDD.n3866 VSS 0.012131f
C21415 VDD.n3867 VSS 0.012131f
C21416 VDD.n3868 VSS 0.012131f
C21417 VDD.n3869 VSS 0.012131f
C21418 VDD.n3870 VSS 0.012131f
C21419 VDD.n3871 VSS 0.012131f
C21420 VDD.n3872 VSS 0.012131f
C21421 VDD.n3873 VSS 0.012131f
C21422 VDD.n3874 VSS 0.012131f
C21423 VDD.n3875 VSS 0.012131f
C21424 VDD.n3876 VSS 0.012131f
C21425 VDD.n3877 VSS 0.012131f
C21426 VDD.n3878 VSS 0.012131f
C21427 VDD.n3879 VSS 0.012131f
C21428 VDD.n3880 VSS 0.012131f
C21429 VDD.n3881 VSS 0.012131f
C21430 VDD.n3882 VSS 0.012131f
C21431 VDD.n3883 VSS 0.012131f
C21432 VDD.n3884 VSS 0.012131f
C21433 VDD.n3885 VSS 0.012131f
C21434 VDD.n3886 VSS 0.012131f
C21435 VDD.n3887 VSS 0.012131f
C21436 VDD.n3888 VSS 0.012131f
C21437 VDD.n3889 VSS 0.012131f
C21438 VDD.n3890 VSS 0.012131f
C21439 VDD.n3891 VSS 0.012131f
C21440 VDD.n3892 VSS 0.012131f
C21441 VDD.n3893 VSS 0.012131f
C21442 VDD.n3894 VSS 0.012131f
C21443 VDD.n3895 VSS 0.012131f
C21444 VDD.n3896 VSS 0.012131f
C21445 VDD.n3897 VSS 0.012131f
C21446 VDD.n3898 VSS 0.012131f
C21447 VDD.n3899 VSS 0.012131f
C21448 VDD.n3900 VSS 0.012131f
C21449 VDD.n3901 VSS 0.012131f
C21450 VDD.n3902 VSS 0.012131f
C21451 VDD.n3903 VSS 0.012131f
C21452 VDD.n3904 VSS 0.012131f
C21453 VDD.n3905 VSS 0.012131f
C21454 VDD.n3906 VSS 0.012131f
C21455 VDD.n3907 VSS 0.012131f
C21456 VDD.n3908 VSS 0.012131f
C21457 VDD.n3909 VSS 0.012131f
C21458 VDD.n3910 VSS 0.012131f
C21459 VDD.n3911 VSS 0.012131f
C21460 VDD.n3912 VSS 0.012131f
C21461 VDD.n3913 VSS 0.012131f
C21462 VDD.n3914 VSS 0.012131f
C21463 VDD.n3915 VSS 0.012131f
C21464 VDD.n3916 VSS 0.012131f
C21465 VDD.n3917 VSS 0.012131f
C21466 VDD.n3918 VSS 0.012131f
C21467 VDD.n3919 VSS 0.012131f
C21468 VDD.n3920 VSS 0.012131f
C21469 VDD.n3921 VSS 0.012131f
C21470 VDD.n3922 VSS 0.012131f
C21471 VDD.n3923 VSS 0.012131f
C21472 VDD.n3924 VSS 0.012131f
C21473 VDD.n3925 VSS 0.012131f
C21474 VDD.n3926 VSS 0.012131f
C21475 VDD.n3927 VSS 0.012131f
C21476 VDD.n3928 VSS 0.012131f
C21477 VDD.n3929 VSS 0.012131f
C21478 VDD.n3930 VSS 0.012131f
C21479 VDD.n3931 VSS 0.012131f
C21480 VDD.n3932 VSS 0.012131f
C21481 VDD.n3933 VSS 0.012131f
C21482 VDD.n3934 VSS 0.012131f
C21483 VDD.n3935 VSS 0.012131f
C21484 VDD.n3936 VSS 0.012131f
C21485 VDD.n3937 VSS 0.012131f
C21486 VDD.n3938 VSS 0.012131f
C21487 VDD.n3939 VSS 0.012131f
C21488 VDD.n3940 VSS 0.012131f
C21489 VDD.n3941 VSS 0.012131f
C21490 VDD.n3942 VSS 0.012131f
C21491 VDD.n3943 VSS 0.012131f
C21492 VDD.n3944 VSS 0.012131f
C21493 VDD.n3945 VSS 0.012131f
C21494 VDD.n3946 VSS 0.012131f
C21495 VDD.n3947 VSS 0.012131f
C21496 VDD.n3948 VSS 0.012131f
C21497 VDD.n3949 VSS 0.012131f
C21498 VDD.n3950 VSS 0.012131f
C21499 VDD.n3951 VSS 0.012131f
C21500 VDD.n3952 VSS 0.012131f
C21501 VDD.n3953 VSS 0.012131f
C21502 VDD.n3954 VSS 0.012131f
C21503 VDD.n3955 VSS 0.012131f
C21504 VDD.n3956 VSS 0.012131f
C21505 VDD.n3957 VSS 0.012131f
C21506 VDD.n3958 VSS 0.012131f
C21507 VDD.n3959 VSS 0.012131f
C21508 VDD.n3960 VSS 0.012131f
C21509 VDD.n3961 VSS 0.012131f
C21510 VDD.n3962 VSS 0.012131f
C21511 VDD.n3963 VSS 0.012131f
C21512 VDD.n3964 VSS 0.012131f
C21513 VDD.n3965 VSS 0.012131f
C21514 VDD.n3966 VSS 0.012131f
C21515 VDD.n3967 VSS 0.012131f
C21516 VDD.n3968 VSS 0.012131f
C21517 VDD.n3969 VSS 0.012131f
C21518 VDD.n3970 VSS 0.012131f
C21519 VDD.n3971 VSS 0.012131f
C21520 VDD.n3972 VSS 0.012131f
C21521 VDD.n3973 VSS 0.012131f
C21522 VDD.n3974 VSS 0.012131f
C21523 VDD.n3975 VSS 0.012131f
C21524 VDD.n3976 VSS 0.012131f
C21525 VDD.n3977 VSS 0.012131f
C21526 VDD.n3978 VSS 0.012131f
C21527 VDD.n3979 VSS 0.012131f
C21528 VDD.n3980 VSS 0.012131f
C21529 VDD.n3981 VSS 0.012131f
C21530 VDD.n3982 VSS 0.012131f
C21531 VDD.n3983 VSS 0.012131f
C21532 VDD.n3984 VSS 0.012131f
C21533 VDD.n3985 VSS 0.012131f
C21534 VDD.n3986 VSS 0.012131f
C21535 VDD.n3987 VSS 0.012131f
C21536 VDD.n3988 VSS 0.012131f
C21537 VDD.n3989 VSS 0.012131f
C21538 VDD.n3990 VSS 0.012131f
C21539 VDD.n3991 VSS 0.012131f
C21540 VDD.n3992 VSS 0.012131f
C21541 VDD.n3993 VSS 0.012131f
C21542 VDD.n3994 VSS 0.012131f
C21543 VDD.n3995 VSS 0.012131f
C21544 VDD.n3996 VSS 0.012131f
C21545 VDD.n3997 VSS 0.012131f
C21546 VDD.n3998 VSS 0.012131f
C21547 VDD.n3999 VSS 0.012131f
C21548 VDD.n4000 VSS 0.012131f
C21549 VDD.n4001 VSS 0.012131f
C21550 VDD.n4002 VSS 0.012131f
C21551 VDD.n4003 VSS 0.012131f
C21552 VDD.n4004 VSS 0.012131f
C21553 VDD.n4005 VSS 0.012131f
C21554 VDD.n4006 VSS 0.012131f
C21555 VDD.n4007 VSS 0.012131f
C21556 VDD.n4008 VSS 0.012131f
C21557 VDD.n4009 VSS 0.012131f
C21558 VDD.n4010 VSS 0.012131f
C21559 VDD.n4011 VSS 0.012131f
C21560 VDD.n4012 VSS 0.012131f
C21561 VDD.n4013 VSS 0.012131f
C21562 VDD.n4014 VSS 0.012131f
C21563 VDD.n4015 VSS 0.012131f
C21564 VDD.n4016 VSS 0.012131f
C21565 VDD.n4017 VSS 0.012131f
C21566 VDD.n4018 VSS 0.012131f
C21567 VDD.n4019 VSS 0.012131f
C21568 VDD.n4020 VSS 0.012131f
C21569 VDD.n4021 VSS 0.012131f
C21570 VDD.n4022 VSS 0.012131f
C21571 VDD.n4023 VSS 0.012131f
C21572 VDD.n4024 VSS 0.012131f
C21573 VDD.n4025 VSS 0.012131f
C21574 VDD.n4026 VSS 0.012131f
C21575 VDD.n4027 VSS 0.012131f
C21576 VDD.n4028 VSS 0.012131f
C21577 VDD.n4029 VSS 0.012131f
C21578 VDD.n4030 VSS 0.012131f
C21579 VDD.n4031 VSS 0.012131f
C21580 VDD.n4032 VSS 0.012131f
C21581 VDD.n4033 VSS 0.012131f
C21582 VDD.n4034 VSS 0.012131f
C21583 VDD.n4035 VSS 0.012131f
C21584 VDD.n4036 VSS 0.012131f
C21585 VDD.n4037 VSS 0.012131f
C21586 VDD.n4038 VSS 0.012131f
C21587 VDD.n4039 VSS 0.012131f
C21588 VDD.n4040 VSS 0.012131f
C21589 VDD.n4041 VSS 0.012131f
C21590 VDD.n4042 VSS 0.012131f
C21591 VDD.n4043 VSS 0.012131f
C21592 VDD.n4044 VSS 0.012131f
C21593 VDD.n4045 VSS 0.012131f
C21594 VDD.n4046 VSS 0.012131f
C21595 VDD.n4047 VSS 0.012131f
C21596 VDD.n4048 VSS 0.012131f
C21597 VDD.n4049 VSS 0.012131f
C21598 VDD.n4050 VSS 0.012131f
C21599 VDD.n4051 VSS 0.012131f
C21600 VDD.n4052 VSS 0.012131f
C21601 VDD.n4053 VSS 0.012131f
C21602 VDD.n4054 VSS 0.012131f
C21603 VDD.n4055 VSS 0.012131f
C21604 VDD.n4056 VSS 0.012131f
C21605 VDD.n4057 VSS 0.012131f
C21606 VDD.n4058 VSS 0.012131f
C21607 VDD.n4059 VSS 0.012131f
C21608 VDD.n4060 VSS 0.012131f
C21609 VDD.n4061 VSS 0.012131f
C21610 VDD.n4062 VSS 0.012131f
C21611 VDD.n4063 VSS 0.012131f
C21612 VDD.n4064 VSS 0.012131f
C21613 VDD.n4065 VSS 0.012131f
C21614 VDD.n4066 VSS 0.012131f
C21615 VDD.n4067 VSS 0.012131f
C21616 VDD.n4068 VSS 0.012131f
C21617 VDD.n4069 VSS 0.012131f
C21618 VDD.n4070 VSS 0.012131f
C21619 VDD.n4071 VSS 0.012131f
C21620 VDD.n4072 VSS 0.012131f
C21621 VDD.n4073 VSS 0.012131f
C21622 VDD.n4074 VSS 0.012131f
C21623 VDD.n4075 VSS 0.012131f
C21624 VDD.n4076 VSS 0.012131f
C21625 VDD.n4077 VSS 0.012131f
C21626 VDD.n4078 VSS 0.012131f
C21627 VDD.n4079 VSS 0.012131f
C21628 VDD.n4080 VSS 0.012131f
C21629 VDD.n4081 VSS 0.012131f
C21630 VDD.n4082 VSS 0.012131f
C21631 VDD.n4083 VSS 0.012131f
C21632 VDD.n4084 VSS 0.012131f
C21633 VDD.n4085 VSS 0.012131f
C21634 VDD.n4086 VSS 0.012131f
C21635 VDD.n4087 VSS 0.012131f
C21636 VDD.n4088 VSS 0.012131f
C21637 VDD.n4089 VSS 0.012131f
C21638 VDD.n4090 VSS 0.012131f
C21639 VDD.n4091 VSS 0.012131f
C21640 VDD.n4092 VSS 0.012131f
C21641 VDD.n4093 VSS 0.012131f
C21642 VDD.n4094 VSS 0.012131f
C21643 VDD.n4095 VSS 0.012131f
C21644 VDD.n4096 VSS 0.012131f
C21645 VDD.n4097 VSS 0.012131f
C21646 VDD.n4098 VSS 0.012131f
C21647 VDD.n4099 VSS 0.012131f
C21648 VDD.n4100 VSS 0.012131f
C21649 VDD.n4101 VSS 0.012131f
C21650 VDD.n4102 VSS 0.012131f
C21651 VDD.n4103 VSS 0.012131f
C21652 VDD.n4104 VSS 0.012131f
C21653 VDD.n4105 VSS 0.012131f
C21654 VDD.n4106 VSS 0.012131f
C21655 VDD.n4107 VSS 0.012131f
C21656 VDD.n4108 VSS 0.012131f
C21657 VDD.n4109 VSS 0.012131f
C21658 VDD.n4110 VSS 0.012131f
C21659 VDD.n4111 VSS 0.012131f
C21660 VDD.n4112 VSS 0.012131f
C21661 VDD.n4113 VSS 0.012131f
C21662 VDD.n4114 VSS 0.012131f
C21663 VDD.n4115 VSS 0.012131f
C21664 VDD.n4116 VSS 0.012131f
C21665 VDD.n4117 VSS 0.012131f
C21666 VDD.n4118 VSS 0.012131f
C21667 VDD.n4119 VSS 0.012131f
C21668 VDD.n4120 VSS 0.012131f
C21669 VDD.n4121 VSS 0.012131f
C21670 VDD.n4122 VSS 0.012131f
C21671 VDD.n4123 VSS 0.012131f
C21672 VDD.n4124 VSS 0.012131f
C21673 VDD.n4125 VSS 0.012131f
C21674 VDD.n4126 VSS 0.012131f
C21675 VDD.n4127 VSS 0.012131f
C21676 VDD.n4128 VSS 0.012131f
C21677 VDD.n4129 VSS 0.012131f
C21678 VDD.n4130 VSS 0.012131f
C21679 VDD.n4131 VSS 0.012131f
C21680 VDD.n4132 VSS 0.012131f
C21681 VDD.n4133 VSS 0.012131f
C21682 VDD.n4134 VSS 0.012131f
C21683 VDD.n4135 VSS 0.012131f
C21684 VDD.n4136 VSS 0.012131f
C21685 VDD.n4137 VSS 0.012131f
C21686 VDD.n4138 VSS 0.012131f
C21687 VDD.n4139 VSS 0.012131f
C21688 VDD.n4140 VSS 0.012131f
C21689 VDD.n4141 VSS 0.012131f
C21690 VDD.n4142 VSS 0.012131f
C21691 VDD.n4143 VSS 0.012131f
C21692 VDD.n4144 VSS 0.012131f
C21693 VDD.n4145 VSS 0.012131f
C21694 VDD.n4146 VSS 0.012131f
C21695 VDD.n4147 VSS 0.012131f
C21696 VDD.n4148 VSS 0.012131f
C21697 VDD.n4149 VSS 0.012131f
C21698 VDD.n4150 VSS 0.012131f
C21699 VDD.n4151 VSS 0.012131f
C21700 VDD.n4152 VSS 0.012131f
C21701 VDD.n4153 VSS 0.012131f
C21702 VDD.n4154 VSS 0.012131f
C21703 VDD.n4155 VSS 0.012131f
C21704 VDD.n4156 VSS 0.012131f
C21705 VDD.n4157 VSS 0.012131f
C21706 VDD.n4158 VSS 0.012131f
C21707 VDD.n4159 VSS 0.012131f
C21708 VDD.n4160 VSS 0.012131f
C21709 VDD.n4161 VSS 0.012131f
C21710 VDD.n4162 VSS 0.012131f
C21711 VDD.n4163 VSS 0.012131f
C21712 VDD.n4164 VSS 0.012131f
C21713 VDD.n4165 VSS 0.012131f
C21714 VDD.n4166 VSS 0.012131f
C21715 VDD.n4167 VSS 0.012131f
C21716 VDD.n4168 VSS 0.012131f
C21717 VDD.n4169 VSS 0.012131f
C21718 VDD.n4170 VSS 0.012131f
C21719 VDD.n4171 VSS 0.012131f
C21720 VDD.n4172 VSS 0.012131f
C21721 VDD.n4173 VSS 0.012131f
C21722 VDD.n4174 VSS 0.012131f
C21723 VDD.n4175 VSS 0.012131f
C21724 VDD.n4176 VSS 0.012131f
C21725 VDD.n4177 VSS 0.012131f
C21726 VDD.n4178 VSS 0.012131f
C21727 VDD.n4179 VSS 0.012131f
C21728 VDD.n4180 VSS 0.012131f
C21729 VDD.n4181 VSS 0.012131f
C21730 VDD.n4182 VSS 0.012131f
C21731 VDD.n4183 VSS 0.012131f
C21732 VDD.n4184 VSS 0.012131f
C21733 VDD.n4185 VSS 0.012131f
C21734 VDD.n4186 VSS 0.012131f
C21735 VDD.n4187 VSS 0.012131f
C21736 VDD.n4188 VSS 0.012131f
C21737 VDD.n4189 VSS 0.012131f
C21738 VDD.n4190 VSS 0.012131f
C21739 VDD.n4191 VSS 0.012131f
C21740 VDD.n4192 VSS 0.012131f
C21741 VDD.n4193 VSS 0.012131f
C21742 VDD.n4194 VSS 0.012131f
C21743 VDD.n4195 VSS 0.012131f
C21744 VDD.n4196 VSS 0.012131f
C21745 VDD.n4197 VSS 0.012131f
C21746 VDD.n4198 VSS 0.012131f
C21747 VDD.n4199 VSS 0.012131f
C21748 VDD.n4200 VSS 0.012131f
C21749 VDD.n4201 VSS 0.012131f
C21750 VDD.n4202 VSS 0.012131f
C21751 VDD.n4203 VSS 0.012131f
C21752 VDD.n4204 VSS 0.012131f
C21753 VDD.n4205 VSS 0.012131f
C21754 VDD.n4206 VSS 0.012131f
C21755 VDD.n4207 VSS 0.012131f
C21756 VDD.n4208 VSS 0.012131f
C21757 VDD.n4209 VSS 0.012131f
C21758 VDD.n4210 VSS 0.012131f
C21759 VDD.n4211 VSS 0.012131f
C21760 VDD.n4212 VSS 0.012131f
C21761 VDD.n4213 VSS 0.012131f
C21762 VDD.n4214 VSS 0.012131f
C21763 VDD.n4215 VSS 0.012131f
C21764 VDD.n4216 VSS 0.012131f
C21765 VDD.n4217 VSS 0.012131f
C21766 VDD.n4218 VSS 0.012131f
C21767 VDD.n4219 VSS 0.012131f
C21768 VDD.n4220 VSS 0.012131f
C21769 VDD.n4221 VSS 0.012131f
C21770 VDD.n4222 VSS 0.012131f
C21771 VDD.n4223 VSS 0.012131f
C21772 VDD.n4224 VSS 0.012131f
C21773 VDD.n4225 VSS 0.012131f
C21774 VDD.n4226 VSS 0.012131f
C21775 VDD.n4227 VSS 0.012131f
C21776 VDD.n4228 VSS 0.012131f
C21777 VDD.n4229 VSS 0.012131f
C21778 VDD.n4230 VSS 0.012131f
C21779 VDD.n4231 VSS 0.012131f
C21780 VDD.n4232 VSS 0.012131f
C21781 VDD.n4233 VSS 0.012131f
C21782 VDD.n4234 VSS 0.012131f
C21783 VDD.n4235 VSS 0.012131f
C21784 VDD.n4236 VSS 0.012131f
C21785 VDD.n4237 VSS 0.012131f
C21786 VDD.n4238 VSS 0.012131f
C21787 VDD.n4239 VSS 0.012131f
C21788 VDD.n4240 VSS 0.012131f
C21789 VDD.n4241 VSS 0.012131f
C21790 VDD.n4242 VSS 0.012131f
C21791 VDD.n4243 VSS 0.012131f
C21792 VDD.n4244 VSS 0.012131f
C21793 VDD.n4245 VSS 0.012131f
C21794 VDD.n4246 VSS 0.012131f
C21795 VDD.n4247 VSS 0.012131f
C21796 VDD.n4248 VSS 0.012131f
C21797 VDD.n4249 VSS 0.012131f
C21798 VDD.n4250 VSS 0.012131f
C21799 VDD.n4251 VSS 0.012131f
C21800 VDD.n4252 VSS 0.012131f
C21801 VDD.n4253 VSS 0.012131f
C21802 VDD.n4254 VSS 0.012131f
C21803 VDD.n4255 VSS 0.012131f
C21804 VDD.n4256 VSS 0.012131f
C21805 VDD.n4257 VSS 0.012131f
C21806 VDD.n4258 VSS 0.012131f
C21807 VDD.n4259 VSS 0.012131f
C21808 VDD.n4260 VSS 0.012131f
C21809 VDD.n4261 VSS 0.012131f
C21810 VDD.n4262 VSS 0.012131f
C21811 VDD.n4263 VSS 0.012131f
C21812 VDD.n4264 VSS 0.012131f
C21813 VDD.n4265 VSS 0.012131f
C21814 VDD.n4266 VSS 0.012131f
C21815 VDD.n4267 VSS 0.012131f
C21816 VDD.n4268 VSS 0.012131f
C21817 VDD.n4269 VSS 0.012131f
C21818 VDD.n4270 VSS 0.012131f
C21819 VDD.n4271 VSS 0.012131f
C21820 VDD.n4272 VSS 0.012131f
C21821 VDD.n4273 VSS 0.012131f
C21822 VDD.n4274 VSS 0.012131f
C21823 VDD.n4275 VSS 0.012131f
C21824 VDD.n4276 VSS 0.012131f
C21825 VDD.n4277 VSS 0.012131f
C21826 VDD.n4278 VSS 0.012131f
C21827 VDD.n4279 VSS 0.012131f
C21828 VDD.n4280 VSS 0.012131f
C21829 VDD.n4281 VSS 0.012131f
C21830 VDD.n4282 VSS 0.012131f
C21831 VDD.n4283 VSS 0.012131f
C21832 VDD.n4284 VSS 0.012131f
C21833 VDD.n4285 VSS 0.012131f
C21834 VDD.n4286 VSS 0.012131f
C21835 VDD.n4287 VSS 0.012131f
C21836 VDD.n4288 VSS 0.012131f
C21837 VDD.n4289 VSS 0.012131f
C21838 VDD.n4290 VSS 0.012131f
C21839 VDD.n4291 VSS 0.012131f
C21840 VDD.n4292 VSS 0.012131f
C21841 VDD.n4293 VSS 0.012131f
C21842 VDD.n4294 VSS 0.012131f
C21843 VDD.n4295 VSS 0.012131f
C21844 VDD.n4296 VSS 0.012131f
C21845 VDD.n4297 VSS 0.012131f
C21846 VDD.n4298 VSS 0.012131f
C21847 VDD.n4299 VSS 0.012131f
C21848 VDD.n4300 VSS 0.012131f
C21849 VDD.n4301 VSS 0.012131f
C21850 VDD.n4302 VSS 0.012131f
C21851 VDD.n4303 VSS 0.012131f
C21852 VDD.n4304 VSS 0.012131f
C21853 VDD.n4305 VSS 0.012131f
C21854 VDD.n4306 VSS 0.012131f
C21855 VDD.n4307 VSS 0.012131f
C21856 VDD.n4308 VSS 0.012131f
C21857 VDD.n4309 VSS 0.012131f
C21858 VDD.n4310 VSS 0.012131f
C21859 VDD.n4311 VSS 0.012131f
C21860 VDD.n4312 VSS 0.012131f
C21861 VDD.n4313 VSS 0.012131f
C21862 VDD.n4314 VSS 0.012131f
C21863 VDD.n4315 VSS 0.012131f
C21864 VDD.n4316 VSS 0.012131f
C21865 VDD.n4317 VSS 0.012131f
C21866 VDD.n4318 VSS 0.012131f
C21867 VDD.n4319 VSS 0.012131f
C21868 VDD.n4320 VSS 0.012131f
C21869 VDD.n4321 VSS 0.012131f
C21870 VDD.n4322 VSS 0.012131f
C21871 VDD.n4323 VSS 0.012131f
C21872 VDD.n4324 VSS 0.012131f
C21873 VDD.n4325 VSS 0.012131f
C21874 VDD.n4326 VSS 0.012131f
C21875 VDD.n4327 VSS 0.012131f
C21876 VDD.n4328 VSS 0.012131f
C21877 VDD.n4329 VSS 0.012131f
C21878 VDD.n4330 VSS 0.012131f
C21879 VDD.n4331 VSS 0.012131f
C21880 VDD.n4332 VSS 0.012131f
C21881 VDD.n4333 VSS 0.012131f
C21882 VDD.n4334 VSS 0.012131f
C21883 VDD.n4335 VSS 0.012131f
C21884 VDD.n4336 VSS 0.012131f
C21885 VDD.n4337 VSS 0.012131f
C21886 VDD.n4338 VSS 0.012131f
C21887 VDD.n4339 VSS 0.012131f
C21888 VDD.n4340 VSS 0.012131f
C21889 VDD.n4341 VSS 0.012131f
C21890 VDD.n4342 VSS 0.012131f
C21891 VDD.n4343 VSS 0.012131f
C21892 VDD.n4344 VSS 0.012131f
C21893 VDD.n4345 VSS 0.012131f
C21894 VDD.n4346 VSS 0.012131f
C21895 VDD.n4347 VSS 0.012131f
C21896 VDD.n4348 VSS 0.012131f
C21897 VDD.n4349 VSS 0.012131f
C21898 VDD.n4350 VSS 0.012131f
C21899 VDD.n4351 VSS 0.012131f
C21900 VDD.n4352 VSS 0.012131f
C21901 VDD.n4353 VSS 0.012131f
C21902 VDD.n4354 VSS 0.012131f
C21903 VDD.n4355 VSS 0.012131f
C21904 VDD.n4356 VSS 0.012131f
C21905 VDD.n4357 VSS 0.012131f
C21906 VDD.n4358 VSS 0.012131f
C21907 VDD.n4359 VSS 0.012131f
C21908 VDD.n4360 VSS 0.012131f
C21909 VDD.n4361 VSS 0.012131f
C21910 VDD.n4362 VSS 0.012131f
C21911 VDD.n4363 VSS 0.012131f
C21912 VDD.n4364 VSS 0.012131f
C21913 VDD.n4365 VSS 0.012131f
C21914 VDD.n4366 VSS 0.012131f
C21915 VDD.n4367 VSS 0.012131f
C21916 VDD.n4368 VSS 0.012131f
C21917 VDD.n4369 VSS 0.012131f
C21918 VDD.n4370 VSS 0.012131f
C21919 VDD.n4371 VSS 0.012131f
C21920 VDD.n4372 VSS 0.012131f
C21921 VDD.n4373 VSS 0.012131f
C21922 VDD.n4374 VSS 0.012131f
C21923 VDD.n4375 VSS 0.012131f
C21924 VDD.n4376 VSS 0.012131f
C21925 VDD.n4377 VSS 0.012131f
C21926 VDD.n4378 VSS 0.012131f
C21927 VDD.n4379 VSS 0.012131f
C21928 VDD.n4380 VSS 0.012131f
C21929 VDD.n4381 VSS 0.012131f
C21930 VDD.n4382 VSS 0.012131f
C21931 VDD.n4383 VSS 0.012131f
C21932 VDD.n4384 VSS 0.012131f
C21933 VDD.n4385 VSS 0.012131f
C21934 VDD.n4386 VSS 0.012131f
C21935 VDD.n4387 VSS 0.012131f
C21936 VDD.n4388 VSS 0.012131f
C21937 VDD.n4389 VSS 0.012131f
C21938 VDD.n4390 VSS 0.012131f
C21939 VDD.n4391 VSS 0.012131f
C21940 VDD.n4392 VSS 0.012131f
C21941 VDD.n4393 VSS 0.012131f
C21942 VDD.n4394 VSS 0.012131f
C21943 VDD.n4395 VSS 0.012131f
C21944 VDD.n4396 VSS 0.012131f
C21945 VDD.n4397 VSS 0.012131f
C21946 VDD.n4398 VSS 0.012131f
C21947 VDD.n4399 VSS 0.012131f
C21948 VDD.n4400 VSS 0.012131f
C21949 VDD.n4401 VSS 0.012131f
C21950 VDD.n4402 VSS 0.012131f
C21951 VDD.n4403 VSS 0.012131f
C21952 VDD.n4404 VSS 0.012131f
C21953 VDD.n4405 VSS 0.012131f
C21954 VDD.n4406 VSS 0.012131f
C21955 VDD.n4407 VSS 0.012131f
C21956 VDD.n4408 VSS 0.012131f
C21957 VDD.n4409 VSS 0.012131f
C21958 VDD.n4410 VSS 0.012131f
C21959 VDD.n4411 VSS 0.012131f
C21960 VDD.n4412 VSS 0.012131f
C21961 VDD.n4413 VSS 0.012131f
C21962 VDD.n4414 VSS 0.012131f
C21963 VDD.n4415 VSS 0.012131f
C21964 VDD.n4416 VSS 0.012131f
C21965 VDD.n4417 VSS 0.012131f
C21966 VDD.n4418 VSS 0.012131f
C21967 VDD.n4419 VSS 0.012131f
C21968 VDD.n4420 VSS 0.012131f
C21969 VDD.n4421 VSS 0.012131f
C21970 VDD.n4422 VSS 0.012131f
C21971 VDD.n4423 VSS 0.012131f
C21972 VDD.n4424 VSS 0.012131f
C21973 VDD.n4425 VSS 0.012131f
C21974 VDD.n4426 VSS 0.012131f
C21975 VDD.n4427 VSS 0.012131f
C21976 VDD.n4428 VSS 0.012131f
C21977 VDD.n4429 VSS 0.012131f
C21978 VDD.n4430 VSS 0.012131f
C21979 VDD.n4431 VSS 0.012131f
C21980 VDD.n4432 VSS 0.012131f
C21981 VDD.n4433 VSS 0.012131f
C21982 VDD.n4434 VSS 0.012131f
C21983 VDD.n4435 VSS 0.012131f
C21984 VDD.n4436 VSS 0.012131f
C21985 VDD.n4437 VSS 0.012131f
C21986 VDD.n4438 VSS 0.012131f
C21987 VDD.n4439 VSS 0.012131f
C21988 VDD.n4440 VSS 0.012131f
C21989 VDD.n4441 VSS 0.012131f
C21990 VDD.n4442 VSS 0.012131f
C21991 VDD.n4443 VSS 0.012131f
C21992 VDD.n4444 VSS 0.012131f
C21993 VDD.n4445 VSS 0.012131f
C21994 VDD.n4446 VSS 0.012131f
C21995 VDD.n4447 VSS 0.012131f
C21996 VDD.n4448 VSS 0.012131f
C21997 VDD.n4449 VSS 0.012131f
C21998 VDD.n4450 VSS 0.012131f
C21999 VDD.n4451 VSS 0.012131f
C22000 VDD.n4452 VSS 0.012131f
C22001 VDD.n4453 VSS 0.012131f
C22002 VDD.n4454 VSS 0.012131f
C22003 VDD.n4455 VSS 0.012131f
C22004 VDD.n4456 VSS 0.012131f
C22005 VDD.n4457 VSS 0.012131f
C22006 VDD.n4458 VSS 0.012131f
C22007 VDD.n4459 VSS 0.012131f
C22008 VDD.n4460 VSS 0.012131f
C22009 VDD.n4461 VSS 0.012131f
C22010 VDD.n4462 VSS 0.012131f
C22011 VDD.n4463 VSS 0.012131f
C22012 VDD.n4464 VSS 0.012131f
C22013 VDD.n4465 VSS 0.012131f
C22014 VDD.n4466 VSS 0.012131f
C22015 VDD.n4467 VSS 0.012131f
C22016 VDD.n4468 VSS 0.012131f
C22017 VDD.n4469 VSS 0.012131f
C22018 VDD.n4470 VSS 0.012131f
C22019 VDD.n4471 VSS 0.012131f
C22020 VDD.n4472 VSS 0.012131f
C22021 VDD.n4473 VSS 0.012131f
C22022 VDD.n4474 VSS 0.012131f
C22023 VDD.n4475 VSS 0.012131f
C22024 VDD.n4476 VSS 0.012131f
C22025 VDD.n4477 VSS 0.012131f
C22026 VDD.n4478 VSS 0.012131f
C22027 VDD.n4479 VSS 0.012131f
C22028 VDD.n4480 VSS 0.012131f
C22029 VDD.n4481 VSS 0.012131f
C22030 VDD.n4482 VSS 0.012131f
C22031 VDD.n4483 VSS 0.012131f
C22032 VDD.n4484 VSS 0.012131f
C22033 VDD.n4485 VSS 0.012131f
C22034 VDD.n4486 VSS 0.012131f
C22035 VDD.n4487 VSS 0.012131f
C22036 VDD.n4488 VSS 0.012131f
C22037 VDD.n4489 VSS 0.012131f
C22038 VDD.n4490 VSS 0.012131f
C22039 VDD.n4491 VSS 0.012131f
C22040 VDD.n4492 VSS 0.012131f
C22041 VDD.n4493 VSS 0.012131f
C22042 VDD.n4494 VSS 0.012131f
C22043 VDD.n4495 VSS 0.012131f
C22044 VDD.n4496 VSS 0.012131f
C22045 VDD.n4497 VSS 0.012131f
C22046 VDD.n4498 VSS 0.012131f
C22047 VDD.n4499 VSS 0.012131f
C22048 VDD.n4500 VSS 0.012131f
C22049 VDD.n4501 VSS 0.012131f
C22050 VDD.n4502 VSS 0.012131f
C22051 VDD.n4503 VSS 0.012131f
C22052 VDD.n4504 VSS 0.012131f
C22053 VDD.n4505 VSS 0.012131f
C22054 VDD.n4506 VSS 0.012131f
C22055 VDD.n4507 VSS 0.012131f
C22056 VDD.n4508 VSS 0.012131f
C22057 VDD.n4509 VSS 0.012131f
C22058 VDD.n4510 VSS 0.012131f
C22059 VDD.n4511 VSS 0.012131f
C22060 VDD.n4512 VSS 0.012131f
C22061 VDD.n4513 VSS 0.012131f
C22062 VDD.n4514 VSS 0.012131f
C22063 VDD.n4515 VSS 0.012131f
C22064 VDD.n4516 VSS 0.012131f
C22065 VDD.n4517 VSS 0.012131f
C22066 VDD.n4518 VSS 0.012131f
C22067 VDD.n4519 VSS 0.012131f
C22068 VDD.n4520 VSS 0.012131f
C22069 VDD.n4521 VSS 0.012131f
C22070 VDD.n4522 VSS 0.012131f
C22071 VDD.n4523 VSS 0.012131f
C22072 VDD.n4524 VSS 0.012131f
C22073 VDD.n4525 VSS 0.012131f
C22074 VDD.n4526 VSS 0.012131f
C22075 VDD.n4527 VSS 0.012131f
C22076 VDD.n4528 VSS 0.012131f
C22077 VDD.n4529 VSS 0.012131f
C22078 VDD.n4530 VSS 0.012131f
C22079 VDD.n4531 VSS 0.012131f
C22080 VDD.n4532 VSS 0.012131f
C22081 VDD.n4533 VSS 0.012131f
C22082 VDD.n4534 VSS 0.012131f
C22083 VDD.n4535 VSS 0.012131f
C22084 VDD.n4536 VSS 0.012131f
C22085 VDD.n4537 VSS 0.012131f
C22086 VDD.n4538 VSS 0.012131f
C22087 VDD.n4539 VSS 0.012131f
C22088 VDD.n4540 VSS 0.012131f
C22089 VDD.n4541 VSS 0.012131f
C22090 VDD.n4542 VSS 0.012131f
C22091 VDD.n4543 VSS 0.012131f
C22092 VDD.n4544 VSS 0.012131f
C22093 VDD.n4545 VSS 0.012131f
C22094 VDD.n4546 VSS 0.012131f
C22095 VDD.n4547 VSS 0.012131f
C22096 VDD.n4548 VSS 0.012131f
C22097 VDD.n4549 VSS 0.012131f
C22098 VDD.n4550 VSS 0.012131f
C22099 VDD.n4551 VSS 0.012131f
C22100 VDD.n4552 VSS 0.012131f
C22101 VDD.n4553 VSS 0.012131f
C22102 VDD.n4554 VSS 0.012131f
C22103 VDD.n4555 VSS 0.012131f
C22104 VDD.n4556 VSS 0.012131f
C22105 VDD.n4557 VSS 0.012131f
C22106 VDD.n4558 VSS 0.012131f
C22107 VDD.n4559 VSS 0.012131f
C22108 VDD.n4560 VSS 0.012131f
C22109 VDD.n4561 VSS 0.012131f
C22110 VDD.n4562 VSS 0.012131f
C22111 VDD.n4563 VSS 0.012131f
C22112 VDD.n4564 VSS 0.012131f
C22113 VDD.n4565 VSS 0.012131f
C22114 VDD.n4566 VSS 0.012131f
C22115 VDD.n4567 VSS 0.012131f
C22116 VDD.n4568 VSS 0.012131f
C22117 VDD.n4569 VSS 0.012131f
C22118 VDD.n4570 VSS 0.012131f
C22119 VDD.n4571 VSS 0.012131f
C22120 VDD.n4572 VSS 0.012131f
C22121 VDD.n4573 VSS 0.012131f
C22122 VDD.n4574 VSS 0.012131f
C22123 VDD.n4575 VSS 0.012131f
C22124 VDD.n4576 VSS 0.012131f
C22125 VDD.n4577 VSS 0.012131f
C22126 VDD.n4578 VSS 0.012131f
C22127 VDD.n4579 VSS 0.012131f
C22128 VDD.n4580 VSS 0.012131f
C22129 VDD.n4581 VSS 0.012131f
C22130 VDD.n4582 VSS 0.012131f
C22131 VDD.n4583 VSS 0.012131f
C22132 VDD.n4584 VSS 0.012131f
C22133 VDD.n4585 VSS 0.012131f
C22134 VDD.n4586 VSS 0.012131f
C22135 VDD.n4587 VSS 0.012131f
C22136 VDD.n4588 VSS 0.012131f
C22137 VDD.n4589 VSS 0.008526f
C22138 VDD.n4590 VSS 0.008222f
C22139 VDD.n4591 VSS 0.010165f
C22140 VDD.n4592 VSS 0.012131f
C22141 VDD.n4593 VSS 0.012131f
C22142 VDD.n4594 VSS 0.012131f
C22143 VDD.n4595 VSS 0.012131f
C22144 VDD.n4596 VSS 0.012131f
C22145 VDD.n4597 VSS 0.006065f
C22146 VDD.n4598 VSS 0.012131f
C22147 VDD.n4599 VSS 0.012131f
C22148 VDD.n4600 VSS 0.012131f
C22149 VDD.n4601 VSS 0.012131f
C22150 VDD.n4602 VSS 0.012131f
C22151 VDD.n4603 VSS 0.012131f
C22152 VDD.n4604 VSS 0.012131f
C22153 VDD.n4605 VSS 0.012131f
C22154 VDD.n4606 VSS 0.012131f
C22155 VDD.n4607 VSS 0.012131f
C22156 VDD.n4608 VSS 0.012131f
C22157 VDD.n4609 VSS 0.012131f
C22158 VDD.n4610 VSS 0.012131f
C22159 VDD.n4611 VSS 0.012131f
C22160 VDD.n4612 VSS 0.012131f
C22161 VDD.n4613 VSS 0.012131f
C22162 VDD.n4614 VSS 0.012131f
C22163 VDD.n4615 VSS 0.012131f
C22164 VDD.n4616 VSS 0.012131f
C22165 VDD.n4617 VSS 0.012131f
C22166 VDD.n4618 VSS 0.012131f
C22167 VDD.n4619 VSS 0.012131f
C22168 VDD.n4620 VSS 0.012131f
C22169 VDD.n4621 VSS 0.012131f
C22170 VDD.n4622 VSS 0.012131f
C22171 VDD.n4623 VSS 0.012131f
C22172 VDD.n4624 VSS 0.012131f
C22173 VDD.n4625 VSS 0.012131f
C22174 VDD.n4626 VSS 0.012131f
C22175 VDD.n4627 VSS 0.012131f
C22176 VDD.n4628 VSS 0.012131f
C22177 VDD.n4629 VSS 0.012131f
C22178 VDD.n4630 VSS 0.012131f
C22179 VDD.n4631 VSS 0.012131f
C22180 VDD.n4632 VSS 0.012131f
C22181 VDD.n4633 VSS 0.012131f
C22182 VDD.n4634 VSS 0.012131f
C22183 VDD.n4635 VSS 0.012131f
C22184 VDD.n4636 VSS 0.012131f
C22185 VDD.n4637 VSS 0.012131f
C22186 VDD.n4638 VSS 0.012131f
C22187 VDD.n4639 VSS 0.012131f
C22188 VDD.n4640 VSS 0.012131f
C22189 VDD.n4641 VSS 0.012131f
C22190 VDD.n4642 VSS 0.012131f
C22191 VDD.n4643 VSS 0.012131f
C22192 VDD.n4644 VSS 0.012131f
C22193 VDD.n4645 VSS 0.012131f
C22194 VDD.n4646 VSS 0.012131f
C22195 VDD.n4647 VSS 0.012131f
C22196 VDD.n4648 VSS 0.012131f
C22197 VDD.n4649 VSS 0.012131f
C22198 VDD.n4650 VSS 0.012131f
C22199 VDD.n4651 VSS 0.012131f
C22200 VDD.n4652 VSS 0.012131f
C22201 VDD.n4653 VSS 0.012131f
C22202 VDD.n4654 VSS 0.012131f
C22203 VDD.n4655 VSS 0.012131f
C22204 VDD.n4656 VSS 0.012131f
C22205 VDD.n4657 VSS 0.012131f
C22206 VDD.n4658 VSS 0.012131f
C22207 VDD.n4659 VSS 0.012131f
C22208 VDD.n4660 VSS 0.012131f
C22209 VDD.n4661 VSS 0.012131f
C22210 VDD.n4662 VSS 0.012131f
C22211 VDD.n4663 VSS 0.012131f
C22212 VDD.n4664 VSS 0.012131f
C22213 VDD.n4665 VSS 0.012131f
C22214 VDD.n4666 VSS 0.012131f
C22215 VDD.n4667 VSS 0.012131f
C22216 VDD.n4668 VSS 0.012131f
C22217 VDD.n4669 VSS 0.012131f
C22218 VDD.n4670 VSS 0.012131f
C22219 VDD.n4671 VSS 0.012131f
C22220 VDD.n4672 VSS 0.012131f
C22221 VDD.n4673 VSS 0.012131f
C22222 VDD.n4674 VSS 0.012131f
C22223 VDD.n4675 VSS 0.012131f
C22224 VDD.n4676 VSS 0.012131f
C22225 VDD.n4677 VSS 0.012131f
C22226 VDD.n4678 VSS 0.012131f
C22227 VDD.n4679 VSS 0.012131f
C22228 VDD.n4680 VSS 0.012131f
C22229 VDD.n4681 VSS 0.012131f
C22230 VDD.n4682 VSS 0.012131f
C22231 VDD.n4683 VSS 0.012131f
C22232 VDD.n4684 VSS 0.012131f
C22233 VDD.n4685 VSS 0.012131f
C22234 VDD.n4686 VSS 0.012131f
C22235 VDD.n4687 VSS 0.012131f
C22236 VDD.n4688 VSS 0.012131f
C22237 VDD.n4689 VSS 0.012131f
C22238 VDD.n4690 VSS 0.012131f
C22239 VDD.n4691 VSS 0.012131f
C22240 VDD.n4692 VSS 0.012131f
C22241 VDD.n4693 VSS 0.012131f
C22242 VDD.n4694 VSS 0.012131f
C22243 VDD.n4695 VSS 0.012131f
C22244 VDD.n4696 VSS 0.012131f
C22245 VDD.n4697 VSS 0.032533f
C22246 VDD.n4698 VSS 0.012131f
C22247 VDD.n4699 VSS 0.012131f
C22248 VDD.n4700 VSS 0.012131f
C22249 VDD.n4701 VSS 0.012131f
C22250 VDD.n4702 VSS 0.012131f
C22251 VDD.n4703 VSS 0.012131f
C22252 VDD.n4704 VSS 0.012131f
C22253 VDD.n4705 VSS 0.012131f
C22254 VDD.n4706 VSS 0.012131f
C22255 VDD.n4707 VSS 0.012131f
C22256 VDD.n4708 VSS 0.012131f
C22257 VDD.n4709 VSS 0.012131f
C22258 VDD.n4710 VSS 0.012131f
C22259 VDD.n4711 VSS 0.012131f
C22260 VDD.n4712 VSS 0.012131f
C22261 VDD.n4713 VSS 0.012131f
C22262 VDD.n4714 VSS 0.012131f
C22263 VDD.n4715 VSS 0.012131f
C22264 VDD.n4716 VSS 0.012131f
C22265 VDD.n4717 VSS 0.012131f
C22266 VDD.n4718 VSS 0.012131f
C22267 VDD.n4719 VSS 0.012131f
C22268 VDD.n4720 VSS 0.012131f
C22269 VDD.n4721 VSS 0.012131f
C22270 VDD.n4722 VSS 0.012131f
C22271 VDD.n4723 VSS 0.012131f
C22272 VDD.n4724 VSS 0.012131f
C22273 VDD.n4725 VSS 0.012131f
C22274 VDD.n4726 VSS 0.012131f
C22275 VDD.n4727 VSS 0.012131f
C22276 VDD.n4728 VSS 0.012131f
C22277 VDD.n4729 VSS 0.012131f
C22278 VDD.n4730 VSS 0.012131f
C22279 VDD.n4731 VSS 0.012131f
C22280 VDD.n4732 VSS 0.012131f
C22281 VDD.n4733 VSS 0.012131f
C22282 VDD.n4734 VSS 0.012131f
C22283 VDD.n4735 VSS 0.012131f
C22284 VDD.n4736 VSS 0.012131f
C22285 VDD.n4737 VSS 0.012131f
C22286 VDD.n4738 VSS 0.012131f
C22287 VDD.n4739 VSS 0.012131f
C22288 VDD.n4740 VSS 0.012131f
C22289 VDD.n4741 VSS 0.012131f
C22290 VDD.n4742 VSS 0.012131f
C22291 VDD.n4743 VSS 0.012131f
C22292 VDD.n4744 VSS 0.012131f
C22293 VDD.n4745 VSS 0.012131f
C22294 VDD.n4746 VSS 0.012131f
C22295 VDD.n4747 VSS 0.012131f
C22296 VDD.n4748 VSS 0.012131f
C22297 VDD.n4749 VSS 0.012131f
C22298 VDD.n4750 VSS 0.012131f
C22299 VDD.n4751 VSS 0.012131f
C22300 VDD.n4752 VSS 0.012131f
C22301 VDD.n4753 VSS 0.012131f
C22302 VDD.n4754 VSS 0.012131f
C22303 VDD.n4755 VSS 0.012131f
C22304 VDD.n4756 VSS 0.012131f
C22305 VDD.n4757 VSS 0.012131f
C22306 VDD.n4758 VSS 0.012131f
C22307 VDD.n4759 VSS 0.012131f
C22308 VDD.n4760 VSS 0.012131f
C22309 VDD.n4761 VSS 0.012131f
C22310 VDD.n4762 VSS 0.012131f
C22311 VDD.n4763 VSS 0.012131f
C22312 VDD.n4764 VSS 0.012131f
C22313 VDD.n4765 VSS 0.012131f
C22314 VDD.n4766 VSS 0.012131f
C22315 VDD.n4767 VSS 0.012131f
C22316 VDD.n4768 VSS 0.012131f
C22317 VDD.n4769 VSS 0.012131f
C22318 VDD.n4770 VSS 0.012131f
C22319 VDD.n4771 VSS 0.012131f
C22320 VDD.n4772 VSS 0.012131f
C22321 VDD.n4773 VSS 0.012131f
C22322 VDD.n4774 VSS 0.012131f
C22323 VDD.n4775 VSS 0.012131f
C22324 VDD.n4776 VSS 0.012131f
C22325 VDD.n4777 VSS 0.012131f
C22326 VDD.n4778 VSS 0.012131f
C22327 VDD.n4779 VSS 0.012131f
C22328 VDD.n4780 VSS 0.012131f
C22329 VDD.n4781 VSS 0.012131f
C22330 VDD.n4782 VSS 0.012131f
C22331 VDD.n4783 VSS 0.012131f
C22332 VDD.n4784 VSS 0.012131f
C22333 VDD.n4785 VSS 0.012131f
C22334 VDD.n4786 VSS 0.012131f
C22335 VDD.n4787 VSS 0.012131f
C22336 VDD.n4788 VSS 0.012131f
C22337 VDD.n4789 VSS 0.012131f
C22338 VDD.n4790 VSS 0.012131f
C22339 VDD.n4791 VSS 0.012131f
C22340 VDD.n4792 VSS 0.012131f
C22341 VDD.n4793 VSS 0.012131f
C22342 VDD.n4794 VSS 0.012131f
C22343 VDD.n4795 VSS 0.012131f
C22344 VDD.n4796 VSS 0.012131f
C22345 VDD.n4797 VSS 0.012131f
C22346 VDD.n4798 VSS 0.012131f
C22347 VDD.n4799 VSS 0.012131f
C22348 VDD.n4800 VSS 0.012131f
C22349 VDD.n4801 VSS 0.012131f
C22350 VDD.n4802 VSS 0.012131f
C22351 VDD.n4803 VSS 0.012131f
C22352 VDD.n4804 VSS 0.012131f
C22353 VDD.n4805 VSS 0.012131f
C22354 VDD.n4806 VSS 0.012131f
C22355 VDD.n4807 VSS 0.012131f
C22356 VDD.n4808 VSS 0.012131f
C22357 VDD.n4809 VSS 0.012131f
C22358 VDD.n4810 VSS 0.012131f
C22359 VDD.n4811 VSS 0.012131f
C22360 VDD.n4812 VSS 0.012131f
C22361 VDD.n4813 VSS 0.012131f
C22362 VDD.n4814 VSS 0.012131f
C22363 VDD.n4815 VSS 0.012131f
C22364 VDD.n4816 VSS 0.012131f
C22365 VDD.n4817 VSS 0.012131f
C22366 VDD.n4818 VSS 0.012131f
C22367 VDD.n4819 VSS 0.012131f
C22368 VDD.n4820 VSS 0.012131f
C22369 VDD.n4821 VSS 0.012131f
C22370 VDD.n4822 VSS 0.012131f
C22371 VDD.n4823 VSS 0.012131f
C22372 VDD.n4824 VSS 0.012131f
C22373 VDD.n4825 VSS 0.012131f
C22374 VDD.n4826 VSS 0.012131f
C22375 VDD.n4827 VSS 0.012131f
C22376 VDD.n4828 VSS 0.012131f
C22377 VDD.n4829 VSS 0.012131f
C22378 VDD.n4830 VSS 0.012131f
C22379 VDD.n4831 VSS 0.012131f
C22380 VDD.n4832 VSS 0.012131f
C22381 VDD.n4833 VSS 0.012131f
C22382 VDD.n4834 VSS 0.012131f
C22383 VDD.n4835 VSS 0.012131f
C22384 VDD.n4836 VSS 0.012131f
C22385 VDD.n4837 VSS 0.012131f
C22386 VDD.n4838 VSS 0.012131f
C22387 VDD.n4839 VSS 0.012131f
C22388 VDD.n4840 VSS 0.012131f
C22389 VDD.n4841 VSS 0.012131f
C22390 VDD.n4842 VSS 0.012131f
C22391 VDD.n4843 VSS 0.012131f
C22392 VDD.n4844 VSS 0.012131f
C22393 VDD.n4845 VSS 0.012131f
C22394 VDD.n4846 VSS 0.012131f
C22395 VDD.n4847 VSS 0.012131f
C22396 VDD.n4848 VSS 0.012131f
C22397 VDD.n4849 VSS 0.012131f
C22398 VDD.n4850 VSS 0.012131f
C22399 VDD.n4851 VSS 0.012131f
C22400 VDD.n4852 VSS 0.012131f
C22401 VDD.n4853 VSS 0.012131f
C22402 VDD.n4854 VSS 0.012131f
C22403 VDD.n4855 VSS 0.012131f
C22404 VDD.n4856 VSS 0.012131f
C22405 VDD.n4857 VSS 0.012131f
C22406 VDD.n4858 VSS 0.012131f
C22407 VDD.n4859 VSS 0.012131f
C22408 VDD.n4860 VSS 0.012131f
C22409 VDD.n4861 VSS 0.012131f
C22410 VDD.n4862 VSS 0.012131f
C22411 VDD.n4863 VSS 0.012131f
C22412 VDD.n4864 VSS 0.012131f
C22413 VDD.n4865 VSS 0.012131f
C22414 VDD.n4866 VSS 0.012131f
C22415 VDD.n4867 VSS 0.012131f
C22416 VDD.n4868 VSS 0.012131f
C22417 VDD.n4869 VSS 0.012131f
C22418 VDD.n4870 VSS 0.012131f
C22419 VDD.n4871 VSS 0.012131f
C22420 VDD.n4872 VSS 0.012131f
C22421 VDD.n4873 VSS 0.012131f
C22422 VDD.n4874 VSS 0.012131f
C22423 VDD.n4875 VSS 0.012131f
C22424 VDD.n4876 VSS 0.012131f
C22425 VDD.n4877 VSS 0.012131f
C22426 VDD.n4878 VSS 0.012131f
C22427 VDD.n4879 VSS 0.012131f
C22428 VDD.n4880 VSS 0.012131f
C22429 VDD.n4881 VSS 0.012131f
C22430 VDD.n4882 VSS 0.012131f
C22431 VDD.n4883 VSS 0.012131f
C22432 VDD.n4884 VSS 0.012131f
C22433 VDD.n4885 VSS 0.012131f
C22434 VDD.n4886 VSS 0.012131f
C22435 VDD.n4887 VSS 0.012131f
C22436 VDD.n4888 VSS 0.012131f
C22437 VDD.n4889 VSS 0.012131f
C22438 VDD.n4890 VSS 0.012131f
C22439 VDD.n4891 VSS 0.012131f
C22440 VDD.n4892 VSS 0.012131f
C22441 VDD.n4893 VSS 0.012131f
C22442 VDD.n4894 VSS 0.012131f
C22443 VDD.n4895 VSS 0.012131f
C22444 VDD.n4896 VSS 0.012131f
C22445 VDD.n4897 VSS 0.012131f
C22446 VDD.n4898 VSS 0.012131f
C22447 VDD.n4899 VSS 0.012131f
C22448 VDD.n4900 VSS 0.012131f
C22449 VDD.n4901 VSS 0.012131f
C22450 VDD.n4902 VSS 0.012131f
C22451 VDD.n4903 VSS 0.012131f
C22452 VDD.n4904 VSS 0.032533f
C22453 VDD.n4905 VSS 0.026861f
C22454 VDD.n4906 VSS 0.026861f
C22455 VDD.n4907 VSS 0.012131f
C22456 VDD.n4908 VSS 0.012131f
C22457 VDD.n4909 VSS 0.012131f
C22458 VDD.n4910 VSS 0.012131f
C22459 VDD.n4911 VSS 0.012131f
C22460 VDD.n4912 VSS 0.012131f
C22461 VDD.n4913 VSS 0.012131f
C22462 VDD.n4914 VSS 0.012131f
C22463 VDD.n4915 VSS 0.012131f
C22464 VDD.n4916 VSS 0.012131f
C22465 VDD.n4917 VSS 0.012131f
C22466 VDD.n4918 VSS 0.012131f
C22467 VDD.n4919 VSS 0.012131f
C22468 VDD.n4920 VSS 0.012131f
C22469 VDD.n4921 VSS 0.012131f
C22470 VDD.n4922 VSS 0.012131f
C22471 VDD.n4923 VSS 0.012131f
C22472 VDD.n4924 VSS 0.012131f
C22473 VDD.n4925 VSS 0.012131f
C22474 VDD.n4926 VSS 0.012131f
C22475 VDD.n4927 VSS 0.012131f
C22476 VDD.n4928 VSS 0.012131f
C22477 VDD.n4929 VSS 0.012131f
C22478 VDD.n4930 VSS 0.012131f
C22479 VDD.n4931 VSS 0.012131f
C22480 VDD.n4932 VSS 0.012131f
C22481 VDD.n4933 VSS 0.012131f
C22482 VDD.n4934 VSS 0.012131f
C22483 VDD.n4935 VSS 0.012131f
C22484 VDD.n4936 VSS 0.012131f
C22485 VDD.n4937 VSS 0.012131f
C22486 VDD.n4938 VSS 0.012131f
C22487 VDD.n4939 VSS 0.012131f
C22488 VDD.n4940 VSS 0.012131f
C22489 VDD.n4941 VSS 0.012131f
C22490 VDD.n4942 VSS 0.012131f
C22491 VDD.n4943 VSS 0.012131f
C22492 VDD.n4944 VSS 0.012131f
C22493 VDD.n4945 VSS 0.012131f
C22494 VDD.n4946 VSS 0.012131f
C22495 VDD.n4947 VSS 0.012131f
C22496 VDD.n4948 VSS 0.012131f
C22497 VDD.n4949 VSS 0.012131f
C22498 VDD.n4950 VSS 0.012131f
C22499 VDD.n4951 VSS 0.012131f
C22500 VDD.n4952 VSS 0.012131f
C22501 VDD.n4953 VSS 0.012131f
C22502 VDD.n4954 VSS 0.012131f
C22503 VDD.n4955 VSS 0.012131f
C22504 VDD.n4956 VSS 0.012131f
C22505 VDD.n4957 VSS 0.012131f
C22506 VDD.n4958 VSS 0.012131f
C22507 VDD.n4959 VSS 0.012131f
C22508 VDD.n4960 VSS 0.012131f
C22509 VDD.n4961 VSS 0.012131f
C22510 VDD.n4962 VSS 0.012131f
C22511 VDD.n4963 VSS 0.012131f
C22512 VDD.n4964 VSS 0.012131f
C22513 VDD.n4965 VSS 0.012131f
C22514 VDD.n4966 VSS 0.012131f
C22515 VDD.n4967 VSS 0.012131f
C22516 VDD.n4968 VSS 0.012131f
C22517 VDD.n4969 VSS 0.012131f
C22518 VDD.n4970 VSS 0.012131f
C22519 VDD.n4971 VSS 0.012131f
C22520 VDD.n4972 VSS 0.012131f
C22521 VDD.n4973 VSS 0.012131f
C22522 VDD.n4974 VSS 0.012131f
C22523 VDD.n4975 VSS 0.012131f
C22524 VDD.n4976 VSS 0.012131f
C22525 VDD.n4977 VSS 0.012131f
C22526 VDD.n4978 VSS 0.012131f
C22527 VDD.n4979 VSS 0.012131f
C22528 VDD.n4980 VSS 0.012131f
C22529 VDD.n4981 VSS 0.012131f
C22530 VDD.n4982 VSS 0.012131f
C22531 VDD.n4983 VSS 0.012131f
C22532 VDD.n4984 VSS 0.012131f
C22533 VDD.n4985 VSS 0.012131f
C22534 VDD.n4986 VSS 0.012131f
C22535 VDD.n4987 VSS 0.012131f
C22536 VDD.n4988 VSS 0.012131f
C22537 VDD.n4989 VSS 0.012131f
C22538 VDD.n4990 VSS 0.012131f
C22539 VDD.n4991 VSS 0.012131f
C22540 VDD.n4992 VSS 0.012131f
C22541 VDD.n4993 VSS 0.012131f
C22542 VDD.n4994 VSS 0.012131f
C22543 VDD.n4995 VSS 0.012131f
C22544 VDD.n4996 VSS 0.012131f
C22545 VDD.n4997 VSS 0.012131f
C22546 VDD.n4998 VSS 0.012131f
C22547 VDD.n4999 VSS 0.012131f
C22548 VDD.n5000 VSS 0.012131f
C22549 VDD.n5001 VSS 0.012131f
C22550 VDD.n5002 VSS 0.012131f
C22551 VDD.n5003 VSS 0.012131f
C22552 VDD.n5004 VSS 0.012131f
C22553 VDD.n5005 VSS 0.012131f
C22554 VDD.n5006 VSS 0.012131f
C22555 VDD.n5007 VSS 0.012131f
C22556 VDD.n5008 VSS 0.012131f
C22557 VDD.n5009 VSS 0.012131f
C22558 VDD.n5010 VSS 0.012131f
C22559 VDD.n5011 VSS 0.012131f
C22560 VDD.n5012 VSS 0.012131f
C22561 VDD.n5013 VSS 0.012131f
C22562 VDD.n5014 VSS 0.012131f
C22563 VDD.n5015 VSS 0.012131f
C22564 VDD.n5016 VSS 0.012131f
C22565 VDD.n5017 VSS 0.012131f
C22566 VDD.n5018 VSS 0.012131f
C22567 VDD.n5019 VSS 0.012131f
C22568 VDD.n5020 VSS 0.012131f
C22569 VDD.n5021 VSS 0.012131f
C22570 VDD.n5022 VSS 0.012131f
C22571 VDD.n5023 VSS 0.012131f
C22572 VDD.n5024 VSS 0.012131f
C22573 VDD.n5025 VSS 0.012131f
C22574 VDD.n5026 VSS 0.012131f
C22575 VDD.n5027 VSS 0.012131f
C22576 VDD.n5028 VSS 0.012131f
C22577 VDD.n5029 VSS 0.012131f
C22578 VDD.n5030 VSS 0.012131f
C22579 VDD.n5031 VSS 0.012131f
C22580 VDD.n5032 VSS 0.012131f
C22581 VDD.n5033 VSS 0.012131f
C22582 VDD.n5034 VSS 0.012131f
C22583 VDD.n5035 VSS 0.012131f
C22584 VDD.n5036 VSS 0.012131f
C22585 VDD.n5037 VSS 0.012131f
C22586 VDD.n5038 VSS 0.012131f
C22587 VDD.n5039 VSS 0.012131f
C22588 VDD.n5040 VSS 0.012131f
C22589 VDD.n5041 VSS 0.012131f
C22590 VDD.n5042 VSS 0.012131f
C22591 VDD.n5043 VSS 0.012131f
C22592 VDD.n5044 VSS 0.012131f
C22593 VDD.n5045 VSS 0.012131f
C22594 VDD.n5046 VSS 0.012131f
C22595 VDD.n5047 VSS 0.012131f
C22596 VDD.n5048 VSS 0.012131f
C22597 VDD.n5049 VSS 0.012131f
C22598 VDD.n5050 VSS 0.012131f
C22599 VDD.n5051 VSS 0.012131f
C22600 VDD.n5052 VSS 0.012131f
C22601 VDD.n5053 VSS 0.012131f
C22602 VDD.n5054 VSS 0.012131f
C22603 VDD.n5055 VSS 0.012131f
C22604 VDD.n5056 VSS 0.012131f
C22605 VDD.n5057 VSS 0.012131f
C22606 VDD.n5058 VSS 0.012131f
C22607 VDD.n5059 VSS 0.012131f
C22608 VDD.n5060 VSS 0.012131f
C22609 VDD.n5061 VSS 0.012131f
C22610 VDD.n5062 VSS 0.012131f
C22611 VDD.n5063 VSS 0.012131f
C22612 VDD.n5064 VSS 0.012131f
C22613 VDD.n5065 VSS 0.012131f
C22614 VDD.n5066 VSS 0.012131f
C22615 VDD.n5067 VSS 0.012131f
C22616 VDD.n5068 VSS 0.012131f
C22617 VDD.n5069 VSS 0.012131f
C22618 VDD.n5070 VSS 0.012131f
C22619 VDD.n5071 VSS 0.012131f
C22620 VDD.n5072 VSS 0.012131f
C22621 VDD.n5073 VSS 0.012131f
C22622 VDD.n5074 VSS 0.012131f
C22623 VDD.n5075 VSS 0.012131f
C22624 VDD.n5076 VSS 0.012131f
C22625 VDD.n5077 VSS 0.012131f
C22626 VDD.n5078 VSS 0.012131f
C22627 VDD.n5079 VSS 0.012131f
C22628 VDD.n5080 VSS 0.012131f
C22629 VDD.n5081 VSS 0.012131f
C22630 VDD.n5082 VSS 0.012131f
C22631 VDD.n5083 VSS 0.012131f
C22632 VDD.n5084 VSS 0.012131f
C22633 VDD.n5085 VSS 0.012131f
C22634 VDD.n5086 VSS 0.012131f
C22635 VDD.n5087 VSS 0.012131f
C22636 VDD.n5088 VSS 0.012131f
C22637 VDD.n5089 VSS 0.012131f
C22638 VDD.n5090 VSS 0.012131f
C22639 VDD.n5091 VSS 0.012131f
C22640 VDD.n5092 VSS 0.012131f
C22641 VDD.n5093 VSS 0.012131f
C22642 VDD.n5094 VSS 0.012131f
C22643 VDD.n5095 VSS 0.012131f
C22644 VDD.n5096 VSS 0.012131f
C22645 VDD.n5097 VSS 0.012131f
C22646 VDD.n5098 VSS 0.012131f
C22647 VDD.n5099 VSS 0.012131f
C22648 VDD.n5100 VSS 0.012131f
C22649 VDD.n5101 VSS 0.012131f
C22650 VDD.n5102 VSS 0.012131f
C22651 VDD.n5103 VSS 0.012131f
C22652 VDD.n5104 VSS 0.012131f
C22653 VDD.n5105 VSS 0.012131f
C22654 VDD.n5106 VSS 0.012131f
C22655 VDD.n5107 VSS 0.012131f
C22656 VDD.n5108 VSS 0.012131f
C22657 VDD.n5109 VSS 0.012131f
C22658 VDD.n5110 VSS 0.012131f
C22659 VDD.n5111 VSS 0.012131f
C22660 VDD.n5112 VSS 0.012131f
C22661 VDD.n5113 VSS 0.012131f
C22662 VDD.n5114 VSS 0.012131f
C22663 VDD.n5115 VSS 0.012131f
C22664 VDD.n5116 VSS 0.012131f
C22665 VDD.n5117 VSS 0.012131f
C22666 VDD.n5118 VSS 0.012131f
C22667 VDD.n5119 VSS 0.012131f
C22668 VDD.n5120 VSS 0.012131f
C22669 VDD.n5121 VSS 0.012131f
C22670 VDD.n5122 VSS 0.012131f
C22671 VDD.n5123 VSS 0.012131f
C22672 VDD.n5124 VSS 0.012131f
C22673 VDD.n5125 VSS 0.012131f
C22674 VDD.n5126 VSS 0.012131f
C22675 VDD.n5127 VSS 0.012131f
C22676 VDD.n5128 VSS 0.012131f
C22677 VDD.n5129 VSS 0.012131f
C22678 VDD.n5130 VSS 0.012131f
C22679 VDD.n5131 VSS 0.012131f
C22680 VDD.n5132 VSS 0.012131f
C22681 VDD.n5133 VSS 0.012131f
C22682 VDD.n5134 VSS 0.012131f
C22683 VDD.n5135 VSS 0.012131f
C22684 VDD.n5136 VSS 0.012131f
C22685 VDD.n5137 VSS 0.012131f
C22686 VDD.n5138 VSS 0.012131f
C22687 VDD.n5139 VSS 0.012131f
C22688 VDD.n5140 VSS 0.012131f
C22689 VDD.n5141 VSS 0.012131f
C22690 VDD.n5142 VSS 0.012131f
C22691 VDD.n5143 VSS 0.012131f
C22692 VDD.n5144 VSS 0.012131f
C22693 VDD.n5145 VSS 0.012131f
C22694 VDD.n5146 VSS 0.012131f
C22695 VDD.n5147 VSS 0.012131f
C22696 VDD.n5148 VSS 0.012131f
C22697 VDD.n5149 VSS 0.012131f
C22698 VDD.n5150 VSS 0.012131f
C22699 VDD.n5151 VSS 0.012131f
C22700 VDD.n5152 VSS 0.012131f
C22701 VDD.n5153 VSS 0.012131f
C22702 VDD.n5154 VSS 0.012131f
C22703 VDD.n5155 VSS 0.012131f
C22704 VDD.n5156 VSS 0.012131f
C22705 VDD.n5157 VSS 0.012131f
C22706 VDD.n5158 VSS 0.012131f
C22707 VDD.n5159 VSS 0.012131f
C22708 VDD.n5160 VSS 0.012131f
C22709 VDD.n5161 VSS 0.012131f
C22710 VDD.n5162 VSS 0.012131f
C22711 VDD.n5163 VSS 0.012131f
C22712 VDD.n5164 VSS 0.012131f
C22713 VDD.n5165 VSS 0.012131f
C22714 VDD.n5166 VSS 0.012131f
C22715 VDD.n5167 VSS 0.012131f
C22716 VDD.n5168 VSS 0.012131f
C22717 VDD.n5169 VSS 0.012131f
C22718 VDD.n5170 VSS 0.012131f
C22719 VDD.n5171 VSS 0.012131f
C22720 VDD.n5172 VSS 0.012131f
C22721 VDD.n5173 VSS 0.012131f
C22722 VDD.n5174 VSS 0.012131f
C22723 VDD.n5175 VSS 0.012131f
C22724 VDD.n5176 VSS 0.012131f
C22725 VDD.n5177 VSS 0.012131f
C22726 VDD.n5178 VSS 0.012131f
C22727 VDD.n5179 VSS 0.012131f
C22728 VDD.n5180 VSS 0.012131f
C22729 VDD.n5181 VSS 0.012131f
C22730 VDD.n5182 VSS 0.012131f
C22731 VDD.n5183 VSS 0.012131f
C22732 VDD.n5184 VSS 0.012131f
C22733 VDD.n5185 VSS 0.012131f
C22734 VDD.n5186 VSS 0.012131f
C22735 VDD.n5187 VSS 0.012131f
C22736 VDD.n5188 VSS 0.012131f
C22737 VDD.n5189 VSS 0.012131f
C22738 VDD.n5190 VSS 0.012131f
C22739 VDD.n5191 VSS 0.012131f
C22740 VDD.n5192 VSS 0.012131f
C22741 VDD.n5193 VSS 0.012131f
C22742 VDD.n5194 VSS 0.012131f
C22743 VDD.n5195 VSS 0.012131f
C22744 VDD.n5196 VSS 0.012131f
C22745 VDD.n5197 VSS 0.012131f
C22746 VDD.n5198 VSS 0.012131f
C22747 VDD.n5199 VSS 0.012131f
C22748 VDD.n5200 VSS 0.009899f
C22749 VDD.n5201 VSS 0.015408f
C22750 VDD.n5202 VSS 0.020419f
C22751 VDD.n5203 VSS 0.006065f
C22752 VDD.n5204 VSS 0.012131f
C22753 VDD.n5205 VSS 0.006065f
C22754 VDD.n5206 VSS 0.012131f
C22755 VDD.n5207 VSS 0.012131f
C22756 VDD.n5208 VSS 0.012131f
C22757 VDD.n5209 VSS 0.012131f
C22758 VDD.n5210 VSS 0.012131f
C22759 VDD.n5211 VSS 0.012131f
C22760 VDD.n5212 VSS 0.012131f
C22761 VDD.n5213 VSS 0.012131f
C22762 VDD.n5214 VSS 0.012131f
C22763 VDD.n5215 VSS 0.012131f
C22764 VDD.n5216 VSS 0.012131f
C22765 VDD.n5217 VSS 0.006065f
C22766 VDD.n5218 VSS 0.166738f
C22767 VDD.n5219 VSS 0.012131f
C22768 VDD.n5220 VSS 0.698912f
C22769 VDD.t2873 VSS 0.034186f
C22770 VDD.t708 VSS 0.034186f
C22771 VDD.t707 VSS 0.066856f
C22772 VDD.t4425 VSS 0.034186f
C22773 VDD.t2448 VSS 0.034186f
C22774 VDD.t2447 VSS 0.066856f
C22775 VDD.t2000 VSS 0.066856f
C22776 VDD.t4091 VSS 0.034186f
C22777 VDD.t2001 VSS 0.034186f
C22778 VDD.n5221 VSS 0.283088f
C22779 VDD.t993 VSS 0.034186f
C22780 VDD.t3111 VSS 0.034186f
C22781 VDD.t3110 VSS 0.066856f
C22782 VDD.t2781 VSS 0.066856f
C22783 VDD.t4741 VSS 0.034186f
C22784 VDD.t2782 VSS 0.034186f
C22785 VDD.t4330 VSS 0.066856f
C22786 VDD.t2294 VSS 0.034186f
C22787 VDD.t4331 VSS 0.034186f
C22788 VDD.t2594 VSS 0.025104f
C22789 VDD.t2593 VSS 0.066856f
C22790 VDD.t4572 VSS 0.066856f
C22791 VDD.n5222 VSS 0.256005f
C22792 VDD.t3692 VSS 0.016021f
C22793 VDD.n5223 VSS 0.016021f
C22794 VDD.t1576 VSS 0.066856f
C22795 VDD.t1577 VSS 0.016021f
C22796 VDD.n5224 VSS 0.016021f
C22797 VDD.t4364 VSS 0.066856f
C22798 VDD.t2391 VSS 0.066856f
C22799 VDD.n5225 VSS 0.256005f
C22800 VDD.t1048 VSS 0.025104f
C22801 VDD.t4365 VSS 0.016021f
C22802 VDD.n5226 VSS 0.016021f
C22803 VDD.t3162 VSS 0.066856f
C22804 VDD.t3163 VSS 0.025104f
C22805 VDD.t3623 VSS 0.025104f
C22806 VDD.t3622 VSS 0.066856f
C22807 VDD.t1533 VSS 0.066856f
C22808 VDD.n5227 VSS 0.256005f
C22809 VDD.t4341 VSS 0.016021f
C22810 VDD.n5228 VSS 0.016021f
C22811 VDD.t2280 VSS 0.066856f
C22812 VDD.t2281 VSS 0.016021f
C22813 VDD.n5229 VSS 0.016021f
C22814 VDD.t4102 VSS 0.066856f
C22815 VDD.t2041 VSS 0.066856f
C22816 VDD.n5230 VSS 0.256005f
C22817 VDD.t4103 VSS 0.025104f
C22818 VDD.t4579 VSS 0.025104f
C22819 VDD.t4578 VSS 0.066856f
C22820 VDD.t2637 VSS 0.066856f
C22821 VDD.n5231 VSS 0.256005f
C22822 VDD.t811 VSS 0.016021f
C22823 VDD.n5232 VSS 0.016021f
C22824 VDD.t2956 VSS 0.066856f
C22825 VDD.t2957 VSS 0.016021f
C22826 VDD.n5233 VSS 0.016021f
C22827 VDD.t1948 VSS 0.066856f
C22828 VDD.t4058 VSS 0.066856f
C22829 VDD.n5234 VSS 0.256005f
C22830 VDD.t2764 VSS 0.025104f
C22831 VDD.t1949 VSS 0.016021f
C22832 VDD.t4727 VSS 0.025104f
C22833 VDD.n5235 VSS 0.016021f
C22834 VDD.t4726 VSS 0.066856f
C22835 VDD.t2763 VSS 0.066856f
C22836 VDD.n5236 VSS 0.256005f
C22837 VDD.n5237 VSS 0.208141f
C22838 VDD.n5238 VSS 0.016021f
C22839 VDD.t4059 VSS 0.016021f
C22840 VDD.n5239 VSS 0.016021f
C22841 VDD.n5240 VSS 0.208141f
C22842 VDD.t810 VSS 0.066856f
C22843 VDD.n5241 VSS 0.256005f
C22844 VDD.n5242 VSS 0.208141f
C22845 VDD.n5243 VSS 0.016021f
C22846 VDD.t2638 VSS 0.025104f
C22847 VDD.n5244 VSS 0.218415f
C22848 VDD.n5245 VSS 0.218415f
C22849 VDD.t2042 VSS 0.025104f
C22850 VDD.n5246 VSS 0.016021f
C22851 VDD.n5247 VSS 0.208141f
C22852 VDD.t4340 VSS 0.066856f
C22853 VDD.n5248 VSS 0.163661f
C22854 VDD.n5249 VSS 0.10407f
C22855 VDD.n5250 VSS 0.196415f
C22856 VDD.n5251 VSS 0.016021f
C22857 VDD.t1534 VSS 0.025104f
C22858 VDD.n5252 VSS 0.218415f
C22859 VDD.n5253 VSS 0.218415f
C22860 VDD.t1047 VSS 0.066856f
C22861 VDD.n5254 VSS 0.256005f
C22862 VDD.n5255 VSS 0.208141f
C22863 VDD.n5256 VSS 0.016021f
C22864 VDD.t2392 VSS 0.016021f
C22865 VDD.n5257 VSS 0.016021f
C22866 VDD.n5258 VSS 0.208141f
C22867 VDD.t3691 VSS 0.066856f
C22868 VDD.n5259 VSS 0.256005f
C22869 VDD.n5260 VSS 0.208141f
C22870 VDD.n5261 VSS 0.016021f
C22871 VDD.t4573 VSS 0.025104f
C22872 VDD.n5262 VSS 0.225377f
C22873 VDD.n5263 VSS 0.225377f
C22874 VDD.t4309 VSS 0.034186f
C22875 VDD.t2260 VSS 0.034186f
C22876 VDD.t2259 VSS 0.066856f
C22877 VDD.t2017 VSS 0.034186f
C22878 VDD.t4113 VSS 0.034186f
C22879 VDD.t4112 VSS 0.066856f
C22880 VDD.t3731 VSS 0.066856f
C22881 VDD.t1640 VSS 0.034186f
C22882 VDD.t3732 VSS 0.034186f
C22883 VDD.n5264 VSS 0.283088f
C22884 VDD.t3929 VSS 0.034186f
C22885 VDD.t1818 VSS 0.034186f
C22886 VDD.t1817 VSS 0.066856f
C22887 VDD.t1451 VSS 0.066856f
C22888 VDD.t3561 VSS 0.034186f
C22889 VDD.t1452 VSS 0.034186f
C22890 VDD.t3188 VSS 0.066856f
C22891 VDD.t1062 VSS 0.034186f
C22892 VDD.t3189 VSS 0.034186f
C22893 VDD.n5265 VSS 0.385214f
C22894 VDD.t1076 VSS 0.034186f
C22895 VDD.t3207 VSS 0.034186f
C22896 VDD.t3206 VSS 0.066856f
C22897 VDD.t2808 VSS 0.034186f
C22898 VDD.t618 VSS 0.034186f
C22899 VDD.t616 VSS 0.066856f
C22900 VDD.t4410 VSS 0.066856f
C22901 VDD.t2438 VSS 0.034186f
C22902 VDD.t4411 VSS 0.034186f
C22903 VDD.n5266 VSS 0.283088f
C22904 VDD.t2691 VSS 0.034186f
C22905 VDD.t4679 VSS 0.034186f
C22906 VDD.n5267 VSS 0.715132f
C22907 VDD.n5268 VSS 12.0304f
C22908 VDD.t2169 VSS 0.034186f
C22909 VDD.t4243 VSS 0.034186f
C22910 VDD.n5269 VSS 0.652605f
C22911 VDD.n5270 VSS 0.283088f
C22912 VDD.t2220 VSS 0.034186f
C22913 VDD.t4275 VSS 0.034186f
C22914 VDD.t4274 VSS 0.066856f
C22915 VDD.t3920 VSS 0.066856f
C22916 VDD.t1808 VSS 0.034186f
C22917 VDD.t3921 VSS 0.034186f
C22918 VDD.t1594 VSS 0.066856f
C22919 VDD.t3686 VSS 0.034186f
C22920 VDD.t1595 VSS 0.034186f
C22921 VDD.t2460 VSS 0.066856f
C22922 VDD.n5271 VSS 0.129831f
C22923 VDD.t3759 VSS 0.016021f
C22924 VDD.t4648 VSS 0.066856f
C22925 VDD.n5272 VSS 0.129831f
C22926 VDD.t2285 VSS 0.025104f
C22927 VDD.t1701 VSS 0.066856f
C22928 VDD.n5273 VSS 0.129831f
C22929 VDD.t4053 VSS 0.016021f
C22930 VDD.n5274 VSS 0.099933f
C22931 VDD.n5275 VSS 0.280759f
C22932 VDD.t403 VSS 9.213929f
C22933 VDD.n5276 VSS 0.283109f
C22934 VDD.n5277 VSS 0.283109f
C22935 VDD.n5278 VSS 0.283109f
C22936 VDD.t617 VSS 9.19382f
C22937 VDD.t397 VSS 9.81076f
C22938 VDD.t410 VSS 7.61793f
C22939 VDD.t407 VSS 7.61793f
C22940 VDD.t399 VSS 9.428519f
C22941 VDD.t395 VSS 9.428519f
C22942 VDD.t408 VSS 4.02355f
C22943 VDD.n5279 VSS 0.279865f
C22944 VDD.n5280 VSS 0.279865f
C22945 VDD.n5281 VSS 0.279865f
C22946 VDD.n5282 VSS 0.280759f
C22947 VDD.n5283 VSS 0.096993f
C22948 VDD.t852 VSS 0.066856f
C22949 VDD.n5284 VSS 0.126716f
C22950 VDD.t3211 VSS 0.016021f
C22951 VDD.t1320 VSS 0.066856f
C22952 VDD.n5285 VSS 0.126716f
C22953 VDD.t3769 VSS 0.016021f
C22954 VDD.t2948 VSS 0.066856f
C22955 VDD.n5286 VSS 0.126716f
C22956 VDD.t1454 VSS 0.025104f
C22957 VDD.t1453 VSS 0.066856f
C22958 VDD.n5287 VSS 0.057673f
C22959 VDD.n5288 VSS 0.05157f
C22960 VDD.n5289 VSS 0.32091f
C22961 VDD.t4882 VSS 0.008011f
C22962 VDD.t4941 VSS 0.008011f
C22963 VDD.n5290 VSS 0.04401f
C22964 VDD.t4881 VSS 0.008011f
C22965 VDD.t4833 VSS 0.008011f
C22966 VDD.n5291 VSS 0.029389f
C22967 VDD.n5292 VSS 0.144542f
C22968 VDD.t4892 VSS 0.008011f
C22969 VDD.t4974 VSS 0.008011f
C22970 VDD.n5293 VSS 0.029389f
C22971 VDD.n5294 VSS 0.102512f
C22972 VDD.t4914 VSS 0.008011f
C22973 VDD.t4898 VSS 0.008011f
C22974 VDD.n5295 VSS 0.029389f
C22975 VDD.n5296 VSS 0.041173f
C22976 VDD.n5297 VSS 0.041824f
C22977 VDD.t1110 VSS 0.066856f
C22978 VDD.n5298 VSS 0.057673f
C22979 VDD.n5299 VSS 0.437712f
C22980 VDD.t1420 VSS 0.016021f
C22981 VDD.t2900 VSS 0.066856f
C22982 VDD.n5300 VSS 0.126716f
C22983 VDD.t1006 VSS 0.025104f
C22984 VDD.t4596 VSS 0.066856f
C22985 VDD.n5301 VSS 0.126716f
C22986 VDD.t2861 VSS 0.016021f
C22987 VDD.n5302 VSS 0.096993f
C22988 VDD.n5303 VSS 0.280759f
C22989 VDD.n5304 VSS 0.283088f
C22990 VDD.t409 VSS 9.213929f
C22991 VDD.n5305 VSS 0.283109f
C22992 VDD.n5306 VSS 0.283109f
C22993 VDD.n5307 VSS 0.283109f
C22994 VDD.n5308 VSS 0.283109f
C22995 VDD.t412 VSS 4.02355f
C22996 VDD.n5309 VSS 0.279865f
C22997 VDD.n5310 VSS 0.279865f
C22998 VDD.n5311 VSS 0.280759f
C22999 VDD.n5312 VSS 0.283088f
C23000 VDD.n5313 VSS 0.196415f
C23001 VDD.t4296 VSS 0.066856f
C23002 VDD.n5314 VSS 0.016021f
C23003 VDD.t1979 VSS 0.066856f
C23004 VDD.t4094 VSS 0.066856f
C23005 VDD.n5315 VSS 0.256005f
C23006 VDD.t2273 VSS 0.016021f
C23007 VDD.t1980 VSS 0.025104f
C23008 VDD.t2592 VSS 0.025104f
C23009 VDD.t2591 VSS 0.066856f
C23010 VDD.t4570 VSS 0.066856f
C23011 VDD.n5316 VSS 0.256005f
C23012 VDD.t2343 VSS 0.016021f
C23013 VDD.n5317 VSS 0.016021f
C23014 VDD.t4342 VSS 0.066856f
C23015 VDD.t4343 VSS 0.016021f
C23016 VDD.n5318 VSS 0.016021f
C23017 VDD.t3044 VSS 0.066856f
C23018 VDD.t930 VSS 0.066856f
C23019 VDD.n5319 VSS 0.256005f
C23020 VDD.t4721 VSS 0.025104f
C23021 VDD.t3045 VSS 0.016021f
C23022 VDD.n5320 VSS 0.016021f
C23023 VDD.t2718 VSS 0.066856f
C23024 VDD.t2719 VSS 0.025104f
C23025 VDD.t2204 VSS 0.025104f
C23026 VDD.t2203 VSS 0.066856f
C23027 VDD.t4278 VSS 0.066856f
C23028 VDD.n5321 VSS 0.256005f
C23029 VDD.t1962 VSS 0.016021f
C23030 VDD.n5322 VSS 0.016021f
C23031 VDD.t4040 VSS 0.066856f
C23032 VDD.t4041 VSS 0.016021f
C23033 VDD.n5323 VSS 0.016021f
C23034 VDD.t2737 VSS 0.066856f
C23035 VDD.t4732 VSS 0.066856f
C23036 VDD.n5324 VSS 0.256005f
C23037 VDD.t717 VSS 0.025104f
C23038 VDD.t2738 VSS 0.016021f
C23039 VDD.n5325 VSS 0.016021f
C23040 VDD.t2862 VSS 0.066856f
C23041 VDD.t2863 VSS 0.025104f
C23042 VDD.t1874 VSS 0.025104f
C23043 VDD.t1873 VSS 0.066856f
C23044 VDD.t3998 VSS 0.066856f
C23045 VDD.n5326 VSS 0.256005f
C23046 VDD.t2697 VSS 0.016021f
C23047 VDD.n5327 VSS 0.016021f
C23048 VDD.t4662 VSS 0.066856f
C23049 VDD.t4663 VSS 0.016021f
C23050 VDD.n5328 VSS 0.016021f
C23051 VDD.t2433 VSS 0.066856f
C23052 VDD.t4442 VSS 0.066856f
C23053 VDD.n5329 VSS 0.256005f
C23054 VDD.t2434 VSS 0.025104f
C23055 VDD.t2963 VSS 0.025104f
C23056 VDD.t2962 VSS 0.066856f
C23057 VDD.t823 VSS 0.066856f
C23058 VDD.n5330 VSS 0.256005f
C23059 VDD.t3279 VSS 0.016021f
C23060 VDD.n5331 VSS 0.016021f
C23061 VDD.t1125 VSS 0.066856f
C23062 VDD.t1126 VSS 0.016021f
C23063 VDD.n5332 VSS 0.016021f
C23064 VDD.t4370 VSS 0.066856f
C23065 VDD.t2395 VSS 0.066856f
C23066 VDD.n5333 VSS 0.256005f
C23067 VDD.t963 VSS 0.025104f
C23068 VDD.t4371 VSS 0.016021f
C23069 VDD.t3079 VSS 0.025104f
C23070 VDD.n5334 VSS 0.016021f
C23071 VDD.t3078 VSS 0.066856f
C23072 VDD.t962 VSS 0.066856f
C23073 VDD.n5335 VSS 0.256005f
C23074 VDD.n5336 VSS 0.208141f
C23075 VDD.n5337 VSS 0.016021f
C23076 VDD.t2396 VSS 0.016021f
C23077 VDD.n5338 VSS 0.016021f
C23078 VDD.n5339 VSS 0.208141f
C23079 VDD.t3278 VSS 0.066856f
C23080 VDD.n5340 VSS 0.256005f
C23081 VDD.n5341 VSS 0.208141f
C23082 VDD.n5342 VSS 0.016021f
C23083 VDD.t824 VSS 0.025104f
C23084 VDD.n5343 VSS 0.218415f
C23085 VDD.n5344 VSS 0.218415f
C23086 VDD.t4443 VSS 0.025104f
C23087 VDD.n5345 VSS 0.016021f
C23088 VDD.n5346 VSS 0.208141f
C23089 VDD.t2696 VSS 0.066856f
C23090 VDD.n5347 VSS 0.163661f
C23091 VDD.n5348 VSS 0.10407f
C23092 VDD.n5349 VSS 0.196415f
C23093 VDD.n5350 VSS 0.016021f
C23094 VDD.t3999 VSS 0.025104f
C23095 VDD.n5351 VSS 0.218415f
C23096 VDD.n5352 VSS 0.218415f
C23097 VDD.t716 VSS 0.066856f
C23098 VDD.n5353 VSS 0.256005f
C23099 VDD.n5354 VSS 0.208141f
C23100 VDD.n5355 VSS 0.016021f
C23101 VDD.t4733 VSS 0.016021f
C23102 VDD.n5356 VSS 0.016021f
C23103 VDD.n5357 VSS 0.208141f
C23104 VDD.t1961 VSS 0.066856f
C23105 VDD.n5358 VSS 0.256005f
C23106 VDD.n5359 VSS 0.208141f
C23107 VDD.n5360 VSS 0.016021f
C23108 VDD.t4279 VSS 0.025104f
C23109 VDD.n5361 VSS 0.225377f
C23110 VDD.t2559 VSS 0.034186f
C23111 VDD.t3473 VSS 0.034186f
C23112 VDD.n5362 VSS 0.172271f
C23113 VDD.t3472 VSS 0.066856f
C23114 VDD.t2558 VSS 0.066856f
C23115 VDD.n5363 VSS 0.58882f
C23116 VDD.t4139 VSS 0.034186f
C23117 VDD.t977 VSS 0.034186f
C23118 VDD.n5364 VSS 0.571765f
C23119 VDD.t976 VSS 0.066856f
C23120 VDD.t4138 VSS 0.066856f
C23121 VDD.n5365 VSS 0.333277f
C23122 VDD.t4734 VSS 0.066856f
C23123 VDD.t3764 VSS 0.066856f
C23124 VDD.n5366 VSS 0.333277f
C23125 VDD.t3765 VSS 0.034186f
C23126 VDD.t4735 VSS 0.034186f
C23127 VDD.n5367 VSS 0.402094f
C23128 VDD.n5368 VSS 0.532659f
C23129 VDD.t621 VSS 0.034186f
C23130 VDD.t1611 VSS 0.034186f
C23131 VDD.n5369 VSS 0.43943f
C23132 VDD.t1610 VSS 0.066856f
C23133 VDD.t619 VSS 0.066856f
C23134 VDD.n5370 VSS 0.333277f
C23135 VDD.t1251 VSS 0.066856f
C23136 VDD.t4422 VSS 0.066856f
C23137 VDD.n5371 VSS 0.333277f
C23138 VDD.t4423 VSS 0.034186f
C23139 VDD.t1252 VSS 0.034186f
C23140 VDD.n5372 VSS 0.571765f
C23141 VDD.t3010 VSS 0.066856f
C23142 VDD.t1923 VSS 0.066856f
C23143 VDD.n5373 VSS 0.58882f
C23144 VDD.t1924 VSS 0.034186f
C23145 VDD.t3011 VSS 0.034186f
C23146 VDD.n5374 VSS 0.33406f
C23147 VDD.t4007 VSS 0.034186f
C23148 VDD.t843 VSS 0.034186f
C23149 VDD.t841 VSS 0.066856f
C23150 VDD.t1674 VSS 0.034186f
C23151 VDD.t2774 VSS 0.034186f
C23152 VDD.t2773 VSS 0.066856f
C23153 VDD.t2397 VSS 0.066856f
C23154 VDD.t1309 VSS 0.034186f
C23155 VDD.t2398 VSS 0.034186f
C23156 VDD.t3598 VSS 0.034186f
C23157 VDD.t4547 VSS 0.034186f
C23158 VDD.n5375 VSS 0.43943f
C23159 VDD.t400 VSS 9.428519f
C23160 VDD.t396 VSS 9.428519f
C23161 VDD.t411 VSS 7.61793f
C23162 VDD.t398 VSS 7.61793f
C23163 VDD.t394 VSS 9.81076f
C23164 VDD.t842 VSS 9.19382f
C23165 VDD.n5376 VSS 4.15767f
C23166 VDD.t402 VSS 9.428519f
C23167 VDD.t391 VSS 7.61793f
C23168 VDD.t414 VSS 7.61793f
C23169 VDD.t390 VSS 9.81076f
C23170 VDD.t620 VSS 9.19382f
C23171 VDD.t2051 VSS 0.034186f
C23172 VDD.t3091 VSS 0.034186f
C23173 VDD.n5377 VSS 0.402094f
C23174 VDD.n5378 VSS 0.283088f
C23175 VDD.t2345 VSS 0.034186f
C23176 VDD.t3305 VSS 0.034186f
C23177 VDD.t3304 VSS 0.066856f
C23178 VDD.t3002 VSS 0.066856f
C23179 VDD.t1911 VSS 0.034186f
C23180 VDD.t3003 VSS 0.034186f
C23181 VDD.t2708 VSS 0.066856f
C23182 VDD.t1624 VSS 0.034186f
C23183 VDD.t2709 VSS 0.034186f
C23184 VDD.t2973 VSS 0.025104f
C23185 VDD.t2972 VSS 0.066856f
C23186 VDD.t3994 VSS 0.066856f
C23187 VDD.n5379 VSS 0.256005f
C23188 VDD.t1653 VSS 0.016021f
C23189 VDD.n5380 VSS 0.016021f
C23190 VDD.t4714 VSS 0.066856f
C23191 VDD.t4715 VSS 0.016021f
C23192 VDD.n5381 VSS 0.016021f
C23193 VDD.t3359 VSS 0.066856f
C23194 VDD.t4438 VSS 0.066856f
C23195 VDD.n5382 VSS 0.256005f
C23196 VDD.t4543 VSS 0.025104f
C23197 VDD.t3360 VSS 0.016021f
C23198 VDD.n5383 VSS 0.016021f
C23199 VDD.t3500 VSS 0.066856f
C23200 VDD.t3501 VSS 0.025104f
C23201 VDD.t2680 VSS 0.025104f
C23202 VDD.t2679 VSS 0.066856f
C23203 VDD.t3689 VSS 0.066856f
C23204 VDD.n5384 VSS 0.256005f
C23205 VDD.t2390 VSS 0.016021f
C23206 VDD.n5385 VSS 0.016021f
C23207 VDD.t1195 VSS 0.066856f
C23208 VDD.t1196 VSS 0.016021f
C23209 VDD.n5386 VSS 0.016021f
C23210 VDD.t3122 VSS 0.066856f
C23211 VDD.t4176 VSS 0.066856f
C23212 VDD.n5387 VSS 0.256005f
C23213 VDD.t3123 VSS 0.025104f
C23214 VDD.t3584 VSS 0.025104f
C23215 VDD.t3583 VSS 0.066856f
C23216 VDD.t4668 VSS 0.066856f
C23217 VDD.n5388 VSS 0.256005f
C23218 VDD.t3019 VSS 0.016021f
C23219 VDD.n5389 VSS 0.016021f
C23220 VDD.t1811 VSS 0.066856f
C23221 VDD.t1812 VSS 0.016021f
C23222 VDD.n5390 VSS 0.016021f
C23223 VDD.t951 VSS 0.066856f
C23224 VDD.t2039 VSS 0.066856f
C23225 VDD.n5391 VSS 0.256005f
C23226 VDD.t632 VSS 0.025104f
C23227 VDD.t952 VSS 0.016021f
C23228 VDD.n5392 VSS 0.016021f
C23229 VDD.t3701 VSS 0.066856f
C23230 VDD.t3702 VSS 0.025104f
C23231 VDD.t3263 VSS 0.025104f
C23232 VDD.t3262 VSS 0.066856f
C23233 VDD.t4302 VSS 0.066856f
C23234 VDD.n5393 VSS 0.256005f
C23235 VDD.t3418 VSS 0.016021f
C23236 VDD.n5394 VSS 0.016021f
C23237 VDD.t2372 VSS 0.066856f
C23238 VDD.t2373 VSS 0.016021f
C23239 VDD.n5395 VSS 0.016021f
C23240 VDD.t949 VSS 0.066856f
C23241 VDD.t2031 VSS 0.066856f
C23242 VDD.n5396 VSS 0.256005f
C23243 VDD.t769 VSS 0.025104f
C23244 VDD.t950 VSS 0.016021f
C23245 VDD.n5397 VSS 0.016021f
C23246 VDD.t3808 VSS 0.066856f
C23247 VDD.t3809 VSS 0.025104f
C23248 VDD.t4319 VSS 0.025104f
C23249 VDD.t4318 VSS 0.066856f
C23250 VDD.t1247 VSS 0.066856f
C23251 VDD.n5398 VSS 0.256005f
C23252 VDD.t4055 VSS 0.016021f
C23253 VDD.n5399 VSS 0.016021f
C23254 VDD.t3026 VSS 0.066856f
C23255 VDD.t3027 VSS 0.016021f
C23256 VDD.n5400 VSS 0.016021f
C23257 VDD.t604 VSS 0.066856f
C23258 VDD.t1703 VSS 0.066856f
C23259 VDD.n5401 VSS 0.256005f
C23260 VDD.t605 VSS 0.025104f
C23261 VDD.t1137 VSS 0.025104f
C23262 VDD.t1136 VSS 0.066856f
C23263 VDD.t2286 VSS 0.066856f
C23264 VDD.n5402 VSS 0.256005f
C23265 VDD.t4651 VSS 0.016021f
C23266 VDD.n5403 VSS 0.016021f
C23267 VDD.t3575 VSS 0.066856f
C23268 VDD.t3576 VSS 0.016021f
C23269 VDD.n5404 VSS 0.016021f
C23270 VDD.t2751 VSS 0.066856f
C23271 VDD.t3762 VSS 0.066856f
C23272 VDD.n5405 VSS 0.256005f
C23273 VDD.t2463 VSS 0.025104f
C23274 VDD.t2752 VSS 0.016021f
C23275 VDD.t1261 VSS 0.025104f
C23276 VDD.n5406 VSS 0.016021f
C23277 VDD.t1260 VSS 0.066856f
C23278 VDD.t2462 VSS 0.066856f
C23279 VDD.n5407 VSS 0.256005f
C23280 VDD.n5408 VSS 0.208141f
C23281 VDD.n5409 VSS 0.016021f
C23282 VDD.t3763 VSS 0.016021f
C23283 VDD.n5410 VSS 0.016021f
C23284 VDD.n5411 VSS 0.208141f
C23285 VDD.t4650 VSS 0.066856f
C23286 VDD.n5412 VSS 0.256005f
C23287 VDD.n5413 VSS 0.208141f
C23288 VDD.n5414 VSS 0.016021f
C23289 VDD.t2287 VSS 0.025104f
C23290 VDD.n5415 VSS 0.218415f
C23291 VDD.n5416 VSS 0.218415f
C23292 VDD.t1704 VSS 0.025104f
C23293 VDD.n5417 VSS 0.016021f
C23294 VDD.n5418 VSS 0.208141f
C23295 VDD.t4054 VSS 0.066856f
C23296 VDD.n5419 VSS 0.163661f
C23297 VDD.n5420 VSS 0.10407f
C23298 VDD.n5421 VSS 0.196415f
C23299 VDD.n5422 VSS 0.016021f
C23300 VDD.t1248 VSS 0.025104f
C23301 VDD.n5423 VSS 0.218415f
C23302 VDD.n5424 VSS 0.218415f
C23303 VDD.t768 VSS 0.066856f
C23304 VDD.n5425 VSS 0.256005f
C23305 VDD.n5426 VSS 0.208141f
C23306 VDD.n5427 VSS 0.016021f
C23307 VDD.t2032 VSS 0.016021f
C23308 VDD.n5428 VSS 0.016021f
C23309 VDD.n5429 VSS 0.208141f
C23310 VDD.t3417 VSS 0.066856f
C23311 VDD.n5430 VSS 0.256005f
C23312 VDD.n5431 VSS 0.208141f
C23313 VDD.n5432 VSS 0.016021f
C23314 VDD.t4303 VSS 0.025104f
C23315 VDD.n5433 VSS 0.225377f
C23316 VDD.t4678 VSS 0.066856f
C23317 VDD.t2690 VSS 0.066856f
C23318 VDD.n5434 VSS 0.525848f
C23319 VDD.t4316 VSS 0.066856f
C23320 VDD.t2276 VSS 0.066856f
C23321 VDD.n5435 VSS 0.525848f
C23322 VDD.t2277 VSS 0.034186f
C23323 VDD.t4317 VSS 0.034186f
C23324 VDD.n5436 VSS 0.936755f
C23325 VDD.t4050 VSS 0.066856f
C23326 VDD.t1954 VSS 0.066856f
C23327 VDD.n5437 VSS 0.95381f
C23328 VDD.t1955 VSS 0.034186f
C23329 VDD.t4051 VSS 0.034186f
C23330 VDD.n5438 VSS 0.538667f
C23331 VDD.t890 VSS 0.034186f
C23332 VDD.t3023 VSS 0.034186f
C23333 VDD.t3022 VSS 0.066856f
C23334 VDD.t2606 VSS 0.034186f
C23335 VDD.t4559 VSS 0.034186f
C23336 VDD.t4558 VSS 0.066856f
C23337 VDD.t4242 VSS 0.066856f
C23338 VDD.t2168 VSS 0.066856f
C23339 VDD.n5439 VSS 0.525848f
C23340 VDD.t2605 VSS 0.066856f
C23341 VDD.n5440 VSS 0.525848f
C23342 VDD.n5441 VSS 0.936755f
C23343 VDD.t888 VSS 0.066856f
C23344 VDD.n5442 VSS 0.95381f
C23345 VDD.n5443 VSS 0.537972f
C23346 VDD.n5444 VSS 0.812758f
C23347 VDD.n5445 VSS 0.225377f
C23348 VDD.t631 VSS 0.066856f
C23349 VDD.n5446 VSS 0.256005f
C23350 VDD.n5447 VSS 0.208141f
C23351 VDD.n5448 VSS 0.016021f
C23352 VDD.t2040 VSS 0.016021f
C23353 VDD.n5449 VSS 0.016021f
C23354 VDD.n5450 VSS 0.208141f
C23355 VDD.t3018 VSS 0.066856f
C23356 VDD.n5451 VSS 0.256005f
C23357 VDD.n5452 VSS 0.208141f
C23358 VDD.n5453 VSS 0.016021f
C23359 VDD.t4669 VSS 0.025104f
C23360 VDD.n5454 VSS 0.218415f
C23361 VDD.n5455 VSS 0.218415f
C23362 VDD.t4177 VSS 0.025104f
C23363 VDD.n5456 VSS 0.016021f
C23364 VDD.n5457 VSS 0.208141f
C23365 VDD.t2389 VSS 0.066856f
C23366 VDD.n5458 VSS 0.163661f
C23367 VDD.n5459 VSS 0.10407f
C23368 VDD.n5460 VSS 0.196415f
C23369 VDD.n5461 VSS 0.016021f
C23370 VDD.t3690 VSS 0.025104f
C23371 VDD.n5462 VSS 0.218415f
C23372 VDD.n5463 VSS 0.218415f
C23373 VDD.t4542 VSS 0.066856f
C23374 VDD.n5464 VSS 0.256005f
C23375 VDD.n5465 VSS 0.208141f
C23376 VDD.n5466 VSS 0.016021f
C23377 VDD.t4439 VSS 0.016021f
C23378 VDD.n5467 VSS 0.016021f
C23379 VDD.n5468 VSS 0.208141f
C23380 VDD.t1652 VSS 0.066856f
C23381 VDD.n5469 VSS 0.256005f
C23382 VDD.n5470 VSS 0.208141f
C23383 VDD.n5471 VSS 0.016021f
C23384 VDD.t3995 VSS 0.025104f
C23385 VDD.n5472 VSS 0.225377f
C23386 VDD.t4691 VSS 0.034186f
C23387 VDD.t1502 VSS 0.034186f
C23388 VDD.n5473 VSS 0.333645f
C23389 VDD.t3338 VSS 0.066856f
C23390 VDD.t4418 VSS 0.066856f
C23391 VDD.n5474 VSS 0.256005f
C23392 VDD.t3339 VSS 0.025104f
C23393 VDD.t570 VSS 0.016021f
C23394 VDD.t3660 VSS 0.066856f
C23395 VDD.t569 VSS 0.066856f
C23396 VDD.n5475 VSS 0.256005f
C23397 VDD.t918 VSS 0.016021f
C23398 VDD.t917 VSS 0.066856f
C23399 VDD.t1987 VSS 0.066856f
C23400 VDD.n5476 VSS 0.256005f
C23401 VDD.t4301 VSS 0.025104f
C23402 VDD.t3264 VSS 0.066856f
C23403 VDD.t4300 VSS 0.066856f
C23404 VDD.n5477 VSS 0.256005f
C23405 VDD.t2787 VSS 0.066856f
C23406 VDD.t3788 VSS 0.066856f
C23407 VDD.n5478 VSS 0.256005f
C23408 VDD.t2788 VSS 0.025104f
C23409 VDD.t1936 VSS 0.016021f
C23410 VDD.t875 VSS 0.066856f
C23411 VDD.t1935 VSS 0.066856f
C23412 VDD.n5479 VSS 0.163661f
C23413 VDD.t1170 VSS 0.025104f
C23414 VDD.t1169 VSS 0.066856f
C23415 VDD.t2336 VSS 0.066856f
C23416 VDD.n5480 VSS 0.256005f
C23417 VDD.n5481 VSS 0.10407f
C23418 VDD.t2088 VSS 0.066856f
C23419 VDD.t3230 VSS 0.066856f
C23420 VDD.n5482 VSS 0.256005f
C23421 VDD.t2089 VSS 0.025104f
C23422 VDD.t4089 VSS 0.016021f
C23423 VDD.t3052 VSS 0.066856f
C23424 VDD.t4088 VSS 0.066856f
C23425 VDD.n5483 VSS 0.256005f
C23426 VDD.t4351 VSS 0.016021f
C23427 VDD.t4350 VSS 0.066856f
C23428 VDD.t1274 VSS 0.066856f
C23429 VDD.n5484 VSS 0.256005f
C23430 VDD.t4097 VSS 0.025104f
C23431 VDD.t3056 VSS 0.066856f
C23432 VDD.t4096 VSS 0.066856f
C23433 VDD.n5485 VSS 0.256005f
C23434 VDD.t3310 VSS 0.066856f
C23435 VDD.t4372 VSS 0.066856f
C23436 VDD.n5486 VSS 0.234752f
C23437 VDD.t3311 VSS 0.034186f
C23438 VDD.n5487 VSS 0.610844f
C23439 VDD.n5488 VSS 1.75925f
C23440 VDD.n5489 VSS 0.009688f
C23441 VDD.t3547 VSS 0.028519f
C23442 VDD.t1201 VSS 0.028519f
C23443 VDD.n5491 VSS 0.009191f
C23444 VDD.t3443 VSS 0.028519f
C23445 VDD.t3557 VSS 0.028519f
C23446 VDD.n5492 VSS 0.009191f
C23447 VDD.n5493 VSS 0.413155f
C23448 VDD.t3546 VSS 0.066856f
C23449 VDD.t3442 VSS 0.066856f
C23450 VDD.t3556 VSS 0.066856f
C23451 VDD.t1200 VSS 0.066856f
C23452 VDD.n5494 VSS 0.690489f
C23453 VDD.t3224 VSS 0.066856f
C23454 VDD.t3112 VSS 0.066856f
C23455 VDD.t3240 VSS 0.066856f
C23456 VDD.t877 VSS 0.066856f
C23457 VDD.n5495 VSS 0.690489f
C23458 VDD.t3225 VSS 0.028519f
C23459 VDD.t879 VSS 0.028519f
C23460 VDD.n5496 VSS 0.009191f
C23461 VDD.t3113 VSS 0.028519f
C23462 VDD.t3241 VSS 0.028519f
C23463 VDD.n5497 VSS 0.009191f
C23464 VDD.n5498 VSS 0.644755f
C23465 VDD.t3884 VSS 0.066856f
C23466 VDD.t3403 VSS 0.066856f
C23467 VDD.t2115 VSS 0.066856f
C23468 VDD.t4710 VSS 0.066856f
C23469 VDD.n5499 VSS 0.709674f
C23470 VDD.t3885 VSS 0.028519f
C23471 VDD.t4711 VSS 0.028519f
C23472 VDD.n5500 VSS 0.009191f
C23473 VDD.t3404 VSS 0.028519f
C23474 VDD.t2116 VSS 0.028519f
C23475 VDD.n5501 VSS 0.009191f
C23476 VDD.n5502 VSS 0.28091f
C23477 VDD.n5503 VSS 0.074002f
C23478 VDD.t1380 VSS 0.066856f
C23479 VDD.n5504 VSS 0.14405f
C23480 VDD.t2262 VSS 0.025104f
C23481 VDD.n5505 VSS 0.105404f
C23482 VDD.t2261 VSS 0.066856f
C23483 VDD.n5506 VSS 0.14405f
C23484 VDD.n5507 VSS 0.120118f
C23485 VDD.n5508 VSS 0.016021f
C23486 VDD.t1382 VSS 0.025104f
C23487 VDD.n5509 VSS 0.116823f
C23488 VDD.t4562 VSS 0.066856f
C23489 VDD.n5510 VSS 0.14405f
C23490 VDD.t3400 VSS 0.025104f
C23491 VDD.t2974 VSS 0.066856f
C23492 VDD.n5511 VSS 0.14405f
C23493 VDD.t612 VSS 0.025104f
C23494 VDD.n5512 VSS 0.033925f
C23495 VDD.t4784 VSS 0.019767f
C23496 VDD.t4782 VSS 0.018805f
C23497 VDD.n5513 VSS 0.054793f
C23498 VDD.t4783 VSS 0.018792f
C23499 VDD.t4785 VSS 0.019781f
C23500 VDD.n5514 VSS 0.077486f
C23501 VDD.n5515 VSS 0.252514f
C23502 VDD.n5516 VSS 0.199549f
C23503 VDD.n5517 VSS 0.060108f
C23504 VDD.t611 VSS 0.066856f
C23505 VDD.n5518 VSS 0.131361f
C23506 VDD.n5519 VSS 0.120118f
C23507 VDD.n5520 VSS 0.016021f
C23508 VDD.t2975 VSS 0.025104f
C23509 VDD.n5521 VSS 0.105404f
C23510 VDD.n5522 VSS 0.057098f
C23511 VDD.n5523 VSS 0.087217f
C23512 VDD.t3399 VSS 0.066856f
C23513 VDD.n5524 VSS 0.14405f
C23514 VDD.n5525 VSS 0.120118f
C23515 VDD.n5526 VSS 0.016021f
C23516 VDD.t4563 VSS 0.025104f
C23517 VDD.n5527 VSS 0.116823f
C23518 VDD.n5528 VSS 0.173497f
C23519 VDD.n5529 VSS 0.122652f
C23520 VDD.n5531 VSS 0.018625f
C23521 VDD.n5533 VSS 0.01502f
C23522 VDD.n5534 VSS 0.437162f
C23523 VDD.n5535 VSS 0.01487f
C23524 VDD.n5537 VSS 0.018249f
C23525 VDD.n5538 VSS 0.203639f
C23526 VDD.n5539 VSS 0.77149f
C23527 VDD.n5540 VSS 0.009688f
C23528 VDD.t3214 VSS 0.066856f
C23529 VDD.n5542 VSS 0.125227f
C23530 VDD.t870 VSS 0.025104f
C23531 VDD.t1340 VSS 0.066856f
C23532 VDD.n5543 VSS 0.125227f
C23533 VDD.t2819 VSS 0.025104f
C23534 VDD.n5544 VSS 0.006598f
C23535 VDD.t2818 VSS 0.066856f
C23536 VDD.n5545 VSS 0.045867f
C23537 VDD.n5546 VSS 0.015693f
C23538 VDD.t1514 VSS 0.066856f
C23539 VDD.n5547 VSS 0.125227f
C23540 VDD.t3392 VSS 0.025104f
C23541 VDD.t3906 VSS 0.066856f
C23542 VDD.n5548 VSS 0.125227f
C23543 VDD.t2985 VSS 0.025104f
C23544 VDD.t3747 VSS 0.066856f
C23545 VDD.n5549 VSS 0.125227f
C23546 VDD.t2924 VSS 0.025104f
C23547 VDD.t3365 VSS 0.066856f
C23548 VDD.n5550 VSS 0.125227f
C23549 VDD.t4725 VSS 0.025104f
C23550 VDD.t3266 VSS 0.066856f
C23551 VDD.n5551 VSS 0.125227f
C23552 VDD.t2381 VSS 0.025104f
C23553 VDD.t1393 VSS 0.066856f
C23554 VDD.n5552 VSS 0.125227f
C23555 VDD.t4211 VSS 0.025104f
C23556 VDD.n5553 VSS 0.006598f
C23557 VDD.t4210 VSS 0.066856f
C23558 VDD.n5554 VSS 0.045867f
C23559 VDD.n5555 VSS 0.015693f
C23560 VDD.n5556 VSS 0.035132f
C23561 VDD.n5557 VSS 0.010188f
C23562 VDD.t515 VSS 0.020392f
C23563 VDD.t516 VSS 0.022133f
C23564 VDD.n5558 VSS 0.069721f
C23565 VDD.n5559 VSS 0.040089f
C23566 VDD.t518 VSS 0.020371f
C23567 VDD.n5560 VSS 0.027146f
C23568 VDD.t519 VSS 0.022106f
C23569 VDD.n5561 VSS 0.036568f
C23570 VDD.n5562 VSS 0.044801f
C23571 VDD.n5563 VSS 0.278297f
C23572 VDD.n5564 VSS 0.040089f
C23573 VDD.t517 VSS 0.020371f
C23574 VDD.n5565 VSS 0.027146f
C23575 VDD.t514 VSS 0.020392f
C23576 VDD.n5566 VSS 0.049654f
C23577 VDD.t499 VSS 0.017093f
C23578 VDD.n5567 VSS 0.042096f
C23579 VDD.n5568 VSS 0.069466f
C23580 VDD.t513 VSS 0.017093f
C23581 VDD.n5569 VSS 0.035464f
C23582 VDD.n5570 VSS 0.016538f
C23583 VDD.n5571 VSS 0.027213f
C23584 VDD.n5572 VSS 0.204333f
C23585 VDD.n5573 VSS 0.030906f
C23586 VDD.n5574 VSS 0.010881f
C23587 VDD.n5575 VSS 0.044227f
C23588 VDD.n5576 VSS 0.094696f
C23589 VDD.n5577 VSS 0.016021f
C23590 VDD.t1394 VSS 0.025104f
C23591 VDD.n5578 VSS 0.083673f
C23592 VDD.n5579 VSS 0.048151f
C23593 VDD.n5580 VSS 0.081176f
C23594 VDD.t2380 VSS 0.066856f
C23595 VDD.n5581 VSS 0.125227f
C23596 VDD.n5582 VSS 0.101294f
C23597 VDD.n5583 VSS 0.016021f
C23598 VDD.t3267 VSS 0.025104f
C23599 VDD.n5584 VSS 0.099723f
C23600 VDD.t2750 VSS 0.028519f
C23601 VDD.t2405 VSS 0.028519f
C23602 VDD.n5585 VSS 0.009191f
C23603 VDD.t2749 VSS 0.066856f
C23604 VDD.t2152 VSS 0.066856f
C23605 VDD.t2377 VSS 0.028519f
C23606 VDD.t1972 VSS 0.028519f
C23607 VDD.n5586 VSS 0.009191f
C23608 VDD.t2376 VSS 0.066856f
C23609 VDD.t1757 VSS 0.066856f
C23610 VDD.t676 VSS 0.066856f
C23611 VDD.t4322 VSS 0.066856f
C23612 VDD.t2012 VSS 0.066856f
C23613 VDD.t4488 VSS 0.066856f
C23614 VDD.n5587 VSS 0.690489f
C23615 VDD.t3624 VSS 0.066856f
C23616 VDD.t1971 VSS 0.066856f
C23617 VDD.n5588 VSS 0.690489f
C23618 VDD.t1758 VSS 0.028519f
C23619 VDD.t3625 VSS 0.028519f
C23620 VDD.n5589 VSS 0.009191f
C23621 VDD.n5590 VSS 0.644755f
C23622 VDD.t3988 VSS 0.066856f
C23623 VDD.t2404 VSS 0.066856f
C23624 VDD.n5591 VSS 0.709674f
C23625 VDD.t2153 VSS 0.028519f
C23626 VDD.t3989 VSS 0.028519f
C23627 VDD.n5592 VSS 0.009191f
C23628 VDD.n5593 VSS 0.261039f
C23629 VDD.n5594 VSS 0.62132f
C23630 VDD.n5595 VSS 0.099723f
C23631 VDD.t4724 VSS 0.066856f
C23632 VDD.n5596 VSS 0.125227f
C23633 VDD.n5597 VSS 0.101294f
C23634 VDD.n5598 VSS 0.016021f
C23635 VDD.t3366 VSS 0.025104f
C23636 VDD.n5599 VSS 0.083673f
C23637 VDD.n5600 VSS 0.048151f
C23638 VDD.n5601 VSS 0.081176f
C23639 VDD.t2922 VSS 0.066856f
C23640 VDD.n5602 VSS 0.125227f
C23641 VDD.n5603 VSS 0.101294f
C23642 VDD.n5604 VSS 0.016021f
C23643 VDD.t3749 VSS 0.025104f
C23644 VDD.n5605 VSS 0.099723f
C23645 VDD.t829 VSS 0.028519f
C23646 VDD.t4625 VSS 0.028519f
C23647 VDD.n5606 VSS 0.009191f
C23648 VDD.t828 VSS 0.066856f
C23649 VDD.t4448 VSS 0.066856f
C23650 VDD.t4601 VSS 0.028519f
C23651 VDD.t4289 VSS 0.028519f
C23652 VDD.n5607 VSS 0.009191f
C23653 VDD.t4600 VSS 0.066856f
C23654 VDD.t4122 VSS 0.066856f
C23655 VDD.t3080 VSS 0.066856f
C23656 VDD.t2574 VSS 0.066856f
C23657 VDD.t4324 VSS 0.066856f
C23658 VDD.t2759 VSS 0.066856f
C23659 VDD.n5608 VSS 0.690489f
C23660 VDD.t1759 VSS 0.066856f
C23661 VDD.t4288 VSS 0.066856f
C23662 VDD.n5609 VSS 0.690489f
C23663 VDD.t4123 VSS 0.028519f
C23664 VDD.t1760 VSS 0.028519f
C23665 VDD.n5610 VSS 0.009191f
C23666 VDD.n5611 VSS 0.644755f
C23667 VDD.t2154 VSS 0.066856f
C23668 VDD.t4624 VSS 0.066856f
C23669 VDD.n5612 VSS 0.709674f
C23670 VDD.t4449 VSS 0.028519f
C23671 VDD.t2155 VSS 0.028519f
C23672 VDD.n5613 VSS 0.009191f
C23673 VDD.n5614 VSS 0.261039f
C23674 VDD.n5615 VSS 0.62132f
C23675 VDD.n5616 VSS 0.099723f
C23676 VDD.t2984 VSS 0.066856f
C23677 VDD.n5617 VSS 0.125227f
C23678 VDD.n5618 VSS 0.101294f
C23679 VDD.n5619 VSS 0.016021f
C23680 VDD.t3907 VSS 0.025104f
C23681 VDD.n5620 VSS 0.083673f
C23682 VDD.n5621 VSS 0.048151f
C23683 VDD.n5622 VSS 0.081176f
C23684 VDD.t3391 VSS 0.066856f
C23685 VDD.n5623 VSS 0.125227f
C23686 VDD.n5624 VSS 0.101294f
C23687 VDD.n5625 VSS 0.016021f
C23688 VDD.t1515 VSS 0.025104f
C23689 VDD.n5626 VSS 0.099723f
C23690 VDD.t2851 VSS 0.028519f
C23691 VDD.t1031 VSS 0.028519f
C23692 VDD.n5627 VSS 0.009191f
C23693 VDD.t2850 VSS 0.066856f
C23694 VDD.t3294 VSS 0.066856f
C23695 VDD.t2495 VSS 0.028519f
C23696 VDD.t663 VSS 0.028519f
C23697 VDD.n5628 VSS 0.009191f
C23698 VDD.t2494 VSS 0.066856f
C23699 VDD.t2988 VSS 0.066856f
C23700 VDD.t800 VSS 0.066856f
C23701 VDD.t1264 VSS 0.066856f
C23702 VDD.t4186 VSS 0.066856f
C23703 VDD.t3274 VSS 0.066856f
C23704 VDD.n5629 VSS 0.696076f
C23705 VDD.t1606 VSS 0.066856f
C23706 VDD.t662 VSS 0.066856f
C23707 VDD.n5630 VSS 0.696076f
C23708 VDD.t2989 VSS 0.028519f
C23709 VDD.t1607 VSS 0.028519f
C23710 VDD.n5631 VSS 0.009191f
C23711 VDD.n5632 VSS 0.650522f
C23712 VDD.t1975 VSS 0.066856f
C23713 VDD.t1030 VSS 0.066856f
C23714 VDD.n5633 VSS 0.715442f
C23715 VDD.t3295 VSS 0.028519f
C23716 VDD.t1976 VSS 0.028519f
C23717 VDD.n5634 VSS 0.009191f
C23718 VDD.n5635 VSS 0.263202f
C23719 VDD.n5636 VSS 0.62638f
C23720 VDD.n5637 VSS 0.08403f
C23721 VDD.n5638 VSS 0.035132f
C23722 VDD.n5639 VSS 0.010188f
C23723 VDD.t4749 VSS 0.020392f
C23724 VDD.t4750 VSS 0.022133f
C23725 VDD.n5640 VSS 0.069721f
C23726 VDD.n5641 VSS 0.040089f
C23727 VDD.t4754 VSS 0.020371f
C23728 VDD.n5642 VSS 0.027146f
C23729 VDD.t4755 VSS 0.022106f
C23730 VDD.n5643 VSS 0.036568f
C23731 VDD.n5644 VSS 0.044801f
C23732 VDD.n5645 VSS 0.278297f
C23733 VDD.n5646 VSS 0.040089f
C23734 VDD.t4753 VSS 0.020371f
C23735 VDD.n5647 VSS 0.027146f
C23736 VDD.t4748 VSS 0.020392f
C23737 VDD.n5648 VSS 0.049654f
C23738 VDD.t4752 VSS 0.017093f
C23739 VDD.n5649 VSS 0.042096f
C23740 VDD.n5650 VSS 0.069466f
C23741 VDD.t4751 VSS 0.017093f
C23742 VDD.n5651 VSS 0.035464f
C23743 VDD.n5652 VSS 0.016538f
C23744 VDD.n5653 VSS 0.027213f
C23745 VDD.n5654 VSS 0.204333f
C23746 VDD.n5655 VSS 0.030906f
C23747 VDD.n5656 VSS 0.010881f
C23748 VDD.n5657 VSS 0.044227f
C23749 VDD.n5658 VSS 0.094696f
C23750 VDD.n5659 VSS 0.016021f
C23751 VDD.t1342 VSS 0.025104f
C23752 VDD.n5660 VSS 0.083673f
C23753 VDD.n5661 VSS 0.048151f
C23754 VDD.n5662 VSS 0.081176f
C23755 VDD.t868 VSS 0.066856f
C23756 VDD.n5663 VSS 0.125227f
C23757 VDD.n5664 VSS 0.101294f
C23758 VDD.n5665 VSS 0.016021f
C23759 VDD.t3215 VSS 0.025104f
C23760 VDD.n5666 VSS 0.099723f
C23761 VDD.t4676 VSS 0.066856f
C23762 VDD.n5667 VSS 0.125227f
C23763 VDD.t1889 VSS 0.025104f
C23764 VDD.t935 VSS 0.066856f
C23765 VDD.n5668 VSS 0.125227f
C23766 VDD.t3698 VSS 0.025104f
C23767 VDD.t4445 VSS 0.028519f
C23768 VDD.t2142 VSS 0.028519f
C23769 VDD.n5669 VSS 0.009191f
C23770 VDD.t4444 VSS 0.066856f
C23771 VDD.t1946 VSS 0.066856f
C23772 VDD.t4119 VSS 0.028519f
C23773 VDD.t1754 VSS 0.028519f
C23774 VDD.n5670 VSS 0.009191f
C23775 VDD.t4118 VSS 0.066856f
C23776 VDD.t1582 VSS 0.066856f
C23777 VDD.t2571 VSS 0.066856f
C23778 VDD.t4160 VSS 0.066856f
C23779 VDD.t3814 VSS 0.066856f
C23780 VDD.t4320 VSS 0.066856f
C23781 VDD.n5671 VSS 0.690489f
C23782 VDD.t1241 VSS 0.066856f
C23783 VDD.t1753 VSS 0.066856f
C23784 VDD.n5672 VSS 0.690489f
C23785 VDD.t1583 VSS 0.028519f
C23786 VDD.t1242 VSS 0.028519f
C23787 VDD.n5673 VSS 0.009191f
C23788 VDD.n5674 VSS 0.644755f
C23789 VDD.t1602 VSS 0.066856f
C23790 VDD.t2141 VSS 0.066856f
C23791 VDD.n5675 VSS 0.709674f
C23792 VDD.t1947 VSS 0.028519f
C23793 VDD.t1603 VSS 0.028519f
C23794 VDD.n5676 VSS 0.009191f
C23795 VDD.n5677 VSS 0.261039f
C23796 VDD.t2925 VSS 0.066856f
C23797 VDD.n5678 VSS 0.125227f
C23798 VDD.t3751 VSS 0.025104f
C23799 VDD.t4626 VSS 0.066856f
C23800 VDD.n5679 VSS 0.125227f
C23801 VDD.t1844 VSS 0.025104f
C23802 VDD.n5680 VSS 0.035132f
C23803 VDD.t3594 VSS 0.025104f
C23804 VDD.t3458 VSS 0.066856f
C23805 VDD.n5681 VSS 0.125227f
C23806 VDD.t648 VSS 0.025104f
C23807 VDD.t2543 VSS 0.028519f
C23808 VDD.t1520 VSS 0.028519f
C23809 VDD.n5682 VSS 0.009191f
C23810 VDD.t2542 VSS 0.066856f
C23811 VDD.t4130 VSS 0.066856f
C23812 VDD.t2108 VSS 0.028519f
C23813 VDD.t1174 VSS 0.028519f
C23814 VDD.n5683 VSS 0.009191f
C23815 VDD.t2107 VSS 0.066856f
C23816 VDD.t3760 VSS 0.066856f
C23817 VDD.t4628 VSS 0.066856f
C23818 VDD.t2156 VSS 0.066856f
C23819 VDD.t782 VSS 0.066856f
C23820 VDD.t3737 VSS 0.066856f
C23821 VDD.n5684 VSS 0.690489f
C23822 VDD.t2458 VSS 0.066856f
C23823 VDD.t1173 VSS 0.066856f
C23824 VDD.n5685 VSS 0.690489f
C23825 VDD.t3761 VSS 0.028519f
C23826 VDD.t2459 VSS 0.028519f
C23827 VDD.n5686 VSS 0.009191f
C23828 VDD.n5687 VSS 0.644755f
C23829 VDD.t2816 VSS 0.066856f
C23830 VDD.t1519 VSS 0.066856f
C23831 VDD.n5688 VSS 0.709674f
C23832 VDD.t4131 VSS 0.028519f
C23833 VDD.t2817 VSS 0.028519f
C23834 VDD.n5689 VSS 0.009191f
C23835 VDD.n5690 VSS 0.261039f
C23836 VDD.t871 VSS 0.066856f
C23837 VDD.n5691 VSS 0.125227f
C23838 VDD.t1729 VSS 0.025104f
C23839 VDD.t3984 VSS 0.066856f
C23840 VDD.n5692 VSS 0.125227f
C23841 VDD.t1178 VSS 0.025104f
C23842 VDD.t1363 VSS 0.066856f
C23843 VDD.n5693 VSS 0.125227f
C23844 VDD.t2367 VSS 0.025104f
C23845 VDD.t2143 VSS 0.066856f
C23846 VDD.n5694 VSS 0.125227f
C23847 VDD.t3525 VSS 0.025104f
C23848 VDD.t1141 VSS 0.028519f
C23849 VDD.t3949 VSS 0.028519f
C23850 VDD.n5695 VSS 0.009191f
C23851 VDD.t1140 VSS 0.066856f
C23852 VDD.t946 VSS 0.066856f
C23853 VDD.t807 VSS 0.028519f
C23854 VDD.t3586 VSS 0.028519f
C23855 VDD.n5696 VSS 0.009191f
C23856 VDD.t806 VSS 0.066856f
C23857 VDD.t4712 VSS 0.066856f
C23858 VDD.t3352 VSS 0.066856f
C23859 VDD.t3168 VSS 0.066856f
C23860 VDD.t3012 VSS 0.066856f
C23861 VDD.t1969 VSS 0.066856f
C23862 VDD.n5697 VSS 0.696076f
C23863 VDD.t4508 VSS 0.066856f
C23864 VDD.t3585 VSS 0.066856f
C23865 VDD.n5698 VSS 0.696076f
C23866 VDD.t4713 VSS 0.028519f
C23867 VDD.t4509 VSS 0.028519f
C23868 VDD.n5699 VSS 0.009191f
C23869 VDD.n5700 VSS 0.650522f
C23870 VDD.t747 VSS 0.066856f
C23871 VDD.t3948 VSS 0.066856f
C23872 VDD.n5701 VSS 0.715442f
C23873 VDD.t948 VSS 0.028519f
C23874 VDD.t749 VSS 0.028519f
C23875 VDD.n5702 VSS 0.009191f
C23876 VDD.n5703 VSS 0.263202f
C23877 VDD.n5704 VSS 0.035132f
C23878 VDD.t1663 VSS 0.025104f
C23879 VDD.t2657 VSS 0.066856f
C23880 VDD.n5705 VSS 0.125227f
C23881 VDD.t3491 VSS 0.025104f
C23882 VDD.t3648 VSS 0.066856f
C23883 VDD.n5706 VSS 0.125227f
C23884 VDD.t1228 VSS 0.025104f
C23885 VDD.t732 VSS 0.066856f
C23886 VDD.n5707 VSS 0.125227f
C23887 VDD.t1618 VSS 0.025104f
C23888 VDD.t2129 VSS 0.028519f
C23889 VDD.t2614 VSS 0.028519f
C23890 VDD.n5708 VSS 0.009191f
C23891 VDD.t2128 VSS 0.066856f
C23892 VDD.t4706 VSS 0.066856f
C23893 VDD.t1741 VSS 0.028519f
C23894 VDD.t2187 VSS 0.028519f
C23895 VDD.n5709 VSS 0.009191f
C23896 VDD.t1740 VSS 0.066856f
C23897 VDD.t4358 VSS 0.066856f
C23898 VDD.t4306 VSS 0.066856f
C23899 VDD.t2836 VSS 0.066856f
C23900 VDD.t4560 VSS 0.066856f
C23901 VDD.t4702 VSS 0.066856f
C23902 VDD.n5710 VSS 0.690489f
C23903 VDD.t2068 VSS 0.066856f
C23904 VDD.t2186 VSS 0.066856f
C23905 VDD.n5711 VSS 0.690489f
C23906 VDD.t4359 VSS 0.028519f
C23907 VDD.t2069 VSS 0.028519f
C23908 VDD.n5712 VSS 0.009191f
C23909 VDD.n5713 VSS 0.644755f
C23910 VDD.t2490 VSS 0.066856f
C23911 VDD.t2613 VSS 0.066856f
C23912 VDD.n5714 VSS 0.709674f
C23913 VDD.t4707 VSS 0.028519f
C23914 VDD.t2491 VSS 0.028519f
C23915 VDD.n5715 VSS 0.009191f
C23916 VDD.n5716 VSS 0.261039f
C23917 VDD.t4222 VSS 0.066856f
C23918 VDD.n5717 VSS 0.125227f
C23919 VDD.t1756 VSS 0.025104f
C23920 VDD.t1755 VSS 0.066856f
C23921 VDD.n5718 VSS 0.125227f
C23922 VDD.n5719 VSS 0.101294f
C23923 VDD.n5720 VSS 0.016021f
C23924 VDD.t4223 VSS 0.025104f
C23925 VDD.n5721 VSS 0.099723f
C23926 VDD.n5722 VSS 0.62132f
C23927 VDD.n5723 VSS 0.099723f
C23928 VDD.t1617 VSS 0.066856f
C23929 VDD.n5724 VSS 0.125227f
C23930 VDD.n5725 VSS 0.101294f
C23931 VDD.n5726 VSS 0.016021f
C23932 VDD.t733 VSS 0.025104f
C23933 VDD.n5727 VSS 0.081176f
C23934 VDD.n5728 VSS 0.048151f
C23935 VDD.n5729 VSS 0.083673f
C23936 VDD.t1227 VSS 0.066856f
C23937 VDD.n5730 VSS 0.125227f
C23938 VDD.n5731 VSS 0.101294f
C23939 VDD.n5732 VSS 0.016021f
C23940 VDD.t3649 VSS 0.025104f
C23941 VDD.n5733 VSS 0.099723f
C23942 VDD.t1560 VSS 0.028519f
C23943 VDD.t4357 VSS 0.028519f
C23944 VDD.n5734 VSS 0.009191f
C23945 VDD.t1559 VSS 0.066856f
C23946 VDD.t4190 VSS 0.066856f
C23947 VDD.t1203 VSS 0.028519f
C23948 VDD.t4021 VSS 0.028519f
C23949 VDD.n5735 VSS 0.009191f
C23950 VDD.t1202 VSS 0.066856f
C23951 VDD.t3824 VSS 0.066856f
C23952 VDD.t3778 VSS 0.066856f
C23953 VDD.t2236 VSS 0.066856f
C23954 VDD.t4056 VSS 0.066856f
C23955 VDD.t2487 VSS 0.066856f
C23956 VDD.n5736 VSS 0.690489f
C23957 VDD.t1481 VSS 0.066856f
C23958 VDD.t4020 VSS 0.066856f
C23959 VDD.n5737 VSS 0.690489f
C23960 VDD.t3825 VSS 0.028519f
C23961 VDD.t1482 VSS 0.028519f
C23962 VDD.n5738 VSS 0.009191f
C23963 VDD.n5739 VSS 0.644755f
C23964 VDD.t1847 VSS 0.066856f
C23965 VDD.t4356 VSS 0.066856f
C23966 VDD.n5740 VSS 0.709674f
C23967 VDD.t4191 VSS 0.028519f
C23968 VDD.t1848 VSS 0.028519f
C23969 VDD.n5741 VSS 0.009191f
C23970 VDD.n5742 VSS 0.261039f
C23971 VDD.n5743 VSS 0.62132f
C23972 VDD.n5744 VSS 0.099723f
C23973 VDD.t3490 VSS 0.066856f
C23974 VDD.n5745 VSS 0.125227f
C23975 VDD.n5746 VSS 0.101294f
C23976 VDD.n5747 VSS 0.016021f
C23977 VDD.t2658 VSS 0.025104f
C23978 VDD.n5748 VSS 0.081176f
C23979 VDD.n5749 VSS 0.048151f
C23980 VDD.n5750 VSS 0.083673f
C23981 VDD.t1662 VSS 0.066856f
C23982 VDD.n5751 VSS 0.125227f
C23983 VDD.n5752 VSS 0.006598f
C23984 VDD.t1318 VSS 0.066856f
C23985 VDD.n5753 VSS 0.045867f
C23986 VDD.n5754 VSS 0.015693f
C23987 VDD.n5755 VSS 0.010188f
C23988 VDD.t326 VSS 0.020392f
C23989 VDD.t367 VSS 0.022133f
C23990 VDD.n5756 VSS 0.069721f
C23991 VDD.n5757 VSS 0.040089f
C23992 VDD.t418 VSS 0.020371f
C23993 VDD.n5758 VSS 0.027146f
C23994 VDD.t302 VSS 0.022106f
C23995 VDD.n5759 VSS 0.036568f
C23996 VDD.n5760 VSS 0.044801f
C23997 VDD.n5761 VSS 0.278297f
C23998 VDD.n5762 VSS 0.040089f
C23999 VDD.t419 VSS 0.020371f
C24000 VDD.n5763 VSS 0.027146f
C24001 VDD.t368 VSS 0.020392f
C24002 VDD.n5764 VSS 0.049654f
C24003 VDD.t369 VSS 0.017093f
C24004 VDD.n5765 VSS 0.042096f
C24005 VDD.n5766 VSS 0.069466f
C24006 VDD.t421 VSS 0.017093f
C24007 VDD.n5767 VSS 0.035464f
C24008 VDD.n5768 VSS 0.016538f
C24009 VDD.n5769 VSS 0.027213f
C24010 VDD.n5770 VSS 0.204333f
C24011 VDD.n5771 VSS 0.030906f
C24012 VDD.n5772 VSS 0.010881f
C24013 VDD.n5773 VSS 0.044227f
C24014 VDD.n5774 VSS 0.094696f
C24015 VDD.n5775 VSS 0.016021f
C24016 VDD.t1319 VSS 0.025104f
C24017 VDD.n5776 VSS 0.08403f
C24018 VDD.n5777 VSS 0.62638f
C24019 VDD.n5778 VSS 0.099723f
C24020 VDD.t3524 VSS 0.066856f
C24021 VDD.n5779 VSS 0.125227f
C24022 VDD.n5780 VSS 0.101294f
C24023 VDD.n5781 VSS 0.016021f
C24024 VDD.t2144 VSS 0.025104f
C24025 VDD.n5782 VSS 0.081176f
C24026 VDD.n5783 VSS 0.048151f
C24027 VDD.n5784 VSS 0.083673f
C24028 VDD.t2366 VSS 0.066856f
C24029 VDD.n5785 VSS 0.125227f
C24030 VDD.n5786 VSS 0.101294f
C24031 VDD.n5787 VSS 0.016021f
C24032 VDD.t1364 VSS 0.025104f
C24033 VDD.n5788 VSS 0.099723f
C24034 VDD.t3069 VSS 0.028519f
C24035 VDD.t1599 VSS 0.028519f
C24036 VDD.n5789 VSS 0.009191f
C24037 VDD.t3068 VSS 0.066856f
C24038 VDD.t4642 VSS 0.066856f
C24039 VDD.t2729 VSS 0.028519f
C24040 VDD.t1238 VSS 0.028519f
C24041 VDD.n5790 VSS 0.009191f
C24042 VDD.t2728 VSS 0.066856f
C24043 VDD.t4292 VSS 0.066856f
C24044 VDD.t1032 VSS 0.066856f
C24045 VDD.t2778 VSS 0.066856f
C24046 VDD.t1284 VSS 0.066856f
C24047 VDD.t3804 VSS 0.066856f
C24048 VDD.n5791 VSS 0.690489f
C24049 VDD.t3008 VSS 0.066856f
C24050 VDD.t1237 VSS 0.066856f
C24051 VDD.n5792 VSS 0.690489f
C24052 VDD.t4293 VSS 0.028519f
C24053 VDD.t3009 VSS 0.028519f
C24054 VDD.n5793 VSS 0.009191f
C24055 VDD.n5794 VSS 0.644755f
C24056 VDD.t3306 VSS 0.066856f
C24057 VDD.t1598 VSS 0.066856f
C24058 VDD.n5795 VSS 0.709674f
C24059 VDD.t4643 VSS 0.028519f
C24060 VDD.t3307 VSS 0.028519f
C24061 VDD.n5796 VSS 0.009191f
C24062 VDD.n5797 VSS 0.261039f
C24063 VDD.n5798 VSS 0.62132f
C24064 VDD.n5799 VSS 0.099723f
C24065 VDD.t1177 VSS 0.066856f
C24066 VDD.n5800 VSS 0.125227f
C24067 VDD.n5801 VSS 0.101294f
C24068 VDD.n5802 VSS 0.016021f
C24069 VDD.t3985 VSS 0.025104f
C24070 VDD.n5803 VSS 0.081176f
C24071 VDD.n5804 VSS 0.048151f
C24072 VDD.n5805 VSS 0.083673f
C24073 VDD.t1728 VSS 0.066856f
C24074 VDD.n5806 VSS 0.125227f
C24075 VDD.n5807 VSS 0.101294f
C24076 VDD.n5808 VSS 0.016021f
C24077 VDD.t872 VSS 0.025104f
C24078 VDD.n5809 VSS 0.099723f
C24079 VDD.n5810 VSS 0.62132f
C24080 VDD.n5811 VSS 0.099723f
C24081 VDD.t646 VSS 0.066856f
C24082 VDD.n5812 VSS 0.125227f
C24083 VDD.n5813 VSS 0.101294f
C24084 VDD.n5814 VSS 0.016021f
C24085 VDD.t3459 VSS 0.025104f
C24086 VDD.n5815 VSS 0.081176f
C24087 VDD.n5816 VSS 0.048151f
C24088 VDD.n5817 VSS 0.083673f
C24089 VDD.t3593 VSS 0.066856f
C24090 VDD.n5818 VSS 0.125227f
C24091 VDD.n5819 VSS 0.006598f
C24092 VDD.t2775 VSS 0.066856f
C24093 VDD.n5820 VSS 0.045867f
C24094 VDD.n5821 VSS 0.015693f
C24095 VDD.n5822 VSS 0.010188f
C24096 VDD.t4795 VSS 0.020392f
C24097 VDD.t4797 VSS 0.022133f
C24098 VDD.n5823 VSS 0.069721f
C24099 VDD.n5824 VSS 0.040089f
C24100 VDD.t4793 VSS 0.020371f
C24101 VDD.n5825 VSS 0.027146f
C24102 VDD.t4796 VSS 0.022106f
C24103 VDD.n5826 VSS 0.036568f
C24104 VDD.n5827 VSS 0.044801f
C24105 VDD.n5828 VSS 0.278297f
C24106 VDD.n5829 VSS 0.040089f
C24107 VDD.t4792 VSS 0.020371f
C24108 VDD.n5830 VSS 0.027146f
C24109 VDD.t4794 VSS 0.020392f
C24110 VDD.n5831 VSS 0.049654f
C24111 VDD.t4799 VSS 0.017093f
C24112 VDD.n5832 VSS 0.042096f
C24113 VDD.n5833 VSS 0.069466f
C24114 VDD.t4798 VSS 0.017093f
C24115 VDD.n5834 VSS 0.035464f
C24116 VDD.n5835 VSS 0.016538f
C24117 VDD.n5836 VSS 0.027213f
C24118 VDD.n5837 VSS 0.204333f
C24119 VDD.n5838 VSS 0.030906f
C24120 VDD.n5839 VSS 0.010881f
C24121 VDD.n5840 VSS 0.044227f
C24122 VDD.n5841 VSS 0.094696f
C24123 VDD.n5842 VSS 0.016021f
C24124 VDD.t2777 VSS 0.025104f
C24125 VDD.n5843 VSS 0.08403f
C24126 VDD.t859 VSS 0.028519f
C24127 VDD.t4105 VSS 0.028519f
C24128 VDD.n5844 VSS 0.009191f
C24129 VDD.t857 VSS 0.066856f
C24130 VDD.t1769 VSS 0.066856f
C24131 VDD.t4623 VSS 0.028519f
C24132 VDD.t3730 VSS 0.028519f
C24133 VDD.n5845 VSS 0.009191f
C24134 VDD.t4622 VSS 0.066856f
C24135 VDD.t1413 VSS 0.066856f
C24136 VDD.t3094 VSS 0.066856f
C24137 VDD.t3992 VSS 0.066856f
C24138 VDD.t2681 VSS 0.066856f
C24139 VDD.t2121 VSS 0.066856f
C24140 VDD.n5846 VSS 0.696076f
C24141 VDD.t4234 VSS 0.066856f
C24142 VDD.t3729 VSS 0.066856f
C24143 VDD.n5847 VSS 0.696076f
C24144 VDD.t1414 VSS 0.028519f
C24145 VDD.t4235 VSS 0.028519f
C24146 VDD.n5848 VSS 0.009191f
C24147 VDD.n5849 VSS 0.650522f
C24148 VDD.t4538 VSS 0.066856f
C24149 VDD.t4104 VSS 0.066856f
C24150 VDD.n5850 VSS 0.715442f
C24151 VDD.t1770 VSS 0.028519f
C24152 VDD.t4539 VSS 0.028519f
C24153 VDD.n5851 VSS 0.009191f
C24154 VDD.n5852 VSS 0.263202f
C24155 VDD.n5853 VSS 0.62638f
C24156 VDD.n5854 VSS 0.099723f
C24157 VDD.t1842 VSS 0.066856f
C24158 VDD.n5855 VSS 0.125227f
C24159 VDD.n5856 VSS 0.101294f
C24160 VDD.n5857 VSS 0.016021f
C24161 VDD.t4627 VSS 0.025104f
C24162 VDD.n5858 VSS 0.081176f
C24163 VDD.n5859 VSS 0.048151f
C24164 VDD.n5860 VSS 0.083673f
C24165 VDD.t3750 VSS 0.066856f
C24166 VDD.n5861 VSS 0.125227f
C24167 VDD.n5862 VSS 0.101294f
C24168 VDD.n5863 VSS 0.016021f
C24169 VDD.t2927 VSS 0.025104f
C24170 VDD.n5864 VSS 0.099723f
C24171 VDD.n5865 VSS 0.62132f
C24172 VDD.n5866 VSS 0.099723f
C24173 VDD.t3697 VSS 0.066856f
C24174 VDD.n5867 VSS 0.125227f
C24175 VDD.n5868 VSS 0.101294f
C24176 VDD.n5869 VSS 0.016021f
C24177 VDD.t936 VSS 0.025104f
C24178 VDD.n5870 VSS 0.081176f
C24179 VDD.n5871 VSS 0.048151f
C24180 VDD.n5872 VSS 0.083673f
C24181 VDD.t1888 VSS 0.066856f
C24182 VDD.n5873 VSS 0.125227f
C24183 VDD.n5874 VSS 0.101294f
C24184 VDD.n5875 VSS 0.016021f
C24185 VDD.t4677 VSS 0.025104f
C24186 VDD.n5876 VSS 0.099723f
C24187 VDD.t3923 VSS 0.028519f
C24188 VDD.t1579 VSS 0.028519f
C24189 VDD.n5877 VSS 0.009191f
C24190 VDD.t3922 VSS 0.066856f
C24191 VDD.t3796 VSS 0.066856f
C24192 VDD.t3565 VSS 0.028519f
C24193 VDD.t1226 VSS 0.028519f
C24194 VDD.n5878 VSS 0.009191f
C24195 VDD.t3564 VSS 0.066856f
C24196 VDD.t3462 VSS 0.066856f
C24197 VDD.t1937 VSS 0.066856f
C24198 VDD.t1800 VSS 0.066856f
C24199 VDD.t1939 VSS 0.028519f
C24200 VDD.t3791 VSS 0.028519f
C24201 VDD.n5879 VSS 0.009191f
C24202 VDD.n5880 VSS 0.018249f
C24203 VDD.n5881 VSS 0.018625f
C24204 VDD.n5883 VSS 0.01502f
C24205 VDD.n5885 VSS 0.01487f
C24206 VDD.n5886 VSS 0.009312f
C24207 VDD.n5888 VSS 0.009688f
C24208 VDD.n5890 VSS 0.271342f
C24209 VDD.t1802 VSS 0.028519f
C24210 VDD.t1960 VSS 0.028519f
C24211 VDD.n5891 VSS 0.009191f
C24212 VDD.n5892 VSS 0.43097f
C24213 VDD.t1958 VSS 0.066856f
C24214 VDD.t3790 VSS 0.066856f
C24215 VDD.n5893 VSS 0.690489f
C24216 VDD.t3579 VSS 0.066856f
C24217 VDD.t1225 VSS 0.066856f
C24218 VDD.n5894 VSS 0.690489f
C24219 VDD.t3463 VSS 0.028519f
C24220 VDD.t3580 VSS 0.028519f
C24221 VDD.n5895 VSS 0.009191f
C24222 VDD.n5896 VSS 0.644755f
C24223 VDD.t3940 VSS 0.066856f
C24224 VDD.t1578 VSS 0.066856f
C24225 VDD.n5897 VSS 0.709674f
C24226 VDD.t3797 VSS 0.028519f
C24227 VDD.t3941 VSS 0.028519f
C24228 VDD.n5898 VSS 0.009191f
C24229 VDD.n5899 VSS 0.261039f
C24230 VDD.n5900 VSS 0.14099f
C24231 VDD.n5901 VSS 0.107577f
C24232 VDD.n5902 VSS 0.150746f
C24233 VDD.n5904 VSS 0.018625f
C24234 VDD.n5905 VSS 1.2e-19
C24235 VDD.n5906 VSS 0.0149f
C24236 VDD.n5907 VSS 0.222007f
C24237 VDD.n5908 VSS 0.01487f
C24238 VDD.n5910 VSS 0.018249f
C24239 VDD.n5911 VSS 0.009312f
C24240 VDD.n5912 VSS 2.44316f
C24241 VDD.n5913 VSS 0.009688f
C24242 VDD.n5914 VSS 0.030573f
C24243 VDD.t1646 VSS 0.066856f
C24244 VDD.n5916 VSS 0.129831f
C24245 VDD.t3099 VSS 0.016021f
C24246 VDD.t1637 VSS 0.066856f
C24247 VDD.n5917 VSS 0.129831f
C24248 VDD.t765 VSS 0.025104f
C24249 VDD.t4024 VSS 0.066856f
C24250 VDD.n5918 VSS 0.129831f
C24251 VDD.t3675 VSS 0.016021f
C24252 VDD.t1338 VSS 0.066856f
C24253 VDD.n5919 VSS 0.129831f
C24254 VDD.t1864 VSS 0.066856f
C24255 VDD.n5920 VSS 0.129831f
C24256 VDD.t3722 VSS 0.016021f
C24257 VDD.t2418 VSS 0.066856f
C24258 VDD.n5921 VSS 0.129831f
C24259 VDD.t2011 VSS 0.025104f
C24260 VDD.t1529 VSS 0.066856f
C24261 VDD.n5922 VSS 0.129831f
C24262 VDD.t3414 VSS 0.016021f
C24263 VDD.t2029 VSS 0.066856f
C24264 VDD.n5923 VSS 0.129831f
C24265 VDD.t2175 VSS 0.025104f
C24266 VDD.t1245 VSS 0.066856f
C24267 VDD.n5924 VSS 0.129831f
C24268 VDD.n5925 VSS 0.016021f
C24269 VDD.t1246 VSS 0.025104f
C24270 VDD.n5926 VSS 0.110991f
C24271 VDD.n5927 VSS 0.110991f
C24272 VDD.t2174 VSS 0.066856f
C24273 VDD.n5928 VSS 0.129831f
C24274 VDD.n5929 VSS 0.105899f
C24275 VDD.n5930 VSS 0.016021f
C24276 VDD.t2030 VSS 0.016021f
C24277 VDD.n5931 VSS 0.016021f
C24278 VDD.n5932 VSS 0.105899f
C24279 VDD.t3413 VSS 0.066856f
C24280 VDD.n5933 VSS 0.129831f
C24281 VDD.n5934 VSS 0.105899f
C24282 VDD.n5935 VSS 0.016021f
C24283 VDD.t1530 VSS 0.025104f
C24284 VDD.n5936 VSS 0.114533f
C24285 VDD.t1501 VSS 0.066856f
C24286 VDD.t4690 VSS 0.066856f
C24287 VDD.n5937 VSS 0.58882f
C24288 VDD.t2216 VSS 0.034186f
C24289 VDD.t3239 VSS 0.034186f
C24290 VDD.n5938 VSS 0.571765f
C24291 VDD.t3238 VSS 0.066856f
C24292 VDD.t2215 VSS 0.066856f
C24293 VDD.n5939 VSS 0.333277f
C24294 VDD.t2898 VSS 0.066856f
C24295 VDD.t1803 VSS 0.066856f
C24296 VDD.n5940 VSS 0.333277f
C24297 VDD.t1804 VSS 0.034186f
C24298 VDD.t2899 VSS 0.034186f
C24299 VDD.n5941 VSS 0.402094f
C24300 VDD.n5942 VSS 0.283088f
C24301 VDD.n5943 VSS 0.532659f
C24302 VDD.t1857 VSS 0.034186f
C24303 VDD.t2953 VSS 0.034186f
C24304 VDD.n5944 VSS 0.43943f
C24305 VDD.t2952 VSS 0.066856f
C24306 VDD.t1856 VSS 0.066856f
C24307 VDD.n5945 VSS 0.333277f
C24308 VDD.t2585 VSS 0.066856f
C24309 VDD.t1486 VSS 0.066856f
C24310 VDD.n5946 VSS 0.333277f
C24311 VDD.t1487 VSS 0.034186f
C24312 VDD.t2586 VSS 0.034186f
C24313 VDD.n5947 VSS 0.571765f
C24314 VDD.t4352 VSS 0.066856f
C24315 VDD.t3381 VSS 0.066856f
C24316 VDD.n5948 VSS 0.58882f
C24317 VDD.t3382 VSS 0.034186f
C24318 VDD.t4353 VSS 0.034186f
C24319 VDD.n5949 VSS 0.177249f
C24320 VDD.n5950 VSS 0.454987f
C24321 VDD.n5951 VSS 0.114533f
C24322 VDD.t2010 VSS 0.066856f
C24323 VDD.n5952 VSS 0.129831f
C24324 VDD.n5953 VSS 0.105899f
C24325 VDD.n5954 VSS 0.016021f
C24326 VDD.t2419 VSS 0.016021f
C24327 VDD.n5955 VSS 0.016021f
C24328 VDD.n5956 VSS 0.105899f
C24329 VDD.t3721 VSS 0.066856f
C24330 VDD.n5957 VSS 0.129831f
C24331 VDD.n5958 VSS 0.105899f
C24332 VDD.n5959 VSS 0.016021f
C24333 VDD.t1865 VSS 0.025104f
C24334 VDD.n5960 VSS 0.110991f
C24335 VDD.n5961 VSS 0.110991f
C24336 VDD.t1339 VSS 0.025104f
C24337 VDD.n5962 VSS 0.016021f
C24338 VDD.n5963 VSS 0.105899f
C24339 VDD.t3674 VSS 0.066856f
C24340 VDD.n5964 VSS 0.082848f
C24341 VDD.n5965 VSS 0.052949f
C24342 VDD.n5966 VSS 0.099933f
C24343 VDD.n5967 VSS 0.016021f
C24344 VDD.t4025 VSS 0.025104f
C24345 VDD.n5968 VSS 0.110991f
C24346 VDD.n5969 VSS 0.110991f
C24347 VDD.t764 VSS 0.066856f
C24348 VDD.n5970 VSS 0.129831f
C24349 VDD.n5971 VSS 0.105899f
C24350 VDD.n5972 VSS 0.016021f
C24351 VDD.t1638 VSS 0.016021f
C24352 VDD.n5973 VSS 0.016021f
C24353 VDD.n5974 VSS 0.105899f
C24354 VDD.t3098 VSS 0.066856f
C24355 VDD.n5975 VSS 0.129831f
C24356 VDD.n5976 VSS 0.105899f
C24357 VDD.n5977 VSS 0.016021f
C24358 VDD.t1647 VSS 0.025104f
C24359 VDD.n5978 VSS 0.114533f
C24360 VDD.t1951 VSS 0.034186f
C24361 VDD.n5979 VSS 0.031606f
C24362 VDD.n5980 VSS 0.080796f
C24363 VDD.n5981 VSS 0.01487f
C24364 VDD.n5983 VSS 0.018625f
C24365 VDD.t790 VSS 0.034186f
C24366 VDD.n5984 VSS 0.346215f
C24367 VDD.t789 VSS 0.066856f
C24368 VDD.n5985 VSS 0.203709f
C24369 VDD.t4536 VSS 0.066856f
C24370 VDD.n5986 VSS 0.203709f
C24371 VDD.t4537 VSS 0.034186f
C24372 VDD.n5987 VSS 0.249272f
C24373 VDD.t405 VSS 9.428519f
C24374 VDD.t393 VSS 7.61793f
C24375 VDD.t415 VSS 7.61793f
C24376 VDD.t392 VSS 9.81076f
C24377 VDD.t590 VSS 9.19382f
C24378 VDD.n5988 VSS 0.049953f
C24379 VDD.t2667 VSS 0.066856f
C24380 VDD.t2668 VSS 0.034186f
C24381 VDD.t2341 VSS 0.025104f
C24382 VDD.t2340 VSS 0.066856f
C24383 VDD.t4368 VSS 0.066856f
C24384 VDD.n5989 VSS 0.256005f
C24385 VDD.t1568 VSS 0.016021f
C24386 VDD.n5990 VSS 0.016021f
C24387 VDD.t3640 VSS 0.066856f
C24388 VDD.t3641 VSS 0.016021f
C24389 VDD.n5991 VSS 0.016021f
C24390 VDD.t2330 VSS 0.066856f
C24391 VDD.t4362 VSS 0.066856f
C24392 VDD.n5992 VSS 0.256005f
C24393 VDD.t3483 VSS 0.025104f
C24394 VDD.t2331 VSS 0.016021f
C24395 VDD.n5993 VSS 0.016021f
C24396 VDD.t1345 VSS 0.066856f
C24397 VDD.t1346 VSS 0.025104f
C24398 VDD.t4297 VSS 0.016021f
C24399 VDD.n5994 VSS 0.016021f
C24400 VDD.t4615 VSS 0.025104f
C24401 VDD.t4614 VSS 0.066856f
C24402 VDD.t2661 VSS 0.066856f
C24403 VDD.n5995 VSS 0.256005f
C24404 VDD.n5996 VSS 0.016021f
C24405 VDD.t2662 VSS 0.025104f
C24406 VDD.n5997 VSS 0.218415f
C24407 VDD.n5998 VSS 0.218415f
C24408 VDD.t3482 VSS 0.066856f
C24409 VDD.n5999 VSS 0.256005f
C24410 VDD.n6000 VSS 0.208141f
C24411 VDD.n6001 VSS 0.016021f
C24412 VDD.t4363 VSS 0.016021f
C24413 VDD.n6002 VSS 0.016021f
C24414 VDD.n6003 VSS 0.208141f
C24415 VDD.t1567 VSS 0.066856f
C24416 VDD.n6004 VSS 0.256005f
C24417 VDD.n6005 VSS 0.208141f
C24418 VDD.n6006 VSS 0.016021f
C24419 VDD.t4369 VSS 0.025104f
C24420 VDD.n6007 VSS 0.239302f
C24421 VDD.n6008 VSS 0.38869f
C24422 VDD.t4673 VSS 0.034186f
C24423 VDD.n6009 VSS 0.239302f
C24424 VDD.t4672 VSS 0.066856f
C24425 VDD.n6010 VSS 0.234752f
C24426 VDD.n6011 VSS 0.018249f
C24427 VDD.n6012 VSS 0.018625f
C24428 VDD.n6013 VSS 1.84672f
C24429 VDD.n6014 VSS 0.643547f
C24430 VDD.n6015 VSS 0.009688f
C24431 VDD.n6016 VSS 1.2e-19
C24432 VDD.t778 VSS 0.066856f
C24433 VDD.n6018 VSS 0.111632f
C24434 VDD.t2136 VSS 0.016021f
C24435 VDD.n6019 VSS 0.309204f
C24436 VDD.t4886 VSS 0.061518f
C24437 VDD.t4859 VSS 0.008011f
C24438 VDD.t4810 VSS 0.008011f
C24439 VDD.n6020 VSS 0.032022f
C24440 VDD.n6021 VSS 0.216759f
C24441 VDD.t649 VSS 0.066856f
C24442 VDD.n6022 VSS 0.111632f
C24443 VDD.t2583 VSS 0.066856f
C24444 VDD.n6023 VSS 0.126716f
C24445 VDD.n6024 VSS 0.111391f
C24446 VDD.t650 VSS 0.025104f
C24447 VDD.t1122 VSS 0.016021f
C24448 VDD.t1233 VSS 0.066856f
C24449 VDD.n6025 VSS 0.126716f
C24450 VDD.t4500 VSS 0.066856f
C24451 VDD.n6026 VSS 0.126716f
C24452 VDD.n6027 VSS 0.016021f
C24453 VDD.t4501 VSS 0.025104f
C24454 VDD.n6028 VSS 0.107953f
C24455 VDD.n6029 VSS 0.107953f
C24456 VDD.t1234 VSS 0.025104f
C24457 VDD.n6030 VSS 0.016021f
C24458 VDD.n6031 VSS 0.102784f
C24459 VDD.t1121 VSS 0.066856f
C24460 VDD.n6032 VSS 0.126716f
C24461 VDD.n6033 VSS 0.102784f
C24462 VDD.n6034 VSS 0.016021f
C24463 VDD.t2584 VSS 0.016021f
C24464 VDD.n6035 VSS 0.016021f
C24465 VDD.n6036 VSS 0.087513f
C24466 VDD.n6037 VSS 0.050646f
C24467 VDD.n6038 VSS 0.339165f
C24468 VDD.n6039 VSS 0.00473f
C24469 VDD.n6040 VSS 0.00473f
C24470 VDD.n6041 VSS 0.096376f
C24471 VDD.t4843 VSS 0.008011f
C24472 VDD.t4976 VSS 0.008011f
C24473 VDD.n6042 VSS 0.024025f
C24474 VDD.t4950 VSS 0.008011f
C24475 VDD.t4889 VSS 0.008011f
C24476 VDD.n6043 VSS 0.018621f
C24477 VDD.n6044 VSS 0.077103f
C24478 VDD.t4967 VSS 0.008011f
C24479 VDD.t4890 VSS 0.008011f
C24480 VDD.n6045 VSS 0.024025f
C24481 VDD.t4885 VSS 0.008011f
C24482 VDD.t4815 VSS 0.008011f
C24483 VDD.n6046 VSS 0.018621f
C24484 VDD.n6047 VSS 0.055299f
C24485 VDD.n6048 VSS 0.111411f
C24486 VDD.t4959 VSS 0.008011f
C24487 VDD.t4965 VSS 0.008011f
C24488 VDD.n6049 VSS 0.024025f
C24489 VDD.t4873 VSS 0.008011f
C24490 VDD.t4879 VSS 0.008011f
C24491 VDD.n6050 VSS 0.018621f
C24492 VDD.n6051 VSS 0.055299f
C24493 VDD.n6052 VSS 0.086287f
C24494 VDD.t4935 VSS 0.008011f
C24495 VDD.t4831 VSS 0.008011f
C24496 VDD.n6053 VSS 0.024025f
C24497 VDD.t4847 VSS 0.008011f
C24498 VDD.t4934 VSS 0.008011f
C24499 VDD.n6054 VSS 0.018621f
C24500 VDD.n6055 VSS 0.055299f
C24501 VDD.n6056 VSS 0.022927f
C24502 VDD.n6057 VSS 0.00473f
C24503 VDD.n6058 VSS 0.00473f
C24504 VDD.t4946 VSS 0.020865f
C24505 VDD.n6059 VSS 0.028664f
C24506 VDD.n6060 VSS 0.010511f
C24507 VDD.n6061 VSS 0.019257f
C24508 VDD.n6062 VSS 0.019243f
C24509 VDD.t4930 VSS 0.008011f
C24510 VDD.t4826 VSS 0.008011f
C24511 VDD.n6063 VSS 0.020046f
C24512 VDD.n6064 VSS 0.020708f
C24513 VDD.n6065 VSS 0.010511f
C24514 VDD.n6066 VSS 0.111886f
C24515 VDD.n6067 VSS 0.00473f
C24516 VDD.t4825 VSS 0.020865f
C24517 VDD.n6068 VSS 0.028664f
C24518 VDD.t4948 VSS 0.008011f
C24519 VDD.t4839 VSS 0.008011f
C24520 VDD.n6069 VSS 0.069277f
C24521 VDD.n6070 VSS 0.149006f
C24522 VDD.n6071 VSS 0.010511f
C24523 VDD.n6072 VSS 0.040406f
C24524 VDD.n6073 VSS 0.212121f
C24525 VDD.n6074 VSS 0.472695f
C24526 VDD.n6075 VSS 0.067373f
C24527 VDD.t4972 VSS 0.008011f
C24528 VDD.t4956 VSS 0.008011f
C24529 VDD.n6076 VSS 0.024025f
C24530 VDD.t4888 VSS 0.008011f
C24531 VDD.t4871 VSS 0.008011f
C24532 VDD.n6077 VSS 0.018621f
C24533 VDD.n6078 VSS 0.055299f
C24534 VDD.n6079 VSS 0.085099f
C24535 VDD.t4951 VSS 0.008011f
C24536 VDD.t4842 VSS 0.008011f
C24537 VDD.n6080 VSS 0.024025f
C24538 VDD.t4865 VSS 0.008011f
C24539 VDD.t4949 VSS 0.008011f
C24540 VDD.n6081 VSS 0.018621f
C24541 VDD.n6082 VSS 0.055299f
C24542 VDD.n6083 VSS 0.086289f
C24543 VDD.t4938 VSS 0.008011f
C24544 VDD.t4903 VSS 0.008011f
C24545 VDD.n6084 VSS 0.024025f
C24546 VDD.t4850 VSS 0.008011f
C24547 VDD.t4820 VSS 0.008011f
C24548 VDD.n6085 VSS 0.018621f
C24549 VDD.n6086 VSS 0.055299f
C24550 VDD.n6087 VSS 0.086287f
C24551 VDD.t4940 VSS 0.008011f
C24552 VDD.t4821 VSS 0.008011f
C24553 VDD.n6088 VSS 0.024025f
C24554 VDD.t4851 VSS 0.008011f
C24555 VDD.t4919 VSS 0.008011f
C24556 VDD.n6089 VSS 0.018621f
C24557 VDD.n6090 VSS 0.055299f
C24558 VDD.n6091 VSS 0.047999f
C24559 VDD.n6092 VSS 0.535333f
C24560 VDD.t4962 VSS 0.061518f
C24561 VDD.t4937 VSS 0.008011f
C24562 VDD.t4878 VSS 0.008011f
C24563 VDD.n6093 VSS 0.032022f
C24564 VDD.n6094 VSS 0.216759f
C24565 VDD.n6095 VSS 0.152023f
C24566 VDD.t4944 VSS 0.031728f
C24567 VDD.n6096 VSS 0.151284f
C24568 VDD.t4876 VSS 0.008011f
C24569 VDD.t4857 VSS 0.008011f
C24570 VDD.n6097 VSS 0.032022f
C24571 VDD.n6098 VSS 0.116906f
C24572 VDD.n6099 VSS 0.388663f
C24573 VDD.n6100 VSS 0.334665f
C24574 VDD.n6101 VSS 0.061022f
C24575 VDD.t4817 VSS 0.020865f
C24576 VDD.n6102 VSS 0.028664f
C24577 VDD.n6103 VSS 0.010511f
C24578 VDD.n6104 VSS 0.019257f
C24579 VDD.n6105 VSS 0.019243f
C24580 VDD.t4982 VSS 0.008011f
C24581 VDD.t4884 VSS 0.008011f
C24582 VDD.n6106 VSS 0.020046f
C24583 VDD.n6107 VSS 0.020708f
C24584 VDD.n6108 VSS 0.010511f
C24585 VDD.n6109 VSS 0.111886f
C24586 VDD.n6110 VSS 0.00473f
C24587 VDD.t4877 VSS 0.020865f
C24588 VDD.n6111 VSS 0.028664f
C24589 VDD.t4819 VSS 0.008011f
C24590 VDD.t4902 VSS 0.008011f
C24591 VDD.n6112 VSS 0.069277f
C24592 VDD.n6113 VSS 0.149006f
C24593 VDD.n6114 VSS 0.010511f
C24594 VDD.n6115 VSS 0.040406f
C24595 VDD.n6116 VSS 0.147417f
C24596 VDD.n6117 VSS 0.303879f
C24597 VDD.t4863 VSS 0.008011f
C24598 VDD.t4925 VSS 0.008011f
C24599 VDD.n6118 VSS 0.024025f
C24600 VDD.t4912 VSS 0.008011f
C24601 VDD.t4971 VSS 0.008011f
C24602 VDD.n6119 VSS 0.018621f
C24603 VDD.n6120 VSS 0.055299f
C24604 VDD.n6121 VSS 0.047999f
C24605 VDD.t4861 VSS 0.008011f
C24606 VDD.t4824 VSS 0.008011f
C24607 VDD.n6122 VSS 0.024025f
C24608 VDD.t4911 VSS 0.008011f
C24609 VDD.t4869 VSS 0.008011f
C24610 VDD.n6123 VSS 0.018621f
C24611 VDD.n6124 VSS 0.055299f
C24612 VDD.n6125 VSS 0.086287f
C24613 VDD.t4874 VSS 0.008011f
C24614 VDD.t4955 VSS 0.008011f
C24615 VDD.n6126 VSS 0.024025f
C24616 VDD.t4921 VSS 0.008011f
C24617 VDD.t4822 VSS 0.008011f
C24618 VDD.n6127 VSS 0.018621f
C24619 VDD.n6128 VSS 0.055299f
C24620 VDD.n6129 VSS 0.086289f
C24621 VDD.t4897 VSS 0.008011f
C24622 VDD.t4880 VSS 0.008011f
C24623 VDD.n6130 VSS 0.024025f
C24624 VDD.t4939 VSS 0.008011f
C24625 VDD.t4926 VSS 0.008011f
C24626 VDD.n6131 VSS 0.018621f
C24627 VDD.n6132 VSS 0.055299f
C24628 VDD.n6133 VSS 0.085099f
C24629 VDD.t4960 VSS 0.008011f
C24630 VDD.t4899 VSS 0.008011f
C24631 VDD.n6134 VSS 0.024025f
C24632 VDD.t4823 VSS 0.008011f
C24633 VDD.t4943 VSS 0.008011f
C24634 VDD.n6135 VSS 0.018621f
C24635 VDD.n6136 VSS 0.077103f
C24636 VDD.t4893 VSS 0.008011f
C24637 VDD.t4816 VSS 0.008011f
C24638 VDD.n6137 VSS 0.024025f
C24639 VDD.t4936 VSS 0.008011f
C24640 VDD.t4853 VSS 0.008011f
C24641 VDD.n6138 VSS 0.018621f
C24642 VDD.n6139 VSS 0.055299f
C24643 VDD.n6140 VSS 0.111411f
C24644 VDD.t4883 VSS 0.008011f
C24645 VDD.t4887 VSS 0.008011f
C24646 VDD.n6141 VSS 0.024025f
C24647 VDD.t4928 VSS 0.008011f
C24648 VDD.t4932 VSS 0.008011f
C24649 VDD.n6142 VSS 0.018621f
C24650 VDD.n6143 VSS 0.055299f
C24651 VDD.n6144 VSS 0.086287f
C24652 VDD.t4854 VSS 0.008011f
C24653 VDD.t4942 VSS 0.008011f
C24654 VDD.n6145 VSS 0.024025f
C24655 VDD.t4908 VSS 0.008011f
C24656 VDD.t4813 VSS 0.008011f
C24657 VDD.n6146 VSS 0.018621f
C24658 VDD.n6147 VSS 0.055299f
C24659 VDD.n6148 VSS 0.022927f
C24660 VDD.n6149 VSS 0.067373f
C24661 VDD.n6150 VSS 0.306702f
C24662 VDD.n6151 VSS 0.27523f
C24663 VDD.n6152 VSS 0.152023f
C24664 VDD.t4866 VSS 0.031728f
C24665 VDD.n6153 VSS 0.151284f
C24666 VDD.t4983 VSS 0.008011f
C24667 VDD.t4969 VSS 0.008011f
C24668 VDD.n6154 VSS 0.032022f
C24669 VDD.n6155 VSS 0.116906f
C24670 VDD.n6156 VSS 0.324728f
C24671 VDD.n6157 VSS 0.050646f
C24672 VDD.t770 VSS 0.066856f
C24673 VDD.n6158 VSS 0.126716f
C24674 VDD.t4015 VSS 0.025104f
C24675 VDD.t3170 VSS 0.066856f
C24676 VDD.n6159 VSS 0.126716f
C24677 VDD.n6160 VSS 0.016021f
C24678 VDD.t3171 VSS 0.025104f
C24679 VDD.n6161 VSS 0.107953f
C24680 VDD.n6162 VSS 0.107953f
C24681 VDD.t4014 VSS 0.066856f
C24682 VDD.n6163 VSS 0.126716f
C24683 VDD.n6164 VSS 0.102784f
C24684 VDD.n6165 VSS 0.016021f
C24685 VDD.t771 VSS 0.016021f
C24686 VDD.n6166 VSS 0.016021f
C24687 VDD.n6167 VSS 0.102784f
C24688 VDD.t2135 VSS 0.066856f
C24689 VDD.n6168 VSS 0.126716f
C24690 VDD.n6169 VSS 0.087513f
C24691 VDD.n6170 VSS 0.016021f
C24692 VDD.t779 VSS 0.025104f
C24693 VDD.n6171 VSS 0.111391f
C24694 VDD.n6172 VSS 0.0149f
C24695 VDD.n6173 VSS 0.182651f
C24696 VDD.n6174 VSS 0.079472f
C24697 VDD.t1068 VSS 0.034186f
C24698 VDD.n6175 VSS 0.028209f
C24699 VDD.n6177 VSS 0.030311f
C24700 VDD.n6178 VSS 0.01487f
C24701 VDD.n6179 VSS 0.076301f
C24702 VDD.t1067 VSS 0.066856f
C24703 VDD.n6180 VSS 0.334361f
C24704 VDD.t2798 VSS 0.034186f
C24705 VDD.n6181 VSS 0.356145f
C24706 VDD.t2797 VSS 0.066856f
C24707 VDD.n6182 VSS 0.203709f
C24708 VDD.t2420 VSS 0.066856f
C24709 VDD.n6183 VSS 0.203709f
C24710 VDD.t2421 VSS 0.034186f
C24711 VDD.n6184 VSS 0.249272f
C24712 VDD.n6185 VSS 0.335514f
C24713 VDD.t3406 VSS 0.034186f
C24714 VDD.n6186 VSS 0.272789f
C24715 VDD.t3405 VSS 0.066856f
C24716 VDD.n6187 VSS 0.203709f
C24717 VDD.t3092 VSS 0.066856f
C24718 VDD.n6188 VSS 0.203709f
C24719 VDD.t3093 VSS 0.034186f
C24720 VDD.n6189 VSS 0.346215f
C24721 VDD.n6190 VSS 0.610826f
C24722 VDD.t4421 VSS 0.034186f
C24723 VDD.n6191 VSS 0.346215f
C24724 VDD.t4420 VSS 0.066856f
C24725 VDD.n6192 VSS 0.203709f
C24726 VDD.t4086 VSS 0.066856f
C24727 VDD.n6193 VSS 0.203709f
C24728 VDD.t4087 VSS 0.034186f
C24729 VDD.n6194 VSS 0.249272f
C24730 VDD.n6195 VSS 0.335514f
C24731 VDD.t2210 VSS 0.034186f
C24732 VDD.n6196 VSS 0.272789f
C24733 VDD.t2209 VSS 0.066856f
C24734 VDD.n6197 VSS 0.203709f
C24735 VDD.t1793 VSS 0.066856f
C24736 VDD.n6198 VSS 0.203709f
C24737 VDD.t1794 VSS 0.034186f
C24738 VDD.n6199 VSS 0.346215f
C24739 VDD.t3502 VSS 0.066856f
C24740 VDD.t3492 VSS 0.066856f
C24741 VDD.n6200 VSS 0.377014f
C24742 VDD.t3503 VSS 0.034186f
C24743 VDD.t3249 VSS 0.025104f
C24744 VDD.t3248 VSS 0.066856f
C24745 VDD.t3234 VSS 0.066856f
C24746 VDD.n6201 VSS 0.414447f
C24747 VDD.t4521 VSS 0.016021f
C24748 VDD.n6202 VSS 0.016021f
C24749 VDD.t4526 VSS 0.066856f
C24750 VDD.t4527 VSS 0.016021f
C24751 VDD.n6203 VSS 0.016021f
C24752 VDD.t3242 VSS 0.066856f
C24753 VDD.t3228 VSS 0.066856f
C24754 VDD.n6204 VSS 0.414447f
C24755 VDD.t2312 VSS 0.025104f
C24756 VDD.t3243 VSS 0.016021f
C24757 VDD.n6205 VSS 0.016021f
C24758 VDD.t2334 VSS 0.066856f
C24759 VDD.t2335 VSS 0.025104f
C24760 VDD.t1366 VSS 0.025104f
C24761 VDD.t1365 VSS 0.066856f
C24762 VDD.t1349 VSS 0.066856f
C24763 VDD.n6206 VSS 0.414447f
C24764 VDD.t1041 VSS 0.016021f
C24765 VDD.n6207 VSS 0.016021f
C24766 VDD.t1065 VSS 0.066856f
C24767 VDD.t1066 VSS 0.016021f
C24768 VDD.n6208 VSS 0.016021f
C24769 VDD.t2980 VSS 0.066856f
C24770 VDD.t2964 VSS 0.066856f
C24771 VDD.n6209 VSS 0.414447f
C24772 VDD.t2981 VSS 0.025104f
C24773 VDD.t3433 VSS 0.025104f
C24774 VDD.t3432 VSS 0.066856f
C24775 VDD.t3411 VSS 0.066856f
C24776 VDD.n6210 VSS 0.414447f
C24777 VDD.t1087 VSS 0.016021f
C24778 VDD.n6211 VSS 0.016021f
C24779 VDD.t1104 VSS 0.066856f
C24780 VDD.t1105 VSS 0.016021f
C24781 VDD.n6212 VSS 0.016021f
C24782 VDD.t3876 VSS 0.066856f
C24783 VDD.t3862 VSS 0.066856f
C24784 VDD.n6213 VSS 0.414447f
C24785 VDD.t3535 VSS 0.025104f
C24786 VDD.t3877 VSS 0.016021f
C24787 VDD.n6214 VSS 0.016021f
C24788 VDD.t3544 VSS 0.066856f
C24789 VDD.t3545 VSS 0.025104f
C24790 VDD.t1708 VSS 0.034186f
C24791 VDD.t1707 VSS 0.066856f
C24792 VDD.t1691 VSS 0.066856f
C24793 VDD.n6215 VSS 0.414447f
C24794 VDD.t4546 VSS 0.066856f
C24795 VDD.t3597 VSS 0.066856f
C24796 VDD.n6216 VSS 0.333277f
C24797 VDD.t4238 VSS 0.066856f
C24798 VDD.t3288 VSS 0.066856f
C24799 VDD.n6217 VSS 0.333277f
C24800 VDD.t3289 VSS 0.034186f
C24801 VDD.t4239 VSS 0.034186f
C24802 VDD.n6218 VSS 0.556001f
C24803 VDD.t763 VSS 0.034186f
C24804 VDD.t762 VSS 0.066856f
C24805 VDD.t736 VSS 0.066856f
C24806 VDD.n6219 VSS 0.414447f
C24807 VDD.t3157 VSS 0.025104f
C24808 VDD.t3156 VSS 0.066856f
C24809 VDD.t3142 VSS 0.066856f
C24810 VDD.n6220 VSS 0.414447f
C24811 VDD.t777 VSS 0.016021f
C24812 VDD.n6221 VSS 0.016021f
C24813 VDD.t787 VSS 0.066856f
C24814 VDD.t788 VSS 0.016021f
C24815 VDD.n6222 VSS 0.016021f
C24816 VDD.t3552 VSS 0.066856f
C24817 VDD.t3540 VSS 0.066856f
C24818 VDD.n6223 VSS 0.414447f
C24819 VDD.t3665 VSS 0.025104f
C24820 VDD.t3553 VSS 0.016021f
C24821 VDD.n6224 VSS 0.016021f
C24822 VDD.t3683 VSS 0.066856f
C24823 VDD.t3684 VSS 0.025104f
C24824 VDD.t2879 VSS 0.025104f
C24825 VDD.t2878 VSS 0.066856f
C24826 VDD.t2866 VSS 0.066856f
C24827 VDD.n6225 VSS 0.414447f
C24828 VDD.t1392 VSS 0.016021f
C24829 VDD.n6226 VSS 0.016021f
C24830 VDD.t1403 VSS 0.066856f
C24831 VDD.t1404 VSS 0.016021f
C24832 VDD.n6227 VSS 0.016021f
C24833 VDD.t3300 VSS 0.066856f
C24834 VDD.t3292 VSS 0.066856f
C24835 VDD.n6228 VSS 0.414447f
C24836 VDD.t3301 VSS 0.025104f
C24837 VDD.t3787 VSS 0.025104f
C24838 VDD.t3786 VSS 0.066856f
C24839 VDD.t3770 VSS 0.066856f
C24840 VDD.n6229 VSS 0.414447f
C24841 VDD.t2038 VSS 0.016021f
C24842 VDD.n6230 VSS 0.016021f
C24843 VDD.t2058 VSS 0.066856f
C24844 VDD.t2059 VSS 0.016021f
C24845 VDD.n6231 VSS 0.016021f
C24846 VDD.t1127 VSS 0.066856f
C24847 VDD.t1117 VSS 0.066856f
C24848 VDD.n6232 VSS 0.414447f
C24849 VDD.t3901 VSS 0.025104f
C24850 VDD.t1128 VSS 0.016021f
C24851 VDD.t3919 VSS 0.025104f
C24852 VDD.n6233 VSS 0.016021f
C24853 VDD.t3918 VSS 0.066856f
C24854 VDD.t3900 VSS 0.066856f
C24855 VDD.n6234 VSS 0.414447f
C24856 VDD.n6235 VSS 0.366582f
C24857 VDD.n6236 VSS 0.016021f
C24858 VDD.t1118 VSS 0.016021f
C24859 VDD.n6237 VSS 0.016021f
C24860 VDD.n6238 VSS 0.366582f
C24861 VDD.t2037 VSS 0.066856f
C24862 VDD.n6239 VSS 0.414447f
C24863 VDD.n6240 VSS 0.366582f
C24864 VDD.n6241 VSS 0.016021f
C24865 VDD.t3771 VSS 0.025104f
C24866 VDD.n6242 VSS 0.372952f
C24867 VDD.n6243 VSS 0.372952f
C24868 VDD.t3293 VSS 0.025104f
C24869 VDD.n6244 VSS 0.016021f
C24870 VDD.n6245 VSS 0.366582f
C24871 VDD.t1391 VSS 0.066856f
C24872 VDD.n6246 VSS 0.251808f
C24873 VDD.n6247 VSS 0.183291f
C24874 VDD.n6248 VSS 0.34593f
C24875 VDD.n6249 VSS 0.016021f
C24876 VDD.t2867 VSS 0.025104f
C24877 VDD.n6250 VSS 0.372952f
C24878 VDD.n6251 VSS 0.372952f
C24879 VDD.t3664 VSS 0.066856f
C24880 VDD.n6252 VSS 0.414447f
C24881 VDD.n6253 VSS 0.366582f
C24882 VDD.n6254 VSS 0.016021f
C24883 VDD.t3541 VSS 0.016021f
C24884 VDD.n6255 VSS 0.016021f
C24885 VDD.n6256 VSS 0.366582f
C24886 VDD.t776 VSS 0.066856f
C24887 VDD.n6257 VSS 0.414447f
C24888 VDD.n6258 VSS 0.366582f
C24889 VDD.n6259 VSS 0.016021f
C24890 VDD.t3143 VSS 0.025104f
C24891 VDD.n6260 VSS 0.409739f
C24892 VDD.n6261 VSS 0.409739f
C24893 VDD.t737 VSS 0.034186f
C24894 VDD.n6262 VSS 0.369079f
C24895 VDD.t2482 VSS 0.034186f
C24896 VDD.t3390 VSS 0.034186f
C24897 VDD.t3389 VSS 0.066856f
C24898 VDD.t3090 VSS 0.066856f
C24899 VDD.t2050 VSS 0.066856f
C24900 VDD.n6263 VSS 0.333277f
C24901 VDD.t2481 VSS 0.066856f
C24902 VDD.n6264 VSS 0.333277f
C24903 VDD.n6265 VSS 0.556001f
C24904 VDD.n6266 VSS 1.1439f
C24905 VDD.n6267 VSS 0.369079f
C24906 VDD.t1692 VSS 0.034186f
C24907 VDD.n6268 VSS 0.409739f
C24908 VDD.n6269 VSS 0.409739f
C24909 VDD.t3534 VSS 0.066856f
C24910 VDD.n6270 VSS 0.414447f
C24911 VDD.n6271 VSS 0.366582f
C24912 VDD.n6272 VSS 0.016021f
C24913 VDD.t3863 VSS 0.016021f
C24914 VDD.n6273 VSS 0.016021f
C24915 VDD.n6274 VSS 0.366582f
C24916 VDD.t1086 VSS 0.066856f
C24917 VDD.n6275 VSS 0.414447f
C24918 VDD.n6276 VSS 0.366582f
C24919 VDD.n6277 VSS 0.016021f
C24920 VDD.t3412 VSS 0.025104f
C24921 VDD.n6278 VSS 0.372952f
C24922 VDD.n6279 VSS 0.372952f
C24923 VDD.t2965 VSS 0.025104f
C24924 VDD.n6280 VSS 0.016021f
C24925 VDD.n6281 VSS 0.366582f
C24926 VDD.t1040 VSS 0.066856f
C24927 VDD.n6282 VSS 0.251808f
C24928 VDD.n6283 VSS 0.183291f
C24929 VDD.n6284 VSS 0.34593f
C24930 VDD.n6285 VSS 0.016021f
C24931 VDD.t1350 VSS 0.025104f
C24932 VDD.n6286 VSS 0.372952f
C24933 VDD.n6287 VSS 0.372952f
C24934 VDD.t2311 VSS 0.066856f
C24935 VDD.n6288 VSS 0.414447f
C24936 VDD.n6289 VSS 0.366582f
C24937 VDD.n6290 VSS 0.016021f
C24938 VDD.t3229 VSS 0.016021f
C24939 VDD.n6291 VSS 0.016021f
C24940 VDD.n6292 VSS 0.366582f
C24941 VDD.t4520 VSS 0.066856f
C24942 VDD.n6293 VSS 0.414447f
C24943 VDD.n6294 VSS 0.366582f
C24944 VDD.n6295 VSS 0.016021f
C24945 VDD.t3235 VSS 0.025104f
C24946 VDD.n6296 VSS 0.409739f
C24947 VDD.n6297 VSS 0.409739f
C24948 VDD.t3493 VSS 0.034186f
C24949 VDD.n6298 VSS 0.678315f
C24950 VDD.n6299 VSS 0.050127f
C24951 VDD.n6300 VSS 0.690048f
C24952 VDD.t1010 VSS 0.034186f
C24953 VDD.n6301 VSS 0.346215f
C24954 VDD.t1009 VSS 0.066856f
C24955 VDD.n6302 VSS 0.203709f
C24956 VDD.t589 VSS 0.066856f
C24957 VDD.n6303 VSS 0.203709f
C24958 VDD.t591 VSS 0.034186f
C24959 VDD.n6304 VSS 0.249272f
C24960 VDD.t899 VSS 0.034186f
C24961 VDD.t4653 VSS 0.034186f
C24962 VDD.n6305 VSS 0.346215f
C24963 VDD.t4652 VSS 0.066856f
C24964 VDD.n6306 VSS 0.203709f
C24965 VDD.t898 VSS 0.066856f
C24966 VDD.n6307 VSS 0.203709f
C24967 VDD.n6308 VSS 0.272789f
C24968 VDD.n6309 VSS 0.335514f
C24969 VDD.n6310 VSS 0.280759f
C24970 VDD.n6311 VSS 4.50638f
C24971 VDD.n6312 VSS 0.280759f
C24972 VDD.n6313 VSS 0.335514f
C24973 VDD.t4595 VSS 0.034186f
C24974 VDD.n6314 VSS 0.272789f
C24975 VDD.t4594 VSS 0.066856f
C24976 VDD.n6315 VSS 0.203709f
C24977 VDD.t4262 VSS 0.066856f
C24978 VDD.n6316 VSS 0.203709f
C24979 VDD.t4263 VSS 0.034186f
C24980 VDD.n6317 VSS 0.356145f
C24981 VDD.t1950 VSS 0.066856f
C24982 VDD.n6318 VSS 0.3341f
C24983 VDD.n6320 VSS 0.076039f
C24984 VDD.n6322 VSS 0.01502f
C24985 VDD.n6323 VSS 0.191797f
C24986 VDD.n6324 VSS 0.018249f
C24987 VDD.n6325 VSS 0.009312f
C24988 VDD.n6326 VSS 2.86995f
C24989 VDD.n6327 VSS 1.64177f
C24990 VDD.n6328 VSS 0.049886f
C24991 VDD.n6329 VSS 0.388695f
C24992 VDD.t4373 VSS 0.034186f
C24993 VDD.n6330 VSS 0.239302f
C24994 VDD.n6331 VSS 0.239302f
C24995 VDD.t3057 VSS 0.025104f
C24996 VDD.n6332 VSS 0.016021f
C24997 VDD.n6333 VSS 0.208141f
C24998 VDD.n6334 VSS 0.016021f
C24999 VDD.t1275 VSS 0.016021f
C25000 VDD.n6335 VSS 0.016021f
C25001 VDD.n6336 VSS 0.208141f
C25002 VDD.n6337 VSS 0.016021f
C25003 VDD.t3053 VSS 0.016021f
C25004 VDD.n6338 VSS 0.016021f
C25005 VDD.n6339 VSS 0.208141f
C25006 VDD.n6340 VSS 0.016021f
C25007 VDD.t3231 VSS 0.025104f
C25008 VDD.n6341 VSS 0.218415f
C25009 VDD.n6342 VSS 0.218415f
C25010 VDD.t2337 VSS 0.025104f
C25011 VDD.n6343 VSS 0.016021f
C25012 VDD.n6344 VSS 0.196415f
C25013 VDD.n6345 VSS 0.016021f
C25014 VDD.t876 VSS 0.016021f
C25015 VDD.n6346 VSS 0.016021f
C25016 VDD.n6347 VSS 0.208141f
C25017 VDD.n6348 VSS 0.016021f
C25018 VDD.t3789 VSS 0.025104f
C25019 VDD.n6349 VSS 0.218415f
C25020 VDD.n6350 VSS 0.218415f
C25021 VDD.t3265 VSS 0.025104f
C25022 VDD.n6351 VSS 0.016021f
C25023 VDD.n6352 VSS 0.208141f
C25024 VDD.n6353 VSS 0.016021f
C25025 VDD.t1988 VSS 0.016021f
C25026 VDD.n6354 VSS 0.016021f
C25027 VDD.n6355 VSS 0.208141f
C25028 VDD.n6356 VSS 0.016021f
C25029 VDD.t3661 VSS 0.016021f
C25030 VDD.n6357 VSS 0.016021f
C25031 VDD.n6358 VSS 0.208141f
C25032 VDD.n6359 VSS 0.016021f
C25033 VDD.t4419 VSS 0.025104f
C25034 VDD.n6360 VSS 0.225377f
C25035 VDD.n6361 VSS 0.570644f
C25036 VDD.n6362 VSS 0.33406f
C25037 VDD.t1623 VSS 0.066856f
C25038 VDD.n6363 VSS 0.58882f
C25039 VDD.n6364 VSS 0.571765f
C25040 VDD.t1910 VSS 0.066856f
C25041 VDD.n6365 VSS 0.333277f
C25042 VDD.t2344 VSS 0.066856f
C25043 VDD.n6366 VSS 0.333277f
C25044 VDD.n6367 VSS 0.43943f
C25045 VDD.n6368 VSS 0.532659f
C25046 VDD.n6369 VSS 0.280759f
C25047 VDD.n6370 VSS 4.15767f
C25048 VDD.n6371 VSS 0.280759f
C25049 VDD.n6372 VSS 0.532659f
C25050 VDD.n6373 VSS 0.402094f
C25051 VDD.t1308 VSS 0.066856f
C25052 VDD.n6374 VSS 0.333277f
C25053 VDD.t1673 VSS 0.066856f
C25054 VDD.n6375 VSS 0.333277f
C25055 VDD.n6376 VSS 0.571765f
C25056 VDD.t4006 VSS 0.066856f
C25057 VDD.n6377 VSS 0.58882f
C25058 VDD.n6378 VSS 0.333645f
C25059 VDD.n6379 VSS 0.570644f
C25060 VDD.n6380 VSS 0.225377f
C25061 VDD.t4720 VSS 0.066856f
C25062 VDD.n6381 VSS 0.256005f
C25063 VDD.n6382 VSS 0.208141f
C25064 VDD.n6383 VSS 0.016021f
C25065 VDD.t931 VSS 0.016021f
C25066 VDD.n6384 VSS 0.016021f
C25067 VDD.n6385 VSS 0.208141f
C25068 VDD.t2342 VSS 0.066856f
C25069 VDD.n6386 VSS 0.256005f
C25070 VDD.n6387 VSS 0.208141f
C25071 VDD.n6388 VSS 0.016021f
C25072 VDD.t4571 VSS 0.025104f
C25073 VDD.n6389 VSS 0.218415f
C25074 VDD.n6390 VSS 0.218415f
C25075 VDD.t4095 VSS 0.025104f
C25076 VDD.n6391 VSS 0.016021f
C25077 VDD.n6392 VSS 0.208141f
C25078 VDD.t2272 VSS 0.066856f
C25079 VDD.n6393 VSS 0.163661f
C25080 VDD.n6394 VSS 0.10407f
C25081 VDD.n6395 VSS 0.279865f
C25082 VDD.n6396 VSS 3.80896f
C25083 VDD.n6397 VSS 0.279865f
C25084 VDD.n6398 VSS 0.051392f
C25085 VDD.t2860 VSS 0.066856f
C25086 VDD.n6399 VSS 0.081115f
C25087 VDD.n6400 VSS 0.102784f
C25088 VDD.n6401 VSS 0.016021f
C25089 VDD.t4597 VSS 0.025104f
C25090 VDD.n6402 VSS 0.107953f
C25091 VDD.n6403 VSS 0.107953f
C25092 VDD.t1005 VSS 0.066856f
C25093 VDD.n6404 VSS 0.126716f
C25094 VDD.n6405 VSS 0.102784f
C25095 VDD.n6406 VSS 0.016021f
C25096 VDD.t2901 VSS 0.016021f
C25097 VDD.n6407 VSS 0.016021f
C25098 VDD.n6408 VSS 0.102784f
C25099 VDD.t1419 VSS 0.066856f
C25100 VDD.n6409 VSS 0.126716f
C25101 VDD.n6410 VSS 0.084772f
C25102 VDD.n6411 VSS 0.016021f
C25103 VDD.t1111 VSS 0.025104f
C25104 VDD.n6412 VSS 0.105419f
C25105 VDD.n6413 VSS 0.05157f
C25106 VDD.n6414 VSS 0.041023f
C25107 VDD.n6415 VSS 0.339165f
C25108 VDD.n6416 VSS 0.00473f
C25109 VDD.n6417 VSS 0.00473f
C25110 VDD.n6418 VSS 0.00473f
C25111 VDD.t4896 VSS 0.008011f
C25112 VDD.t4954 VSS 0.008011f
C25113 VDD.n6419 VSS 0.042109f
C25114 VDD.n6420 VSS 0.063057f
C25115 VDD.t4895 VSS 0.008011f
C25116 VDD.t4848 VSS 0.008011f
C25117 VDD.n6421 VSS 0.018495f
C25118 VDD.n6422 VSS 0.016425f
C25119 VDD.n6423 VSS 0.010511f
C25120 VDD.n6424 VSS 0.062181f
C25121 VDD.n6425 VSS 0.062177f
C25122 VDD.t4906 VSS 0.008011f
C25123 VDD.t4809 VSS 0.008011f
C25124 VDD.n6426 VSS 0.018495f
C25125 VDD.n6427 VSS 0.016425f
C25126 VDD.n6428 VSS 0.010511f
C25127 VDD.n6429 VSS 0.019381f
C25128 VDD.n6430 VSS 0.019376f
C25129 VDD.t4924 VSS 0.008011f
C25130 VDD.t4910 VSS 0.008011f
C25131 VDD.n6431 VSS 0.018495f
C25132 VDD.n6432 VSS 0.016425f
C25133 VDD.n6433 VSS 0.010511f
C25134 VDD.n6434 VSS 0.00416f
C25135 VDD.n6435 VSS 0.00473f
C25136 VDD.t4891 VSS 0.008011f
C25137 VDD.t4973 VSS 0.008011f
C25138 VDD.n6436 VSS 0.018495f
C25139 VDD.n6437 VSS 0.016425f
C25140 VDD.n6438 VSS 0.00473f
C25141 VDD.t4913 VSS 0.008011f
C25142 VDD.t4918 VSS 0.008011f
C25143 VDD.n6439 VSS 0.018495f
C25144 VDD.n6440 VSS 0.016425f
C25145 VDD.n6441 VSS 0.00473f
C25146 VDD.t4922 VSS 0.008011f
C25147 VDD.t4837 VSS 0.008011f
C25148 VDD.n6442 VSS 0.018495f
C25149 VDD.n6443 VSS 0.016425f
C25150 VDD.n6444 VSS 0.00473f
C25151 VDD.t4812 VSS 0.008011f
C25152 VDD.t4927 VSS 0.008011f
C25153 VDD.n6445 VSS 0.018495f
C25154 VDD.n6446 VSS 0.016425f
C25155 VDD.n6447 VSS 0.093664f
C25156 VDD.t4856 VSS 0.008011f
C25157 VDD.t4840 VSS 0.008011f
C25158 VDD.n6448 VSS 0.0221f
C25159 VDD.t4963 VSS 0.008011f
C25160 VDD.t4947 VSS 0.008011f
C25161 VDD.n6449 VSS 0.020181f
C25162 VDD.n6450 VSS 0.124159f
C25163 VDD.t4929 VSS 0.022609f
C25164 VDD.t4838 VSS 0.02098f
C25165 VDD.n6451 VSS 0.071904f
C25166 VDD.n6452 VSS 0.142473f
C25167 VDD.n6453 VSS 0.00473f
C25168 VDD.n6454 VSS 0.00473f
C25169 VDD.n6455 VSS 0.00473f
C25170 VDD.t4836 VSS 0.008011f
C25171 VDD.t4904 VSS 0.008011f
C25172 VDD.n6456 VSS 0.042109f
C25173 VDD.n6457 VSS 0.063057f
C25174 VDD.t4835 VSS 0.008011f
C25175 VDD.t4808 VSS 0.008011f
C25176 VDD.n6458 VSS 0.018495f
C25177 VDD.n6459 VSS 0.016425f
C25178 VDD.n6460 VSS 0.010511f
C25179 VDD.n6461 VSS 0.062181f
C25180 VDD.n6462 VSS 0.062177f
C25181 VDD.t4845 VSS 0.008011f
C25182 VDD.t4931 VSS 0.008011f
C25183 VDD.n6463 VSS 0.018495f
C25184 VDD.n6464 VSS 0.016425f
C25185 VDD.n6465 VSS 0.010511f
C25186 VDD.n6466 VSS 0.019381f
C25187 VDD.n6467 VSS 0.019376f
C25188 VDD.t4870 VSS 0.008011f
C25189 VDD.t4849 VSS 0.008011f
C25190 VDD.n6468 VSS 0.018495f
C25191 VDD.n6469 VSS 0.016425f
C25192 VDD.n6470 VSS 0.010511f
C25193 VDD.n6471 VSS 0.00416f
C25194 VDD.n6472 VSS 0.00473f
C25195 VDD.t4832 VSS 0.008011f
C25196 VDD.t4920 VSS 0.008011f
C25197 VDD.n6473 VSS 0.018495f
C25198 VDD.n6474 VSS 0.016425f
C25199 VDD.n6475 VSS 0.00473f
C25200 VDD.t4852 VSS 0.008011f
C25201 VDD.t4860 VSS 0.008011f
C25202 VDD.n6476 VSS 0.018495f
C25203 VDD.n6477 VSS 0.016425f
C25204 VDD.n6478 VSS 0.00473f
C25205 VDD.t4867 VSS 0.008011f
C25206 VDD.t4979 VSS 0.008011f
C25207 VDD.n6479 VSS 0.018495f
C25208 VDD.n6480 VSS 0.016425f
C25209 VDD.n6481 VSS 0.00473f
C25210 VDD.t4933 VSS 0.008011f
C25211 VDD.t4872 VSS 0.008011f
C25212 VDD.n6482 VSS 0.018495f
C25213 VDD.n6483 VSS 0.016425f
C25214 VDD.n6484 VSS 0.010511f
C25215 VDD.n6485 VSS 0.019376f
C25216 VDD.n6486 VSS 0.019381f
C25217 VDD.n6487 VSS 0.010511f
C25218 VDD.n6488 VSS 0.062177f
C25219 VDD.n6489 VSS 0.062181f
C25220 VDD.n6490 VSS 0.010511f
C25221 VDD.n6491 VSS 0.019376f
C25222 VDD.n6492 VSS 0.019381f
C25223 VDD.n6493 VSS 0.010511f
C25224 VDD.n6494 VSS 0.061871f
C25225 VDD.n6495 VSS 0.132226f
C25226 VDD.n6496 VSS 0.466322f
C25227 VDD.n6497 VSS 0.152036f
C25228 VDD.t4923 VSS 0.008011f
C25229 VDD.t4858 VSS 0.008011f
C25230 VDD.n6498 VSS 0.0221f
C25231 VDD.t4834 VSS 0.008011f
C25232 VDD.t4964 VSS 0.008011f
C25233 VDD.n6499 VSS 0.020181f
C25234 VDD.n6500 VSS 0.055665f
C25235 VDD.n6501 VSS 0.1321f
C25236 VDD.t4945 VSS 0.022609f
C25237 VDD.t4855 VSS 0.02098f
C25238 VDD.n6502 VSS 0.071904f
C25239 VDD.n6503 VSS 0.086055f
C25240 VDD.n6504 VSS 0.507601f
C25241 VDD.t4958 VSS 0.008011f
C25242 VDD.t4830 VSS 0.008011f
C25243 VDD.n6505 VSS 0.04401f
C25244 VDD.t4957 VSS 0.008011f
C25245 VDD.t4917 VSS 0.008011f
C25246 VDD.n6506 VSS 0.029389f
C25247 VDD.n6507 VSS 0.144542f
C25248 VDD.t4966 VSS 0.008011f
C25249 VDD.t4862 VSS 0.008011f
C25250 VDD.n6508 VSS 0.029389f
C25251 VDD.n6509 VSS 0.102512f
C25252 VDD.t4811 VSS 0.008011f
C25253 VDD.t4975 VSS 0.008011f
C25254 VDD.n6510 VSS 0.029389f
C25255 VDD.n6511 VSS 0.041173f
C25256 VDD.n6512 VSS 0.066805f
C25257 VDD.t4952 VSS 0.008011f
C25258 VDD.t4844 VSS 0.008011f
C25259 VDD.n6513 VSS 0.029389f
C25260 VDD.n6514 VSS 0.099866f
C25261 VDD.t4977 VSS 0.008011f
C25262 VDD.t4980 VSS 0.008011f
C25263 VDD.n6515 VSS 0.029389f
C25264 VDD.n6516 VSS 0.10251f
C25265 VDD.t4981 VSS 0.008011f
C25266 VDD.t4907 VSS 0.008011f
C25267 VDD.n6517 VSS 0.029389f
C25268 VDD.n6518 VSS 0.102512f
C25269 VDD.t4864 VSS 0.008011f
C25270 VDD.t4814 VSS 0.008011f
C25271 VDD.n6519 VSS 0.029389f
C25272 VDD.n6520 VSS 0.063034f
C25273 VDD.n6521 VSS 0.342598f
C25274 VDD.n6522 VSS 0.328043f
C25275 VDD.n6523 VSS 0.025494f
C25276 VDD.n6524 VSS 0.010511f
C25277 VDD.n6525 VSS 0.019376f
C25278 VDD.n6526 VSS 0.019381f
C25279 VDD.n6527 VSS 0.010511f
C25280 VDD.n6528 VSS 0.062177f
C25281 VDD.n6529 VSS 0.062181f
C25282 VDD.n6530 VSS 0.010511f
C25283 VDD.n6531 VSS 0.019376f
C25284 VDD.n6532 VSS 0.019381f
C25285 VDD.n6533 VSS 0.010511f
C25286 VDD.n6534 VSS 0.061871f
C25287 VDD.n6535 VSS 0.061149f
C25288 VDD.n6536 VSS 0.326603f
C25289 VDD.t4968 VSS 0.008011f
C25290 VDD.t4953 VSS 0.008011f
C25291 VDD.n6537 VSS 0.0221f
C25292 VDD.t4828 VSS 0.008011f
C25293 VDD.t4818 VSS 0.008011f
C25294 VDD.n6538 VSS 0.020181f
C25295 VDD.n6539 VSS 0.124159f
C25296 VDD.t4846 VSS 0.022609f
C25297 VDD.t4901 VSS 0.02098f
C25298 VDD.n6540 VSS 0.071904f
C25299 VDD.n6541 VSS 0.142473f
C25300 VDD.t4868 VSS 0.022609f
C25301 VDD.t4916 VSS 0.02098f
C25302 VDD.n6542 VSS 0.071904f
C25303 VDD.n6543 VSS 0.086055f
C25304 VDD.t4841 VSS 0.008011f
C25305 VDD.t4970 VSS 0.008011f
C25306 VDD.n6544 VSS 0.0221f
C25307 VDD.t4894 VSS 0.008011f
C25308 VDD.t4829 VSS 0.008011f
C25309 VDD.n6545 VSS 0.020181f
C25310 VDD.n6546 VSS 0.055665f
C25311 VDD.n6547 VSS 0.1321f
C25312 VDD.n6548 VSS 0.152036f
C25313 VDD.n6549 VSS 0.283978f
C25314 VDD.n6550 VSS 0.25413f
C25315 VDD.n6551 VSS 0.066805f
C25316 VDD.t4875 VSS 0.008011f
C25317 VDD.t4961 VSS 0.008011f
C25318 VDD.n6552 VSS 0.029389f
C25319 VDD.n6553 VSS 0.099866f
C25320 VDD.t4900 VSS 0.008011f
C25321 VDD.t4905 VSS 0.008011f
C25322 VDD.n6554 VSS 0.029389f
C25323 VDD.n6555 VSS 0.10251f
C25324 VDD.t4909 VSS 0.008011f
C25325 VDD.t4827 VSS 0.008011f
C25326 VDD.n6556 VSS 0.029389f
C25327 VDD.n6557 VSS 0.102512f
C25328 VDD.t4978 VSS 0.008011f
C25329 VDD.t4915 VSS 0.008011f
C25330 VDD.n6558 VSS 0.029389f
C25331 VDD.n6559 VSS 0.063034f
C25332 VDD.n6560 VSS 0.257563f
C25333 VDD.n6561 VSS 0.041023f
C25334 VDD.n6562 VSS 0.041824f
C25335 VDD.n6563 VSS 0.084772f
C25336 VDD.n6564 VSS 0.016021f
C25337 VDD.t2949 VSS 0.016021f
C25338 VDD.n6565 VSS 0.016021f
C25339 VDD.n6566 VSS 0.102784f
C25340 VDD.t3768 VSS 0.066856f
C25341 VDD.n6567 VSS 0.126716f
C25342 VDD.n6568 VSS 0.102784f
C25343 VDD.n6569 VSS 0.016021f
C25344 VDD.t1321 VSS 0.025104f
C25345 VDD.n6570 VSS 0.107953f
C25346 VDD.n6571 VSS 0.107953f
C25347 VDD.t853 VSS 0.025104f
C25348 VDD.n6572 VSS 0.016021f
C25349 VDD.n6573 VSS 0.102784f
C25350 VDD.t3210 VSS 0.066856f
C25351 VDD.n6574 VSS 0.081115f
C25352 VDD.n6575 VSS 0.051392f
C25353 VDD.n6576 VSS 0.279865f
C25354 VDD.n6577 VSS 3.80896f
C25355 VDD.n6578 VSS 0.283109f
C25356 VDD.n6579 VSS 0.052949f
C25357 VDD.t4052 VSS 0.066856f
C25358 VDD.n6580 VSS 0.082848f
C25359 VDD.n6581 VSS 0.105899f
C25360 VDD.n6582 VSS 0.016021f
C25361 VDD.t1702 VSS 0.025104f
C25362 VDD.n6583 VSS 0.110991f
C25363 VDD.n6584 VSS 0.110991f
C25364 VDD.t2284 VSS 0.066856f
C25365 VDD.n6585 VSS 0.129831f
C25366 VDD.n6586 VSS 0.105899f
C25367 VDD.n6587 VSS 0.016021f
C25368 VDD.t4649 VSS 0.016021f
C25369 VDD.n6588 VSS 0.016021f
C25370 VDD.n6589 VSS 0.105899f
C25371 VDD.t3758 VSS 0.066856f
C25372 VDD.n6590 VSS 0.129831f
C25373 VDD.n6591 VSS 0.105899f
C25374 VDD.n6592 VSS 0.016021f
C25375 VDD.t2461 VSS 0.025104f
C25376 VDD.n6593 VSS 0.114533f
C25377 VDD.t1866 VSS 0.066856f
C25378 VDD.n6594 VSS 0.129831f
C25379 VDD.t1002 VSS 0.016021f
C25380 VDD.t3754 VSS 0.066856f
C25381 VDD.n6595 VSS 0.129831f
C25382 VDD.t2566 VSS 0.025104f
C25383 VDD.t3072 VSS 0.066856f
C25384 VDD.n6596 VSS 0.129831f
C25385 VDD.t1605 VSS 0.016021f
C25386 VDD.t3480 VSS 0.066856f
C25387 VDD.n6597 VSS 0.129831f
C25388 VDD.t3990 VSS 0.066856f
C25389 VDD.n6598 VSS 0.129831f
C25390 VDD.t2269 VSS 0.016021f
C25391 VDD.t1306 VSS 0.066856f
C25392 VDD.n6599 VSS 0.354366f
C25393 VDD.n6600 VSS 0.016021f
C25394 VDD.n6601 VSS 0.158321f
C25395 VDD.t2268 VSS 0.066856f
C25396 VDD.n6602 VSS 0.129831f
C25397 VDD.n6603 VSS 0.105899f
C25398 VDD.n6604 VSS 0.016021f
C25399 VDD.t3991 VSS 0.025104f
C25400 VDD.n6605 VSS 0.110991f
C25401 VDD.n6606 VSS 0.110991f
C25402 VDD.t3481 VSS 0.025104f
C25403 VDD.n6607 VSS 0.016021f
C25404 VDD.n6608 VSS 0.105899f
C25405 VDD.t1604 VSS 0.066856f
C25406 VDD.n6609 VSS 0.082848f
C25407 VDD.n6610 VSS 0.052949f
C25408 VDD.n6611 VSS 0.099933f
C25409 VDD.n6612 VSS 0.016021f
C25410 VDD.t3073 VSS 0.025104f
C25411 VDD.n6613 VSS 0.110991f
C25412 VDD.n6614 VSS 0.110991f
C25413 VDD.t2565 VSS 0.066856f
C25414 VDD.n6615 VSS 0.129831f
C25415 VDD.n6616 VSS 0.105899f
C25416 VDD.n6617 VSS 0.016021f
C25417 VDD.t3755 VSS 0.016021f
C25418 VDD.n6618 VSS 0.016021f
C25419 VDD.n6619 VSS 0.105899f
C25420 VDD.t1001 VSS 0.066856f
C25421 VDD.n6620 VSS 0.129831f
C25422 VDD.n6621 VSS 0.105899f
C25423 VDD.n6622 VSS 0.016021f
C25424 VDD.t1867 VSS 0.025104f
C25425 VDD.n6623 VSS 0.114533f
C25426 VDD.n6624 VSS 0.689263f
C25427 VDD.n6625 VSS 0.276054f
C25428 VDD.t3685 VSS 0.066856f
C25429 VDD.n6626 VSS 0.95381f
C25430 VDD.n6627 VSS 0.936755f
C25431 VDD.t1807 VSS 0.066856f
C25432 VDD.n6628 VSS 0.525848f
C25433 VDD.t2219 VSS 0.066856f
C25434 VDD.n6629 VSS 0.525848f
C25435 VDD.n6630 VSS 0.715132f
C25436 VDD.n6631 VSS 0.892051f
C25437 VDD.n6632 VSS 0.280759f
C25438 VDD.t63 VSS 9.428519f
C25439 VDD.t71 VSS 7.61793f
C25440 VDD.t140 VSS 7.61793f
C25441 VDD.t85 VSS 9.81076f
C25442 VDD.t889 VSS 9.19382f
C25443 VDD.n6633 VSS 12.0304f
C25444 VDD.n6634 VSS 0.280759f
C25445 VDD.n6635 VSS 0.892051f
C25446 VDD.n6636 VSS 0.652605f
C25447 VDD.t2437 VSS 0.066856f
C25448 VDD.n6637 VSS 0.525848f
C25449 VDD.t2807 VSS 0.066856f
C25450 VDD.n6638 VSS 0.525848f
C25451 VDD.n6639 VSS 0.936755f
C25452 VDD.t1075 VSS 0.066856f
C25453 VDD.n6640 VSS 0.95381f
C25454 VDD.n6641 VSS 0.944397f
C25455 VDD.t3431 VSS 0.025104f
C25456 VDD.t3430 VSS 0.066856f
C25457 VDD.t3415 VSS 0.066856f
C25458 VDD.n6642 VSS 0.414447f
C25459 VDD.t2578 VSS 0.016021f
C25460 VDD.n6643 VSS 0.016021f
C25461 VDD.t2595 VSS 0.066856f
C25462 VDD.t2596 VSS 0.016021f
C25463 VDD.n6644 VSS 0.016021f
C25464 VDD.t1123 VSS 0.066856f
C25465 VDD.t1112 VSS 0.066856f
C25466 VDD.n6645 VSS 0.414447f
C25467 VDD.t4013 VSS 0.025104f
C25468 VDD.t1124 VSS 0.016021f
C25469 VDD.n6646 VSS 0.016021f
C25470 VDD.t4026 VSS 0.066856f
C25471 VDD.t4027 VSS 0.025104f
C25472 VDD.t4507 VSS 0.025104f
C25473 VDD.t4506 VSS 0.066856f
C25474 VDD.t4492 VSS 0.066856f
C25475 VDD.n6647 VSS 0.414447f
C25476 VDD.t3193 VSS 0.016021f
C25477 VDD.t861 VSS 0.025104f
C25478 VDD.t3212 VSS 0.066856f
C25479 VDD.t3192 VSS 0.066856f
C25480 VDD.n6648 VSS 0.251808f
C25481 VDD.t860 VSS 0.066856f
C25482 VDD.t833 VSS 0.066856f
C25483 VDD.n6649 VSS 0.414447f
C25484 VDD.t1330 VSS 0.025104f
C25485 VDD.t1329 VSS 0.066856f
C25486 VDD.t1316 VSS 0.066856f
C25487 VDD.n6650 VSS 0.414447f
C25488 VDD.t3757 VSS 0.016021f
C25489 VDD.n6651 VSS 0.016021f
C25490 VDD.t3776 VSS 0.066856f
C25491 VDD.t3777 VSS 0.016021f
C25492 VDD.n6652 VSS 0.016021f
C25493 VDD.t2958 VSS 0.066856f
C25494 VDD.t2930 VSS 0.066856f
C25495 VDD.n6653 VSS 0.414447f
C25496 VDD.t1438 VSS 0.025104f
C25497 VDD.t2959 VSS 0.016021f
C25498 VDD.n6654 VSS 0.016021f
C25499 VDD.t1469 VSS 0.066856f
C25500 VDD.t1470 VSS 0.025104f
C25501 VDD.t719 VSS 0.034186f
C25502 VDD.t718 VSS 0.066856f
C25503 VDD.t697 VSS 0.066856f
C25504 VDD.n6655 VSS 0.414447f
C25505 VDD.t698 VSS 0.034186f
C25506 VDD.n6656 VSS 0.409739f
C25507 VDD.n6657 VSS 0.409739f
C25508 VDD.t1437 VSS 0.066856f
C25509 VDD.n6658 VSS 0.414447f
C25510 VDD.n6659 VSS 0.366582f
C25511 VDD.n6660 VSS 0.016021f
C25512 VDD.t2931 VSS 0.016021f
C25513 VDD.n6661 VSS 0.016021f
C25514 VDD.n6662 VSS 0.366582f
C25515 VDD.t3756 VSS 0.066856f
C25516 VDD.n6663 VSS 0.414447f
C25517 VDD.n6664 VSS 0.366582f
C25518 VDD.n6665 VSS 0.016021f
C25519 VDD.t1317 VSS 0.025104f
C25520 VDD.n6666 VSS 0.372952f
C25521 VDD.n6667 VSS 0.372952f
C25522 VDD.t834 VSS 0.025104f
C25523 VDD.n6668 VSS 0.016021f
C25524 VDD.n6669 VSS 0.366582f
C25525 VDD.n6670 VSS 0.016021f
C25526 VDD.t3213 VSS 0.016021f
C25527 VDD.n6671 VSS 0.016021f
C25528 VDD.n6672 VSS 0.34593f
C25529 VDD.n6673 VSS 0.016021f
C25530 VDD.t4493 VSS 0.025104f
C25531 VDD.n6674 VSS 0.372952f
C25532 VDD.n6675 VSS 0.372952f
C25533 VDD.t4012 VSS 0.066856f
C25534 VDD.n6676 VSS 0.414447f
C25535 VDD.n6677 VSS 0.366582f
C25536 VDD.n6678 VSS 0.016021f
C25537 VDD.t1113 VSS 0.016021f
C25538 VDD.n6679 VSS 0.016021f
C25539 VDD.n6680 VSS 0.366582f
C25540 VDD.t2577 VSS 0.066856f
C25541 VDD.n6681 VSS 0.414447f
C25542 VDD.n6682 VSS 0.366582f
C25543 VDD.n6683 VSS 0.016021f
C25544 VDD.t3416 VSS 0.025104f
C25545 VDD.n6684 VSS 0.385214f
C25546 VDD.n6685 VSS 1.78684f
C25547 VDD.n6686 VSS 0.945092f
C25548 VDD.t1061 VSS 0.066856f
C25549 VDD.n6687 VSS 0.95381f
C25550 VDD.n6688 VSS 0.936755f
C25551 VDD.t3560 VSS 0.066856f
C25552 VDD.n6689 VSS 0.525848f
C25553 VDD.t3928 VSS 0.066856f
C25554 VDD.n6690 VSS 0.525848f
C25555 VDD.n6691 VSS 0.715132f
C25556 VDD.n6692 VSS 0.892051f
C25557 VDD.n6693 VSS 0.652605f
C25558 VDD.t1639 VSS 0.066856f
C25559 VDD.n6694 VSS 0.525848f
C25560 VDD.t2016 VSS 0.066856f
C25561 VDD.n6695 VSS 0.525848f
C25562 VDD.n6696 VSS 0.936755f
C25563 VDD.t4308 VSS 0.066856f
C25564 VDD.n6697 VSS 0.95381f
C25565 VDD.n6698 VSS 0.537972f
C25566 VDD.n6699 VSS 0.812758f
C25567 VDD.n6700 VSS 0.538667f
C25568 VDD.t2293 VSS 0.066856f
C25569 VDD.n6701 VSS 0.95381f
C25570 VDD.n6702 VSS 0.936755f
C25571 VDD.t4740 VSS 0.066856f
C25572 VDD.n6703 VSS 0.525848f
C25573 VDD.t992 VSS 0.066856f
C25574 VDD.n6704 VSS 0.525848f
C25575 VDD.n6705 VSS 0.715132f
C25576 VDD.n6706 VSS 0.892051f
C25577 VDD.n6707 VSS 0.652605f
C25578 VDD.t4090 VSS 0.066856f
C25579 VDD.n6708 VSS 0.525848f
C25580 VDD.t4424 VSS 0.066856f
C25581 VDD.n6709 VSS 0.525848f
C25582 VDD.n6710 VSS 0.936755f
C25583 VDD.t2872 VSS 0.066856f
C25584 VDD.n6711 VSS 0.95381f
C25585 VDD.n6712 VSS 0.749174f
C25586 VDD.n6713 VSS 1.39946f
C25587 VDD.n6714 VSS 0.186728f
C25588 VDD.t1008 VSS 0.025329f
C25589 VDD.t2947 VSS 0.016021f
C25590 VDD.t1553 VSS 0.066856f
C25591 VDD.n6715 VSS 0.126716f
C25592 VDD.t2105 VSS 0.066856f
C25593 VDD.n6716 VSS 0.126716f
C25594 VDD.n6717 VSS 0.016021f
C25595 VDD.t2106 VSS 0.025104f
C25596 VDD.n6718 VSS 0.107953f
C25597 VDD.n6719 VSS 0.107953f
C25598 VDD.t1554 VSS 0.025104f
C25599 VDD.n6720 VSS 0.016021f
C25600 VDD.n6721 VSS 0.102784f
C25601 VDD.t2946 VSS 0.066856f
C25602 VDD.n6722 VSS 0.126716f
C25603 VDD.n6723 VSS 0.102784f
C25604 VDD.n6724 VSS 0.016021f
C25605 VDD.t4245 VSS 0.016021f
C25606 VDD.n6725 VSS 0.016021f
C25607 VDD.n6726 VSS 0.087513f
C25608 VDD.n6727 VSS 0.050646f
C25609 VDD.n6728 VSS 0.388663f
C25610 VDD.n6729 VSS 0.00473f
C25611 VDD.t103 VSS 0.020865f
C25612 VDD.n6730 VSS 0.028664f
C25613 VDD.n6731 VSS 0.00473f
C25614 VDD.t182 VSS 0.008011f
C25615 VDD.t68 VSS 0.008011f
C25616 VDD.n6732 VSS 0.020046f
C25617 VDD.n6733 VSS 0.020708f
C25618 VDD.n6734 VSS 0.00473f
C25619 VDD.t80 VSS 0.020865f
C25620 VDD.n6735 VSS 0.028664f
C25621 VDD.t161 VSS 0.008011f
C25622 VDD.t258 VSS 0.008011f
C25623 VDD.n6736 VSS 0.069277f
C25624 VDD.n6737 VSS 0.149006f
C25625 VDD.n6738 VSS 0.010511f
C25626 VDD.n6739 VSS 0.040406f
C25627 VDD.n6740 VSS 0.00473f
C25628 VDD.t153 VSS 0.020865f
C25629 VDD.n6741 VSS 0.028664f
C25630 VDD.t226 VSS 0.008011f
C25631 VDD.t92 VSS 0.008011f
C25632 VDD.n6742 VSS 0.069277f
C25633 VDD.n6743 VSS 0.149006f
C25634 VDD.n6744 VSS 0.010511f
C25635 VDD.n6745 VSS 0.040406f
C25636 VDD.n6746 VSS 0.212121f
C25637 VDD.n6747 VSS 0.00473f
C25638 VDD.t171 VSS 0.020865f
C25639 VDD.n6748 VSS 0.028664f
C25640 VDD.n6749 VSS 0.00473f
C25641 VDD.t246 VSS 0.008011f
C25642 VDD.t149 VSS 0.008011f
C25643 VDD.n6750 VSS 0.020046f
C25644 VDD.n6751 VSS 0.020708f
C25645 VDD.n6752 VSS 0.111886f
C25646 VDD.n6753 VSS 0.010511f
C25647 VDD.n6754 VSS 0.019243f
C25648 VDD.n6755 VSS 0.019257f
C25649 VDD.n6756 VSS 0.010511f
C25650 VDD.n6757 VSS 0.096376f
C25651 VDD.n6758 VSS 0.535333f
C25652 VDD.t108 VSS 0.008011f
C25653 VDD.t160 VSS 0.008011f
C25654 VDD.n6759 VSS 0.024025f
C25655 VDD.t212 VSS 0.008011f
C25656 VDD.t263 VSS 0.008011f
C25657 VDD.n6760 VSS 0.018621f
C25658 VDD.n6761 VSS 0.055299f
C25659 VDD.n6762 VSS 0.047999f
C25660 VDD.t235 VSS 0.008011f
C25661 VDD.t64 VSS 0.008011f
C25662 VDD.n6763 VSS 0.024025f
C25663 VDD.t110 VSS 0.008011f
C25664 VDD.t181 VSS 0.008011f
C25665 VDD.n6764 VSS 0.018621f
C25666 VDD.n6765 VSS 0.055299f
C25667 VDD.n6766 VSS 0.086287f
C25668 VDD.t225 VSS 0.008011f
C25669 VDD.t87 VSS 0.008011f
C25670 VDD.n6767 VSS 0.024025f
C25671 VDD.t94 VSS 0.008011f
C25672 VDD.t191 VSS 0.008011f
C25673 VDD.n6768 VSS 0.018621f
C25674 VDD.n6769 VSS 0.055299f
C25675 VDD.n6770 VSS 0.086289f
C25676 VDD.t142 VSS 0.008011f
C25677 VDD.t218 VSS 0.008011f
C25678 VDD.n6771 VSS 0.024025f
C25679 VDD.t242 VSS 0.008011f
C25680 VDD.t89 VSS 0.008011f
C25681 VDD.n6772 VSS 0.018621f
C25682 VDD.n6773 VSS 0.055299f
C25683 VDD.n6774 VSS 0.085099f
C25684 VDD.t148 VSS 0.008011f
C25685 VDD.t192 VSS 0.008011f
C25686 VDD.n6775 VSS 0.024025f
C25687 VDD.t248 VSS 0.008011f
C25688 VDD.t59 VSS 0.008011f
C25689 VDD.n6776 VSS 0.018621f
C25690 VDD.n6777 VSS 0.077103f
C25691 VDD.t147 VSS 0.008011f
C25692 VDD.t55 VSS 0.008011f
C25693 VDD.n6778 VSS 0.024025f
C25694 VDD.t247 VSS 0.008011f
C25695 VDD.t172 VSS 0.008011f
C25696 VDD.n6779 VSS 0.018621f
C25697 VDD.n6780 VSS 0.055299f
C25698 VDD.n6781 VSS 0.111411f
C25699 VDD.t158 VSS 0.008011f
C25700 VDD.t231 VSS 0.008011f
C25701 VDD.n6782 VSS 0.024025f
C25702 VDD.t262 VSS 0.008011f
C25703 VDD.t107 VSS 0.008011f
C25704 VDD.n6783 VSS 0.018621f
C25705 VDD.n6784 VSS 0.055299f
C25706 VDD.n6785 VSS 0.086287f
C25707 VDD.t240 VSS 0.008011f
C25708 VDD.t70 VSS 0.008011f
C25709 VDD.n6786 VSS 0.024025f
C25710 VDD.t114 VSS 0.008011f
C25711 VDD.t187 VSS 0.008011f
C25712 VDD.n6787 VSS 0.018621f
C25713 VDD.n6788 VSS 0.055299f
C25714 VDD.n6789 VSS 0.022927f
C25715 VDD.n6790 VSS 0.067373f
C25716 VDD.n6791 VSS 0.472695f
C25717 VDD.t257 VSS 0.008011f
C25718 VDD.t100 VSS 0.008011f
C25719 VDD.n6792 VSS 0.032022f
C25720 VDD.n6793 VSS 0.116906f
C25721 VDD.t228 VSS 0.031728f
C25722 VDD.n6794 VSS 0.151284f
C25723 VDD.t180 VSS 0.061518f
C25724 VDD.t236 VSS 0.008011f
C25725 VDD.t77 VSS 0.008011f
C25726 VDD.n6795 VSS 0.032022f
C25727 VDD.n6796 VSS 0.216759f
C25728 VDD.n6797 VSS 0.152023f
C25729 VDD.n6798 VSS 0.339165f
C25730 VDD.n6799 VSS 0.303879f
C25731 VDD.n6800 VSS 0.147417f
C25732 VDD.n6801 VSS 0.111886f
C25733 VDD.n6802 VSS 0.010511f
C25734 VDD.n6803 VSS 0.019243f
C25735 VDD.n6804 VSS 0.019257f
C25736 VDD.n6805 VSS 0.010511f
C25737 VDD.n6806 VSS 0.061022f
C25738 VDD.n6807 VSS 0.334665f
C25739 VDD.t241 VSS 0.008011f
C25740 VDD.t283 VSS 0.008011f
C25741 VDD.n6808 VSS 0.024025f
C25742 VDD.t184 VSS 0.008011f
C25743 VDD.t230 VSS 0.008011f
C25744 VDD.n6809 VSS 0.018621f
C25745 VDD.n6810 VSS 0.077103f
C25746 VDD.t239 VSS 0.008011f
C25747 VDD.t164 VSS 0.008011f
C25748 VDD.n6811 VSS 0.024025f
C25749 VDD.t183 VSS 0.008011f
C25750 VDD.t106 VSS 0.008011f
C25751 VDD.n6812 VSS 0.018621f
C25752 VDD.n6813 VSS 0.055299f
C25753 VDD.n6814 VSS 0.111411f
C25754 VDD.t252 VSS 0.008011f
C25755 VDD.t95 VSS 0.008011f
C25756 VDD.n6815 VSS 0.024025f
C25757 VDD.t193 VSS 0.008011f
C25758 VDD.t268 VSS 0.008011f
C25759 VDD.n6816 VSS 0.018621f
C25760 VDD.n6817 VSS 0.055299f
C25761 VDD.n6818 VSS 0.086287f
C25762 VDD.t104 VSS 0.008011f
C25763 VDD.t176 VSS 0.008011f
C25764 VDD.n6819 VSS 0.024025f
C25765 VDD.t274 VSS 0.008011f
C25766 VDD.t117 VSS 0.008011f
C25767 VDD.n6820 VSS 0.018621f
C25768 VDD.n6821 VSS 0.055299f
C25769 VDD.n6822 VSS 0.022927f
C25770 VDD.n6823 VSS 0.067373f
C25771 VDD.t234 VSS 0.008011f
C25772 VDD.t74 VSS 0.008011f
C25773 VDD.n6824 VSS 0.024025f
C25774 VDD.t177 VSS 0.008011f
C25775 VDD.t254 VSS 0.008011f
C25776 VDD.n6825 VSS 0.018621f
C25777 VDD.n6826 VSS 0.055299f
C25778 VDD.n6827 VSS 0.085099f
C25779 VDD.t84 VSS 0.008011f
C25780 VDD.t186 VSS 0.008011f
C25781 VDD.n6828 VSS 0.024025f
C25782 VDD.t261 VSS 0.008011f
C25783 VDD.t129 VSS 0.008011f
C25784 VDD.n6829 VSS 0.018621f
C25785 VDD.n6830 VSS 0.055299f
C25786 VDD.n6831 VSS 0.086289f
C25787 VDD.t96 VSS 0.008011f
C25788 VDD.t170 VSS 0.008011f
C25789 VDD.n6832 VSS 0.024025f
C25790 VDD.t270 VSS 0.008011f
C25791 VDD.t113 VSS 0.008011f
C25792 VDD.n6833 VSS 0.018621f
C25793 VDD.n6834 VSS 0.055299f
C25794 VDD.n6835 VSS 0.086287f
C25795 VDD.t206 VSS 0.008011f
C25796 VDD.t255 VSS 0.008011f
C25797 VDD.n6836 VSS 0.024025f
C25798 VDD.t150 VSS 0.008011f
C25799 VDD.t195 VSS 0.008011f
C25800 VDD.n6837 VSS 0.018621f
C25801 VDD.n6838 VSS 0.055299f
C25802 VDD.n6839 VSS 0.047999f
C25803 VDD.n6840 VSS 0.309204f
C25804 VDD.n6841 VSS 0.324728f
C25805 VDD.t121 VSS 0.008011f
C25806 VDD.t199 VSS 0.008011f
C25807 VDD.n6842 VSS 0.032022f
C25808 VDD.n6843 VSS 0.116906f
C25809 VDD.t93 VSS 0.031728f
C25810 VDD.n6844 VSS 0.151284f
C25811 VDD.t272 VSS 0.061518f
C25812 VDD.t97 VSS 0.008011f
C25813 VDD.t179 VSS 0.008011f
C25814 VDD.n6845 VSS 0.032022f
C25815 VDD.n6846 VSS 0.216759f
C25816 VDD.n6847 VSS 0.152023f
C25817 VDD.n6848 VSS 0.27523f
C25818 VDD.n6849 VSS 0.050646f
C25819 VDD.n6850 VSS 0.087513f
C25820 VDD.n6851 VSS 0.016021f
C25821 VDD.t1464 VSS 0.016021f
C25822 VDD.n6852 VSS 0.016021f
C25823 VDD.n6853 VSS 0.102784f
C25824 VDD.t4268 VSS 0.066856f
C25825 VDD.n6854 VSS 0.126716f
C25826 VDD.n6855 VSS 0.102784f
C25827 VDD.n6856 VSS 0.016021f
C25828 VDD.t2977 VSS 0.025104f
C25829 VDD.n6857 VSS 0.107953f
C25830 VDD.n6858 VSS 0.107953f
C25831 VDD.t2557 VSS 0.025104f
C25832 VDD.n6859 VSS 0.016021f
C25833 VDD.n6860 VSS 0.096993f
C25834 VDD.n6861 VSS 0.051392f
C25835 VDD.t1095 VSS 0.066856f
C25836 VDD.n6862 VSS 0.081115f
C25837 VDD.n6863 VSS 0.102784f
C25838 VDD.n6864 VSS 0.016021f
C25839 VDD.t3515 VSS 0.025104f
C25840 VDD.n6865 VSS 0.107953f
C25841 VDD.n6866 VSS 0.107953f
C25842 VDD.t4478 VSS 0.066856f
C25843 VDD.n6867 VSS 0.126716f
C25844 VDD.n6868 VSS 0.102784f
C25845 VDD.n6869 VSS 0.016021f
C25846 VDD.t1690 VSS 0.016021f
C25847 VDD.n6870 VSS 0.016021f
C25848 VDD.n6871 VSS 0.102784f
C25849 VDD.t4474 VSS 0.066856f
C25850 VDD.n6872 VSS 0.126716f
C25851 VDD.n6873 VSS 0.084772f
C25852 VDD.n6874 VSS 0.016021f
C25853 VDD.t3590 VSS 0.025104f
C25854 VDD.n6875 VSS 0.1306f
C25855 VDD.n6876 VSS 0.05157f
C25856 VDD.n6877 VSS 0.041023f
C25857 VDD.n6878 VSS 0.342598f
C25858 VDD.n6879 VSS 0.00473f
C25859 VDD.n6880 VSS 0.00473f
C25860 VDD.n6881 VSS 0.00473f
C25861 VDD.n6882 VSS 0.00473f
C25862 VDD.n6883 VSS 0.00473f
C25863 VDD.n6884 VSS 0.00473f
C25864 VDD.n6885 VSS 0.00473f
C25865 VDD.t167 VSS 0.008011f
C25866 VDD.t219 VSS 0.008011f
C25867 VDD.n6886 VSS 0.042109f
C25868 VDD.n6887 VSS 0.063057f
C25869 VDD.t287 VSS 0.008011f
C25870 VDD.t135 VSS 0.008011f
C25871 VDD.n6888 VSS 0.018495f
C25872 VDD.n6889 VSS 0.016425f
C25873 VDD.n6890 VSS 0.010511f
C25874 VDD.n6891 VSS 0.062181f
C25875 VDD.n6892 VSS 0.062177f
C25876 VDD.t276 VSS 0.008011f
C25877 VDD.t151 VSS 0.008011f
C25878 VDD.n6893 VSS 0.018495f
C25879 VDD.n6894 VSS 0.016425f
C25880 VDD.n6895 VSS 0.010511f
C25881 VDD.n6896 VSS 0.019381f
C25882 VDD.n6897 VSS 0.019376f
C25883 VDD.t196 VSS 0.008011f
C25884 VDD.t271 VSS 0.008011f
C25885 VDD.n6898 VSS 0.018495f
C25886 VDD.n6899 VSS 0.016425f
C25887 VDD.n6900 VSS 0.010511f
C25888 VDD.n6901 VSS 0.00416f
C25889 VDD.n6902 VSS 0.00473f
C25890 VDD.n6903 VSS 0.00473f
C25891 VDD.n6904 VSS 0.00473f
C25892 VDD.t232 VSS 0.008011f
C25893 VDD.t278 VSS 0.008011f
C25894 VDD.n6905 VSS 0.042109f
C25895 VDD.n6906 VSS 0.063057f
C25896 VDD.t132 VSS 0.008011f
C25897 VDD.t201 VSS 0.008011f
C25898 VDD.n6907 VSS 0.018495f
C25899 VDD.n6908 VSS 0.016425f
C25900 VDD.n6909 VSS 0.010511f
C25901 VDD.n6910 VSS 0.062181f
C25902 VDD.n6911 VSS 0.062177f
C25903 VDD.t116 VSS 0.008011f
C25904 VDD.t213 VSS 0.008011f
C25905 VDD.n6912 VSS 0.018495f
C25906 VDD.n6913 VSS 0.016425f
C25907 VDD.n6914 VSS 0.010511f
C25908 VDD.n6915 VSS 0.019381f
C25909 VDD.n6916 VSS 0.019376f
C25910 VDD.t264 VSS 0.008011f
C25911 VDD.t111 VSS 0.008011f
C25912 VDD.n6917 VSS 0.018495f
C25913 VDD.n6918 VSS 0.016425f
C25914 VDD.n6919 VSS 0.010511f
C25915 VDD.n6920 VSS 0.00416f
C25916 VDD.n6921 VSS 0.132226f
C25917 VDD.t273 VSS 0.008011f
C25918 VDD.t122 VSS 0.008011f
C25919 VDD.n6922 VSS 0.0221f
C25920 VDD.t155 VSS 0.008011f
C25921 VDD.t227 VSS 0.008011f
C25922 VDD.n6923 VSS 0.020181f
C25923 VDD.n6924 VSS 0.124159f
C25924 VDD.t250 VSS 0.022609f
C25925 VDD.t127 VSS 0.02098f
C25926 VDD.n6925 VSS 0.071904f
C25927 VDD.n6926 VSS 0.142473f
C25928 VDD.n6927 VSS 0.00473f
C25929 VDD.n6928 VSS 0.00473f
C25930 VDD.n6929 VSS 0.00473f
C25931 VDD.n6930 VSS 0.00473f
C25932 VDD.n6931 VSS 0.061871f
C25933 VDD.t136 VSS 0.008011f
C25934 VDD.t207 VSS 0.008011f
C25935 VDD.n6932 VSS 0.018495f
C25936 VDD.n6933 VSS 0.016425f
C25937 VDD.n6934 VSS 0.010511f
C25938 VDD.n6935 VSS 0.019381f
C25939 VDD.n6936 VSS 0.019376f
C25940 VDD.t277 VSS 0.008011f
C25941 VDD.t130 VSS 0.008011f
C25942 VDD.n6937 VSS 0.018495f
C25943 VDD.n6938 VSS 0.016425f
C25944 VDD.n6939 VSS 0.010511f
C25945 VDD.n6940 VSS 0.062181f
C25946 VDD.n6941 VSS 0.062177f
C25947 VDD.t265 VSS 0.008011f
C25948 VDD.t190 VSS 0.008011f
C25949 VDD.n6942 VSS 0.018495f
C25950 VDD.n6943 VSS 0.016425f
C25951 VDD.n6944 VSS 0.010511f
C25952 VDD.n6945 VSS 0.019381f
C25953 VDD.n6946 VSS 0.019376f
C25954 VDD.t266 VSS 0.008011f
C25955 VDD.t88 VSS 0.008011f
C25956 VDD.n6947 VSS 0.018495f
C25957 VDD.n6948 VSS 0.016425f
C25958 VDD.n6949 VSS 0.010511f
C25959 VDD.n6950 VSS 0.093664f
C25960 VDD.n6951 VSS 0.507601f
C25961 VDD.t200 VSS 0.022609f
C25962 VDD.t62 VSS 0.02098f
C25963 VDD.n6952 VSS 0.071904f
C25964 VDD.n6953 VSS 0.086055f
C25965 VDD.t256 VSS 0.008011f
C25966 VDD.t98 VSS 0.008011f
C25967 VDD.n6954 VSS 0.0221f
C25968 VDD.t133 VSS 0.008011f
C25969 VDD.t208 VSS 0.008011f
C25970 VDD.n6955 VSS 0.020181f
C25971 VDD.n6956 VSS 0.055665f
C25972 VDD.n6957 VSS 0.1321f
C25973 VDD.n6958 VSS 0.152036f
C25974 VDD.n6959 VSS 0.466322f
C25975 VDD.t86 VSS 0.008011f
C25976 VDD.t141 VSS 0.008011f
C25977 VDD.n6960 VSS 0.04401f
C25978 VDD.t216 VSS 0.008011f
C25979 VDD.t279 VSS 0.008011f
C25980 VDD.n6961 VSS 0.029389f
C25981 VDD.n6962 VSS 0.144542f
C25982 VDD.t203 VSS 0.008011f
C25983 VDD.t57 VSS 0.008011f
C25984 VDD.n6963 VSS 0.029389f
C25985 VDD.n6964 VSS 0.102512f
C25986 VDD.t119 VSS 0.008011f
C25987 VDD.t194 VSS 0.008011f
C25988 VDD.n6965 VSS 0.029389f
C25989 VDD.n6966 VSS 0.041173f
C25990 VDD.t126 VSS 0.008011f
C25991 VDD.t173 VSS 0.008011f
C25992 VDD.n6967 VSS 0.029389f
C25993 VDD.n6968 VSS 0.063034f
C25994 VDD.t124 VSS 0.008011f
C25995 VDD.t275 VSS 0.008011f
C25996 VDD.n6969 VSS 0.029389f
C25997 VDD.n6970 VSS 0.102512f
C25998 VDD.t138 VSS 0.008011f
C25999 VDD.t211 VSS 0.008011f
C26000 VDD.n6971 VSS 0.029389f
C26001 VDD.n6972 VSS 0.10251f
C26002 VDD.t222 VSS 0.008011f
C26003 VDD.t284 VSS 0.008011f
C26004 VDD.n6973 VSS 0.029389f
C26005 VDD.n6974 VSS 0.099866f
C26006 VDD.n6975 VSS 0.066805f
C26007 VDD.n6976 VSS 0.339165f
C26008 VDD.n6977 VSS 0.326603f
C26009 VDD.n6978 VSS 0.061149f
C26010 VDD.n6979 VSS 0.061871f
C26011 VDD.t53 VSS 0.008011f
C26012 VDD.t139 VSS 0.008011f
C26013 VDD.n6980 VSS 0.018495f
C26014 VDD.n6981 VSS 0.016425f
C26015 VDD.n6982 VSS 0.010511f
C26016 VDD.n6983 VSS 0.019381f
C26017 VDD.n6984 VSS 0.019376f
C26018 VDD.t215 VSS 0.008011f
C26019 VDD.t286 VSS 0.008011f
C26020 VDD.n6985 VSS 0.018495f
C26021 VDD.n6986 VSS 0.016425f
C26022 VDD.n6987 VSS 0.010511f
C26023 VDD.n6988 VSS 0.062181f
C26024 VDD.n6989 VSS 0.062177f
C26025 VDD.t202 VSS 0.008011f
C26026 VDD.t128 VSS 0.008011f
C26027 VDD.n6990 VSS 0.018495f
C26028 VDD.n6991 VSS 0.016425f
C26029 VDD.n6992 VSS 0.010511f
C26030 VDD.n6993 VSS 0.019381f
C26031 VDD.n6994 VSS 0.019376f
C26032 VDD.t204 VSS 0.008011f
C26033 VDD.t253 VSS 0.008011f
C26034 VDD.n6995 VSS 0.018495f
C26035 VDD.n6996 VSS 0.016425f
C26036 VDD.n6997 VSS 0.010511f
C26037 VDD.n6998 VSS 0.025494f
C26038 VDD.n6999 VSS 0.328043f
C26039 VDD.t145 VSS 0.008011f
C26040 VDD.t220 VSS 0.008011f
C26041 VDD.n7000 VSS 0.0221f
C26042 VDD.t82 VSS 0.008011f
C26043 VDD.t162 VSS 0.008011f
C26044 VDD.n7001 VSS 0.020181f
C26045 VDD.n7002 VSS 0.124159f
C26046 VDD.t115 VSS 0.022609f
C26047 VDD.t282 VSS 0.02098f
C26048 VDD.n7003 VSS 0.071904f
C26049 VDD.n7004 VSS 0.142473f
C26050 VDD.n7005 VSS 0.152036f
C26051 VDD.t120 VSS 0.008011f
C26052 VDD.t198 VSS 0.008011f
C26053 VDD.n7006 VSS 0.0221f
C26054 VDD.t288 VSS 0.008011f
C26055 VDD.t144 VSS 0.008011f
C26056 VDD.n7007 VSS 0.020181f
C26057 VDD.n7008 VSS 0.055665f
C26058 VDD.n7009 VSS 0.1321f
C26059 VDD.t289 VSS 0.022609f
C26060 VDD.t237 VSS 0.02098f
C26061 VDD.n7010 VSS 0.071904f
C26062 VDD.n7011 VSS 0.086055f
C26063 VDD.n7012 VSS 0.32091f
C26064 VDD.n7013 VSS 0.257563f
C26065 VDD.t223 VSS 0.008011f
C26066 VDD.t267 VSS 0.008011f
C26067 VDD.n7014 VSS 0.029389f
C26068 VDD.n7015 VSS 0.063034f
C26069 VDD.t221 VSS 0.008011f
C26070 VDD.t146 VSS 0.008011f
C26071 VDD.n7016 VSS 0.029389f
C26072 VDD.n7017 VSS 0.102512f
C26073 VDD.t229 VSS 0.008011f
C26074 VDD.t66 VSS 0.008011f
C26075 VDD.n7018 VSS 0.029389f
C26076 VDD.n7019 VSS 0.10251f
C26077 VDD.t83 VSS 0.008011f
C26078 VDD.t157 VSS 0.008011f
C26079 VDD.n7020 VSS 0.029389f
C26080 VDD.n7021 VSS 0.099866f
C26081 VDD.n7022 VSS 0.066805f
C26082 VDD.n7023 VSS 0.25413f
C26083 VDD.n7024 VSS 0.041023f
C26084 VDD.n7025 VSS 0.041824f
C26085 VDD.n7026 VSS 0.084772f
C26086 VDD.n7027 VSS 0.016021f
C26087 VDD.t4555 VSS 0.016021f
C26088 VDD.n7028 VSS 0.016021f
C26089 VDD.n7029 VSS 0.102784f
C26090 VDD.t1314 VSS 0.066856f
C26091 VDD.n7030 VSS 0.126716f
C26092 VDD.n7031 VSS 0.102784f
C26093 VDD.n7032 VSS 0.016021f
C26094 VDD.t3151 VSS 0.025104f
C26095 VDD.n7033 VSS 0.107953f
C26096 VDD.n7034 VSS 0.107953f
C26097 VDD.t2652 VSS 0.025104f
C26098 VDD.n7035 VSS 0.016021f
C26099 VDD.n7036 VSS 0.102784f
C26100 VDD.t725 VSS 0.066856f
C26101 VDD.n7037 VSS 0.081115f
C26102 VDD.n7038 VSS 0.051392f
C26103 VDD.n7039 VSS 0.279865f
C26104 VDD.n7040 VSS 3.80896f
C26105 VDD.n7041 VSS 0.283109f
C26106 VDD.n7042 VSS 0.283088f
C26107 VDD.n7043 VSS 0.532659f
C26108 VDD.t3931 VSS 0.034186f
C26109 VDD.t3578 VSS 0.034186f
C26110 VDD.n7044 VSS 0.43943f
C26111 VDD.t3577 VSS 0.066856f
C26112 VDD.t3930 VSS 0.066856f
C26113 VDD.n7045 VSS 0.333277f
C26114 VDD.t3268 VSS 0.066856f
C26115 VDD.t3562 VSS 0.066856f
C26116 VDD.n7046 VSS 0.333277f
C26117 VDD.t3563 VSS 0.034186f
C26118 VDD.t3269 VSS 0.034186f
C26119 VDD.n7047 VSS 0.556001f
C26120 VDD.n7048 VSS 1.1439f
C26121 VDD.n7049 VSS 0.369079f
C26122 VDD.t1064 VSS 0.034186f
C26123 VDD.n7050 VSS 0.409739f
C26124 VDD.n7051 VSS 0.409739f
C26125 VDD.t1037 VSS 0.025104f
C26126 VDD.n7052 VSS 0.016021f
C26127 VDD.n7053 VSS 0.366582f
C26128 VDD.n7054 VSS 0.016021f
C26129 VDD.t3909 VSS 0.016021f
C26130 VDD.n7055 VSS 0.016021f
C26131 VDD.n7056 VSS 0.366582f
C26132 VDD.n7057 VSS 0.016021f
C26133 VDD.t2634 VSS 0.016021f
C26134 VDD.n7058 VSS 0.016021f
C26135 VDD.n7059 VSS 0.366582f
C26136 VDD.n7060 VSS 0.016021f
C26137 VDD.t1135 VSS 0.025104f
C26138 VDD.n7061 VSS 0.372952f
C26139 VDD.t3533 VSS 0.016021f
C26140 VDD.n7062 VSS 0.016021f
C26141 VDD.t761 VSS 0.025104f
C26142 VDD.t760 VSS 0.066856f
C26143 VDD.t734 VSS 0.066856f
C26144 VDD.n7063 VSS 0.414447f
C26145 VDD.n7064 VSS 0.372952f
C26146 VDD.t735 VSS 0.025104f
C26147 VDD.n7065 VSS 0.016021f
C26148 VDD.t3521 VSS 0.016021f
C26149 VDD.t1752 VSS 0.025104f
C26150 VDD.t2855 VSS 0.025104f
C26151 VDD.t2854 VSS 0.066856f
C26152 VDD.t2840 VSS 0.066856f
C26153 VDD.n7066 VSS 0.414447f
C26154 VDD.t4143 VSS 0.016021f
C26155 VDD.n7067 VSS 0.016021f
C26156 VDD.t4158 VSS 0.066856f
C26157 VDD.t4159 VSS 0.016021f
C26158 VDD.n7068 VSS 0.016021f
C26159 VDD.t2848 VSS 0.066856f
C26160 VDD.t2832 VSS 0.066856f
C26161 VDD.n7069 VSS 0.414447f
C26162 VDD.t1816 VSS 0.025104f
C26163 VDD.t2849 VSS 0.016021f
C26164 VDD.t1835 VSS 0.025104f
C26165 VDD.n7070 VSS 0.016021f
C26166 VDD.t1834 VSS 0.066856f
C26167 VDD.t1815 VSS 0.066856f
C26168 VDD.n7071 VSS 0.414447f
C26169 VDD.n7072 VSS 0.366582f
C26170 VDD.n7073 VSS 0.016021f
C26171 VDD.t2833 VSS 0.016021f
C26172 VDD.n7074 VSS 0.016021f
C26173 VDD.n7075 VSS 0.366582f
C26174 VDD.t4142 VSS 0.066856f
C26175 VDD.n7076 VSS 0.414447f
C26176 VDD.n7077 VSS 0.366582f
C26177 VDD.n7078 VSS 0.016021f
C26178 VDD.t2841 VSS 0.025104f
C26179 VDD.n7079 VSS 0.372952f
C26180 VDD.n7080 VSS 0.372952f
C26181 VDD.t1737 VSS 0.025104f
C26182 VDD.n7081 VSS 0.016021f
C26183 VDD.n7082 VSS 0.366582f
C26184 VDD.t3520 VSS 0.066856f
C26185 VDD.n7083 VSS 0.251808f
C26186 VDD.n7084 VSS 0.183291f
C26187 VDD.n7085 VSS 0.279865f
C26188 VDD.n7086 VSS 3.80896f
C26189 VDD.n7087 VSS 0.279865f
C26190 VDD.t2702 VSS 0.066856f
C26191 VDD.t2703 VSS 0.016021f
C26192 VDD.n7088 VSS 0.016021f
C26193 VDD.t903 VSS 0.066856f
C26194 VDD.t3046 VSS 0.066856f
C26195 VDD.n7089 VSS 0.256005f
C26196 VDD.t904 VSS 0.025104f
C26197 VDD.t1841 VSS 0.025104f
C26198 VDD.t1840 VSS 0.066856f
C26199 VDD.t3970 VSS 0.066856f
C26200 VDD.n7090 VSS 0.256005f
C26201 VDD.t1150 VSS 0.016021f
C26202 VDD.n7091 VSS 0.016021f
C26203 VDD.t3282 VSS 0.066856f
C26204 VDD.t3283 VSS 0.016021f
C26205 VDD.n7092 VSS 0.016021f
C26206 VDD.t1832 VSS 0.066856f
C26207 VDD.t3964 VSS 0.066856f
C26208 VDD.n7093 VSS 0.256005f
C26209 VDD.t3109 VSS 0.025104f
C26210 VDD.t1833 VSS 0.016021f
C26211 VDD.n7094 VSS 0.016021f
C26212 VDD.t972 VSS 0.066856f
C26213 VDD.t973 VSS 0.025104f
C26214 VDD.t4337 VSS 0.034186f
C26215 VDD.t2333 VSS 0.034186f
C26216 VDD.n7095 VSS 0.239302f
C26217 VDD.n7096 VSS 0.239302f
C26218 VDD.t3108 VSS 0.066856f
C26219 VDD.n7097 VSS 0.256005f
C26220 VDD.n7098 VSS 0.208141f
C26221 VDD.n7099 VSS 0.016021f
C26222 VDD.t3965 VSS 0.016021f
C26223 VDD.n7100 VSS 0.016021f
C26224 VDD.n7101 VSS 0.208141f
C26225 VDD.t1149 VSS 0.066856f
C26226 VDD.n7102 VSS 0.256005f
C26227 VDD.n7103 VSS 0.208141f
C26228 VDD.n7104 VSS 0.016021f
C26229 VDD.t3971 VSS 0.025104f
C26230 VDD.n7105 VSS 0.218415f
C26231 VDD.n7106 VSS 0.218415f
C26232 VDD.t3047 VSS 0.025104f
C26233 VDD.n7107 VSS 0.016021f
C26234 VDD.n7108 VSS 0.208141f
C26235 VDD.t4700 VSS 0.066856f
C26236 VDD.n7109 VSS 0.163661f
C26237 VDD.n7110 VSS 0.10407f
C26238 VDD.n7111 VSS 0.196415f
C26239 VDD.n7112 VSS 0.016021f
C26240 VDD.t1922 VSS 0.025104f
C26241 VDD.n7113 VSS 0.218415f
C26242 VDD.n7114 VSS 0.218415f
C26243 VDD.t2427 VSS 0.066856f
C26244 VDD.n7115 VSS 0.256005f
C26245 VDD.n7116 VSS 0.208141f
C26246 VDD.n7117 VSS 0.016021f
C26247 VDD.t3726 VSS 0.016021f
C26248 VDD.n7118 VSS 0.016021f
C26249 VDD.n7119 VSS 0.208141f
C26250 VDD.t974 VSS 0.066856f
C26251 VDD.n7120 VSS 0.256005f
C26252 VDD.n7121 VSS 0.208141f
C26253 VDD.n7122 VSS 0.016021f
C26254 VDD.t2250 VSS 0.025104f
C26255 VDD.n7123 VSS 0.225377f
C26256 VDD.n7124 VSS 0.570644f
C26257 VDD.n7125 VSS 0.33406f
C26258 VDD.t2295 VSS 0.066856f
C26259 VDD.n7126 VSS 0.58882f
C26260 VDD.n7127 VSS 0.571765f
C26261 VDD.t4742 VSS 0.066856f
C26262 VDD.n7128 VSS 0.333277f
C26263 VDD.t994 VSS 0.066856f
C26264 VDD.n7129 VSS 0.333277f
C26265 VDD.n7130 VSS 0.43943f
C26266 VDD.n7131 VSS 0.532659f
C26267 VDD.n7132 VSS 0.280759f
C26268 VDD.n7133 VSS 4.15767f
C26269 VDD.n7134 VSS 0.280759f
C26270 VDD.n7135 VSS 0.532659f
C26271 VDD.n7136 VSS 0.402094f
C26272 VDD.t2166 VSS 0.066856f
C26273 VDD.n7137 VSS 0.333277f
C26274 VDD.t2603 VSS 0.066856f
C26275 VDD.n7138 VSS 0.333277f
C26276 VDD.n7139 VSS 0.571765f
C26277 VDD.t885 VSS 0.066856f
C26278 VDD.n7140 VSS 0.58882f
C26279 VDD.n7141 VSS 0.333645f
C26280 VDD.n7142 VSS 0.570644f
C26281 VDD.n7143 VSS 0.225377f
C26282 VDD.t851 VSS 0.025104f
C26283 VDD.n7144 VSS 0.016021f
C26284 VDD.n7145 VSS 0.208141f
C26285 VDD.n7146 VSS 0.016021f
C26286 VDD.t645 VSS 0.016021f
C26287 VDD.n7147 VSS 0.016021f
C26288 VDD.n7148 VSS 0.208141f
C26289 VDD.n7149 VSS 0.016021f
C26290 VDD.t2415 VSS 0.016021f
C26291 VDD.n7150 VSS 0.016021f
C26292 VDD.n7151 VSS 0.208141f
C26293 VDD.n7152 VSS 0.016021f
C26294 VDD.t2077 VSS 0.025104f
C26295 VDD.n7153 VSS 0.218415f
C26296 VDD.n7154 VSS 0.218415f
C26297 VDD.t1622 VSS 0.025104f
C26298 VDD.n7155 VSS 0.016021f
C26299 VDD.n7156 VSS 0.196415f
C26300 VDD.n7157 VSS 0.016021f
C26301 VDD.t3333 VSS 0.016021f
C26302 VDD.n7158 VSS 0.016021f
C26303 VDD.n7159 VSS 0.208141f
C26304 VDD.n7160 VSS 0.016021f
C26305 VDD.t2762 VSS 0.025104f
C26306 VDD.n7161 VSS 0.218415f
C26307 VDD.n7162 VSS 0.218415f
C26308 VDD.t2656 VSS 0.025104f
C26309 VDD.n7163 VSS 0.016021f
C26310 VDD.n7164 VSS 0.208141f
C26311 VDD.n7165 VSS 0.016021f
C26312 VDD.t911 VSS 0.016021f
C26313 VDD.n7166 VSS 0.016021f
C26314 VDD.n7167 VSS 0.208141f
C26315 VDD.n7168 VSS 0.016021f
C26316 VDD.t2644 VSS 0.016021f
C26317 VDD.n7169 VSS 0.016021f
C26318 VDD.n7170 VSS 0.208141f
C26319 VDD.n7171 VSS 0.016021f
C26320 VDD.t2835 VSS 0.025104f
C26321 VDD.n7172 VSS 0.239302f
C26322 VDD.n7173 VSS 0.239302f
C26323 VDD.t1978 VSS 0.034186f
C26324 VDD.n7174 VSS 0.266053f
C26325 VDD.n7175 VSS 0.501023f
C26326 VDD.n7176 VSS 0.274982f
C26327 VDD.t2315 VSS 0.066856f
C26328 VDD.n7177 VSS 0.14839f
C26329 VDD.n7178 VSS 0.012131f
C26330 VDD.n7179 VSS 0.012131f
C26331 VDD.n7180 VSS 0.012131f
C26332 VDD.n7181 VSS 0.012131f
C26333 VDD.n7182 VSS 0.012131f
C26334 VDD.n7183 VSS 0.012131f
C26335 VDD.n7184 VSS 0.012131f
C26336 VDD.n7185 VSS 0.012131f
C26337 VDD.n7186 VSS 0.012131f
C26338 VDD.n7187 VSS 0.012131f
C26339 VDD.n7188 VSS 0.012131f
C26340 VDD.n7189 VSS 0.012131f
C26341 VDD.n7190 VSS 0.012131f
C26342 VDD.n7191 VSS 0.012131f
C26343 VDD.n7192 VSS 0.012131f
C26344 VDD.n7193 VSS 0.012131f
C26345 VDD.n7194 VSS 0.012131f
C26346 VDD.n7195 VSS 0.012131f
C26347 VDD.n7196 VSS 0.012131f
C26348 VDD.n7197 VSS 0.012131f
C26349 VDD.n7198 VSS 0.012131f
C26350 VDD.n7199 VSS 0.012131f
C26351 VDD.n7200 VSS 0.012131f
C26352 VDD.n7201 VSS 0.012131f
C26353 VDD.n7202 VSS 0.012131f
C26354 VDD.n7203 VSS 0.012131f
C26355 VDD.n7204 VSS 0.012131f
C26356 VDD.n7205 VSS 0.012131f
C26357 VDD.n7206 VSS 0.012131f
C26358 VDD.n7207 VSS 0.012131f
C26359 VDD.n7208 VSS 0.012131f
C26360 VDD.n7209 VSS 0.012131f
C26361 VDD.n7210 VSS 0.012131f
C26362 VDD.n7211 VSS 0.012131f
C26363 VDD.n7212 VSS 0.012131f
C26364 VDD.n7213 VSS 0.012131f
C26365 VDD.n7214 VSS 0.012131f
C26366 VDD.n7215 VSS 0.012131f
C26367 VDD.n7216 VSS 0.012131f
C26368 VDD.n7217 VSS 0.012131f
C26369 VDD.n7218 VSS 0.012131f
C26370 VDD.n7219 VSS 0.012131f
C26371 VDD.n7220 VSS 0.012131f
C26372 VDD.n7221 VSS 0.012131f
C26373 VDD.n7222 VSS 0.012131f
C26374 VDD.n7223 VSS 0.012131f
C26375 VDD.n7224 VSS 0.012131f
C26376 VDD.n7225 VSS 0.012131f
C26377 VDD.n7226 VSS 0.012131f
C26378 VDD.n7227 VSS 0.012131f
C26379 VDD.n7228 VSS 0.012131f
C26380 VDD.n7229 VSS 0.012131f
C26381 VDD.n7230 VSS 0.012131f
C26382 VDD.n7231 VSS 0.012131f
C26383 VDD.n7232 VSS 0.012131f
C26384 VDD.n7233 VSS 0.012131f
C26385 VDD.n7234 VSS 0.012131f
C26386 VDD.n7235 VSS 0.012131f
C26387 VDD.n7236 VSS 0.012131f
C26388 VDD.n7237 VSS 0.012131f
C26389 VDD.n7238 VSS 0.012131f
C26390 VDD.n7239 VSS 0.012131f
C26391 VDD.n7240 VSS 0.012131f
C26392 VDD.n7241 VSS 0.012131f
C26393 VDD.n7242 VSS 0.012131f
C26394 VDD.n7243 VSS 0.012131f
C26395 VDD.n7244 VSS 0.012131f
C26396 VDD.n7245 VSS 0.012131f
C26397 VDD.n7246 VSS 0.012131f
C26398 VDD.n7247 VSS 0.012131f
C26399 VDD.n7248 VSS 0.012131f
C26400 VDD.n7249 VSS 0.012131f
C26401 VDD.n7250 VSS 0.012131f
C26402 VDD.n7251 VSS 0.012131f
C26403 VDD.n7252 VSS 0.012131f
C26404 VDD.n7253 VSS 0.012131f
C26405 VDD.n7254 VSS 0.012131f
C26406 VDD.n7255 VSS 0.012131f
C26407 VDD.n7256 VSS 0.012131f
C26408 VDD.n7257 VSS 0.012131f
C26409 VDD.n7258 VSS 0.012131f
C26410 VDD.n7259 VSS 0.012131f
C26411 VDD.n7260 VSS 0.012131f
C26412 VDD.n7261 VSS 0.012131f
C26413 VDD.n7262 VSS 0.012131f
C26414 VDD.n7263 VSS 0.012131f
C26415 VDD.n7264 VSS 0.012131f
C26416 VDD.n7265 VSS 0.012131f
C26417 VDD.n7266 VSS 0.012131f
C26418 VDD.n7267 VSS 0.012131f
C26419 VDD.n7268 VSS 0.012131f
C26420 VDD.n7269 VSS 0.012131f
C26421 VDD.n7270 VSS 0.012131f
C26422 VDD.n7271 VSS 0.012131f
C26423 VDD.n7272 VSS 0.012131f
C26424 VDD.n7273 VSS 0.012131f
C26425 VDD.n7274 VSS 0.012131f
C26426 VDD.n7275 VSS 0.012131f
C26427 VDD.n7276 VSS 0.012131f
C26428 VDD.n7277 VSS 0.012131f
C26429 VDD.n7278 VSS 0.012131f
C26430 VDD.n7279 VSS 0.012131f
C26431 VDD.n7280 VSS 0.012131f
C26432 VDD.n7281 VSS 0.012131f
C26433 VDD.n7282 VSS 0.012131f
C26434 VDD.n7283 VSS 0.012131f
C26435 VDD.n7284 VSS 0.012131f
C26436 VDD.n7285 VSS 0.012131f
C26437 VDD.n7286 VSS 0.012131f
C26438 VDD.n7287 VSS 0.012131f
C26439 VDD.n7288 VSS 0.012131f
C26440 VDD.n7289 VSS 0.012131f
C26441 VDD.n7290 VSS 0.012131f
C26442 VDD.n7291 VSS 0.012131f
C26443 VDD.n7292 VSS 0.012131f
C26444 VDD.n7293 VSS 0.012131f
C26445 VDD.n7294 VSS 0.012131f
C26446 VDD.n7295 VSS 0.012131f
C26447 VDD.n7296 VSS 0.012131f
C26448 VDD.n7297 VSS 0.012131f
C26449 VDD.n7298 VSS 0.012131f
C26450 VDD.n7299 VSS 0.012131f
C26451 VDD.n7300 VSS 0.012131f
C26452 VDD.n7301 VSS 0.012131f
C26453 VDD.n7302 VSS 0.084561f
C26454 VDD.n7303 VSS 0.012131f
C26455 VDD.n7304 VSS 0.106951f
C26456 VDD.n7305 VSS 0.106951f
C26457 VDD.n7306 VSS 0.012131f
C26458 VDD.n7307 VSS 0.012131f
C26459 VDD.n7308 VSS 0.012131f
C26460 VDD.n7309 VSS 0.011263f
C26461 VDD.n7310 VSS 0.012131f
C26462 VDD.n7311 VSS 0.012131f
C26463 VDD.n7312 VSS 0.012131f
C26464 VDD.n7313 VSS 0.012131f
C26465 VDD.n7314 VSS 0.012131f
C26466 VDD.n7315 VSS 0.012131f
C26467 VDD.n7316 VSS 0.012131f
C26468 VDD.n7317 VSS 0.012131f
C26469 VDD.n7318 VSS 0.012131f
C26470 VDD.n7319 VSS 0.012131f
C26471 VDD.n7320 VSS 0.012131f
C26472 VDD.n7321 VSS 0.012131f
C26473 VDD.n7322 VSS 0.012131f
C26474 VDD.n7323 VSS 0.012131f
C26475 VDD.n7324 VSS 0.012131f
C26476 VDD.n7325 VSS 0.012131f
C26477 VDD.n7326 VSS 0.012131f
C26478 VDD.n7327 VSS 0.012131f
C26479 VDD.n7328 VSS 0.012131f
C26480 VDD.n7329 VSS 0.012131f
C26481 VDD.n7330 VSS 0.012131f
C26482 VDD.n7331 VSS 0.012131f
C26483 VDD.n7332 VSS 0.012131f
C26484 VDD.n7333 VSS 0.012131f
C26485 VDD.n7334 VSS 0.012131f
C26486 VDD.n7335 VSS 0.012131f
C26487 VDD.n7336 VSS 0.012131f
C26488 VDD.n7337 VSS 0.012131f
C26489 VDD.n7338 VSS 0.012131f
C26490 VDD.n7339 VSS 0.012131f
C26491 VDD.n7340 VSS 0.012131f
C26492 VDD.n7341 VSS 0.012131f
C26493 VDD.n7342 VSS 0.012131f
C26494 VDD.n7343 VSS 0.012131f
C26495 VDD.n7344 VSS 0.012131f
C26496 VDD.n7345 VSS 0.012131f
C26497 VDD.n7346 VSS 0.012131f
C26498 VDD.n7347 VSS 0.012131f
C26499 VDD.n7348 VSS 0.012131f
C26500 VDD.n7349 VSS 0.012131f
C26501 VDD.n7350 VSS 0.012131f
C26502 VDD.n7351 VSS 0.012131f
C26503 VDD.n7352 VSS 0.012131f
C26504 VDD.n7353 VSS 0.012131f
C26505 VDD.n7354 VSS 0.012131f
C26506 VDD.n7355 VSS 0.012131f
C26507 VDD.n7356 VSS 0.012131f
C26508 VDD.n7357 VSS 0.012131f
C26509 VDD.n7358 VSS 0.012131f
C26510 VDD.n7359 VSS 0.012131f
C26511 VDD.n7360 VSS 0.012131f
C26512 VDD.n7361 VSS 0.012131f
C26513 VDD.n7362 VSS 0.012131f
C26514 VDD.n7363 VSS 0.012131f
C26515 VDD.n7364 VSS 0.012131f
C26516 VDD.n7365 VSS 0.012131f
C26517 VDD.n7366 VSS 0.012131f
C26518 VDD.n7367 VSS 0.012131f
C26519 VDD.n7368 VSS 0.012131f
C26520 VDD.n7369 VSS 0.012131f
C26521 VDD.n7370 VSS 0.012131f
C26522 VDD.n7371 VSS 0.012131f
C26523 VDD.n7372 VSS 0.012131f
C26524 VDD.n7373 VSS 0.012131f
C26525 VDD.n7374 VSS 0.012131f
C26526 VDD.n7375 VSS 0.012131f
C26527 VDD.n7376 VSS 0.012131f
C26528 VDD.n7377 VSS 0.012131f
C26529 VDD.n7378 VSS 0.012131f
C26530 VDD.n7379 VSS 0.012131f
C26531 VDD.n7380 VSS 0.012131f
C26532 VDD.n7381 VSS 0.012131f
C26533 VDD.n7382 VSS 0.012131f
C26534 VDD.n7383 VSS 0.012131f
C26535 VDD.n7384 VSS 0.012131f
C26536 VDD.n7385 VSS 0.012131f
C26537 VDD.n7386 VSS 0.012131f
C26538 VDD.n7387 VSS 0.012131f
C26539 VDD.n7388 VSS 0.012131f
C26540 VDD.n7389 VSS 0.012131f
C26541 VDD.n7390 VSS 0.012131f
C26542 VDD.n7391 VSS 0.012131f
C26543 VDD.n7392 VSS 0.012131f
C26544 VDD.n7393 VSS 0.012131f
C26545 VDD.n7394 VSS 0.012131f
C26546 VDD.n7395 VSS 0.012131f
C26547 VDD.n7396 VSS 0.012131f
C26548 VDD.n7397 VSS 0.012131f
C26549 VDD.n7398 VSS 0.012131f
C26550 VDD.n7399 VSS 0.012131f
C26551 VDD.n7400 VSS 0.012131f
C26552 VDD.n7401 VSS 0.012131f
C26553 VDD.n7402 VSS 0.012131f
C26554 VDD.n7403 VSS 0.012131f
C26555 VDD.n7404 VSS 0.012131f
C26556 VDD.n7405 VSS 0.012131f
C26557 VDD.n7406 VSS 0.012131f
C26558 VDD.n7407 VSS 0.012131f
C26559 VDD.n7408 VSS 0.012131f
C26560 VDD.n7409 VSS 0.012131f
C26561 VDD.n7410 VSS 0.012131f
C26562 VDD.n7411 VSS 0.012131f
C26563 VDD.n7412 VSS 0.012131f
C26564 VDD.n7413 VSS 0.012131f
C26565 VDD.n7414 VSS 0.012131f
C26566 VDD.n7415 VSS 0.012131f
C26567 VDD.n7416 VSS 0.012131f
C26568 VDD.n7417 VSS 0.012131f
C26569 VDD.n7418 VSS 0.012131f
C26570 VDD.n7419 VSS 0.012131f
C26571 VDD.n7420 VSS 0.012131f
C26572 VDD.n7421 VSS 0.012131f
C26573 VDD.n7422 VSS 0.012131f
C26574 VDD.n7423 VSS 0.012131f
C26575 VDD.n7424 VSS 0.012131f
C26576 VDD.n7425 VSS 0.012131f
C26577 VDD.n7426 VSS 0.012131f
C26578 VDD.n7427 VSS 0.012131f
C26579 VDD.n7428 VSS 0.012131f
C26580 VDD.n7429 VSS 0.012131f
C26581 VDD.n7430 VSS 0.012131f
C26582 VDD.n7431 VSS 0.012131f
C26583 VDD.n7432 VSS 0.012131f
C26584 VDD.n7433 VSS 0.012131f
C26585 VDD.n7434 VSS 0.012131f
C26586 VDD.n7435 VSS 0.012131f
C26587 VDD.n7436 VSS 0.012131f
C26588 VDD.n7437 VSS 0.012131f
C26589 VDD.n7438 VSS 0.012131f
C26590 VDD.n7439 VSS 0.012131f
C26591 VDD.n7440 VSS 0.012131f
C26592 VDD.n7441 VSS 0.012131f
C26593 VDD.n7442 VSS 0.012131f
C26594 VDD.n7443 VSS 0.012131f
C26595 VDD.n7444 VSS 0.012131f
C26596 VDD.n7445 VSS 0.012131f
C26597 VDD.n7446 VSS 0.012131f
C26598 VDD.n7447 VSS 0.012131f
C26599 VDD.n7448 VSS 0.012131f
C26600 VDD.n7449 VSS 0.012131f
C26601 VDD.n7450 VSS 0.012131f
C26602 VDD.n7451 VSS 0.012131f
C26603 VDD.n7452 VSS 0.012131f
C26604 VDD.n7453 VSS 0.012131f
C26605 VDD.n7454 VSS 0.012131f
C26606 VDD.n7455 VSS 0.012131f
C26607 VDD.n7456 VSS 0.012131f
C26608 VDD.n7457 VSS 0.012131f
C26609 VDD.n7458 VSS 0.012131f
C26610 VDD.n7459 VSS 0.012131f
C26611 VDD.n7460 VSS 0.012131f
C26612 VDD.n7461 VSS 0.012131f
C26613 VDD.n7462 VSS 0.012131f
C26614 VDD.n7463 VSS 0.012131f
C26615 VDD.n7464 VSS 0.012131f
C26616 VDD.n7465 VSS 0.012131f
C26617 VDD.n7466 VSS 0.012131f
C26618 VDD.n7467 VSS 0.012131f
C26619 VDD.n7468 VSS 0.012131f
C26620 VDD.n7469 VSS 0.012131f
C26621 VDD.n7470 VSS 0.012131f
C26622 VDD.n7471 VSS 0.012131f
C26623 VDD.n7472 VSS 0.012131f
C26624 VDD.n7473 VSS 0.012131f
C26625 VDD.n7474 VSS 0.012131f
C26626 VDD.n7475 VSS 0.012131f
C26627 VDD.n7476 VSS 0.012131f
C26628 VDD.n7477 VSS 0.012131f
C26629 VDD.n7478 VSS 0.012131f
C26630 VDD.n7479 VSS 0.012131f
C26631 VDD.n7480 VSS 0.012131f
C26632 VDD.n7481 VSS 0.012131f
C26633 VDD.n7482 VSS 0.012131f
C26634 VDD.n7483 VSS 0.012131f
C26635 VDD.n7484 VSS 0.012131f
C26636 VDD.n7485 VSS 0.012131f
C26637 VDD.n7486 VSS 0.012131f
C26638 VDD.n7487 VSS 0.012131f
C26639 VDD.n7488 VSS 0.012131f
C26640 VDD.n7489 VSS 0.012131f
C26641 VDD.n7490 VSS 0.012131f
C26642 VDD.n7491 VSS 0.012131f
C26643 VDD.n7492 VSS 0.012131f
C26644 VDD.n7493 VSS 0.012131f
C26645 VDD.n7494 VSS 0.012131f
C26646 VDD.n7495 VSS 0.012131f
C26647 VDD.n7496 VSS 0.012131f
C26648 VDD.n7497 VSS 0.012131f
C26649 VDD.n7498 VSS 0.012131f
C26650 VDD.n7499 VSS 0.012131f
C26651 VDD.n7500 VSS 0.012131f
C26652 VDD.n7501 VSS 0.012131f
C26653 VDD.n7502 VSS 0.012131f
C26654 VDD.n7503 VSS 0.012131f
C26655 VDD.n7504 VSS 0.012131f
C26656 VDD.n7505 VSS 0.012131f
C26657 VDD.n7506 VSS 0.012131f
C26658 VDD.n7507 VSS 0.012131f
C26659 VDD.n7508 VSS 0.012131f
C26660 VDD.n7509 VSS 0.012131f
C26661 VDD.n7510 VSS 0.012131f
C26662 VDD.n7511 VSS 0.012131f
C26663 VDD.n7512 VSS 0.012131f
C26664 VDD.n7513 VSS 0.012131f
C26665 VDD.n7514 VSS 0.012131f
C26666 VDD.n7515 VSS 0.012131f
C26667 VDD.n7516 VSS 0.012131f
C26668 VDD.n7517 VSS 0.012131f
C26669 VDD.n7518 VSS 0.012131f
C26670 VDD.n7519 VSS 0.012131f
C26671 VDD.n7520 VSS 0.012131f
C26672 VDD.n7521 VSS 0.012131f
C26673 VDD.n7522 VSS 0.012131f
C26674 VDD.n7523 VSS 0.012131f
C26675 VDD.n7524 VSS 0.012131f
C26676 VDD.n7525 VSS 0.012131f
C26677 VDD.n7526 VSS 0.012131f
C26678 VDD.n7527 VSS 0.012131f
C26679 VDD.n7528 VSS 0.012131f
C26680 VDD.n7529 VSS 0.012131f
C26681 VDD.n7530 VSS 0.012131f
C26682 VDD.n7531 VSS 0.012131f
C26683 VDD.n7532 VSS 0.012131f
C26684 VDD.n7533 VSS 0.012131f
C26685 VDD.n7534 VSS 0.012131f
C26686 VDD.n7535 VSS 0.012131f
C26687 VDD.n7536 VSS 0.012131f
C26688 VDD.n7537 VSS 0.012131f
C26689 VDD.n7538 VSS 0.012131f
C26690 VDD.n7539 VSS 0.012131f
C26691 VDD.n7540 VSS 0.012131f
C26692 VDD.n7541 VSS 0.012131f
C26693 VDD.n7542 VSS 0.012131f
C26694 VDD.n7543 VSS 0.012131f
C26695 VDD.n7544 VSS 0.012131f
C26696 VDD.n7545 VSS 0.012131f
C26697 VDD.n7546 VSS 0.012131f
C26698 VDD.n7547 VSS 0.012131f
C26699 VDD.n7548 VSS 0.012131f
C26700 VDD.n7549 VSS 0.012131f
C26701 VDD.n7550 VSS 0.012131f
C26702 VDD.n7551 VSS 0.012131f
C26703 VDD.n7552 VSS 0.012131f
C26704 VDD.n7553 VSS 0.012131f
C26705 VDD.n7554 VSS 0.012131f
C26706 VDD.n7555 VSS 0.012131f
C26707 VDD.n7556 VSS 0.012131f
C26708 VDD.n7557 VSS 0.012131f
C26709 VDD.n7558 VSS 0.012131f
C26710 VDD.n7559 VSS 0.012131f
C26711 VDD.n7560 VSS 0.012131f
C26712 VDD.n7561 VSS 0.012131f
C26713 VDD.n7562 VSS 0.012131f
C26714 VDD.n7563 VSS 0.012131f
C26715 VDD.n7564 VSS 0.012131f
C26716 VDD.n7565 VSS 0.012131f
C26717 VDD.n7566 VSS 0.012131f
C26718 VDD.n7567 VSS 0.012131f
C26719 VDD.n7568 VSS 0.012131f
C26720 VDD.n7569 VSS 0.012131f
C26721 VDD.n7570 VSS 0.012131f
C26722 VDD.n7571 VSS 0.012131f
C26723 VDD.n7572 VSS 0.012131f
C26724 VDD.n7573 VSS 0.012131f
C26725 VDD.n7574 VSS 0.012131f
C26726 VDD.n7575 VSS 0.012131f
C26727 VDD.n7576 VSS 0.012131f
C26728 VDD.n7577 VSS 0.012131f
C26729 VDD.n7578 VSS 0.012131f
C26730 VDD.n7579 VSS 0.012131f
C26731 VDD.n7580 VSS 0.012131f
C26732 VDD.n7581 VSS 0.012131f
C26733 VDD.n7582 VSS 0.012131f
C26734 VDD.n7583 VSS 0.012131f
C26735 VDD.n7584 VSS 0.012131f
C26736 VDD.n7585 VSS 0.012131f
C26737 VDD.n7586 VSS 0.012131f
C26738 VDD.n7587 VSS 0.012131f
C26739 VDD.n7588 VSS 0.012131f
C26740 VDD.n7589 VSS 0.012131f
C26741 VDD.n7590 VSS 0.012131f
C26742 VDD.n7591 VSS 0.012131f
C26743 VDD.n7592 VSS 0.012131f
C26744 VDD.n7593 VSS 0.012131f
C26745 VDD.n7594 VSS 0.012131f
C26746 VDD.n7595 VSS 0.012131f
C26747 VDD.n7596 VSS 0.012131f
C26748 VDD.n7597 VSS 0.012131f
C26749 VDD.n7598 VSS 0.012131f
C26750 VDD.n7599 VSS 0.012131f
C26751 VDD.n7600 VSS 0.012131f
C26752 VDD.n7601 VSS 0.012131f
C26753 VDD.n7602 VSS 0.012131f
C26754 VDD.n7603 VSS 0.012131f
C26755 VDD.n7604 VSS 0.012131f
C26756 VDD.n7605 VSS 0.012131f
C26757 VDD.n7606 VSS 0.012131f
C26758 VDD.n7607 VSS 0.012131f
C26759 VDD.n7608 VSS 0.012131f
C26760 VDD.n7609 VSS 0.012131f
C26761 VDD.n7610 VSS 0.012131f
C26762 VDD.n7611 VSS 0.012131f
C26763 VDD.n7612 VSS 0.012131f
C26764 VDD.n7613 VSS 0.012131f
C26765 VDD.n7614 VSS 0.012131f
C26766 VDD.n7615 VSS 0.012131f
C26767 VDD.n7616 VSS 0.012131f
C26768 VDD.n7617 VSS 0.012131f
C26769 VDD.n7618 VSS 0.012131f
C26770 VDD.n7619 VSS 0.012131f
C26771 VDD.n7620 VSS 0.012131f
C26772 VDD.n7621 VSS 0.012131f
C26773 VDD.n7622 VSS 0.012131f
C26774 VDD.n7623 VSS 0.012131f
C26775 VDD.n7624 VSS 0.012131f
C26776 VDD.n7625 VSS 0.012131f
C26777 VDD.n7626 VSS 0.012131f
C26778 VDD.n7627 VSS 0.012131f
C26779 VDD.n7628 VSS 0.012131f
C26780 VDD.n7629 VSS 0.012131f
C26781 VDD.n7630 VSS 0.012131f
C26782 VDD.n7631 VSS 0.012131f
C26783 VDD.n7632 VSS 0.012131f
C26784 VDD.n7633 VSS 0.012131f
C26785 VDD.n7634 VSS 0.012131f
C26786 VDD.n7635 VSS 0.012131f
C26787 VDD.n7636 VSS 0.012131f
C26788 VDD.n7637 VSS 0.012131f
C26789 VDD.n7638 VSS 0.012131f
C26790 VDD.n7639 VSS 0.012131f
C26791 VDD.n7640 VSS 0.012131f
C26792 VDD.n7641 VSS 0.012131f
C26793 VDD.n7642 VSS 0.012131f
C26794 VDD.n7643 VSS 0.012131f
C26795 VDD.n7644 VSS 0.012131f
C26796 VDD.n7645 VSS 0.012131f
C26797 VDD.n7646 VSS 0.012131f
C26798 VDD.n7647 VSS 0.012131f
C26799 VDD.n7648 VSS 0.012131f
C26800 VDD.n7649 VSS 0.012131f
C26801 VDD.n7650 VSS 0.012131f
C26802 VDD.n7651 VSS 0.012131f
C26803 VDD.n7652 VSS 0.012131f
C26804 VDD.n7653 VSS 0.012131f
C26805 VDD.n7654 VSS 0.012131f
C26806 VDD.n7655 VSS 0.012131f
C26807 VDD.n7656 VSS 0.012131f
C26808 VDD.n7657 VSS 0.012131f
C26809 VDD.n7658 VSS 0.012131f
C26810 VDD.n7659 VSS 0.012131f
C26811 VDD.n7660 VSS 0.012131f
C26812 VDD.n7661 VSS 0.012131f
C26813 VDD.n7662 VSS 0.012131f
C26814 VDD.n7663 VSS 0.012131f
C26815 VDD.n7664 VSS 0.012131f
C26816 VDD.n7665 VSS 0.012131f
C26817 VDD.n7666 VSS 0.012131f
C26818 VDD.n7667 VSS 0.012131f
C26819 VDD.n7668 VSS 0.012131f
C26820 VDD.n7669 VSS 0.012131f
C26821 VDD.n7670 VSS 0.012131f
C26822 VDD.n7671 VSS 0.012131f
C26823 VDD.n7672 VSS 0.012131f
C26824 VDD.n7673 VSS 0.012131f
C26825 VDD.n7674 VSS 0.012131f
C26826 VDD.n7675 VSS 0.012131f
C26827 VDD.n7676 VSS 0.012131f
C26828 VDD.n7677 VSS 0.012131f
C26829 VDD.n7678 VSS 0.012131f
C26830 VDD.n7679 VSS 0.012131f
C26831 VDD.n7680 VSS 0.012131f
C26832 VDD.n7681 VSS 0.012131f
C26833 VDD.n7682 VSS 0.010414f
C26834 VDD.n7683 VSS 0.104583f
C26835 VDD.n7684 VSS 0.099571f
C26836 VDD.n7685 VSS 0.012131f
C26837 VDD.n7686 VSS 0.012131f
C26838 VDD.n7687 VSS 0.197913f
C26839 VDD.n7688 VSS 0.260606f
C26840 VDD.n7689 VSS 0.16841f
C26841 VDD.n7690 VSS 0.012131f
C26842 VDD.n7691 VSS 0.012131f
C26843 VDD.n7692 VSS 0.012131f
C26844 VDD.n7693 VSS 0.260606f
C26845 VDD.n7694 VSS 0.260606f
C26846 VDD.n7695 VSS 0.260606f
C26847 VDD.n7696 VSS 0.012131f
C26848 VDD.n7697 VSS 0.012131f
C26849 VDD.n7698 VSS 0.012131f
C26850 VDD.n7699 VSS 0.231103f
C26851 VDD.n7700 VSS 0.130303f
C26852 VDD.n7701 VSS 0.159805f
C26853 VDD.n7702 VSS 0.260606f
C26854 VDD.n7703 VSS 0.012131f
C26855 VDD.n7704 VSS 0.012131f
C26856 VDD.n7705 VSS 0.012131f
C26857 VDD.n7706 VSS 0.260606f
C26858 VDD.n7707 VSS 0.260606f
C26859 VDD.n7708 VSS 0.183161f
C26860 VDD.n7709 VSS 0.012131f
C26861 VDD.n7710 VSS 0.012131f
C26862 VDD.n7711 VSS 0.207747f
C26863 VDD.n7712 VSS 0.260606f
C26864 VDD.n7713 VSS 0.158576f
C26865 VDD.n7714 VSS 0.012131f
C26866 VDD.n7715 VSS 0.012131f
C26867 VDD.n7716 VSS 0.012131f
C26868 VDD.n7717 VSS 0.260606f
C26869 VDD.n7718 VSS 0.247084f
C26870 VDD.t2828 VSS 0.066856f
C26871 VDD.n7719 VSS 0.154235f
C26872 VDD.n7720 VSS 0.143825f
C26873 VDD.n7721 VSS 0.012131f
C26874 VDD.n7722 VSS 0.012131f
C26875 VDD.n7723 VSS 0.012131f
C26876 VDD.n7724 VSS 0.222498f
C26877 VDD.n7725 VSS 0.145708f
C26878 VDD.n7726 VSS 0.16841f
C26879 VDD.n7727 VSS 0.260606f
C26880 VDD.n7728 VSS 0.012131f
C26881 VDD.n7729 VSS 0.012131f
C26882 VDD.n7730 VSS 0.012131f
C26883 VDD.n7731 VSS 0.260606f
C26884 VDD.n7732 VSS 0.260606f
C26885 VDD.n7733 VSS 0.260606f
C26886 VDD.n7734 VSS 0.012131f
C26887 VDD.n7735 VSS 0.012131f
C26888 VDD.n7736 VSS 0.012131f
C26889 VDD.n7737 VSS 0.260606f
C26890 VDD.n7738 VSS 0.260606f
C26891 VDD.n7739 VSS 0.156118f
C26892 VDD.n7740 VSS 0.012131f
C26893 VDD.n7741 VSS 0.012131f
C26894 VDD.n7742 VSS 0.234791f
C26895 VDD.n7743 VSS 0.260606f
C26896 VDD.n7744 VSS 0.131532f
C26897 VDD.n7745 VSS 0.012131f
C26898 VDD.n7746 VSS 0.012131f
C26899 VDD.n7747 VSS 0.259376f
C26900 VDD.n7748 VSS 0.260606f
C26901 VDD.n7749 VSS 0.260606f
C26902 VDD.n7750 VSS 0.012131f
C26903 VDD.n7751 VSS 0.012131f
C26904 VDD.n7752 VSS 0.012131f
C26905 VDD.n7753 VSS 0.260606f
C26906 VDD.n7754 VSS 0.260606f
C26907 VDD.n7755 VSS 0.260606f
C26908 VDD.n7756 VSS 0.012131f
C26909 VDD.n7757 VSS 0.012131f
C26910 VDD.n7758 VSS 0.012131f
C26911 VDD.n7759 VSS 0.208976f
C26912 VDD.n7760 VSS 0.316821f
C26913 VDD.n7761 VSS 0.181932f
C26914 VDD.n7762 VSS 0.260606f
C26915 VDD.n7763 VSS 0.012131f
C26916 VDD.n7764 VSS 0.012131f
C26917 VDD.n7765 VSS 0.012131f
C26918 VDD.n7766 VSS 0.260606f
C26919 VDD.n7767 VSS 0.260606f
C26920 VDD.n7768 VSS 0.260606f
C26921 VDD.n7769 VSS 0.012131f
C26922 VDD.n7770 VSS 0.012131f
C26923 VDD.n7771 VSS 0.012131f
C26924 VDD.n7772 VSS 0.260606f
C26925 VDD.n7773 VSS 0.260606f
C26926 VDD.n7774 VSS 0.157347f
C26927 VDD.n7775 VSS 0.012131f
C26928 VDD.n7776 VSS 0.012131f
C26929 VDD.n7777 VSS 0.012131f
C26930 VDD.n7778 VSS 0.260606f
C26931 VDD.n7779 VSS 0.132761f
C26932 VDD.t1081 VSS 0.066856f
C26933 VDD.n7780 VSS 0.154235f
C26934 VDD.n7781 VSS 0.258147f
C26935 VDD.n7782 VSS 0.012131f
C26936 VDD.n7783 VSS 0.012131f
C26937 VDD.n7784 VSS 0.012131f
C26938 VDD.n7785 VSS 0.260606f
C26939 VDD.n7786 VSS 0.260606f
C26940 VDD.n7787 VSS 0.260606f
C26941 VDD.n7788 VSS 0.012131f
C26942 VDD.n7789 VSS 0.012131f
C26943 VDD.n7790 VSS 0.012131f
C26944 VDD.n7791 VSS 0.260606f
C26945 VDD.n7792 VSS 0.260606f
C26946 VDD.n7793 VSS 0.196683f
C26947 VDD.n7794 VSS 0.012131f
C26948 VDD.n7795 VSS 0.012131f
C26949 VDD.n7796 VSS 0.194225f
C26950 VDD.n7797 VSS 0.260606f
C26951 VDD.n7798 VSS 0.172098f
C26952 VDD.n7799 VSS 0.012131f
C26953 VDD.n7800 VSS 0.012131f
C26954 VDD.n7801 VSS 0.21881f
C26955 VDD.n7802 VSS 0.260606f
C26956 VDD.n7803 VSS 0.260606f
C26957 VDD.n7804 VSS 0.012131f
C26958 VDD.n7805 VSS 0.012131f
C26959 VDD.n7806 VSS 0.012131f
C26960 VDD.n7807 VSS 0.260606f
C26961 VDD.n7808 VSS 0.23602f
C26962 VDD.n7809 VSS 0.145708f
C26963 VDD.n7810 VSS 0.154888f
C26964 VDD.n7811 VSS 0.012131f
C26965 VDD.n7812 VSS 0.012131f
C26966 VDD.n7813 VSS 0.012131f
C26967 VDD.n7814 VSS 0.260606f
C26968 VDD.n7815 VSS 0.260606f
C26969 VDD.n7816 VSS 0.260606f
C26970 VDD.n7817 VSS 0.012131f
C26971 VDD.n7818 VSS 0.012131f
C26972 VDD.n7819 VSS 0.012131f
C26973 VDD.n7820 VSS 0.16841f
C26974 VDD.n7821 VSS 0.089737f
C26975 VDD.n7822 VSS 0.167314f
C26976 VDD.n7823 VSS 0.190302f
C26977 VDD.t1664 VSS 0.066856f
C26978 VDD.n7824 VSS 0.164998f
C26979 VDD.t2054 VSS 0.066856f
C26980 VDD.n7825 VSS 0.164998f
C26981 VDD.n7826 VSS 0.274982f
C26982 VDD.n7827 VSS 0.501023f
C26983 VDD.n7828 VSS 0.274982f
C26984 VDD.t596 VSS 0.066856f
C26985 VDD.n7829 VSS 0.164998f
C26986 VDD.t1011 VSS 0.066856f
C26987 VDD.n7830 VSS 0.164998f
C26988 VDD.n7831 VSS 0.217367f
C26989 VDD.n7832 VSS 0.263268f
C26990 VDD.n7833 VSS 0.283088f
C26991 VDD.n7834 VSS 4.4125f
C26992 VDD.n7835 VSS 0.283088f
C26993 VDD.n7836 VSS 0.263268f
C26994 VDD.t2246 VSS 0.034186f
C26995 VDD.n7837 VSS 0.217367f
C26996 VDD.t2245 VSS 0.066856f
C26997 VDD.n7838 VSS 0.164998f
C26998 VDD.t1836 VSS 0.066856f
C26999 VDD.n7839 VSS 0.164998f
C27000 VDD.t1837 VSS 0.034186f
C27001 VDD.n7840 VSS 0.282774f
C27002 VDD.t3711 VSS 0.066856f
C27003 VDD.n7841 VSS 0.291301f
C27004 VDD.t3712 VSS 0.034186f
C27005 VDD.n7842 VSS 0.280015f
C27006 VDD.n7843 VSS 0.147799f
C27007 VDD.t4466 VSS 0.066856f
C27008 VDD.n7844 VSS 0.129831f
C27009 VDD.n7845 VSS 0.105899f
C27010 VDD.n7846 VSS 0.016021f
C27011 VDD.t1205 VSS 0.016021f
C27012 VDD.n7847 VSS 0.016021f
C27013 VDD.t2695 VSS 0.016021f
C27014 VDD.n7848 VSS 0.016021f
C27015 VDD.n7849 VSS 0.248157f
C27016 VDD.n7850 VSS 0.25586f
C27017 VDD.t2786 VSS 0.034186f
C27018 VDD.n7851 VSS 0.25586f
C27019 VDD.t2694 VSS 0.066856f
C27020 VDD.n7852 VSS 0.182089f
C27021 VDD.n7853 VSS 0.311521f
C27022 VDD.t1398 VSS 0.034186f
C27023 VDD.t3987 VSS 0.034186f
C27024 VDD.t2338 VSS 0.066856f
C27025 VDD.n7854 VSS 0.154441f
C27026 VDD.n7855 VSS 0.00473f
C27027 VDD.n7856 VSS 0.00473f
C27028 VDD.n7857 VSS 0.00473f
C27029 VDD.n7858 VSS 0.00473f
C27030 VDD.n7859 VSS 0.00473f
C27031 VDD.n7860 VSS 0.00473f
C27032 VDD.t1383 VSS 0.066856f
C27033 VDD.n7861 VSS 0.164014f
C27034 VDD.t3966 VSS 0.066856f
C27035 VDD.n7862 VSS 0.164014f
C27036 VDD.t3967 VSS 0.034186f
C27037 VDD.n7863 VSS 0.14612f
C27038 VDD.t2308 VSS 0.034186f
C27039 VDD.n7864 VSS 0.116748f
C27040 VDD.n7865 VSS 0.00473f
C27041 VDD.t245 VSS 0.008011f
C27042 VDD.t49 VSS 0.008011f
C27043 VDD.n7866 VSS 0.018711f
C27044 VDD.n7867 VSS 0.017079f
C27045 VDD.t75 VSS 0.008011f
C27046 VDD.t134 VSS 0.008011f
C27047 VDD.n7868 VSS 0.020036f
C27048 VDD.n7869 VSS 0.00473f
C27049 VDD.t224 VSS 0.008011f
C27050 VDD.t269 VSS 0.008011f
C27051 VDD.n7870 VSS 0.018711f
C27052 VDD.n7871 VSS 0.017079f
C27053 VDD.t280 VSS 0.008011f
C27054 VDD.t105 VSS 0.008011f
C27055 VDD.n7872 VSS 0.020036f
C27056 VDD.n7873 VSS 0.00473f
C27057 VDD.t34 VSS 0.019712f
C27058 VDD.n7874 VSS 0.024851f
C27059 VDD.t31 VSS 0.020856f
C27060 VDD.n7875 VSS 0.00473f
C27061 VDD.t27 VSS 0.008011f
C27062 VDD.t18 VSS 0.008011f
C27063 VDD.n7876 VSS 0.018711f
C27064 VDD.n7877 VSS 0.017079f
C27065 VDD.t45 VSS 0.008011f
C27066 VDD.t39 VSS 0.008011f
C27067 VDD.n7878 VSS 0.020036f
C27068 VDD.n7879 VSS 0.00473f
C27069 VDD.t112 VSS 0.008011f
C27070 VDD.t188 VSS 0.008011f
C27071 VDD.n7880 VSS 0.018711f
C27072 VDD.n7881 VSS 0.017079f
C27073 VDD.t175 VSS 0.008011f
C27074 VDD.t251 VSS 0.008011f
C27075 VDD.n7882 VSS 0.020036f
C27076 VDD.n7883 VSS 0.00473f
C27077 VDD.t259 VSS 0.008011f
C27078 VDD.t101 VSS 0.008011f
C27079 VDD.n7884 VSS 0.018711f
C27080 VDD.n7885 VSS 0.017079f
C27081 VDD.t90 VSS 0.008011f
C27082 VDD.t168 VSS 0.008011f
C27083 VDD.n7886 VSS 0.020036f
C27084 VDD.t2339 VSS 0.034186f
C27085 VDD.n7887 VSS 0.157262f
C27086 VDD.t1120 VSS 0.034186f
C27087 VDD.n7888 VSS 0.172056f
C27088 VDD.n7889 VSS 0.110446f
C27089 VDD.n7890 VSS 0.105916f
C27090 VDD.n7891 VSS 0.034447f
C27091 VDD.n7892 VSS 0.029907f
C27092 VDD.n7893 VSS 0.019376f
C27093 VDD.n7894 VSS 0.019381f
C27094 VDD.n7895 VSS 0.029907f
C27095 VDD.n7896 VSS 0.024526f
C27096 VDD.n7897 VSS 0.024531f
C27097 VDD.n7898 VSS 0.029907f
C27098 VDD.n7899 VSS 0.019376f
C27099 VDD.n7900 VSS 0.019381f
C27100 VDD.n7901 VSS 0.03786f
C27101 VDD.n7902 VSS 0.013692f
C27102 VDD.n7903 VSS 0.013697f
C27103 VDD.n7904 VSS 0.029907f
C27104 VDD.n7905 VSS 0.019376f
C27105 VDD.n7906 VSS 0.019381f
C27106 VDD.n7907 VSS 0.029907f
C27107 VDD.n7908 VSS 0.03416f
C27108 VDD.n7909 VSS 0.106152f
C27109 VDD.n7910 VSS 0.15793f
C27110 VDD.t2307 VSS 0.066856f
C27111 VDD.n7911 VSS 0.155055f
C27112 VDD.n7912 VSS 0.150553f
C27113 VDD.n7913 VSS 0.034182f
C27114 VDD.t156 VSS 0.008011f
C27115 VDD.t205 VSS 0.008011f
C27116 VDD.n7914 VSS 0.018207f
C27117 VDD.n7915 VSS 0.015517f
C27118 VDD.n7916 VSS 0.010511f
C27119 VDD.n7917 VSS 0.019382f
C27120 VDD.n7918 VSS 0.019375f
C27121 VDD.t131 VSS 0.008011f
C27122 VDD.t178 VSS 0.008011f
C27123 VDD.n7919 VSS 0.018207f
C27124 VDD.n7920 VSS 0.015517f
C27125 VDD.n7921 VSS 0.010511f
C27126 VDD.n7922 VSS 0.013698f
C27127 VDD.n7923 VSS 0.013691f
C27128 VDD.t60 VSS 0.019268f
C27129 VDD.n7924 VSS 0.02323f
C27130 VDD.n7925 VSS 0.010511f
C27131 VDD.n7926 VSS 0.019382f
C27132 VDD.n7927 VSS 0.019375f
C27133 VDD.t152 VSS 0.008011f
C27134 VDD.t197 VSS 0.008011f
C27135 VDD.n7928 VSS 0.018207f
C27136 VDD.n7929 VSS 0.015517f
C27137 VDD.n7930 VSS 0.010511f
C27138 VDD.n7931 VSS 0.024532f
C27139 VDD.n7932 VSS 0.024525f
C27140 VDD.t243 VSS 0.008011f
C27141 VDD.t91 VSS 0.008011f
C27142 VDD.n7933 VSS 0.018207f
C27143 VDD.n7934 VSS 0.015517f
C27144 VDD.n7935 VSS 0.010511f
C27145 VDD.n7936 VSS 0.019382f
C27146 VDD.n7937 VSS 0.019375f
C27147 VDD.t163 VSS 0.008011f
C27148 VDD.t238 VSS 0.008011f
C27149 VDD.n7938 VSS 0.018207f
C27150 VDD.n7939 VSS 0.015517f
C27151 VDD.n7940 VSS 0.010511f
C27152 VDD.n7941 VSS 0.03438f
C27153 VDD.n7942 VSS 0.150048f
C27154 VDD.n7943 VSS 0.145508f
C27155 VDD.t3986 VSS 0.066856f
C27156 VDD.n7944 VSS 0.163358f
C27157 VDD.t1397 VSS 0.066856f
C27158 VDD.n7945 VSS 0.163358f
C27159 VDD.n7946 VSS 0.154425f
C27160 VDD.n7947 VSS 0.208309f
C27161 VDD.t46 VSS 0.008011f
C27162 VDD.t38 VSS 0.008011f
C27163 VDD.n7948 VSS 0.029324f
C27164 VDD.n7949 VSS 0.072806f
C27165 VDD.t36 VSS 0.008011f
C27166 VDD.t29 VSS 0.008011f
C27167 VDD.n7950 VSS 0.029324f
C27168 VDD.n7951 VSS 0.053965f
C27169 VDD.t109 VSS 0.029515f
C27170 VDD.n7952 VSS 0.062674f
C27171 VDD.t210 VSS 0.008011f
C27172 VDD.t281 VSS 0.008011f
C27173 VDD.n7953 VSS 0.029389f
C27174 VDD.n7954 VSS 0.06486f
C27175 VDD.t22 VSS 0.008011f
C27176 VDD.t44 VSS 0.008011f
C27177 VDD.n7955 VSS 0.029324f
C27178 VDD.n7956 VSS 0.064798f
C27179 VDD.t16 VSS 0.008011f
C27180 VDD.t42 VSS 0.008011f
C27181 VDD.n7957 VSS 0.029324f
C27182 VDD.n7958 VSS 0.072559f
C27183 VDD.n7959 VSS 0.209012f
C27184 VDD.n7960 VSS 0.347026f
C27185 VDD.t4132 VSS 0.066856f
C27186 VDD.n7961 VSS 0.27209f
C27187 VDD.t2757 VSS 0.066856f
C27188 VDD.n7962 VSS 0.27209f
C27189 VDD.n7963 VSS 0.091748f
C27190 VDD.n7964 VSS 0.016021f
C27191 VDD.t4133 VSS 0.025104f
C27192 VDD.n7965 VSS 0.293433f
C27193 VDD.n7966 VSS 0.293433f
C27194 VDD.t1883 VSS 0.066856f
C27195 VDD.n7967 VSS 0.27209f
C27196 VDD.n7968 VSS 0.25586f
C27197 VDD.t3351 VSS 0.034186f
C27198 VDD.n7969 VSS 0.25586f
C27199 VDD.n7970 VSS 0.248157f
C27200 VDD.n7971 VSS 0.016021f
C27201 VDD.t1014 VSS 0.016021f
C27202 VDD.n7972 VSS 0.016021f
C27203 VDD.n7973 VSS 0.230682f
C27204 VDD.t2441 VSS 0.066856f
C27205 VDD.n7974 VSS 0.27209f
C27206 VDD.n7975 VSS 0.25586f
C27207 VDD.t3688 VSS 0.034186f
C27208 VDD.n7976 VSS 0.25586f
C27209 VDD.n7977 VSS 0.248157f
C27210 VDD.n7978 VSS 0.016021f
C27211 VDD.t1432 VSS 0.025104f
C27212 VDD.n7979 VSS 0.255859f
C27213 VDD.n7980 VSS 0.255859f
C27214 VDD.t3647 VSS 0.025104f
C27215 VDD.n7981 VSS 0.016021f
C27216 VDD.n7982 VSS 0.248157f
C27217 VDD.n7983 VSS 0.255859f
C27218 VDD.t3402 VSS 0.025104f
C27219 VDD.n7984 VSS 0.016021f
C27220 VDD.t2009 VSS 0.016021f
C27221 VDD.n7985 VSS 0.016021f
C27222 VDD.t1109 VSS 0.025104f
C27223 VDD.n7986 VSS 0.247995f
C27224 VDD.t3792 VSS 0.066856f
C27225 VDD.n7987 VSS 0.272089f
C27226 VDD.t1108 VSS 0.066856f
C27227 VDD.n7988 VSS 0.272089f
C27228 VDD.n7989 VSS 0.248157f
C27229 VDD.n7990 VSS 0.016021f
C27230 VDD.t1021 VSS 0.016021f
C27231 VDD.n7991 VSS 0.016021f
C27232 VDD.n7992 VSS 0.034078f
C27233 VDD.n7993 VSS 0.243788f
C27234 VDD.n7994 VSS 0.311265f
C27235 VDD.n7995 VSS 1.4234f
C27236 VDD.n7996 VSS 0.312066f
C27237 VDD.n7997 VSS 0.051391f
C27238 VDD.n7998 VSS 0.095726f
C27239 VDD.n7999 VSS 0.016021f
C27240 VDD.t1587 VSS 0.025104f
C27241 VDD.n8000 VSS 0.107953f
C27242 VDD.n8001 VSS 0.107953f
C27243 VDD.t3834 VSS 0.066856f
C27244 VDD.n8002 VSS 0.126716f
C27245 VDD.n8003 VSS 0.102784f
C27246 VDD.n8004 VSS 0.016021f
C27247 VDD.t4729 VSS 0.016021f
C27248 VDD.n8005 VSS 0.016021f
C27249 VDD.n8006 VSS 0.102784f
C27250 VDD.t3377 VSS 0.066856f
C27251 VDD.n8007 VSS 0.126716f
C27252 VDD.n8008 VSS 0.102784f
C27253 VDD.n8009 VSS 0.016021f
C27254 VDD.t4277 VSS 0.025104f
C27255 VDD.n8010 VSS 0.111391f
C27256 VDD.n8011 VSS 0.085484f
C27257 VDD.n8012 VSS 0.090906f
C27258 VDD.t4686 VSS 0.043485f
C27259 VDD.n8013 VSS 0.14041f
C27260 VDD.t912 VSS 0.066856f
C27261 VDD.n8014 VSS 0.197337f
C27262 VDD.n8015 VSS 0.207237f
C27263 VDD.t2429 VSS 0.043485f
C27264 VDD.n8016 VSS 0.17899f
C27265 VDD.n8017 VSS 0.129987f
C27266 VDD.n8018 VSS 0.034227f
C27267 VDD.t25 VSS 0.008011f
C27268 VDD.t47 VSS 0.008011f
C27269 VDD.n8019 VSS 0.018285f
C27270 VDD.n8020 VSS 0.015766f
C27271 VDD.n8021 VSS 0.010511f
C27272 VDD.n8022 VSS 0.019381f
C27273 VDD.n8023 VSS 0.019376f
C27274 VDD.t32 VSS 0.008011f
C27275 VDD.t20 VSS 0.008011f
C27276 VDD.n8024 VSS 0.018285f
C27277 VDD.n8025 VSS 0.015766f
C27278 VDD.n8026 VSS 0.010511f
C27279 VDD.n8027 VSS 0.013697f
C27280 VDD.n8028 VSS 0.013692f
C27281 VDD.t169 VSS 0.019337f
C27282 VDD.n8029 VSS 0.023488f
C27283 VDD.n8030 VSS 0.010511f
C27284 VDD.n8031 VSS 0.019381f
C27285 VDD.n8032 VSS 0.019376f
C27286 VDD.t244 VSS 0.008011f
C27287 VDD.t48 VSS 0.008011f
C27288 VDD.n8033 VSS 0.018285f
C27289 VDD.n8034 VSS 0.015766f
C27290 VDD.n8035 VSS 0.010511f
C27291 VDD.n8036 VSS 0.024531f
C27292 VDD.n8037 VSS 0.024526f
C27293 VDD.t40 VSS 0.008011f
C27294 VDD.t33 VSS 0.008011f
C27295 VDD.n8038 VSS 0.018285f
C27296 VDD.n8039 VSS 0.015766f
C27297 VDD.n8040 VSS 0.010511f
C27298 VDD.n8041 VSS 0.019381f
C27299 VDD.n8042 VSS 0.019376f
C27300 VDD.t24 VSS 0.008011f
C27301 VDD.t43 VSS 0.008011f
C27302 VDD.n8043 VSS 0.018285f
C27303 VDD.n8044 VSS 0.015766f
C27304 VDD.n8045 VSS 0.010511f
C27305 VDD.n8046 VSS 0.034424f
C27306 VDD.n8047 VSS 0.214117f
C27307 VDD.n8048 VSS 0.148143f
C27308 VDD.t2199 VSS 0.066856f
C27309 VDD.n8049 VSS 0.163358f
C27310 VDD.t3780 VSS 0.066856f
C27311 VDD.n8050 VSS 0.163358f
C27312 VDD.n8051 VSS 0.148953f
C27313 VDD.n8052 VSS 0.155735f
C27314 VDD.t174 VSS 0.008011f
C27315 VDD.t249 VSS 0.008011f
C27316 VDD.n8053 VSS 0.028899f
C27317 VDD.n8054 VSS 0.072165f
C27318 VDD.t260 VSS 0.008011f
C27319 VDD.t102 VSS 0.008011f
C27320 VDD.n8055 VSS 0.028899f
C27321 VDD.n8056 VSS 0.053429f
C27322 VDD.t209 VSS 0.029106f
C27323 VDD.n8057 VSS 0.061996f
C27324 VDD.t78 VSS 0.008011f
C27325 VDD.t159 VSS 0.008011f
C27326 VDD.n8058 VSS 0.028899f
C27327 VDD.n8059 VSS 0.064263f
C27328 VDD.t143 VSS 0.008011f
C27329 VDD.t189 VSS 0.008011f
C27330 VDD.n8060 VSS 0.028899f
C27331 VDD.n8061 VSS 0.064263f
C27332 VDD.t166 VSS 0.008011f
C27333 VDD.t217 VSS 0.008011f
C27334 VDD.n8062 VSS 0.028899f
C27335 VDD.n8063 VSS 0.071961f
C27336 VDD.n8064 VSS 0.180708f
C27337 VDD.t1099 VSS 0.066856f
C27338 VDD.n8065 VSS 0.172861f
C27339 VDD.t571 VSS 0.043485f
C27340 VDD.n8066 VSS 0.111785f
C27341 VDD.n8067 VSS 0.117631f
C27342 VDD.n8068 VSS 0.069759f
C27343 VDD.n8069 VSS 0.086443f
C27344 VDD.t1361 VSS 0.043485f
C27345 VDD.n8070 VSS 0.097632f
C27346 VDD.n8071 VSS 0.080846f
C27347 VDD.n8072 VSS 0.009613f
C27348 VDD.t2843 VSS 0.009613f
C27349 VDD.n8073 VSS 0.009613f
C27350 VDD.n8074 VSS 0.056791f
C27351 VDD.n8075 VSS 0.040422f
C27352 VDD.n8076 VSS 0.154413f
C27353 VDD.n8077 VSS 1.4234f
C27354 VDD.n8078 VSS 0.154999f
C27355 VDD.n8079 VSS 0.040084f
C27356 VDD.t2771 VSS 0.043485f
C27357 VDD.n8080 VSS 0.088711f
C27358 VDD.n8081 VSS 0.056316f
C27359 VDD.n8082 VSS 0.009613f
C27360 VDD.t2772 VSS 0.009613f
C27361 VDD.n8083 VSS 0.009613f
C27362 VDD.t1279 VSS 0.014798f
C27363 VDD.n8084 VSS 0.099647f
C27364 VDD.t1278 VSS 0.043485f
C27365 VDD.n8085 VSS 0.078673f
C27366 VDD.n8086 VSS 0.031734f
C27367 VDD.n8087 VSS 0.848485f
C27368 VDD.n8088 VSS 0.495896f
C27369 VDD.n8089 VSS 1.8928f
C27370 VDD.n8090 VSS 0.009312f
C27371 VDD.n8091 VSS 0.009688f
C27372 VDD.n8092 VSS 0.202652f
C27373 VDD.n8094 VSS 0.01502f
C27374 VDD.n8095 VSS 0.079539f
C27375 VDD.t653 VSS 0.028519f
C27376 VDD.t3465 VSS 0.028519f
C27377 VDD.n8096 VSS 0.009191f
C27378 VDD.n8097 VSS 0.06055f
C27379 VDD.n8098 VSS 0.15537f
C27380 VDD.n8099 VSS 0.099723f
C27381 VDD.t2084 VSS 0.066856f
C27382 VDD.n8100 VSS 0.125227f
C27383 VDD.n8101 VSS 0.101294f
C27384 VDD.n8102 VSS 0.016021f
C27385 VDD.t675 VSS 0.025104f
C27386 VDD.n8103 VSS 0.081176f
C27387 VDD.n8104 VSS 0.048151f
C27388 VDD.n8105 VSS 0.083673f
C27389 VDD.t864 VSS 0.066856f
C27390 VDD.n8106 VSS 0.125227f
C27391 VDD.n8107 VSS 0.101294f
C27392 VDD.n8108 VSS 0.016021f
C27393 VDD.t4107 VSS 0.025104f
C27394 VDD.n8109 VSS 0.099723f
C27395 VDD.n8110 VSS 0.62132f
C27396 VDD.n8111 VSS 0.099723f
C27397 VDD.t1496 VSS 0.066856f
C27398 VDD.n8112 VSS 0.125227f
C27399 VDD.n8113 VSS 0.101294f
C27400 VDD.n8114 VSS 0.016021f
C27401 VDD.t4299 VSS 0.025104f
C27402 VDD.n8115 VSS 0.081176f
C27403 VDD.n8116 VSS 0.048151f
C27404 VDD.n8117 VSS 0.083673f
C27405 VDD.t4450 VSS 0.066856f
C27406 VDD.n8118 VSS 0.125227f
C27407 VDD.n8119 VSS 0.101294f
C27408 VDD.n8120 VSS 0.016021f
C27409 VDD.t3551 VSS 0.025104f
C27410 VDD.n8121 VSS 0.099723f
C27411 VDD.t1016 VSS 0.028519f
C27412 VDD.t4259 VSS 0.028519f
C27413 VDD.n8122 VSS 0.009191f
C27414 VDD.t1015 VSS 0.066856f
C27415 VDD.t2753 VSS 0.066856f
C27416 VDD.t637 VSS 0.028519f
C27417 VDD.t3903 VSS 0.028519f
C27418 VDD.n8123 VSS 0.009191f
C27419 VDD.t636 VSS 0.066856f
C27420 VDD.t2382 VSS 0.066856f
C27421 VDD.t3250 VSS 0.066856f
C27422 VDD.t679 VSS 0.066856f
C27423 VDD.t3488 VSS 0.066856f
C27424 VDD.t2351 VSS 0.066856f
C27425 VDD.n8124 VSS 0.690489f
C27426 VDD.t955 VSS 0.066856f
C27427 VDD.t3902 VSS 0.066856f
C27428 VDD.n8125 VSS 0.690489f
C27429 VDD.t2383 VSS 0.028519f
C27430 VDD.t956 VSS 0.028519f
C27431 VDD.n8126 VSS 0.009191f
C27432 VDD.n8127 VSS 0.644755f
C27433 VDD.t1262 VSS 0.066856f
C27434 VDD.t4258 VSS 0.066856f
C27435 VDD.n8128 VSS 0.709674f
C27436 VDD.t2754 VSS 0.028519f
C27437 VDD.t1263 VSS 0.028519f
C27438 VDD.n8129 VSS 0.009191f
C27439 VDD.n8130 VSS 0.261039f
C27440 VDD.n8131 VSS 0.62132f
C27441 VDD.n8132 VSS 0.099723f
C27442 VDD.t3367 VSS 0.066856f
C27443 VDD.n8133 VSS 0.125227f
C27444 VDD.n8134 VSS 0.101294f
C27445 VDD.n8135 VSS 0.016021f
C27446 VDD.t1982 VSS 0.025104f
C27447 VDD.n8136 VSS 0.081176f
C27448 VDD.n8137 VSS 0.048151f
C27449 VDD.n8138 VSS 0.083673f
C27450 VDD.t2150 VSS 0.066856f
C27451 VDD.n8139 VSS 0.125227f
C27452 VDD.n8140 VSS 0.006598f
C27453 VDD.t1206 VSS 0.066856f
C27454 VDD.n8141 VSS 0.045867f
C27455 VDD.n8142 VSS 0.015693f
C27456 VDD.n8143 VSS 0.010188f
C27457 VDD.t339 VSS 0.020392f
C27458 VDD.t305 VSS 0.022133f
C27459 VDD.n8144 VSS 0.069721f
C27460 VDD.n8145 VSS 0.040089f
C27461 VDD.t365 VSS 0.020371f
C27462 VDD.n8146 VSS 0.027146f
C27463 VDD.t303 VSS 0.022106f
C27464 VDD.n8147 VSS 0.036568f
C27465 VDD.n8148 VSS 0.044801f
C27466 VDD.n8149 VSS 0.278297f
C27467 VDD.n8150 VSS 0.040089f
C27468 VDD.t14 VSS 0.020371f
C27469 VDD.n8151 VSS 0.027146f
C27470 VDD.t366 VSS 0.020392f
C27471 VDD.n8152 VSS 0.049654f
C27472 VDD.t4767 VSS 0.017093f
C27473 VDD.n8153 VSS 0.042096f
C27474 VDD.n8154 VSS 0.069466f
C27475 VDD.t4766 VSS 0.017093f
C27476 VDD.n8155 VSS 0.035464f
C27477 VDD.n8156 VSS 0.016538f
C27478 VDD.n8157 VSS 0.027213f
C27479 VDD.n8158 VSS 0.204333f
C27480 VDD.n8159 VSS 0.030906f
C27481 VDD.n8160 VSS 0.010881f
C27482 VDD.n8161 VSS 0.044227f
C27483 VDD.n8162 VSS 0.094696f
C27484 VDD.n8163 VSS 0.016021f
C27485 VDD.t1207 VSS 0.025104f
C27486 VDD.n8164 VSS 0.08403f
C27487 VDD.n8165 VSS 0.075174f
C27488 VDD.t2125 VSS 0.028519f
C27489 VDD.t759 VSS 0.028519f
C27490 VDD.n8166 VSS 0.009191f
C27491 VDD.n8167 VSS 0.05425f
C27492 VDD.n8168 VSS 0.073151f
C27493 VDD.n8169 VSS 0.012131f
C27494 VDD.n8170 VSS 0.012131f
C27495 VDD.n8171 VSS 0.012131f
C27496 VDD.n8172 VSS 0.077187f
C27497 VDD.t2124 VSS 0.066856f
C27498 VDD.t757 VSS 0.066856f
C27499 VDD.n8173 VSS 0.10134f
C27500 VDD.n8174 VSS 0.083241f
C27501 VDD.n8175 VSS 0.106951f
C27502 VDD.n8176 VSS 0.012131f
C27503 VDD.n8177 VSS 0.012131f
C27504 VDD.n8178 VSS 0.012131f
C27505 VDD.n8179 VSS 0.106951f
C27506 VDD.n8180 VSS 0.106951f
C27507 VDD.t1735 VSS 0.028519f
C27508 VDD.t4519 VSS 0.028519f
C27509 VDD.n8181 VSS 0.009191f
C27510 VDD.n8182 VSS 0.06888f
C27511 VDD.n8183 VSS 0.058016f
C27512 VDD.n8184 VSS 0.012131f
C27513 VDD.n8185 VSS 0.012131f
C27514 VDD.n8186 VSS 0.012131f
C27515 VDD.n8187 VSS 0.101402f
C27516 VDD.t1734 VSS 0.066856f
C27517 VDD.t4518 VSS 0.066856f
C27518 VDD.n8188 VSS 0.10134f
C27519 VDD.n8189 VSS 0.059025f
C27520 VDD.n8190 VSS 0.106951f
C27521 VDD.n8191 VSS 0.012131f
C27522 VDD.n8192 VSS 0.012131f
C27523 VDD.n8193 VSS 0.012131f
C27524 VDD.n8194 VSS 0.106951f
C27525 VDD.n8195 VSS 0.106951f
C27526 VDD.n8196 VSS 0.068106f
C27527 VDD.n8197 VSS 0.012131f
C27528 VDD.n8198 VSS 0.012131f
C27529 VDD.n8199 VSS 0.092321f
C27530 VDD.n8200 VSS 0.106951f
C27531 VDD.t4305 VSS 0.028519f
C27532 VDD.t3021 VSS 0.028519f
C27533 VDD.n8201 VSS 0.009191f
C27534 VDD.n8202 VSS 0.06888f
C27535 VDD.n8203 VSS 0.058016f
C27536 VDD.n8204 VSS 0.012131f
C27537 VDD.n8205 VSS 0.012131f
C27538 VDD.n8206 VSS 0.012131f
C27539 VDD.n8207 VSS 0.106951f
C27540 VDD.n8208 VSS 0.106951f
C27541 VDD.n8209 VSS 0.056503f
C27542 VDD.n8210 VSS 0.012131f
C27543 VDD.n8211 VSS 0.012131f
C27544 VDD.n8212 VSS 0.103924f
C27545 VDD.n8213 VSS 0.106951f
C27546 VDD.t1721 VSS 0.028519f
C27547 VDD.t4505 VSS 0.028519f
C27548 VDD.n8214 VSS 0.009191f
C27549 VDD.n8215 VSS 0.06888f
C27550 VDD.n8216 VSS 0.070124f
C27551 VDD.n8217 VSS 0.012131f
C27552 VDD.n8218 VSS 0.012131f
C27553 VDD.n8219 VSS 0.012131f
C27554 VDD.n8220 VSS 0.106951f
C27555 VDD.n8221 VSS 0.060034f
C27556 VDD.t1720 VSS 0.066856f
C27557 VDD.t4504 VSS 0.066856f
C27558 VDD.n8222 VSS 0.10134f
C27559 VDD.n8223 VSS 0.100393f
C27560 VDD.n8224 VSS 0.012131f
C27561 VDD.n8225 VSS 0.012131f
C27562 VDD.n8226 VSS 0.012131f
C27563 VDD.n8227 VSS 0.106951f
C27564 VDD.n8228 VSS 0.106951f
C27565 VDD.t1351 VSS 0.066856f
C27566 VDD.t4174 VSS 0.066856f
C27567 VDD.n8229 VSS 0.10134f
C27568 VDD.n8230 VSS 0.080214f
C27569 VDD.n8231 VSS 0.012131f
C27570 VDD.n8232 VSS 0.012131f
C27571 VDD.n8233 VSS 0.012131f
C27572 VDD.n8234 VSS 0.106951f
C27573 VDD.n8235 VSS 0.070124f
C27574 VDD.t1353 VSS 0.028519f
C27575 VDD.t4175 VSS 0.028519f
C27576 VDD.n8236 VSS 0.009191f
C27577 VDD.n8237 VSS 0.06888f
C27578 VDD.n8238 VSS 0.090303f
C27579 VDD.n8239 VSS 0.012131f
C27580 VDD.n8240 VSS 0.012131f
C27581 VDD.n8241 VSS 0.012131f
C27582 VDD.n8242 VSS 0.106951f
C27583 VDD.n8243 VSS 0.106951f
C27584 VDD.n8244 VSS 0.104429f
C27585 VDD.n8245 VSS 0.012131f
C27586 VDD.n8246 VSS 0.012131f
C27587 VDD.n8247 VSS 0.055998f
C27588 VDD.n8248 VSS 0.106951f
C27589 VDD.t3037 VSS 0.028519f
C27590 VDD.t4185 VSS 0.028519f
C27591 VDD.n8249 VSS 0.009191f
C27592 VDD.n8250 VSS 0.06888f
C27593 VDD.n8251 VSS 0.094339f
C27594 VDD.n8252 VSS 0.012131f
C27595 VDD.n8253 VSS 0.012131f
C27596 VDD.n8254 VSS 0.012131f
C27597 VDD.n8255 VSS 0.012131f
C27598 VDD.n8256 VSS 0.012131f
C27599 VDD.n8257 VSS 0.012131f
C27600 VDD.n8258 VSS 0.012131f
C27601 VDD.n8259 VSS 0.012131f
C27602 VDD.n8260 VSS 0.012131f
C27603 VDD.n8261 VSS 0.012131f
C27604 VDD.n8262 VSS 0.012131f
C27605 VDD.n8263 VSS 0.012131f
C27606 VDD.n8264 VSS 0.012131f
C27607 VDD.n8265 VSS 0.012131f
C27608 VDD.n8266 VSS 0.012131f
C27609 VDD.n8267 VSS 0.012131f
C27610 VDD.n8268 VSS 0.012131f
C27611 VDD.n8269 VSS 0.012131f
C27612 VDD.n8270 VSS 0.012131f
C27613 VDD.n8271 VSS 0.012131f
C27614 VDD.n8272 VSS 0.012131f
C27615 VDD.n8273 VSS 0.012131f
C27616 VDD.n8274 VSS 0.012131f
C27617 VDD.n8275 VSS 0.012131f
C27618 VDD.n8276 VSS 0.012131f
C27619 VDD.n8277 VSS 0.012131f
C27620 VDD.n8278 VSS 0.012131f
C27621 VDD.n8279 VSS 0.012131f
C27622 VDD.n8280 VSS 0.012131f
C27623 VDD.n8281 VSS 0.012131f
C27624 VDD.n8282 VSS 0.012131f
C27625 VDD.n8283 VSS 0.012131f
C27626 VDD.n8284 VSS 0.012131f
C27627 VDD.n8285 VSS 0.012131f
C27628 VDD.n8286 VSS 0.012131f
C27629 VDD.n8287 VSS 0.012131f
C27630 VDD.n8288 VSS 0.012131f
C27631 VDD.n8289 VSS 0.012131f
C27632 VDD.n8290 VSS 0.012131f
C27633 VDD.n8291 VSS 0.012131f
C27634 VDD.n8292 VSS 0.012131f
C27635 VDD.n8293 VSS 0.012131f
C27636 VDD.n8294 VSS 0.012131f
C27637 VDD.n8295 VSS 0.012131f
C27638 VDD.n8296 VSS 0.012131f
C27639 VDD.n8297 VSS 0.012131f
C27640 VDD.n8298 VSS 0.012131f
C27641 VDD.n8299 VSS 0.012131f
C27642 VDD.n8300 VSS 0.012131f
C27643 VDD.n8301 VSS 0.012131f
C27644 VDD.n8302 VSS 0.012131f
C27645 VDD.n8303 VSS 0.012131f
C27646 VDD.n8304 VSS 0.012131f
C27647 VDD.n8305 VSS 0.012131f
C27648 VDD.n8306 VSS 0.012131f
C27649 VDD.n8307 VSS 0.012131f
C27650 VDD.n8308 VSS 0.012131f
C27651 VDD.n8309 VSS 0.012131f
C27652 VDD.n8310 VSS 0.012131f
C27653 VDD.n8311 VSS 0.012131f
C27654 VDD.n8312 VSS 0.012131f
C27655 VDD.n8313 VSS 0.012131f
C27656 VDD.n8314 VSS 0.012131f
C27657 VDD.n8315 VSS 0.012131f
C27658 VDD.n8316 VSS 0.012131f
C27659 VDD.n8317 VSS 0.012131f
C27660 VDD.n8318 VSS 0.012131f
C27661 VDD.n8319 VSS 0.012131f
C27662 VDD.n8320 VSS 0.012131f
C27663 VDD.n8321 VSS 0.012131f
C27664 VDD.n8322 VSS 0.012131f
C27665 VDD.n8323 VSS 0.012131f
C27666 VDD.n8324 VSS 0.012131f
C27667 VDD.n8325 VSS 0.012131f
C27668 VDD.n8326 VSS 0.012131f
C27669 VDD.n8327 VSS 0.012131f
C27670 VDD.n8328 VSS 0.012131f
C27671 VDD.n8329 VSS 0.012131f
C27672 VDD.n8330 VSS 0.012131f
C27673 VDD.n8331 VSS 0.012131f
C27674 VDD.n8332 VSS 0.012131f
C27675 VDD.n8333 VSS 0.012131f
C27676 VDD.n8334 VSS 0.012131f
C27677 VDD.n8335 VSS 0.012131f
C27678 VDD.n8336 VSS 0.012131f
C27679 VDD.n8337 VSS 0.012131f
C27680 VDD.n8338 VSS 0.012131f
C27681 VDD.n8339 VSS 0.012131f
C27682 VDD.n8340 VSS 0.012131f
C27683 VDD.n8341 VSS 0.012131f
C27684 VDD.n8342 VSS 0.012131f
C27685 VDD.n8343 VSS 0.012131f
C27686 VDD.n8344 VSS 0.012131f
C27687 VDD.n8345 VSS 0.012131f
C27688 VDD.n8346 VSS 0.012131f
C27689 VDD.n8347 VSS 0.012131f
C27690 VDD.n8348 VSS 0.012131f
C27691 VDD.n8349 VSS 0.012131f
C27692 VDD.n8350 VSS 0.012131f
C27693 VDD.n8351 VSS 0.012131f
C27694 VDD.n8352 VSS 0.012131f
C27695 VDD.n8353 VSS 0.012131f
C27696 VDD.n8354 VSS 0.012131f
C27697 VDD.n8355 VSS 0.012131f
C27698 VDD.n8356 VSS 0.012131f
C27699 VDD.n8357 VSS 0.012131f
C27700 VDD.n8358 VSS 0.012131f
C27701 VDD.n8359 VSS 0.012131f
C27702 VDD.n8360 VSS 0.012131f
C27703 VDD.n8361 VSS 0.012131f
C27704 VDD.n8362 VSS 0.012131f
C27705 VDD.n8363 VSS 0.012131f
C27706 VDD.n8364 VSS 0.012131f
C27707 VDD.n8365 VSS 0.012131f
C27708 VDD.n8366 VSS 0.012131f
C27709 VDD.n8367 VSS 0.012131f
C27710 VDD.n8368 VSS 0.012131f
C27711 VDD.n8369 VSS 0.012131f
C27712 VDD.n8370 VSS 0.012131f
C27713 VDD.n8371 VSS 0.012131f
C27714 VDD.n8372 VSS 0.012131f
C27715 VDD.n8373 VSS 0.012131f
C27716 VDD.n8374 VSS 0.012131f
C27717 VDD.n8375 VSS 0.012131f
C27718 VDD.n8376 VSS 0.012131f
C27719 VDD.n8377 VSS 0.012131f
C27720 VDD.n8378 VSS 0.012131f
C27721 VDD.n8379 VSS 0.012131f
C27722 VDD.n8380 VSS 0.012131f
C27723 VDD.n8381 VSS 0.012131f
C27724 VDD.n8382 VSS 0.012131f
C27725 VDD.n8383 VSS 0.012131f
C27726 VDD.n8384 VSS 0.012131f
C27727 VDD.n8385 VSS 0.012131f
C27728 VDD.n8386 VSS 0.012131f
C27729 VDD.n8387 VSS 0.012131f
C27730 VDD.n8388 VSS 0.012131f
C27731 VDD.n8389 VSS 0.012131f
C27732 VDD.n8390 VSS 0.012131f
C27733 VDD.n8391 VSS 0.012131f
C27734 VDD.n8392 VSS 0.012131f
C27735 VDD.n8393 VSS 0.012131f
C27736 VDD.n8394 VSS 0.012131f
C27737 VDD.n8395 VSS 0.012131f
C27738 VDD.n8396 VSS 0.012131f
C27739 VDD.n8397 VSS 0.012131f
C27740 VDD.n8398 VSS 0.012131f
C27741 VDD.n8399 VSS 0.012131f
C27742 VDD.n8400 VSS 0.012131f
C27743 VDD.n8401 VSS 0.012131f
C27744 VDD.n8402 VSS 0.012131f
C27745 VDD.n8403 VSS 0.012131f
C27746 VDD.n8404 VSS 0.012131f
C27747 VDD.n8405 VSS 0.012131f
C27748 VDD.n8406 VSS 0.012131f
C27749 VDD.n8407 VSS 0.012131f
C27750 VDD.n8408 VSS 0.012131f
C27751 VDD.n8409 VSS 0.012131f
C27752 VDD.n8410 VSS 0.012131f
C27753 VDD.n8411 VSS 0.012131f
C27754 VDD.n8412 VSS 0.012131f
C27755 VDD.n8413 VSS 0.012131f
C27756 VDD.n8414 VSS 0.012131f
C27757 VDD.n8415 VSS 0.012131f
C27758 VDD.n8416 VSS 0.012131f
C27759 VDD.n8417 VSS 0.012131f
C27760 VDD.n8418 VSS 0.012131f
C27761 VDD.n8419 VSS 0.012131f
C27762 VDD.n8420 VSS 0.012131f
C27763 VDD.n8421 VSS 0.012131f
C27764 VDD.n8422 VSS 0.012131f
C27765 VDD.n8423 VSS 0.012131f
C27766 VDD.n8424 VSS 0.012131f
C27767 VDD.n8425 VSS 0.012131f
C27768 VDD.n8426 VSS 0.012131f
C27769 VDD.n8427 VSS 0.012131f
C27770 VDD.n8428 VSS 0.012131f
C27771 VDD.n8429 VSS 0.012131f
C27772 VDD.n8430 VSS 0.012131f
C27773 VDD.n8431 VSS 0.012131f
C27774 VDD.n8432 VSS 0.012131f
C27775 VDD.n8433 VSS 0.012131f
C27776 VDD.n8434 VSS 0.012131f
C27777 VDD.n8435 VSS 0.012131f
C27778 VDD.n8436 VSS 0.012131f
C27779 VDD.n8437 VSS 0.012131f
C27780 VDD.n8438 VSS 0.012131f
C27781 VDD.n8439 VSS 0.012131f
C27782 VDD.n8440 VSS 0.012131f
C27783 VDD.n8441 VSS 0.012131f
C27784 VDD.n8442 VSS 0.012131f
C27785 VDD.n8443 VSS 0.012131f
C27786 VDD.n8444 VSS 0.012131f
C27787 VDD.n8445 VSS 0.012131f
C27788 VDD.n8446 VSS 0.012131f
C27789 VDD.n8447 VSS 0.012131f
C27790 VDD.n8448 VSS 0.012131f
C27791 VDD.n8449 VSS 0.012131f
C27792 VDD.n8450 VSS 0.012131f
C27793 VDD.n8451 VSS 0.012131f
C27794 VDD.n8452 VSS 0.012131f
C27795 VDD.n8453 VSS 0.012131f
C27796 VDD.n8454 VSS 0.012131f
C27797 VDD.n8455 VSS 0.012131f
C27798 VDD.n8456 VSS 0.012131f
C27799 VDD.n8457 VSS 0.012131f
C27800 VDD.n8458 VSS 0.012131f
C27801 VDD.n8459 VSS 0.179614f
C27802 VDD.n8460 VSS 0.208771f
C27803 VDD.n8461 VSS 0.206947f
C27804 VDD.n8462 VSS 0.865258f
C27805 VDD.t4657 VSS 0.028519f
C27806 VDD.t3167 VSS 0.028519f
C27807 VDD.n8463 VSS 0.009191f
C27808 VDD.t3261 VSS 0.028519f
C27809 VDD.t3441 VSS 0.028519f
C27810 VDD.n8464 VSS 0.009191f
C27811 VDD.n8465 VSS 0.471397f
C27812 VDD.n8466 VSS 0.207221f
C27813 VDD.t4077 VSS 0.028519f
C27814 VDD.t2602 VSS 0.028519f
C27815 VDD.n8467 VSS 0.009191f
C27816 VDD.t4076 VSS 0.066856f
C27817 VDD.t2686 VSS 0.066856f
C27818 VDD.t4434 VSS 0.066856f
C27819 VDD.t3054 VSS 0.066856f
C27820 VDD.t4435 VSS 0.028519f
C27821 VDD.t2971 VSS 0.028519f
C27822 VDD.n8468 VSS 0.009191f
C27823 VDD.t1868 VSS 0.066856f
C27824 VDD.t4540 VSS 0.066856f
C27825 VDD.t1870 VSS 0.028519f
C27826 VDD.t4465 VSS 0.028519f
C27827 VDD.n8469 VSS 0.009191f
C27828 VDD.n8470 VSS 0.099723f
C27829 VDD.t3102 VSS 0.066856f
C27830 VDD.n8471 VSS 0.125227f
C27831 VDD.t4569 VSS 0.025104f
C27832 VDD.n8472 VSS 0.081176f
C27833 VDD.n8473 VSS 0.208534f
C27834 VDD.t2131 VSS 1.36988f
C27835 VDD.t607 VSS 1.45794f
C27836 VDD.t2257 VSS 1.96535f
C27837 VDD.t683 VSS 1.96535f
C27838 VDD.t2305 VSS 1.31955f
C27839 VDD.t2130 VSS 0.066856f
C27840 VDD.n8474 VSS 0.14405f
C27841 VDD.t1896 VSS 0.025104f
C27842 VDD.n8475 VSS 0.033925f
C27843 VDD.n8476 VSS 0.116823f
C27844 VDD.t1920 VSS 0.028519f
C27845 VDD.t2160 VSS 0.028519f
C27846 VDD.n8477 VSS 0.009191f
C27847 VDD.t1918 VSS 0.066856f
C27848 VDD.t2163 VSS 0.066856f
C27849 VDD.t2355 VSS 0.028519f
C27850 VDD.t2588 VSS 0.028519f
C27851 VDD.n8478 VSS 0.009191f
C27852 VDD.t2354 VSS 0.066856f
C27853 VDD.t2589 VSS 0.066856f
C27854 VDD.t2990 VSS 0.066856f
C27855 VDD.t3178 VSS 0.066856f
C27856 VDD.t2991 VSS 0.028519f
C27857 VDD.t3177 VSS 0.028519f
C27858 VDD.n8479 VSS 0.009191f
C27859 VDD.n8480 VSS 0.207221f
C27860 VDD.t2375 VSS 0.028519f
C27861 VDD.t2610 VSS 0.028519f
C27862 VDD.n8481 VSS 0.009191f
C27863 VDD.t2374 VSS 0.066856f
C27864 VDD.t2611 VSS 0.066856f
C27865 VDD.t2769 VSS 0.066856f
C27866 VDD.t2986 VSS 0.066856f
C27867 VDD.t2770 VSS 0.028519f
C27868 VDD.t2983 VSS 0.028519f
C27869 VDD.n8482 VSS 0.009191f
C27870 VDD.t4270 VSS 0.066856f
C27871 VDD.t4472 VSS 0.066856f
C27872 VDD.t4271 VSS 0.028519f
C27873 VDD.t4469 VSS 0.028519f
C27874 VDD.n8483 VSS 0.009191f
C27875 VDD.t4256 VSS 0.066856f
C27876 VDD.n8484 VSS 0.125227f
C27877 VDD.t4461 VSS 0.025104f
C27878 VDD.t4460 VSS 0.066856f
C27879 VDD.n8485 VSS 0.125227f
C27880 VDD.n8486 VSS 0.101294f
C27881 VDD.n8487 VSS 0.016021f
C27882 VDD.t4257 VSS 0.025104f
C27883 VDD.n8488 VSS 0.099723f
C27884 VDD.t3024 VSS 0.066856f
C27885 VDD.n8489 VSS 0.125227f
C27886 VDD.t4487 VSS 0.025104f
C27887 VDD.n8490 VSS 0.081176f
C27888 VDD.n8491 VSS 0.208534f
C27889 VDD.t2064 VSS 1.36988f
C27890 VDD.t1895 VSS 1.96535f
C27891 VDD.t2159 VSS 1.96535f
C27892 VDD.t1919 VSS 1.45794f
C27893 VDD.n8492 VSS 0.865258f
C27894 VDD.n8493 VSS 0.865258f
C27895 VDD.t2450 VSS 1.45794f
C27896 VDD.t2164 VSS 1.96535f
C27897 VDD.t564 VSS 1.96535f
C27898 VDD.t2193 VSS 1.31955f
C27899 VDD.t2063 VSS 0.066856f
C27900 VDD.n8494 VSS 0.14405f
C27901 VDD.t1799 VSS 0.025104f
C27902 VDD.t1827 VSS 0.028519f
C27903 VDD.t2083 VSS 0.028519f
C27904 VDD.n8495 VSS 0.009191f
C27905 VDD.t2734 VSS 0.028519f
C27906 VDD.t2951 VSS 0.028519f
C27907 VDD.n8496 VSS 0.009191f
C27908 VDD.n8497 VSS 0.310925f
C27909 VDD.t4290 VSS 0.066856f
C27910 VDD.n8498 VSS 0.14405f
C27911 VDD.t4083 VSS 0.025104f
C27912 VDD.n8499 VSS 0.105404f
C27913 VDD.n8500 VSS 0.208534f
C27914 VDD.n8501 VSS 0.207221f
C27915 VDD.t710 VSS 1.36988f
C27916 VDD.t709 VSS 0.066856f
C27917 VDD.n8502 VSS 0.125227f
C27918 VDD.t2329 VSS 0.025104f
C27919 VDD.t3612 VSS 0.028519f
C27920 VDD.t2507 VSS 0.028519f
C27921 VDD.n8503 VSS 0.009191f
C27922 VDD.t2067 VSS 0.028519f
C27923 VDD.t983 VSS 0.028519f
C27924 VDD.n8504 VSS 0.009191f
C27925 VDD.n8505 VSS 0.261039f
C27926 VDD.t2469 VSS 0.066856f
C27927 VDD.n8506 VSS 0.125227f
C27928 VDD.t1678 VSS 0.025104f
C27929 VDD.n8507 VSS 0.081176f
C27930 VDD.n8508 VSS 0.208534f
C27931 VDD.n8509 VSS 0.207221f
C27932 VDD.t296 VSS 1.36988f
C27933 VDD.t2328 VSS 1.96535f
C27934 VDD.t845 VSS 1.96535f
C27935 VDD.t1254 VSS 1.45794f
C27936 VDD.n8510 VSS 0.865258f
C27937 VDD.n8511 VSS 0.865258f
C27938 VDD.t982 VSS 1.45794f
C27939 VDD.t670 VSS 1.96535f
C27940 VDD.t322 VSS 1.96535f
C27941 VDD.t420 VSS 1.31955f
C27942 VDD.t2530 VSS 0.066856f
C27943 VDD.n8512 VSS 0.14405f
C27944 VDD.t4019 VSS 0.025104f
C27945 VDD.n8513 VSS 0.033925f
C27946 VDD.t3651 VSS 0.028519f
C27947 VDD.t2555 VSS 0.028519f
C27948 VDD.n8514 VSS 0.009191f
C27949 VDD.t2104 VSS 0.028519f
C27950 VDD.t1019 VSS 0.028519f
C27951 VDD.n8515 VSS 0.009191f
C27952 VDD.n8516 VSS 0.308318f
C27953 VDD.t2522 VSS 0.066856f
C27954 VDD.n8517 VSS 0.14405f
C27955 VDD.t3447 VSS 0.025104f
C27956 VDD.n8518 VSS 0.105404f
C27957 VDD.n8519 VSS 0.208534f
C27958 VDD.n8520 VSS 0.207221f
C27959 VDD.t545 VSS 1.36988f
C27960 VDD.t4692 VSS 0.066856f
C27961 VDD.n8521 VSS 0.125227f
C27962 VDD.t1620 VSS 0.025104f
C27963 VDD.t1269 VSS 0.028519f
C27964 VDD.t4709 VSS 0.028519f
C27965 VDD.n8522 VSS 0.009191f
C27966 VDD.t3867 VSS 0.028519f
C27967 VDD.t1337 VSS 0.028519f
C27968 VDD.n8523 VSS 0.009191f
C27969 VDD.n8524 VSS 0.263202f
C27970 VDD.n8525 VSS 0.035132f
C27971 VDD.t2112 VSS 0.025104f
C27972 VDD.n8526 VSS 0.081176f
C27973 VDD.n8527 VSS 0.208534f
C27974 VDD.n8528 VSS 0.207221f
C27975 VDD.t6 VSS 1.36988f
C27976 VDD.t547 VSS 1.96535f
C27977 VDD.t2467 VSS 1.96535f
C27978 VDD.t1268 VSS 1.45794f
C27979 VDD.n8529 VSS 0.902999f
C27980 VDD.n8530 VSS 0.902999f
C27981 VDD.t1336 VSS 1.45794f
C27982 VDD.t1492 VSS 1.96535f
C27983 VDD.t0 VSS 1.96535f
C27984 VDD.t1 VSS 1.31955f
C27985 VDD.t2942 VSS 0.066856f
C27986 VDD.n8531 VSS 0.14405f
C27987 VDD.t3959 VSS 0.025104f
C27988 VDD.t1199 VSS 0.028519f
C27989 VDD.t4283 VSS 0.028519f
C27990 VDD.n8532 VSS 0.009191f
C27991 VDD.t1197 VSS 0.066856f
C27992 VDD.t1410 VSS 0.066856f
C27993 VDD.t1540 VSS 0.028519f
C27994 VDD.t4619 VSS 0.028519f
C27995 VDD.n8533 VSS 0.009191f
C27996 VDD.t1539 VSS 0.066856f
C27997 VDD.t1763 VSS 0.066856f
C27998 VDD.t2211 VSS 0.066856f
C27999 VDD.t2492 VSS 0.066856f
C28000 VDD.t2212 VSS 0.028519f
C28001 VDD.t1098 VSS 0.028519f
C28002 VDD.n8534 VSS 0.009191f
C28003 VDD.t795 VSS 1.96535f
C28004 VDD.t2061 VSS 1.96535f
C28005 VDD.t2814 VSS 1.36988f
C28006 VDD.n8535 VSS 0.645798f
C28007 VDD.n8536 VSS 0.595476f
C28008 VDD.t2023 VSS 1.31955f
C28009 VDD.t2254 VSS 1.96535f
C28010 VDD.t1411 VSS 1.96535f
C28011 VDD.t813 VSS 1.45794f
C28012 VDD.t3 VSS 1.96535f
C28013 VDD.t901 VSS 1.96535f
C28014 VDD.t1198 VSS 1.45794f
C28015 VDD.n8537 VSS 0.865258f
C28016 VDD.n8538 VSS 0.865258f
C28017 VDD.n8539 VSS 0.207221f
C28018 VDD.t1564 VSS 0.028519f
C28019 VDD.t4645 VSS 0.028519f
C28020 VDD.n8540 VSS 0.009191f
C28021 VDD.t1563 VSS 0.066856f
C28022 VDD.t1779 VSS 0.066856f
C28023 VDD.t1965 VSS 0.066856f
C28024 VDD.t2205 VSS 0.066856f
C28025 VDD.t1966 VSS 0.028519f
C28026 VDD.t902 VSS 0.028519f
C28027 VDD.n8541 VSS 0.009191f
C28028 VDD.t3558 VSS 0.066856f
C28029 VDD.t3782 VSS 0.066856f
C28030 VDD.t3559 VSS 0.028519f
C28031 VDD.t2551 VSS 0.028519f
C28032 VDD.n8542 VSS 0.009191f
C28033 VDD.t2133 VSS 0.066856f
C28034 VDD.n8543 VSS 0.125227f
C28035 VDD.t1035 VSS 0.025104f
C28036 VDD.t1034 VSS 0.066856f
C28037 VDD.n8544 VSS 0.125227f
C28038 VDD.n8545 VSS 0.101294f
C28039 VDD.n8546 VSS 0.016021f
C28040 VDD.t2134 VSS 0.025104f
C28041 VDD.n8547 VSS 0.099723f
C28042 VDD.t2253 VSS 0.066856f
C28043 VDD.n8548 VSS 0.125227f
C28044 VDD.t2024 VSS 0.025104f
C28045 VDD.t2813 VSS 0.066856f
C28046 VDD.n8549 VSS 0.125227f
C28047 VDD.t2062 VSS 0.025104f
C28048 VDD.t2060 VSS 0.066856f
C28049 VDD.n8550 VSS 0.125227f
C28050 VDD.n8551 VSS 0.101294f
C28051 VDD.n8552 VSS 0.016021f
C28052 VDD.t2815 VSS 0.025104f
C28053 VDD.n8553 VSS 0.081176f
C28054 VDD.n8554 VSS 0.048151f
C28055 VDD.n8555 VSS 0.083673f
C28056 VDD.t2022 VSS 0.066856f
C28057 VDD.n8556 VSS 0.125227f
C28058 VDD.n8557 VSS 0.101294f
C28059 VDD.n8558 VSS 0.016021f
C28060 VDD.t2255 VSS 0.025104f
C28061 VDD.n8559 VSS 0.099723f
C28062 VDD.n8560 VSS 0.62132f
C28063 VDD.t3783 VSS 0.028519f
C28064 VDD.t814 VSS 0.028519f
C28065 VDD.n8561 VSS 0.009191f
C28066 VDD.n8562 VSS 0.261039f
C28067 VDD.t812 VSS 0.066856f
C28068 VDD.t2550 VSS 0.066856f
C28069 VDD.n8563 VSS 0.709674f
C28070 VDD.t2206 VSS 0.028519f
C28071 VDD.t3384 VSS 0.028519f
C28072 VDD.n8564 VSS 0.009191f
C28073 VDD.n8565 VSS 0.644755f
C28074 VDD.t3383 VSS 0.066856f
C28075 VDD.t900 VSS 0.066856f
C28076 VDD.n8566 VSS 0.690489f
C28077 VDD.t3066 VSS 0.066856f
C28078 VDD.t4644 VSS 0.066856f
C28079 VDD.n8567 VSS 0.690489f
C28080 VDD.t1780 VSS 0.028519f
C28081 VDD.t3067 VSS 0.028519f
C28082 VDD.n8568 VSS 0.009191f
C28083 VDD.n8569 VSS 0.523473f
C28084 VDD.n8570 VSS 0.524869f
C28085 VDD.t2493 VSS 0.028519f
C28086 VDD.t3596 VSS 0.028519f
C28087 VDD.n8571 VSS 0.009191f
C28088 VDD.n8572 VSS 0.471397f
C28089 VDD.t3595 VSS 0.066856f
C28090 VDD.t1097 VSS 0.066856f
C28091 VDD.n8573 VSS 0.690489f
C28092 VDD.t3048 VSS 0.066856f
C28093 VDD.t4618 VSS 0.066856f
C28094 VDD.n8574 VSS 0.690489f
C28095 VDD.t1764 VSS 0.028519f
C28096 VDD.t3049 VSS 0.028519f
C28097 VDD.n8575 VSS 0.009191f
C28098 VDD.n8576 VSS 0.644755f
C28099 VDD.t2704 VSS 0.066856f
C28100 VDD.t4282 VSS 0.066856f
C28101 VDD.n8577 VSS 0.709674f
C28102 VDD.t1412 VSS 0.028519f
C28103 VDD.t2705 VSS 0.028519f
C28104 VDD.n8578 VSS 0.009191f
C28105 VDD.n8579 VSS 0.308318f
C28106 VDD.t4060 VSS 0.066856f
C28107 VDD.n8580 VSS 0.14405f
C28108 VDD.t3841 VSS 0.025104f
C28109 VDD.t4516 VSS 0.066856f
C28110 VDD.n8581 VSS 0.14405f
C28111 VDD.t3861 VSS 0.025104f
C28112 VDD.n8582 VSS 0.033925f
C28113 VDD.t1131 VSS 0.028519f
C28114 VDD.t4219 VSS 0.028519f
C28115 VDD.n8583 VSS 0.009191f
C28116 VDD.t1129 VSS 0.066856f
C28117 VDD.t3826 VSS 0.066856f
C28118 VDD.t1462 VSS 0.028519f
C28119 VDD.t4525 VSS 0.028519f
C28120 VDD.n8584 VSS 0.009191f
C28121 VDD.t1461 VSS 0.066856f
C28122 VDD.t4194 VSS 0.066856f
C28123 VDD.t2109 VSS 0.066856f
C28124 VDD.t613 VSS 0.066856f
C28125 VDD.t3601 VSS 0.066856f
C28126 VDD.t1022 VSS 0.066856f
C28127 VDD.n8585 VSS 0.690489f
C28128 VDD.t3058 VSS 0.066856f
C28129 VDD.t4524 VSS 0.066856f
C28130 VDD.n8586 VSS 0.690489f
C28131 VDD.t4195 VSS 0.028519f
C28132 VDD.t3059 VSS 0.028519f
C28133 VDD.n8587 VSS 0.009191f
C28134 VDD.n8588 VSS 0.644755f
C28135 VDD.t2716 VSS 0.066856f
C28136 VDD.t4218 VSS 0.066856f
C28137 VDD.n8589 VSS 0.709674f
C28138 VDD.t3827 VSS 0.028519f
C28139 VDD.t2717 VSS 0.028519f
C28140 VDD.n8590 VSS 0.009191f
C28141 VDD.n8591 VSS 0.308318f
C28142 VDD.t2346 VSS 0.066856f
C28143 VDD.n8592 VSS 0.14405f
C28144 VDD.t3851 VSS 0.025104f
C28145 VDD.t2384 VSS 0.066856f
C28146 VDD.n8593 VSS 0.14405f
C28147 VDD.t2101 VSS 0.025104f
C28148 VDD.t4454 VSS 0.066856f
C28149 VDD.n8594 VSS 0.14405f
C28150 VDD.t1853 VSS 0.025104f
C28151 VDD.t1709 VSS 0.066856f
C28152 VDD.n8595 VSS 0.14405f
C28153 VDD.t1490 VSS 0.025104f
C28154 VDD.t1509 VSS 0.028519f
C28155 VDD.t4149 VSS 0.028519f
C28156 VDD.n8596 VSS 0.009191f
C28157 VDD.t1507 VSS 0.066856f
C28158 VDD.t4246 VSS 0.066856f
C28159 VDD.t1876 VSS 0.028519f
C28160 VDD.t4471 VSS 0.028519f
C28161 VDD.n8597 VSS 0.009191f
C28162 VDD.t1875 VSS 0.066856f
C28163 VDD.t4548 VSS 0.066856f
C28164 VDD.t2599 VSS 0.066856f
C28165 VDD.t1049 VSS 0.066856f
C28166 VDD.t1235 VSS 0.066856f
C28167 VDD.t970 VSS 0.066856f
C28168 VDD.n8598 VSS 0.690489f
C28169 VDD.t622 VSS 0.066856f
C28170 VDD.t4470 VSS 0.066856f
C28171 VDD.n8599 VSS 0.690489f
C28172 VDD.t4549 VSS 0.028519f
C28173 VDD.t624 VSS 0.028519f
C28174 VDD.n8600 VSS 0.009191f
C28175 VDD.n8601 VSS 0.644755f
C28176 VDD.t4440 VSS 0.066856f
C28177 VDD.t4148 VSS 0.066856f
C28178 VDD.n8602 VSS 0.709674f
C28179 VDD.t4247 VSS 0.028519f
C28180 VDD.t4441 VSS 0.028519f
C28181 VDD.n8603 VSS 0.009191f
C28182 VDD.n8604 VSS 0.308318f
C28183 VDD.t2789 VSS 0.066856f
C28184 VDD.n8605 VSS 0.14405f
C28185 VDD.t4261 VSS 0.025104f
C28186 VDD.t1633 VSS 0.066856f
C28187 VDD.n8606 VSS 0.14405f
C28188 VDD.t1406 VSS 0.025104f
C28189 VDD.n8607 VSS 0.033925f
C28190 VDD.t2684 VSS 0.066856f
C28191 VDD.n8608 VSS 0.14405f
C28192 VDD.t4183 VSS 0.025104f
C28193 VDD.t4048 VSS 0.066856f
C28194 VDD.n8609 VSS 0.14405f
C28195 VDD.t3819 VSS 0.025104f
C28196 VDD.t3843 VSS 0.028519f
C28197 VDD.t4065 VSS 0.028519f
C28198 VDD.n8610 VSS 0.009191f
C28199 VDD.t3842 VSS 0.066856f
C28200 VDD.t3468 VSS 0.066856f
C28201 VDD.t4213 VSS 0.028519f
C28202 VDD.t4391 VSS 0.028519f
C28203 VDD.n8611 VSS 0.009191f
C28204 VDD.t4212 VSS 0.066856f
C28205 VDD.t3800 VSS 0.066856f
C28206 VDD.t638 VSS 0.066856f
C28207 VDD.t4400 VSS 0.066856f
C28208 VDD.t1650 VSS 0.066856f
C28209 VDD.t893 VSS 0.066856f
C28210 VDD.n8612 VSS 0.696076f
C28211 VDD.t1059 VSS 0.066856f
C28212 VDD.t4390 VSS 0.066856f
C28213 VDD.n8613 VSS 0.696076f
C28214 VDD.t3801 VSS 0.028519f
C28215 VDD.t1060 VSS 0.028519f
C28216 VDD.n8614 VSS 0.009191f
C28217 VDD.n8615 VSS 0.650522f
C28218 VDD.t688 VSS 0.066856f
C28219 VDD.t4064 VSS 0.066856f
C28220 VDD.n8616 VSS 0.715442f
C28221 VDD.t3469 VSS 0.028519f
C28222 VDD.t690 VSS 0.028519f
C28223 VDD.n8617 VSS 0.009191f
C28224 VDD.n8618 VSS 0.310925f
C28225 VDD.t3681 VSS 0.066856f
C28226 VDD.n8619 VSS 0.14405f
C28227 VDD.t731 VSS 0.025104f
C28228 VDD.t3346 VSS 0.066856f
C28229 VDD.n8620 VSS 0.14405f
C28230 VDD.t767 VSS 0.025104f
C28231 VDD.t1905 VSS 0.066856f
C28232 VDD.n8621 VSS 0.14405f
C28233 VDD.t2736 VSS 0.025104f
C28234 VDD.t1541 VSS 0.066856f
C28235 VDD.n8622 VSS 0.14405f
C28236 VDD.t3191 VSS 0.025104f
C28237 VDD.n8623 VSS 0.033925f
C28238 VDD.t3125 VSS 0.028519f
C28239 VDD.t1573 VSS 0.028519f
C28240 VDD.n8624 VSS 0.009191f
C28241 VDD.t3124 VSS 0.066856f
C28242 VDD.t2996 VSS 0.066856f
C28243 VDD.t3439 VSS 0.028519f
C28244 VDD.t1941 VSS 0.028519f
C28245 VDD.n8625 VSS 0.009191f
C28246 VDD.t3438 VSS 0.066856f
C28247 VDD.t3298 VSS 0.066856f
C28248 VDD.t4044 VSS 0.066856f
C28249 VDD.t3872 VSS 0.066856f
C28250 VDD.t2864 VSS 0.066856f
C28251 VDD.t2653 VSS 0.066856f
C28252 VDD.n8626 VSS 0.690489f
C28253 VDD.t2184 VSS 0.066856f
C28254 VDD.t1940 VSS 0.066856f
C28255 VDD.n8627 VSS 0.690489f
C28256 VDD.t3299 VSS 0.028519f
C28257 VDD.t2185 VSS 0.028519f
C28258 VDD.n8628 VSS 0.009191f
C28259 VDD.n8629 VSS 0.644755f
C28260 VDD.t1781 VSS 0.066856f
C28261 VDD.t1571 VSS 0.066856f
C28262 VDD.n8630 VSS 0.709674f
C28263 VDD.t2997 VSS 0.028519f
C28264 VDD.t1783 VSS 0.028519f
C28265 VDD.n8631 VSS 0.009191f
C28266 VDD.n8632 VSS 0.308318f
C28267 VDD.t1809 VSS 0.066856f
C28268 VDD.n8633 VSS 0.14405f
C28269 VDD.t2642 VSS 0.025104f
C28270 VDD.t2641 VSS 0.066856f
C28271 VDD.n8634 VSS 0.14405f
C28272 VDD.n8635 VSS 0.120118f
C28273 VDD.n8636 VSS 0.016021f
C28274 VDD.t1810 VSS 0.025104f
C28275 VDD.n8637 VSS 0.116823f
C28276 VDD.n8638 VSS 0.766371f
C28277 VDD.n8639 VSS 0.04911f
C28278 VDD.t543 VSS 0.018805f
C28279 VDD.t541 VSS 0.019767f
C28280 VDD.n8640 VSS 0.054793f
C28281 VDD.t540 VSS 0.019781f
C28282 VDD.t542 VSS 0.018792f
C28283 VDD.n8641 VSS 0.077486f
C28284 VDD.n8642 VSS 0.252514f
C28285 VDD.n8643 VSS 0.199549f
C28286 VDD.n8644 VSS 0.060108f
C28287 VDD.t3190 VSS 0.066856f
C28288 VDD.n8645 VSS 0.131361f
C28289 VDD.n8646 VSS 0.120118f
C28290 VDD.n8647 VSS 0.016021f
C28291 VDD.t1543 VSS 0.025104f
C28292 VDD.n8648 VSS 0.105404f
C28293 VDD.n8649 VSS 0.057098f
C28294 VDD.n8650 VSS 0.087217f
C28295 VDD.t2735 VSS 0.066856f
C28296 VDD.n8651 VSS 0.14405f
C28297 VDD.n8652 VSS 0.120118f
C28298 VDD.n8653 VSS 0.016021f
C28299 VDD.t1907 VSS 0.025104f
C28300 VDD.n8654 VSS 0.116823f
C28301 VDD.t3209 VSS 0.028519f
C28302 VDD.t3372 VSS 0.028519f
C28303 VDD.n8655 VSS 0.009191f
C28304 VDD.t3208 VSS 0.066856f
C28305 VDD.t3064 VSS 0.066856f
C28306 VDD.t3509 VSS 0.028519f
C28307 VDD.t3720 VSS 0.028519f
C28308 VDD.n8656 VSS 0.009191f
C28309 VDD.t3508 VSS 0.066856f
C28310 VDD.t3357 VSS 0.066856f
C28311 VDD.t4134 VSS 0.066856f
C28312 VDD.t3974 VSS 0.066856f
C28313 VDD.t2960 VSS 0.066856f
C28314 VDD.t4328 VSS 0.066856f
C28315 VDD.n8657 VSS 0.690489f
C28316 VDD.t2288 VSS 0.066856f
C28317 VDD.t3719 VSS 0.066856f
C28318 VDD.n8658 VSS 0.690489f
C28319 VDD.t3358 VSS 0.028519f
C28320 VDD.t2289 VSS 0.028519f
C28321 VDD.n8659 VSS 0.009191f
C28322 VDD.n8660 VSS 0.644755f
C28323 VDD.t1885 VSS 0.066856f
C28324 VDD.t3371 VSS 0.066856f
C28325 VDD.n8661 VSS 0.709674f
C28326 VDD.t3065 VSS 0.028519f
C28327 VDD.t1887 VSS 0.028519f
C28328 VDD.n8662 VSS 0.009191f
C28329 VDD.n8663 VSS 0.308318f
C28330 VDD.n8664 VSS 0.779905f
C28331 VDD.n8665 VSS 0.116823f
C28332 VDD.t766 VSS 0.066856f
C28333 VDD.n8666 VSS 0.14405f
C28334 VDD.n8667 VSS 0.120118f
C28335 VDD.n8668 VSS 0.016021f
C28336 VDD.t3347 VSS 0.025104f
C28337 VDD.n8669 VSS 0.105404f
C28338 VDD.n8670 VSS 0.057098f
C28339 VDD.n8671 VSS 0.087217f
C28340 VDD.t730 VSS 0.066856f
C28341 VDD.n8672 VSS 0.14405f
C28342 VDD.n8673 VSS 0.120118f
C28343 VDD.n8674 VSS 0.016021f
C28344 VDD.t3682 VSS 0.025104f
C28345 VDD.n8675 VSS 0.116823f
C28346 VDD.n8676 VSS 0.78631f
C28347 VDD.n8677 VSS 0.116823f
C28348 VDD.t3818 VSS 0.066856f
C28349 VDD.n8678 VSS 0.14405f
C28350 VDD.n8679 VSS 0.120118f
C28351 VDD.n8680 VSS 0.016021f
C28352 VDD.t4049 VSS 0.025104f
C28353 VDD.n8681 VSS 0.105404f
C28354 VDD.n8682 VSS 0.057098f
C28355 VDD.n8683 VSS 0.087217f
C28356 VDD.t4182 VSS 0.066856f
C28357 VDD.n8684 VSS 0.14405f
C28358 VDD.n8685 VSS 0.120118f
C28359 VDD.n8686 VSS 0.016021f
C28360 VDD.t2685 VSS 0.025104f
C28361 VDD.n8687 VSS 0.116823f
C28362 VDD.t1428 VSS 0.028519f
C28363 VDD.t1656 VSS 0.028519f
C28364 VDD.n8688 VSS 0.009191f
C28365 VDD.t1426 VSS 0.066856f
C28366 VDD.t4166 VSS 0.066856f
C28367 VDD.t1778 VSS 0.028519f
C28368 VDD.t2036 VSS 0.028519f
C28369 VDD.n8689 VSS 0.009191f
C28370 VDD.t1777 VSS 0.066856f
C28371 VDD.t4482 VSS 0.066856f
C28372 VDD.t2512 VSS 0.066856f
C28373 VDD.t986 VSS 0.066856f
C28374 VDD.t1155 VSS 0.066856f
C28375 VDD.t2724 VSS 0.066856f
C28376 VDD.n8690 VSS 0.690489f
C28377 VDD.t4704 VSS 0.066856f
C28378 VDD.t2035 VSS 0.066856f
C28379 VDD.n8691 VSS 0.690489f
C28380 VDD.t4483 VSS 0.028519f
C28381 VDD.t4705 VSS 0.028519f
C28382 VDD.n8692 VSS 0.009191f
C28383 VDD.n8693 VSS 0.644755f
C28384 VDD.t4354 VSS 0.066856f
C28385 VDD.t1654 VSS 0.066856f
C28386 VDD.n8694 VSS 0.709674f
C28387 VDD.t4167 VSS 0.028519f
C28388 VDD.t4355 VSS 0.028519f
C28389 VDD.n8695 VSS 0.009191f
C28390 VDD.n8696 VSS 0.308318f
C28391 VDD.n8697 VSS 0.766371f
C28392 VDD.n8698 VSS 0.04911f
C28393 VDD.t4787 VSS 0.018805f
C28394 VDD.t4788 VSS 0.019767f
C28395 VDD.n8699 VSS 0.054793f
C28396 VDD.t4786 VSS 0.019781f
C28397 VDD.t4789 VSS 0.018792f
C28398 VDD.n8700 VSS 0.077486f
C28399 VDD.n8701 VSS 0.252514f
C28400 VDD.n8702 VSS 0.199549f
C28401 VDD.n8703 VSS 0.060108f
C28402 VDD.t1405 VSS 0.066856f
C28403 VDD.n8704 VSS 0.131361f
C28404 VDD.n8705 VSS 0.120118f
C28405 VDD.n8706 VSS 0.016021f
C28406 VDD.t1634 VSS 0.025104f
C28407 VDD.n8707 VSS 0.105404f
C28408 VDD.n8708 VSS 0.057098f
C28409 VDD.n8709 VSS 0.087217f
C28410 VDD.t4260 VSS 0.066856f
C28411 VDD.n8710 VSS 0.14405f
C28412 VDD.n8711 VSS 0.120118f
C28413 VDD.n8712 VSS 0.016021f
C28414 VDD.t2790 VSS 0.025104f
C28415 VDD.n8713 VSS 0.116823f
C28416 VDD.n8714 VSS 0.779905f
C28417 VDD.n8715 VSS 0.116823f
C28418 VDD.t1488 VSS 0.066856f
C28419 VDD.n8716 VSS 0.14405f
C28420 VDD.n8717 VSS 0.120118f
C28421 VDD.n8718 VSS 0.016021f
C28422 VDD.t1711 VSS 0.025104f
C28423 VDD.n8719 VSS 0.105404f
C28424 VDD.n8720 VSS 0.057098f
C28425 VDD.n8721 VSS 0.087217f
C28426 VDD.t1851 VSS 0.066856f
C28427 VDD.n8722 VSS 0.14405f
C28428 VDD.n8723 VSS 0.120118f
C28429 VDD.n8724 VSS 0.016021f
C28430 VDD.t4455 VSS 0.025104f
C28431 VDD.n8725 VSS 0.116823f
C28432 VDD.t1056 VSS 0.028519f
C28433 VDD.t3631 VSS 0.028519f
C28434 VDD.n8726 VSS 0.009191f
C28435 VDD.t1054 VSS 0.066856f
C28436 VDD.t1822 VSS 0.066856f
C28437 VDD.t1386 VSS 0.028519f
C28438 VDD.t4009 VSS 0.028519f
C28439 VDD.n8727 VSS 0.009191f
C28440 VDD.t1385 VSS 0.066856f
C28441 VDD.t2221 VSS 0.066856f
C28442 VDD.t2014 VSS 0.066856f
C28443 VDD.t2892 VSS 0.066856f
C28444 VDD.t3096 VSS 0.066856f
C28445 VDD.t4586 VSS 0.066856f
C28446 VDD.n8728 VSS 0.696076f
C28447 VDD.t2496 VSS 0.066856f
C28448 VDD.t4008 VSS 0.066856f
C28449 VDD.n8729 VSS 0.696076f
C28450 VDD.t2222 VSS 0.028519f
C28451 VDD.t2497 VSS 0.028519f
C28452 VDD.n8730 VSS 0.009191f
C28453 VDD.n8731 VSS 0.650522f
C28454 VDD.t2078 VSS 0.066856f
C28455 VDD.t3630 VSS 0.066856f
C28456 VDD.n8732 VSS 0.715442f
C28457 VDD.t1824 VSS 0.028519f
C28458 VDD.t2080 VSS 0.028519f
C28459 VDD.n8733 VSS 0.009191f
C28460 VDD.n8734 VSS 0.310925f
C28461 VDD.n8735 VSS 0.78631f
C28462 VDD.n8736 VSS 0.116823f
C28463 VDD.t2099 VSS 0.066856f
C28464 VDD.n8737 VSS 0.14405f
C28465 VDD.n8738 VSS 0.120118f
C28466 VDD.n8739 VSS 0.016021f
C28467 VDD.t2386 VSS 0.025104f
C28468 VDD.n8740 VSS 0.105404f
C28469 VDD.n8741 VSS 0.057098f
C28470 VDD.n8742 VSS 0.087217f
C28471 VDD.t3850 VSS 0.066856f
C28472 VDD.n8743 VSS 0.14405f
C28473 VDD.n8744 VSS 0.120118f
C28474 VDD.n8745 VSS 0.016021f
C28475 VDD.t2348 VSS 0.025104f
C28476 VDD.n8746 VSS 0.116823f
C28477 VDD.n8747 VSS 0.766371f
C28478 VDD.n8748 VSS 0.04911f
C28479 VDD.t300 VSS 0.018805f
C28480 VDD.t298 VSS 0.019767f
C28481 VDD.n8749 VSS 0.054793f
C28482 VDD.t299 VSS 0.019781f
C28483 VDD.t297 VSS 0.018792f
C28484 VDD.n8750 VSS 0.077486f
C28485 VDD.n8751 VSS 0.252514f
C28486 VDD.n8752 VSS 0.199549f
C28487 VDD.n8753 VSS 0.060108f
C28488 VDD.t3860 VSS 0.066856f
C28489 VDD.n8754 VSS 0.131361f
C28490 VDD.n8755 VSS 0.120118f
C28491 VDD.n8756 VSS 0.016021f
C28492 VDD.t4517 VSS 0.025104f
C28493 VDD.n8757 VSS 0.105404f
C28494 VDD.n8758 VSS 0.057098f
C28495 VDD.n8759 VSS 0.087217f
C28496 VDD.t3840 VSS 0.066856f
C28497 VDD.n8760 VSS 0.14405f
C28498 VDD.n8761 VSS 0.120118f
C28499 VDD.n8762 VSS 0.016021f
C28500 VDD.t4061 VSS 0.025104f
C28501 VDD.n8763 VSS 0.116823f
C28502 VDD.n8764 VSS 0.779905f
C28503 VDD.n8765 VSS 0.116823f
C28504 VDD.t3958 VSS 0.066856f
C28505 VDD.n8766 VSS 0.14405f
C28506 VDD.n8767 VSS 0.120118f
C28507 VDD.n8768 VSS 0.016021f
C28508 VDD.t2943 VSS 0.025104f
C28509 VDD.n8769 VSS 0.105404f
C28510 VDD.t3934 VSS 0.066856f
C28511 VDD.n8770 VSS 0.14405f
C28512 VDD.t4585 VSS 0.025104f
C28513 VDD.t3470 VSS 0.066856f
C28514 VDD.n8771 VSS 0.14405f
C28515 VDD.t2440 VSS 0.025104f
C28516 VDD.t2439 VSS 0.066856f
C28517 VDD.n8772 VSS 0.14405f
C28518 VDD.n8773 VSS 0.120118f
C28519 VDD.n8774 VSS 0.016021f
C28520 VDD.t3471 VSS 0.025104f
C28521 VDD.n8775 VSS 0.116823f
C28522 VDD.t3165 VSS 0.028519f
C28523 VDD.t2468 VSS 0.028519f
C28524 VDD.n8776 VSS 0.009191f
C28525 VDD.t3164 VSS 0.066856f
C28526 VDD.t1491 VSS 0.066856f
C28527 VDD.t3477 VSS 0.028519f
C28528 VDD.t2823 VSS 0.028519f
C28529 VDD.n8777 VSS 0.009191f
C28530 VDD.t3476 VSS 0.066856f
C28531 VDD.t1858 VSS 0.066856f
C28532 VDD.t4084 VSS 0.066856f
C28533 VDD.t2579 VSS 0.066856f
C28534 VDD.t4085 VSS 0.028519f
C28535 VDD.t3362 VSS 0.028519f
C28536 VDD.n8778 VSS 0.009191f
C28537 VDD.t3497 VSS 0.028519f
C28538 VDD.t2839 VSS 0.028519f
C28539 VDD.n8779 VSS 0.009191f
C28540 VDD.t3496 VSS 0.066856f
C28541 VDD.t1879 VSS 0.066856f
C28542 VDD.t3854 VSS 0.066856f
C28543 VDD.t2319 VSS 0.066856f
C28544 VDD.t3855 VSS 0.028519f
C28545 VDD.t3187 VSS 0.028519f
C28546 VDD.n8780 VSS 0.009191f
C28547 VDD.t1267 VSS 0.066856f
C28548 VDD.t3866 VSS 0.066856f
C28549 VDD.t1335 VSS 0.066856f
C28550 VDD.t4708 VSS 0.066856f
C28551 VDD.n8781 VSS 0.715442f
C28552 VDD.t2320 VSS 0.028519f
C28553 VDD.t3937 VSS 0.028519f
C28554 VDD.n8782 VSS 0.009191f
C28555 VDD.n8783 VSS 0.650522f
C28556 VDD.t3936 VSS 0.066856f
C28557 VDD.t3186 VSS 0.066856f
C28558 VDD.n8784 VSS 0.696076f
C28559 VDD.t3548 VSS 0.066856f
C28560 VDD.t2838 VSS 0.066856f
C28561 VDD.n8785 VSS 0.696076f
C28562 VDD.t1880 VSS 0.028519f
C28563 VDD.t3549 VSS 0.028519f
C28564 VDD.n8786 VSS 0.009191f
C28565 VDD.n8787 VSS 0.528101f
C28566 VDD.n8788 VSS 0.529799f
C28567 VDD.t2580 VSS 0.028519f
C28568 VDD.t4171 VSS 0.028519f
C28569 VDD.n8789 VSS 0.009191f
C28570 VDD.n8790 VSS 0.475536f
C28571 VDD.t4170 VSS 0.066856f
C28572 VDD.t3361 VSS 0.066856f
C28573 VDD.n8791 VSS 0.696076f
C28574 VDD.t3538 VSS 0.066856f
C28575 VDD.t2822 VSS 0.066856f
C28576 VDD.n8792 VSS 0.696076f
C28577 VDD.t1859 VSS 0.028519f
C28578 VDD.t3539 VSS 0.028519f
C28579 VDD.n8793 VSS 0.009191f
C28580 VDD.n8794 VSS 0.650522f
C28581 VDD.t3236 VSS 0.066856f
C28582 VDD.t2466 VSS 0.066856f
C28583 VDD.n8795 VSS 0.715442f
C28584 VDD.t1493 VSS 0.028519f
C28585 VDD.t3237 VSS 0.028519f
C28586 VDD.n8796 VSS 0.009191f
C28587 VDD.n8797 VSS 0.310925f
C28588 VDD.n8798 VSS 0.78631f
C28589 VDD.n8799 VSS 0.116823f
C28590 VDD.t4584 VSS 0.066856f
C28591 VDD.n8800 VSS 0.14405f
C28592 VDD.n8801 VSS 0.120118f
C28593 VDD.n8802 VSS 0.016021f
C28594 VDD.t3935 VSS 0.025104f
C28595 VDD.n8803 VSS 0.087217f
C28596 VDD.n8804 VSS 0.057098f
C28597 VDD.n8805 VSS 0.208771f
C28598 VDD.n8806 VSS 0.595476f
C28599 VDD.n8807 VSS 0.645798f
C28600 VDD.n8808 VSS 0.206947f
C28601 VDD.n8809 VSS 0.048151f
C28602 VDD.n8810 VSS 0.083673f
C28603 VDD.t2111 VSS 0.066856f
C28604 VDD.n8811 VSS 0.125227f
C28605 VDD.n8812 VSS 0.006598f
C28606 VDD.n8813 VSS 0.010188f
C28607 VDD.t7 VSS 0.020387f
C28608 VDD.t10 VSS 0.022137f
C28609 VDD.n8814 VSS 0.069721f
C28610 VDD.n8815 VSS 0.040089f
C28611 VDD.t5 VSS 0.022115f
C28612 VDD.t11 VSS 0.020371f
C28613 VDD.n8816 VSS 0.027128f
C28614 VDD.n8817 VSS 0.036577f
C28615 VDD.n8818 VSS 0.044801f
C28616 VDD.n8819 VSS 0.278297f
C28617 VDD.n8820 VSS 0.040089f
C28618 VDD.t8 VSS 0.020387f
C28619 VDD.n8821 VSS 0.049653f
C28620 VDD.t9 VSS 0.017093f
C28621 VDD.n8822 VSS 0.042104f
C28622 VDD.n8823 VSS 0.069461f
C28623 VDD.t4 VSS 0.017093f
C28624 VDD.n8824 VSS 0.035483f
C28625 VDD.t2 VSS 0.020371f
C28626 VDD.n8825 VSS 0.027128f
C28627 VDD.n8826 VSS 0.016538f
C28628 VDD.n8827 VSS 0.027213f
C28629 VDD.n8828 VSS 0.204333f
C28630 VDD.n8829 VSS 0.030906f
C28631 VDD.t2870 VSS 0.066856f
C28632 VDD.n8830 VSS 0.045867f
C28633 VDD.n8831 VSS 0.015693f
C28634 VDD.n8832 VSS 0.010881f
C28635 VDD.n8833 VSS 0.044227f
C28636 VDD.n8834 VSS 0.094696f
C28637 VDD.n8835 VSS 0.016021f
C28638 VDD.t2871 VSS 0.025104f
C28639 VDD.n8836 VSS 0.08403f
C28640 VDD.n8837 VSS 0.62638f
C28641 VDD.n8838 VSS 0.099723f
C28642 VDD.t1619 VSS 0.066856f
C28643 VDD.n8839 VSS 0.125227f
C28644 VDD.n8840 VSS 0.101294f
C28645 VDD.n8841 VSS 0.016021f
C28646 VDD.t4693 VSS 0.025104f
C28647 VDD.n8842 VSS 0.081176f
C28648 VDD.t1592 VSS 0.066856f
C28649 VDD.n8843 VSS 0.125227f
C28650 VDD.t581 VSS 0.025104f
C28651 VDD.t2213 VSS 0.066856f
C28652 VDD.n8844 VSS 0.125227f
C28653 VDD.t600 VSS 0.025104f
C28654 VDD.t599 VSS 0.066856f
C28655 VDD.n8845 VSS 0.125227f
C28656 VDD.n8846 VSS 0.101294f
C28657 VDD.n8847 VSS 0.016021f
C28658 VDD.t2214 VSS 0.025104f
C28659 VDD.n8848 VSS 0.099723f
C28660 VDD.t3650 VSS 0.066856f
C28661 VDD.t2102 VSS 0.066856f
C28662 VDD.t1017 VSS 0.066856f
C28663 VDD.t2554 VSS 0.066856f
C28664 VDD.n8849 VSS 0.709674f
C28665 VDD.t4033 VSS 0.028519f
C28666 VDD.t2903 VSS 0.028519f
C28667 VDD.n8850 VSS 0.009191f
C28668 VDD.t2535 VSS 0.028519f
C28669 VDD.t1334 VSS 0.028519f
C28670 VDD.n8851 VSS 0.009191f
C28671 VDD.n8852 VSS 0.644755f
C28672 VDD.t4032 VSS 0.066856f
C28673 VDD.t2534 VSS 0.066856f
C28674 VDD.t1333 VSS 0.066856f
C28675 VDD.t2902 VSS 0.066856f
C28676 VDD.n8853 VSS 0.690489f
C28677 VDD.t4612 VSS 0.066856f
C28678 VDD.t3130 VSS 0.066856f
C28679 VDD.t1973 VSS 0.066856f
C28680 VDD.t3460 VSS 0.066856f
C28681 VDD.n8854 VSS 0.690489f
C28682 VDD.t4613 VSS 0.028519f
C28683 VDD.t3461 VSS 0.028519f
C28684 VDD.n8855 VSS 0.009191f
C28685 VDD.t3131 VSS 0.028519f
C28686 VDD.t1974 VSS 0.028519f
C28687 VDD.n8856 VSS 0.009191f
C28688 VDD.n8857 VSS 0.471397f
C28689 VDD.n8858 VSS 0.524869f
C28690 VDD.t4047 VSS 0.028519f
C28691 VDD.t2915 VSS 0.028519f
C28692 VDD.n8859 VSS 0.009191f
C28693 VDD.t2553 VSS 0.028519f
C28694 VDD.t1355 VSS 0.028519f
C28695 VDD.n8860 VSS 0.009191f
C28696 VDD.n8861 VSS 0.523473f
C28697 VDD.t4046 VSS 0.066856f
C28698 VDD.t2552 VSS 0.066856f
C28699 VDD.t1354 VSS 0.066856f
C28700 VDD.t2914 VSS 0.066856f
C28701 VDD.n8862 VSS 0.690489f
C28702 VDD.t4388 VSS 0.066856f
C28703 VDD.t2920 VSS 0.066856f
C28704 VDD.t1726 VSS 0.066856f
C28705 VDD.t3276 VSS 0.066856f
C28706 VDD.n8863 VSS 0.690489f
C28707 VDD.t4389 VSS 0.028519f
C28708 VDD.t3277 VSS 0.028519f
C28709 VDD.n8864 VSS 0.009191f
C28710 VDD.t2921 VSS 0.028519f
C28711 VDD.t1727 VSS 0.028519f
C28712 VDD.n8865 VSS 0.009191f
C28713 VDD.n8866 VSS 0.644755f
C28714 VDD.t1819 VSS 0.066856f
C28715 VDD.t4416 VSS 0.066856f
C28716 VDD.t3348 VSS 0.066856f
C28717 VDD.t633 VSS 0.066856f
C28718 VDD.n8867 VSS 0.709674f
C28719 VDD.t1821 VSS 0.028519f
C28720 VDD.t635 VSS 0.028519f
C28721 VDD.n8868 VSS 0.009191f
C28722 VDD.t4417 VSS 0.028519f
C28723 VDD.t3349 VSS 0.028519f
C28724 VDD.n8869 VSS 0.009191f
C28725 VDD.n8870 VSS 0.261039f
C28726 VDD.n8871 VSS 0.62132f
C28727 VDD.n8872 VSS 0.099723f
C28728 VDD.t580 VSS 0.066856f
C28729 VDD.n8873 VSS 0.125227f
C28730 VDD.n8874 VSS 0.101294f
C28731 VDD.n8875 VSS 0.016021f
C28732 VDD.t1593 VSS 0.025104f
C28733 VDD.n8876 VSS 0.083673f
C28734 VDD.n8877 VSS 0.048151f
C28735 VDD.n8878 VSS 0.206947f
C28736 VDD.n8879 VSS 0.645798f
C28737 VDD.t334 VSS 1.96535f
C28738 VDD.t634 VSS 1.96535f
C28739 VDD.t1820 VSS 1.45794f
C28740 VDD.n8880 VSS 0.865258f
C28741 VDD.n8881 VSS 0.865258f
C28742 VDD.t1018 VSS 1.45794f
C28743 VDD.t2103 VSS 1.96535f
C28744 VDD.t544 VSS 1.96535f
C28745 VDD.t546 VSS 1.31955f
C28746 VDD.n8882 VSS 0.595476f
C28747 VDD.n8883 VSS 0.208771f
C28748 VDD.n8884 VSS 0.057098f
C28749 VDD.n8885 VSS 0.087217f
C28750 VDD.t3446 VSS 0.066856f
C28751 VDD.n8886 VSS 0.14405f
C28752 VDD.n8887 VSS 0.120118f
C28753 VDD.n8888 VSS 0.016021f
C28754 VDD.t2523 VSS 0.025104f
C28755 VDD.n8889 VSS 0.116823f
C28756 VDD.n8890 VSS 0.766371f
C28757 VDD.n8891 VSS 0.04911f
C28758 VDD.t522 VSS 0.018805f
C28759 VDD.t520 VSS 0.019767f
C28760 VDD.n8892 VSS 0.054793f
C28761 VDD.t523 VSS 0.019781f
C28762 VDD.t521 VSS 0.018792f
C28763 VDD.n8893 VSS 0.077486f
C28764 VDD.n8894 VSS 0.252514f
C28765 VDD.n8895 VSS 0.199549f
C28766 VDD.n8896 VSS 0.060108f
C28767 VDD.t4018 VSS 0.066856f
C28768 VDD.n8897 VSS 0.131361f
C28769 VDD.n8898 VSS 0.120118f
C28770 VDD.n8899 VSS 0.016021f
C28771 VDD.t2531 VSS 0.025104f
C28772 VDD.n8900 VSS 0.105404f
C28773 VDD.t3526 VSS 0.066856f
C28774 VDD.n8901 VSS 0.14405f
C28775 VDD.t4227 VSS 0.025104f
C28776 VDD.t4110 VSS 0.066856f
C28777 VDD.n8902 VSS 0.14405f
C28778 VDD.t2626 VSS 0.025104f
C28779 VDD.t2625 VSS 0.066856f
C28780 VDD.n8903 VSS 0.14405f
C28781 VDD.n8904 VSS 0.120118f
C28782 VDD.n8905 VSS 0.016021f
C28783 VDD.t4111 VSS 0.025104f
C28784 VDD.n8906 VSS 0.116823f
C28785 VDD.t1255 VSS 0.028519f
C28786 VDD.t4251 VSS 0.028519f
C28787 VDD.n8907 VSS 0.009191f
C28788 VDD.t1253 VSS 0.066856f
C28789 VDD.t3868 VSS 0.066856f
C28790 VDD.t1609 VSS 0.028519f
C28791 VDD.t4557 VSS 0.028519f
C28792 VDD.n8908 VSS 0.009191f
C28793 VDD.t1608 VSS 0.066856f
C28794 VDD.t4236 VSS 0.066856f
C28795 VDD.t2270 VSS 0.066856f
C28796 VDD.t669 VSS 0.066856f
C28797 VDD.t2271 VSS 0.028519f
C28798 VDD.t1058 VSS 0.028519f
C28799 VDD.n8909 VSS 0.009191f
C28800 VDD.t1628 VSS 0.028519f
C28801 VDD.t4581 VSS 0.028519f
C28802 VDD.n8910 VSS 0.009191f
C28803 VDD.t1627 VSS 0.066856f
C28804 VDD.t4248 VSS 0.066856f
C28805 VDD.t2020 VSS 0.066856f
C28806 VDD.t4590 VSS 0.066856f
C28807 VDD.t2021 VSS 0.028519f
C28808 VDD.t846 VSS 0.028519f
C28809 VDD.n8911 VSS 0.009191f
C28810 VDD.t3611 VSS 0.066856f
C28811 VDD.t2066 VSS 0.066856f
C28812 VDD.t981 VSS 0.066856f
C28813 VDD.t2506 VSS 0.066856f
C28814 VDD.n8912 VSS 0.709674f
C28815 VDD.t4591 VSS 0.028519f
C28816 VDD.t3531 VSS 0.028519f
C28817 VDD.n8913 VSS 0.009191f
C28818 VDD.n8914 VSS 0.644755f
C28819 VDD.t3530 VSS 0.066856f
C28820 VDD.t844 VSS 0.066856f
C28821 VDD.n8915 VSS 0.690489f
C28822 VDD.t3198 VSS 0.066856f
C28823 VDD.t4580 VSS 0.066856f
C28824 VDD.n8916 VSS 0.690489f
C28825 VDD.t4249 VSS 0.028519f
C28826 VDD.t3199 VSS 0.028519f
C28827 VDD.n8917 VSS 0.009191f
C28828 VDD.n8918 VSS 0.523473f
C28829 VDD.n8919 VSS 0.524869f
C28830 VDD.t671 VSS 0.028519f
C28831 VDD.t3746 VSS 0.028519f
C28832 VDD.n8920 VSS 0.009191f
C28833 VDD.n8921 VSS 0.471397f
C28834 VDD.t3745 VSS 0.066856f
C28835 VDD.t1057 VSS 0.066856f
C28836 VDD.n8922 VSS 0.690489f
C28837 VDD.t3184 VSS 0.066856f
C28838 VDD.t4556 VSS 0.066856f
C28839 VDD.n8923 VSS 0.690489f
C28840 VDD.t4237 VSS 0.028519f
C28841 VDD.t3185 VSS 0.028519f
C28842 VDD.n8924 VSS 0.009191f
C28843 VDD.n8925 VSS 0.644755f
C28844 VDD.t2856 VSS 0.066856f
C28845 VDD.t4250 VSS 0.066856f
C28846 VDD.n8926 VSS 0.709674f
C28847 VDD.t3869 VSS 0.028519f
C28848 VDD.t2857 VSS 0.028519f
C28849 VDD.n8927 VSS 0.009191f
C28850 VDD.n8928 VSS 0.308318f
C28851 VDD.n8929 VSS 0.779905f
C28852 VDD.n8930 VSS 0.116823f
C28853 VDD.t4226 VSS 0.066856f
C28854 VDD.n8931 VSS 0.14405f
C28855 VDD.n8932 VSS 0.120118f
C28856 VDD.n8933 VSS 0.016021f
C28857 VDD.t3527 VSS 0.025104f
C28858 VDD.n8934 VSS 0.087217f
C28859 VDD.n8935 VSS 0.057098f
C28860 VDD.n8936 VSS 0.208771f
C28861 VDD.n8937 VSS 0.595476f
C28862 VDD.n8938 VSS 0.645798f
C28863 VDD.n8939 VSS 0.206947f
C28864 VDD.n8940 VSS 0.048151f
C28865 VDD.n8941 VSS 0.083673f
C28866 VDD.t1677 VSS 0.066856f
C28867 VDD.n8942 VSS 0.125227f
C28868 VDD.n8943 VSS 0.101294f
C28869 VDD.n8944 VSS 0.016021f
C28870 VDD.t2470 VSS 0.025104f
C28871 VDD.n8945 VSS 0.099723f
C28872 VDD.n8946 VSS 0.62132f
C28873 VDD.n8947 VSS 0.099723f
C28874 VDD.t2327 VSS 0.066856f
C28875 VDD.n8948 VSS 0.125227f
C28876 VDD.n8949 VSS 0.101294f
C28877 VDD.n8950 VSS 0.016021f
C28878 VDD.t711 VSS 0.025104f
C28879 VDD.n8951 VSS 0.081176f
C28880 VDD.t2290 VSS 0.066856f
C28881 VDD.n8952 VSS 0.125227f
C28882 VDD.t2562 VSS 0.025104f
C28883 VDD.n8953 VSS 0.006598f
C28884 VDD.t4802 VSS 0.020387f
C28885 VDD.t4805 VSS 0.022137f
C28886 VDD.n8954 VSS 0.069721f
C28887 VDD.n8955 VSS 0.040089f
C28888 VDD.t4801 VSS 0.022115f
C28889 VDD.t4806 VSS 0.020371f
C28890 VDD.n8956 VSS 0.027128f
C28891 VDD.n8957 VSS 0.036577f
C28892 VDD.n8958 VSS 0.044801f
C28893 VDD.n8959 VSS 0.278297f
C28894 VDD.n8960 VSS 0.040089f
C28895 VDD.t4803 VSS 0.020387f
C28896 VDD.n8961 VSS 0.049653f
C28897 VDD.t4804 VSS 0.017093f
C28898 VDD.n8962 VSS 0.042104f
C28899 VDD.n8963 VSS 0.069461f
C28900 VDD.t4800 VSS 0.017093f
C28901 VDD.n8964 VSS 0.035483f
C28902 VDD.t4807 VSS 0.020371f
C28903 VDD.n8965 VSS 0.027128f
C28904 VDD.n8966 VSS 0.016538f
C28905 VDD.n8967 VSS 0.027213f
C28906 VDD.n8968 VSS 0.204333f
C28907 VDD.n8969 VSS 0.030906f
C28908 VDD.t2560 VSS 0.066856f
C28909 VDD.n8970 VSS 0.045867f
C28910 VDD.t4178 VSS 0.066856f
C28911 VDD.n8971 VSS 0.125227f
C28912 VDD.t4367 VSS 0.025104f
C28913 VDD.t4366 VSS 0.066856f
C28914 VDD.n8972 VSS 0.125227f
C28915 VDD.n8973 VSS 0.101294f
C28916 VDD.n8974 VSS 0.016021f
C28917 VDD.t4179 VSS 0.025104f
C28918 VDD.n8975 VSS 0.099723f
C28919 VDD.t1825 VSS 0.066856f
C28920 VDD.t2733 VSS 0.066856f
C28921 VDD.t2950 VSS 0.066856f
C28922 VDD.t2081 VSS 0.066856f
C28923 VDD.n8976 VSS 0.715442f
C28924 VDD.t2226 VSS 0.028519f
C28925 VDD.t2505 VSS 0.028519f
C28926 VDD.n8977 VSS 0.009191f
C28927 VDD.t3071 VSS 0.028519f
C28928 VDD.t3273 VSS 0.028519f
C28929 VDD.n8978 VSS 0.009191f
C28930 VDD.n8979 VSS 0.650522f
C28931 VDD.t2225 VSS 0.066856f
C28932 VDD.t3070 VSS 0.066856f
C28933 VDD.t3272 VSS 0.066856f
C28934 VDD.t2504 VSS 0.066856f
C28935 VDD.n8980 VSS 0.696076f
C28936 VDD.t2894 VSS 0.066856f
C28937 VDD.t3616 VSS 0.066856f
C28938 VDD.t3832 VSS 0.066856f
C28939 VDD.t3100 VSS 0.066856f
C28940 VDD.n8981 VSS 0.696076f
C28941 VDD.t2895 VSS 0.028519f
C28942 VDD.t3101 VSS 0.028519f
C28943 VDD.n8982 VSS 0.009191f
C28944 VDD.t3617 VSS 0.028519f
C28945 VDD.t3833 VSS 0.028519f
C28946 VDD.n8983 VSS 0.009191f
C28947 VDD.n8984 VSS 0.475536f
C28948 VDD.n8985 VSS 0.529799f
C28949 VDD.t2241 VSS 0.028519f
C28950 VDD.t2519 VSS 0.028519f
C28951 VDD.n8986 VSS 0.009191f
C28952 VDD.t3085 VSS 0.028519f
C28953 VDD.t3281 VSS 0.028519f
C28954 VDD.n8987 VSS 0.009191f
C28955 VDD.n8988 VSS 0.528101f
C28956 VDD.t2240 VSS 0.066856f
C28957 VDD.t3084 VSS 0.066856f
C28958 VDD.t3280 VSS 0.066856f
C28959 VDD.t2518 VSS 0.066856f
C28960 VDD.n8989 VSS 0.696076f
C28961 VDD.t2677 VSS 0.066856f
C28962 VDD.t3407 VSS 0.066856f
C28963 VDD.t3605 VSS 0.066856f
C28964 VDD.t2884 VSS 0.066856f
C28965 VDD.n8990 VSS 0.696076f
C28966 VDD.t2678 VSS 0.028519f
C28967 VDD.t2885 VSS 0.028519f
C28968 VDD.n8991 VSS 0.009191f
C28969 VDD.t3408 VSS 0.028519f
C28970 VDD.t3606 VSS 0.028519f
C28971 VDD.n8992 VSS 0.009191f
C28972 VDD.n8993 VSS 0.650522f
C28973 VDD.t4202 VSS 0.066856f
C28974 VDD.t838 VSS 0.066856f
C28975 VDD.t1044 VSS 0.066856f
C28976 VDD.t4384 VSS 0.066856f
C28977 VDD.n8994 VSS 0.715442f
C28978 VDD.t4203 VSS 0.028519f
C28979 VDD.t4385 VSS 0.028519f
C28980 VDD.n8995 VSS 0.009191f
C28981 VDD.t840 VSS 0.028519f
C28982 VDD.t1046 VSS 0.028519f
C28983 VDD.n8996 VSS 0.009191f
C28984 VDD.n8997 VSS 0.263202f
C28985 VDD.n8998 VSS 0.62638f
C28986 VDD.n8999 VSS 0.08403f
C28987 VDD.n9000 VSS 0.010188f
C28988 VDD.n9001 VSS 0.035132f
C28989 VDD.n9002 VSS 0.015693f
C28990 VDD.n9003 VSS 0.010881f
C28991 VDD.n9004 VSS 0.044227f
C28992 VDD.n9005 VSS 0.094696f
C28993 VDD.n9006 VSS 0.016021f
C28994 VDD.t2292 VSS 0.025104f
C28995 VDD.n9007 VSS 0.083673f
C28996 VDD.n9008 VSS 0.048151f
C28997 VDD.n9009 VSS 0.206947f
C28998 VDD.n9010 VSS 0.645798f
C28999 VDD.t1798 VSS 1.96535f
C29000 VDD.t2082 VSS 1.96535f
C29001 VDD.t1826 VSS 1.45794f
C29002 VDD.n9011 VSS 0.902999f
C29003 VDD.n9012 VSS 0.902999f
C29004 VDD.t1045 VSS 1.45794f
C29005 VDD.t839 VSS 1.96535f
C29006 VDD.t2561 VSS 1.96535f
C29007 VDD.t2291 VSS 1.31955f
C29008 VDD.n9013 VSS 0.595476f
C29009 VDD.n9014 VSS 0.208771f
C29010 VDD.n9015 VSS 0.057098f
C29011 VDD.n9016 VSS 0.087217f
C29012 VDD.t4082 VSS 0.066856f
C29013 VDD.n9017 VSS 0.14405f
C29014 VDD.n9018 VSS 0.120118f
C29015 VDD.n9019 VSS 0.016021f
C29016 VDD.t4291 VSS 0.025104f
C29017 VDD.n9020 VSS 0.116823f
C29018 VDD.n9021 VSS 0.78631f
C29019 VDD.n9022 VSS 0.116823f
C29020 VDD.t1797 VSS 0.066856f
C29021 VDD.n9023 VSS 0.14405f
C29022 VDD.n9024 VSS 0.120118f
C29023 VDD.n9025 VSS 0.016021f
C29024 VDD.t2065 VSS 0.025104f
C29025 VDD.n9026 VSS 0.105404f
C29026 VDD.t2192 VSS 0.066856f
C29027 VDD.n9027 VSS 0.14405f
C29028 VDD.t565 VSS 0.025104f
C29029 VDD.t563 VSS 0.066856f
C29030 VDD.n9028 VSS 0.14405f
C29031 VDD.n9029 VSS 0.120118f
C29032 VDD.n9030 VSS 0.016021f
C29033 VDD.t2194 VSS 0.025104f
C29034 VDD.n9031 VSS 0.087217f
C29035 VDD.n9032 VSS 0.057098f
C29036 VDD.n9033 VSS 0.208771f
C29037 VDD.n9034 VSS 0.595476f
C29038 VDD.n9035 VSS 0.645798f
C29039 VDD.n9036 VSS 0.206947f
C29040 VDD.n9037 VSS 0.048151f
C29041 VDD.n9038 VSS 0.083673f
C29042 VDD.t4486 VSS 0.066856f
C29043 VDD.n9039 VSS 0.125227f
C29044 VDD.n9040 VSS 0.101294f
C29045 VDD.n9041 VSS 0.016021f
C29046 VDD.t3025 VSS 0.025104f
C29047 VDD.n9042 VSS 0.099723f
C29048 VDD.n9043 VSS 0.62132f
C29049 VDD.t4473 VSS 0.028519f
C29050 VDD.t4695 VSS 0.028519f
C29051 VDD.n9044 VSS 0.009191f
C29052 VDD.n9045 VSS 0.261039f
C29053 VDD.t4694 VSS 0.066856f
C29054 VDD.t4468 VSS 0.066856f
C29055 VDD.n9046 VSS 0.709674f
C29056 VDD.t2987 VSS 0.028519f
C29057 VDD.t3173 VSS 0.028519f
C29058 VDD.n9047 VSS 0.009191f
C29059 VDD.n9048 VSS 0.644755f
C29060 VDD.t3172 VSS 0.066856f
C29061 VDD.t2982 VSS 0.066856f
C29062 VDD.n9049 VSS 0.690489f
C29063 VDD.t2824 VSS 0.066856f
C29064 VDD.t2609 VSS 0.066856f
C29065 VDD.n9050 VSS 0.690489f
C29066 VDD.t2612 VSS 0.028519f
C29067 VDD.t2825 VSS 0.028519f
C29068 VDD.n9051 VSS 0.009191f
C29069 VDD.n9052 VSS 0.523473f
C29070 VDD.n9053 VSS 0.524869f
C29071 VDD.t3179 VSS 0.028519f
C29072 VDD.t3337 VSS 0.028519f
C29073 VDD.n9054 VSS 0.009191f
C29074 VDD.n9055 VSS 0.471397f
C29075 VDD.t3336 VSS 0.066856f
C29076 VDD.t3176 VSS 0.066856f
C29077 VDD.n9056 VSS 0.690489f
C29078 VDD.t2809 VSS 0.066856f
C29079 VDD.t2587 VSS 0.066856f
C29080 VDD.n9057 VSS 0.690489f
C29081 VDD.t2590 VSS 0.028519f
C29082 VDD.t2810 VSS 0.028519f
C29083 VDD.n9058 VSS 0.009191f
C29084 VDD.n9059 VSS 0.644755f
C29085 VDD.t2449 VSS 0.066856f
C29086 VDD.t2158 VSS 0.066856f
C29087 VDD.n9060 VSS 0.709674f
C29088 VDD.t2165 VSS 0.028519f
C29089 VDD.t2451 VSS 0.028519f
C29090 VDD.n9061 VSS 0.009191f
C29091 VDD.n9062 VSS 0.308318f
C29092 VDD.n9063 VSS 0.766371f
C29093 VDD.n9064 VSS 0.04911f
C29094 VDD.t4772 VSS 0.018805f
C29095 VDD.t4774 VSS 0.019767f
C29096 VDD.n9065 VSS 0.054793f
C29097 VDD.t4775 VSS 0.019781f
C29098 VDD.t4773 VSS 0.018792f
C29099 VDD.n9066 VSS 0.077486f
C29100 VDD.n9067 VSS 0.252514f
C29101 VDD.n9068 VSS 0.199549f
C29102 VDD.n9069 VSS 0.060108f
C29103 VDD.t1894 VSS 0.066856f
C29104 VDD.n9070 VSS 0.131361f
C29105 VDD.n9071 VSS 0.120118f
C29106 VDD.n9072 VSS 0.016021f
C29107 VDD.t2132 VSS 0.025104f
C29108 VDD.n9073 VSS 0.105404f
C29109 VDD.t2304 VSS 0.066856f
C29110 VDD.n9074 VSS 0.14405f
C29111 VDD.t684 VSS 0.025104f
C29112 VDD.t3696 VSS 0.028519f
C29113 VDD.t2147 VSS 0.028519f
C29114 VDD.n9075 VSS 0.009191f
C29115 VDD.t3695 VSS 0.066856f
C29116 VDD.t2256 VSS 0.066856f
C29117 VDD.t4063 VSS 0.028519f
C29118 VDD.t2582 VSS 0.028519f
C29119 VDD.n9076 VSS 0.009191f
C29120 VDD.t4062 VSS 0.066856f
C29121 VDD.t2675 VSS 0.066856f
C29122 VDD.t4656 VSS 0.066856f
C29123 VDD.t3260 VSS 0.066856f
C29124 VDD.t3440 VSS 0.066856f
C29125 VDD.t3166 VSS 0.066856f
C29126 VDD.n9077 VSS 0.690489f
C29127 VDD.t2882 VSS 0.066856f
C29128 VDD.t2581 VSS 0.066856f
C29129 VDD.n9078 VSS 0.690489f
C29130 VDD.t2676 VSS 0.028519f
C29131 VDD.t2883 VSS 0.028519f
C29132 VDD.n9079 VSS 0.009191f
C29133 VDD.n9080 VSS 0.644755f
C29134 VDD.t2538 VSS 0.066856f
C29135 VDD.t2145 VSS 0.066856f
C29136 VDD.n9081 VSS 0.709674f
C29137 VDD.t2258 VSS 0.028519f
C29138 VDD.t2539 VSS 0.028519f
C29139 VDD.n9082 VSS 0.009191f
C29140 VDD.n9083 VSS 0.308318f
C29141 VDD.t3672 VSS 0.066856f
C29142 VDD.n9084 VSS 0.14405f
C29143 VDD.t3899 VSS 0.025104f
C29144 VDD.t4042 VSS 0.066856f
C29145 VDD.n9085 VSS 0.14405f
C29146 VDD.t2549 VSS 0.025104f
C29147 VDD.t2403 VSS 0.028519f
C29148 VDD.t2632 VSS 0.028519f
C29149 VDD.n9086 VSS 0.009191f
C29150 VDD.t2401 VSS 0.066856f
C29151 VDD.t2768 VSS 0.028519f
C29152 VDD.t2979 VSS 0.028519f
C29153 VDD.n9087 VSS 0.009191f
C29154 VDD.t2767 VSS 0.066856f
C29155 VDD.t3134 VSS 0.066856f
C29156 VDD.t3135 VSS 0.028519f
C29157 VDD.t3315 VSS 0.028519f
C29158 VDD.n9088 VSS 0.009191f
C29159 VDD.t4646 VSS 0.066856f
C29160 VDD.t4647 VSS 0.028519f
C29161 VDD.t724 VSS 0.028519f
C29162 VDD.n9089 VSS 0.009191f
C29163 VDD.n9090 VSS 0.035132f
C29164 VDD.t2232 VSS 0.025104f
C29165 VDD.t2090 VSS 0.066856f
C29166 VDD.n9091 VSS 0.125227f
C29167 VDD.t1839 VSS 0.025104f
C29168 VDD.t1838 VSS 0.066856f
C29169 VDD.n9092 VSS 0.125227f
C29170 VDD.n9093 VSS 0.101294f
C29171 VDD.n9094 VSS 0.016021f
C29172 VDD.t2092 VSS 0.025104f
C29173 VDD.n9095 VSS 0.081176f
C29174 VDD.n9096 VSS 0.048151f
C29175 VDD.n9097 VSS 0.083673f
C29176 VDD.t2231 VSS 0.066856f
C29177 VDD.n9098 VSS 0.125227f
C29178 VDD.n9099 VSS 0.006598f
C29179 VDD.n9100 VSS 0.010188f
C29180 VDD.t4756 VSS 0.020387f
C29181 VDD.t4747 VSS 0.022137f
C29182 VDD.n9101 VSS 0.069721f
C29183 VDD.n9102 VSS 0.040089f
C29184 VDD.t4757 VSS 0.022115f
C29185 VDD.t555 VSS 0.020371f
C29186 VDD.n9103 VSS 0.027128f
C29187 VDD.n9104 VSS 0.036577f
C29188 VDD.n9105 VSS 0.044801f
C29189 VDD.n9106 VSS 0.278297f
C29190 VDD.n9107 VSS 0.040089f
C29191 VDD.t4746 VSS 0.020387f
C29192 VDD.n9108 VSS 0.049653f
C29193 VDD.t4790 VSS 0.017093f
C29194 VDD.n9109 VSS 0.042104f
C29195 VDD.n9110 VSS 0.069461f
C29196 VDD.t4791 VSS 0.017093f
C29197 VDD.n9111 VSS 0.035483f
C29198 VDD.t553 VSS 0.020371f
C29199 VDD.n9112 VSS 0.027128f
C29200 VDD.n9113 VSS 0.016538f
C29201 VDD.n9114 VSS 0.027213f
C29202 VDD.n9115 VSS 0.204333f
C29203 VDD.n9116 VSS 0.030906f
C29204 VDD.t625 VSS 0.066856f
C29205 VDD.n9117 VSS 0.045867f
C29206 VDD.n9118 VSS 0.015693f
C29207 VDD.n9119 VSS 0.010881f
C29208 VDD.n9120 VSS 0.044227f
C29209 VDD.n9121 VSS 0.094696f
C29210 VDD.n9122 VSS 0.016021f
C29211 VDD.t627 VSS 0.025104f
C29212 VDD.n9123 VSS 0.108446f
C29213 VDD.n9124 VSS 0.413821f
C29214 VDD.t722 VSS 0.066856f
C29215 VDD.n9125 VSS 0.352487f
C29216 VDD.n9126 VSS 0.320028f
C29217 VDD.t3314 VSS 0.066856f
C29218 VDD.n9127 VSS 0.317129f
C29219 VDD.t2795 VSS 0.066856f
C29220 VDD.t3322 VSS 0.066856f
C29221 VDD.n9128 VSS 0.244224f
C29222 VDD.t3001 VSS 0.025104f
C29223 VDD.n9129 VSS 0.016021f
C29224 VDD.t2796 VSS 0.025104f
C29225 VDD.n9130 VSS 0.139858f
C29226 VDD.t3323 VSS 0.025104f
C29227 VDD.t3519 VSS 0.025104f
C29228 VDD.n9131 VSS 0.016021f
C29229 VDD.n9132 VSS 0.13517f
C29230 VDD.t3000 VSS 0.066856f
C29231 VDD.t3518 VSS 0.066856f
C29232 VDD.n9133 VSS 0.207234f
C29233 VDD.n9134 VSS 0.45584f
C29234 VDD.t2978 VSS 0.066856f
C29235 VDD.n9135 VSS 0.338888f
C29236 VDD.n9136 VSS 0.320028f
C29237 VDD.t2631 VSS 0.066856f
C29238 VDD.n9137 VSS 0.352487f
C29239 VDD.n9138 VSS 0.454091f
C29240 VDD.n9139 VSS 0.203172f
C29241 VDD.t2548 VSS 0.066856f
C29242 VDD.n9140 VSS 0.14405f
C29243 VDD.n9141 VSS 0.120118f
C29244 VDD.n9142 VSS 0.016021f
C29245 VDD.t4043 VSS 0.025104f
C29246 VDD.n9143 VSS 0.087217f
C29247 VDD.n9144 VSS 0.057098f
C29248 VDD.n9145 VSS 0.105404f
C29249 VDD.t3898 VSS 0.066856f
C29250 VDD.n9146 VSS 0.14405f
C29251 VDD.n9147 VSS 0.120118f
C29252 VDD.n9148 VSS 0.016021f
C29253 VDD.t3673 VSS 0.025104f
C29254 VDD.n9149 VSS 0.116823f
C29255 VDD.n9150 VSS 0.779905f
C29256 VDD.n9151 VSS 0.116823f
C29257 VDD.t682 VSS 0.066856f
C29258 VDD.n9152 VSS 0.14405f
C29259 VDD.n9153 VSS 0.120118f
C29260 VDD.n9154 VSS 0.016021f
C29261 VDD.t2306 VSS 0.025104f
C29262 VDD.n9155 VSS 0.087217f
C29263 VDD.n9156 VSS 0.057098f
C29264 VDD.n9157 VSS 0.208771f
C29265 VDD.n9158 VSS 0.595476f
C29266 VDD.n9159 VSS 0.645798f
C29267 VDD.n9160 VSS 0.206947f
C29268 VDD.n9161 VSS 0.048151f
C29269 VDD.n9162 VSS 0.083673f
C29270 VDD.t4568 VSS 0.066856f
C29271 VDD.n9163 VSS 0.125227f
C29272 VDD.n9164 VSS 0.101294f
C29273 VDD.n9165 VSS 0.016021f
C29274 VDD.t3103 VSS 0.025104f
C29275 VDD.n9166 VSS 0.099723f
C29276 VDD.n9167 VSS 0.62132f
C29277 VDD.t4541 VSS 0.028519f
C29278 VDD.t608 VSS 0.028519f
C29279 VDD.n9168 VSS 0.009191f
C29280 VDD.n9169 VSS 0.261039f
C29281 VDD.t606 VSS 0.066856f
C29282 VDD.t4464 VSS 0.066856f
C29283 VDD.n9170 VSS 0.709674f
C29284 VDD.t3055 VSS 0.028519f
C29285 VDD.t3255 VSS 0.028519f
C29286 VDD.n9171 VSS 0.009191f
C29287 VDD.n9172 VSS 0.644755f
C29288 VDD.t3254 VSS 0.066856f
C29289 VDD.t2970 VSS 0.066856f
C29290 VDD.n9173 VSS 0.690489f
C29291 VDD.t2904 VSS 0.066856f
C29292 VDD.t2601 VSS 0.066856f
C29293 VDD.n9174 VSS 0.690489f
C29294 VDD.t2687 VSS 0.028519f
C29295 VDD.t2905 VSS 0.028519f
C29296 VDD.n9175 VSS 0.009191f
C29297 VDD.n9176 VSS 0.523473f
C29298 VDD.n9177 VSS 0.524869f
C29299 VDD.n9178 VSS 0.208534f
C29300 VDD.n9179 VSS 0.865258f
C29301 VDD.t1869 VSS 1.45794f
C29302 VDD.t2146 VSS 1.96535f
C29303 VDD.t554 VSS 1.96535f
C29304 VDD.t2091 VSS 1.36988f
C29305 VDD.n9180 VSS 0.645798f
C29306 VDD.n9181 VSS 0.595476f
C29307 VDD.t552 VSS 1.31955f
C29308 VDD.t626 VSS 1.96535f
C29309 VDD.t2402 VSS 1.96535f
C29310 VDD.t723 VSS 1.45905f
C29311 VDD.n9182 VSS 1.049f
C29312 VDD.n9183 VSS 0.265846f
C29313 VDD.n9184 VSS 0.218139f
C29314 VDD.n9185 VSS 0.064646f
C29315 VDD.n9186 VSS 0.012131f
C29316 VDD.n9187 VSS 0.006065f
C29317 VDD.n9188 VSS 0.012131f
C29318 VDD.n9189 VSS 0.012131f
C29319 VDD.n9190 VSS 0.012131f
C29320 VDD.n9191 VSS 0.012131f
C29321 VDD.n9192 VSS 0.012131f
C29322 VDD.n9193 VSS 0.012131f
C29323 VDD.n9194 VSS 0.012131f
C29324 VDD.n9195 VSS 0.012131f
C29325 VDD.n9196 VSS 0.012131f
C29326 VDD.n9197 VSS 0.012131f
C29327 VDD.n9198 VSS 0.012131f
C29328 VDD.n9199 VSS 0.006065f
C29329 VDD.n9200 VSS 0.012131f
C29330 VDD.n9201 VSS 0.012131f
C29331 VDD.n9202 VSS 0.012131f
C29332 VDD.n9203 VSS 0.012131f
C29333 VDD.n9204 VSS 0.012131f
C29334 VDD.n9205 VSS 0.012131f
C29335 VDD.n9206 VSS 0.012131f
C29336 VDD.n9207 VSS 0.012131f
C29337 VDD.n9208 VSS 0.012131f
C29338 VDD.n9209 VSS 0.012131f
C29339 VDD.n9210 VSS 0.012131f
C29340 VDD.n9211 VSS 0.012131f
C29341 VDD.n9212 VSS 0.012131f
C29342 VDD.n9213 VSS 0.012131f
C29343 VDD.n9214 VSS 0.032509f
C29344 VDD.n9215 VSS 0.012131f
C29345 VDD.n9216 VSS 0.012131f
C29346 VDD.n9217 VSS 0.012131f
C29347 VDD.n9218 VSS 0.012131f
C29348 VDD.n9219 VSS 0.012131f
C29349 VDD.n9220 VSS 0.012131f
C29350 VDD.n9221 VSS 0.012131f
C29351 VDD.n9222 VSS 0.012131f
C29352 VDD.n9223 VSS 0.012131f
C29353 VDD.n9224 VSS 0.012131f
C29354 VDD.n9225 VSS 0.012131f
C29355 VDD.n9226 VSS 0.012131f
C29356 VDD.n9227 VSS 0.012131f
C29357 VDD.n9228 VSS 0.012131f
C29358 VDD.n9229 VSS 0.012131f
C29359 VDD.n9230 VSS 0.012131f
C29360 VDD.n9231 VSS 0.012131f
C29361 VDD.n9232 VSS 0.012131f
C29362 VDD.n9233 VSS 0.012131f
C29363 VDD.n9234 VSS 0.012131f
C29364 VDD.n9235 VSS 0.012131f
C29365 VDD.n9236 VSS 0.012131f
C29366 VDD.n9237 VSS 0.012131f
C29367 VDD.n9238 VSS 0.012131f
C29368 VDD.n9239 VSS 0.012131f
C29369 VDD.n9240 VSS 0.012131f
C29370 VDD.n9241 VSS 0.012131f
C29371 VDD.n9242 VSS 0.012131f
C29372 VDD.n9243 VSS 0.012131f
C29373 VDD.n9244 VSS 0.012131f
C29374 VDD.n9245 VSS 0.012131f
C29375 VDD.n9246 VSS 0.012131f
C29376 VDD.n9247 VSS 0.012131f
C29377 VDD.n9248 VSS 0.012131f
C29378 VDD.n9249 VSS 0.012131f
C29379 VDD.n9250 VSS 0.012131f
C29380 VDD.n9251 VSS 0.012131f
C29381 VDD.n9252 VSS 0.012131f
C29382 VDD.n9253 VSS 0.012131f
C29383 VDD.n9254 VSS 0.012131f
C29384 VDD.n9255 VSS 0.012131f
C29385 VDD.n9256 VSS 0.012131f
C29386 VDD.n9257 VSS 0.012131f
C29387 VDD.n9258 VSS 0.012131f
C29388 VDD.n9259 VSS 0.012131f
C29389 VDD.n9260 VSS 0.012131f
C29390 VDD.n9261 VSS 0.012131f
C29391 VDD.n9262 VSS 0.012131f
C29392 VDD.n9263 VSS 0.012131f
C29393 VDD.n9264 VSS 0.012131f
C29394 VDD.n9265 VSS 0.012131f
C29395 VDD.n9266 VSS 0.012131f
C29396 VDD.n9267 VSS 0.012131f
C29397 VDD.n9268 VSS 0.012131f
C29398 VDD.n9269 VSS 0.012131f
C29399 VDD.n9270 VSS 0.012131f
C29400 VDD.n9271 VSS 0.012131f
C29401 VDD.n9272 VSS 0.012131f
C29402 VDD.n9273 VSS 0.012131f
C29403 VDD.n9274 VSS 0.012131f
C29404 VDD.n9275 VSS 0.012131f
C29405 VDD.n9276 VSS 0.012131f
C29406 VDD.n9277 VSS 0.012131f
C29407 VDD.n9278 VSS 0.012131f
C29408 VDD.n9279 VSS 0.012131f
C29409 VDD.n9280 VSS 0.012131f
C29410 VDD.n9281 VSS 0.012131f
C29411 VDD.n9282 VSS 0.012131f
C29412 VDD.n9283 VSS 0.012131f
C29413 VDD.n9284 VSS 0.012131f
C29414 VDD.n9285 VSS 0.012131f
C29415 VDD.n9286 VSS 0.012131f
C29416 VDD.n9287 VSS 0.012131f
C29417 VDD.n9288 VSS 0.012131f
C29418 VDD.n9289 VSS 0.012131f
C29419 VDD.n9290 VSS 0.012131f
C29420 VDD.n9291 VSS 0.012131f
C29421 VDD.n9292 VSS 0.012131f
C29422 VDD.n9293 VSS 0.012131f
C29423 VDD.n9294 VSS 0.012131f
C29424 VDD.n9295 VSS 0.012131f
C29425 VDD.n9296 VSS 0.012131f
C29426 VDD.n9297 VSS 0.012131f
C29427 VDD.n9298 VSS 0.012131f
C29428 VDD.n9299 VSS 0.012131f
C29429 VDD.n9300 VSS 0.012131f
C29430 VDD.n9301 VSS 0.012131f
C29431 VDD.n9302 VSS 0.012131f
C29432 VDD.n9303 VSS 0.012131f
C29433 VDD.n9304 VSS 0.012131f
C29434 VDD.n9305 VSS 0.012131f
C29435 VDD.n9306 VSS 0.012131f
C29436 VDD.n9307 VSS 0.012131f
C29437 VDD.n9308 VSS 0.012131f
C29438 VDD.n9309 VSS 0.012131f
C29439 VDD.n9310 VSS 0.012131f
C29440 VDD.n9311 VSS 0.012131f
C29441 VDD.n9312 VSS 0.012131f
C29442 VDD.n9313 VSS 0.012131f
C29443 VDD.n9314 VSS 0.012131f
C29444 VDD.n9315 VSS 0.012131f
C29445 VDD.n9316 VSS 0.012131f
C29446 VDD.n9317 VSS 0.012131f
C29447 VDD.n9318 VSS 0.012131f
C29448 VDD.n9319 VSS 0.012131f
C29449 VDD.n9320 VSS 0.012131f
C29450 VDD.n9321 VSS 0.012131f
C29451 VDD.n9322 VSS 0.012131f
C29452 VDD.n9323 VSS 0.012131f
C29453 VDD.n9324 VSS 0.012131f
C29454 VDD.n9325 VSS 0.012131f
C29455 VDD.n9326 VSS 0.012131f
C29456 VDD.n9327 VSS 0.012131f
C29457 VDD.n9328 VSS 0.012131f
C29458 VDD.n9329 VSS 0.012131f
C29459 VDD.n9330 VSS 0.012131f
C29460 VDD.n9331 VSS 0.012131f
C29461 VDD.n9332 VSS 0.012131f
C29462 VDD.n9333 VSS 0.012131f
C29463 VDD.n9334 VSS 0.012131f
C29464 VDD.n9335 VSS 0.012131f
C29465 VDD.n9336 VSS 0.012131f
C29466 VDD.n9337 VSS 0.012131f
C29467 VDD.n9338 VSS 0.012131f
C29468 VDD.n9339 VSS 0.012131f
C29469 VDD.n9340 VSS 0.012131f
C29470 VDD.n9341 VSS 0.012131f
C29471 VDD.n9342 VSS 0.012131f
C29472 VDD.n9343 VSS 0.012131f
C29473 VDD.n9344 VSS 0.012131f
C29474 VDD.n9345 VSS 0.012131f
C29475 VDD.n9346 VSS 0.012131f
C29476 VDD.n9347 VSS 0.012131f
C29477 VDD.n9348 VSS 0.012131f
C29478 VDD.n9349 VSS 0.012131f
C29479 VDD.n9350 VSS 0.012131f
C29480 VDD.n9351 VSS 0.012131f
C29481 VDD.n9352 VSS 0.012131f
C29482 VDD.n9353 VSS 0.012131f
C29483 VDD.n9354 VSS 0.012131f
C29484 VDD.n9355 VSS 0.012131f
C29485 VDD.n9356 VSS 0.012131f
C29486 VDD.n9357 VSS 0.012131f
C29487 VDD.n9358 VSS 0.012131f
C29488 VDD.n9359 VSS 0.012131f
C29489 VDD.n9360 VSS 0.012131f
C29490 VDD.n9361 VSS 0.012131f
C29491 VDD.n9362 VSS 0.012131f
C29492 VDD.n9363 VSS 0.012131f
C29493 VDD.n9364 VSS 0.012131f
C29494 VDD.n9365 VSS 0.012131f
C29495 VDD.n9366 VSS 0.012131f
C29496 VDD.n9367 VSS 0.012131f
C29497 VDD.n9368 VSS 0.012131f
C29498 VDD.n9369 VSS 0.012131f
C29499 VDD.n9370 VSS 0.012131f
C29500 VDD.n9371 VSS 0.012131f
C29501 VDD.n9372 VSS 0.012131f
C29502 VDD.n9373 VSS 0.012131f
C29503 VDD.n9374 VSS 0.012131f
C29504 VDD.n9375 VSS 0.012131f
C29505 VDD.n9376 VSS 0.012131f
C29506 VDD.n9377 VSS 0.012131f
C29507 VDD.n9378 VSS 0.012131f
C29508 VDD.n9379 VSS 0.012131f
C29509 VDD.n9380 VSS 0.012131f
C29510 VDD.n9381 VSS 0.012131f
C29511 VDD.n9382 VSS 0.012131f
C29512 VDD.n9383 VSS 0.012131f
C29513 VDD.n9384 VSS 0.012131f
C29514 VDD.n9385 VSS 0.012131f
C29515 VDD.n9386 VSS 0.012131f
C29516 VDD.n9387 VSS 0.012131f
C29517 VDD.n9388 VSS 0.012131f
C29518 VDD.n9389 VSS 0.012131f
C29519 VDD.n9390 VSS 0.012131f
C29520 VDD.n9391 VSS 0.012131f
C29521 VDD.n9392 VSS 0.012131f
C29522 VDD.n9393 VSS 0.012131f
C29523 VDD.n9394 VSS 0.012131f
C29524 VDD.n9395 VSS 0.012131f
C29525 VDD.n9396 VSS 0.012131f
C29526 VDD.n9397 VSS 0.012131f
C29527 VDD.n9398 VSS 0.012131f
C29528 VDD.n9399 VSS 0.012131f
C29529 VDD.n9400 VSS 0.012131f
C29530 VDD.n9401 VSS 0.012131f
C29531 VDD.n9402 VSS 0.012131f
C29532 VDD.n9403 VSS 0.012131f
C29533 VDD.n9404 VSS 0.012131f
C29534 VDD.n9405 VSS 0.012131f
C29535 VDD.n9406 VSS 0.012131f
C29536 VDD.n9407 VSS 0.012131f
C29537 VDD.n9408 VSS 0.012131f
C29538 VDD.n9409 VSS 0.012131f
C29539 VDD.n9410 VSS 0.012131f
C29540 VDD.n9411 VSS 0.012131f
C29541 VDD.n9412 VSS 0.012131f
C29542 VDD.n9413 VSS 0.012131f
C29543 VDD.n9414 VSS 0.012131f
C29544 VDD.n9415 VSS 0.012131f
C29545 VDD.n9416 VSS 0.012131f
C29546 VDD.n9417 VSS 0.012131f
C29547 VDD.n9418 VSS 0.012131f
C29548 VDD.n9419 VSS 0.012131f
C29549 VDD.n9420 VSS 0.012131f
C29550 VDD.n9421 VSS 0.012131f
C29551 VDD.n9422 VSS 0.012131f
C29552 VDD.n9423 VSS 0.012131f
C29553 VDD.n9424 VSS 0.012131f
C29554 VDD.n9425 VSS 0.012131f
C29555 VDD.n9426 VSS 0.012131f
C29556 VDD.n9427 VSS 0.012131f
C29557 VDD.n9428 VSS 0.012131f
C29558 VDD.n9429 VSS 0.012131f
C29559 VDD.n9430 VSS 0.012131f
C29560 VDD.n9431 VSS 0.012131f
C29561 VDD.n9432 VSS 0.012131f
C29562 VDD.n9433 VSS 0.012131f
C29563 VDD.n9434 VSS 0.012131f
C29564 VDD.n9435 VSS 0.012131f
C29565 VDD.n9436 VSS 0.009956f
C29566 VDD.n9437 VSS 0.012131f
C29567 VDD.n9438 VSS 0.012131f
C29568 VDD.n9439 VSS 0.012131f
C29569 VDD.n9440 VSS 0.012131f
C29570 VDD.n9441 VSS 0.012131f
C29571 VDD.n9442 VSS 0.012131f
C29572 VDD.n9443 VSS 0.012131f
C29573 VDD.n9444 VSS 0.012131f
C29574 VDD.n9445 VSS 0.012131f
C29575 VDD.n9446 VSS 0.012131f
C29576 VDD.n9447 VSS 0.012131f
C29577 VDD.n9448 VSS 0.012131f
C29578 VDD.n9449 VSS 0.012131f
C29579 VDD.n9450 VSS 0.012131f
C29580 VDD.n9451 VSS 0.012131f
C29581 VDD.n9452 VSS 0.012131f
C29582 VDD.n9453 VSS 0.012131f
C29583 VDD.n9454 VSS 0.012131f
C29584 VDD.n9455 VSS 0.012131f
C29585 VDD.n9456 VSS 0.012131f
C29586 VDD.n9457 VSS 0.012131f
C29587 VDD.n9458 VSS 0.012131f
C29588 VDD.n9459 VSS 0.012131f
C29589 VDD.n9460 VSS 0.012131f
C29590 VDD.n9461 VSS 0.012131f
C29591 VDD.n9462 VSS 0.012131f
C29592 VDD.n9463 VSS 0.012131f
C29593 VDD.n9464 VSS 0.012131f
C29594 VDD.n9465 VSS 0.012131f
C29595 VDD.n9466 VSS 0.012131f
C29596 VDD.n9467 VSS 0.012131f
C29597 VDD.n9468 VSS 0.012131f
C29598 VDD.n9469 VSS 0.012131f
C29599 VDD.n9470 VSS 0.012131f
C29600 VDD.n9471 VSS 0.012131f
C29601 VDD.n9472 VSS 0.012131f
C29602 VDD.n9473 VSS 0.012131f
C29603 VDD.n9474 VSS 0.012131f
C29604 VDD.n9475 VSS 0.012131f
C29605 VDD.n9476 VSS 0.012131f
C29606 VDD.n9477 VSS 0.012131f
C29607 VDD.n9478 VSS 0.012131f
C29608 VDD.n9479 VSS 0.012131f
C29609 VDD.n9480 VSS 0.012131f
C29610 VDD.n9481 VSS 0.012131f
C29611 VDD.n9482 VSS 0.012131f
C29612 VDD.n9483 VSS 0.012131f
C29613 VDD.n9484 VSS 0.012131f
C29614 VDD.n9485 VSS 0.012131f
C29615 VDD.n9486 VSS 0.012131f
C29616 VDD.n9487 VSS 0.012131f
C29617 VDD.n9488 VSS 0.012131f
C29618 VDD.n9489 VSS 0.012131f
C29619 VDD.n9490 VSS 0.012131f
C29620 VDD.n9491 VSS 0.012131f
C29621 VDD.n9492 VSS 0.012131f
C29622 VDD.n9493 VSS 0.012131f
C29623 VDD.n9494 VSS 0.012131f
C29624 VDD.n9495 VSS 0.012131f
C29625 VDD.n9496 VSS 0.012131f
C29626 VDD.n9497 VSS 0.012131f
C29627 VDD.n9498 VSS 0.012131f
C29628 VDD.n9499 VSS 0.012131f
C29629 VDD.n9500 VSS 0.012131f
C29630 VDD.n9501 VSS 0.012131f
C29631 VDD.n9502 VSS 0.012131f
C29632 VDD.n9503 VSS 0.012131f
C29633 VDD.n9504 VSS 0.012131f
C29634 VDD.n9505 VSS 0.012131f
C29635 VDD.n9506 VSS 0.012131f
C29636 VDD.n9507 VSS 0.012131f
C29637 VDD.n9508 VSS 0.012131f
C29638 VDD.n9509 VSS 0.012131f
C29639 VDD.n9510 VSS 0.012131f
C29640 VDD.n9511 VSS 0.012131f
C29641 VDD.n9512 VSS 0.012131f
C29642 VDD.n9513 VSS 0.012131f
C29643 VDD.n9514 VSS 0.012131f
C29644 VDD.n9515 VSS 0.012131f
C29645 VDD.n9516 VSS 0.012131f
C29646 VDD.n9517 VSS 0.012131f
C29647 VDD.n9518 VSS 0.012131f
C29648 VDD.n9519 VSS 0.012131f
C29649 VDD.n9520 VSS 0.012131f
C29650 VDD.n9521 VSS 0.012131f
C29651 VDD.n9522 VSS 0.012131f
C29652 VDD.n9523 VSS 0.012131f
C29653 VDD.n9524 VSS 0.012131f
C29654 VDD.n9525 VSS 0.012131f
C29655 VDD.n9526 VSS 0.012131f
C29656 VDD.n9527 VSS 0.012131f
C29657 VDD.n9528 VSS 0.012131f
C29658 VDD.n9529 VSS 0.012131f
C29659 VDD.n9530 VSS 0.012131f
C29660 VDD.n9531 VSS 0.012131f
C29661 VDD.n9532 VSS 0.012131f
C29662 VDD.n9533 VSS 0.012131f
C29663 VDD.n9534 VSS 0.012131f
C29664 VDD.n9535 VSS 0.012131f
C29665 VDD.n9536 VSS 0.012131f
C29666 VDD.n9537 VSS 0.012131f
C29667 VDD.n9538 VSS 0.012131f
C29668 VDD.n9539 VSS 0.012131f
C29669 VDD.n9540 VSS 0.012131f
C29670 VDD.n9541 VSS 0.012131f
C29671 VDD.n9542 VSS 0.012131f
C29672 VDD.n9543 VSS 0.012131f
C29673 VDD.n9544 VSS 0.012131f
C29674 VDD.n9545 VSS 0.012131f
C29675 VDD.n9546 VSS 0.012131f
C29676 VDD.n9547 VSS 0.012131f
C29677 VDD.n9548 VSS 0.012131f
C29678 VDD.n9549 VSS 0.012131f
C29679 VDD.n9550 VSS 0.012131f
C29680 VDD.n9551 VSS 0.012131f
C29681 VDD.n9552 VSS 0.012131f
C29682 VDD.n9553 VSS 0.012131f
C29683 VDD.n9554 VSS 0.012131f
C29684 VDD.n9555 VSS 0.012131f
C29685 VDD.n9556 VSS 0.012131f
C29686 VDD.n9557 VSS 0.012131f
C29687 VDD.n9558 VSS 0.012131f
C29688 VDD.n9559 VSS 0.012131f
C29689 VDD.n9560 VSS 0.012131f
C29690 VDD.n9561 VSS 0.012131f
C29691 VDD.n9562 VSS 0.012131f
C29692 VDD.n9563 VSS 0.012131f
C29693 VDD.n9564 VSS 0.012131f
C29694 VDD.n9565 VSS 0.012131f
C29695 VDD.n9566 VSS 0.012131f
C29696 VDD.n9567 VSS 0.012131f
C29697 VDD.n9568 VSS 0.012131f
C29698 VDD.n9569 VSS 0.012131f
C29699 VDD.n9570 VSS 0.012131f
C29700 VDD.n9571 VSS 0.012131f
C29701 VDD.n9572 VSS 0.012131f
C29702 VDD.n9573 VSS 0.012131f
C29703 VDD.n9574 VSS 0.012131f
C29704 VDD.n9575 VSS 0.012131f
C29705 VDD.n9576 VSS 0.012131f
C29706 VDD.n9577 VSS 0.012131f
C29707 VDD.n9578 VSS 0.012131f
C29708 VDD.n9579 VSS 0.012131f
C29709 VDD.n9580 VSS 0.012131f
C29710 VDD.n9581 VSS 0.012131f
C29711 VDD.n9582 VSS 0.012131f
C29712 VDD.n9583 VSS 0.012131f
C29713 VDD.n9584 VSS 0.012131f
C29714 VDD.n9585 VSS 0.012131f
C29715 VDD.n9586 VSS 0.012131f
C29716 VDD.n9587 VSS 0.012131f
C29717 VDD.n9588 VSS 0.012131f
C29718 VDD.n9589 VSS 0.012131f
C29719 VDD.n9590 VSS 0.012131f
C29720 VDD.n9591 VSS 0.012131f
C29721 VDD.n9592 VSS 0.012131f
C29722 VDD.n9593 VSS 0.012131f
C29723 VDD.n9594 VSS 0.012131f
C29724 VDD.n9595 VSS 0.012131f
C29725 VDD.n9596 VSS 0.012131f
C29726 VDD.n9597 VSS 0.012131f
C29727 VDD.n9598 VSS 0.012131f
C29728 VDD.n9599 VSS 0.012131f
C29729 VDD.n9600 VSS 0.012131f
C29730 VDD.n9601 VSS 0.012131f
C29731 VDD.n9602 VSS 0.012131f
C29732 VDD.n9603 VSS 0.012131f
C29733 VDD.n9604 VSS 0.012131f
C29734 VDD.n9605 VSS 0.012131f
C29735 VDD.n9606 VSS 0.012131f
C29736 VDD.n9607 VSS 0.012131f
C29737 VDD.n9608 VSS 0.012131f
C29738 VDD.n9609 VSS 0.012131f
C29739 VDD.n9610 VSS 0.012131f
C29740 VDD.n9611 VSS 0.012131f
C29741 VDD.n9612 VSS 0.012131f
C29742 VDD.n9613 VSS 0.012131f
C29743 VDD.n9614 VSS 0.012131f
C29744 VDD.n9615 VSS 0.012131f
C29745 VDD.n9616 VSS 0.012131f
C29746 VDD.n9617 VSS 0.012131f
C29747 VDD.n9618 VSS 0.012131f
C29748 VDD.n9619 VSS 0.012131f
C29749 VDD.n9620 VSS 0.012131f
C29750 VDD.n9621 VSS 0.012131f
C29751 VDD.n9622 VSS 0.012131f
C29752 VDD.n9623 VSS 0.012131f
C29753 VDD.n9624 VSS 0.012131f
C29754 VDD.n9625 VSS 0.012131f
C29755 VDD.n9626 VSS 0.012131f
C29756 VDD.n9627 VSS 0.012131f
C29757 VDD.n9628 VSS 0.012131f
C29758 VDD.n9629 VSS 0.012131f
C29759 VDD.n9630 VSS 0.012131f
C29760 VDD.n9631 VSS 0.012131f
C29761 VDD.n9632 VSS 0.012131f
C29762 VDD.n9633 VSS 0.012131f
C29763 VDD.n9634 VSS 0.012131f
C29764 VDD.n9635 VSS 0.012131f
C29765 VDD.n9636 VSS 0.012131f
C29766 VDD.n9637 VSS 0.012131f
C29767 VDD.n9638 VSS 0.012131f
C29768 VDD.n9639 VSS 0.012131f
C29769 VDD.n9640 VSS 0.012131f
C29770 VDD.n9641 VSS 0.012131f
C29771 VDD.n9642 VSS 0.012131f
C29772 VDD.n9643 VSS 0.012131f
C29773 VDD.n9644 VSS 0.012131f
C29774 VDD.n9645 VSS 0.012131f
C29775 VDD.n9646 VSS 0.012131f
C29776 VDD.n9647 VSS 0.012131f
C29777 VDD.n9648 VSS 0.012131f
C29778 VDD.n9649 VSS 0.012131f
C29779 VDD.n9650 VSS 0.012131f
C29780 VDD.n9651 VSS 0.012131f
C29781 VDD.n9652 VSS 0.012131f
C29782 VDD.n9653 VSS 0.012131f
C29783 VDD.n9654 VSS 0.012131f
C29784 VDD.n9655 VSS 0.012131f
C29785 VDD.n9656 VSS 0.012131f
C29786 VDD.n9657 VSS 0.012131f
C29787 VDD.n9658 VSS 0.012131f
C29788 VDD.n9659 VSS 0.012131f
C29789 VDD.n9660 VSS 0.012131f
C29790 VDD.n9661 VSS 0.012131f
C29791 VDD.n9662 VSS 0.012131f
C29792 VDD.n9663 VSS 0.012131f
C29793 VDD.n9664 VSS 0.012131f
C29794 VDD.n9665 VSS 0.012131f
C29795 VDD.n9666 VSS 0.012131f
C29796 VDD.n9667 VSS 0.012131f
C29797 VDD.n9668 VSS 0.012131f
C29798 VDD.n9669 VSS 0.012131f
C29799 VDD.n9670 VSS 0.012131f
C29800 VDD.n9671 VSS 0.012131f
C29801 VDD.n9672 VSS 0.012131f
C29802 VDD.n9673 VSS 0.012131f
C29803 VDD.n9674 VSS 0.012131f
C29804 VDD.n9675 VSS 0.012131f
C29805 VDD.n9676 VSS 0.012131f
C29806 VDD.n9677 VSS 0.012131f
C29807 VDD.n9678 VSS 0.012131f
C29808 VDD.n9679 VSS 0.012131f
C29809 VDD.n9680 VSS 0.012131f
C29810 VDD.n9681 VSS 0.012131f
C29811 VDD.n9682 VSS 0.012131f
C29812 VDD.n9683 VSS 0.012131f
C29813 VDD.n9684 VSS 0.012131f
C29814 VDD.n9685 VSS 0.012131f
C29815 VDD.n9686 VSS 0.012131f
C29816 VDD.n9687 VSS 0.012131f
C29817 VDD.n9688 VSS 0.012131f
C29818 VDD.n9689 VSS 0.012131f
C29819 VDD.n9690 VSS 0.012131f
C29820 VDD.n9691 VSS 0.012131f
C29821 VDD.n9692 VSS 0.012131f
C29822 VDD.n9693 VSS 0.012131f
C29823 VDD.n9694 VSS 0.012131f
C29824 VDD.n9695 VSS 0.012131f
C29825 VDD.n9696 VSS 0.012131f
C29826 VDD.n9697 VSS 0.012131f
C29827 VDD.n9698 VSS 0.012131f
C29828 VDD.n9699 VSS 0.012131f
C29829 VDD.n9700 VSS 0.012131f
C29830 VDD.n9701 VSS 0.012131f
C29831 VDD.n9702 VSS 0.012131f
C29832 VDD.n9703 VSS 0.012131f
C29833 VDD.n9704 VSS 0.012131f
C29834 VDD.n9705 VSS 0.012131f
C29835 VDD.n9706 VSS 0.012131f
C29836 VDD.n9707 VSS 0.012131f
C29837 VDD.n9708 VSS 0.012131f
C29838 VDD.n9709 VSS 0.012131f
C29839 VDD.n9710 VSS 0.012131f
C29840 VDD.n9711 VSS 0.012131f
C29841 VDD.n9712 VSS 0.012131f
C29842 VDD.n9713 VSS 0.012131f
C29843 VDD.n9714 VSS 0.012131f
C29844 VDD.n9715 VSS 0.012131f
C29845 VDD.n9716 VSS 0.012131f
C29846 VDD.n9717 VSS 0.012131f
C29847 VDD.n9718 VSS 0.012131f
C29848 VDD.n9719 VSS 0.012131f
C29849 VDD.n9720 VSS 0.012131f
C29850 VDD.n9721 VSS 0.012131f
C29851 VDD.n9722 VSS 0.012131f
C29852 VDD.n9723 VSS 0.012131f
C29853 VDD.n9724 VSS 0.012131f
C29854 VDD.n9725 VSS 0.012131f
C29855 VDD.n9726 VSS 0.012131f
C29856 VDD.n9727 VSS 0.012131f
C29857 VDD.n9728 VSS 0.012131f
C29858 VDD.n9729 VSS 0.012131f
C29859 VDD.n9730 VSS 0.012131f
C29860 VDD.n9731 VSS 0.012131f
C29861 VDD.n9732 VSS 0.012131f
C29862 VDD.n9733 VSS 0.012131f
C29863 VDD.n9734 VSS 0.012131f
C29864 VDD.n9735 VSS 0.012131f
C29865 VDD.n9736 VSS 0.012131f
C29866 VDD.n9737 VSS 0.012131f
C29867 VDD.n9738 VSS 0.012131f
C29868 VDD.n9739 VSS 0.012131f
C29869 VDD.n9740 VSS 0.012131f
C29870 VDD.n9741 VSS 0.012131f
C29871 VDD.n9742 VSS 0.012131f
C29872 VDD.n9743 VSS 0.012131f
C29873 VDD.n9744 VSS 0.012131f
C29874 VDD.n9745 VSS 0.012131f
C29875 VDD.n9746 VSS 0.012131f
C29876 VDD.n9747 VSS 0.012131f
C29877 VDD.n9748 VSS 0.012131f
C29878 VDD.n9749 VSS 0.012131f
C29879 VDD.n9750 VSS 0.012131f
C29880 VDD.n9751 VSS 0.012131f
C29881 VDD.n9752 VSS 0.012131f
C29882 VDD.n9753 VSS 0.012131f
C29883 VDD.n9754 VSS 0.012131f
C29884 VDD.n9755 VSS 0.012131f
C29885 VDD.n9756 VSS 0.012131f
C29886 VDD.n9757 VSS 0.012131f
C29887 VDD.n9758 VSS 0.012131f
C29888 VDD.n9759 VSS 0.012131f
C29889 VDD.n9760 VSS 0.012131f
C29890 VDD.n9761 VSS 0.012131f
C29891 VDD.n9762 VSS 0.012131f
C29892 VDD.n9763 VSS 0.012131f
C29893 VDD.n9764 VSS 0.012131f
C29894 VDD.n9765 VSS 0.012131f
C29895 VDD.n9766 VSS 0.012131f
C29896 VDD.n9767 VSS 0.012131f
C29897 VDD.n9768 VSS 0.012131f
C29898 VDD.n9769 VSS 0.012131f
C29899 VDD.n9770 VSS 0.012131f
C29900 VDD.n9771 VSS 0.012131f
C29901 VDD.n9772 VSS 0.012131f
C29902 VDD.n9773 VSS 0.012131f
C29903 VDD.n9774 VSS 0.012131f
C29904 VDD.n9775 VSS 0.012131f
C29905 VDD.n9776 VSS 0.012131f
C29906 VDD.n9777 VSS 0.012131f
C29907 VDD.n9778 VSS 0.012131f
C29908 VDD.n9779 VSS 0.012131f
C29909 VDD.n9780 VSS 0.012131f
C29910 VDD.n9781 VSS 0.012131f
C29911 VDD.n9782 VSS 0.012131f
C29912 VDD.n9783 VSS 0.012131f
C29913 VDD.n9784 VSS 0.012131f
C29914 VDD.n9785 VSS 0.012131f
C29915 VDD.n9786 VSS 0.012131f
C29916 VDD.n9787 VSS 0.012131f
C29917 VDD.n9788 VSS 0.012131f
C29918 VDD.n9789 VSS 0.012131f
C29919 VDD.n9790 VSS 0.012131f
C29920 VDD.n9791 VSS 0.012131f
C29921 VDD.n9792 VSS 0.012131f
C29922 VDD.n9793 VSS 0.012131f
C29923 VDD.n9794 VSS 0.012131f
C29924 VDD.n9795 VSS 0.012131f
C29925 VDD.n9796 VSS 0.012131f
C29926 VDD.n9797 VSS 0.012131f
C29927 VDD.n9798 VSS 0.012131f
C29928 VDD.n9799 VSS 0.012131f
C29929 VDD.n9800 VSS 0.012131f
C29930 VDD.n9801 VSS 0.012131f
C29931 VDD.n9802 VSS 0.012131f
C29932 VDD.n9803 VSS 0.012131f
C29933 VDD.n9804 VSS 0.012131f
C29934 VDD.n9805 VSS 0.012131f
C29935 VDD.n9806 VSS 0.012131f
C29936 VDD.n9807 VSS 0.012131f
C29937 VDD.n9808 VSS 0.012131f
C29938 VDD.n9809 VSS 0.012131f
C29939 VDD.n9810 VSS 0.012131f
C29940 VDD.n9811 VSS 0.012131f
C29941 VDD.n9812 VSS 0.012131f
C29942 VDD.n9813 VSS 0.012131f
C29943 VDD.n9814 VSS 0.012131f
C29944 VDD.n9815 VSS 0.012131f
C29945 VDD.n9816 VSS 0.012131f
C29946 VDD.n9817 VSS 0.012131f
C29947 VDD.n9818 VSS 0.012131f
C29948 VDD.n9819 VSS 0.012131f
C29949 VDD.n9820 VSS 0.012131f
C29950 VDD.n9821 VSS 0.012131f
C29951 VDD.n9822 VSS 0.012131f
C29952 VDD.n9823 VSS 0.012131f
C29953 VDD.n9824 VSS 0.012131f
C29954 VDD.n9825 VSS 0.012131f
C29955 VDD.n9826 VSS 0.012131f
C29956 VDD.n9827 VSS 0.012131f
C29957 VDD.n9828 VSS 0.012131f
C29958 VDD.n9829 VSS 0.012131f
C29959 VDD.n9830 VSS 0.012131f
C29960 VDD.n9831 VSS 0.012131f
C29961 VDD.n9832 VSS 0.012131f
C29962 VDD.n9833 VSS 0.012131f
C29963 VDD.n9834 VSS 0.012131f
C29964 VDD.n9835 VSS 0.012131f
C29965 VDD.n9836 VSS 0.012131f
C29966 VDD.n9837 VSS 0.012131f
C29967 VDD.n9838 VSS 0.012131f
C29968 VDD.n9839 VSS 0.012131f
C29969 VDD.n9840 VSS 0.012131f
C29970 VDD.n9841 VSS 0.012131f
C29971 VDD.n9842 VSS 0.012131f
C29972 VDD.n9843 VSS 0.012131f
C29973 VDD.n9844 VSS 0.012131f
C29974 VDD.n9845 VSS 0.012131f
C29975 VDD.n9846 VSS 0.012131f
C29976 VDD.n9847 VSS 0.012131f
C29977 VDD.n9848 VSS 0.012131f
C29978 VDD.n9849 VSS 0.012131f
C29979 VDD.n9850 VSS 0.012131f
C29980 VDD.n9851 VSS 0.012131f
C29981 VDD.n9852 VSS 0.012131f
C29982 VDD.n9853 VSS 0.012131f
C29983 VDD.n9854 VSS 0.012131f
C29984 VDD.n9855 VSS 0.012131f
C29985 VDD.n9856 VSS 0.012131f
C29986 VDD.n9857 VSS 0.012131f
C29987 VDD.n9858 VSS 0.012131f
C29988 VDD.n9859 VSS 0.012131f
C29989 VDD.n9860 VSS 0.012131f
C29990 VDD.n9861 VSS 0.012131f
C29991 VDD.n9862 VSS 0.012131f
C29992 VDD.n9863 VSS 0.012131f
C29993 VDD.n9864 VSS 0.012131f
C29994 VDD.n9865 VSS 0.012131f
C29995 VDD.n9866 VSS 0.012131f
C29996 VDD.n9867 VSS 0.012131f
C29997 VDD.n9868 VSS 0.012131f
C29998 VDD.n9869 VSS 0.012131f
C29999 VDD.n9870 VSS 0.012131f
C30000 VDD.n9871 VSS 0.012131f
C30001 VDD.n9872 VSS 0.012131f
C30002 VDD.n9873 VSS 0.012131f
C30003 VDD.n9874 VSS 0.012131f
C30004 VDD.n9875 VSS 0.012131f
C30005 VDD.n9876 VSS 0.012131f
C30006 VDD.n9877 VSS 0.012131f
C30007 VDD.n9878 VSS 0.012131f
C30008 VDD.n9879 VSS 0.012131f
C30009 VDD.n9880 VSS 0.012131f
C30010 VDD.n9881 VSS 0.012131f
C30011 VDD.n9882 VSS 0.012131f
C30012 VDD.n9883 VSS 0.012131f
C30013 VDD.n9884 VSS 0.012131f
C30014 VDD.n9885 VSS 0.012131f
C30015 VDD.n9886 VSS 0.012131f
C30016 VDD.n9887 VSS 0.012131f
C30017 VDD.n9888 VSS 0.012131f
C30018 VDD.n9889 VSS 0.012131f
C30019 VDD.n9890 VSS 0.012131f
C30020 VDD.n9891 VSS 0.012131f
C30021 VDD.n9892 VSS 0.012131f
C30022 VDD.n9893 VSS 0.012131f
C30023 VDD.n9894 VSS 0.012131f
C30024 VDD.n9895 VSS 0.012131f
C30025 VDD.n9896 VSS 0.012131f
C30026 VDD.n9897 VSS 0.012131f
C30027 VDD.n9898 VSS 0.012131f
C30028 VDD.n9899 VSS 0.012131f
C30029 VDD.n9900 VSS 0.012131f
C30030 VDD.n9901 VSS 0.012131f
C30031 VDD.n9902 VSS 0.012131f
C30032 VDD.n9903 VSS 0.012131f
C30033 VDD.n9904 VSS 0.012131f
C30034 VDD.n9905 VSS 0.012131f
C30035 VDD.n9906 VSS 0.012131f
C30036 VDD.n9907 VSS 0.012131f
C30037 VDD.n9908 VSS 0.012131f
C30038 VDD.n9909 VSS 0.012131f
C30039 VDD.n9910 VSS 0.012131f
C30040 VDD.n9911 VSS 0.012131f
C30041 VDD.n9912 VSS 0.012131f
C30042 VDD.n9913 VSS 0.012131f
C30043 VDD.n9914 VSS 0.012131f
C30044 VDD.n9915 VSS 0.012131f
C30045 VDD.n9916 VSS 0.012131f
C30046 VDD.n9917 VSS 0.012131f
C30047 VDD.n9918 VSS 0.012131f
C30048 VDD.n9919 VSS 0.012131f
C30049 VDD.n9920 VSS 0.012131f
C30050 VDD.n9921 VSS 0.012131f
C30051 VDD.n9922 VSS 0.012131f
C30052 VDD.n9923 VSS 0.012131f
C30053 VDD.n9924 VSS 0.012131f
C30054 VDD.n9925 VSS 0.012131f
C30055 VDD.n9926 VSS 0.012131f
C30056 VDD.n9927 VSS 0.012131f
C30057 VDD.n9928 VSS 0.012131f
C30058 VDD.n9929 VSS 0.012131f
C30059 VDD.n9930 VSS 0.012131f
C30060 VDD.n9931 VSS 0.012131f
C30061 VDD.n9932 VSS 0.012131f
C30062 VDD.n9933 VSS 0.012131f
C30063 VDD.n9934 VSS 0.012131f
C30064 VDD.n9935 VSS 0.012131f
C30065 VDD.n9936 VSS 0.012131f
C30066 VDD.n9937 VSS 0.012131f
C30067 VDD.n9938 VSS 0.012131f
C30068 VDD.n9939 VSS 0.012131f
C30069 VDD.n9940 VSS 0.012131f
C30070 VDD.n9941 VSS 0.012131f
C30071 VDD.n9942 VSS 0.012131f
C30072 VDD.n9943 VSS 0.012131f
C30073 VDD.n9944 VSS 0.012131f
C30074 VDD.n9945 VSS 0.012131f
C30075 VDD.n9946 VSS 0.012131f
C30076 VDD.n9947 VSS 0.012131f
C30077 VDD.n9948 VSS 0.012131f
C30078 VDD.n9949 VSS 0.012131f
C30079 VDD.n9950 VSS 0.012131f
C30080 VDD.n9951 VSS 0.012131f
C30081 VDD.n9952 VSS 0.012131f
C30082 VDD.n9953 VSS 0.012131f
C30083 VDD.n9954 VSS 0.012131f
C30084 VDD.n9955 VSS 0.012131f
C30085 VDD.n9956 VSS 0.012131f
C30086 VDD.n9957 VSS 0.012131f
C30087 VDD.n9958 VSS 0.012131f
C30088 VDD.n9959 VSS 0.012131f
C30089 VDD.n9960 VSS 0.012131f
C30090 VDD.n9961 VSS 0.012131f
C30091 VDD.n9962 VSS 0.012131f
C30092 VDD.n9963 VSS 0.012131f
C30093 VDD.n9964 VSS 0.012131f
C30094 VDD.n9965 VSS 0.012131f
C30095 VDD.n9966 VSS 0.012131f
C30096 VDD.n9967 VSS 0.012131f
C30097 VDD.n9968 VSS 0.012131f
C30098 VDD.n9969 VSS 0.012131f
C30099 VDD.n9970 VSS 0.012131f
C30100 VDD.n9971 VSS 0.012131f
C30101 VDD.n9972 VSS 0.012131f
C30102 VDD.n9973 VSS 0.012131f
C30103 VDD.n9974 VSS 0.012131f
C30104 VDD.n9975 VSS 0.012131f
C30105 VDD.n9976 VSS 0.012131f
C30106 VDD.n9977 VSS 0.012131f
C30107 VDD.n9978 VSS 0.012131f
C30108 VDD.n9979 VSS 0.012131f
C30109 VDD.n9980 VSS 0.012131f
C30110 VDD.n9981 VSS 0.012131f
C30111 VDD.n9982 VSS 0.012131f
C30112 VDD.n9983 VSS 0.012131f
C30113 VDD.n9984 VSS 0.012131f
C30114 VDD.n9985 VSS 0.012131f
C30115 VDD.n9986 VSS 0.012131f
C30116 VDD.n9987 VSS 0.012131f
C30117 VDD.n9988 VSS 0.012131f
C30118 VDD.n9989 VSS 0.012131f
C30119 VDD.n9990 VSS 0.012131f
C30120 VDD.n9991 VSS 0.012131f
C30121 VDD.n9992 VSS 0.012131f
C30122 VDD.n9993 VSS 0.012131f
C30123 VDD.n9994 VSS 0.012131f
C30124 VDD.n9995 VSS 0.012131f
C30125 VDD.n9996 VSS 0.012131f
C30126 VDD.n9997 VSS 0.012131f
C30127 VDD.n9998 VSS 0.012131f
C30128 VDD.n9999 VSS 0.012131f
C30129 VDD.n10000 VSS 0.012131f
C30130 VDD.n10001 VSS 0.012131f
C30131 VDD.n10002 VSS 0.012131f
C30132 VDD.n10003 VSS 0.012131f
C30133 VDD.n10004 VSS 0.012131f
C30134 VDD.n10005 VSS 0.012131f
C30135 VDD.n10006 VSS 0.012131f
C30136 VDD.n10007 VSS 0.012131f
C30137 VDD.n10008 VSS 0.012131f
C30138 VDD.n10009 VSS 0.012131f
C30139 VDD.n10010 VSS 0.012131f
C30140 VDD.n10011 VSS 0.012131f
C30141 VDD.n10012 VSS 0.012131f
C30142 VDD.n10013 VSS 0.012131f
C30143 VDD.n10014 VSS 0.012131f
C30144 VDD.n10015 VSS 0.012131f
C30145 VDD.n10016 VSS 0.012131f
C30146 VDD.n10017 VSS 0.012131f
C30147 VDD.n10018 VSS 0.012131f
C30148 VDD.n10019 VSS 0.012131f
C30149 VDD.n10020 VSS 0.012131f
C30150 VDD.n10021 VSS 0.012131f
C30151 VDD.n10022 VSS 0.012131f
C30152 VDD.n10023 VSS 0.012131f
C30153 VDD.n10024 VSS 0.012131f
C30154 VDD.n10025 VSS 0.012131f
C30155 VDD.n10026 VSS 0.012131f
C30156 VDD.n10027 VSS 0.012131f
C30157 VDD.n10028 VSS 0.012131f
C30158 VDD.n10029 VSS 0.012131f
C30159 VDD.n10030 VSS 0.012131f
C30160 VDD.n10031 VSS 0.012131f
C30161 VDD.n10032 VSS 0.012131f
C30162 VDD.n10033 VSS 0.012131f
C30163 VDD.n10034 VSS 0.012131f
C30164 VDD.n10035 VSS 0.012131f
C30165 VDD.n10036 VSS 0.012131f
C30166 VDD.n10037 VSS 0.012131f
C30167 VDD.n10038 VSS 0.012131f
C30168 VDD.n10039 VSS 0.012131f
C30169 VDD.n10040 VSS 0.012131f
C30170 VDD.n10041 VSS 0.012131f
C30171 VDD.n10042 VSS 0.012131f
C30172 VDD.n10043 VSS 0.012131f
C30173 VDD.n10044 VSS 0.012131f
C30174 VDD.n10045 VSS 0.012131f
C30175 VDD.n10046 VSS 0.012131f
C30176 VDD.n10047 VSS 0.012131f
C30177 VDD.n10048 VSS 0.012131f
C30178 VDD.n10049 VSS 0.012131f
C30179 VDD.n10050 VSS 0.012131f
C30180 VDD.n10051 VSS 0.012131f
C30181 VDD.n10052 VSS 0.012131f
C30182 VDD.n10053 VSS 0.012131f
C30183 VDD.n10054 VSS 0.012131f
C30184 VDD.n10055 VSS 0.012131f
C30185 VDD.n10056 VSS 0.012131f
C30186 VDD.n10057 VSS 0.012131f
C30187 VDD.n10058 VSS 0.012131f
C30188 VDD.n10059 VSS 0.012131f
C30189 VDD.n10060 VSS 0.012131f
C30190 VDD.n10061 VSS 0.012131f
C30191 VDD.n10062 VSS 0.012131f
C30192 VDD.n10063 VSS 0.012131f
C30193 VDD.n10064 VSS 0.012131f
C30194 VDD.n10065 VSS 0.012131f
C30195 VDD.n10066 VSS 0.012131f
C30196 VDD.n10067 VSS 0.012131f
C30197 VDD.n10068 VSS 0.012131f
C30198 VDD.n10069 VSS 0.012131f
C30199 VDD.n10070 VSS 0.012131f
C30200 VDD.n10071 VSS 0.012131f
C30201 VDD.n10072 VSS 0.012131f
C30202 VDD.n10073 VSS 0.012131f
C30203 VDD.n10074 VSS 0.012131f
C30204 VDD.n10075 VSS 0.012131f
C30205 VDD.n10076 VSS 0.012131f
C30206 VDD.n10077 VSS 0.012131f
C30207 VDD.n10078 VSS 0.012131f
C30208 VDD.n10079 VSS 0.012131f
C30209 VDD.n10080 VSS 0.012131f
C30210 VDD.n10081 VSS 0.012131f
C30211 VDD.n10082 VSS 0.012131f
C30212 VDD.n10083 VSS 0.012131f
C30213 VDD.n10084 VSS 0.012131f
C30214 VDD.n10085 VSS 0.012131f
C30215 VDD.n10086 VSS 0.012131f
C30216 VDD.n10087 VSS 0.012131f
C30217 VDD.n10088 VSS 0.012131f
C30218 VDD.n10089 VSS 0.012131f
C30219 VDD.n10090 VSS 0.012131f
C30220 VDD.n10091 VSS 0.012131f
C30221 VDD.n10092 VSS 0.012131f
C30222 VDD.n10093 VSS 0.012131f
C30223 VDD.n10094 VSS 0.012131f
C30224 VDD.n10095 VSS 0.012131f
C30225 VDD.n10096 VSS 0.012131f
C30226 VDD.n10097 VSS 0.012131f
C30227 VDD.n10098 VSS 0.012131f
C30228 VDD.n10099 VSS 0.012131f
C30229 VDD.n10100 VSS 0.012131f
C30230 VDD.n10101 VSS 0.026771f
C30231 VDD.n10102 VSS 0.026771f
C30232 VDD.n10103 VSS 0.032509f
C30233 VDD.n10104 VSS 0.012131f
C30234 VDD.n10105 VSS 0.012131f
C30235 VDD.n10106 VSS 0.012131f
C30236 VDD.n10107 VSS 0.012131f
C30237 VDD.n10108 VSS 0.012131f
C30238 VDD.n10109 VSS 0.012131f
C30239 VDD.n10110 VSS 0.012131f
C30240 VDD.n10111 VSS 0.012131f
C30241 VDD.n10112 VSS 0.012131f
C30242 VDD.n10113 VSS 0.012131f
C30243 VDD.n10114 VSS 0.012131f
C30244 VDD.n10115 VSS 0.012131f
C30245 VDD.n10116 VSS 0.012131f
C30246 VDD.n10117 VSS 0.012131f
C30247 VDD.n10118 VSS 0.012131f
C30248 VDD.n10119 VSS 0.012131f
C30249 VDD.n10120 VSS 0.012131f
C30250 VDD.n10121 VSS 0.012131f
C30251 VDD.n10122 VSS 0.012131f
C30252 VDD.n10123 VSS 0.012131f
C30253 VDD.n10124 VSS 0.012131f
C30254 VDD.n10125 VSS 0.012131f
C30255 VDD.n10126 VSS 0.012131f
C30256 VDD.n10127 VSS 0.012131f
C30257 VDD.n10128 VSS 0.012131f
C30258 VDD.n10129 VSS 0.012131f
C30259 VDD.n10130 VSS 0.012131f
C30260 VDD.n10131 VSS 0.012131f
C30261 VDD.n10132 VSS 0.012131f
C30262 VDD.n10133 VSS 0.012131f
C30263 VDD.n10134 VSS 0.012131f
C30264 VDD.n10135 VSS 0.012131f
C30265 VDD.n10136 VSS 0.012131f
C30266 VDD.n10137 VSS 0.012131f
C30267 VDD.n10138 VSS 0.012131f
C30268 VDD.n10139 VSS 0.012131f
C30269 VDD.n10140 VSS 0.012131f
C30270 VDD.n10141 VSS 0.012131f
C30271 VDD.n10142 VSS 0.012131f
C30272 VDD.n10143 VSS 0.012131f
C30273 VDD.n10144 VSS 0.012131f
C30274 VDD.n10145 VSS 0.012131f
C30275 VDD.n10146 VSS 0.012131f
C30276 VDD.n10147 VSS 0.01173f
C30277 VDD.n10148 VSS 0.044655f
C30278 VDD.n10149 VSS 0.008411f
C30279 VDD.n10150 VSS 0.012131f
C30280 VDD.n10151 VSS 0.012131f
C30281 VDD.n10152 VSS 0.012131f
C30282 VDD.n10153 VSS 0.012131f
C30283 VDD.n10154 VSS 0.012131f
C30284 VDD.n10155 VSS 0.012131f
C30285 VDD.n10156 VSS 0.012131f
C30286 VDD.n10157 VSS 0.012131f
C30287 VDD.n10158 VSS 0.012131f
C30288 VDD.n10159 VSS 0.012131f
C30289 VDD.n10160 VSS 0.012131f
C30290 VDD.n10161 VSS 0.012131f
C30291 VDD.n10162 VSS 0.012131f
C30292 VDD.n10163 VSS 0.012131f
C30293 VDD.n10164 VSS 0.012131f
C30294 VDD.n10165 VSS 0.012131f
C30295 VDD.n10166 VSS 0.012131f
C30296 VDD.n10167 VSS 0.012131f
C30297 VDD.n10168 VSS 0.012131f
C30298 VDD.n10169 VSS 0.012131f
C30299 VDD.n10170 VSS 0.012131f
C30300 VDD.n10171 VSS 0.012131f
C30301 VDD.n10172 VSS 0.012131f
C30302 VDD.n10173 VSS 0.012131f
C30303 VDD.n10174 VSS 0.012131f
C30304 VDD.n10175 VSS 0.012131f
C30305 VDD.n10176 VSS 0.012131f
C30306 VDD.n10177 VSS 0.012131f
C30307 VDD.n10178 VSS 0.012131f
C30308 VDD.n10179 VSS 0.012131f
C30309 VDD.n10180 VSS 0.012131f
C30310 VDD.n10181 VSS 0.012131f
C30311 VDD.n10182 VSS 0.012131f
C30312 VDD.n10183 VSS 0.012131f
C30313 VDD.n10184 VSS 0.012131f
C30314 VDD.n10185 VSS 0.012131f
C30315 VDD.n10186 VSS 0.012131f
C30316 VDD.n10187 VSS 0.012131f
C30317 VDD.n10188 VSS 0.012131f
C30318 VDD.n10189 VSS 0.012131f
C30319 VDD.n10190 VSS 0.012131f
C30320 VDD.n10191 VSS 0.012131f
C30321 VDD.n10192 VSS 0.012131f
C30322 VDD.n10193 VSS 0.012131f
C30323 VDD.n10194 VSS 0.012131f
C30324 VDD.n10195 VSS 0.012131f
C30325 VDD.n10196 VSS 0.012131f
C30326 VDD.n10197 VSS 0.012131f
C30327 VDD.n10198 VSS 0.012131f
C30328 VDD.n10199 VSS 0.012131f
C30329 VDD.n10200 VSS 0.012131f
C30330 VDD.n10201 VSS 0.012131f
C30331 VDD.n10202 VSS 0.012131f
C30332 VDD.n10203 VSS 0.012131f
C30333 VDD.n10204 VSS 0.012131f
C30334 VDD.n10205 VSS 0.012131f
C30335 VDD.n10206 VSS 0.012131f
C30336 VDD.n10207 VSS 0.012131f
C30337 VDD.n10208 VSS 0.012131f
C30338 VDD.n10209 VSS 0.012131f
C30339 VDD.n10210 VSS 0.012131f
C30340 VDD.n10211 VSS 0.012131f
C30341 VDD.n10212 VSS 0.012131f
C30342 VDD.n10213 VSS 0.012131f
C30343 VDD.n10214 VSS 0.012131f
C30344 VDD.n10215 VSS 0.012131f
C30345 VDD.n10216 VSS 0.012131f
C30346 VDD.n10217 VSS 0.012131f
C30347 VDD.n10218 VSS 0.012131f
C30348 VDD.n10219 VSS 0.012131f
C30349 VDD.n10220 VSS 0.012131f
C30350 VDD.n10221 VSS 0.012131f
C30351 VDD.n10222 VSS 0.012131f
C30352 VDD.n10223 VSS 0.012131f
C30353 VDD.n10224 VSS 0.012131f
C30354 VDD.n10225 VSS 0.012131f
C30355 VDD.n10226 VSS 0.012131f
C30356 VDD.n10227 VSS 0.012131f
C30357 VDD.n10228 VSS 0.012131f
C30358 VDD.n10229 VSS 0.012131f
C30359 VDD.n10230 VSS 0.012131f
C30360 VDD.n10231 VSS 0.012131f
C30361 VDD.n10232 VSS 0.012131f
C30362 VDD.n10233 VSS 0.012131f
C30363 VDD.n10234 VSS 0.012131f
C30364 VDD.n10235 VSS 0.012131f
C30365 VDD.n10236 VSS 0.012131f
C30366 VDD.n10237 VSS 0.012131f
C30367 VDD.n10238 VSS 0.012131f
C30368 VDD.n10239 VSS 0.012131f
C30369 VDD.n10240 VSS 0.012131f
C30370 VDD.n10241 VSS 0.012131f
C30371 VDD.n10242 VSS 0.012131f
C30372 VDD.n10243 VSS 0.012131f
C30373 VDD.n10244 VSS 0.012131f
C30374 VDD.n10245 VSS 0.012131f
C30375 VDD.n10246 VSS 0.012131f
C30376 VDD.n10247 VSS 0.012131f
C30377 VDD.n10248 VSS 0.012131f
C30378 VDD.n10249 VSS 0.012131f
C30379 VDD.n10250 VSS 0.012131f
C30380 VDD.n10251 VSS 0.012131f
C30381 VDD.n10252 VSS 0.012131f
C30382 VDD.n10253 VSS 0.012131f
C30383 VDD.n10254 VSS 0.012131f
C30384 VDD.n10255 VSS 0.012131f
C30385 VDD.n10256 VSS 0.012131f
C30386 VDD.n10257 VSS 0.012131f
C30387 VDD.n10258 VSS 0.012131f
C30388 VDD.n10259 VSS 0.012131f
C30389 VDD.n10260 VSS 0.012131f
C30390 VDD.n10261 VSS 0.012131f
C30391 VDD.n10262 VSS 0.012131f
C30392 VDD.n10263 VSS 0.012131f
C30393 VDD.n10264 VSS 0.012131f
C30394 VDD.n10265 VSS 0.012131f
C30395 VDD.n10266 VSS 0.012131f
C30396 VDD.n10267 VSS 0.012131f
C30397 VDD.n10268 VSS 0.012131f
C30398 VDD.n10269 VSS 0.012131f
C30399 VDD.n10270 VSS 0.012131f
C30400 VDD.n10271 VSS 0.012131f
C30401 VDD.n10272 VSS 0.012131f
C30402 VDD.n10273 VSS 0.012131f
C30403 VDD.n10274 VSS 0.012131f
C30404 VDD.n10275 VSS 0.012131f
C30405 VDD.n10276 VSS 0.012131f
C30406 VDD.n10277 VSS 0.012131f
C30407 VDD.n10278 VSS 0.012131f
C30408 VDD.n10279 VSS 0.012131f
C30409 VDD.n10280 VSS 0.012131f
C30410 VDD.n10281 VSS 0.012131f
C30411 VDD.n10282 VSS 0.012131f
C30412 VDD.n10283 VSS 0.012131f
C30413 VDD.n10284 VSS 0.012131f
C30414 VDD.n10285 VSS 0.012131f
C30415 VDD.n10286 VSS 0.012131f
C30416 VDD.n10287 VSS 0.012131f
C30417 VDD.n10288 VSS 0.012131f
C30418 VDD.n10289 VSS 0.012131f
C30419 VDD.n10290 VSS 0.012131f
C30420 VDD.n10291 VSS 0.012131f
C30421 VDD.n10292 VSS 0.012131f
C30422 VDD.n10293 VSS 0.012131f
C30423 VDD.n10294 VSS 0.012131f
C30424 VDD.n10295 VSS 0.012131f
C30425 VDD.n10296 VSS 0.012131f
C30426 VDD.n10297 VSS 0.012131f
C30427 VDD.n10298 VSS 0.012131f
C30428 VDD.n10299 VSS 0.012131f
C30429 VDD.n10300 VSS 0.012131f
C30430 VDD.n10301 VSS 0.012131f
C30431 VDD.n10302 VSS 0.012131f
C30432 VDD.n10303 VSS 0.012131f
C30433 VDD.n10304 VSS 0.012131f
C30434 VDD.n10305 VSS 0.012131f
C30435 VDD.n10306 VSS 0.012131f
C30436 VDD.n10307 VSS 0.012131f
C30437 VDD.n10308 VSS 0.012131f
C30438 VDD.n10309 VSS 0.012131f
C30439 VDD.n10310 VSS 0.012131f
C30440 VDD.n10311 VSS 0.012131f
C30441 VDD.n10312 VSS 0.012131f
C30442 VDD.n10313 VSS 0.012131f
C30443 VDD.n10314 VSS 0.012131f
C30444 VDD.n10315 VSS 0.012131f
C30445 VDD.n10316 VSS 0.012131f
C30446 VDD.n10317 VSS 0.012131f
C30447 VDD.n10318 VSS 0.012131f
C30448 VDD.n10319 VSS 0.012131f
C30449 VDD.n10320 VSS 0.012131f
C30450 VDD.n10321 VSS 0.012131f
C30451 VDD.n10322 VSS 0.012131f
C30452 VDD.n10323 VSS 0.012131f
C30453 VDD.n10324 VSS 0.012131f
C30454 VDD.n10325 VSS 0.012131f
C30455 VDD.n10326 VSS 0.012131f
C30456 VDD.n10327 VSS 0.012131f
C30457 VDD.n10328 VSS 0.012131f
C30458 VDD.n10329 VSS 0.012131f
C30459 VDD.n10330 VSS 0.012131f
C30460 VDD.n10331 VSS 0.012131f
C30461 VDD.n10332 VSS 0.012131f
C30462 VDD.n10333 VSS 0.012131f
C30463 VDD.n10334 VSS 0.012131f
C30464 VDD.n10335 VSS 0.012131f
C30465 VDD.n10336 VSS 0.012131f
C30466 VDD.n10337 VSS 0.012131f
C30467 VDD.n10338 VSS 0.012131f
C30468 VDD.n10339 VSS 0.012131f
C30469 VDD.n10340 VSS 0.012131f
C30470 VDD.n10341 VSS 0.012131f
C30471 VDD.n10342 VSS 0.012131f
C30472 VDD.n10343 VSS 0.012131f
C30473 VDD.n10344 VSS 0.012131f
C30474 VDD.n10345 VSS 0.012131f
C30475 VDD.n10346 VSS 0.012131f
C30476 VDD.n10347 VSS 0.012131f
C30477 VDD.n10348 VSS 0.012131f
C30478 VDD.n10349 VSS 0.012131f
C30479 VDD.n10350 VSS 0.012131f
C30480 VDD.n10351 VSS 0.012131f
C30481 VDD.n10352 VSS 0.012131f
C30482 VDD.n10353 VSS 0.012131f
C30483 VDD.n10354 VSS 0.012131f
C30484 VDD.n10355 VSS 0.012131f
C30485 VDD.n10356 VSS 0.012131f
C30486 VDD.n10357 VSS 0.012131f
C30487 VDD.n10358 VSS 0.012131f
C30488 VDD.n10359 VSS 0.012131f
C30489 VDD.n10360 VSS 0.012131f
C30490 VDD.n10361 VSS 0.012131f
C30491 VDD.n10362 VSS 0.012131f
C30492 VDD.n10363 VSS 0.012131f
C30493 VDD.n10364 VSS 0.012131f
C30494 VDD.n10365 VSS 0.012131f
C30495 VDD.n10366 VSS 0.012131f
C30496 VDD.n10367 VSS 0.012131f
C30497 VDD.n10368 VSS 0.012131f
C30498 VDD.n10369 VSS 0.012131f
C30499 VDD.n10370 VSS 0.012131f
C30500 VDD.n10371 VSS 0.012131f
C30501 VDD.n10372 VSS 0.012131f
C30502 VDD.n10373 VSS 0.012131f
C30503 VDD.n10374 VSS 0.012131f
C30504 VDD.n10375 VSS 0.012131f
C30505 VDD.n10376 VSS 0.012131f
C30506 VDD.n10377 VSS 0.012131f
C30507 VDD.n10378 VSS 0.012131f
C30508 VDD.n10379 VSS 0.012131f
C30509 VDD.n10380 VSS 0.012131f
C30510 VDD.n10381 VSS 0.012131f
C30511 VDD.n10382 VSS 0.012131f
C30512 VDD.n10383 VSS 0.012131f
C30513 VDD.n10384 VSS 0.012131f
C30514 VDD.n10385 VSS 0.012131f
C30515 VDD.n10386 VSS 0.012131f
C30516 VDD.n10387 VSS 0.012131f
C30517 VDD.n10388 VSS 0.012131f
C30518 VDD.n10389 VSS 0.012131f
C30519 VDD.n10390 VSS 0.012131f
C30520 VDD.n10391 VSS 0.012131f
C30521 VDD.n10392 VSS 0.012131f
C30522 VDD.n10393 VSS 0.012131f
C30523 VDD.n10394 VSS 0.012131f
C30524 VDD.n10395 VSS 0.012131f
C30525 VDD.n10396 VSS 0.012131f
C30526 VDD.n10397 VSS 0.012131f
C30527 VDD.n10398 VSS 0.012131f
C30528 VDD.n10399 VSS 0.012131f
C30529 VDD.n10400 VSS 0.012131f
C30530 VDD.n10401 VSS 0.012131f
C30531 VDD.n10402 VSS 0.012131f
C30532 VDD.n10403 VSS 0.012131f
C30533 VDD.n10404 VSS 0.012131f
C30534 VDD.n10405 VSS 0.012131f
C30535 VDD.n10406 VSS 0.012131f
C30536 VDD.n10407 VSS 0.012131f
C30537 VDD.n10408 VSS 0.012131f
C30538 VDD.n10409 VSS 0.012131f
C30539 VDD.n10410 VSS 0.012131f
C30540 VDD.n10411 VSS 0.012131f
C30541 VDD.n10412 VSS 0.012131f
C30542 VDD.n10413 VSS 0.012131f
C30543 VDD.n10414 VSS 0.012131f
C30544 VDD.n10415 VSS 0.012131f
C30545 VDD.n10416 VSS 0.012131f
C30546 VDD.n10417 VSS 0.012131f
C30547 VDD.n10418 VSS 0.012131f
C30548 VDD.n10419 VSS 0.012131f
C30549 VDD.n10420 VSS 0.012131f
C30550 VDD.n10421 VSS 0.012131f
C30551 VDD.n10422 VSS 0.012131f
C30552 VDD.n10423 VSS 0.012131f
C30553 VDD.n10424 VSS 0.012131f
C30554 VDD.n10425 VSS 0.012131f
C30555 VDD.n10426 VSS 0.012131f
C30556 VDD.n10427 VSS 0.012131f
C30557 VDD.n10428 VSS 0.012131f
C30558 VDD.n10429 VSS 0.012131f
C30559 VDD.n10430 VSS 0.012131f
C30560 VDD.n10431 VSS 0.012131f
C30561 VDD.n10432 VSS 0.012131f
C30562 VDD.n10433 VSS 0.012131f
C30563 VDD.n10434 VSS 0.012131f
C30564 VDD.n10435 VSS 0.012131f
C30565 VDD.n10436 VSS 0.012131f
C30566 VDD.n10437 VSS 0.012131f
C30567 VDD.n10438 VSS 0.012131f
C30568 VDD.n10439 VSS 0.012131f
C30569 VDD.n10440 VSS 0.012131f
C30570 VDD.n10441 VSS 0.012131f
C30571 VDD.n10442 VSS 0.012131f
C30572 VDD.n10443 VSS 0.012131f
C30573 VDD.n10444 VSS 0.012131f
C30574 VDD.n10445 VSS 0.012131f
C30575 VDD.n10446 VSS 0.012131f
C30576 VDD.n10447 VSS 0.012131f
C30577 VDD.n10448 VSS 0.012131f
C30578 VDD.n10449 VSS 0.012131f
C30579 VDD.n10450 VSS 0.012131f
C30580 VDD.n10451 VSS 0.012131f
C30581 VDD.n10452 VSS 0.012131f
C30582 VDD.n10453 VSS 0.012131f
C30583 VDD.n10454 VSS 0.012131f
C30584 VDD.n10455 VSS 0.012131f
C30585 VDD.n10456 VSS 0.012131f
C30586 VDD.n10457 VSS 0.012131f
C30587 VDD.n10458 VSS 0.012131f
C30588 VDD.n10459 VSS 0.012131f
C30589 VDD.n10460 VSS 0.012131f
C30590 VDD.n10461 VSS 0.012131f
C30591 VDD.n10462 VSS 0.012131f
C30592 VDD.n10463 VSS 0.012131f
C30593 VDD.n10464 VSS 0.012131f
C30594 VDD.n10465 VSS 0.012131f
C30595 VDD.n10466 VSS 0.012131f
C30596 VDD.n10467 VSS 0.012131f
C30597 VDD.n10468 VSS 0.012131f
C30598 VDD.n10469 VSS 0.012131f
C30599 VDD.n10470 VSS 0.012131f
C30600 VDD.n10471 VSS 0.012131f
C30601 VDD.n10472 VSS 0.012131f
C30602 VDD.n10473 VSS 0.012131f
C30603 VDD.n10474 VSS 0.012131f
C30604 VDD.n10475 VSS 0.012131f
C30605 VDD.n10476 VSS 0.012131f
C30606 VDD.n10477 VSS 0.012131f
C30607 VDD.n10478 VSS 0.012131f
C30608 VDD.n10479 VSS 0.012131f
C30609 VDD.n10480 VSS 0.012131f
C30610 VDD.n10481 VSS 0.012131f
C30611 VDD.n10482 VSS 0.012131f
C30612 VDD.n10483 VSS 0.012131f
C30613 VDD.n10484 VSS 0.012131f
C30614 VDD.n10485 VSS 0.012131f
C30615 VDD.n10486 VSS 0.012131f
C30616 VDD.n10487 VSS 0.012131f
C30617 VDD.n10488 VSS 0.012131f
C30618 VDD.n10489 VSS 0.012131f
C30619 VDD.n10490 VSS 0.012131f
C30620 VDD.n10491 VSS 0.012131f
C30621 VDD.n10492 VSS 0.012131f
C30622 VDD.n10493 VSS 0.012131f
C30623 VDD.n10494 VSS 0.012131f
C30624 VDD.n10495 VSS 0.012131f
C30625 VDD.n10496 VSS 0.012131f
C30626 VDD.n10497 VSS 0.012131f
C30627 VDD.n10498 VSS 0.012131f
C30628 VDD.n10499 VSS 0.012131f
C30629 VDD.n10500 VSS 0.012131f
C30630 VDD.n10501 VSS 0.012131f
C30631 VDD.n10502 VSS 0.012131f
C30632 VDD.n10503 VSS 0.012131f
C30633 VDD.n10504 VSS 0.012131f
C30634 VDD.n10505 VSS 0.012131f
C30635 VDD.n10506 VSS 0.012131f
C30636 VDD.n10507 VSS 0.012131f
C30637 VDD.n10508 VSS 0.012131f
C30638 VDD.n10509 VSS 0.012131f
C30639 VDD.n10510 VSS 0.012131f
C30640 VDD.n10511 VSS 0.012131f
C30641 VDD.n10512 VSS 0.012131f
C30642 VDD.n10513 VSS 0.012131f
C30643 VDD.n10514 VSS 0.012131f
C30644 VDD.n10515 VSS 0.012131f
C30645 VDD.n10516 VSS 0.012131f
C30646 VDD.n10517 VSS 0.012131f
C30647 VDD.n10518 VSS 0.012131f
C30648 VDD.n10519 VSS 0.012131f
C30649 VDD.n10520 VSS 0.012131f
C30650 VDD.n10521 VSS 0.012131f
C30651 VDD.n10522 VSS 0.012131f
C30652 VDD.n10523 VSS 0.012131f
C30653 VDD.n10524 VSS 0.012131f
C30654 VDD.n10525 VSS 0.012131f
C30655 VDD.n10526 VSS 0.012131f
C30656 VDD.n10527 VSS 0.012131f
C30657 VDD.n10528 VSS 0.012131f
C30658 VDD.n10529 VSS 0.012131f
C30659 VDD.n10530 VSS 0.012131f
C30660 VDD.n10531 VSS 0.012131f
C30661 VDD.n10532 VSS 0.012131f
C30662 VDD.n10533 VSS 0.012131f
C30663 VDD.n10534 VSS 0.012131f
C30664 VDD.n10535 VSS 0.012131f
C30665 VDD.n10536 VSS 0.012131f
C30666 VDD.n10537 VSS 0.012131f
C30667 VDD.n10538 VSS 0.012131f
C30668 VDD.n10539 VSS 0.012131f
C30669 VDD.n10540 VSS 0.012131f
C30670 VDD.n10541 VSS 0.012131f
C30671 VDD.n10542 VSS 0.012131f
C30672 VDD.n10543 VSS 0.012131f
C30673 VDD.n10544 VSS 0.012131f
C30674 VDD.n10545 VSS 0.012131f
C30675 VDD.n10546 VSS 0.012131f
C30676 VDD.n10547 VSS 0.012131f
C30677 VDD.n10548 VSS 0.012131f
C30678 VDD.n10549 VSS 0.012131f
C30679 VDD.n10550 VSS 0.012131f
C30680 VDD.n10551 VSS 0.012131f
C30681 VDD.n10552 VSS 0.012131f
C30682 VDD.n10553 VSS 0.012131f
C30683 VDD.n10554 VSS 0.012131f
C30684 VDD.n10555 VSS 0.012131f
C30685 VDD.n10556 VSS 0.012131f
C30686 VDD.n10557 VSS 0.012131f
C30687 VDD.n10558 VSS 0.012131f
C30688 VDD.n10559 VSS 0.012131f
C30689 VDD.n10560 VSS 0.012131f
C30690 VDD.n10561 VSS 0.012131f
C30691 VDD.n10562 VSS 0.012131f
C30692 VDD.n10563 VSS 0.012131f
C30693 VDD.n10564 VSS 0.012131f
C30694 VDD.n10565 VSS 0.012131f
C30695 VDD.n10566 VSS 0.012131f
C30696 VDD.n10567 VSS 0.012131f
C30697 VDD.n10568 VSS 0.012131f
C30698 VDD.n10569 VSS 0.012131f
C30699 VDD.n10570 VSS 0.012131f
C30700 VDD.n10571 VSS 0.012131f
C30701 VDD.n10572 VSS 0.012131f
C30702 VDD.n10573 VSS 0.012131f
C30703 VDD.n10574 VSS 0.012131f
C30704 VDD.n10575 VSS 0.012131f
C30705 VDD.n10576 VSS 0.012131f
C30706 VDD.n10577 VSS 0.012131f
C30707 VDD.n10578 VSS 0.012131f
C30708 VDD.n10579 VSS 0.012131f
C30709 VDD.n10580 VSS 0.012131f
C30710 VDD.n10581 VSS 0.012131f
C30711 VDD.n10582 VSS 0.012131f
C30712 VDD.n10583 VSS 0.012131f
C30713 VDD.n10584 VSS 0.012131f
C30714 VDD.n10585 VSS 0.012131f
C30715 VDD.n10586 VSS 0.012131f
C30716 VDD.n10587 VSS 0.012131f
C30717 VDD.n10588 VSS 0.012131f
C30718 VDD.n10589 VSS 0.012131f
C30719 VDD.n10590 VSS 0.012131f
C30720 VDD.n10591 VSS 0.012131f
C30721 VDD.n10592 VSS 0.012131f
C30722 VDD.n10593 VSS 0.012131f
C30723 VDD.n10594 VSS 0.012131f
C30724 VDD.n10595 VSS 0.012131f
C30725 VDD.n10596 VSS 0.012131f
C30726 VDD.n10597 VSS 0.012131f
C30727 VDD.n10598 VSS 0.012131f
C30728 VDD.n10599 VSS 0.012131f
C30729 VDD.n10600 VSS 0.012131f
C30730 VDD.n10601 VSS 0.012131f
C30731 VDD.n10602 VSS 0.012131f
C30732 VDD.n10603 VSS 0.012131f
C30733 VDD.n10604 VSS 0.012131f
C30734 VDD.n10605 VSS 0.012131f
C30735 VDD.n10606 VSS 0.012131f
C30736 VDD.n10607 VSS 0.012131f
C30737 VDD.n10608 VSS 0.012131f
C30738 VDD.n10609 VSS 0.012131f
C30739 VDD.n10610 VSS 0.012131f
C30740 VDD.n10611 VSS 0.012131f
C30741 VDD.n10612 VSS 0.012131f
C30742 VDD.n10613 VSS 0.012131f
C30743 VDD.n10614 VSS 0.012131f
C30744 VDD.n10615 VSS 0.012131f
C30745 VDD.n10616 VSS 0.012131f
C30746 VDD.n10617 VSS 0.012131f
C30747 VDD.n10618 VSS 0.012131f
C30748 VDD.n10619 VSS 0.012131f
C30749 VDD.n10620 VSS 0.012131f
C30750 VDD.n10621 VSS 0.012131f
C30751 VDD.n10622 VSS 0.012131f
C30752 VDD.n10623 VSS 0.012131f
C30753 VDD.n10624 VSS 0.012131f
C30754 VDD.n10625 VSS 0.012131f
C30755 VDD.n10626 VSS 0.012131f
C30756 VDD.n10627 VSS 0.012131f
C30757 VDD.n10628 VSS 0.012131f
C30758 VDD.n10629 VSS 0.012131f
C30759 VDD.n10630 VSS 0.012131f
C30760 VDD.n10631 VSS 0.012131f
C30761 VDD.n10632 VSS 0.012131f
C30762 VDD.n10633 VSS 0.012131f
C30763 VDD.n10634 VSS 0.012131f
C30764 VDD.n10635 VSS 0.012131f
C30765 VDD.n10636 VSS 0.012131f
C30766 VDD.n10637 VSS 0.012131f
C30767 VDD.n10638 VSS 0.012131f
C30768 VDD.n10639 VSS 0.012131f
C30769 VDD.n10640 VSS 0.012131f
C30770 VDD.n10641 VSS 0.012131f
C30771 VDD.n10642 VSS 0.012131f
C30772 VDD.n10643 VSS 0.012131f
C30773 VDD.n10644 VSS 0.012131f
C30774 VDD.n10645 VSS 0.012131f
C30775 VDD.n10646 VSS 0.012131f
C30776 VDD.n10647 VSS 0.012131f
C30777 VDD.n10648 VSS 0.012131f
C30778 VDD.n10649 VSS 0.012131f
C30779 VDD.n10650 VSS 0.012131f
C30780 VDD.n10651 VSS 0.012131f
C30781 VDD.n10652 VSS 0.012131f
C30782 VDD.n10653 VSS 0.012131f
C30783 VDD.n10654 VSS 0.012131f
C30784 VDD.n10655 VSS 0.012131f
C30785 VDD.n10656 VSS 0.012131f
C30786 VDD.n10657 VSS 0.012131f
C30787 VDD.n10658 VSS 0.012131f
C30788 VDD.n10659 VSS 0.012131f
C30789 VDD.n10660 VSS 0.012131f
C30790 VDD.n10661 VSS 0.012131f
C30791 VDD.n10662 VSS 0.012131f
C30792 VDD.n10663 VSS 0.012131f
C30793 VDD.n10664 VSS 0.012131f
C30794 VDD.n10665 VSS 0.012131f
C30795 VDD.n10666 VSS 0.012131f
C30796 VDD.n10667 VSS 0.012131f
C30797 VDD.n10668 VSS 0.012131f
C30798 VDD.n10669 VSS 0.012131f
C30799 VDD.n10670 VSS 0.012131f
C30800 VDD.n10671 VSS 0.012131f
C30801 VDD.n10672 VSS 0.012131f
C30802 VDD.n10673 VSS 0.012131f
C30803 VDD.n10674 VSS 0.012131f
C30804 VDD.n10675 VSS 0.012131f
C30805 VDD.n10676 VSS 0.012131f
C30806 VDD.n10677 VSS 0.012131f
C30807 VDD.n10678 VSS 0.012131f
C30808 VDD.n10679 VSS 0.012131f
C30809 VDD.n10680 VSS 0.012131f
C30810 VDD.n10681 VSS 0.012131f
C30811 VDD.n10682 VSS 0.012131f
C30812 VDD.n10683 VSS 0.012131f
C30813 VDD.n10684 VSS 0.012131f
C30814 VDD.n10685 VSS 0.012131f
C30815 VDD.n10686 VSS 0.012131f
C30816 VDD.n10687 VSS 0.012131f
C30817 VDD.n10688 VSS 0.012131f
C30818 VDD.n10689 VSS 0.012131f
C30819 VDD.n10690 VSS 0.012131f
C30820 VDD.n10691 VSS 0.012131f
C30821 VDD.n10692 VSS 0.012131f
C30822 VDD.n10693 VSS 0.012131f
C30823 VDD.n10694 VSS 0.012131f
C30824 VDD.n10695 VSS 0.012131f
C30825 VDD.n10696 VSS 0.012131f
C30826 VDD.n10697 VSS 0.012131f
C30827 VDD.n10698 VSS 0.012131f
C30828 VDD.n10699 VSS 0.012131f
C30829 VDD.n10700 VSS 0.012131f
C30830 VDD.n10701 VSS 0.012131f
C30831 VDD.n10702 VSS 0.012131f
C30832 VDD.n10703 VSS 0.012131f
C30833 VDD.n10704 VSS 0.012131f
C30834 VDD.n10705 VSS 0.012131f
C30835 VDD.n10706 VSS 0.012131f
C30836 VDD.n10707 VSS 0.012131f
C30837 VDD.n10708 VSS 0.012131f
C30838 VDD.n10709 VSS 0.012131f
C30839 VDD.n10710 VSS 0.012131f
C30840 VDD.n10711 VSS 0.012131f
C30841 VDD.n10712 VSS 0.012131f
C30842 VDD.n10713 VSS 0.012131f
C30843 VDD.n10714 VSS 0.012131f
C30844 VDD.n10715 VSS 0.012131f
C30845 VDD.n10716 VSS 0.012131f
C30846 VDD.n10717 VSS 0.012131f
C30847 VDD.n10718 VSS 0.012131f
C30848 VDD.n10719 VSS 0.012131f
C30849 VDD.n10720 VSS 0.012131f
C30850 VDD.n10721 VSS 0.012131f
C30851 VDD.n10722 VSS 0.012131f
C30852 VDD.n10723 VSS 0.012131f
C30853 VDD.n10724 VSS 0.012131f
C30854 VDD.n10725 VSS 0.012131f
C30855 VDD.n10726 VSS 0.012131f
C30856 VDD.n10727 VSS 0.012131f
C30857 VDD.n10728 VSS 0.012131f
C30858 VDD.n10729 VSS 0.012131f
C30859 VDD.n10730 VSS 0.012131f
C30860 VDD.n10731 VSS 0.012131f
C30861 VDD.n10732 VSS 0.012131f
C30862 VDD.n10733 VSS 0.012131f
C30863 VDD.n10734 VSS 0.012131f
C30864 VDD.n10735 VSS 0.012131f
C30865 VDD.n10736 VSS 0.012131f
C30866 VDD.n10737 VSS 0.012131f
C30867 VDD.n10738 VSS 0.012131f
C30868 VDD.n10739 VSS 0.012131f
C30869 VDD.n10740 VSS 0.012131f
C30870 VDD.n10741 VSS 0.012131f
C30871 VDD.n10742 VSS 0.012131f
C30872 VDD.n10743 VSS 0.012131f
C30873 VDD.n10744 VSS 0.012131f
C30874 VDD.n10745 VSS 0.012131f
C30875 VDD.n10746 VSS 0.012131f
C30876 VDD.n10747 VSS 0.012131f
C30877 VDD.n10748 VSS 0.012131f
C30878 VDD.n10749 VSS 0.012131f
C30879 VDD.n10750 VSS 0.012131f
C30880 VDD.n10751 VSS 0.012131f
C30881 VDD.n10752 VSS 0.012131f
C30882 VDD.n10753 VSS 0.012131f
C30883 VDD.n10754 VSS 0.012131f
C30884 VDD.n10755 VSS 0.012131f
C30885 VDD.n10756 VSS 0.012131f
C30886 VDD.n10757 VSS 0.012131f
C30887 VDD.n10758 VSS 0.012131f
C30888 VDD.n10759 VSS 0.044701f
C30889 VDD.n10760 VSS 0.118213f
C30890 VDD.n10761 VSS 0.106951f
C30891 VDD.n10762 VSS 0.012131f
C30892 VDD.n10763 VSS 0.012131f
C30893 VDD.n10764 VSS 0.012131f
C30894 VDD.n10765 VSS 0.065079f
C30895 VDD.n10766 VSS 0.102538f
C30896 VDD.n10767 VSS 0.116823f
C30897 VDD.t4616 VSS 0.066856f
C30898 VDD.n10768 VSS 0.14405f
C30899 VDD.n10769 VSS 0.120118f
C30900 VDD.n10770 VSS 0.016021f
C30901 VDD.t673 VSS 0.025104f
C30902 VDD.n10771 VSS 0.087217f
C30903 VDD.n10772 VSS 0.057098f
C30904 VDD.t602 VSS 1.45794f
C30905 VDD.t2352 VSS 1.96535f
C30906 VDD.t12 VSS 1.96535f
C30907 VDD.t304 VSS 1.36988f
C30908 VDD.n10773 VSS 0.645798f
C30909 VDD.t758 VSS 1.45905f
C30910 VDD.t1352 VSS 1.96535f
C30911 VDD.t351 VSS 1.96535f
C30912 VDD.t13 VSS 1.31955f
C30913 VDD.n10774 VSS 0.595476f
C30914 VDD.n10775 VSS 0.208771f
C30915 VDD.n10776 VSS 0.208534f
C30916 VDD.n10777 VSS 0.524869f
C30917 VDD.n10778 VSS 0.207221f
C30918 VDD.n10779 VSS 0.865258f
C30919 VDD.t933 VSS 1.45794f
C30920 VDD.t680 VSS 1.96535f
C30921 VDD.t3424 VSS 1.96535f
C30922 VDD.t3614 VSS 1.31955f
C30923 VDD.n10780 VSS 0.595476f
C30924 VDD.n10781 VSS 0.645798f
C30925 VDD.t1713 VSS 1.36988f
C30926 VDD.t1497 VSS 1.96535f
C30927 VDD.t1180 VSS 1.96535f
C30928 VDD.t1325 VSS 1.45794f
C30929 VDD.n10782 VSS 0.865258f
C30930 VDD.n10783 VSS 0.208534f
C30931 VDD.n10784 VSS 0.524869f
C30932 VDD.t3029 VSS 0.028519f
C30933 VDD.t1545 VSS 0.028519f
C30934 VDD.n10785 VSS 0.009191f
C30935 VDD.t2909 VSS 0.028519f
C30936 VDD.t1425 VSS 0.028519f
C30937 VDD.n10786 VSS 0.009191f
C30938 VDD.n10787 VSS 0.471397f
C30939 VDD.t3028 VSS 0.066856f
C30940 VDD.t2908 VSS 0.066856f
C30941 VDD.t1424 VSS 0.066856f
C30942 VDD.t1544 VSS 0.066856f
C30943 VDD.n10788 VSS 0.690489f
C30944 VDD.t2663 VSS 0.066856f
C30945 VDD.t2540 VSS 0.066856f
C30946 VDD.t1083 VSS 0.066856f
C30947 VDD.t1179 VSS 0.066856f
C30948 VDD.n10789 VSS 0.690489f
C30949 VDD.t2664 VSS 0.028519f
C30950 VDD.t1181 VSS 0.028519f
C30951 VDD.n10790 VSS 0.009191f
C30952 VDD.t2541 VSS 0.028519f
C30953 VDD.t1085 VSS 0.028519f
C30954 VDD.n10791 VSS 0.009191f
C30955 VDD.n10792 VSS 0.644755f
C30956 VDD.t1927 VSS 0.066856f
C30957 VDD.t1415 VSS 0.066856f
C30958 VDD.t2743 VSS 0.066856f
C30959 VDD.t3204 VSS 0.066856f
C30960 VDD.n10793 VSS 0.709674f
C30961 VDD.t1928 VSS 0.028519f
C30962 VDD.t3205 VSS 0.028519f
C30963 VDD.n10794 VSS 0.009191f
C30964 VDD.t1416 VSS 0.028519f
C30965 VDD.t2744 VSS 0.028519f
C30966 VDD.n10795 VSS 0.009191f
C30967 VDD.n10796 VSS 0.309003f
C30968 VDD.n10797 VSS 0.765686f
C30969 VDD.n10798 VSS 0.116823f
C30970 VDD.t2741 VSS 0.066856f
C30971 VDD.n10799 VSS 0.14405f
C30972 VDD.n10800 VSS 0.120118f
C30973 VDD.n10801 VSS 0.016021f
C30974 VDD.t2939 VSS 0.025104f
C30975 VDD.n10802 VSS 0.087217f
C30976 VDD.n10803 VSS 0.057098f
C30977 VDD.n10804 VSS 0.105404f
C30978 VDD.t1003 VSS 0.066856f
C30979 VDD.n10805 VSS 0.14405f
C30980 VDD.n10806 VSS 0.120118f
C30981 VDD.n10807 VSS 0.016021f
C30982 VDD.t3939 VSS 0.025104f
C30983 VDD.n10808 VSS 0.116823f
C30984 VDD.t4436 VSS 0.066856f
C30985 VDD.n10809 VSS 0.14405f
C30986 VDD.t3291 VSS 0.025104f
C30987 VDD.n10810 VSS 0.087217f
C30988 VDD.t3290 VSS 0.066856f
C30989 VDD.n10811 VSS 0.14405f
C30990 VDD.n10812 VSS 0.120118f
C30991 VDD.n10813 VSS 0.016021f
C30992 VDD.t4437 VSS 0.025104f
C30993 VDD.n10814 VSS 0.116823f
C30994 VDD.n10815 VSS 0.174205f
C30995 VDD.n10817 VSS 0.604497f
C30996 VDD.n10819 VSS 0.01487f
C30997 VDD.n10820 VSS 0.20611f
C30998 VDD.t1956 VSS 0.066856f
C30999 VDD.t2471 VSS 0.066856f
C31000 VDD.n10821 VSS 0.646278f
C31001 VDD.t4075 VSS 0.028519f
C31002 VDD.t2794 VSS 0.028519f
C31003 VDD.n10822 VSS 0.009191f
C31004 VDD.n10823 VSS 0.650522f
C31005 VDD.t2793 VSS 0.066856f
C31006 VDD.t1715 VSS 0.066856f
C31007 VDD.n10824 VSS 0.696076f
C31008 VDD.t3132 VSS 0.066856f
C31009 VDD.t2117 VSS 0.066856f
C31010 VDD.n10825 VSS 0.696076f
C31011 VDD.t4431 VSS 0.028519f
C31012 VDD.t3133 VSS 0.028519f
C31013 VDD.n10826 VSS 0.009191f
C31014 VDD.n10827 VSS 0.475536f
C31015 VDD.n10828 VSS 0.529799f
C31016 VDD.n10829 VSS 0.208534f
C31017 VDD.n10830 VSS 0.902999f
C31018 VDD.n10831 VSS 0.902999f
C31019 VDD.t1442 VSS 1.45794f
C31020 VDD.t652 VSS 1.96535f
C31021 VDD.t497 VSS 1.96535f
C31022 VDD.t512 VSS 1.31955f
C31023 VDD.n10832 VSS 0.595476f
C31024 VDD.n10833 VSS 0.208771f
C31025 VDD.n10834 VSS 0.208534f
C31026 VDD.n10835 VSS 0.524869f
C31027 VDD.n10836 VSS 0.207221f
C31028 VDD.n10837 VSS 0.865258f
C31029 VDD.t1183 VSS 1.45794f
C31030 VDD.t1373 VSS 1.96535f
C31031 VDD.t3679 VSS 1.96535f
C31032 VDD.t1408 VSS 1.31955f
C31033 VDD.n10838 VSS 0.595476f
C31034 VDD.n10839 VSS 0.645798f
C31035 VDD.t2923 VSS 1.36988f
C31036 VDD.t3748 VSS 1.96535f
C31037 VDD.t958 VSS 1.96535f
C31038 VDD.t816 VSS 1.45794f
C31039 VDD.n10840 VSS 0.865258f
C31040 VDD.n10841 VSS 0.208534f
C31041 VDD.n10842 VSS 0.524869f
C31042 VDD.t4577 VSS 0.028519f
C31043 VDD.t4273 VSS 0.028519f
C31044 VDD.n10843 VSS 0.009191f
C31045 VDD.t4101 VSS 0.028519f
C31046 VDD.t1745 VSS 0.028519f
C31047 VDD.n10844 VSS 0.009191f
C31048 VDD.n10845 VSS 0.471397f
C31049 VDD.t4576 VSS 0.066856f
C31050 VDD.t4100 VSS 0.066856f
C31051 VDD.t1744 VSS 0.066856f
C31052 VDD.t4272 VSS 0.066856f
C31053 VDD.n10846 VSS 0.690489f
C31054 VDD.t4240 VSS 0.066856f
C31055 VDD.t3709 VSS 0.066856f
C31056 VDD.t1375 VSS 0.066856f
C31057 VDD.t3896 VSS 0.066856f
C31058 VDD.n10847 VSS 0.690489f
C31059 VDD.t4241 VSS 0.028519f
C31060 VDD.t3897 VSS 0.028519f
C31061 VDD.n10848 VSS 0.009191f
C31062 VDD.t3710 VSS 0.028519f
C31063 VDD.t1377 VSS 0.028519f
C31064 VDD.n10849 VSS 0.009191f
C31065 VDD.n10850 VSS 0.644755f
C31066 VDD.t815 VSS 0.066856f
C31067 VDD.t3320 VSS 0.066856f
C31068 VDD.t4144 VSS 0.066856f
C31069 VDD.t957 VSS 0.066856f
C31070 VDD.n10851 VSS 0.709674f
C31071 VDD.t817 VSS 0.028519f
C31072 VDD.t959 VSS 0.028519f
C31073 VDD.n10852 VSS 0.009191f
C31074 VDD.t3321 VSS 0.028519f
C31075 VDD.t4145 VSS 0.028519f
C31076 VDD.n10853 VSS 0.009191f
C31077 VDD.n10854 VSS 0.309003f
C31078 VDD.n10855 VSS 0.765686f
C31079 VDD.n10856 VSS 0.116823f
C31080 VDD.t2544 VSS 0.066856f
C31081 VDD.n10857 VSS 0.14405f
C31082 VDD.n10858 VSS 0.120118f
C31083 VDD.n10859 VSS 0.016021f
C31084 VDD.t668 VSS 0.025104f
C31085 VDD.n10860 VSS 0.087217f
C31086 VDD.n10861 VSS 0.057098f
C31087 VDD.n10862 VSS 0.105404f
C31088 VDD.t3014 VSS 0.066856f
C31089 VDD.n10863 VSS 0.14405f
C31090 VDD.n10864 VSS 0.120118f
C31091 VDD.n10865 VSS 0.016021f
C31092 VDD.t2098 VSS 0.025104f
C31093 VDD.n10866 VSS 0.116823f
C31094 VDD.t2263 VSS 0.066856f
C31095 VDD.n10867 VSS 0.14405f
C31096 VDD.t4165 VSS 0.025104f
C31097 VDD.n10868 VSS 0.087217f
C31098 VDD.t4164 VSS 0.066856f
C31099 VDD.n10869 VSS 0.14405f
C31100 VDD.n10870 VSS 0.120118f
C31101 VDD.n10871 VSS 0.016021f
C31102 VDD.t2265 VSS 0.025104f
C31103 VDD.n10872 VSS 0.116823f
C31104 VDD.n10873 VSS 0.785619f
C31105 VDD.t4169 VSS 0.028519f
C31106 VDD.t3913 VSS 0.028519f
C31107 VDD.n10874 VSS 0.009191f
C31108 VDD.n10875 VSS 0.311617f
C31109 VDD.t3912 VSS 0.066856f
C31110 VDD.t4332 VSS 0.066856f
C31111 VDD.n10876 VSS 0.715442f
C31112 VDD.t2598 VSS 0.028519f
C31113 VDD.t1213 VSS 0.028519f
C31114 VDD.n10877 VSS 0.009191f
C31115 VDD.n10878 VSS 0.650522f
C31116 VDD.t1211 VSS 0.066856f
C31117 VDD.t4412 VSS 0.066856f
C31118 VDD.n10879 VSS 0.696076f
C31119 VDD.t1590 VSS 0.066856f
C31120 VDD.t641 VSS 0.066856f
C31121 VDD.n10880 VSS 0.696076f
C31122 VDD.t2967 VSS 0.028519f
C31123 VDD.t1591 VSS 0.028519f
C31124 VDD.n10881 VSS 0.009191f
C31125 VDD.n10882 VSS 0.475536f
C31126 VDD.n10883 VSS 0.529799f
C31127 VDD.n10884 VSS 0.208534f
C31128 VDD.n10885 VSS 0.902999f
C31129 VDD.n10886 VSS 0.902999f
C31130 VDD.t1212 VSS 1.45794f
C31131 VDD.t1265 VSS 1.96535f
C31132 VDD.t2264 VSS 1.96535f
C31133 VDD.t1341 VSS 1.31955f
C31134 VDD.n10887 VSS 0.595476f
C31135 VDD.n10888 VSS 0.208771f
C31136 VDD.n10889 VSS 0.208534f
C31137 VDD.n10890 VSS 0.075373f
C31138 VDD.n10891 VSS 0.207221f
C31139 VDD.n10892 VSS 0.865258f
C31140 VDD.t1959 VSS 1.45794f
C31141 VDD.t1801 VSS 1.96535f
C31142 VDD.t488 VSS 1.96535f
C31143 VDD.t489 VSS 1.31955f
C31144 VDD.n10893 VSS 0.595476f
C31145 VDD.n10894 VSS 0.645798f
C31146 VDD.t491 VSS 1.36988f
C31147 VDD.t490 VSS 1.96535f
C31148 VDD.t1368 VSS 1.96535f
C31149 VDD.t2572 VSS 1.45794f
C31150 VDD.n10895 VSS 0.865258f
C31151 VDD.n10896 VSS 0.208534f
C31152 VDD.n10897 VSS 0.524869f
C31153 VDD.t4099 VSS 0.028519f
C31154 VDD.t1739 VSS 0.028519f
C31155 VDD.n10898 VSS 0.009191f
C31156 VDD.t1558 VSS 0.028519f
C31157 VDD.t1232 VSS 0.028519f
C31158 VDD.n10899 VSS 0.009191f
C31159 VDD.n10900 VSS 0.471397f
C31160 VDD.t4098 VSS 0.066856f
C31161 VDD.t1557 VSS 0.066856f
C31162 VDD.t1231 VSS 0.066856f
C31163 VDD.t1738 VSS 0.066856f
C31164 VDD.n10901 VSS 0.690489f
C31165 VDD.t3703 VSS 0.066856f
C31166 VDD.t1185 VSS 0.066856f
C31167 VDD.t907 VSS 0.066856f
C31168 VDD.t1367 VSS 0.066856f
C31169 VDD.n10902 VSS 0.690489f
C31170 VDD.t3704 VSS 0.028519f
C31171 VDD.t1369 VSS 0.028519f
C31172 VDD.n10903 VSS 0.009191f
C31173 VDD.t1187 VSS 0.028519f
C31174 VDD.t909 VSS 0.028519f
C31175 VDD.n10904 VSS 0.009191f
C31176 VDD.n10905 VSS 0.644755f
C31177 VDD.t3182 VSS 0.066856f
C31178 VDD.t2176 VSS 0.066856f
C31179 VDD.t2358 VSS 0.066856f
C31180 VDD.t3976 VSS 0.066856f
C31181 VDD.n10906 VSS 0.709674f
C31182 VDD.t3183 VSS 0.028519f
C31183 VDD.t3977 VSS 0.028519f
C31184 VDD.n10907 VSS 0.009191f
C31185 VDD.t2177 VSS 0.028519f
C31186 VDD.t2359 VSS 0.028519f
C31187 VDD.n10908 VSS 0.009191f
C31188 VDD.n10909 VSS 0.309003f
C31189 VDD.n10910 VSS 0.765686f
C31190 VDD.n10911 VSS 0.116823f
C31191 VDD.t3369 VSS 0.066856f
C31192 VDD.n10912 VSS 0.14405f
C31193 VDD.n10913 VSS 0.120118f
C31194 VDD.n10914 VSS 0.016021f
C31195 VDD.t3572 VSS 0.025104f
C31196 VDD.n10915 VSS 0.087217f
C31197 VDD.n10916 VSS 0.057098f
C31198 VDD.n10917 VSS 0.105404f
C31199 VDD.t574 VSS 0.066856f
C31200 VDD.n10918 VSS 0.14405f
C31201 VDD.n10919 VSS 0.120118f
C31202 VDD.n10920 VSS 0.016021f
C31203 VDD.t3569 VSS 0.025104f
C31204 VDD.n10921 VSS 0.116823f
C31205 VDD.t3200 VSS 0.066856f
C31206 VDD.n10922 VSS 0.14405f
C31207 VDD.t3356 VSS 0.025104f
C31208 VDD.n10923 VSS 0.087217f
C31209 VDD.t3354 VSS 0.066856f
C31210 VDD.n10924 VSS 0.14405f
C31211 VDD.n10925 VSS 0.120118f
C31212 VDD.n10926 VSS 0.016021f
C31213 VDD.t3201 VSS 0.025104f
C31214 VDD.n10927 VSS 0.116823f
C31215 VDD.n10928 VSS 0.785619f
C31216 VDD.t1926 VSS 0.028519f
C31217 VDD.t3203 VSS 0.028519f
C31218 VDD.n10929 VSS 0.009191f
C31219 VDD.n10930 VSS 0.311617f
C31220 VDD.t3202 VSS 0.066856f
C31221 VDD.t2178 VSS 0.066856f
C31222 VDD.n10931 VSS 0.715442f
C31223 VDD.t1053 VSS 0.028519f
C31224 VDD.t3831 VSS 0.028519f
C31225 VDD.n10932 VSS 0.009191f
C31226 VDD.n10933 VSS 0.650522f
C31227 VDD.t3830 VSS 0.066856f
C31228 VDD.t3340 VSS 0.066856f
C31229 VDD.n10934 VSS 0.696076f
C31230 VDD.t4224 VSS 0.066856f
C31231 VDD.t3717 VSS 0.066856f
C31232 VDD.n10935 VSS 0.696076f
C31233 VDD.t1402 VSS 0.028519f
C31234 VDD.t4225 VSS 0.028519f
C31235 VDD.n10936 VSS 0.009191f
C31236 VDD.n10937 VSS 0.475536f
C31237 VDD.n10938 VSS 0.529799f
C31238 VDD.n10939 VSS 0.208534f
C31239 VDD.n10940 VSS 0.902999f
C31240 VDD.n10941 VSS 0.902999f
C31241 VDD.t2682 VSS 1.45794f
C31242 VDD.t1052 VSS 1.96535f
C31243 VDD.t2776 VSS 1.96535f
C31244 VDD.t3355 VSS 1.31955f
C31245 VDD.n10942 VSS 0.595476f
C31246 VDD.n10943 VSS 0.208771f
C31247 VDD.n10944 VSS 0.208534f
C31248 VDD.n10945 VSS 0.524869f
C31249 VDD.n10946 VSS 0.207221f
C31250 VDD.n10947 VSS 0.865258f
C31251 VDD.t783 VSS 1.45794f
C31252 VDD.t700 VSS 1.96535f
C31253 VDD.t556 VSS 1.96535f
C31254 VDD.t558 VSS 1.31955f
C31255 VDD.n10948 VSS 0.595476f
C31256 VDD.n10949 VSS 0.645798f
C31257 VDD.t559 VSS 1.36988f
C31258 VDD.t557 VSS 1.96535f
C31259 VDD.t896 VSS 1.96535f
C31260 VDD.t938 VSS 1.45794f
C31261 VDD.n10950 VSS 0.865258f
C31262 VDD.n10951 VSS 0.208534f
C31263 VDD.n10952 VSS 0.524869f
C31264 VDD.t2707 VSS 0.028519f
C31265 VDD.t1230 VSS 0.028519f
C31266 VDD.n10953 VSS 0.009191f
C31267 VDD.t4281 VSS 0.028519f
C31268 VDD.t2993 VSS 0.028519f
C31269 VDD.n10954 VSS 0.009191f
C31270 VDD.n10955 VSS 0.471397f
C31271 VDD.t2706 VSS 0.066856f
C31272 VDD.t4280 VSS 0.066856f
C31273 VDD.t2992 VSS 0.066856f
C31274 VDD.t1229 VSS 0.066856f
C31275 VDD.n10956 VSS 0.690489f
C31276 VDD.t2282 VSS 0.066856f
C31277 VDD.t3910 VSS 0.066856f
C31278 VDD.t2619 VSS 0.066856f
C31279 VDD.t895 VSS 0.066856f
C31280 VDD.n10957 VSS 0.690489f
C31281 VDD.t2283 VSS 0.028519f
C31282 VDD.t897 VSS 0.028519f
C31283 VDD.n10958 VSS 0.009191f
C31284 VDD.t3911 VSS 0.028519f
C31285 VDD.t2620 VSS 0.028519f
C31286 VDD.n10959 VSS 0.009191f
C31287 VDD.n10960 VSS 0.644755f
C31288 VDD.t937 VSS 0.066856f
C31289 VDD.t4126 VSS 0.066856f
C31290 VDD.t1144 VSS 0.066856f
C31291 VDD.t2126 VSS 0.066856f
C31292 VDD.n10961 VSS 0.709674f
C31293 VDD.t939 VSS 0.028519f
C31294 VDD.t2127 VSS 0.028519f
C31295 VDD.n10962 VSS 0.009191f
C31296 VDD.t4127 VSS 0.028519f
C31297 VDD.t1146 VSS 0.028519f
C31298 VDD.n10963 VSS 0.009191f
C31299 VDD.n10964 VSS 0.309003f
C31300 VDD.n10965 VSS 0.765686f
C31301 VDD.n10966 VSS 0.116823f
C31302 VDD.t1138 VSS 0.066856f
C31303 VDD.n10967 VSS 0.14405f
C31304 VDD.n10968 VSS 0.120118f
C31305 VDD.n10969 VSS 0.016021f
C31306 VDD.t1332 VSS 0.025104f
C31307 VDD.n10970 VSS 0.087217f
C31308 VDD.n10971 VSS 0.057098f
C31309 VDD.n10972 VSS 0.105404f
C31310 VDD.t3628 VSS 0.066856f
C31311 VDD.n10973 VSS 0.14405f
C31312 VDD.n10974 VSS 0.120118f
C31313 VDD.n10975 VSS 0.016021f
C31314 VDD.t2521 VSS 0.025104f
C31315 VDD.n10976 VSS 0.116823f
C31316 VDD.t1503 VSS 0.066856f
C31317 VDD.n10977 VSS 0.14405f
C31318 VDD.t1388 VSS 0.025104f
C31319 VDD.n10978 VSS 0.087217f
C31320 VDD.t1387 VSS 0.066856f
C31321 VDD.n10979 VSS 0.14405f
C31322 VDD.n10980 VSS 0.120118f
C31323 VDD.n10981 VSS 0.016021f
C31324 VDD.t1504 VSS 0.025104f
C31325 VDD.n10982 VSS 0.116823f
C31326 VDD.n10983 VSS 0.785619f
C31327 VDD.t3141 VSS 0.028519f
C31328 VDD.t4607 VSS 0.028519f
C31329 VDD.n10984 VSS 0.009191f
C31330 VDD.n10985 VSS 0.311617f
C31331 VDD.t4606 VSS 0.066856f
C31332 VDD.t919 VSS 0.066856f
C31333 VDD.n10986 VSS 0.715442f
C31334 VDD.t4327 VSS 0.028519f
C31335 VDD.t4163 VSS 0.028519f
C31336 VDD.n10987 VSS 0.009191f
C31337 VDD.n10988 VSS 0.650522f
C31338 VDD.t4162 VSS 0.066856f
C31339 VDD.t3246 VSS 0.066856f
C31340 VDD.n10989 VSS 0.696076f
C31341 VDD.t4496 VSS 0.066856f
C31342 VDD.t3566 VSS 0.066856f
C31343 VDD.n10990 VSS 0.696076f
C31344 VDD.t4699 VSS 0.028519f
C31345 VDD.t4497 VSS 0.028519f
C31346 VDD.n10991 VSS 0.009191f
C31347 VDD.n10992 VSS 0.475536f
C31348 VDD.n10993 VSS 0.529799f
C31349 VDD.n10994 VSS 0.208534f
C31350 VDD.n10995 VSS 0.902999f
C31351 VDD.n10996 VSS 0.902999f
C31352 VDD.t748 VSS 1.45794f
C31353 VDD.t947 VSS 1.96535f
C31354 VDD.t323 VSS 1.96535f
C31355 VDD.t301 VSS 1.31955f
C31356 VDD.n10997 VSS 0.595476f
C31357 VDD.n10998 VSS 0.208771f
C31358 VDD.n10999 VSS 0.208534f
C31359 VDD.n11000 VSS 0.524869f
C31360 VDD.n11001 VSS 0.207221f
C31361 VDD.n11002 VSS 0.865258f
C31362 VDD.t1115 VSS 1.45794f
C31363 VDD.t2234 VSS 1.96535f
C31364 VDD.t527 VSS 1.96535f
C31365 VDD.t524 VSS 1.31955f
C31366 VDD.n11003 VSS 0.595476f
C31367 VDD.n11004 VSS 0.645798f
C31368 VDD.t525 VSS 1.36988f
C31369 VDD.t526 VSS 1.96535f
C31370 VDD.t1749 VSS 1.96535f
C31371 VDD.t1357 VSS 1.45794f
C31372 VDD.n11005 VSS 0.865258f
C31373 VDD.n11006 VSS 0.208534f
C31374 VDD.n11007 VSS 0.524869f
C31375 VDD.t1731 VSS 0.028519f
C31376 VDD.t2171 VSS 0.028519f
C31377 VDD.n11008 VSS 0.009191f
C31378 VDD.t4349 VSS 0.028519f
C31379 VDD.t2049 VSS 0.028519f
C31380 VDD.n11009 VSS 0.009191f
C31381 VDD.n11010 VSS 0.471397f
C31382 VDD.t1730 VSS 0.066856f
C31383 VDD.t4348 VSS 0.066856f
C31384 VDD.t2048 VSS 0.066856f
C31385 VDD.t2170 VSS 0.066856f
C31386 VDD.n11011 VSS 0.690489f
C31387 VDD.t1356 VSS 0.066856f
C31388 VDD.t3982 VSS 0.066856f
C31389 VDD.t1643 VSS 0.066856f
C31390 VDD.t1748 VSS 0.066856f
C31391 VDD.n11012 VSS 0.690489f
C31392 VDD.t1358 VSS 0.028519f
C31393 VDD.t1750 VSS 0.028519f
C31394 VDD.n11013 VSS 0.009191f
C31395 VDD.t3983 VSS 0.028519f
C31396 VDD.t1645 VSS 0.028519f
C31397 VDD.n11014 VSS 0.009191f
C31398 VDD.n11015 VSS 0.644755f
C31399 VDD.t2070 VSS 0.066856f
C31400 VDD.t1421 VSS 0.066856f
C31401 VDD.t2364 VSS 0.066856f
C31402 VDD.t2868 VSS 0.066856f
C31403 VDD.n11016 VSS 0.709674f
C31404 VDD.t2071 VSS 0.028519f
C31405 VDD.t2869 VSS 0.028519f
C31406 VDD.n11017 VSS 0.009191f
C31407 VDD.t1423 VSS 0.028519f
C31408 VDD.t2365 VSS 0.028519f
C31409 VDD.n11018 VSS 0.009191f
C31410 VDD.n11019 VSS 0.309003f
C31411 VDD.n11020 VSS 0.765686f
C31412 VDD.n11021 VSS 0.116823f
C31413 VDD.t3693 VSS 0.066856f
C31414 VDD.n11022 VSS 0.14405f
C31415 VDD.n11023 VSS 0.120118f
C31416 VDD.n11024 VSS 0.016021f
C31417 VDD.t2616 VSS 0.025104f
C31418 VDD.n11025 VSS 0.087217f
C31419 VDD.n11026 VSS 0.057098f
C31420 VDD.n11027 VSS 0.208771f
C31421 VDD.n11028 VSS 0.595476f
C31422 VDD.n11029 VSS 0.645798f
C31423 VDD.n11030 VSS 0.206947f
C31424 VDD.n11031 VSS 0.048151f
C31425 VDD.n11032 VSS 0.081176f
C31426 VDD.t1243 VSS 0.066856f
C31427 VDD.n11033 VSS 0.125227f
C31428 VDD.n11034 VSS 0.101294f
C31429 VDD.n11035 VSS 0.016021f
C31430 VDD.t3592 VSS 0.025104f
C31431 VDD.n11036 VSS 0.099723f
C31432 VDD.n11037 VSS 0.126402f
C31433 VDD.n11038 VSS 0.171327f
C31434 VDD.n11039 VSS 0.012131f
C31435 VDD.n11040 VSS 0.012131f
C31436 VDD.n11041 VSS 0.012131f
C31437 VDD.n11042 VSS 0.012131f
C31438 VDD.n11043 VSS 0.106603f
C31439 VDD.n11044 VSS 0.134523f
C31440 VDD.n11045 VSS 0.01487f
C31441 VDD.n11046 VSS 0.134523f
C31442 VDD.n11047 VSS 0.01502f
C31443 VDD.n11048 VSS 0.074876f
C31444 VDD.n11049 VSS 0.201785f
C31445 VDD.n11050 VSS 0.269046f
C31446 VDD.n11051 VSS 0.012131f
C31447 VDD.n11052 VSS 0.012131f
C31448 VDD.n11053 VSS 0.012131f
C31449 VDD.n11054 VSS 0.269046f
C31450 VDD.n11055 VSS 0.269046f
C31451 VDD.t1313 VSS 0.028519f
C31452 VDD.t2800 VSS 0.028519f
C31453 VDD.n11056 VSS 0.009191f
C31454 VDD.n11057 VSS 0.149927f
C31455 VDD.n11058 VSS 0.145945f
C31456 VDD.n11059 VSS 0.012131f
C31457 VDD.n11060 VSS 0.012131f
C31458 VDD.n11061 VSS 0.012131f
C31459 VDD.n11062 VSS 0.255086f
C31460 VDD.t1312 VSS 0.066856f
C31461 VDD.t2799 VSS 0.066856f
C31462 VDD.n11063 VSS 0.182387f
C31463 VDD.n11064 VSS 0.148483f
C31464 VDD.n11065 VSS 0.269046f
C31465 VDD.n11066 VSS 0.012131f
C31466 VDD.n11067 VSS 0.012131f
C31467 VDD.n11068 VSS 0.012131f
C31468 VDD.n11069 VSS 0.269046f
C31469 VDD.n11070 VSS 0.269046f
C31470 VDD.n11071 VSS 0.171327f
C31471 VDD.n11072 VSS 0.012131f
C31472 VDD.n11073 VSS 0.012131f
C31473 VDD.n11074 VSS 0.232243f
C31474 VDD.n11075 VSS 0.269046f
C31475 VDD.t3883 VSS 0.028519f
C31476 VDD.t1103 VSS 0.028519f
C31477 VDD.n11076 VSS 0.009191f
C31478 VDD.n11077 VSS 0.149927f
C31479 VDD.n11078 VSS 0.145945f
C31480 VDD.n11079 VSS 0.012131f
C31481 VDD.n11080 VSS 0.012131f
C31482 VDD.n11081 VSS 0.012131f
C31483 VDD.n11082 VSS 0.269046f
C31484 VDD.n11083 VSS 0.269046f
C31485 VDD.n11084 VSS 0.142138f
C31486 VDD.n11085 VSS 0.012131f
C31487 VDD.n11086 VSS 0.012131f
C31488 VDD.n11087 VSS 0.261432f
C31489 VDD.n11088 VSS 0.269046f
C31490 VDD.t1296 VSS 0.028519f
C31491 VDD.t2792 VSS 0.028519f
C31492 VDD.n11089 VSS 0.009191f
C31493 VDD.n11090 VSS 0.149927f
C31494 VDD.n11091 VSS 0.176403f
C31495 VDD.n11092 VSS 0.012131f
C31496 VDD.n11093 VSS 0.012131f
C31497 VDD.n11094 VSS 0.012131f
C31498 VDD.n11095 VSS 0.269046f
C31499 VDD.n11096 VSS 0.151021f
C31500 VDD.t1295 VSS 0.066856f
C31501 VDD.t2791 VSS 0.066856f
C31502 VDD.n11097 VSS 0.182387f
C31503 VDD.n11098 VSS 0.252548f
C31504 VDD.n11099 VSS 0.012131f
C31505 VDD.n11100 VSS 0.012131f
C31506 VDD.n11101 VSS 0.012131f
C31507 VDD.n11102 VSS 0.269046f
C31508 VDD.n11103 VSS 0.269046f
C31509 VDD.n11104 VSS 0.201785f
C31510 VDD.n11105 VSS 0.012131f
C31511 VDD.n11106 VSS 0.012131f
C31512 VDD.n11107 VSS 0.201785f
C31513 VDD.n11108 VSS 0.269046f
C31514 VDD.n11109 VSS 0.176403f
C31515 VDD.n11110 VSS 0.012131f
C31516 VDD.n11111 VSS 0.012131f
C31517 VDD.n11112 VSS 0.227166f
C31518 VDD.n11113 VSS 0.269046f
C31519 VDD.n11114 VSS 0.269046f
C31520 VDD.n11115 VSS 0.012131f
C31521 VDD.n11116 VSS 0.012131f
C31522 VDD.n11117 VSS 0.012131f
C31523 VDD.n11118 VSS 0.262701f
C31524 VDD.t3942 VSS 0.066856f
C31525 VDD.t2043 VSS 0.066856f
C31526 VDD.n11119 VSS 0.182387f
C31527 VDD.n11120 VSS 0.140868f
C31528 VDD.n11121 VSS 0.261432f
C31529 VDD.n11122 VSS 0.012131f
C31530 VDD.n11123 VSS 0.11041f
C31531 VDD.n11124 VSS 0.012131f
C31532 VDD.n11125 VSS 0.012131f
C31533 VDD.n11126 VSS 0.107872f
C31534 VDD.n11127 VSS 0.031727f
C31535 VDD.n11129 VSS 0.018249f
C31536 VDD.n11130 VSS 0.134523f
C31537 VDD.n11131 VSS 0.266508f
C31538 VDD.n11132 VSS 0.012131f
C31539 VDD.n11133 VSS 0.012131f
C31540 VDD.n11134 VSS 0.012131f
C31541 VDD.n11135 VSS 0.324292f
C31542 VDD.n11136 VSS 0.075648f
C31543 VDD.n11137 VSS 0.012131f
C31544 VDD.n11138 VSS 0.012131f
C31545 VDD.n11139 VSS 0.012131f
C31546 VDD.n11140 VSS 0.012131f
C31547 VDD.n11141 VSS 0.012131f
C31548 VDD.n11142 VSS 0.012131f
C31549 VDD.n11143 VSS 0.012131f
C31550 VDD.n11144 VSS 0.012131f
C31551 VDD.n11145 VSS 0.012131f
C31552 VDD.n11146 VSS 0.012131f
C31553 VDD.n11147 VSS 0.012131f
C31554 VDD.n11148 VSS 0.012131f
C31555 VDD.n11149 VSS 0.012131f
C31556 VDD.n11150 VSS 0.012131f
C31557 VDD.n11151 VSS 0.012131f
C31558 VDD.n11152 VSS 0.012131f
C31559 VDD.n11153 VSS 0.012131f
C31560 VDD.n11154 VSS 0.012131f
C31561 VDD.n11155 VSS 0.012131f
C31562 VDD.n11156 VSS 0.012131f
C31563 VDD.n11157 VSS 0.012131f
C31564 VDD.n11158 VSS 0.012131f
C31565 VDD.n11159 VSS 0.012131f
C31566 VDD.n11160 VSS 0.012131f
C31567 VDD.n11161 VSS 0.012131f
C31568 VDD.n11162 VSS 0.012131f
C31569 VDD.n11163 VSS 0.012131f
C31570 VDD.n11164 VSS 0.012131f
C31571 VDD.n11165 VSS 0.012131f
C31572 VDD.n11166 VSS 0.012131f
C31573 VDD.n11167 VSS 0.012131f
C31574 VDD.n11168 VSS 0.012131f
C31575 VDD.n11169 VSS 0.012131f
C31576 VDD.n11170 VSS 0.012131f
C31577 VDD.n11171 VSS 0.012131f
C31578 VDD.n11172 VSS 0.012131f
C31579 VDD.n11173 VSS 0.012131f
C31580 VDD.n11174 VSS 0.012131f
C31581 VDD.n11175 VSS 0.012131f
C31582 VDD.n11176 VSS 0.012131f
C31583 VDD.n11177 VSS 0.012131f
C31584 VDD.n11178 VSS 0.012131f
C31585 VDD.n11179 VSS 0.012131f
C31586 VDD.n11180 VSS 0.012131f
C31587 VDD.n11181 VSS 0.012131f
C31588 VDD.n11182 VSS 0.012131f
C31589 VDD.n11183 VSS 0.012131f
C31590 VDD.n11184 VSS 0.012131f
C31591 VDD.n11185 VSS 0.012131f
C31592 VDD.n11186 VSS 0.012131f
C31593 VDD.n11187 VSS 0.012131f
C31594 VDD.n11188 VSS 0.012131f
C31595 VDD.n11189 VSS 0.012131f
C31596 VDD.n11190 VSS 0.012131f
C31597 VDD.n11191 VSS 0.012131f
C31598 VDD.n11192 VSS 0.012131f
C31599 VDD.n11193 VSS 0.012131f
C31600 VDD.n11194 VSS 0.012131f
C31601 VDD.n11195 VSS 0.012131f
C31602 VDD.n11196 VSS 0.012131f
C31603 VDD.n11197 VSS 0.012131f
C31604 VDD.n11198 VSS 0.012131f
C31605 VDD.n11199 VSS 0.012131f
C31606 VDD.n11200 VSS 0.012131f
C31607 VDD.n11201 VSS 0.012131f
C31608 VDD.n11202 VSS 0.012131f
C31609 VDD.n11203 VSS 0.012131f
C31610 VDD.n11204 VSS 0.012131f
C31611 VDD.n11205 VSS 0.012131f
C31612 VDD.n11206 VSS 0.012131f
C31613 VDD.n11207 VSS 0.012131f
C31614 VDD.n11208 VSS 0.012131f
C31615 VDD.n11209 VSS 0.012131f
C31616 VDD.n11210 VSS 0.012131f
C31617 VDD.n11211 VSS 0.012131f
C31618 VDD.n11212 VSS 0.012131f
C31619 VDD.n11213 VSS 0.012131f
C31620 VDD.n11214 VSS 0.012131f
C31621 VDD.n11215 VSS 0.012131f
C31622 VDD.n11216 VSS 0.012131f
C31623 VDD.n11217 VSS 0.012131f
C31624 VDD.n11218 VSS 0.012131f
C31625 VDD.n11219 VSS 0.012131f
C31626 VDD.n11220 VSS 0.012131f
C31627 VDD.n11221 VSS 0.012131f
C31628 VDD.n11222 VSS 0.012131f
C31629 VDD.n11223 VSS 0.012131f
C31630 VDD.n11224 VSS 0.012131f
C31631 VDD.n11225 VSS 0.012131f
C31632 VDD.n11226 VSS 0.012131f
C31633 VDD.n11227 VSS 0.012131f
C31634 VDD.n11228 VSS 0.012131f
C31635 VDD.n11229 VSS 0.012131f
C31636 VDD.n11230 VSS 0.012131f
C31637 VDD.n11231 VSS 0.012131f
C31638 VDD.n11232 VSS 0.012131f
C31639 VDD.n11233 VSS 0.012131f
C31640 VDD.n11234 VSS 0.012131f
C31641 VDD.n11235 VSS 0.012131f
C31642 VDD.n11236 VSS 0.012131f
C31643 VDD.n11237 VSS 0.012131f
C31644 VDD.n11238 VSS 0.012131f
C31645 VDD.n11239 VSS 0.012131f
C31646 VDD.n11240 VSS 0.012131f
C31647 VDD.n11241 VSS 0.012131f
C31648 VDD.n11242 VSS 0.012131f
C31649 VDD.n11243 VSS 0.012131f
C31650 VDD.n11244 VSS 0.012131f
C31651 VDD.n11245 VSS 0.012131f
C31652 VDD.n11246 VSS 0.012131f
C31653 VDD.n11247 VSS 0.012131f
C31654 VDD.n11248 VSS 0.012131f
C31655 VDD.n11249 VSS 0.012131f
C31656 VDD.n11250 VSS 0.012131f
C31657 VDD.n11251 VSS 0.012131f
C31658 VDD.n11252 VSS 0.012131f
C31659 VDD.n11253 VSS 0.012131f
C31660 VDD.n11254 VSS 0.012131f
C31661 VDD.n11255 VSS 0.012131f
C31662 VDD.n11256 VSS 0.012131f
C31663 VDD.n11257 VSS 0.012131f
C31664 VDD.n11258 VSS 0.012131f
C31665 VDD.n11259 VSS 0.012131f
C31666 VDD.n11260 VSS 0.012131f
C31667 VDD.n11261 VSS 0.012131f
C31668 VDD.n11262 VSS 0.012131f
C31669 VDD.n11263 VSS 0.012131f
C31670 VDD.n11264 VSS 0.012131f
C31671 VDD.n11265 VSS 0.012131f
C31672 VDD.n11266 VSS 0.012131f
C31673 VDD.n11267 VSS 0.012131f
C31674 VDD.n11268 VSS 0.012131f
C31675 VDD.n11269 VSS 0.012131f
C31676 VDD.n11270 VSS 0.012131f
C31677 VDD.n11271 VSS 0.012131f
C31678 VDD.n11272 VSS 0.012131f
C31679 VDD.n11273 VSS 0.012131f
C31680 VDD.n11274 VSS 0.012131f
C31681 VDD.n11275 VSS 0.012131f
C31682 VDD.n11276 VSS 0.012131f
C31683 VDD.n11277 VSS 0.012131f
C31684 VDD.n11278 VSS 0.012131f
C31685 VDD.n11279 VSS 0.012131f
C31686 VDD.n11280 VSS 0.012131f
C31687 VDD.n11281 VSS 0.012131f
C31688 VDD.n11282 VSS 0.012131f
C31689 VDD.n11283 VSS 0.012131f
C31690 VDD.n11284 VSS 0.012131f
C31691 VDD.n11285 VSS 0.012131f
C31692 VDD.n11286 VSS 0.012131f
C31693 VDD.n11287 VSS 0.012131f
C31694 VDD.n11288 VSS 0.012131f
C31695 VDD.n11289 VSS 0.012131f
C31696 VDD.n11290 VSS 0.012131f
C31697 VDD.n11291 VSS 0.012131f
C31698 VDD.n11292 VSS 0.012131f
C31699 VDD.n11293 VSS 0.012131f
C31700 VDD.n11294 VSS 0.012131f
C31701 VDD.n11295 VSS 0.012131f
C31702 VDD.n11296 VSS 0.012131f
C31703 VDD.n11297 VSS 0.012131f
C31704 VDD.n11298 VSS 0.012131f
C31705 VDD.n11299 VSS 0.012131f
C31706 VDD.n11300 VSS 0.012131f
C31707 VDD.n11301 VSS 0.012131f
C31708 VDD.n11302 VSS 0.012131f
C31709 VDD.n11303 VSS 0.012131f
C31710 VDD.n11304 VSS 0.012131f
C31711 VDD.n11305 VSS 0.012131f
C31712 VDD.n11306 VSS 0.012131f
C31713 VDD.n11307 VSS 0.012131f
C31714 VDD.n11308 VSS 0.012131f
C31715 VDD.n11309 VSS 0.012131f
C31716 VDD.n11310 VSS 0.012131f
C31717 VDD.n11311 VSS 0.012131f
C31718 VDD.n11312 VSS 0.012131f
C31719 VDD.n11313 VSS 0.012131f
C31720 VDD.n11314 VSS 0.012131f
C31721 VDD.n11315 VSS 0.012131f
C31722 VDD.n11316 VSS 0.012131f
C31723 VDD.n11317 VSS 0.012131f
C31724 VDD.n11318 VSS 0.012131f
C31725 VDD.n11319 VSS 0.012131f
C31726 VDD.n11320 VSS 0.012131f
C31727 VDD.n11321 VSS 0.012131f
C31728 VDD.n11322 VSS 0.012131f
C31729 VDD.n11323 VSS 0.012131f
C31730 VDD.n11324 VSS 0.012131f
C31731 VDD.n11325 VSS 0.012131f
C31732 VDD.n11326 VSS 0.012131f
C31733 VDD.n11327 VSS 0.012131f
C31734 VDD.n11328 VSS 0.012131f
C31735 VDD.n11329 VSS 0.012131f
C31736 VDD.n11330 VSS 0.012131f
C31737 VDD.n11331 VSS 0.012131f
C31738 VDD.n11332 VSS 0.012131f
C31739 VDD.n11333 VSS 0.012131f
C31740 VDD.n11334 VSS 0.012131f
C31741 VDD.n11335 VSS 0.012131f
C31742 VDD.n11336 VSS 0.012131f
C31743 VDD.n11337 VSS 0.012131f
C31744 VDD.n11338 VSS 0.012131f
C31745 VDD.n11339 VSS 0.012131f
C31746 VDD.n11340 VSS 0.012131f
C31747 VDD.n11341 VSS 0.012131f
C31748 VDD.n11342 VSS 0.012131f
C31749 VDD.n11343 VSS 0.012131f
C31750 VDD.n11344 VSS 0.012131f
C31751 VDD.n11345 VSS 0.012131f
C31752 VDD.n11346 VSS 0.012131f
C31753 VDD.n11347 VSS 0.012131f
C31754 VDD.n11348 VSS 0.012131f
C31755 VDD.n11349 VSS 0.012131f
C31756 VDD.n11350 VSS 0.012131f
C31757 VDD.n11351 VSS 0.012131f
C31758 VDD.n11352 VSS 0.012131f
C31759 VDD.n11353 VSS 0.012131f
C31760 VDD.n11354 VSS 0.012131f
C31761 VDD.n11355 VSS 0.012131f
C31762 VDD.n11356 VSS 0.012131f
C31763 VDD.n11357 VSS 0.012131f
C31764 VDD.n11358 VSS 0.012131f
C31765 VDD.n11359 VSS 0.012131f
C31766 VDD.n11360 VSS 0.012131f
C31767 VDD.n11361 VSS 0.012131f
C31768 VDD.n11362 VSS 0.012131f
C31769 VDD.n11363 VSS 0.012131f
C31770 VDD.n11364 VSS 0.012131f
C31771 VDD.n11365 VSS 0.012131f
C31772 VDD.n11366 VSS 0.012131f
C31773 VDD.n11367 VSS 0.012131f
C31774 VDD.n11368 VSS 0.012131f
C31775 VDD.n11369 VSS 0.012131f
C31776 VDD.n11370 VSS 0.012131f
C31777 VDD.n11371 VSS 0.012131f
C31778 VDD.n11372 VSS 0.012131f
C31779 VDD.n11373 VSS 0.012131f
C31780 VDD.n11374 VSS 0.012131f
C31781 VDD.n11375 VSS 0.012131f
C31782 VDD.n11376 VSS 0.012131f
C31783 VDD.n11377 VSS 0.012131f
C31784 VDD.n11378 VSS 0.012131f
C31785 VDD.n11379 VSS 0.012131f
C31786 VDD.n11380 VSS 0.012131f
C31787 VDD.n11381 VSS 0.012131f
C31788 VDD.n11382 VSS 0.012131f
C31789 VDD.n11383 VSS 0.012131f
C31790 VDD.n11384 VSS 0.012131f
C31791 VDD.n11385 VSS 0.012131f
C31792 VDD.n11386 VSS 0.012131f
C31793 VDD.n11387 VSS 0.012131f
C31794 VDD.n11388 VSS 0.012131f
C31795 VDD.n11389 VSS 0.012131f
C31796 VDD.n11390 VSS 0.012131f
C31797 VDD.n11391 VSS 0.012131f
C31798 VDD.n11392 VSS 0.012131f
C31799 VDD.n11393 VSS 0.012131f
C31800 VDD.n11394 VSS 0.012131f
C31801 VDD.n11395 VSS 0.012131f
C31802 VDD.n11396 VSS 0.012131f
C31803 VDD.n11397 VSS 0.012131f
C31804 VDD.n11398 VSS 0.012131f
C31805 VDD.n11399 VSS 0.012131f
C31806 VDD.n11400 VSS 0.012131f
C31807 VDD.n11401 VSS 0.012131f
C31808 VDD.n11402 VSS 0.012131f
C31809 VDD.n11403 VSS 0.012131f
C31810 VDD.n11404 VSS 0.012131f
C31811 VDD.n11405 VSS 0.012131f
C31812 VDD.n11406 VSS 0.012131f
C31813 VDD.n11407 VSS 0.012131f
C31814 VDD.n11408 VSS 0.012131f
C31815 VDD.n11409 VSS 0.012131f
C31816 VDD.n11410 VSS 0.012131f
C31817 VDD.n11411 VSS 0.012131f
C31818 VDD.n11412 VSS 0.012131f
C31819 VDD.n11413 VSS 0.012131f
C31820 VDD.n11414 VSS 0.012131f
C31821 VDD.n11415 VSS 0.012131f
C31822 VDD.n11416 VSS 0.012131f
C31823 VDD.n11417 VSS 0.012131f
C31824 VDD.n11418 VSS 0.012131f
C31825 VDD.n11419 VSS 0.012131f
C31826 VDD.n11420 VSS 0.012131f
C31827 VDD.n11421 VSS 0.012131f
C31828 VDD.n11422 VSS 0.012131f
C31829 VDD.n11423 VSS 0.012131f
C31830 VDD.n11424 VSS 0.012131f
C31831 VDD.n11425 VSS 0.012131f
C31832 VDD.n11426 VSS 0.012131f
C31833 VDD.n11427 VSS 0.012131f
C31834 VDD.n11428 VSS 0.012131f
C31835 VDD.n11429 VSS 0.012131f
C31836 VDD.n11430 VSS 0.012131f
C31837 VDD.n11431 VSS 0.012131f
C31838 VDD.n11432 VSS 0.012131f
C31839 VDD.n11433 VSS 0.012131f
C31840 VDD.n11434 VSS 0.012131f
C31841 VDD.n11435 VSS 0.012131f
C31842 VDD.n11436 VSS 0.012131f
C31843 VDD.n11437 VSS 0.012131f
C31844 VDD.n11438 VSS 0.012131f
C31845 VDD.n11439 VSS 0.012131f
C31846 VDD.n11440 VSS 0.012131f
C31847 VDD.n11441 VSS 0.012131f
C31848 VDD.n11442 VSS 0.012131f
C31849 VDD.n11443 VSS 0.012131f
C31850 VDD.n11444 VSS 0.012131f
C31851 VDD.n11445 VSS 0.012131f
C31852 VDD.n11446 VSS 0.012131f
C31853 VDD.n11447 VSS 0.012131f
C31854 VDD.n11448 VSS 0.012131f
C31855 VDD.n11449 VSS 0.012131f
C31856 VDD.n11450 VSS 0.012131f
C31857 VDD.n11451 VSS 0.012131f
C31858 VDD.n11452 VSS 0.012131f
C31859 VDD.n11453 VSS 0.012131f
C31860 VDD.n11454 VSS 0.012131f
C31861 VDD.n11455 VSS 0.012131f
C31862 VDD.n11456 VSS 0.012131f
C31863 VDD.n11457 VSS 0.012131f
C31864 VDD.n11458 VSS 0.012131f
C31865 VDD.n11459 VSS 0.012131f
C31866 VDD.n11460 VSS 0.012131f
C31867 VDD.n11461 VSS 0.012131f
C31868 VDD.n11462 VSS 0.012131f
C31869 VDD.n11463 VSS 0.012131f
C31870 VDD.n11464 VSS 0.012131f
C31871 VDD.n11465 VSS 0.012131f
C31872 VDD.n11466 VSS 0.012131f
C31873 VDD.n11467 VSS 0.012131f
C31874 VDD.n11468 VSS 0.012131f
C31875 VDD.n11469 VSS 0.012131f
C31876 VDD.n11470 VSS 0.012131f
C31877 VDD.n11471 VSS 0.012131f
C31878 VDD.n11472 VSS 0.012131f
C31879 VDD.n11473 VSS 0.012131f
C31880 VDD.n11474 VSS 0.012131f
C31881 VDD.n11475 VSS 0.012131f
C31882 VDD.n11476 VSS 0.012131f
C31883 VDD.n11477 VSS 0.012131f
C31884 VDD.n11478 VSS 0.012131f
C31885 VDD.n11479 VSS 0.012131f
C31886 VDD.n11480 VSS 0.012131f
C31887 VDD.n11481 VSS 0.012131f
C31888 VDD.n11482 VSS 0.012131f
C31889 VDD.n11483 VSS 0.012131f
C31890 VDD.n11484 VSS 0.012131f
C31891 VDD.n11485 VSS 0.012131f
C31892 VDD.n11486 VSS 0.012131f
C31893 VDD.n11487 VSS 0.012131f
C31894 VDD.n11488 VSS 0.012131f
C31895 VDD.n11489 VSS 0.012131f
C31896 VDD.n11490 VSS 0.012131f
C31897 VDD.n11491 VSS 0.012131f
C31898 VDD.n11492 VSS 0.012131f
C31899 VDD.n11493 VSS 0.012131f
C31900 VDD.n11494 VSS 0.012131f
C31901 VDD.n11495 VSS 0.012131f
C31902 VDD.n11496 VSS 0.012131f
C31903 VDD.n11497 VSS 0.012131f
C31904 VDD.n11498 VSS 0.012131f
C31905 VDD.n11499 VSS 0.012131f
C31906 VDD.n11500 VSS 0.012131f
C31907 VDD.n11501 VSS 0.012131f
C31908 VDD.n11502 VSS 0.012131f
C31909 VDD.n11503 VSS 0.012131f
C31910 VDD.n11504 VSS 0.012131f
C31911 VDD.n11505 VSS 0.012131f
C31912 VDD.n11506 VSS 0.012131f
C31913 VDD.n11507 VSS 0.012131f
C31914 VDD.n11508 VSS 0.012131f
C31915 VDD.n11509 VSS 0.012131f
C31916 VDD.n11510 VSS 0.012131f
C31917 VDD.n11511 VSS 0.012131f
C31918 VDD.n11512 VSS 0.012131f
C31919 VDD.n11513 VSS 0.012131f
C31920 VDD.n11514 VSS 0.012131f
C31921 VDD.n11515 VSS 0.012131f
C31922 VDD.n11516 VSS 0.012131f
C31923 VDD.n11517 VSS 0.012131f
C31924 VDD.n11518 VSS 0.012131f
C31925 VDD.n11519 VSS 0.012131f
C31926 VDD.n11520 VSS 0.012131f
C31927 VDD.n11521 VSS 0.012131f
C31928 VDD.n11522 VSS 0.012131f
C31929 VDD.n11523 VSS 0.012131f
C31930 VDD.n11524 VSS 0.012131f
C31931 VDD.n11525 VSS 0.012131f
C31932 VDD.n11526 VSS 0.012131f
C31933 VDD.n11527 VSS 0.012131f
C31934 VDD.n11528 VSS 0.012131f
C31935 VDD.n11529 VSS 0.012131f
C31936 VDD.n11530 VSS 0.012131f
C31937 VDD.n11531 VSS 0.012131f
C31938 VDD.n11532 VSS 0.012131f
C31939 VDD.n11533 VSS 0.012131f
C31940 VDD.n11534 VSS 0.012131f
C31941 VDD.n11535 VSS 0.012131f
C31942 VDD.n11536 VSS 0.012131f
C31943 VDD.n11537 VSS 0.012131f
C31944 VDD.n11538 VSS 0.012131f
C31945 VDD.n11539 VSS 0.012131f
C31946 VDD.n11540 VSS 0.012131f
C31947 VDD.n11541 VSS 0.012131f
C31948 VDD.n11542 VSS 0.012131f
C31949 VDD.n11543 VSS 0.012131f
C31950 VDD.n11544 VSS 0.012131f
C31951 VDD.n11545 VSS 0.012131f
C31952 VDD.n11546 VSS 0.012131f
C31953 VDD.n11547 VSS 0.012131f
C31954 VDD.n11548 VSS 0.012131f
C31955 VDD.n11549 VSS 0.012131f
C31956 VDD.n11550 VSS 0.012131f
C31957 VDD.n11551 VSS 0.012131f
C31958 VDD.n11552 VSS 0.012131f
C31959 VDD.n11553 VSS 0.012131f
C31960 VDD.n11554 VSS 0.012131f
C31961 VDD.n11555 VSS 0.012131f
C31962 VDD.n11556 VSS 0.012131f
C31963 VDD.n11557 VSS 0.012131f
C31964 VDD.n11558 VSS 0.012131f
C31965 VDD.n11559 VSS 0.012131f
C31966 VDD.n11560 VSS 0.012131f
C31967 VDD.n11561 VSS 0.012131f
C31968 VDD.n11562 VSS 0.012131f
C31969 VDD.n11563 VSS 0.012131f
C31970 VDD.n11564 VSS 0.012131f
C31971 VDD.n11565 VSS 0.012131f
C31972 VDD.n11566 VSS 0.012131f
C31973 VDD.n11567 VSS 0.012131f
C31974 VDD.n11568 VSS 0.012131f
C31975 VDD.n11569 VSS 0.012131f
C31976 VDD.n11570 VSS 0.012131f
C31977 VDD.n11571 VSS 0.012131f
C31978 VDD.n11572 VSS 0.012131f
C31979 VDD.n11573 VSS 0.012131f
C31980 VDD.n11574 VSS 0.012131f
C31981 VDD.n11575 VSS 0.012131f
C31982 VDD.n11576 VSS 0.012131f
C31983 VDD.n11577 VSS 0.012131f
C31984 VDD.n11578 VSS 0.012131f
C31985 VDD.n11579 VSS 0.012131f
C31986 VDD.n11580 VSS 0.012131f
C31987 VDD.n11581 VSS 0.012131f
C31988 VDD.n11582 VSS 0.012131f
C31989 VDD.n11583 VSS 0.012131f
C31990 VDD.n11584 VSS 0.012131f
C31991 VDD.n11585 VSS 0.012131f
C31992 VDD.n11586 VSS 0.012131f
C31993 VDD.n11587 VSS 0.012131f
C31994 VDD.n11588 VSS 0.012131f
C31995 VDD.n11589 VSS 0.012131f
C31996 VDD.n11590 VSS 0.012131f
C31997 VDD.n11591 VSS 0.012131f
C31998 VDD.n11592 VSS 0.012131f
C31999 VDD.n11593 VSS 0.012131f
C32000 VDD.n11594 VSS 0.012131f
C32001 VDD.n11595 VSS 0.012131f
C32002 VDD.n11596 VSS 0.012131f
C32003 VDD.n11597 VSS 0.012131f
C32004 VDD.n11598 VSS 0.012131f
C32005 VDD.n11599 VSS 0.012131f
C32006 VDD.n11600 VSS 0.012131f
C32007 VDD.n11601 VSS 0.012131f
C32008 VDD.n11602 VSS 0.012131f
C32009 VDD.n11603 VSS 0.012131f
C32010 VDD.n11604 VSS 0.012131f
C32011 VDD.n11605 VSS 0.012131f
C32012 VDD.n11606 VSS 0.012131f
C32013 VDD.n11607 VSS 0.012131f
C32014 VDD.n11608 VSS 0.012131f
C32015 VDD.n11609 VSS 0.012131f
C32016 VDD.n11610 VSS 0.012131f
C32017 VDD.n11611 VSS 0.012131f
C32018 VDD.n11612 VSS 0.012131f
C32019 VDD.n11613 VSS 0.012131f
C32020 VDD.n11614 VSS 0.012131f
C32021 VDD.n11615 VSS 0.012131f
C32022 VDD.n11616 VSS 0.012131f
C32023 VDD.n11617 VSS 0.012131f
C32024 VDD.n11618 VSS 0.012131f
C32025 VDD.n11619 VSS 0.012131f
C32026 VDD.n11620 VSS 0.012131f
C32027 VDD.n11621 VSS 0.012131f
C32028 VDD.n11622 VSS 0.012131f
C32029 VDD.n11623 VSS 0.012131f
C32030 VDD.n11624 VSS 0.012131f
C32031 VDD.n11625 VSS 0.012131f
C32032 VDD.n11626 VSS 0.012131f
C32033 VDD.n11627 VSS 0.012131f
C32034 VDD.n11628 VSS 0.012131f
C32035 VDD.n11629 VSS 0.012131f
C32036 VDD.n11630 VSS 0.012131f
C32037 VDD.n11631 VSS 0.012131f
C32038 VDD.n11632 VSS 0.012131f
C32039 VDD.n11633 VSS 0.012131f
C32040 VDD.n11634 VSS 0.012131f
C32041 VDD.n11635 VSS 0.012131f
C32042 VDD.n11636 VSS 0.012131f
C32043 VDD.n11637 VSS 0.012131f
C32044 VDD.n11638 VSS 0.012131f
C32045 VDD.n11639 VSS 0.012131f
C32046 VDD.n11640 VSS 0.012131f
C32047 VDD.n11641 VSS 0.012131f
C32048 VDD.n11642 VSS 0.012131f
C32049 VDD.n11643 VSS 0.012131f
C32050 VDD.n11644 VSS 0.012131f
C32051 VDD.n11645 VSS 0.012131f
C32052 VDD.n11646 VSS 0.012131f
C32053 VDD.n11647 VSS 0.012131f
C32054 VDD.n11648 VSS 0.012131f
C32055 VDD.n11649 VSS 0.012131f
C32056 VDD.n11650 VSS 0.012131f
C32057 VDD.n11651 VSS 0.012131f
C32058 VDD.n11652 VSS 0.012131f
C32059 VDD.n11653 VSS 0.012131f
C32060 VDD.n11654 VSS 0.012131f
C32061 VDD.n11655 VSS 0.012131f
C32062 VDD.n11656 VSS 0.012131f
C32063 VDD.n11657 VSS 0.012131f
C32064 VDD.n11658 VSS 0.012131f
C32065 VDD.n11659 VSS 0.012131f
C32066 VDD.n11660 VSS 0.012131f
C32067 VDD.n11661 VSS 0.012131f
C32068 VDD.n11662 VSS 0.012131f
C32069 VDD.n11663 VSS 0.012131f
C32070 VDD.n11664 VSS 0.012131f
C32071 VDD.n11665 VSS 0.012131f
C32072 VDD.n11666 VSS 0.012131f
C32073 VDD.n11667 VSS 0.012131f
C32074 VDD.n11668 VSS 0.012131f
C32075 VDD.n11669 VSS 0.012131f
C32076 VDD.n11670 VSS 0.012131f
C32077 VDD.n11671 VSS 0.012131f
C32078 VDD.n11672 VSS 0.012131f
C32079 VDD.n11673 VSS 0.012131f
C32080 VDD.n11674 VSS 0.012131f
C32081 VDD.n11675 VSS 0.012131f
C32082 VDD.n11676 VSS 0.012131f
C32083 VDD.n11677 VSS 0.012131f
C32084 VDD.n11678 VSS 0.012131f
C32085 VDD.n11679 VSS 0.012131f
C32086 VDD.n11680 VSS 0.012131f
C32087 VDD.n11681 VSS 0.012131f
C32088 VDD.n11682 VSS 0.012131f
C32089 VDD.n11683 VSS 0.012131f
C32090 VDD.n11684 VSS 0.012131f
C32091 VDD.n11685 VSS 0.012131f
C32092 VDD.n11686 VSS 0.012131f
C32093 VDD.n11687 VSS 0.012131f
C32094 VDD.n11688 VSS 0.012131f
C32095 VDD.n11689 VSS 0.012131f
C32096 VDD.n11690 VSS 0.012131f
C32097 VDD.n11691 VSS 0.012131f
C32098 VDD.n11692 VSS 0.012131f
C32099 VDD.n11693 VSS 0.012131f
C32100 VDD.n11694 VSS 0.012131f
C32101 VDD.n11695 VSS 0.012131f
C32102 VDD.n11696 VSS 0.012131f
C32103 VDD.n11697 VSS 0.012131f
C32104 VDD.n11698 VSS 0.012131f
C32105 VDD.n11699 VSS 0.012131f
C32106 VDD.n11700 VSS 0.012131f
C32107 VDD.n11701 VSS 0.012131f
C32108 VDD.n11702 VSS 0.012131f
C32109 VDD.n11703 VSS 0.012131f
C32110 VDD.n11704 VSS 0.012131f
C32111 VDD.n11705 VSS 0.012131f
C32112 VDD.n11706 VSS 0.012131f
C32113 VDD.n11707 VSS 0.012131f
C32114 VDD.n11708 VSS 0.012131f
C32115 VDD.n11709 VSS 0.012131f
C32116 VDD.n11710 VSS 0.012131f
C32117 VDD.n11711 VSS 0.012131f
C32118 VDD.n11712 VSS 0.012131f
C32119 VDD.n11713 VSS 0.012131f
C32120 VDD.n11714 VSS 0.012131f
C32121 VDD.n11715 VSS 0.012131f
C32122 VDD.n11716 VSS 0.012131f
C32123 VDD.n11717 VSS 0.012131f
C32124 VDD.n11718 VSS 0.012131f
C32125 VDD.n11719 VSS 0.012131f
C32126 VDD.n11720 VSS 0.012131f
C32127 VDD.n11721 VSS 0.012131f
C32128 VDD.n11722 VSS 0.012131f
C32129 VDD.n11723 VSS 0.012131f
C32130 VDD.n11724 VSS 0.012131f
C32131 VDD.n11725 VSS 0.012131f
C32132 VDD.n11726 VSS 0.012131f
C32133 VDD.n11727 VSS 0.012131f
C32134 VDD.n11728 VSS 0.012131f
C32135 VDD.n11729 VSS 0.012131f
C32136 VDD.n11730 VSS 0.012131f
C32137 VDD.n11731 VSS 0.012131f
C32138 VDD.n11732 VSS 0.012131f
C32139 VDD.n11733 VSS 0.012131f
C32140 VDD.n11734 VSS 0.012131f
C32141 VDD.n11735 VSS 0.012131f
C32142 VDD.n11736 VSS 0.012131f
C32143 VDD.n11737 VSS 0.012131f
C32144 VDD.n11738 VSS 0.012131f
C32145 VDD.n11739 VSS 0.012131f
C32146 VDD.n11740 VSS 0.012131f
C32147 VDD.n11741 VSS 0.012131f
C32148 VDD.n11742 VSS 0.012131f
C32149 VDD.n11743 VSS 0.012131f
C32150 VDD.n11744 VSS 0.012131f
C32151 VDD.n11745 VSS 0.012131f
C32152 VDD.n11746 VSS 0.012131f
C32153 VDD.n11747 VSS 0.012131f
C32154 VDD.n11748 VSS 0.012131f
C32155 VDD.n11749 VSS 0.012131f
C32156 VDD.n11750 VSS 0.012131f
C32157 VDD.n11751 VSS 0.012131f
C32158 VDD.n11752 VSS 0.012131f
C32159 VDD.n11753 VSS 0.012131f
C32160 VDD.n11754 VSS 0.012131f
C32161 VDD.n11755 VSS 0.012131f
C32162 VDD.n11756 VSS 0.012131f
C32163 VDD.n11757 VSS 0.012131f
C32164 VDD.n11758 VSS 0.012131f
C32165 VDD.n11759 VSS 0.012131f
C32166 VDD.n11760 VSS 0.012131f
C32167 VDD.n11761 VSS 0.012131f
C32168 VDD.n11762 VSS 0.012131f
C32169 VDD.n11763 VSS 0.012131f
C32170 VDD.n11764 VSS 0.012131f
C32171 VDD.n11765 VSS 0.012131f
C32172 VDD.n11766 VSS 0.012131f
C32173 VDD.n11767 VSS 0.012131f
C32174 VDD.n11768 VSS 0.012131f
C32175 VDD.n11769 VSS 0.012131f
C32176 VDD.n11770 VSS 0.012131f
C32177 VDD.n11771 VSS 0.012131f
C32178 VDD.n11772 VSS 0.012131f
C32179 VDD.n11773 VSS 0.012131f
C32180 VDD.n11774 VSS 0.012131f
C32181 VDD.n11775 VSS 0.012131f
C32182 VDD.n11776 VSS 0.012131f
C32183 VDD.n11777 VSS 0.012131f
C32184 VDD.n11778 VSS 0.012131f
C32185 VDD.n11779 VSS 0.012131f
C32186 VDD.n11780 VSS 0.012131f
C32187 VDD.n11781 VSS 0.012131f
C32188 VDD.n11782 VSS 0.012131f
C32189 VDD.n11783 VSS 0.012131f
C32190 VDD.n11784 VSS 0.012131f
C32191 VDD.n11785 VSS 0.012131f
C32192 VDD.n11786 VSS 0.012131f
C32193 VDD.n11787 VSS 0.012131f
C32194 VDD.n11788 VSS 0.012131f
C32195 VDD.n11789 VSS 0.012131f
C32196 VDD.n11790 VSS 0.012131f
C32197 VDD.n11791 VSS 0.012131f
C32198 VDD.n11792 VSS 0.012131f
C32199 VDD.n11793 VSS 0.012131f
C32200 VDD.n11794 VSS 0.012131f
C32201 VDD.n11795 VSS 0.012131f
C32202 VDD.n11796 VSS 0.012131f
C32203 VDD.n11797 VSS 0.012131f
C32204 VDD.n11798 VSS 0.012131f
C32205 VDD.n11799 VSS 0.012131f
C32206 VDD.n11800 VSS 0.012131f
C32207 VDD.n11801 VSS 0.012131f
C32208 VDD.n11802 VSS 0.012131f
C32209 VDD.n11803 VSS 0.012131f
C32210 VDD.n11804 VSS 0.012131f
C32211 VDD.n11805 VSS 0.012131f
C32212 VDD.n11806 VSS 0.012131f
C32213 VDD.n11807 VSS 0.012131f
C32214 VDD.n11808 VSS 0.012131f
C32215 VDD.n11809 VSS 0.012131f
C32216 VDD.n11810 VSS 0.012131f
C32217 VDD.n11811 VSS 0.032438f
C32218 VDD.n11812 VSS 0.026728f
C32219 VDD.n11813 VSS 0.026728f
C32220 VDD.n11814 VSS 0.012131f
C32221 VDD.n11815 VSS 0.012131f
C32222 VDD.n11816 VSS 0.012131f
C32223 VDD.n11817 VSS 0.012131f
C32224 VDD.n11818 VSS 0.012131f
C32225 VDD.n11819 VSS 0.012131f
C32226 VDD.n11820 VSS 0.012131f
C32227 VDD.n11821 VSS 0.012131f
C32228 VDD.n11822 VSS 0.012131f
C32229 VDD.n11823 VSS 0.012131f
C32230 VDD.n11824 VSS 0.012131f
C32231 VDD.n11825 VSS 0.012131f
C32232 VDD.n11826 VSS 0.012131f
C32233 VDD.n11827 VSS 0.012131f
C32234 VDD.n11828 VSS 0.012131f
C32235 VDD.n11829 VSS 0.012131f
C32236 VDD.n11830 VSS 0.012131f
C32237 VDD.n11831 VSS 0.012131f
C32238 VDD.n11832 VSS 0.012131f
C32239 VDD.n11833 VSS 0.012131f
C32240 VDD.n11834 VSS 0.012131f
C32241 VDD.n11835 VSS 0.012131f
C32242 VDD.n11836 VSS 0.012131f
C32243 VDD.n11837 VSS 0.012131f
C32244 VDD.n11838 VSS 0.012131f
C32245 VDD.n11839 VSS 0.012131f
C32246 VDD.n11840 VSS 0.012131f
C32247 VDD.n11841 VSS 0.012131f
C32248 VDD.n11842 VSS 0.012131f
C32249 VDD.n11843 VSS 0.012131f
C32250 VDD.n11844 VSS 0.012131f
C32251 VDD.n11845 VSS 0.012131f
C32252 VDD.n11846 VSS 0.012131f
C32253 VDD.n11847 VSS 0.012131f
C32254 VDD.n11848 VSS 0.012131f
C32255 VDD.n11849 VSS 0.012131f
C32256 VDD.n11850 VSS 0.012131f
C32257 VDD.n11851 VSS 0.012131f
C32258 VDD.n11852 VSS 0.012131f
C32259 VDD.n11853 VSS 0.012131f
C32260 VDD.n11854 VSS 0.012131f
C32261 VDD.n11855 VSS 0.012131f
C32262 VDD.n11856 VSS 0.012131f
C32263 VDD.n11857 VSS 0.012131f
C32264 VDD.n11858 VSS 0.012131f
C32265 VDD.n11859 VSS 0.012131f
C32266 VDD.n11860 VSS 0.012131f
C32267 VDD.n11861 VSS 0.012131f
C32268 VDD.n11862 VSS 0.012131f
C32269 VDD.n11863 VSS 0.012131f
C32270 VDD.n11864 VSS 0.012131f
C32271 VDD.n11865 VSS 0.012131f
C32272 VDD.n11866 VSS 0.012131f
C32273 VDD.n11867 VSS 0.012131f
C32274 VDD.n11868 VSS 0.012131f
C32275 VDD.n11869 VSS 0.012131f
C32276 VDD.n11870 VSS 0.012131f
C32277 VDD.n11871 VSS 0.012131f
C32278 VDD.n11872 VSS 0.159151f
C32279 VDD.n11873 VSS 0.010242f
C32280 VDD.n11874 VSS 0.012131f
C32281 VDD.n11875 VSS 0.012131f
C32282 VDD.n11876 VSS 0.012131f
C32283 VDD.n11877 VSS 0.012131f
C32284 VDD.n11878 VSS 0.012131f
C32285 VDD.n11879 VSS 0.012131f
C32286 VDD.n11880 VSS 0.012131f
C32287 VDD.n11881 VSS 0.012131f
C32288 VDD.n11882 VSS 0.012131f
C32289 VDD.n11883 VSS 0.012131f
C32290 VDD.n11884 VSS 0.012131f
C32291 VDD.n11885 VSS 0.012131f
C32292 VDD.n11886 VSS 0.012131f
C32293 VDD.n11887 VSS 0.012131f
C32294 VDD.n11888 VSS 0.012131f
C32295 VDD.n11889 VSS 0.012131f
C32296 VDD.n11890 VSS 0.012131f
C32297 VDD.n11891 VSS 0.012131f
C32298 VDD.n11892 VSS 0.012131f
C32299 VDD.n11893 VSS 0.012131f
C32300 VDD.n11894 VSS 0.012131f
C32301 VDD.n11895 VSS 0.012131f
C32302 VDD.n11896 VSS 0.012131f
C32303 VDD.n11897 VSS 0.012131f
C32304 VDD.n11898 VSS 0.012131f
C32305 VDD.n11899 VSS 0.012131f
C32306 VDD.n11900 VSS 0.012131f
C32307 VDD.n11901 VSS 0.012131f
C32308 VDD.n11902 VSS 0.012131f
C32309 VDD.n11903 VSS 0.012131f
C32310 VDD.n11904 VSS 0.012131f
C32311 VDD.n11905 VSS 0.012131f
C32312 VDD.n11906 VSS 0.012131f
C32313 VDD.n11907 VSS 0.012131f
C32314 VDD.n11908 VSS 0.012131f
C32315 VDD.n11909 VSS 0.012131f
C32316 VDD.n11910 VSS 0.012131f
C32317 VDD.n11911 VSS 0.012131f
C32318 VDD.n11912 VSS 0.012131f
C32319 VDD.n11913 VSS 0.012131f
C32320 VDD.n11914 VSS 0.012131f
C32321 VDD.n11915 VSS 0.012131f
C32322 VDD.n11916 VSS 0.012131f
C32323 VDD.n11917 VSS 0.012131f
C32324 VDD.n11918 VSS 0.012131f
C32325 VDD.n11919 VSS 0.012131f
C32326 VDD.n11920 VSS 0.012131f
C32327 VDD.n11921 VSS 0.012131f
C32328 VDD.n11922 VSS 0.012131f
C32329 VDD.n11923 VSS 0.012131f
C32330 VDD.n11924 VSS 0.012131f
C32331 VDD.n11925 VSS 0.012131f
C32332 VDD.n11926 VSS 0.012131f
C32333 VDD.n11927 VSS 0.012131f
C32334 VDD.n11928 VSS 0.012131f
C32335 VDD.n11929 VSS 0.012131f
C32336 VDD.n11930 VSS 0.012131f
C32337 VDD.n11931 VSS 0.012131f
C32338 VDD.n11932 VSS 0.012131f
C32339 VDD.n11933 VSS 0.012131f
C32340 VDD.n11934 VSS 0.012131f
C32341 VDD.n11935 VSS 0.012131f
C32342 VDD.n11936 VSS 0.012131f
C32343 VDD.n11937 VSS 0.012131f
C32344 VDD.n11938 VSS 0.012131f
C32345 VDD.n11939 VSS 0.012131f
C32346 VDD.n11940 VSS 0.012131f
C32347 VDD.n11941 VSS 0.012131f
C32348 VDD.n11942 VSS 0.012131f
C32349 VDD.n11943 VSS 0.012131f
C32350 VDD.n11944 VSS 0.012131f
C32351 VDD.n11945 VSS 0.012131f
C32352 VDD.n11946 VSS 0.012131f
C32353 VDD.n11947 VSS 0.012131f
C32354 VDD.n11948 VSS 0.012131f
C32355 VDD.n11949 VSS 0.012131f
C32356 VDD.n11950 VSS 0.012131f
C32357 VDD.n11951 VSS 0.012131f
C32358 VDD.n11952 VSS 0.012131f
C32359 VDD.n11953 VSS 0.012131f
C32360 VDD.n11954 VSS 0.012131f
C32361 VDD.n11955 VSS 0.012131f
C32362 VDD.n11956 VSS 0.012131f
C32363 VDD.n11957 VSS 0.012131f
C32364 VDD.n11958 VSS 0.012131f
C32365 VDD.n11959 VSS 0.012131f
C32366 VDD.n11960 VSS 0.012131f
C32367 VDD.n11961 VSS 0.012131f
C32368 VDD.n11962 VSS 0.012131f
C32369 VDD.n11963 VSS 0.012131f
C32370 VDD.n11964 VSS 0.012131f
C32371 VDD.n11965 VSS 0.012131f
C32372 VDD.n11966 VSS 0.012131f
C32373 VDD.n11967 VSS 0.012131f
C32374 VDD.n11968 VSS 0.012131f
C32375 VDD.n11969 VSS 0.012131f
C32376 VDD.n11970 VSS 0.012131f
C32377 VDD.n11971 VSS 0.012131f
C32378 VDD.n11972 VSS 0.012131f
C32379 VDD.n11973 VSS 0.012131f
C32380 VDD.n11974 VSS 0.012131f
C32381 VDD.n11975 VSS 0.012131f
C32382 VDD.n11976 VSS 0.012131f
C32383 VDD.n11977 VSS 0.012131f
C32384 VDD.n11978 VSS 0.012131f
C32385 VDD.n11979 VSS 0.012131f
C32386 VDD.n11980 VSS 0.012131f
C32387 VDD.n11981 VSS 0.012131f
C32388 VDD.n11982 VSS 0.012131f
C32389 VDD.n11983 VSS 0.012131f
C32390 VDD.n11984 VSS 0.012131f
C32391 VDD.n11985 VSS 0.012131f
C32392 VDD.n11986 VSS 0.012131f
C32393 VDD.n11987 VSS 0.012131f
C32394 VDD.n11988 VSS 0.012131f
C32395 VDD.n11989 VSS 0.012131f
C32396 VDD.n11990 VSS 0.012131f
C32397 VDD.n11991 VSS 0.012131f
C32398 VDD.n11992 VSS 0.012131f
C32399 VDD.n11993 VSS 0.012131f
C32400 VDD.n11994 VSS 0.012131f
C32401 VDD.n11995 VSS 0.012131f
C32402 VDD.n11996 VSS 0.012131f
C32403 VDD.n11997 VSS 0.012131f
C32404 VDD.n11998 VSS 0.012131f
C32405 VDD.n11999 VSS 0.012131f
C32406 VDD.n12000 VSS 0.012131f
C32407 VDD.n12001 VSS 0.012131f
C32408 VDD.n12002 VSS 0.012131f
C32409 VDD.n12003 VSS 0.012131f
C32410 VDD.n12004 VSS 0.012131f
C32411 VDD.n12005 VSS 0.012131f
C32412 VDD.n12006 VSS 0.012131f
C32413 VDD.n12007 VSS 0.012131f
C32414 VDD.n12008 VSS 0.012131f
C32415 VDD.n12009 VSS 0.012131f
C32416 VDD.n12010 VSS 0.012131f
C32417 VDD.n12011 VSS 0.012131f
C32418 VDD.n12012 VSS 0.012131f
C32419 VDD.n12013 VSS 0.012131f
C32420 VDD.n12014 VSS 0.012131f
C32421 VDD.n12015 VSS 0.012131f
C32422 VDD.n12016 VSS 0.012131f
C32423 VDD.n12017 VSS 0.012131f
C32424 VDD.n12018 VSS 0.012131f
C32425 VDD.n12019 VSS 0.012131f
C32426 VDD.n12020 VSS 0.012131f
C32427 VDD.n12021 VSS 0.012131f
C32428 VDD.n12022 VSS 0.012131f
C32429 VDD.n12023 VSS 0.012131f
C32430 VDD.n12024 VSS 0.012131f
C32431 VDD.n12025 VSS 0.012131f
C32432 VDD.n12026 VSS 0.012131f
C32433 VDD.n12027 VSS 0.012131f
C32434 VDD.n12028 VSS 0.012131f
C32435 VDD.n12029 VSS 0.012131f
C32436 VDD.n12030 VSS 0.012131f
C32437 VDD.n12031 VSS 0.012131f
C32438 VDD.n12032 VSS 0.012131f
C32439 VDD.n12033 VSS 0.012131f
C32440 VDD.n12034 VSS 0.012131f
C32441 VDD.n12035 VSS 0.012131f
C32442 VDD.n12036 VSS 0.012131f
C32443 VDD.n12037 VSS 0.012131f
C32444 VDD.n12038 VSS 0.012131f
C32445 VDD.n12039 VSS 0.012131f
C32446 VDD.n12040 VSS 0.012131f
C32447 VDD.n12041 VSS 0.012131f
C32448 VDD.n12042 VSS 0.012131f
C32449 VDD.n12043 VSS 0.012131f
C32450 VDD.n12044 VSS 0.012131f
C32451 VDD.n12045 VSS 0.012131f
C32452 VDD.n12046 VSS 0.012131f
C32453 VDD.n12047 VSS 0.012131f
C32454 VDD.n12048 VSS 0.012131f
C32455 VDD.n12049 VSS 0.012131f
C32456 VDD.n12050 VSS 0.012131f
C32457 VDD.n12051 VSS 0.012131f
C32458 VDD.n12052 VSS 0.012131f
C32459 VDD.n12053 VSS 0.012131f
C32460 VDD.n12054 VSS 0.012131f
C32461 VDD.n12055 VSS 0.012131f
C32462 VDD.n12056 VSS 0.012131f
C32463 VDD.n12057 VSS 0.012131f
C32464 VDD.n12058 VSS 0.012131f
C32465 VDD.n12059 VSS 0.012131f
C32466 VDD.n12060 VSS 0.012131f
C32467 VDD.n12061 VSS 0.012131f
C32468 VDD.n12062 VSS 0.012131f
C32469 VDD.n12063 VSS 0.012131f
C32470 VDD.n12064 VSS 0.012131f
C32471 VDD.n12065 VSS 0.012131f
C32472 VDD.n12066 VSS 0.012131f
C32473 VDD.n12067 VSS 0.012131f
C32474 VDD.n12068 VSS 0.012131f
C32475 VDD.n12069 VSS 0.012131f
C32476 VDD.n12070 VSS 0.012131f
C32477 VDD.n12071 VSS 0.012131f
C32478 VDD.n12072 VSS 0.012131f
C32479 VDD.n12073 VSS 0.012131f
C32480 VDD.n12074 VSS 0.012131f
C32481 VDD.n12075 VSS 0.012131f
C32482 VDD.n12076 VSS 0.012131f
C32483 VDD.n12077 VSS 0.012131f
C32484 VDD.n12078 VSS 0.012131f
C32485 VDD.n12079 VSS 0.012131f
C32486 VDD.n12080 VSS 0.012131f
C32487 VDD.n12081 VSS 0.012131f
C32488 VDD.n12082 VSS 0.012131f
C32489 VDD.n12083 VSS 0.012131f
C32490 VDD.n12084 VSS 0.012131f
C32491 VDD.n12085 VSS 0.012131f
C32492 VDD.n12086 VSS 0.012131f
C32493 VDD.n12087 VSS 0.012131f
C32494 VDD.n12088 VSS 0.012131f
C32495 VDD.n12089 VSS 0.012131f
C32496 VDD.n12090 VSS 0.012131f
C32497 VDD.n12091 VSS 0.012131f
C32498 VDD.n12092 VSS 0.012131f
C32499 VDD.n12093 VSS 0.012131f
C32500 VDD.n12094 VSS 0.012131f
C32501 VDD.n12095 VSS 0.012131f
C32502 VDD.n12096 VSS 0.012131f
C32503 VDD.n12097 VSS 0.012131f
C32504 VDD.n12098 VSS 0.012131f
C32505 VDD.n12099 VSS 0.012131f
C32506 VDD.n12100 VSS 0.012131f
C32507 VDD.n12101 VSS 0.012131f
C32508 VDD.n12102 VSS 0.012131f
C32509 VDD.n12103 VSS 0.012131f
C32510 VDD.n12104 VSS 0.012131f
C32511 VDD.n12105 VSS 0.012131f
C32512 VDD.n12106 VSS 0.012131f
C32513 VDD.n12107 VSS 0.012131f
C32514 VDD.n12108 VSS 0.012131f
C32515 VDD.n12109 VSS 0.012131f
C32516 VDD.n12110 VSS 0.012131f
C32517 VDD.n12111 VSS 0.012131f
C32518 VDD.n12112 VSS 0.012131f
C32519 VDD.n12113 VSS 0.012131f
C32520 VDD.n12114 VSS 0.012131f
C32521 VDD.n12115 VSS 0.012131f
C32522 VDD.n12116 VSS 0.012131f
C32523 VDD.n12117 VSS 0.012131f
C32524 VDD.n12118 VSS 0.012131f
C32525 VDD.n12119 VSS 0.012131f
C32526 VDD.n12120 VSS 0.012131f
C32527 VDD.n12121 VSS 0.012131f
C32528 VDD.n12122 VSS 0.012131f
C32529 VDD.n12123 VSS 0.012131f
C32530 VDD.n12124 VSS 0.012131f
C32531 VDD.n12125 VSS 0.012131f
C32532 VDD.n12126 VSS 0.012131f
C32533 VDD.n12127 VSS 0.012131f
C32534 VDD.n12128 VSS 0.012131f
C32535 VDD.n12129 VSS 0.012131f
C32536 VDD.n12130 VSS 0.012131f
C32537 VDD.n12131 VSS 0.012131f
C32538 VDD.n12132 VSS 0.012131f
C32539 VDD.n12133 VSS 0.012131f
C32540 VDD.n12134 VSS 0.012131f
C32541 VDD.n12135 VSS 0.012131f
C32542 VDD.n12136 VSS 0.012131f
C32543 VDD.n12137 VSS 0.012131f
C32544 VDD.n12138 VSS 0.012131f
C32545 VDD.n12139 VSS 0.012131f
C32546 VDD.n12140 VSS 0.012131f
C32547 VDD.n12141 VSS 0.012131f
C32548 VDD.n12142 VSS 0.012131f
C32549 VDD.n12143 VSS 0.012131f
C32550 VDD.n12144 VSS 0.012131f
C32551 VDD.n12145 VSS 0.012131f
C32552 VDD.n12146 VSS 0.012131f
C32553 VDD.n12147 VSS 0.012131f
C32554 VDD.n12148 VSS 0.012131f
C32555 VDD.n12149 VSS 0.012131f
C32556 VDD.n12150 VSS 0.012131f
C32557 VDD.n12151 VSS 0.012131f
C32558 VDD.n12152 VSS 0.012131f
C32559 VDD.n12153 VSS 0.012131f
C32560 VDD.n12154 VSS 0.012131f
C32561 VDD.n12155 VSS 0.012131f
C32562 VDD.n12156 VSS 0.012131f
C32563 VDD.n12157 VSS 0.012131f
C32564 VDD.n12158 VSS 0.012131f
C32565 VDD.n12159 VSS 0.012131f
C32566 VDD.n12160 VSS 0.012131f
C32567 VDD.n12161 VSS 0.012131f
C32568 VDD.n12162 VSS 0.012131f
C32569 VDD.n12163 VSS 0.012131f
C32570 VDD.n12164 VSS 0.012131f
C32571 VDD.n12165 VSS 0.012131f
C32572 VDD.n12166 VSS 0.012131f
C32573 VDD.n12167 VSS 0.012131f
C32574 VDD.n12168 VSS 0.012131f
C32575 VDD.n12169 VSS 0.012131f
C32576 VDD.n12170 VSS 0.012131f
C32577 VDD.n12171 VSS 0.012131f
C32578 VDD.n12172 VSS 0.012131f
C32579 VDD.n12173 VSS 0.012131f
C32580 VDD.n12174 VSS 0.012131f
C32581 VDD.n12175 VSS 0.012131f
C32582 VDD.n12176 VSS 0.012131f
C32583 VDD.n12177 VSS 0.012131f
C32584 VDD.n12178 VSS 0.012131f
C32585 VDD.n12179 VSS 0.012131f
C32586 VDD.n12180 VSS 0.012131f
C32587 VDD.n12181 VSS 0.012131f
C32588 VDD.n12182 VSS 0.012131f
C32589 VDD.n12183 VSS 0.012131f
C32590 VDD.n12184 VSS 0.012131f
C32591 VDD.n12185 VSS 0.012131f
C32592 VDD.n12186 VSS 0.012131f
C32593 VDD.n12187 VSS 0.012131f
C32594 VDD.n12188 VSS 0.012131f
C32595 VDD.n12189 VSS 0.012131f
C32596 VDD.n12190 VSS 0.012131f
C32597 VDD.n12191 VSS 0.012131f
C32598 VDD.n12192 VSS 0.012131f
C32599 VDD.n12193 VSS 0.012131f
C32600 VDD.n12194 VSS 0.012131f
C32601 VDD.n12195 VSS 0.012131f
C32602 VDD.n12196 VSS 0.012131f
C32603 VDD.n12197 VSS 0.012131f
C32604 VDD.n12198 VSS 0.012131f
C32605 VDD.n12199 VSS 0.012131f
C32606 VDD.n12200 VSS 0.012131f
C32607 VDD.n12201 VSS 0.012131f
C32608 VDD.n12202 VSS 0.012131f
C32609 VDD.n12203 VSS 0.012131f
C32610 VDD.n12204 VSS 0.012131f
C32611 VDD.n12205 VSS 0.012131f
C32612 VDD.n12206 VSS 0.012131f
C32613 VDD.n12207 VSS 0.012131f
C32614 VDD.n12208 VSS 0.012131f
C32615 VDD.n12209 VSS 0.012131f
C32616 VDD.n12210 VSS 0.012131f
C32617 VDD.n12211 VSS 0.012131f
C32618 VDD.n12212 VSS 0.012131f
C32619 VDD.n12213 VSS 0.012131f
C32620 VDD.n12214 VSS 0.012131f
C32621 VDD.n12215 VSS 0.012131f
C32622 VDD.n12216 VSS 0.012131f
C32623 VDD.n12217 VSS 0.012131f
C32624 VDD.n12218 VSS 0.012131f
C32625 VDD.n12219 VSS 0.012131f
C32626 VDD.n12220 VSS 0.012131f
C32627 VDD.n12221 VSS 0.012131f
C32628 VDD.n12222 VSS 0.012131f
C32629 VDD.n12223 VSS 0.012131f
C32630 VDD.n12224 VSS 0.012131f
C32631 VDD.n12225 VSS 0.012131f
C32632 VDD.n12226 VSS 0.012131f
C32633 VDD.n12227 VSS 0.012131f
C32634 VDD.n12228 VSS 0.012131f
C32635 VDD.n12229 VSS 0.012131f
C32636 VDD.n12230 VSS 0.012131f
C32637 VDD.n12231 VSS 0.012131f
C32638 VDD.n12232 VSS 0.012131f
C32639 VDD.n12233 VSS 0.012131f
C32640 VDD.n12234 VSS 0.012131f
C32641 VDD.n12235 VSS 0.012131f
C32642 VDD.n12236 VSS 0.012131f
C32643 VDD.n12237 VSS 0.012131f
C32644 VDD.n12238 VSS 0.012131f
C32645 VDD.n12239 VSS 0.012131f
C32646 VDD.n12240 VSS 0.012131f
C32647 VDD.n12241 VSS 0.012131f
C32648 VDD.n12242 VSS 0.012131f
C32649 VDD.n12243 VSS 0.012131f
C32650 VDD.n12244 VSS 0.012131f
C32651 VDD.n12245 VSS 0.012131f
C32652 VDD.n12246 VSS 0.012131f
C32653 VDD.n12247 VSS 0.012131f
C32654 VDD.n12248 VSS 0.012131f
C32655 VDD.n12249 VSS 0.012131f
C32656 VDD.n12250 VSS 0.012131f
C32657 VDD.n12251 VSS 0.012131f
C32658 VDD.n12252 VSS 0.012131f
C32659 VDD.n12253 VSS 0.012131f
C32660 VDD.n12254 VSS 0.012131f
C32661 VDD.n12255 VSS 0.012131f
C32662 VDD.n12256 VSS 0.012131f
C32663 VDD.n12257 VSS 0.012131f
C32664 VDD.n12258 VSS 0.012131f
C32665 VDD.n12259 VSS 0.012131f
C32666 VDD.n12260 VSS 0.012131f
C32667 VDD.n12261 VSS 0.012131f
C32668 VDD.n12262 VSS 0.012131f
C32669 VDD.n12263 VSS 0.012131f
C32670 VDD.n12264 VSS 0.012131f
C32671 VDD.n12265 VSS 0.012131f
C32672 VDD.n12266 VSS 0.012131f
C32673 VDD.n12267 VSS 0.012131f
C32674 VDD.n12268 VSS 0.012131f
C32675 VDD.n12269 VSS 0.012131f
C32676 VDD.n12270 VSS 0.012131f
C32677 VDD.n12271 VSS 0.012131f
C32678 VDD.n12272 VSS 0.012131f
C32679 VDD.n12273 VSS 0.012131f
C32680 VDD.n12274 VSS 0.012131f
C32681 VDD.n12275 VSS 0.012131f
C32682 VDD.n12276 VSS 0.012131f
C32683 VDD.n12277 VSS 0.012131f
C32684 VDD.n12278 VSS 0.012131f
C32685 VDD.n12279 VSS 0.012131f
C32686 VDD.n12280 VSS 0.012131f
C32687 VDD.n12281 VSS 0.012131f
C32688 VDD.n12282 VSS 0.012131f
C32689 VDD.n12283 VSS 0.012131f
C32690 VDD.n12284 VSS 0.012131f
C32691 VDD.n12285 VSS 0.012131f
C32692 VDD.n12286 VSS 0.012131f
C32693 VDD.n12287 VSS 0.012131f
C32694 VDD.n12288 VSS 0.012131f
C32695 VDD.n12289 VSS 0.012131f
C32696 VDD.n12290 VSS 0.012131f
C32697 VDD.n12291 VSS 0.012131f
C32698 VDD.n12292 VSS 0.012131f
C32699 VDD.n12293 VSS 0.012131f
C32700 VDD.n12294 VSS 0.012131f
C32701 VDD.n12295 VSS 0.012131f
C32702 VDD.n12296 VSS 0.012131f
C32703 VDD.n12297 VSS 0.012131f
C32704 VDD.n12298 VSS 0.012131f
C32705 VDD.n12299 VSS 0.012131f
C32706 VDD.n12300 VSS 0.012131f
C32707 VDD.n12301 VSS 0.012131f
C32708 VDD.n12302 VSS 0.012131f
C32709 VDD.n12303 VSS 0.012131f
C32710 VDD.n12304 VSS 0.012131f
C32711 VDD.n12305 VSS 0.012131f
C32712 VDD.n12306 VSS 0.012131f
C32713 VDD.n12307 VSS 0.012131f
C32714 VDD.n12308 VSS 0.012131f
C32715 VDD.n12309 VSS 0.012131f
C32716 VDD.n12310 VSS 0.012131f
C32717 VDD.n12311 VSS 0.012131f
C32718 VDD.n12312 VSS 0.012131f
C32719 VDD.n12313 VSS 0.012131f
C32720 VDD.n12314 VSS 0.012131f
C32721 VDD.n12315 VSS 0.012131f
C32722 VDD.n12316 VSS 0.012131f
C32723 VDD.n12317 VSS 0.012131f
C32724 VDD.n12318 VSS 0.012131f
C32725 VDD.n12319 VSS 0.012131f
C32726 VDD.n12320 VSS 0.012131f
C32727 VDD.n12321 VSS 0.012131f
C32728 VDD.n12322 VSS 0.012131f
C32729 VDD.n12323 VSS 0.012131f
C32730 VDD.n12324 VSS 0.012131f
C32731 VDD.n12325 VSS 0.012131f
C32732 VDD.n12326 VSS 0.012131f
C32733 VDD.n12327 VSS 0.012131f
C32734 VDD.n12328 VSS 0.012131f
C32735 VDD.n12329 VSS 0.012131f
C32736 VDD.n12330 VSS 0.012131f
C32737 VDD.n12331 VSS 0.012131f
C32738 VDD.n12332 VSS 0.012131f
C32739 VDD.n12333 VSS 0.012131f
C32740 VDD.n12334 VSS 0.012131f
C32741 VDD.n12335 VSS 0.012131f
C32742 VDD.n12336 VSS 0.012131f
C32743 VDD.n12337 VSS 0.012131f
C32744 VDD.n12338 VSS 0.012131f
C32745 VDD.n12339 VSS 0.012131f
C32746 VDD.n12340 VSS 0.012131f
C32747 VDD.n12341 VSS 0.012131f
C32748 VDD.n12342 VSS 0.012131f
C32749 VDD.n12343 VSS 0.012131f
C32750 VDD.n12344 VSS 0.012131f
C32751 VDD.n12345 VSS 0.012131f
C32752 VDD.n12346 VSS 0.012131f
C32753 VDD.n12347 VSS 0.012131f
C32754 VDD.n12348 VSS 0.012131f
C32755 VDD.n12349 VSS 0.012131f
C32756 VDD.n12350 VSS 0.012131f
C32757 VDD.n12351 VSS 0.012131f
C32758 VDD.n12352 VSS 0.012131f
C32759 VDD.n12353 VSS 0.012131f
C32760 VDD.n12354 VSS 0.012131f
C32761 VDD.n12355 VSS 0.012131f
C32762 VDD.n12356 VSS 0.012131f
C32763 VDD.n12357 VSS 0.012131f
C32764 VDD.n12358 VSS 0.012131f
C32765 VDD.n12359 VSS 0.012131f
C32766 VDD.n12360 VSS 0.012131f
C32767 VDD.n12361 VSS 0.012131f
C32768 VDD.n12362 VSS 0.012131f
C32769 VDD.n12363 VSS 0.012131f
C32770 VDD.n12364 VSS 0.012131f
C32771 VDD.n12365 VSS 0.012131f
C32772 VDD.n12366 VSS 0.012131f
C32773 VDD.n12367 VSS 0.012131f
C32774 VDD.n12368 VSS 0.012131f
C32775 VDD.n12369 VSS 0.012131f
C32776 VDD.n12370 VSS 0.012131f
C32777 VDD.n12371 VSS 0.012131f
C32778 VDD.n12372 VSS 0.012131f
C32779 VDD.n12373 VSS 0.012131f
C32780 VDD.n12374 VSS 0.012131f
C32781 VDD.n12375 VSS 0.012131f
C32782 VDD.n12376 VSS 0.012131f
C32783 VDD.n12377 VSS 0.012131f
C32784 VDD.n12378 VSS 0.012131f
C32785 VDD.n12379 VSS 0.012131f
C32786 VDD.n12380 VSS 0.012131f
C32787 VDD.n12381 VSS 0.012131f
C32788 VDD.n12382 VSS 0.012131f
C32789 VDD.n12383 VSS 0.012131f
C32790 VDD.n12384 VSS 0.012131f
C32791 VDD.n12385 VSS 0.012131f
C32792 VDD.n12386 VSS 0.012131f
C32793 VDD.n12387 VSS 0.012131f
C32794 VDD.n12388 VSS 0.012131f
C32795 VDD.n12389 VSS 0.012131f
C32796 VDD.n12390 VSS 0.012131f
C32797 VDD.n12391 VSS 0.012131f
C32798 VDD.n12392 VSS 0.012131f
C32799 VDD.n12393 VSS 0.012131f
C32800 VDD.n12394 VSS 0.012131f
C32801 VDD.n12395 VSS 0.012131f
C32802 VDD.n12396 VSS 0.012131f
C32803 VDD.n12397 VSS 0.012131f
C32804 VDD.n12398 VSS 0.012131f
C32805 VDD.n12399 VSS 0.012131f
C32806 VDD.n12400 VSS 0.012131f
C32807 VDD.n12401 VSS 0.012131f
C32808 VDD.n12402 VSS 0.012131f
C32809 VDD.n12403 VSS 0.012131f
C32810 VDD.n12404 VSS 0.012131f
C32811 VDD.n12405 VSS 0.012131f
C32812 VDD.n12406 VSS 0.012131f
C32813 VDD.n12407 VSS 0.012131f
C32814 VDD.n12408 VSS 0.012131f
C32815 VDD.n12409 VSS 0.012131f
C32816 VDD.n12410 VSS 0.012131f
C32817 VDD.n12411 VSS 0.012131f
C32818 VDD.n12412 VSS 0.012131f
C32819 VDD.n12413 VSS 0.012131f
C32820 VDD.n12414 VSS 0.012131f
C32821 VDD.n12415 VSS 0.012131f
C32822 VDD.n12416 VSS 0.012131f
C32823 VDD.n12417 VSS 0.012131f
C32824 VDD.n12418 VSS 0.012131f
C32825 VDD.n12419 VSS 0.012131f
C32826 VDD.n12420 VSS 0.012131f
C32827 VDD.n12421 VSS 0.012131f
C32828 VDD.n12422 VSS 0.012131f
C32829 VDD.n12423 VSS 0.012131f
C32830 VDD.n12424 VSS 0.012131f
C32831 VDD.n12425 VSS 0.012131f
C32832 VDD.n12426 VSS 0.012131f
C32833 VDD.n12427 VSS 0.012131f
C32834 VDD.n12428 VSS 0.012131f
C32835 VDD.n12429 VSS 0.012131f
C32836 VDD.n12430 VSS 0.012131f
C32837 VDD.n12431 VSS 0.012131f
C32838 VDD.n12432 VSS 0.012131f
C32839 VDD.n12433 VSS 0.012131f
C32840 VDD.n12434 VSS 0.012131f
C32841 VDD.n12435 VSS 0.012131f
C32842 VDD.n12436 VSS 0.012131f
C32843 VDD.n12437 VSS 0.012131f
C32844 VDD.n12438 VSS 0.012131f
C32845 VDD.n12439 VSS 0.012131f
C32846 VDD.n12440 VSS 0.00864f
C32847 VDD.n12441 VSS 0.012131f
C32848 VDD.n12442 VSS 0.012131f
C32849 VDD.n12443 VSS 0.012131f
C32850 VDD.n12444 VSS 0.006065f
C32851 VDD.n12445 VSS 0.037495f
C32852 VDD.n12446 VSS 0.006065f
C32853 VDD.n12447 VSS 0.012131f
C32854 VDD.n12448 VSS 0.29741f
C32855 VDD.n12449 VSS 0.825781f
C32856 VDD.t2005 VSS 0.028519f
C32857 VDD.t827 VSS 0.028519f
C32858 VDD.n12450 VSS 0.009191f
C32859 VDD.n12451 VSS 0.261039f
C32860 VDD.t825 VSS 0.066856f
C32861 VDD.t2456 VSS 0.066856f
C32862 VDD.n12452 VSS 0.709674f
C32863 VDD.t4535 VSS 0.028519f
C32864 VDD.t3386 VSS 0.028519f
C32865 VDD.n12453 VSS 0.009191f
C32866 VDD.n12454 VSS 0.644755f
C32867 VDD.t3385 VSS 0.066856f
C32868 VDD.t794 VSS 0.066856f
C32869 VDD.n12455 VSS 0.690489f
C32870 VDD.t3076 VSS 0.066856f
C32871 VDD.t4532 VSS 0.066856f
C32872 VDD.n12456 VSS 0.690489f
C32873 VDD.t4217 VSS 0.028519f
C32874 VDD.t3077 VSS 0.028519f
C32875 VDD.n12457 VSS 0.009191f
C32876 VDD.n12458 VSS 0.523473f
C32877 VDD.n12459 VSS 0.524869f
C32878 VDD.n12460 VSS 0.208534f
C32879 VDD.n12461 VSS 0.865258f
C32880 VDD.n12462 VSS 0.865258f
C32881 VDD.t826 VSS 1.45794f
C32882 VDD.t614 VSS 1.96535f
C32883 VDD.t2347 VSS 1.96535f
C32884 VDD.t2046 VSS 1.31955f
C32885 VDD.n12463 VSS 0.595476f
C32886 VDD.n12464 VSS 0.645798f
C32887 VDD.n12465 VSS 0.206947f
C32888 VDD.n12466 VSS 0.208534f
C32889 VDD.n12467 VSS 0.529799f
C32890 VDD.n12468 VSS 0.207221f
C32891 VDD.n12469 VSS 0.902999f
C32892 VDD.t2079 VSS 1.45794f
C32893 VDD.t1823 VSS 1.96535f
C32894 VDD.t2731 VSS 1.96535f
C32895 VDD.t1852 VSS 1.31955f
C32896 VDD.n12470 VSS 0.595476f
C32897 VDD.n12471 VSS 0.645798f
C32898 VDD.t1710 VSS 1.36988f
C32899 VDD.t1489 VSS 1.96535f
C32900 VDD.t728 VSS 1.96535f
C32901 VDD.t1508 VSS 1.45794f
C32902 VDD.n12472 VSS 0.865258f
C32903 VDD.n12473 VSS 0.208534f
C32904 VDD.n12474 VSS 0.524869f
C32905 VDD.t1893 VSS 0.028519f
C32906 VDD.t4485 VSS 0.028519f
C32907 VDD.n12475 VSS 0.009191f
C32908 VDD.t4575 VSS 0.028519f
C32909 VDD.t655 VSS 0.028519f
C32910 VDD.n12476 VSS 0.009191f
C32911 VDD.n12477 VSS 0.523473f
C32912 VDD.t1892 VSS 0.066856f
C32913 VDD.t4574 VSS 0.066856f
C32914 VDD.t654 VSS 0.066856f
C32915 VDD.t4484 VSS 0.066856f
C32916 VDD.n12478 VSS 0.690489f
C32917 VDD.t2349 VSS 0.066856f
C32918 VDD.t830 VSS 0.066856f
C32919 VDD.t1038 VSS 0.066856f
C32920 VDD.t727 VSS 0.066856f
C32921 VDD.n12479 VSS 0.690489f
C32922 VDD.t2350 VSS 0.028519f
C32923 VDD.t729 VSS 0.028519f
C32924 VDD.n12480 VSS 0.009191f
C32925 VDD.t832 VSS 0.028519f
C32926 VDD.t1039 VSS 0.028519f
C32927 VDD.n12481 VSS 0.009191f
C32928 VDD.n12482 VSS 0.644755f
C32929 VDD.t3878 VSS 0.066856f
C32930 VDD.t2498 VSS 0.066856f
C32931 VDD.t2714 VSS 0.066856f
C32932 VDD.t2387 VSS 0.066856f
C32933 VDD.n12483 VSS 0.709674f
C32934 VDD.t3879 VSS 0.028519f
C32935 VDD.t2388 VSS 0.028519f
C32936 VDD.n12484 VSS 0.009191f
C32937 VDD.t2499 VSS 0.028519f
C32938 VDD.t2715 VSS 0.028519f
C32939 VDD.n12485 VSS 0.009191f
C32940 VDD.n12486 VSS 0.261039f
C32941 VDD.n12487 VSS 0.62132f
C32942 VDD.n12488 VSS 0.099723f
C32943 VDD.t905 VSS 0.066856f
C32944 VDD.n12489 VSS 0.125227f
C32945 VDD.n12490 VSS 0.101294f
C32946 VDD.n12491 VSS 0.016021f
C32947 VDD.t2525 VSS 0.025104f
C32948 VDD.n12492 VSS 0.083673f
C32949 VDD.n12493 VSS 0.048151f
C32950 VDD.n12494 VSS 0.081176f
C32951 VDD.t3996 VSS 0.066856f
C32952 VDD.n12495 VSS 0.125227f
C32953 VDD.n12496 VSS 0.101294f
C32954 VDD.n12497 VSS 0.016021f
C32955 VDD.t3773 VSS 0.025104f
C32956 VDD.n12498 VSS 0.099723f
C32957 VDD.t797 VSS 0.066856f
C32958 VDD.n12499 VSS 0.125227f
C32959 VDD.t2426 VSS 0.025104f
C32960 VDD.n12500 VSS 0.083673f
C32961 VDD.t2424 VSS 0.066856f
C32962 VDD.n12501 VSS 0.125227f
C32963 VDD.n12502 VSS 0.101294f
C32964 VDD.n12503 VSS 0.016021f
C32965 VDD.t799 VSS 0.025104f
C32966 VDD.n12504 VSS 0.099723f
C32967 VDD.n12505 VSS 0.62132f
C32968 VDD.t2411 VSS 0.028519f
C32969 VDD.t2636 VSS 0.028519f
C32970 VDD.n12506 VSS 0.009191f
C32971 VDD.n12507 VSS 0.261039f
C32972 VDD.t2635 VSS 0.066856f
C32973 VDD.t4016 VSS 0.066856f
C32974 VDD.n12508 VSS 0.709674f
C32975 VDD.t752 VSS 0.028519f
C32976 VDD.t980 VSS 0.028519f
C32977 VDD.n12509 VSS 0.009191f
C32978 VDD.n12510 VSS 0.644755f
C32979 VDD.t978 VSS 0.066856f
C32980 VDD.t2502 VSS 0.066856f
C32981 VDD.n12511 VSS 0.690489f
C32982 VDD.t4722 VSS 0.066856f
C32983 VDD.t2056 VSS 0.066856f
C32984 VDD.n12512 VSS 0.690489f
C32985 VDD.t4491 VSS 0.028519f
C32986 VDD.t4723 VSS 0.028519f
C32987 VDD.n12513 VSS 0.009191f
C32988 VDD.n12514 VSS 0.523473f
C32989 VDD.n12515 VSS 0.524869f
C32990 VDD.n12516 VSS 0.208534f
C32991 VDD.n12517 VSS 0.865258f
C32992 VDD.n12518 VSS 0.865258f
C32993 VDD.t979 VSS 1.45794f
C32994 VDD.t751 VSS 1.96535f
C32995 VDD.t798 VSS 1.96535f
C32996 VDD.t2425 VSS 1.31955f
C32997 VDD.n12519 VSS 0.595476f
C32998 VDD.n12520 VSS 0.645798f
C32999 VDD.n12521 VSS 0.206947f
C33000 VDD.n12522 VSS 0.208534f
C33001 VDD.n12523 VSS 0.529799f
C33002 VDD.n12524 VSS 0.207221f
C33003 VDD.n12525 VSS 0.902999f
C33004 VDD.t689 VSS 1.45794f
C33005 VDD.t1613 VSS 1.96535f
C33006 VDD.t529 VSS 1.96535f
C33007 VDD.t535 VSS 1.31955f
C33008 VDD.n12526 VSS 0.595476f
C33009 VDD.n12527 VSS 0.645798f
C33010 VDD.t530 VSS 1.36988f
C33011 VDD.t528 VSS 1.96535f
C33012 VDD.t1517 VSS 1.96535f
C33013 VDD.t1302 VSS 1.45794f
C33014 VDD.n12528 VSS 0.865258f
C33015 VDD.n12529 VSS 0.208534f
C33016 VDD.n12530 VSS 0.524869f
C33017 VDD.t3529 VSS 0.028519f
C33018 VDD.t3736 VSS 0.028519f
C33019 VDD.n12531 VSS 0.009191f
C33020 VDD.t3374 VSS 0.028519f
C33021 VDD.t2322 VSS 0.028519f
C33022 VDD.n12532 VSS 0.009191f
C33023 VDD.n12533 VSS 0.523473f
C33024 VDD.t3528 VSS 0.066856f
C33025 VDD.t3373 VSS 0.066856f
C33026 VDD.t2321 VSS 0.066856f
C33027 VDD.t3735 VSS 0.066856f
C33028 VDD.n12534 VSS 0.690489f
C33029 VDD.t3892 VSS 0.066856f
C33030 VDD.t3741 VSS 0.066856f
C33031 VDD.t2739 VSS 0.066856f
C33032 VDD.t4128 VSS 0.066856f
C33033 VDD.n12535 VSS 0.690489f
C33034 VDD.t3893 VSS 0.028519f
C33035 VDD.t4129 VSS 0.028519f
C33036 VDD.n12536 VSS 0.009191f
C33037 VDD.t3742 VSS 0.028519f
C33038 VDD.t2740 VSS 0.028519f
C33039 VDD.n12537 VSS 0.009191f
C33040 VDD.n12538 VSS 0.644755f
C33041 VDD.t1301 VSS 0.066856f
C33042 VDD.t1157 VSS 0.066856f
C33043 VDD.t4252 VSS 0.066856f
C33044 VDD.t1516 VSS 0.066856f
C33045 VDD.n12539 VSS 0.709674f
C33046 VDD.t1303 VSS 0.028519f
C33047 VDD.t1518 VSS 0.028519f
C33048 VDD.n12540 VSS 0.009191f
C33049 VDD.t1159 VSS 0.028519f
C33050 VDD.t4253 VSS 0.028519f
C33051 VDD.n12541 VSS 0.009191f
C33052 VDD.n12542 VSS 0.261039f
C33053 VDD.n12543 VSS 0.62132f
C33054 VDD.n12544 VSS 0.099723f
C33055 VDD.t4266 VSS 0.066856f
C33056 VDD.n12545 VSS 0.125227f
C33057 VDD.n12546 VSS 0.101294f
C33058 VDD.n12547 VSS 0.016021f
C33059 VDD.t849 VSS 0.025104f
C33060 VDD.n12548 VSS 0.083673f
C33061 VDD.n12549 VSS 0.048151f
C33062 VDD.n12550 VSS 0.081176f
C33063 VDD.t3916 VSS 0.066856f
C33064 VDD.n12551 VSS 0.125227f
C33065 VDD.n12552 VSS 0.101294f
C33066 VDD.n12553 VSS 0.016021f
C33067 VDD.t1294 VSS 0.025104f
C33068 VDD.n12554 VSS 0.099723f
C33069 VDD.t4188 VSS 0.066856f
C33070 VDD.n12555 VSS 0.125227f
C33071 VDD.t756 VSS 0.025104f
C33072 VDD.t3828 VSS 0.066856f
C33073 VDD.n12556 VSS 0.125227f
C33074 VDD.t781 VSS 0.025104f
C33075 VDD.t3219 VSS 0.028519f
C33076 VDD.t3853 VSS 0.028519f
C33077 VDD.n12557 VSS 0.009191f
C33078 VDD.n12558 VSS 0.049743f
C33079 VDD.n12559 VSS 0.018625f
C33080 VDD.n12560 VSS 0.014751f
C33081 VDD.n12561 VSS 0.009688f
C33082 VDD.t835 VSS 0.066856f
C33083 VDD.t1483 VSS 0.066856f
C33084 VDD.n12563 VSS 0.343648f
C33085 VDD.t1165 VSS 0.028519f
C33086 VDD.t1850 VSS 0.028519f
C33087 VDD.n12564 VSS 0.009191f
C33088 VDD.n12565 VSS 0.320028f
C33089 VDD.t1164 VSS 0.066856f
C33090 VDD.t1849 VSS 0.066856f
C33091 VDD.n12566 VSS 0.342968f
C33092 VDD.t1767 VSS 0.066856f
C33093 VDD.t2563 VSS 0.066856f
C33094 VDD.n12567 VSS 0.342968f
C33095 VDD.t1768 VSS 0.028519f
C33096 VDD.t2564 VSS 0.028519f
C33097 VDD.n12568 VSS 0.009191f
C33098 VDD.n12569 VSS 0.234012f
C33099 VDD.n12570 VSS 0.260425f
C33100 VDD.t1176 VSS 0.028519f
C33101 VDD.t1863 VSS 0.028519f
C33102 VDD.n12571 VSS 0.009191f
C33103 VDD.n12572 VSS 0.259851f
C33104 VDD.t1175 VSS 0.066856f
C33105 VDD.t1862 VSS 0.066856f
C33106 VDD.n12573 VSS 0.342968f
C33107 VDD.t1537 VSS 0.066856f
C33108 VDD.t2297 VSS 0.066856f
C33109 VDD.n12574 VSS 0.342968f
C33110 VDD.t1538 VSS 0.028519f
C33111 VDD.t2298 VSS 0.028519f
C33112 VDD.n12575 VSS 0.009191f
C33113 VDD.n12576 VSS 0.320028f
C33114 VDD.t3218 VSS 0.066856f
C33115 VDD.t3852 VSS 0.066856f
C33116 VDD.n12577 VSS 0.293671f
C33117 VDD.n12579 VSS 0.009312f
C33118 VDD.n12580 VSS 0.018249f
C33119 VDD.n12581 VSS 0.058817f
C33120 VDD.n12582 VSS 1.19e-19
C33121 VDD.n12583 VSS 0.079896f
C33122 VDD.n12584 VSS 0.01502f
C33123 VDD.n12585 VSS 0.251246f
C33124 VDD.n12586 VSS 0.057353f
C33125 VDD.n12587 VSS 0.099723f
C33126 VDD.t780 VSS 0.066856f
C33127 VDD.n12588 VSS 0.125227f
C33128 VDD.n12589 VSS 0.101294f
C33129 VDD.n12590 VSS 0.016021f
C33130 VDD.t3829 VSS 0.025104f
C33131 VDD.n12591 VSS 0.081176f
C33132 VDD.n12592 VSS 0.206947f
C33133 VDD.n12593 VSS 0.048151f
C33134 VDD.n12594 VSS 0.083673f
C33135 VDD.t755 VSS 0.066856f
C33136 VDD.n12595 VSS 0.125227f
C33137 VDD.n12596 VSS 0.101294f
C33138 VDD.n12597 VSS 0.016021f
C33139 VDD.t4189 VSS 0.025104f
C33140 VDD.n12598 VSS 0.099723f
C33141 VDD.n12599 VSS 0.62132f
C33142 VDD.t1090 VSS 0.028519f
C33143 VDD.t4173 VSS 0.028519f
C33144 VDD.n12600 VSS 0.009191f
C33145 VDD.n12601 VSS 0.261039f
C33146 VDD.t4172 VSS 0.066856f
C33147 VDD.t3944 VSS 0.066856f
C33148 VDD.n12602 VSS 0.709674f
C33149 VDD.t3639 VSS 0.028519f
C33150 VDD.t2646 VSS 0.028519f
C33151 VDD.n12603 VSS 0.009191f
C33152 VDD.n12604 VSS 0.644755f
C33153 VDD.t2645 VSS 0.066856f
C33154 VDD.t2416 VSS 0.066856f
C33155 VDD.n12605 VSS 0.690489f
C33156 VDD.t2207 VSS 0.066856f
C33157 VDD.t1967 VSS 0.066856f
C33158 VDD.n12606 VSS 0.690489f
C33159 VDD.t3309 VSS 0.028519f
C33160 VDD.t2208 VSS 0.028519f
C33161 VDD.n12607 VSS 0.009191f
C33162 VDD.n12608 VSS 0.523473f
C33163 VDD.n12609 VSS 0.524869f
C33164 VDD.n12610 VSS 0.208534f
C33165 VDD.n12611 VSS 0.865258f
C33166 VDD.n12612 VSS 0.865258f
C33167 VDD.t1782 VSS 1.45794f
C33168 VDD.t1089 VSS 1.96535f
C33169 VDD.t328 VSS 1.96535f
C33170 VDD.t330 VSS 1.31955f
C33171 VDD.n12613 VSS 0.595476f
C33172 VDD.n12614 VSS 0.208771f
C33173 VDD.n12615 VSS 0.057098f
C33174 VDD.n12616 VSS 0.105404f
C33175 VDD.t1467 VSS 0.066856f
C33176 VDD.n12617 VSS 0.14405f
C33177 VDD.n12618 VSS 0.120118f
C33178 VDD.n12619 VSS 0.016021f
C33179 VDD.t2666 VSS 0.025104f
C33180 VDD.n12620 VSS 0.116823f
C33181 VDD.n12621 VSS 0.08646f
C33182 VDD.n12623 VSS 0.018625f
C33183 VDD.t837 VSS 0.028519f
C33184 VDD.t1485 VSS 0.028519f
C33185 VDD.n12624 VSS 0.009191f
C33186 VDD.n12625 VSS 0.052803f
C33187 VDD.n12626 VSS 0.272325f
C33188 VDD.n12628 VSS 0.01502f
C33189 VDD.n12629 VSS 0.01487f
C33190 VDD.n12630 VSS 0.036378f
C33191 VDD.n12631 VSS 0.018249f
C33192 VDD.n12632 VSS 0.009312f
C33193 VDD.n12633 VSS 1.76802f
C33194 VDD.n12634 VSS 2.45351f
C33195 VDD.n12635 VSS 0.009312f
C33196 VDD.n12636 VSS 0.009688f
C33197 VDD.n12638 VSS 0.018625f
C33198 VDD.t4001 VSS 0.034186f
C33199 VDD.n12639 VSS 0.203247f
C33200 VDD.n12640 VSS 0.177689f
C33201 VDD.n12641 VSS 0.01502f
C33202 VDD.n12642 VSS 0.118218f
C33203 VDD.n12643 VSS 0.103711f
C33204 VDD.t4000 VSS 0.080376f
C33205 a_52635_34067.n0 VSS 0.968206f
C33206 a_52635_34067.n1 VSS 1.05429f
C33207 a_52635_34067.n2 VSS 0.519869f
C33208 a_52635_34067.n3 VSS 0.968206f
C33209 a_52635_34067.n4 VSS 1.05429f
C33210 a_52635_34067.n5 VSS 0.393308f
C33211 a_52635_34067.n6 VSS 1.04685f
C33212 a_52635_34067.n7 VSS 0.772359f
C33213 a_52635_34067.n8 VSS 0.570135f
C33214 a_52635_34067.n9 VSS 0.772359f
C33215 a_52635_34067.n10 VSS 1.04685f
C33216 a_52635_34067.n11 VSS 0.389035f
C33217 a_52635_34067.n12 VSS 1.05549f
C33218 a_52635_34067.n13 VSS 0.769973f
C33219 a_52635_34067.n14 VSS 0.563421f
C33220 a_52635_34067.n15 VSS 0.294912f
C33221 a_52635_34067.n16 VSS 0.609476f
C33222 a_52635_34067.n17 VSS 0.726532f
C33223 a_52635_34067.n18 VSS 0.988415f
C33224 a_52635_34067.n19 VSS 1.35551f
C33225 a_52635_34067.n20 VSS 0.390166f
C33226 a_52635_34067.n21 VSS 1.35551f
C33227 a_52635_34067.n22 VSS 0.988415f
C33228 a_52635_34067.n23 VSS 0.563421f
C33229 a_52635_34067.n24 VSS 0.769973f
C33230 a_52635_34067.n25 VSS 1.05549f
C33231 a_52635_34067.n26 VSS 0.964177f
C33232 a_52635_34067.n27 VSS 1.05056f
C33233 a_52635_34067.n28 VSS 0.519502f
C33234 a_52635_34067.n29 VSS 0.964177f
C33235 a_52635_34067.n30 VSS 1.05056f
C33236 a_52635_34067.n31 VSS 0.392989f
C33237 a_52635_34067.n32 VSS 0.989056f
C33238 a_52635_34067.n33 VSS 1.34521f
C33239 a_52635_34067.n34 VSS 0.716481f
C33240 a_52635_34067.n35 VSS 0.989056f
C33241 a_52635_34067.n36 VSS 1.34521f
C33242 a_52635_34067.n37 VSS 0.389035f
C33243 a_52635_34067.n38 VSS 0.609476f
C33244 a_52635_34067.n39 VSS 0.744707f
C33245 a_52635_34067.n40 VSS 0.294912f
C33246 a_52635_34067.n41 VSS 0.389035f
C33247 a_52635_34067.n42 VSS 0.744707f
C33248 a_52635_34067.n43 VSS 0.599484f
C33249 a_52635_34067.n44 VSS 1.50271f
C33250 a_52635_34067.n45 VSS 0.599484f
C33251 a_52635_34067.n46 VSS 0.716481f
C33252 a_52635_34067.n47 VSS 0.750489f
C33253 a_52635_34067.n48 VSS 0.393308f
C33254 a_52635_34067.n49 VSS 0.750489f
C33255 a_52635_34067.n50 VSS 0.296169f
C33256 a_52635_34067.n51 VSS 0.393308f
C33257 a_52635_34067.n52 VSS 0.296169f
C33258 a_52635_34067.n53 VSS 0.970844f
C33259 a_52635_34067.n54 VSS 0.94646f
C33260 a_52635_34067.n55 VSS 2.60562f
C33261 a_52635_34067.n56 VSS 0.854303f
C33262 a_52635_34067.n57 VSS 1.10968f
C33263 a_52635_34067.n58 VSS 1.8542f
C33264 a_52635_34067.n59 VSS 0.647472f
C33265 a_52635_34067.n60 VSS 2.60562f
C33266 a_52635_34067.n61 VSS 1.05782f
C33267 a_52635_34067.n62 VSS 0.613009f
C33268 a_52635_34067.n63 VSS 0.854303f
C33269 a_52635_34067.n64 VSS 2.60562f
C33270 a_52635_34067.n65 VSS 0.94646f
C33271 a_52635_34067.n66 VSS 0.667926f
C33272 a_52635_34067.n67 VSS 1.05782f
C33273 a_52635_34067.n68 VSS 2.60562f
C33274 a_52635_34067.n69 VSS 0.970844f
C33275 a_52635_34067.n70 VSS 1.3574f
C33276 a_52635_34067.n71 VSS 1.04844f
C33277 a_52635_34067.n72 VSS 0.879472f
C33278 a_52635_34067.n73 VSS 0.92402f
C33279 a_52635_34067.n74 VSS 2.64985f
C33280 a_52635_34067.n75 VSS 2.65467f
C33281 a_52635_34067.n76 VSS 0.97646f
C33282 a_52635_34067.n77 VSS 0.6236f
C33283 a_52635_34067.n78 VSS 0.654457f
C33284 a_52635_34067.n79 VSS 2.65467f
C33285 a_52635_34067.n80 VSS 1.04847f
C33286 a_52635_34067.n81 VSS 0.879464f
C33287 a_52635_34067.n82 VSS 2.64985f
C33288 a_52635_34067.n83 VSS 0.924019f
C33289 a_52635_34067.n84 VSS 0.976487f
C33290 a_52635_34067.n85 VSS 0.726532f
C33291 a_52635_34067.n86 VSS 1.8542f
C33292 a_52635_34067.n87 VSS 0.647472f
C33293 a_52635_34067.n88 VSS 1.8542f
C33294 a_52635_34067.n89 VSS 0.648333f
C33295 a_52635_34067.n90 VSS 1.8542f
C33296 a_52635_34067.n91 VSS 0.648333f
C33297 a_52635_34067.n92 VSS 2.51871f
C33298 a_52635_34067.n93 VSS 1.36384f
C33299 a_52635_34067.n94 VSS 1.36384f
C33300 a_52635_34067.n95 VSS 2.51871f
C33301 a_52635_34067.n96 VSS 1.93502f
C33302 a_52635_34067.n97 VSS 0.686888f
C33303 a_52635_34067.n98 VSS 1.93502f
C33304 a_52635_34067.n99 VSS 0.638844f
C33305 a_52635_34067.n100 VSS 1.93502f
C33306 a_52635_34067.n101 VSS 0.686973f
C33307 a_52635_34067.n102 VSS 1.93502f
C33308 a_52635_34067.n103 VSS 0.638862f
C33309 a_52635_34067.n104 VSS 2.54563f
C33310 a_52635_34067.n105 VSS 1.38682f
C33311 a_52635_34067.n106 VSS 1.38682f
C33312 a_52635_34067.n107 VSS 2.54563f
C33313 a_52635_34067.n108 VSS 0.667926f
C33314 a_52635_34067.n109 VSS 2.51775f
C33315 a_52635_34067.n110 VSS 1.10968f
C33316 a_52635_34067.n111 VSS 2.51775f
C33317 a_52635_34067.n112 VSS 2.53332f
C33318 a_52635_34067.n113 VSS 1.11217f
C33319 a_52635_34067.n114 VSS 1.38815f
C33320 a_52635_34067.n115 VSS 1.11218f
C33321 a_52635_34067.n116 VSS 2.53332f
C33322 a_52635_34067.n117 VSS 0.613009f
C33323 a_52635_34067.t166 VSS 0.532505f
C33324 a_52635_34067.t90 VSS 0.532505f
C33325 a_52635_34067.n118 VSS 0.812262f
C33326 a_52635_34067.n119 VSS 0.634239f
C33327 a_52635_34067.n120 VSS 0.695643f
C33328 a_52635_34067.n121 VSS 0.557311f
C33329 a_52635_34067.n122 VSS 0.705817f
C33330 a_52635_34067.n123 VSS 0.705816f
C33331 a_52635_34067.n124 VSS 0.456895f
C33332 a_52635_34067.n125 VSS 0.634239f
C33333 a_52635_34067.n126 VSS 0.695643f
C33334 a_52635_34067.n127 VSS 0.910818f
C33335 a_52635_34067.n128 VSS 0.812262f
C33336 a_52635_34067.n129 VSS 0.634239f
C33337 a_52635_34067.n130 VSS 0.695643f
C33338 a_52635_34067.n131 VSS 0.557311f
C33339 a_52635_34067.n132 VSS 0.705817f
C33340 a_52635_34067.n133 VSS 0.705816f
C33341 a_52635_34067.n134 VSS 0.456895f
C33342 a_52635_34067.n135 VSS 0.634239f
C33343 a_52635_34067.n136 VSS 0.695643f
C33344 a_52635_34067.n137 VSS 0.910818f
C33345 a_52635_34067.n138 VSS 1.16767f
C33346 a_52635_34067.t45 VSS 1.50638f
C33347 a_52635_34067.n139 VSS 0.706418f
C33348 a_52635_34067.n140 VSS 2.01071f
C33349 a_52635_34067.n141 VSS 0.815817f
C33350 a_52635_34067.n142 VSS 0.904816f
C33351 a_52635_34067.t60 VSS 0.323218f
C33352 a_52635_34067.t48 VSS 0.283215f
C33353 a_52635_34067.t31 VSS 0.245001f
C33354 a_52635_34067.n143 VSS 0.696281f
C33355 a_52635_34067.t55 VSS 0.242904f
C33356 a_52635_34067.n144 VSS 0.630882f
C33357 a_52635_34067.n145 VSS 2.65583f
C33358 a_52635_34067.n146 VSS 2.3552f
C33359 a_52635_34067.t40 VSS 1.08042f
C33360 a_52635_34067.t17 VSS 3.04611f
C33361 a_52635_34067.n147 VSS 3.51664f
C33362 a_52635_34067.n148 VSS 3.42219f
C33363 a_52635_34067.t216 VSS 0.481804f
C33364 a_52635_34067.t117 VSS 0.481804f
C33365 a_52635_34067.t203 VSS 0.481804f
C33366 a_52635_34067.t240 VSS 0.481804f
C33367 a_52635_34067.t213 VSS 0.481804f
C33368 a_52635_34067.t144 VSS 0.481804f
C33369 a_52635_34067.t212 VSS 0.5311f
C33370 a_52635_34067.n149 VSS 1.45207f
C33371 a_52635_34067.t94 VSS 0.481804f
C33372 a_52635_34067.t152 VSS 0.5311f
C33373 a_52635_34067.t153 VSS 0.481804f
C33374 a_52635_34067.t200 VSS 0.481804f
C33375 a_52635_34067.t220 VSS 0.481804f
C33376 a_52635_34067.n150 VSS 0.390166f
C33377 a_52635_34067.t230 VSS 0.481804f
C33378 a_52635_34067.n151 VSS 0.320807f
C33379 a_52635_34067.t147 VSS 0.481804f
C33380 a_52635_34067.t124 VSS 0.481804f
C33381 a_52635_34067.t138 VSS 0.481804f
C33382 a_52635_34067.t75 VSS 0.481804f
C33383 a_52635_34067.t135 VSS 0.481804f
C33384 a_52635_34067.t130 VSS 0.481804f
C33385 a_52635_34067.t156 VSS 0.481804f
C33386 a_52635_34067.t215 VSS 0.481804f
C33387 a_52635_34067.t107 VSS 0.481804f
C33388 a_52635_34067.t167 VSS 0.481804f
C33389 a_52635_34067.t80 VSS 0.481804f
C33390 a_52635_34067.n152 VSS 0.392989f
C33391 a_52635_34067.t95 VSS 0.481804f
C33392 a_52635_34067.n153 VSS 0.320807f
C33393 a_52635_34067.t202 VSS 0.481804f
C33394 a_52635_34067.t74 VSS 0.481804f
C33395 a_52635_34067.t134 VSS 0.481804f
C33396 a_52635_34067.t150 VSS 0.481804f
C33397 a_52635_34067.t173 VSS 0.481804f
C33398 a_52635_34067.t87 VSS 0.481804f
C33399 a_52635_34067.t148 VSS 0.481804f
C33400 a_52635_34067.t143 VSS 0.481804f
C33401 a_52635_34067.t207 VSS 0.481804f
C33402 a_52635_34067.n154 VSS 0.392989f
C33403 a_52635_34067.t78 VSS 0.481804f
C33404 a_52635_34067.n155 VSS 0.320807f
C33405 a_52635_34067.t180 VSS 0.481804f
C33406 a_52635_34067.t221 VSS 0.481804f
C33407 a_52635_34067.t70 VSS 0.481804f
C33408 a_52635_34067.t133 VSS 0.532581f
C33409 a_52635_34067.t139 VSS 0.481804f
C33410 a_52635_34067.n156 VSS 5.15047f
C33411 a_52635_34067.t126 VSS 0.481804f
C33412 a_52635_34067.t211 VSS 0.481804f
C33413 a_52635_34067.t236 VSS 0.481804f
C33414 a_52635_34067.t121 VSS 0.533512f
C33415 a_52635_34067.t132 VSS 0.481804f
C33416 a_52635_34067.n157 VSS 0.389035f
C33417 a_52635_34067.t219 VSS 0.481804f
C33418 a_52635_34067.n158 VSS 0.320807f
C33419 a_52635_34067.t154 VSS 0.481804f
C33420 a_52635_34067.t157 VSS 0.481804f
C33421 a_52635_34067.t239 VSS 0.481804f
C33422 a_52635_34067.t142 VSS 0.481804f
C33423 a_52635_34067.n159 VSS 5.15047f
C33424 a_52635_34067.t218 VSS 0.481804f
C33425 a_52635_34067.t91 VSS 0.481804f
C33426 a_52635_34067.t131 VSS 0.481804f
C33427 a_52635_34067.t192 VSS 0.481804f
C33428 a_52635_34067.n160 VSS 0.392989f
C33429 a_52635_34067.t208 VSS 0.481804f
C33430 a_52635_34067.n161 VSS 0.320807f
C33431 a_52635_34067.t119 VSS 0.481804f
C33432 a_52635_34067.t186 VSS 0.481804f
C33433 a_52635_34067.t237 VSS 0.481804f
C33434 a_52635_34067.t204 VSS 0.481804f
C33435 a_52635_34067.t71 VSS 0.481804f
C33436 a_52635_34067.t68 VSS 0.481804f
C33437 a_52635_34067.t67 VSS 0.481804f
C33438 a_52635_34067.t141 VSS 0.481804f
C33439 a_52635_34067.t184 VSS 0.481804f
C33440 a_52635_34067.t234 VSS 0.532581f
C33441 a_52635_34067.t103 VSS 0.481804f
C33442 a_52635_34067.n162 VSS 0.393308f
C33443 a_52635_34067.t190 VSS 0.481804f
C33444 a_52635_34067.n163 VSS 0.320807f
C33445 a_52635_34067.t125 VSS 0.481804f
C33446 a_52635_34067.t96 VSS 0.481804f
C33447 a_52635_34067.t73 VSS 0.481804f
C33448 a_52635_34067.t82 VSS 0.481804f
C33449 a_52635_34067.n164 VSS 3.42219f
C33450 a_52635_34067.n165 VSS 3.42219f
C33451 a_52635_34067.t102 VSS 0.481804f
C33452 a_52635_34067.t198 VSS 0.481804f
C33453 a_52635_34067.t129 VSS 0.481804f
C33454 a_52635_34067.t197 VSS 0.481804f
C33455 a_52635_34067.t228 VSS 0.481804f
C33456 a_52635_34067.t118 VSS 0.481804f
C33457 a_52635_34067.t222 VSS 0.481804f
C33458 a_52635_34067.t99 VSS 0.481804f
C33459 a_52635_34067.t160 VSS 0.481804f
C33460 a_52635_34067.t177 VSS 0.481804f
C33461 a_52635_34067.t175 VSS 0.481804f
C33462 a_52635_34067.t171 VSS 0.481804f
C33463 a_52635_34067.t120 VSS 0.481804f
C33464 a_52635_34067.t235 VSS 0.481804f
C33465 a_52635_34067.t109 VSS 0.481804f
C33466 a_52635_34067.t226 VSS 0.481804f
C33467 a_52635_34067.t65 VSS 0.481804f
C33468 a_52635_34067.t185 VSS 0.481804f
C33469 a_52635_34067.t123 VSS 0.481804f
C33470 a_52635_34067.t187 VSS 0.481804f
C33471 a_52635_34067.t224 VSS 0.481804f
C33472 a_52635_34067.t79 VSS 0.481804f
C33473 a_52635_34067.t182 VSS 0.481804f
C33474 a_52635_34067.t174 VSS 0.481804f
C33475 a_52635_34067.t93 VSS 0.481804f
C33476 a_52635_34067.t151 VSS 0.481804f
C33477 a_52635_34067.t168 VSS 0.481804f
C33478 a_52635_34067.t238 VSS 0.481804f
C33479 a_52635_34067.t162 VSS 0.481804f
C33480 a_52635_34067.t155 VSS 0.481804f
C33481 a_52635_34067.t232 VSS 0.481804f
C33482 a_52635_34067.t88 VSS 0.481804f
C33483 a_52635_34067.t149 VSS 0.481804f
C33484 a_52635_34067.t189 VSS 0.481804f
C33485 a_52635_34067.t161 VSS 0.481804f
C33486 a_52635_34067.t165 VSS 0.481804f
C33487 a_52635_34067.t106 VSS 0.481804f
C33488 a_52635_34067.t194 VSS 0.481804f
C33489 a_52635_34067.n166 VSS 5.34875f
C33490 a_52635_34067.t231 VSS 0.481804f
C33491 a_52635_34067.t179 VSS 0.481804f
C33492 a_52635_34067.t137 VSS 0.481804f
C33493 a_52635_34067.t77 VSS 0.481804f
C33494 a_52635_34067.t136 VSS 0.481804f
C33495 a_52635_34067.t66 VSS 0.481804f
C33496 a_52635_34067.t164 VSS 0.481804f
C33497 a_52635_34067.t127 VSS 0.481804f
C33498 a_52635_34067.t122 VSS 0.481804f
C33499 a_52635_34067.t140 VSS 0.481804f
C33500 a_52635_34067.t116 VSS 0.481804f
C33501 a_52635_34067.t229 VSS 0.481804f
C33502 a_52635_34067.t146 VSS 0.481804f
C33503 a_52635_34067.t195 VSS 0.481804f
C33504 a_52635_34067.t225 VSS 0.481804f
C33505 a_52635_34067.t105 VSS 0.481804f
C33506 a_52635_34067.t112 VSS 0.481804f
C33507 a_52635_34067.n167 VSS 5.34875f
C33508 a_52635_34067.t111 VSS 0.481804f
C33509 a_52635_34067.t92 VSS 0.481804f
C33510 a_52635_34067.t206 VSS 0.481804f
C33511 a_52635_34067.t97 VSS 0.481804f
C33512 a_52635_34067.t145 VSS 0.481804f
C33513 a_52635_34067.t227 VSS 0.481804f
C33514 a_52635_34067.t108 VSS 0.481804f
C33515 a_52635_34067.t110 VSS 0.481804f
C33516 a_52635_34067.t191 VSS 0.481804f
C33517 a_52635_34067.t104 VSS 0.481804f
C33518 a_52635_34067.t172 VSS 0.481804f
C33519 a_52635_34067.t76 VSS 0.481804f
C33520 a_52635_34067.t113 VSS 0.481804f
C33521 a_52635_34067.t217 VSS 0.481804f
C33522 a_52635_34067.t89 VSS 0.481804f
C33523 a_52635_34067.t83 VSS 0.481804f
C33524 a_52635_34067.t170 VSS 0.481804f
C33525 a_52635_34067.t86 VSS 0.481804f
C33526 a_52635_34067.t81 VSS 0.481804f
C33527 a_52635_34067.t158 VSS 0.481804f
C33528 a_52635_34067.t205 VSS 0.481804f
C33529 a_52635_34067.t72 VSS 0.481804f
C33530 a_52635_34067.n168 VSS 3.42219f
C33531 a_52635_34067.n169 VSS 3.48946f
C33532 a_52635_34067.t169 VSS 0.481804f
C33533 a_52635_34067.t100 VSS 0.481804f
C33534 a_52635_34067.t209 VSS 0.481804f
C33535 a_52635_34067.t163 VSS 0.481804f
C33536 a_52635_34067.t233 VSS 0.481804f
C33537 a_52635_34067.t98 VSS 0.481804f
C33538 a_52635_34067.t159 VSS 0.481804f
C33539 a_52635_34067.t223 VSS 0.481804f
C33540 a_52635_34067.t114 VSS 0.481804f
C33541 a_52635_34067.t201 VSS 0.481804f
C33542 a_52635_34067.t183 VSS 0.481804f
C33543 a_52635_34067.n170 VSS 3.8813f
C33544 a_52635_34067.n171 VSS 2.83365f
C33545 a_52635_34067.n172 VSS 3.65877f
C33546 a_52635_34067.n173 VSS 0.519869f
C33547 a_52635_34067.t85 VSS 0.481804f
C33548 a_52635_34067.n174 VSS 0.390166f
C33549 a_52635_34067.t101 VSS 0.481804f
C33550 a_52635_34067.n175 VSS 0.320807f
C33551 a_52635_34067.t210 VSS 0.481804f
C33552 a_52635_34067.t178 VSS 0.481804f
C33553 a_52635_34067.t199 VSS 0.481804f
C33554 a_52635_34067.t128 VSS 0.481804f
C33555 a_52635_34067.t196 VSS 0.481804f
C33556 a_52635_34067.t188 VSS 0.481804f
C33557 a_52635_34067.t214 VSS 0.481804f
C33558 a_52635_34067.n176 VSS 0.390166f
C33559 a_52635_34067.t84 VSS 0.481804f
C33560 a_52635_34067.n177 VSS 0.320807f
C33561 a_52635_34067.t193 VSS 0.481804f
C33562 a_52635_34067.t176 VSS 0.533512f
C33563 a_52635_34067.t115 VSS 0.481804f
C33564 a_52635_34067.t69 VSS 0.481804f
C33565 a_52635_34067.t181 VSS 0.481804f
C33566 a_52635_34067.n178 VSS 3.65877f
C33567 a_52635_34067.n179 VSS 2.14406f
C33568 a_52635_34067.t49 VSS 0.32777f
C33569 a_52635_34067.t34 VSS 0.283215f
C33570 a_52635_34067.n180 VSS 2.39757f
C33571 a_52635_34067.n181 VSS 2.73209f
C33572 a_52635_34067.n182 VSS 0.904816f
C33573 a_52635_34067.t10 VSS 0.323218f
C33574 a_52635_34067.t11 VSS 0.283215f
C33575 a_52635_34067.t33 VSS 0.245001f
C33576 a_52635_34067.n183 VSS 0.696281f
C33577 a_52635_34067.t59 VSS 0.242904f
C33578 a_52635_34067.n184 VSS 0.630882f
C33579 a_52635_34067.t2 VSS 0.325302f
C33580 a_52635_34067.t63 VSS 0.278851f
C33581 a_52635_34067.t64 VSS 0.239255f
C33582 a_52635_34067.n185 VSS 0.715351f
C33583 a_52635_34067.t62 VSS 0.322103f
C33584 a_52635_34067.n186 VSS 1.28863f
C33585 a_52635_34067.t4 VSS 2.58185f
C33586 a_52635_34067.t0 VSS 0.550597f
C33587 a_52635_34067.n187 VSS 3.88688f
C33588 a_52635_34067.t61 VSS 0.783671f
C33589 a_52635_34067.t1 VSS 1.9214f
C33590 a_52635_34067.t3 VSS 0.322492f
C33591 a_52635_34067.n188 VSS 0.664421f
C33592 a_52635_34067.n189 VSS 2.80961f
C33593 a_52635_34067.n190 VSS 4.57473f
C33594 a_52635_34067.t28 VSS 0.326259f
C33595 a_52635_34067.t29 VSS 0.282773f
C33596 a_52635_34067.t38 VSS 0.244504f
C33597 a_52635_34067.t26 VSS 0.244187f
C33598 a_52635_34067.t9 VSS 0.282773f
C33599 a_52635_34067.t24 VSS 0.244504f
C33600 a_52635_34067.t32 VSS 0.244504f
C33601 a_52635_34067.t23 VSS 0.282773f
C33602 a_52635_34067.t16 VSS 0.244504f
C33603 a_52635_34067.t14 VSS 0.244187f
C33604 a_52635_34067.t41 VSS 0.282773f
C33605 a_52635_34067.t8 VSS 0.326696f
C33606 a_52635_34067.n191 VSS 3.72315f
C33607 a_52635_34067.n192 VSS 0.160921f
C33608 a_52635_34067.n193 VSS 0.160921f
C33609 a_52635_34067.n194 VSS 3.69214f
C33610 a_52635_34067.t44 VSS 1.08042f
C33611 a_52635_34067.t27 VSS 3.04611f
C33612 a_52635_34067.t18 VSS 0.392987f
C33613 a_52635_34067.t21 VSS 1.21614f
C33614 a_52635_34067.t30 VSS 0.340802f
C33615 a_52635_34067.n195 VSS 1.5238f
C33616 a_52635_34067.n196 VSS 2.37199f
C33617 a_52635_34067.n197 VSS 2.11719f
C33618 a_52635_34067.n198 VSS 0.160928f
C33619 a_52635_34067.t43 VSS 0.283215f
C33620 a_52635_34067.n199 VSS 0.457208f
C33621 a_52635_34067.t56 VSS 0.244933f
C33622 a_52635_34067.n200 VSS 0.706418f
C33623 a_52635_34067.t15 VSS 0.242904f
C33624 a_52635_34067.n201 VSS 0.700675f
C33625 a_52635_34067.t47 VSS 0.283215f
C33626 a_52635_34067.n202 VSS 0.557196f
C33627 a_52635_34067.t53 VSS 0.245001f
C33628 a_52635_34067.n203 VSS 0.696281f
C33629 a_52635_34067.t51 VSS 0.242904f
C33630 a_52635_34067.n204 VSS 0.630882f
C33631 a_52635_34067.n205 VSS 0.815817f
C33632 a_52635_34067.t50 VSS 0.32777f
C33633 a_52635_34067.t35 VSS 0.283215f
C33634 a_52635_34067.n206 VSS 0.160928f
C33635 a_52635_34067.n207 VSS 2.11719f
C33636 a_52635_34067.t19 VSS 0.326259f
C33637 a_52635_34067.t20 VSS 0.282773f
C33638 a_52635_34067.t36 VSS 0.244504f
C33639 a_52635_34067.t12 VSS 0.244187f
C33640 a_52635_34067.n208 VSS 0.160921f
C33641 a_52635_34067.t46 VSS 0.282773f
C33642 a_52635_34067.t7 VSS 0.244504f
C33643 a_52635_34067.t25 VSS 0.244504f
C33644 a_52635_34067.t6 VSS 0.282773f
C33645 a_52635_34067.t58 VSS 0.244504f
C33646 a_52635_34067.t57 VSS 0.244187f
C33647 a_52635_34067.t37 VSS 0.282773f
C33648 a_52635_34067.t54 VSS 0.326696f
C33649 a_52635_34067.n209 VSS 0.160921f
C33650 a_52635_34067.n210 VSS 2.3552f
C33651 a_52635_34067.n211 VSS 2.73209f
C33652 a_52635_34067.t39 VSS 0.392987f
C33653 a_52635_34067.t13 VSS 1.21614f
C33654 a_52635_34067.t22 VSS 0.340802f
C33655 a_52635_34067.n212 VSS 1.5238f
C33656 a_52635_34067.n213 VSS 2.37199f
C33657 a_52635_34067.n214 VSS 2.13513f
C33658 a_52635_34067.n215 VSS 0.160928f
C33659 a_52635_34067.t42 VSS 0.283215f
C33660 a_52635_34067.n216 VSS 0.457208f
C33661 a_52635_34067.t52 VSS 0.244933f
C33662 a_52635_34067.t5 VSS 0.242904f
.ends

