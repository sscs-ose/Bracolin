** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/PRbiased_net.sch
.subckt PRbiased_net VA VB IBN IBP ITN ITP VDD VSS
*.PININFO VA:B VB:B IBN:B IBP:B ITN:B ITP:B VDD:B VSS:B
x1 VA VB net1 net2 IBN IBP vc VDD VSS PR_net
x2 IBN vc net1 ITN VDD VSS DiffN_net
x3 IBP vc net2 ITP VDD VSS DiffP_net
.ends

* expanding   symbol:  PR_net.sym # of pins=9
** sym_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/PR_net.sym
** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/PR_net.sch
.subckt PR_net VA VB VG_N VG_P IB_N IB_P VC VDD VSS
*.PININFO VA:B VB:B VG_N:B VG_P:B IB_N:B IB_P:B VC:B VDD:B VSS:B
x1 VDD net1 IB_N net2 VG_N VC VSS PR_nfets
x2 IB_P VSS VA VB VG_P net1 net2 VDD PR_pfets
.ends


* expanding   symbol:  DiffN_net.sym # of pins=6
** sym_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/DiffN_net.sym
** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/DiffN_net.sch
.subckt DiffN_net VN VP OUT IT VDD VSS
*.PININFO VN:B VP:B OUT:B IT:B VDD:B VSS:B
x1 net1 OUT VP VN IT VSS DiffN_nfets
x2 net1 OUT net1 VDD VDD DiffN_pfets
.ends


* expanding   symbol:  DiffP_net.sym # of pins=6
** sym_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/DiffP_net.sym
** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/DiffP_net.sch
.subckt DiffP_net VN VP OUT IT VDD VSS
*.PININFO VN:B VP:B OUT:B IT:B VDD:B VSS:B
x1 net1 OUT net1 VSS VSS DiffP_nfets
x2 net1 OUT VP VN IT VDD DiffP_pfets
.ends


* expanding   symbol:  PR_nfets.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/PR_nfets.sym
** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/PR_nfets.sch
.subckt PR_nfets VD1 VD2 VS1 VS2 VG VC VB
*.PININFO VD1:B VD2:B VS1:B VS2:B VG:B VC:B VB:B
M5[1] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[2] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[3] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[4] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[5] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[6] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[7] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[8] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[9] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[10] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[11] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[12] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[13] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[14] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[15] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[16] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[17] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[18] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[19] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[20] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[21] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[22] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[23] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[24] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[25] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[26] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[27] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[28] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[29] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[30] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[31] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M5[32] VB VB VB VB nfet_03v3 L=2u W=2u nf=1 m=1
M3 VD2 VG net1 VB nfet_03v3 L=2u W=2u nf=1 m=1
M4 net1 VG VC VB nfet_03v3 L=2u W=2u nf=1 m=1
M6 VD2 VG net2 VB nfet_03v3 L=2u W=2u nf=1 m=1
M8 net2 VG VC VB nfet_03v3 L=2u W=2u nf=1 m=1
M1 VC VG net3 VB nfet_03v3 L=2u W=2u nf=1 m=1
M9 net3 VG VS2 VB nfet_03v3 L=2u W=2u nf=1 m=1
M10 VC VG net4 VB nfet_03v3 L=2u W=2u nf=1 m=1
M11 net4 VG VS2 VB nfet_03v3 L=2u W=2u nf=1 m=1
M2 VD1 VG net5 VB nfet_03v3 L=2u W=2u nf=1 m=1
M12 net5 VG VS1 VB nfet_03v3 L=2u W=2u nf=1 m=1
M13 VD1 VG net6 VB nfet_03v3 L=2u W=2u nf=1 m=1
M14 net6 VG VS1 VB nfet_03v3 L=2u W=2u nf=1 m=1
M7 VD1 VG net7 VB nfet_03v3 L=2u W=2u nf=1 m=1
M15 net7 VG VS1 VB nfet_03v3 L=2u W=2u nf=1 m=1
M16 VD1 VG net8 VB nfet_03v3 L=2u W=2u nf=1 m=1
M17 net8 VG VS1 VB nfet_03v3 L=2u W=2u nf=1 m=1
.ends


* expanding   symbol:  PR_pfets.sym # of pins=8
** sym_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/PR_pfets.sym
** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/PR_pfets.sch
.subckt PR_pfets VD1 VS1 VS2_A VS2_B VG VC_A VC_B VB
*.PININFO VD1:B VS1:B VS2_A:B VS2_B:B VG:B VC_A:B VC_B:B VB:B
M1 net3 VG VS1 VB pfet_03v3 L=2u W=2u nf=1 m=1
M2 VD1 VG net3 VB pfet_03v3 L=2u W=2u nf=1 m=1
M5 net4 VG VS1 VB pfet_03v3 L=2u W=2u nf=1 m=1
M6 VD1 VG net4 VB pfet_03v3 L=2u W=2u nf=1 m=1
M7 net5 VG VS1 VB pfet_03v3 L=2u W=2u nf=1 m=1
M9 VD1 VG net5 VB pfet_03v3 L=2u W=2u nf=1 m=1
M10 net6 VG VS1 VB pfet_03v3 L=2u W=2u nf=1 m=1
M11 VD1 VG net6 VB pfet_03v3 L=2u W=2u nf=1 m=1
M12 net1 VG VS2_A VB pfet_03v3 L=2u W=2u nf=1 m=1
M13 VC_A VG net1 VB pfet_03v3 L=2u W=2u nf=1 m=1
M14 net2 VG VS2_A VB pfet_03v3 L=2u W=2u nf=1 m=1
M15 VC_A VG net2 VB pfet_03v3 L=2u W=2u nf=1 m=1
M16 VC_B VG net7 VB pfet_03v3 L=2u W=2u nf=1 m=1
M17 net7 VG VS2_B VB pfet_03v3 L=2u W=2u nf=1 m=1
M18 VC_B VG net8 VB pfet_03v3 L=2u W=2u nf=1 m=1
M19 net8 VG VS2_B VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[1] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[2] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[3] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[4] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[5] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[6] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[7] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[8] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[9] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[10] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[11] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[12] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[13] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[14] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[15] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[16] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[17] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[18] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[19] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[20] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[21] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[22] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[23] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[24] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[25] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[26] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[27] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[28] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[29] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[30] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[31] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
M3[32] VB VB VB VB pfet_03v3 L=2u W=2u nf=1 m=1
.ends


* expanding   symbol:  DiffN_nfets.sym # of pins=6
** sym_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/DiffN_nfets.sym
** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/DiffN_nfets.sch
.subckt DiffN_nfets D1 D2 G1 G2 S B
*.PININFO D1:B D2:B G1:B G2:B S:B B:B
M1 D1 G1 net1 B nfet_03v3 L=2u W=2u nf=1 m=1
M2 D2 G2 net5 B nfet_03v3 L=2u W=2u nf=1 m=1
M3 D1 G1 net2 B nfet_03v3 L=2u W=2u nf=1 m=1
M4 D1 G1 net3 B nfet_03v3 L=2u W=2u nf=1 m=1
M5 D1 G1 net4 B nfet_03v3 L=2u W=2u nf=1 m=1
M6 net1 G1 S B nfet_03v3 L=2u W=2u nf=1 m=1
M7 net2 G1 S B nfet_03v3 L=2u W=2u nf=1 m=1
M8 net3 G1 S B nfet_03v3 L=2u W=2u nf=1 m=1
M9 net4 G1 S B nfet_03v3 L=2u W=2u nf=1 m=1
M10 D2 G2 net6 B nfet_03v3 L=2u W=2u nf=1 m=1
M11 D2 G2 net7 B nfet_03v3 L=2u W=2u nf=1 m=1
M12 D2 G2 net8 B nfet_03v3 L=2u W=2u nf=1 m=1
M13 net5 G2 S B nfet_03v3 L=2u W=2u nf=1 m=1
M14 net6 G2 S B nfet_03v3 L=2u W=2u nf=1 m=1
M15 net7 G2 S B nfet_03v3 L=2u W=2u nf=1 m=1
M16 net8 G2 S B nfet_03v3 L=2u W=2u nf=1 m=1
M17[1] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[2] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[3] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[4] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[5] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[6] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[7] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[8] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[9] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[10] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[11] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[12] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[13] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[14] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[15] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[16] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[17] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[18] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[19] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[20] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[21] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[22] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[23] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[24] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[25] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[26] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[27] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[28] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[29] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[30] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[31] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M17[32] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
.ends


* expanding   symbol:  DiffN_pfets.sym # of pins=5
** sym_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/DiffN_pfets.sym
** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/DiffN_pfets.sch
.subckt DiffN_pfets D1 D2 G S B
*.PININFO D1:B D2:B G:B S:B B:B
M1 net4 G S B pfet_03v3 L=2u W=2u nf=1 m=1
M2 net5 G S B pfet_03v3 L=2u W=2u nf=1 m=1
M3 net3 G S B pfet_03v3 L=2u W=2u nf=1 m=1
M4 net2 G S B pfet_03v3 L=2u W=2u nf=1 m=1
M5 net1 G S B pfet_03v3 L=2u W=2u nf=1 m=1
M6 D1 G net4 B pfet_03v3 L=2u W=2u nf=1 m=1
M7 D1 G net3 B pfet_03v3 L=2u W=2u nf=1 m=1
M8 D1 G net2 B pfet_03v3 L=2u W=2u nf=1 m=1
M9 D1 G net1 B pfet_03v3 L=2u W=2u nf=1 m=1
M10 net6 G S B pfet_03v3 L=2u W=2u nf=1 m=1
M11 net7 G S B pfet_03v3 L=2u W=2u nf=1 m=1
M12 net8 G S B pfet_03v3 L=2u W=2u nf=1 m=1
M13 D2 G net5 B pfet_03v3 L=2u W=2u nf=1 m=1
M14 D2 G net6 B pfet_03v3 L=2u W=2u nf=1 m=1
M15 D2 G net7 B pfet_03v3 L=2u W=2u nf=1 m=1
M16 D2 G net8 B pfet_03v3 L=2u W=2u nf=1 m=1
M17[1] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[2] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[3] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[4] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[5] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[6] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[7] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[8] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[9] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[10] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[11] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[12] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[13] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[14] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[15] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[16] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[17] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[18] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[19] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[20] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[21] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[22] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[23] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[24] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[25] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[26] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[27] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[28] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[29] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[30] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[31] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M17[32] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
.ends


* expanding   symbol:  DiffP_nfets.sym # of pins=5
** sym_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/DiffP_nfets.sym
** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/DiffP_nfets.sch
.subckt DiffP_nfets D1 D2 G S B
*.PININFO D1:B D2:B G:B S:B B:B
M1 D1 G net4 B nfet_03v3 L=2u W=2u nf=1 m=1
M2 D2 G net5 B nfet_03v3 L=2u W=2u nf=1 m=1
M5 D1 G net3 B nfet_03v3 L=2u W=2u nf=1 m=1
M6 D1 G net2 B nfet_03v3 L=2u W=2u nf=1 m=1
M7 D1 G net1 B nfet_03v3 L=2u W=2u nf=1 m=1
M8 net4 G S B nfet_03v3 L=2u W=2u nf=1 m=1
M9 net3 G S B nfet_03v3 L=2u W=2u nf=1 m=1
M10 net2 G S B nfet_03v3 L=2u W=2u nf=1 m=1
M11 net1 G S B nfet_03v3 L=2u W=2u nf=1 m=1
M12 D2 G net6 B nfet_03v3 L=2u W=2u nf=1 m=1
M13 D2 G net7 B nfet_03v3 L=2u W=2u nf=1 m=1
M14 D2 G net8 B nfet_03v3 L=2u W=2u nf=1 m=1
M15 net5 G S B nfet_03v3 L=2u W=2u nf=1 m=1
M16 net6 G S B nfet_03v3 L=2u W=2u nf=1 m=1
M17 net7 G S B nfet_03v3 L=2u W=2u nf=1 m=1
M18 net8 G S B nfet_03v3 L=2u W=2u nf=1 m=1
M3[1] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[2] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[3] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[4] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[5] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[6] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[7] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[8] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[9] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[10] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[11] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[12] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[13] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[14] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[15] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[16] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[17] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[18] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[19] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[20] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[21] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[22] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[23] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[24] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[25] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[26] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[27] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[28] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[29] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[30] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[31] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[32] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
.ends


* expanding   symbol:  DiffP_pfets.sym # of pins=6
** sym_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/DiffP_pfets.sym
** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/PseudoResistor/DiffP_pfets.sch
.subckt DiffP_pfets D1 D2 G1 G2 S B
*.PININFO D1:B D2:B G1:B G2:B S:B B:B
M1 net4 G1 S B pfet_03v3 L=2u W=2u nf=1 m=1
M2 net5 G2 S B pfet_03v3 L=2u W=2u nf=1 m=1
M5 net3 G1 S B pfet_03v3 L=2u W=2u nf=1 m=1
M6 net2 G1 S B pfet_03v3 L=2u W=2u nf=1 m=1
M7 net1 G1 S B pfet_03v3 L=2u W=2u nf=1 m=1
M8 D1 G1 net4 B pfet_03v3 L=2u W=2u nf=1 m=1
M9 D1 G1 net3 B pfet_03v3 L=2u W=2u nf=1 m=1
M10 D1 G1 net2 B pfet_03v3 L=2u W=2u nf=1 m=1
M11 D1 G1 net1 B pfet_03v3 L=2u W=2u nf=1 m=1
M12 net6 G2 S B pfet_03v3 L=2u W=2u nf=1 m=1
M15 D2 G2 net5 B pfet_03v3 L=2u W=2u nf=1 m=1
M16 D2 G2 net6 B pfet_03v3 L=2u W=2u nf=1 m=1
M19 net7 G2 S B pfet_03v3 L=2u W=2u nf=1 m=1
M20 net8 G2 S B pfet_03v3 L=2u W=2u nf=1 m=1
M21 D2 G2 net7 B pfet_03v3 L=2u W=2u nf=1 m=1
M22 D2 G2 net8 B pfet_03v3 L=2u W=2u nf=1 m=1
M3[1] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[2] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[3] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[4] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[5] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[6] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[7] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[8] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[9] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[10] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[11] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[12] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[13] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[14] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[15] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[16] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[17] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[18] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[19] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[20] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[21] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[22] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[23] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[24] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[25] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[26] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[27] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[28] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[29] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[30] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[31] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[32] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
.ends

.end
