* Extracted by KLayout with GF180MCU LVS runset on : 28/03/2024 15:38

.SUBCKT FC_top AVSS IREF AVDD VOUT VP VN
M$1 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$4 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$5 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$6 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$7 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$8 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$9 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$10 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$11 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$12 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$13 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$14 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$15 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P PS=3.7U
+ PD=2.04U
M$16 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P PS=2.04U
+ PD=2.04U
M$17 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P PS=2.04U
+ PD=3.7U
M$18 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$19 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$20 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$21 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$22 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$23 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$24 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$25 AVDD IREF \$56 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$26 \$56 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$27 AVDD IREF \$56 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$28 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$29 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$30 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$31 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$32 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$33 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$34 \$144 \$24 \$143 AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P PS=3.7U
+ PD=2.04U
M$35 \$145 \$24 \$144 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P PS=2.04U
+ PD=2.04U
M$36 AVDD \$24 \$145 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P PS=2.04U
+ PD=3.7U
M$37 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$38 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$39 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$40 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$41 \$164 \$24 \$143 AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P PS=3.7U
+ PD=2.04U
M$42 \$165 \$24 \$164 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P PS=2.04U
+ PD=2.04U
M$43 \$166 \$24 \$165 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P PS=2.04U
+ PD=3.7U
M$44 \$179 \$24 \$178 AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P PS=3.7U
+ PD=2.04U
M$45 \$180 \$24 \$179 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P PS=2.04U
+ PD=2.04U
M$46 \$166 \$24 \$180 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P PS=2.04U
+ PD=3.7U
M$47 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$48 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$49 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$50 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$51 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$52 AVDD IREF \$56 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$53 \$56 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$54 AVDD IREF \$56 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$55 \$56 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$56 \$30 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$57 AVDD IREF \$30 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$58 \$30 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$59 AVDD IREF \$56 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$60 \$56 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$61 AVDD IREF \$56 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$62 \$56 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$63 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$64 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$65 AVDD IREF \$30 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$66 \$30 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$67 AVDD IREF \$30 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$68 \$30 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$69 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$70 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$71 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$72 AVDD IREF \$30 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$73 \$30 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$74 AVDD IREF \$30 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$75 \$30 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$76 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$77 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$78 \$192 \$24 \$178 AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P PS=3.7U
+ PD=2.04U
M$79 \$193 \$24 \$192 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P PS=2.04U
+ PD=2.04U
M$80 \$194 \$24 \$193 AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P PS=2.04U
+ PD=3.7U
M$81 \$24 \$24 \$194 AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$82 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$83 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$84 AVDD IREF \$30 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$85 \$30 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$86 AVDD IREF \$30 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$87 \$30 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$88 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$89 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$90 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$91 AVDD IREF \$30 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$92 \$30 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$93 AVDD IREF \$30 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$94 \$30 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$95 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$96 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U PD=3.7U
M$97 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.504P PS=3.7U
+ PD=2.04U
M$98 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.504P PS=2.04U
+ PD=2.04U
M$99 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.504P AD=0.78P PS=2.04U
+ PD=3.7U
M$100 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$101 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=1.2U AS=0.78P AD=0.78P PS=3.7U
+ PD=3.7U
M$102 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$103 AVDD IREF \$56 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$104 \$56 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$105 AVDD IREF \$56 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$106 \$56 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$107 AVDD IREF \$30 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$108 \$30 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$109 AVDD IREF \$30 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$110 AVDD IREF \$56 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$111 \$56 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$112 AVDD IREF \$56 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$113 \$56 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$114 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$115 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$116 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$117 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$118 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$119 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$120 \$56 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$121 AVDD IREF \$56 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$122 \$56 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$123 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$124 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$125 AVDD IREF IREF AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$126 IREF IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$127 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$128 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$129 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$130 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$131 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$132 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$133 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$134 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$135 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$136 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$137 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$138 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$139 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$140 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$141 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$142 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$143 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$144 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$145 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$146 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$147 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$148 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$149 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$150 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$151 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$152 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$153 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$154 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$155 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$156 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$157 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$158 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$159 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$160 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$161 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$162 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$163 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$164 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$165 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$166 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$167 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$168 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$169 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$170 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$171 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$172 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$173 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$174 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$175 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$176 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$177 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$178 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$179 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$180 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$181 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$182 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$183 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$184 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$185 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$186 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$187 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$188 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$189 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$190 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$191 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$192 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$193 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$194 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$195 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$196 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$197 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$198 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$199 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$200 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$201 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$202 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$203 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$204 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$205 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$206 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$207 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$208 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$209 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$210 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$211 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$212 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$213 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$214 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$215 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$216 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$217 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$218 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$219 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$220 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$221 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$222 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$223 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$224 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$225 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$226 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$227 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$228 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$229 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$230 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$231 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$232 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$233 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$234 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$235 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$236 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$237 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$238 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$239 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$240 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$241 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$242 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$243 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$244 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$245 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$246 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$247 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$248 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$249 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$250 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$251 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$252 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$253 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$254 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$255 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$256 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$257 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$258 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$259 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$260 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$261 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$262 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$263 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$264 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$265 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$266 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$267 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$268 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$269 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$270 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$271 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$272 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$273 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$274 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$275 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$276 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$277 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$278 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$279 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$280 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$281 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$282 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$283 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$284 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$285 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$286 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$287 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$288 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$289 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$290 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$291 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$292 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$293 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$294 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$295 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$296 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$297 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$298 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$299 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$300 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$301 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$302 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$303 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$304 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$305 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$306 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$307 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$308 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$309 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$310 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$311 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$312 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$313 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$314 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$315 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$316 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$317 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$318 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$319 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$320 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$321 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$322 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$323 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$324 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$325 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$326 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$327 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$328 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$329 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$330 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$331 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$332 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$333 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$334 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$335 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$336 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$337 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$338 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$339 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$340 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$341 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$342 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$343 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$344 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$345 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$346 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$347 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$348 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$349 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$350 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$351 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$352 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$353 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$354 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$355 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$356 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$357 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$358 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$359 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$360 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$361 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$362 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$363 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$364 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$365 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$366 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$367 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$368 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$369 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$370 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$371 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$372 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$373 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$374 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$375 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$376 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$377 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$378 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$379 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$380 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$381 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$382 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$383 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$384 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$385 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$386 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$387 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$388 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$389 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$390 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$391 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$392 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$393 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$394 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$395 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$396 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$397 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$398 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$399 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$400 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$401 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$402 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$403 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$404 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$405 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$406 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$407 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$408 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$409 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$410 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$411 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$412 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$413 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$414 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$415 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$416 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$417 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$418 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$419 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$420 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$421 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$422 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$423 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$424 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$425 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$426 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$427 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$428 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$429 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$430 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$431 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$432 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$433 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$434 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$435 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$436 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$437 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$438 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$439 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$440 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$441 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$442 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$443 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$444 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$445 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$446 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$447 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$448 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$449 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$450 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$451 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$452 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$453 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$454 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$455 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$456 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$457 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$458 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$459 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$460 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$461 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$462 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$463 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$464 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$465 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$466 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$467 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$468 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$469 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$470 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$471 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$472 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$473 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$474 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$475 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$476 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$477 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$478 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$479 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$480 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$481 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$482 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$483 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$484 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$485 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$486 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$487 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$488 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$489 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$490 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$491 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$492 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$493 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$494 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$495 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$496 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$497 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$498 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$499 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$500 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$501 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$502 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$503 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$504 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$505 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$506 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$507 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$508 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$509 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$510 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$511 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$512 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$513 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$514 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$515 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$516 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$517 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$518 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$519 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$520 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$521 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$522 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$523 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$524 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$525 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$526 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$527 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$528 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$529 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$530 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$531 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$532 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$533 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$534 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$535 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$536 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$537 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$538 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$539 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$540 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$541 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$542 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$543 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$544 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$545 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$546 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$547 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$548 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$549 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$550 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$551 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$552 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$553 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$554 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$555 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$556 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$557 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$558 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$559 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$560 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$561 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$562 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$563 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$564 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$565 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$566 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$567 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$568 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$569 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$570 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$571 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$572 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$573 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$574 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$575 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$576 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$577 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$578 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$579 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$580 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$581 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$582 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$583 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$584 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$585 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$586 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$587 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$588 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$589 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$590 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$591 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$592 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$593 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$594 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$595 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$596 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$597 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$598 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$599 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$600 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$601 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$602 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$603 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$604 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$605 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$606 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$607 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$608 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$609 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$610 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$611 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$612 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$613 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$614 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$615 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$616 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$617 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$618 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$619 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$620 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$621 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$622 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$623 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$624 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$625 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$626 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$627 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$628 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$629 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$630 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$631 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$632 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$633 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$634 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$635 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$636 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$637 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$638 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$639 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$640 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$641 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$642 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$643 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$644 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$645 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$646 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$647 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$648 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$649 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$650 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$651 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$652 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$653 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$654 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$655 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$656 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$657 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$658 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$659 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$660 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$661 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$662 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$663 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$664 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$665 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$666 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$667 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$668 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$669 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$670 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$671 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$672 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$673 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$674 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$675 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$676 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$677 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$678 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$679 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$680 \$331 VN \$15 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$681 \$15 VN \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$682 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$683 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$684 \$331 VP \$14 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U PD=2.84U
M$685 \$14 VP \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$686 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$687 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$688 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$689 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$690 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$691 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$692 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$693 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$694 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$695 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$696 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$697 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$698 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$699 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$700 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$701 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$702 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$703 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$704 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$705 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$706 \$326 \$24 VOUT AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$707 VOUT \$24 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$708 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$709 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$710 \$332 \$24 \$211 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$711 \$211 \$24 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$712 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$713 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$714 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$715 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$716 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$717 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$718 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$719 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$720 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$721 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$722 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$723 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$724 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$725 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$726 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$727 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$728 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$729 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$730 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$731 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$732 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$733 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$734 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$735 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$736 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$737 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$738 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$739 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$740 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$741 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$742 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$743 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$744 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$745 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$746 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$747 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$748 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$749 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$750 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$751 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$752 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$753 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$754 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$755 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$756 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$757 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$758 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$759 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$760 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$761 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$762 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$763 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$764 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$765 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$766 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$767 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$768 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$769 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$770 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$771 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$772 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$773 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$774 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$775 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$776 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$777 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$778 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$779 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$780 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$781 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$782 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$783 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$784 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$785 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$786 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$787 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$788 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$789 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$790 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$791 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$792 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$793 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$794 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$795 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$796 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$797 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$798 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$799 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$800 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$801 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$802 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$803 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$804 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$805 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$806 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$807 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$808 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$809 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$810 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$811 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$812 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$813 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$814 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$815 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$816 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$817 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$818 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$819 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$820 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$821 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$822 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$823 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$824 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$825 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$826 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$827 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$828 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$829 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$830 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$831 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$832 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$833 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$834 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$835 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$836 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$837 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$838 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$839 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$840 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$841 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$842 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$843 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$844 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$845 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$846 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$847 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$848 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$849 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$850 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$851 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$852 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$853 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$854 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$855 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$856 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$857 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$858 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$859 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$860 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$861 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$862 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$863 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$864 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$865 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$866 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$867 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$868 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$869 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$870 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$871 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$872 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$873 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$874 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$875 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$876 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$877 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$878 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$879 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$880 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$881 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$882 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$883 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$884 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$885 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$886 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$887 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$888 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$889 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$890 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$891 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$892 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$893 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$894 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$895 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$896 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$897 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$898 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$899 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$900 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$901 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$902 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$903 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$904 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$905 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$906 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$907 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$908 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$909 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$910 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$911 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$912 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$913 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$914 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$915 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$916 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$917 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$918 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$919 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$920 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$921 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$922 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$923 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$924 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$925 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$926 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$927 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$928 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$929 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$930 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$931 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$932 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$933 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$934 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$935 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$936 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$937 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$938 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$939 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$940 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$941 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$942 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$943 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$944 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$945 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$946 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$947 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$948 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$949 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$950 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$951 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$952 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$953 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$954 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$955 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$956 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$957 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$958 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$959 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$960 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$961 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$962 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$963 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$964 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$965 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$966 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$967 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$968 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$969 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$970 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$971 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$972 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$973 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$974 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$975 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$976 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$977 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$978 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$979 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$980 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$981 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$982 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$983 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$984 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$985 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$986 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$987 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$988 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$989 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$990 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$991 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$992 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$993 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$994 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$995 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$996 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$997 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$998 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$999 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1000 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1001 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1002 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1003 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1004 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1005 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1006 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1007 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1008 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1009 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1010 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1011 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1012 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1013 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1014 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1015 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1016 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1017 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1018 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1019 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1020 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1021 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1022 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1023 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1024 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1025 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1026 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1027 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1028 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1029 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1030 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1031 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1032 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1033 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1034 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1035 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1036 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1037 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1038 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1039 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1040 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1041 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1042 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1043 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1044 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1045 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1046 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1047 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1048 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1049 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1050 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1051 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1052 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1053 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1054 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1055 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1056 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1057 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1058 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1059 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1060 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1061 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1062 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1063 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1064 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1065 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1066 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1067 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1068 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1069 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1070 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1071 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1072 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1073 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1074 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1075 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1076 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1077 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1078 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1079 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1080 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1081 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1082 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1083 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1084 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1085 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1086 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1087 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1088 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1089 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1090 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1091 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1092 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1093 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1094 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1095 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1096 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1097 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1098 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1099 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1100 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1101 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1102 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1103 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1104 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1105 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1106 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1107 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1108 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1109 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1110 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1111 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1112 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1113 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1114 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1115 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1116 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1117 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1118 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1119 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1120 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1121 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1122 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1123 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1124 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1125 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1126 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1127 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1128 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1129 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1130 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1131 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1132 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1133 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1134 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1135 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1136 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1137 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1138 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1139 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1140 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1141 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1142 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1143 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1144 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1145 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1146 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1147 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1148 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1149 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1150 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1151 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1152 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1153 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1154 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1155 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1156 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1157 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1158 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1159 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1160 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1161 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1162 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1163 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1164 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1165 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1166 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1167 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1168 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1169 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1170 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1171 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1172 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1173 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1174 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1175 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1176 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1177 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1178 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1179 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1180 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1181 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1182 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1183 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1184 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1185 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1186 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1187 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1188 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1189 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1190 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1191 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1192 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1193 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1194 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1195 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1196 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1197 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1198 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1199 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1200 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1201 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1202 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1203 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1204 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1205 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1206 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1207 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1208 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1209 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1210 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1211 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1212 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1213 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1214 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1215 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1216 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1217 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1218 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1219 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1220 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1221 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1222 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1223 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1224 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1225 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1226 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1227 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1228 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1229 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1230 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1231 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1232 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1233 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1234 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1235 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1236 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1237 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1238 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1239 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1240 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1241 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1242 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1243 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1244 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1245 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1246 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1247 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1248 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1249 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1250 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1251 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1252 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1253 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1254 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1255 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1256 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1257 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1258 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1259 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1260 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1261 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1262 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1263 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1264 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1265 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1266 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1267 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1268 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1269 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1270 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1271 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1272 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1273 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1274 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1275 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1276 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1277 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1278 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1279 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1280 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1281 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1282 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1283 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1284 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1285 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1286 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1287 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1288 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1289 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1290 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1291 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1292 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1293 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1294 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1295 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1296 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1297 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1298 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1299 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1300 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1301 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1302 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1303 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1304 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1305 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1306 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1307 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1308 AVDD IREF \$331 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1309 \$331 IREF AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1310 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1311 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1312 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1313 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1314 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1315 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1316 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1317 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1318 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1319 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1320 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1321 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1322 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1323 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1324 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1325 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1326 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1327 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1328 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1329 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1330 AVDD \$211 \$326 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1331 \$326 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1332 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U
+ PD=2.84U
M$1333 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1334 AVDD \$211 \$332 AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1335 \$332 \$211 AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U
+ PD=5.3U
M$1336 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1337 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1338 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1339 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1340 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1341 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1342 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1343 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1344 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1345 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1346 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1347 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1348 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1349 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1350 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1351 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1352 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1353 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1354 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1355 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1356 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1357 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1358 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1359 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1360 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1361 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1362 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1363 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1364 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1365 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1366 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1367 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1368 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1369 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1370 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1371 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1372 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1373 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1374 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1375 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1376 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1377 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1378 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1379 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1380 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1381 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1382 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1383 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1384 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$1385 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1386 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=0.84P PS=2.84U
+ PD=2.84U
M$1387 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$1388 AVDD AVDD AVDD AVDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$1389 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1390 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1391 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1392 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1393 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1394 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1395 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1396 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1397 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1398 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1399 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1400 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1401 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1402 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1403 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1404 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1405 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1406 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1407 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1408 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1409 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1410 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1411 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P
+ PS=5.72U PD=5.72U
M$1412 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$1413 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$1414 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$1415 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$1416 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P
+ PS=5.72U PD=5.72U
M$1417 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1418 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1419 AVSS \$30 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1420 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1421 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1422 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1423 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1424 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1425 AVSS \$30 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1426 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1427 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1428 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1429 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1430 AVSS \$30 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1431 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1432 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1433 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1434 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1435 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1436 AVSS \$30 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1437 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1438 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1439 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P
+ PS=5.72U PD=5.72U
M$1440 AVSS \$30 \$30 AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$1441 \$30 \$30 AVSS AVSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$1442 AVSS \$30 \$24 AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$1443 \$24 \$30 AVSS AVSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$1444 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P
+ PS=5.72U PD=5.72U
M$1445 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$1446 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P PS=3.62U
+ PD=2U
M$1447 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U
+ PD=3.62U
M$1448 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$1449 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1450 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1451 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1452 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1453 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1454 AVSS \$30 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1455 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1456 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1457 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1458 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1459 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1460 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1461 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1462 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1463 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1464 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1465 AVSS \$30 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1466 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1467 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1468 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1469 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1470 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1471 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P
+ PS=5.72U PD=5.72U
M$1472 AVSS \$30 \$24 AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$1473 \$24 \$30 AVSS AVSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$1474 AVSS \$30 \$30 AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$1475 \$30 \$30 AVSS AVSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$1476 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P
+ PS=5.72U PD=5.72U
M$1477 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$1478 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$1479 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$1480 \$73 \$56 \$48 AVSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P PS=3.62U
+ PD=2U
M$1481 \$74 \$56 \$73 AVSS nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U
+ PD=3.62U
M$1482 \$89 \$56 \$56 AVSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P PS=3.62U
+ PD=2U
M$1483 \$74 \$56 \$89 AVSS nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U
+ PD=3.62U
M$1484 \$49 \$56 \$48 AVSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P PS=3.62U
+ PD=2U
M$1485 AVSS \$56 \$49 AVSS nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U
+ PD=3.62U
M$1486 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$1487 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$1488 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$1489 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1490 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1491 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1492 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1493 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1494 AVSS \$30 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1495 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1496 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1497 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1498 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1499 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1500 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1501 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1502 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1503 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1504 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1505 AVSS \$30 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1506 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1507 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1508 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1509 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1510 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1511 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P
+ PS=5.72U PD=5.72U
M$1512 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$1513 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$1514 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=0.9P PS=5.72U
+ PD=3.05U
M$1515 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=0.9P AD=1.3725P PS=3.05U
+ PD=5.72U
M$1516 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2.25U AS=1.3725P AD=1.3725P
+ PS=5.72U PD=5.72U
M$1517 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$1518 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.48P PS=3.62U
+ PD=2U
M$1519 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=1.2U AS=0.48P AD=0.732P PS=2U
+ PD=3.62U
M$1520 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=1.2U AS=0.732P AD=0.732P PS=3.62U
+ PD=3.62U
M$1521 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1522 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1523 AVSS \$30 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1524 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1525 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1526 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1527 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1528 AVSS \$30 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1529 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1530 AVSS \$30 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1531 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1532 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1533 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1534 AVSS \$30 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1535 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1536 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1537 AVSS \$30 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1538 \$15 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1539 AVSS \$30 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1540 \$14 \$30 AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1541 AVSS \$30 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1542 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1543 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1544 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1545 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1546 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1547 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1548 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1549 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1550 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1551 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1552 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1553 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1554 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1555 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1556 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1557 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1558 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1559 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1560 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1561 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1562 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1563 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1564 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1565 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1566 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1567 \$211 \$56 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1568 \$14 \$56 \$211 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1569 \$211 \$56 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1570 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1571 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1572 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1573 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1574 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1575 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1576 \$15 \$56 VOUT AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1577 VOUT \$56 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1578 \$15 \$56 VOUT AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1579 \$211 \$56 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1580 \$14 \$56 \$211 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1581 \$211 \$56 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1582 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1583 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1584 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1585 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1586 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1587 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1588 VOUT \$56 \$15 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1589 \$15 \$56 VOUT AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1590 VOUT \$56 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1591 \$211 \$56 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1592 \$14 \$56 \$211 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1593 \$211 \$56 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1594 \$15 \$56 VOUT AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1595 VOUT \$56 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1596 \$15 \$56 VOUT AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1597 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1598 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1599 VOUT \$56 \$15 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1600 \$15 \$56 VOUT AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1601 VOUT \$56 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1602 \$211 \$56 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1603 \$14 \$56 \$211 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1604 \$211 \$56 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1605 \$15 \$56 VOUT AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1606 VOUT \$56 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1607 \$15 \$56 VOUT AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1608 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1609 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1610 \$211 \$56 \$14 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1611 \$14 \$56 \$211 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1612 \$211 \$56 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1613 VOUT \$56 \$15 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1614 \$15 \$56 VOUT AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1615 VOUT \$56 \$15 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1616 \$14 \$56 \$211 AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U
+ PD=2.8U
M$1617 \$211 \$56 \$14 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1618 \$14 \$56 \$211 AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U
+ PD=5.22U
M$1619 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1620 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$1621 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1622 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1623 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1624 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1625 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1626 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1627 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$1628 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$1629 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$1630 AVSS AVSS AVSS AVSS nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
.ENDS FC_top
