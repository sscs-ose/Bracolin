* Extracted by KLayout with GF180MCU LVS runset on : 10/04/2024 20:16

.SUBCKT overvoltageProtection GND iref Load vdd vfb vref PowerGate
M$1 \$5 \$6 vfb vdd pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$2 vfb \$6 \$5 vdd pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$3 \$6 \$6 vref vdd pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$4 vref \$6 \$6 vdd pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$5 vdd \$32 \$32 vdd pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$6 PowerGate \$34 vdd vdd pfet_03v3 L=1U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$7 \$5 \$6 vfb vdd pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$8 vfb \$6 \$5 vdd pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$9 \$6 \$6 vref vdd pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$10 vref \$6 \$6 vdd pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$11 PowerGate \$34 vdd vdd pfet_03v3 L=1U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$12 vdd \$34 \$34 vdd pfet_03v3 L=5U W=1U AS=2.12P AD=2.12P PS=6.24U PD=6.24U
M$13 \$5 \$6 vfb vdd pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$14 vfb \$6 \$5 vdd pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$15 \$6 \$6 vref vdd pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$16 vref \$6 \$6 vdd pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$17 vdd \$32 \$29 vdd pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$18 PowerGate \$34 vdd vdd pfet_03v3 L=1U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$19 \$5 \$6 vfb vdd pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$20 vfb \$6 \$5 vdd pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$21 \$6 \$6 vref vdd pfet_03v3 L=2U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$22 vref \$6 \$6 vdd pfet_03v3 L=2U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$23 vdd \$32 \$29 vdd pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$24 PowerGate \$34 vdd vdd pfet_03v3 L=1U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$25 \$7 \$5 GND GND nfet_03v3 L=20U W=0.5U AS=0.305P AD=0.305P PS=2.22U
+ PD=2.22U
M$26 \$7 \$5 \$5 GND nfet_03v3 L=20U W=0.5U AS=0.305P AD=0.305P PS=2.22U
+ PD=2.22U
M$27 \$6 iref GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=0.52P PS=5.22U PD=2.52U
M$28 GND iref \$6 GND nfet_03v3 L=2U W=2U AS=0.52P AD=1.22P PS=2.52U PD=5.22U
M$29 \$5 iref GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=0.52P PS=5.22U PD=2.52U
M$30 GND iref \$5 GND nfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$31 \$5 iref GND GND nfet_03v3 L=2U W=2U AS=0.52P AD=1.22P PS=2.52U PD=5.22U
M$32 \$8 iref GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=0.52P PS=5.22U PD=2.52U
M$33 GND iref \$8 GND nfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$34 \$8 iref GND GND nfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$35 GND iref \$8 GND nfet_03v3 L=2U W=2U AS=0.52P AD=1.22P PS=2.52U PD=5.22U
M$36 GND \$29 \$33 GND nfet_03v3 L=20U W=0.5U AS=0.305P AD=0.305P PS=2.22U
+ PD=2.22U
M$37 \$29 \$29 \$33 GND nfet_03v3 L=20U W=0.5U AS=0.305P AD=0.305P PS=2.22U
+ PD=2.22U
M$38 \$32 iref GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$39 \$8 \$5 \$34 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$40 vdd \$29 \$8 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$41 Load \$5 GND GND nfet_03v3 L=0.45U W=20U AS=12.2P AD=5.2P PS=41.22U
+ PD=20.52U
M$42 GND \$5 Load GND nfet_03v3 L=0.45U W=20U AS=5.2P AD=5.2P PS=20.52U
+ PD=20.52U
M$43 Load \$5 GND GND nfet_03v3 L=0.45U W=20U AS=5.2P AD=5.2P PS=20.52U
+ PD=20.52U
M$44 GND \$5 Load GND nfet_03v3 L=0.45U W=20U AS=5.2P AD=5.2P PS=20.52U
+ PD=20.52U
M$45 Load \$5 GND GND nfet_03v3 L=0.45U W=20U AS=5.2P AD=5.2P PS=20.52U
+ PD=20.52U
M$46 GND \$5 Load GND nfet_03v3 L=0.45U W=20U AS=5.2P AD=5.2P PS=20.52U
+ PD=20.52U
M$47 Load \$5 GND GND nfet_03v3 L=0.45U W=20U AS=5.2P AD=5.2P PS=20.52U
+ PD=20.52U
M$48 GND \$5 Load GND nfet_03v3 L=0.45U W=20U AS=5.2P AD=5.2P PS=20.52U
+ PD=20.52U
M$49 Load \$5 GND GND nfet_03v3 L=0.45U W=20U AS=5.2P AD=5.2P PS=20.52U
+ PD=20.52U
M$50 GND \$5 Load GND nfet_03v3 L=0.45U W=20U AS=5.2P AD=5.2P PS=20.52U
+ PD=20.52U
M$51 Load \$5 GND GND nfet_03v3 L=0.45U W=20U AS=5.2P AD=5.2P PS=20.52U
+ PD=20.52U
M$52 GND \$5 Load GND nfet_03v3 L=0.45U W=20U AS=5.2P AD=5.2P PS=20.52U
+ PD=20.52U
M$53 Load \$5 GND GND nfet_03v3 L=0.45U W=20U AS=5.2P AD=5.2P PS=20.52U
+ PD=20.52U
M$54 GND \$5 Load GND nfet_03v3 L=0.45U W=20U AS=5.2P AD=5.2P PS=20.52U
+ PD=20.52U
M$55 Load \$5 GND GND nfet_03v3 L=0.45U W=20U AS=5.2P AD=5.2P PS=20.52U
+ PD=20.52U
M$56 GND \$5 Load GND nfet_03v3 L=0.45U W=20U AS=5.2P AD=12.2P PS=20.52U
+ PD=41.22U
.ENDS overvoltageProtection
