* NGSPICE file created from Filter_TOP.ext - technology: gf180mcuD

.subckt Filter_TOP IN_NEG IN_POS VCM VSS I1U VDD I1N IBNOUT OUT IBPOUT
X0 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6 a_100820_11614# a_57977_n12421# a_102796_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X7 a_31284_4481# a_30324_4421# a_30724_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X8 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X9 a_102756_12380# a_100820_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X10 a_36032_n36322# a_53829_n36382# a_55635_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X11 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X12 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X13 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X14 a_101350_10448# a_100820_10448# a_100820_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X15 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X16 a_38619_n2651# a_31953_n19727# a_38097_n2651# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X17 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X18 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X19 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X20 VDD a_31699_20742# a_35502_24538# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X21 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X22 a_43817_6405# a_41891_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X23 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X24 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X25 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X26 a_105365_n7865# a_71281_n8397# a_104527_n7865# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X27 VDD a_31699_20742# a_35502_25545# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X28 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X29 a_58851_n7138# a_50751_n19729# a_58329_n8035# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X30 a_53145_n19597# a_50751_n19729# a_52585_n19597# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X31 a_71864_n30339# a_65486_n36322# a_71342_n30339# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X32 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X33 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X34 a_106809_n17715# a_71281_n8397# a_106501_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X35 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X36 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X37 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X38 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X39 a_105933_n2435# a_71281_n8397# a_105365_n2435# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X40 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X41 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X42 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X43 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X44 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X45 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X46 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X47 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X48 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X49 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X50 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X51 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X52 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X53 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X54 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X55 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X56 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X57 VSS VSS VSS VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X58 a_31284_n30339# a_30324_n30399# a_30724_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X59 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X60 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X61 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X62 a_33249_35053# a_35502_24538# OUT VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X63 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X64 a_38097_n5342# a_100992_n29313# a_101392_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X65 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X66 a_101392_6405# a_100992_4421# a_100820_10448# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X67 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X68 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X69 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X70 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X71 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X72 a_100235_n15000# a_71281_n8397# a_99667_n15000# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X73 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X74 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X75 a_73302_13546# a_71496_10388# a_71342_4481# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X76 a_30724_6405# a_30324_4421# a_30152_10448# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X77 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X78 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X79 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X80 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X81 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X82 a_31831_n5342# a_32913_n8930# a_83725_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X83 a_45445_n18698# a_31953_n19727# a_44885_n17801# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X84 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X85 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X86 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X87 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X88 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X89 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X90 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X91 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X92 a_51711_n5344# a_50751_n19729# a_51151_n5344# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X93 a_66551_n17803# a_50751_n19729# a_66029_n18700# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X94 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X95 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X96 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X97 a_98829_n17715# a_71281_n8397# a_98299_n16810# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X98 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X99 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X100 a_73302_11614# a_71496_10388# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X101 a_73268_n29181# a_65486_n36322# a_45445_n19595# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X102 a_90245_n6055# a_71281_n10073# a_60677_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X103 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X104 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X105 a_98829_n15000# a_71281_n8397# a_98299_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X106 a_51711_n14215# a_50751_n19729# a_51151_n14215# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X107 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X108 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X109 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X110 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X111 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X112 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X113 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X114 a_65486_n35156# a_65486_n35156# a_67422_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X115 a_60285_n2653# a_50751_n19729# a_59763_n3550# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X116 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X117 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X118 a_105365_n15000# a_71281_n8397# a_104527_n15000# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X119 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X120 a_106676_n30339# a_100820_n36322# a_108602_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X121 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X122 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X123 a_40613_n8930# a_31953_n19727# a_40053_n8930# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X124 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X125 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X126 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X127 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X128 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X129 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X130 a_110225_n1530# a_71281_n8397# a_109695_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X131 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X132 a_88271_n3340# a_71281_n10073# a_87433_n3340# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X133 VDD a_83153_11614# a_90935_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X134 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X135 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X136 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X137 a_114516_10448# a_86903_n14095# a_89715_n17715# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X138 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X139 a_39179_n8033# a_31953_n19727# a_38619_n8033# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X140 VDD a_31699_20742# a_35502_25545# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X141 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X142 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X143 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X144 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X145 a_84547_n15000# a_71281_n10073# a_83709_n14095# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X146 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X147 a_100235_n20430# a_71281_n8397# a_99667_n20430# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X148 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X149 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X150 VDD a_65486_n35156# a_66016_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X151 a_67111_n2653# a_50751_n19729# a_66551_n1756# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X152 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X153 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X154 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X155 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X156 a_54579_n4447# a_50751_n19729# a_54019_n4447# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X157 a_32353_n7136# a_31953_n19727# a_31831_n7136# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X158 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X159 VSS a_112559_4481# a_113081_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X160 a_30324_n30399# a_30152_n36322# a_36530_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X161 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X162 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X163 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X164 a_34347_n7136# a_31953_n19727# a_33787_n7136# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X165 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X166 a_48349_n35156# a_47819_n35156# a_47819_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X167 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X168 a_51711_n12421# a_83153_11614# a_89531_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X169 a_101350_n34390# a_100820_n35156# a_100820_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X170 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X171 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X172 a_77225_4481# a_77225_4481# a_79151_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X173 a_106676_4481# a_106830_10388# a_107230_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X174 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X175 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X176 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X177 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X178 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X179 a_57417_n8932# a_50751_n19729# a_56895_n8932# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X180 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X181 a_98829_n20430# a_71281_n8397# a_36032_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X182 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X183 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X184 VSS VSS VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X185 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X186 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X187 a_30152_n35156# a_30152_n35156# a_32088_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X188 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X189 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X190 a_89563_13546# a_89163_10388# a_89033_13546# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X191 a_67422_13546# a_65486_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X192 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X193 a_51151_n17803# a_50751_n19729# a_50629_n17803# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X194 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X195 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X196 a_43010_10448# a_36032_11614# a_42442_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X197 VSS VSS VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X198 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X199 a_48349_n33224# a_47819_n35156# a_47819_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X200 a_42047_n19595# a_31953_n19727# a_41487_n19595# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X201 a_30682_10448# a_30152_10448# a_30152_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X202 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X203 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X204 a_32088_n36322# a_30152_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X205 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X206 a_105365_n20430# a_71281_n8397# a_104527_n20430# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X207 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X208 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X209 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X210 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X211 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X212 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X213 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X214 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X215 VDD a_31699_20742# a_31699_20742# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X216 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X217 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X218 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X219 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X220 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X221 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X222 a_89563_11614# a_89163_10388# a_81205_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X223 a_67422_11614# a_65486_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X224 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X225 a_44885_n6239# a_31953_n19727# a_44363_n7136# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X226 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X227 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X228 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X229 a_43010_10448# a_36032_11614# a_42442_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X230 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X231 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X232 VSS a_89163_n36382# a_89563_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X233 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X234 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X235 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X236 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X237 a_47753_n15110# a_31953_n19727# a_47231_n16904# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X238 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X239 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X240 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X241 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X242 a_89531_6405# a_83153_11614# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X243 a_107339_n6055# a_71281_n8397# a_106809_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X244 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X245 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X246 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X247 a_52635_34067# a_35502_24538# a_33249_34067# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X248 VSS a_41891_n29181# a_42413_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X249 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X250 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X251 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X252 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X253 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X254 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X255 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X256 a_89407_n6960# a_71281_n10073# a_88839_n6960# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X257 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X258 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X259 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X260 a_89009_n27257# a_89163_n36382# a_89563_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X261 a_89033_13546# a_89163_10388# a_90969_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X262 a_31699_20742# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X263 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X264 a_53699_n36322# a_71496_n36382# a_73302_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X265 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X266 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X267 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X268 a_100235_n15905# a_71281_n8397# a_99667_n15905# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X269 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X270 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X271 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X272 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X273 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X274 a_40613_n14213# a_31953_n19727# a_40053_n14213# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X275 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X276 a_67462_n29181# a_45445_n19595# a_44363_n16007# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X277 a_31699_20742# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X278 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X279 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X280 a_94537_n9675# a_71281_n10073# a_93969_n9675# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X281 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X282 a_78344_n36322# a_71366_n35156# a_77776_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X283 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X284 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X285 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X286 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X287 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X288 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X289 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X290 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X291 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X292 a_39179_n19595# a_31953_n19727# a_38619_n19595# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X293 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X294 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X295 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X296 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X297 a_60845_n19597# a_50751_n19729# a_60285_n18700# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X298 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X299 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X300 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X301 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X302 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X303 a_71342_n30339# a_71496_n36382# a_71896_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X304 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X305 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X306 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X307 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X308 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X309 a_60285_n19597# a_50751_n19729# a_57977_n19597# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X310 a_98829_n15905# a_71281_n8397# a_98299_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X311 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X312 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X313 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X314 a_61484_4481# a_59558_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X315 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X316 a_54229_n35156# a_53829_n36382# a_53699_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X317 a_82573_n13190# a_71281_n10073# a_81735_n13190# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X318 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X319 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X320 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X321 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X322 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X323 a_105365_n15905# a_71281_n8397# a_104527_n15905# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X324 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X325 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X326 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X327 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X328 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X329 a_39179_n3548# a_31953_n19727# a_38619_n3548# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X330 a_94892_n29181# a_83325_n29313# a_96849_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X331 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X332 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X333 a_54579_n19597# a_50751_n19729# a_54019_n18700# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X334 a_32353_n15110# a_31953_n19727# a_31831_n15110# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X335 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X336 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X337 a_64243_n18700# a_50751_n19729# a_63683_n18700# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X338 a_54019_n4447# a_50751_n19729# a_53497_n6241# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X339 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X340 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X341 a_54229_n33224# a_53829_n36382# a_36032_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X342 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X343 a_88271_n2435# a_71281_n10073# a_87433_n2435# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X344 a_31699_19142# I1U a_30377_18342# VSS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X345 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X346 a_79151_n29181# a_77225_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X347 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X348 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X349 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X350 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X351 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X352 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X353 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X354 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X355 a_81735_n8770# a_71281_n10073# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X356 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X357 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X358 a_48313_n13316# a_31953_n19727# a_47753_n13316# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X359 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X360 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X361 a_63161_n5344# a_64243_n1756# a_66058_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X362 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X363 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X364 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X365 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X366 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X367 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X368 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X369 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X370 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X371 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X372 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X373 a_36008_4481# a_30152_11614# a_37934_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X374 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X375 a_58851_n14215# a_50751_n19729# a_58329_n14215# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X376 a_102796_n30339# a_100992_n29313# a_38097_n5342# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X377 a_96011_n36322# a_83325_n29313# a_95443_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X378 a_98829_n8770# a_71281_n8397# a_89033_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X379 a_83725_n29181# a_83325_n29313# a_83153_n35156# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X380 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X381 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X382 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X383 a_77747_7563# a_77225_4481# a_71496_10388# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X384 a_57977_n18700# a_50751_n19729# a_57417_n18700# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X385 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X386 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X387 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X388 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X389 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X390 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X391 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X392 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X393 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X394 a_108636_13546# a_106830_10388# a_106676_4481# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X395 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X396 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X397 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X398 a_57417_n16009# a_50751_n19729# a_56895_n16009# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X399 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X400 a_87433_n9675# a_71281_n10073# a_86903_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X401 a_33787_n17801# a_31953_n19727# a_33265_n18698# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X402 a_96011_n36322# a_83325_n29313# a_95443_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X403 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X404 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X405 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X406 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X407 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X408 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X409 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X410 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X411 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X412 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X413 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X414 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X415 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X416 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X417 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X418 a_108636_11614# a_106830_10388# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X419 a_64243_n8932# a_50751_n19729# a_63683_n8932# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X420 a_32128_7563# a_30324_4421# a_31284_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X421 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X422 a_66551_n4447# a_50751_n19729# a_66029_n6241# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X423 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X424 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X425 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X426 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X427 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X428 a_30152_n35156# a_30324_n29313# a_32128_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X429 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X430 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X431 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X432 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X433 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X434 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X435 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X436 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X437 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X438 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X439 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X440 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X441 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X442 a_48313_n7136# a_31953_n19727# a_47753_n7136# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X443 a_45706_22884# a_35922_19591# a_45138_22884# VDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X444 VSS a_112559_n29181# a_113081_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X445 a_107339_n6960# a_71281_n8397# a_106501_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X446 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X447 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X448 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X449 a_49755_12380# a_47819_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X450 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X451 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X452 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X453 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X454 a_43848_13546# a_30324_4421# a_43010_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X455 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X456 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X457 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X458 a_47819_n36322# a_39179_n19595# a_49795_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X459 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X460 a_93131_n8770# a_71281_n10073# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X461 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X462 VSS a_53829_n36382# a_54229_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X463 a_35502_25545# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X464 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X465 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X466 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X467 a_84017_n17715# a_83325_4421# a_95443_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X468 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X469 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X470 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X471 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X472 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X473 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X474 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X475 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X476 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X477 a_105365_n1530# a_71281_n8397# a_104527_n1530# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X478 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X479 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X480 a_43848_11614# a_30324_4421# a_43010_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X481 a_35502_25545# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X482 a_38619_n12419# a_31953_n19727# a_38097_n13316# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X483 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X484 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X485 a_105933_n15000# a_71281_n8397# a_105365_n15000# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X486 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X487 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X488 a_90935_n30339# a_83153_n36322# a_83325_n29313# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X489 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X490 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X491 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X492 a_47819_n36322# a_47819_n35156# a_49755_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X493 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X494 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X495 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X496 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X497 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X498 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X499 a_101392_n27257# a_100992_n29313# a_100820_n35156# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X500 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X501 a_41891_n29181# a_41891_n29181# a_43817_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X502 a_83153_10448# a_83153_10448# a_85089_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X503 a_47991_4421# a_47819_11614# a_54197_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X504 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X505 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X506 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X507 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X508 a_63683_n19597# a_50751_n19729# a_63161_n19597# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X509 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X510 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X511 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X512 a_106501_n6960# a_71281_n8397# a_105933_n6960# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X513 a_104527_n17715# a_71281_n8397# a_103997_n16810# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X514 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X515 a_58851_n1756# a_50751_n19729# a_57977_n5344# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X516 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X517 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X518 a_104527_n15000# a_71281_n8397# a_103997_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X519 a_47819_n36322# a_47819_n35156# a_49755_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X520 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X521 a_44885_n5342# a_31953_n19727# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X522 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X523 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X524 a_112199_n18620# a_71281_n8397# a_111631_n18620# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X525 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X526 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X527 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X528 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X529 OUT a_35502_24538# a_33249_35053# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X530 VDD a_47819_n35156# a_48349_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X531 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X532 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X533 a_104527_n8770# a_71281_n8397# a_103997_n8770# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X534 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X535 a_83153_10448# a_83153_10448# a_85089_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X536 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X537 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X538 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X539 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X540 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X541 a_111631_n9675# a_71281_n8397# a_111063_n9675# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X542 a_47753_n14213# a_31953_n19727# a_47231_n14213# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X543 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X544 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X545 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X546 a_46879_n19595# a_31953_n19727# a_46319_n18698# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X547 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X548 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X549 a_49795_4481# a_47991_5507# a_48951_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X550 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X551 a_83709_n19525# a_71281_n10073# a_83141_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X552 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X553 a_101350_n36322# a_100820_n35156# a_100820_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X554 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X555 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X556 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X557 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X558 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X559 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X560 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X561 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X562 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X563 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X564 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X565 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X566 a_42047_n4445# a_31953_n19727# a_41487_n4445# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X567 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X568 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X569 a_106830_10388# a_112559_4481# a_114485_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X570 VDD a_47819_n35156# a_48349_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X571 VSS a_41891_4481# a_42413_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X572 a_114485_n27257# a_112559_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X573 a_30152_n35156# a_30152_n35156# a_32088_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X574 a_54019_n17803# a_50751_n19729# a_53497_n18700# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X575 a_71896_n35156# a_71496_n36382# a_71366_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X576 a_81735_n7865# a_71281_n10073# a_81205_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X577 a_105933_n20430# a_71281_n8397# a_105365_n20430# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X578 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X579 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X580 a_59558_n29181# a_47991_n29313# a_61515_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X581 a_32913_n6239# a_31953_n19727# a_32353_n6239# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X582 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X583 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X584 a_54197_n30339# a_47819_n36322# a_53675_n30339# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X585 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X586 a_98829_n7865# a_71281_n8397# a_98299_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X587 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X588 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X589 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X590 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X591 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X592 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X593 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X594 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X595 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X596 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X597 VSS VSS VSS VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X598 a_71896_n33224# a_71496_n36382# a_53699_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X599 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X600 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X601 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X602 a_96849_n35156# a_89033_n35156# a_96011_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X603 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X604 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X605 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X606 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X607 a_84547_n6960# a_71281_n10073# a_83709_n6960# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X608 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X609 a_104527_n20430# a_71281_n8397# a_53699_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X610 a_93131_n19525# a_71281_n10073# a_92601_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X611 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X612 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X613 a_60677_n36322# a_53699_n35156# a_60109_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X614 a_56895_n16009# a_100992_4421# a_101392_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X615 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X616 a_88271_n19525# a_71281_n10073# a_87433_n19525# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X617 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X618 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X619 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X620 VDD a_30152_n35156# a_30682_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X621 VDD a_47819_n36322# a_55601_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X622 a_108602_n30339# a_100820_n36322# a_100992_n29313# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X623 a_45445_n14213# a_31953_n19727# a_44885_n13316# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X624 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X625 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X626 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X627 a_113081_6405# a_112559_4481# a_112559_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X628 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X629 a_96849_n33224# a_89033_n35156# a_96011_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X630 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X631 a_100235_n14095# a_71281_n8397# a_99667_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X632 a_65486_11614# a_64243_n1756# a_67462_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X633 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X634 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X635 a_66551_n13318# a_50751_n19729# a_66029_n14215# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X636 a_39179_n3548# a_31953_n19727# a_38619_n2651# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X637 a_42413_6405# a_41891_4481# a_41891_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X638 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X639 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X640 a_32353_n14213# a_31953_n19727# a_31831_n15110# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X641 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X642 a_79151_6405# a_77225_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X643 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X644 VDD a_30152_n35156# a_30682_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X645 a_54229_13546# a_53829_10388# a_53699_13546# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X646 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X647 a_53699_n35156# a_53829_n36382# a_55635_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X648 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X649 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X650 a_32353_n1754# a_31953_n19727# a_31831_n2651# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X651 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X652 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X653 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X654 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X655 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X656 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X657 a_34347_n2651# a_31953_n19727# a_33787_n1754# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X658 a_90935_4481# a_83153_11614# a_83325_4421# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X659 a_41487_n16904# a_31953_n19727# a_40965_n16904# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X660 a_35781_n7136# a_31953_n19727# a_35221_n6239# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X661 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X662 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X663 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X664 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X665 a_113037_n17715# a_71281_n8397# a_78344_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X666 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X667 a_98829_n14095# a_71281_n8397# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X668 a_93131_n7865# a_71281_n10073# a_92601_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X669 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X670 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X671 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X672 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X673 a_113037_n15000# a_71281_n8397# a_112199_n15000# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X674 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X675 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X676 a_54229_11614# a_53829_10388# a_53699_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X677 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X678 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X679 a_53699_n36322# a_53829_n36382# a_55635_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X680 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X681 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X682 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X683 a_83141_n18620# a_71281_n10073# a_82573_n18620# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X684 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X685 a_105365_n14095# a_71281_n8397# a_104527_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X686 a_66058_4481# a_65658_4421# a_65486_10448# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X687 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X688 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X689 a_83153_n35156# a_83325_n29313# a_85129_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X690 a_105933_n15905# a_71281_n8397# a_105365_n15905# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X691 a_72603_n10073# I1N a_71281_n10073# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X692 a_95105_n13190# a_71281_n10073# a_94537_n13190# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X693 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X694 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X695 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X696 a_89715_n16810# a_71281_n10073# a_89407_n13190# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X697 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X698 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X699 a_57417_n15112# a_50751_n19729# a_56895_n15112# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X700 a_53829_n36382# a_59558_n29181# a_61484_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X701 a_95943_n6960# a_71281_n10073# a_95105_n6960# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X702 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X703 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X704 a_44885_n16904# a_31953_n19727# a_44363_n17801# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X705 VDD a_31699_20742# a_31699_20742# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X706 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X707 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X708 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X709 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X710 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X711 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X712 a_81735_n18620# a_71281_n10073# a_81205_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X713 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X714 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X715 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X716 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X717 a_57417_n4447# a_50751_n19729# a_56895_n4447# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X718 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X719 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X720 a_93969_n8770# a_71281_n10073# a_93131_n8770# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X721 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X722 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X723 a_104527_n15905# a_71281_n8397# a_103997_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X724 a_112199_n4245# a_71281_n8397# a_111631_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X725 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X726 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X727 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X728 VDD a_30152_10448# a_30682_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X729 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X730 a_51151_n13318# a_50751_n19729# a_50629_n13318# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X731 a_71896_13546# a_71496_10388# a_71366_13546# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X732 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X733 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X734 a_94537_n3340# a_71281_n10073# a_93969_n3340# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X735 a_96849_12380# a_81205_n14095# a_84017_n17715# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X736 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X737 a_42413_n30339# a_41891_n29181# a_36162_n36382# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X738 a_88839_n13190# a_71281_n10073# a_88271_n13190# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X739 a_73302_10448# a_71496_10388# a_71342_7563# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X740 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X741 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X742 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X743 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X744 a_104527_n7865# a_71281_n8397# a_103997_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X745 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X746 a_82573_n9675# a_71281_n10073# a_81735_n9675# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X747 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X748 a_75585_n9297# I1N VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X749 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X750 a_113037_n20430# a_71281_n8397# a_112199_n20430# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X751 a_65486_n36322# a_65486_n35156# a_67422_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X752 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X753 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X754 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X755 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X756 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X757 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X758 a_99667_n9675# a_71281_n8397# a_98829_n9675# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X759 a_71896_11614# a_71496_10388# a_71366_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X760 a_102756_n34390# a_100820_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X761 a_34347_n13316# a_31953_n19727# a_33787_n12419# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X762 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X763 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X764 a_95414_n28415# a_94892_n29181# a_89163_n36382# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X765 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X766 a_94892_n29181# a_94892_n29181# a_96818_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X767 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X768 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X769 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X770 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X771 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X772 a_30152_10448# a_30324_4421# a_32128_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X773 a_35502_25545# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X774 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X775 VDD a_47819_11614# a_55601_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X776 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X777 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X778 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X779 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X780 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X781 a_46319_n17801# a_31953_n19727# a_45797_n18698# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X782 a_65486_n36322# a_65486_n35156# a_67422_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X783 a_40613_n8930# a_31953_n19727# a_40053_n8033# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X784 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X785 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X786 VDD a_65486_n35156# a_66016_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X787 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X788 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X789 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X790 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X791 a_57977_n8932# a_50751_n19729# a_57417_n8932# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X792 a_79182_13546# a_65658_4421# a_78344_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X793 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X794 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X795 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X796 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X797 a_43817_n29181# a_41891_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X798 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X799 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X800 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X801 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X802 VDD a_31699_20742# a_35502_24538# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X803 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X804 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X805 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X806 a_40053_n7136# a_31953_n19727# a_39531_n8033# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X807 a_49795_n29181# a_39179_n19595# a_38097_n16007# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X808 VDD a_65486_n35156# a_66016_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X809 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X810 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X811 a_31831_n5342# a_83325_n29313# a_83725_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X812 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X813 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X814 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X815 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X816 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X817 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X818 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X819 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X820 a_60080_n30339# a_59558_n29181# a_53829_n36382# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X821 a_54197_4481# a_47819_11614# a_53675_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X822 a_112199_n21335# a_71281_n8397# a_111631_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X823 a_102796_5639# a_100992_4421# a_56895_n16009# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X824 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X825 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X826 a_93969_n19525# a_71281_n10073# a_93131_n19525# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X827 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X828 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X829 a_79182_11614# a_65658_4421# a_78344_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X830 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X831 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X832 a_40613_n14213# a_31953_n19727# a_41487_n16007# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X833 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X834 a_41487_n7136# a_31953_n19727# a_40965_n8033# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X835 a_35781_n19595# a_31953_n19727# a_35221_n18698# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X836 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X837 a_32088_n35156# a_30152_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X838 a_35221_n6239# a_31953_n19727# a_34699_n6239# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X839 a_53675_n30339# a_53829_n36382# a_54229_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X840 a_55601_6405# a_47819_11614# a_47991_5507# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X841 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X842 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X843 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X844 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X845 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X846 a_87433_n3340# a_71281_n10073# a_86903_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X847 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X848 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X849 a_106501_n15000# a_71281_n8397# a_105933_n15000# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X850 a_89563_10448# a_89163_10388# a_71366_13546# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X851 a_67422_10448# a_65486_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X852 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X853 a_36162_10388# a_36032_11614# a_43848_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X854 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X855 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X856 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X857 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X858 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X859 a_43010_10448# a_30324_4421# a_42442_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X860 a_101641_n6960# a_71281_n8397# a_100803_n6960# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X861 a_32088_n33224# a_30152_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X862 VSS VSS VSS VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X863 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X864 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X865 a_113037_n18620# a_71281_n8397# a_112199_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X866 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X867 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X868 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X869 a_32913_n5342# a_31953_n19727# a_32353_n5342# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X870 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X871 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X872 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X873 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X874 a_52635_34067# a_35502_24538# a_33249_34067# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X875 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X876 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X877 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X878 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X879 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X880 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X881 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X882 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X883 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X884 a_71366_n35156# a_71496_n36382# a_73302_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X885 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X886 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X887 a_45138_23609# a_35922_19591# a_44608_22884# VDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X888 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X889 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X890 a_41891_4481# a_41891_4481# a_43817_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X891 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X892 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X893 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X894 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X895 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X896 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X897 a_78344_n36322# a_65658_n29313# a_77776_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X898 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X899 a_66058_n29181# a_65658_n29313# a_65486_n35156# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X900 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X901 a_81735_n17715# a_71281_n10073# a_81205_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X902 a_39179_n16007# a_31953_n19727# a_38619_n16007# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X903 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X904 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X905 a_71366_n36322# a_71496_n36382# a_73302_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X906 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X907 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X908 a_93969_n7865# a_71281_n10073# a_93131_n7865# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X909 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X910 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X911 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X912 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X913 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X914 VSS a_71496_n36382# a_71896_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X915 a_48313_n2651# a_31953_n19727# a_47753_n1754# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X916 a_106501_n20430# a_71281_n8397# a_105933_n20430# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X917 a_33787_n13316# a_31953_n19727# a_33265_n14213# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X918 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X919 a_66551_n12421# a_50751_n19729# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X920 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X921 a_60285_n16009# a_50751_n19729# a_59411_n14215# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X922 a_94537_n2435# a_71281_n10073# a_93969_n2435# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X923 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X924 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X925 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X926 a_45445_n6239# a_31953_n19727# a_44885_n4445# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X927 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X928 a_78344_n36322# a_65658_n29313# a_77776_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X929 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X930 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X931 a_59558_n29181# a_47991_n29313# a_61515_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X932 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X933 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X934 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X935 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X936 a_64243_n6241# a_50751_n19729# a_63683_n4447# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X937 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X938 a_51711_n19597# a_50751_n19729# a_51151_n19597# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X939 a_100820_10448# a_100992_4421# a_102796_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X940 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X941 a_31284_4481# a_30324_5507# a_30724_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X942 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X943 VSS VSS VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X944 a_71342_n27257# a_71496_n36382# a_71896_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X945 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X946 a_34347_n3548# a_31953_n19727# a_35221_n5342# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X947 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X948 a_89163_n36382# a_89033_n35156# a_96849_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X949 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X950 a_40613_n3548# a_31953_n19727# a_40053_n3548# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X951 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X952 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X953 a_83141_n21335# a_71281_n10073# a_82573_n21335# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X954 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X955 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X956 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X957 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X958 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X959 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X960 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X961 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X962 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X963 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X964 a_111063_n8770# a_71281_n8397# a_110225_n8770# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X965 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X966 a_85129_5639# a_83325_4421# a_50629_n16009# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X967 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X968 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X969 a_43817_7563# a_41891_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X970 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X971 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X972 a_60677_n36322# a_53699_n35156# a_60109_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X973 a_83709_n4245# a_71281_n10073# a_83141_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X974 a_32088_12380# a_30152_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X975 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X976 a_38097_n5342# a_39179_n8930# a_101392_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X977 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X978 a_111631_n3340# a_71281_n8397# a_111063_n3340# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X979 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X980 a_89163_n36382# a_89033_n35156# a_96849_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X981 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X982 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X983 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X984 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X985 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X986 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X987 a_81735_n21335# a_71281_n10073# a_81205_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X988 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X989 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X990 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X991 a_87433_n19525# a_71281_n10073# a_86903_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X992 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X993 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X994 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X995 a_101392_7563# a_57977_n12421# a_100820_11614# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X996 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X997 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X998 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X999 a_81735_n1530# a_71281_n10073# a_81205_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1000 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1001 a_45445_n19595# a_65486_n36322# a_71864_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1002 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1003 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1004 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1005 a_30724_7563# a_30324_5507# a_30152_11614# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1006 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1007 a_73268_n30339# a_65486_n36322# a_65658_n29313# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1008 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1009 a_98829_n1530# a_71281_n8397# a_98299_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1010 a_51151_n12421# a_50751_n19729# a_50629_n13318# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1011 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1012 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1013 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1014 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1015 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1016 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1017 a_65677_n17803# a_50751_n19729# a_65117_n17803# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1018 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1019 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1020 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1021 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1022 a_105933_n14095# a_71281_n8397# a_105365_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1023 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1024 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1025 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1026 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1027 a_30724_n28415# a_30324_n30399# a_30152_n36322# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1028 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1029 a_106501_n15905# a_71281_n8397# a_105933_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1030 a_61484_n29181# a_59558_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1031 a_108636_10448# a_106830_10388# a_106676_7563# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1032 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1033 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1034 a_87433_n2435# a_71281_n10073# a_53699_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1035 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1036 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1037 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1038 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1039 a_100820_n36322# a_39179_n8930# a_102796_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1040 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1041 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1042 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1043 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1044 a_60285_n8932# a_50751_n19729# a_57977_n8932# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1045 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1046 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1047 a_35221_n17801# a_31953_n19727# a_34699_n18698# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1048 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1049 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1050 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1051 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1052 a_104527_n14095# a_71281_n8397# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1053 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1054 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1055 a_95105_n4245# a_71281_n10073# a_94537_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1056 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1057 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1058 a_30324_n29313# a_30152_n36322# a_36530_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1059 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1060 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1061 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1062 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1063 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1064 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1065 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1066 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1067 a_89407_n13190# a_71281_n10073# a_88839_n13190# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1068 a_54019_n13318# a_50751_n19729# a_53497_n14215# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1069 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1070 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1071 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1072 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1073 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1074 a_103997_n8770# a_106830_n36382# a_108636_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1075 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1076 a_36008_7563# a_36162_10388# a_36562_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1077 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1078 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1079 a_100803_n13190# a_71281_n8397# a_100235_n13190# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1080 a_32913_n8930# a_83153_n36322# a_89531_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1081 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1082 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1083 a_40613_n19595# a_31953_n19727# a_40053_n19595# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1084 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1085 a_93131_n1530# a_71281_n10073# a_92601_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1086 a_43848_10448# a_36032_11614# a_43010_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1087 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1088 a_107198_n29181# a_100820_n36322# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1089 a_83325_4421# a_83153_11614# a_89531_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1090 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1091 a_73268_5639# a_65486_11614# a_64243_n1756# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1092 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1093 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1094 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1095 VSS a_71496_10388# a_71896_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1096 VSS VSS VSS VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1097 VDD a_31699_20742# a_35502_25545# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1098 a_52635_34067# a_35502_24538# a_33249_34067# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1099 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1100 a_102756_n36322# a_100820_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1101 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1102 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1103 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1104 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1105 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1106 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1107 VSS a_36162_10388# a_36562_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1108 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1109 a_48391_n28415# a_39179_n19595# a_47819_n36322# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1110 a_35221_n5342# a_31953_n19727# a_34347_n7136# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1111 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1112 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1113 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1114 a_32913_n16904# a_31953_n19727# a_32353_n16904# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1115 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1116 a_63683_n16009# a_50751_n19729# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1117 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1118 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1119 VDD a_83153_11614# a_90935_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1120 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1121 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1122 VDD a_31699_20742# a_35502_24538# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1123 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1124 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1125 a_95943_n20430# a_71281_n10073# a_95105_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1126 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1127 a_84547_n6055# a_71281_n10073# a_43010_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1128 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1129 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1130 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1131 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1132 a_51151_n8035# a_50751_n19729# a_50629_n8932# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1133 a_30152_n36322# a_30324_n30399# a_32128_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1134 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1135 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1136 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1137 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1138 VSS a_112559_4481# a_113081_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1139 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1140 a_45706_24920# a_35922_19591# a_45138_24920# VDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X1141 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1142 a_83153_11614# a_83153_10448# a_85089_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1143 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1144 a_53145_n8932# a_50751_n19729# a_52585_n8035# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1145 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1146 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1147 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1148 VSS a_112559_n29181# a_113081_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1149 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1150 a_101350_n35156# a_100820_n35156# a_100820_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1151 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1152 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1153 a_111063_n7865# a_71281_n8397# a_110225_n7865# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1154 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1155 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1156 a_71496_10388# a_77225_4481# a_79151_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1157 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1158 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1159 a_41487_n12419# a_31953_n19727# a_39179_n12419# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1160 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1161 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1162 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1163 a_94537_n19525# a_71281_n10073# a_93969_n19525# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1164 a_89531_7563# a_83153_11614# a_89009_7563# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1165 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1166 a_104527_n1530# a_71281_n8397# a_103997_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1167 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1168 a_111631_n2435# a_71281_n8397# a_111063_n2435# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1169 a_82573_n3340# a_71281_n10073# a_81735_n3340# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1170 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1171 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1172 VSS a_35502_25545# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1173 a_71496_10388# a_71366_11614# a_79182_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1174 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1175 a_30152_n36322# a_30152_n35156# a_32088_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1176 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1177 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1178 a_67462_n30339# a_65658_n29313# a_44363_n16007# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1179 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1180 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1181 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1182 a_47753_n4445# a_31953_n19727# a_47231_n6239# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1183 a_99667_n3340# a_71281_n8397# a_98829_n3340# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1184 a_101350_n33224# a_100820_n35156# a_100820_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1185 a_48313_n19595# a_31953_n19727# a_47753_n18698# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1186 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1187 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1188 VDD a_31699_20742# a_35502_25545# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1189 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1190 VSS VSS VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1191 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1192 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1193 a_35502_25545# a_35502_25545# VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X1194 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1195 a_58851_n19597# a_50751_n19729# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1196 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1197 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1198 a_113037_n15000# a_71281_n8397# a_112199_n14095# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1199 a_90245_n8770# a_71281_n10073# a_89407_n8770# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1200 a_63161_n5344# a_65658_4421# a_66058_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1201 a_60845_n15112# a_50751_n19729# a_60285_n14215# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1202 a_63683_n7138# a_50751_n19729# a_63161_n7138# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1203 a_30152_n36322# a_30152_n35156# a_32088_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1204 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1205 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1206 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1207 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1208 a_36008_7563# a_30152_11614# a_37934_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1209 a_65677_n7138# a_50751_n19729# a_65117_n7138# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1210 a_44885_n12419# a_31953_n19727# a_44363_n13316# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1211 a_77747_4481# a_77225_4481# a_77225_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1212 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1213 a_60285_n15112# a_50751_n19729# a_59763_n16906# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1214 a_36162_n36382# a_41891_n29181# a_43817_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1215 a_100803_n4245# a_71281_n8397# a_100235_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1216 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1217 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1218 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1219 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1220 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1221 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1222 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1223 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1224 a_95943_n6055# a_71281_n10073# a_78344_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1225 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1226 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1227 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1228 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1229 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1230 a_84547_n18620# a_71281_n10073# a_83709_n18620# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1231 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1232 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1233 a_40613_n2651# a_31953_n19727# a_40053_n2651# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1234 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1235 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1236 a_54579_n15112# a_50751_n19729# a_54019_n14215# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1237 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1238 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1239 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1240 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1241 a_64243_n14215# a_50751_n19729# a_63683_n14215# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1242 a_79151_n30339# a_77225_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1243 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1244 VSS a_35502_25545# a_33249_34067# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1245 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1246 a_32128_4481# a_30324_5507# a_31284_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1247 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1248 a_32353_n8930# a_31953_n19727# a_31831_n8930# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1249 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1250 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1251 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1252 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1253 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1254 a_34347_n8930# a_31953_n19727# a_33787_n8930# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1255 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1256 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1257 a_45706_24195# a_35922_19591# a_45138_24195# VDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X1258 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1259 a_77747_n28415# a_77225_n29181# a_71496_n36382# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1260 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1261 a_40053_n1754# a_31953_n19727# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1262 a_35502_24538# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1263 a_83725_n30339# a_32913_n8930# a_83153_n36322# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1264 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1265 a_54229_10448# a_53829_10388# a_36032_13546# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1266 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1267 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1268 VDD a_31699_20742# a_31699_20742# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1269 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1270 a_33249_34067# a_35502_24538# a_52635_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1271 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1272 a_46319_n13316# a_31953_n19727# a_45797_n14213# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1273 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1274 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1275 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1276 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1277 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1278 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1279 a_57977_n14215# a_50751_n19729# a_57417_n14215# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1280 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1281 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1282 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1283 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X1284 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1285 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1286 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1287 a_41487_n1754# a_31953_n19727# a_39179_n1754# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1288 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1289 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1290 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1291 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1292 a_89715_n17715# a_100992_4421# a_113110_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1293 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1294 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1295 a_57977_n6241# a_50751_n19729# a_57417_n4447# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1296 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1297 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1298 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1299 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1300 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1301 a_51151_n3550# a_50751_n19729# a_50629_n4447# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1302 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1303 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1304 a_35502_25545# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1305 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1306 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1307 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1308 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1309 a_53145_n3550# a_50751_n19729# a_52585_n3550# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1310 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1311 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1312 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1313 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1314 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1315 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1316 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1317 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1318 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1319 a_110225_n9675# a_71281_n8397# a_109695_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1320 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1321 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1322 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1323 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1324 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1325 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1326 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1327 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1328 a_37968_13546# a_36162_10388# a_36008_4481# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1329 a_47991_4421# a_47819_11614# a_54197_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1330 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1331 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1332 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1333 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1334 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1335 a_85129_n29181# a_32913_n8930# a_31831_n5342# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1336 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1337 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1338 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1339 a_93969_n1530# a_71281_n10073# a_93131_n1530# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1340 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1341 a_99667_n13190# a_71281_n8397# a_98829_n13190# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1342 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1343 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1344 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1345 VSS a_89163_10388# a_89563_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1346 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1347 a_114485_5639# a_112559_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1348 a_47753_n19595# a_31953_n19727# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1349 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1350 a_111063_n13190# a_71281_n8397# a_110225_n13190# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1351 a_71896_10448# a_71496_10388# a_53699_13546# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1352 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1353 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1354 a_113037_n6055# a_71281_n8397# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1355 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1356 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1357 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1358 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1359 a_37968_11614# a_36162_10388# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1360 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1361 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1362 a_82573_n2435# a_71281_n10073# a_81735_n2435# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1363 VSS VSS VSS VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1364 a_54019_n12421# a_50751_n19729# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1365 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1366 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1367 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1368 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1369 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1370 a_89531_n29181# a_83153_n36322# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1371 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1372 a_106501_n14095# a_71281_n8397# a_105933_n14095# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1373 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1374 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1375 a_99667_n2435# a_71281_n8397# a_98829_n2435# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1376 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1377 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1378 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1379 a_65117_n7138# a_50751_n19729# a_64595_n8035# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1380 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1381 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1382 a_101641_n6055# a_71281_n8397# a_101111_n6055# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1383 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1384 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1385 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1386 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1387 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1388 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1389 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1390 a_38097_n16007# a_47991_n29313# a_48391_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1391 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1392 a_90245_n8770# a_71281_n10073# a_89407_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1393 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1394 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1395 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1396 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1397 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1398 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1399 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1400 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1401 a_112559_n29181# a_112559_n29181# a_114485_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1402 a_33379_34007# IN_POS cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
X1403 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1404 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1405 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1406 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1407 a_67111_n8932# a_50751_n19729# a_66551_n8035# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1408 a_67462_5639# a_65658_4421# a_63161_n5344# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1409 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1410 a_63683_n15112# a_50751_n19729# a_63161_n15112# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1411 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1412 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1413 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1414 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1415 a_33249_34067# a_35502_24538# a_52635_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1416 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1417 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1418 a_88839_n4245# a_71281_n10073# a_88271_n4245# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1419 VDD a_30152_n36322# a_37934_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1420 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1421 a_79182_10448# a_71366_11614# a_78344_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1422 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1423 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1424 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1425 a_45445_n18698# a_31953_n19727# a_44885_n18698# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1426 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1427 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1428 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1429 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1430 a_35781_n15110# a_31953_n19727# a_35221_n15110# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1431 a_94892_4481# a_94892_4481# a_96818_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1432 a_84547_n17715# a_71281_n10073# a_84017_n17715# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1433 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X1434 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1435 VSS a_53829_n36382# a_54229_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1436 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1437 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1438 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1439 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1440 OUT a_35502_24538# a_33249_35053# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1441 a_66551_n18700# a_50751_n19729# a_66029_n18700# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1442 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1443 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1444 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1445 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1446 a_46879_n14213# a_31953_n19727# a_46319_n14213# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1447 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1448 a_89033_n36322# a_106830_n36382# a_108636_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1449 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1450 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1451 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1452 a_32353_n19595# a_31953_n19727# a_31831_n19595# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1453 VDD a_31699_20742# a_31699_20742# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1454 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1455 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1456 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1457 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1458 a_95414_n27257# a_94892_n29181# a_94892_n29181# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1459 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X1460 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1461 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1462 a_38619_n4445# a_31953_n19727# a_38097_n4445# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1463 a_53675_n27257# a_53829_n36382# a_54229_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1464 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1465 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1466 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1467 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1468 VDD a_100820_10448# a_101350_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1469 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1470 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1471 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1472 a_112559_4481# a_112559_4481# a_114485_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1473 a_50629_n16009# a_51711_n12421# a_83725_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1474 VSS a_41891_4481# a_42413_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1475 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1476 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1477 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1478 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1479 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1480 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1481 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1482 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1483 a_31699_20742# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1484 a_71281_n8397# I1N a_75585_n10973# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X1485 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1486 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1487 a_63683_n6241# a_50751_n19729# a_63161_n7138# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1488 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1489 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1490 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1491 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1492 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1493 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1494 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1495 a_96818_5639# a_94892_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1496 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1497 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1498 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1499 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1500 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1501 a_53675_n27257# a_47819_n36322# a_55601_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1502 a_113110_13546# a_86903_n14095# a_106830_10388# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1503 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1504 a_83141_n4245# a_71281_n10073# a_82573_n4245# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1505 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1506 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1507 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1508 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1509 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1510 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1511 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1512 a_48349_13546# a_47819_10448# a_47819_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1513 VDD a_71281_n10073# a_83709_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1514 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1515 a_100235_n4245# a_71281_n8397# a_99667_n4245# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1516 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1517 a_56895_n16009# a_57977_n12421# a_101392_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1518 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1519 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1520 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1521 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1522 a_39179_n19595# a_47819_n36322# a_54197_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1523 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1524 a_59411_n7138# a_50751_n19729# a_60285_n5344# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1525 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1526 a_107339_n6960# a_71281_n8397# a_106501_n6960# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1527 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1528 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1529 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1530 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1531 a_65677_n13318# a_50751_n19729# a_65117_n13318# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1532 a_113110_11614# a_86903_n14095# a_106830_10388# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1533 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1534 a_101641_n20430# a_71281_n8397# a_100803_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1535 a_48313_n8930# a_31953_n19727# a_47753_n8930# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1536 a_113081_7563# a_112559_4481# a_106830_10388# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1537 a_51151_n18700# a_50751_n19729# a_50629_n19597# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1538 a_51711_n8035# a_50751_n19729# a_51151_n7138# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1539 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1540 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1541 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1542 a_65486_10448# a_65658_4421# a_67462_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1543 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1544 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1545 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1546 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1547 a_53829_n36382# a_53699_n35156# a_61515_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1548 a_86903_n14095# a_106830_10388# a_108636_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1549 a_48349_11614# a_47819_10448# a_47819_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1550 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1551 a_67422_n34390# a_65486_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1552 a_83725_5639# a_51711_n12421# a_83153_11614# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1553 a_42413_7563# a_41891_4481# a_36162_10388# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1554 a_51711_n16009# a_50751_n19729# a_51151_n16009# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1555 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1556 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1557 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1558 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1559 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1560 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1561 a_79151_7563# a_77225_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1562 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1563 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1564 a_60285_n4447# a_50751_n19729# a_59763_n6241# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1565 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1566 a_113037_n6960# a_71281_n8397# a_112199_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1567 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1568 a_35221_n13316# a_31953_n19727# a_34699_n14213# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1569 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1570 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1571 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1572 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1573 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1574 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1575 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1576 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1577 a_53829_n36382# a_53699_n35156# a_61515_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1578 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1579 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1580 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1581 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1582 a_60677_n36322# a_47991_n29313# a_60109_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1583 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1584 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1585 a_107339_n20430# a_71281_n8397# a_106501_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1586 a_110225_n13190# a_71281_n8397# a_109695_n16810# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1587 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1588 a_67111_n4447# a_50751_n19729# a_66551_n3550# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1589 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1590 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1591 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1592 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1593 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1594 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1595 a_111063_n1530# a_71281_n8397# a_110225_n1530# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1596 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1597 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1598 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1599 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1600 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1601 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1602 OUT a_35502_24538# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1603 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1604 a_82573_n15000# a_71281_n10073# a_81735_n15000# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1605 a_60677_n36322# a_47991_n29313# a_60109_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1606 a_51151_n2653# a_50751_n19729# a_50629_n2653# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1607 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1608 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1609 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1610 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1611 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1612 a_33249_35053# a_35502_24538# OUT VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1613 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1614 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1615 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1616 a_53145_n2653# a_50751_n19729# a_52585_n2653# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1617 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1618 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1619 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1620 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1621 VSS VSS VSS VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1622 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1623 VSS a_59558_n29181# a_60080_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1624 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1625 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1626 VDD a_65486_11614# a_73268_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1627 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1628 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1629 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1630 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1631 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1632 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1633 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1634 a_32913_n12419# a_31953_n19727# a_32353_n12419# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1635 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1636 a_46274_23609# a_35922_19591# a_45706_23609# VDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X1637 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1638 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1639 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1640 VSS a_35502_25545# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1641 VSS a_35502_24538# a_41100_19075# VSS nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X1642 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1643 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1644 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1645 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1646 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1647 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1648 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1649 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1650 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1651 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1652 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1653 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1654 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1655 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1656 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1657 a_67111_n17803# a_50751_n19729# a_66551_n17803# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1658 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1659 a_105365_n9675# a_71281_n8397# a_104527_n9675# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1660 a_63683_n1756# a_50751_n19729# a_63161_n2653# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1661 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1662 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1663 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1664 a_105933_n4245# a_71281_n8397# a_105365_n4245# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1665 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1666 a_82573_n20430# a_71281_n10073# a_81735_n20430# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1667 a_53675_4481# a_47819_11614# a_55601_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1668 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1669 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1670 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1671 a_65677_n2653# a_50751_n19729# a_65117_n1756# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1672 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1673 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1674 a_71864_5639# a_65486_11614# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1675 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1676 a_43817_n30339# a_41891_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1677 a_42442_13546# a_36032_11614# a_36162_10388# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1678 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1679 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1680 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1681 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1682 a_53829_10388# a_53699_11614# a_61515_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1683 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1684 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1685 a_38619_n17801# a_31953_n19727# a_38097_n17801# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1686 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1687 a_100235_n18620# a_71281_n8397# a_99667_n18620# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1688 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1689 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1690 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1691 a_49795_n30339# a_47991_n29313# a_38097_n16007# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1692 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1693 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1694 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1695 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1696 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1697 a_52635_34067# a_35502_24538# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1698 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1699 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1700 a_96818_n28415# a_94892_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1701 a_111631_n13190# a_71281_n8397# a_111063_n13190# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1702 a_65658_n29313# a_65486_n36322# a_71864_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1703 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1704 a_42442_11614# a_36032_11614# a_36162_10388# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1705 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1706 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1707 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1708 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1709 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1710 a_36032_11614# a_36162_10388# a_37968_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1711 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1712 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1713 a_102756_n35156# a_100820_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1714 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1715 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1716 a_36162_10388# a_41891_4481# a_43817_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1717 a_35781_n15110# a_31953_n19727# a_35221_n14213# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1718 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1719 a_36008_4481# a_36162_10388# a_36562_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1720 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1721 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1722 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1723 a_98829_n18620# a_71281_n8397# a_98299_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1724 a_30152_11614# a_30324_5507# a_32128_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1725 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1726 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1727 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1728 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1729 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1730 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1731 a_33787_n18698# a_31953_n19727# a_33265_n18698# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1732 a_30724_n27257# a_30324_n29313# a_30152_n35156# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1733 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1734 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1735 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1736 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1737 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1738 a_105365_n18620# a_71281_n8397# a_104527_n18620# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1739 a_55601_7563# a_47819_11614# a_47991_4421# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1740 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1741 a_102756_n33224# a_100820_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1742 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1743 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1744 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1745 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1746 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1747 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1748 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1749 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1750 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1751 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1752 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1753 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1754 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1755 VDD a_31699_20742# a_31699_20742# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1756 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1757 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1758 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1759 a_110225_n3340# a_71281_n8397# a_109695_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1760 a_100820_11614# a_57977_n12421# a_102796_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1761 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1762 a_31284_4481# a_30324_4421# a_30724_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1763 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1764 a_58851_n8035# a_50751_n19729# a_58329_n8035# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1765 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1766 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1767 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1768 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1769 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1770 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1771 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1772 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1773 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1774 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1775 a_57417_n16906# a_50751_n19729# a_56895_n17803# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1776 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1777 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1778 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1779 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1780 a_102796_6405# a_57977_n12421# a_56895_n16009# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1781 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1782 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1783 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1784 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1785 a_82573_n15905# a_71281_n10073# a_81735_n15905# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1786 a_43817_4481# a_41891_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1787 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1788 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1789 a_66058_n30339# a_45445_n19595# a_65486_n36322# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1790 a_48313_n15110# a_31953_n19727# a_47753_n15110# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1791 a_112199_n6960# a_71281_n8397# a_111631_n6960# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1792 a_83325_n29313# a_83153_n36322# a_89531_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1793 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1794 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1795 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1796 a_89563_n34390# a_89163_n36382# a_89033_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1797 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1798 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1799 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1800 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1801 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1802 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1803 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1804 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1805 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1806 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1807 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1808 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1809 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1810 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1811 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1812 a_41100_19075# a_35502_24538# a_40578_19075# VSS nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X1813 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1814 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1815 a_35502_24538# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1816 a_48391_n27257# a_47991_n29313# a_47819_n35156# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1817 a_101392_4481# a_100992_4421# a_100820_10448# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1818 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1819 a_65677_n13318# a_50751_n19729# a_65117_n12421# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1820 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1821 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1822 a_51711_n6241# a_50751_n19729# a_51151_n6241# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1823 a_89715_n5150# a_71281_n10073# a_89407_n1530# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1824 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1825 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1826 a_65486_n36322# a_45445_n19595# a_67462_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1827 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1828 a_30724_4481# a_30324_4421# a_30152_10448# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1829 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1830 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1831 a_51711_n16906# a_50751_n19729# a_51151_n15112# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1832 a_107198_5639# a_100820_11614# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1833 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1834 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1835 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1836 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1837 a_65117_n1756# a_50751_n19729# a_64243_n5344# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1838 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1839 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1840 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1841 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1842 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1843 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1844 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1845 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1846 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1847 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1848 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1849 a_90969_13546# a_89163_10388# a_89009_4481# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1850 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1851 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1852 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1853 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1854 VSS a_106830_n36382# a_107230_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1855 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1856 a_89407_n8770# a_71281_n10073# a_88839_n8770# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1857 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1858 a_67111_n2653# a_50751_n19729# a_66551_n2653# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1859 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1860 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1861 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1862 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1863 a_32353_n8033# a_31953_n19727# a_31831_n8930# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1864 a_53145_n7138# a_50751_n19729# a_54019_n5344# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1865 a_40053_n8930# a_31953_n19727# a_39179_n5342# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1866 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1867 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1868 a_54019_n18700# a_50751_n19729# a_53497_n18700# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1869 a_40053_n12419# a_31953_n19727# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1870 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1871 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1872 a_90969_11614# a_89163_10388# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1873 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1874 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X1875 a_34347_n8930# a_31953_n19727# a_33787_n8033# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1876 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1877 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1878 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1879 VDD a_47819_10448# a_48349_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1880 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1881 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1882 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1883 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1884 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1885 a_67422_n36322# a_65486_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1886 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1887 a_41487_n8930# a_31953_n19727# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1888 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1889 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1890 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1891 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1892 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1893 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1894 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1895 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1896 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1897 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1898 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1899 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1900 a_61484_n30339# a_59558_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1901 a_83325_4421# a_83153_11614# a_89531_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1902 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1903 a_98829_n17715# a_71281_n8397# a_98299_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1904 VSS VSS VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1905 a_100820_n35156# a_100992_n29313# a_102796_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1906 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1907 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1908 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1909 a_85129_6405# a_51711_n12421# a_50629_n16009# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1910 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1911 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1912 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1913 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1914 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1915 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1916 VDD a_31699_20742# a_35502_25545# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1917 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1918 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1919 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1920 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1921 a_58851_n3550# a_50751_n19729# a_58329_n3550# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1922 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1923 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1924 a_95443_n34390# a_89033_n35156# a_89163_n36382# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1925 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1926 a_95443_12380# a_83325_4421# a_94892_4481# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1927 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1928 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1929 a_44885_n7136# a_31953_n19727# a_44363_n7136# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1930 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1931 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1932 a_34347_n17801# a_31953_n19727# a_33787_n17801# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1933 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1934 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1935 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1936 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1937 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1938 a_90245_n17715# a_71281_n10073# a_89715_n16810# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1939 a_46879_n7136# a_31953_n19727# a_46319_n7136# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1940 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1941 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1942 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1943 VDD a_65486_n36322# a_73268_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1944 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1945 a_95105_n15000# a_71281_n10073# a_94537_n15000# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1946 a_47753_n16007# a_31953_n19727# a_46879_n17801# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1947 a_110225_n2435# a_71281_n8397# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1948 a_88271_n4245# a_71281_n10073# a_87433_n4245# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1949 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1950 a_90245_n15000# a_71281_n10073# a_89407_n15000# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1951 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1952 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1953 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1954 a_37968_10448# a_36162_10388# a_36008_7563# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1955 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1956 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1957 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1958 a_77747_n27257# a_77225_n29181# a_77225_n29181# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1959 a_100235_n21335# a_71281_n8397# a_99667_n21335# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1960 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1961 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1962 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1963 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1964 a_42047_n7136# a_31953_n19727# a_41487_n6239# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1965 VDD a_65486_10448# a_66016_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1966 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1967 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1968 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1969 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1970 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1971 a_112559_n29181# a_100992_n29313# a_114516_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1972 a_60677_10448# a_53699_11614# a_60109_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1973 a_32128_n28415# a_30324_n29313# a_31284_n30339# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1974 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1975 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1976 a_107198_n30339# a_100820_n36322# a_106676_n30339# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1977 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1978 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1979 a_89531_4481# a_83153_11614# a_89009_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1980 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1981 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1982 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1983 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1984 a_88839_n15000# a_71281_n10073# a_88271_n15000# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1985 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1986 a_30324_5507# a_50751_n19729# a_51151_n1756# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1987 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1988 a_98829_n21335# a_71281_n8397# a_98299_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1989 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1990 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1991 VSS a_94892_4481# a_95414_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1992 a_60677_10448# a_53699_11614# a_60109_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1993 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1994 a_60845_n19597# a_50751_n19729# a_60285_n19597# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1995 a_101350_12380# a_100820_10448# a_100820_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1996 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1997 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1998 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1999 a_36530_n28415# a_30152_n36322# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2000 a_106809_n5150# a_103997_n8770# a_113110_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2001 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2002 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2003 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2004 a_105365_n21335# a_71281_n8397# a_104527_n21335# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2005 VDD a_100820_n36322# a_108602_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2006 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2007 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2008 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2009 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2010 a_45445_n16904# a_31953_n19727# a_44885_n15110# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2011 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2012 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2013 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2014 a_95105_n20430# a_71281_n10073# a_94537_n20430# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2015 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2016 OUT a_35502_24538# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2017 a_89009_4481# a_83153_11614# a_90935_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2018 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2019 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2020 a_90245_n20430# a_71281_n10073# a_89407_n20430# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2021 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2022 a_83709_n6960# a_71281_n10073# a_83141_n6960# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2023 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2024 a_39179_n6239# a_31953_n19727# a_38619_n4445# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2025 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2026 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2027 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2028 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2029 a_103997_n8770# a_106830_n36382# a_108636_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2030 a_54579_n19597# a_50751_n19729# a_54019_n19597# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2031 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2032 a_32353_n16007# a_31953_n19727# a_31284_n30339# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2033 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2034 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2035 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2036 VSS a_112559_4481# a_113081_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2037 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2038 a_54019_n5344# a_50751_n19729# a_53145_n3550# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2039 a_64243_n19597# a_50751_n19729# a_63683_n19597# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2040 a_49755_n34390# a_47819_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2041 a_107339_n6055# a_71281_n8397# a_106809_n6055# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2042 a_32353_n3548# a_31953_n19727# a_31831_n4445# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2043 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2044 a_73268_6405# a_65486_11614# a_64243_n1756# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2045 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2046 a_34347_n3548# a_31953_n19727# a_33787_n3548# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2047 a_77225_4481# a_77225_4481# a_79151_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2048 I1U I1U VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X2049 a_88839_n20430# a_71281_n10073# a_88271_n20430# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2050 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2051 a_89407_n7865# a_71281_n10073# a_88839_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2052 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2053 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2054 a_95414_5639# a_94892_4481# a_89163_10388# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2055 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2056 VCM a_106830_n36382# a_108636_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2057 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2058 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2059 a_48313_n15110# a_31953_n19727# a_47753_n14213# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2060 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2061 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2062 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2063 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2064 a_46319_n18698# a_31953_n19727# a_45797_n18698# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2065 a_105933_n18620# a_71281_n8397# a_105365_n18620# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2066 a_105365_n3340# a_71281_n8397# a_104527_n3340# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2067 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X2068 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2069 a_35922_19591# a_35502_25545# VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X2070 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2071 a_57977_n19597# a_50751_n19729# a_57417_n19597# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2072 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2073 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2074 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2075 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2076 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2077 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2078 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2079 a_106830_n36382# a_112559_n29181# a_114485_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2080 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2081 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2082 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2083 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2084 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2085 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2086 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2087 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2088 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2089 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2090 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2091 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2092 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2093 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2094 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2095 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2096 a_36008_n30339# a_30152_n36322# a_37934_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2097 a_106501_n8770# a_71281_n8397# a_105933_n8770# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2098 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2099 a_104527_n18620# a_71281_n8397# a_103997_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2100 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2101 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2102 a_46319_n7136# a_31953_n19727# a_45797_n8033# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2103 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2104 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X2105 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2106 a_82573_n14095# a_71281_n10073# a_81735_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2107 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2108 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2109 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2110 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2111 a_114516_12380# a_86903_n14095# a_89715_n17715# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2112 a_95105_n6960# a_71281_n10073# a_94537_n6960# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2113 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2114 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2115 a_113110_10448# a_100992_4421# a_112559_4481# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2116 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2117 VSS a_41891_n29181# a_42413_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2118 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2119 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2120 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2121 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2122 a_66551_n5344# a_50751_n19729# a_65677_n3550# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2123 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2124 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2125 a_35502_24538# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2126 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2127 a_48349_10448# a_47819_10448# a_47819_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2128 a_95105_n15905# a_71281_n10073# a_94537_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2129 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2130 a_90245_n18620# a_71281_n10073# a_89407_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2131 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2132 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2133 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2134 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2135 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2136 a_48313_n8930# a_31953_n19727# a_47753_n8033# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2137 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2138 a_89563_n36322# a_89163_n36382# a_89033_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2139 OUT a_35502_24538# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2140 a_59411_n7138# a_50751_n19729# a_58851_n7138# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2141 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2142 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2143 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2144 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2145 VSS a_106830_10388# a_107230_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2146 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2147 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2148 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2149 a_30682_n34390# a_30152_n35156# a_30152_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2150 a_67111_n13318# a_50751_n19729# a_66551_n13318# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2151 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2152 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2153 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2154 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2155 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2156 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2157 a_81735_n9675# a_71281_n10073# a_81205_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2158 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X2159 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2160 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2161 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2162 a_72603_n10973# I1N I1N VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X2163 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2164 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2165 a_98829_n9675# a_71281_n8397# a_98299_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2166 a_88839_n15905# a_71281_n10073# a_88271_n15905# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2167 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2168 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2169 a_30682_12380# a_30152_10448# a_30152_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2170 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2171 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2172 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2173 a_42047_n17801# a_31953_n19727# a_41487_n16904# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2174 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2175 a_77225_n29181# a_77225_n29181# a_79151_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2176 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2177 VDD a_83153_n36322# a_90935_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2178 a_55635_n34390# a_53829_n36382# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2179 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2180 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2181 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2182 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2183 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2184 a_38619_n13316# a_31953_n19727# a_38097_n13316# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2185 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2186 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2187 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2188 a_64243_n1756# a_65486_11614# a_71864_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2189 a_52585_n17803# a_50751_n19729# a_52063_n18700# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2190 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2191 VCM a_33379_34007# cap_mim_2f0_m4m5_noshield c_width=9.8u c_length=9.8u
X2192 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2193 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2194 a_84547_n8770# a_71281_n10073# a_83709_n8770# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2195 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2196 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2197 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2198 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2199 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2200 a_60109_n34390# a_53699_n35156# a_53829_n36382# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2201 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2202 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2203 a_47991_n29313# a_47819_n36322# a_54197_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2204 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2205 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2206 a_85129_n30339# a_83325_n29313# a_31831_n5342# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2207 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2208 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2209 a_78344_10448# a_71366_11614# a_77776_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2210 a_36032_13546# a_53829_10388# a_55635_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2211 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2212 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2213 a_58851_n2653# a_50751_n19729# a_58329_n3550# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2214 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2215 a_106676_n30339# a_106830_n36382# a_107230_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2216 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2217 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2218 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2219 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2220 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2221 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2222 a_81205_n14095# a_89163_10388# a_90969_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2223 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2224 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2225 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2226 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2227 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2228 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2229 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2230 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2231 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2232 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2233 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2234 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2235 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2236 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2237 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2238 a_46879_n19595# a_31953_n19727# a_46319_n19595# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2239 a_78344_10448# a_71366_11614# a_77776_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2240 a_53699_11614# a_53829_10388# a_55635_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2241 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2242 a_35922_19591# a_35922_19591# a_46274_24920# VDD pfet_03v3 ad=0.78p pd=3.7u as=0.78p ps=3.7u w=1.2u l=2u
X2243 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2244 a_89531_n30339# a_83153_n36322# a_89009_n30339# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2245 a_113037_n18620# a_71281_n8397# a_112199_n18620# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2246 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2247 a_40613_n3548# a_31953_n19727# a_41487_n5342# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2248 a_93131_n9675# a_71281_n10073# a_92601_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2249 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2250 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2251 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2252 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2253 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2254 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2255 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2256 a_39179_n16904# a_31953_n19727# a_38619_n16904# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2257 a_38097_n16007# a_39179_n19595# a_48391_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2258 a_32913_n8033# a_31953_n19727# a_32353_n7136# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2259 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2260 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2261 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2262 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2263 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2264 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2265 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2266 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2267 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2268 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2269 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2270 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2271 a_100803_n6960# a_71281_n8397# a_100235_n6960# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2272 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2273 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2274 a_105365_n2435# a_71281_n8397# a_104527_n2435# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2275 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2276 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2277 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2278 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2279 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2280 a_60285_n16906# a_50751_n19729# a_59763_n16906# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2281 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2282 a_106830_10388# a_112559_4481# a_114485_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2283 VSS a_41891_4481# a_42413_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2284 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2285 a_95443_n36322# a_89033_n35156# a_89163_n36382# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2286 a_95943_n8770# a_71281_n10073# a_95105_n8770# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2287 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2288 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2289 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2290 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2291 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2292 a_53699_13546# a_71496_10388# a_73302_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2293 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2294 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2295 a_42442_10448# a_30324_4421# a_41891_4481# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2296 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2297 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2298 a_114485_6405# a_112559_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2299 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2300 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2301 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2302 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2303 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2304 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2305 a_106501_n7865# a_71281_n8397# a_105933_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2306 a_45445_n14213# a_31953_n19727# a_44885_n14213# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2307 a_104527_n17715# a_71281_n8397# a_103997_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2308 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2309 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2310 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2311 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2312 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2313 a_48313_n4445# a_31953_n19727# a_47753_n3548# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2314 a_112199_n19525# a_71281_n8397# a_111631_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2315 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2316 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2317 a_66551_n14215# a_50751_n19729# a_66029_n14215# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2318 a_71366_11614# a_71496_10388# a_73302_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2319 a_61515_n34390# a_47991_n29313# a_60677_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2320 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2321 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2322 a_52635_34067# a_35502_24538# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2323 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2324 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2325 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2326 a_104527_n9675# a_71281_n8397# a_103997_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2327 a_65677_n19597# a_50751_n19729# a_65117_n18700# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2328 a_112559_n29181# a_100992_n29313# a_114516_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2329 a_56895_n16009# a_100992_4421# a_101392_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2330 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2331 a_45445_n6239# a_31953_n19727# a_44885_n6239# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2332 a_47819_n36322# a_39179_n19595# a_49795_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2333 a_89407_n15000# a_71281_n10073# a_88839_n15000# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2334 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2335 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2336 a_32353_n2651# a_31953_n19727# a_31831_n2651# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2337 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2338 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2339 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2340 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2341 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2342 a_113081_4481# a_112559_4481# a_112559_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2343 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2344 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2345 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X2346 a_100803_n15000# a_71281_n8397# a_100235_n15000# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2347 a_34347_n2651# a_31953_n19727# a_33787_n2651# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2348 a_65486_11614# a_64243_n1756# a_67462_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2349 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2350 a_41487_n17801# a_31953_n19727# a_40965_n18698# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2351 a_35781_n7136# a_31953_n19727# a_35221_n7136# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2352 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2353 a_57977_n12421# a_100820_11614# a_107198_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2354 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2355 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2356 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2357 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2358 a_42413_4481# a_41891_4481# a_41891_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2359 a_35221_n18698# a_31953_n19727# a_34699_n18698# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2360 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2361 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2362 a_105933_n21335# a_71281_n8397# a_105365_n21335# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2363 a_79151_4481# a_77225_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2364 a_107230_13546# a_106830_10388# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2365 a_106809_n5150# a_103997_n8770# a_113110_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2366 a_67462_6405# a_64243_n1756# a_63161_n5344# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2367 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2368 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X2369 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2370 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2371 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2372 a_35502_25545# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2373 a_101392_n29181# a_100992_n29313# a_100820_n35156# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2374 a_72603_n8397# I1N a_71281_n8397# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X2375 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2376 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2377 a_89163_10388# a_94892_4481# a_96818_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2378 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2379 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2380 a_107230_11614# a_106830_10388# a_86903_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2381 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2382 a_84547_n8770# a_71281_n10073# a_83709_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2383 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2384 a_96818_n27257# a_94892_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2385 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2386 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2387 a_104527_n21335# a_71281_n8397# a_103997_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2388 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2389 a_44885_n17801# a_31953_n19727# a_44363_n17801# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2390 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2391 a_44885_n1754# a_31953_n19727# a_44363_n2651# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2392 a_49755_n36322# a_47819_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2393 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2394 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2395 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2396 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2397 a_57417_n5344# a_50751_n19729# a_48951_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2398 a_46879_n2651# a_31953_n19727# a_46319_n1754# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2399 a_79182_n34390# a_65658_n29313# a_78344_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2400 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2401 a_89407_n20430# a_71281_n10073# a_88839_n20430# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2402 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2403 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2404 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2405 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2406 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2407 a_51151_n14215# a_50751_n19729# a_50629_n15112# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2408 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2409 a_100803_n20430# a_71281_n8397# a_100235_n20430# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2410 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2411 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2412 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2413 a_50629_n16009# a_83325_4421# a_83725_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2414 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2415 a_106501_n18620# a_71281_n8397# a_105933_n18620# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2416 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2417 a_114485_n29181# a_112559_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2418 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2419 a_87433_n6055# a_71281_n10073# a_86903_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2420 OUT a_35502_24538# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2421 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2422 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2423 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2424 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2425 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2426 a_55601_n28415# a_47819_n36322# a_39179_n19595# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2427 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2428 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2429 a_101641_n8770# a_71281_n8397# a_100803_n8770# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2430 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2431 a_77776_n34390# a_71366_n35156# a_71496_n36382# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2432 a_34347_n13316# a_31953_n19727# a_33787_n13316# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2433 a_67111_n13318# a_50751_n19729# a_66551_n12421# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2434 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2435 a_113037_n17715# a_71281_n8397# a_112507_n17715# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2436 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2437 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2438 a_96818_6405# a_94892_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2439 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2440 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2441 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2442 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2443 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2444 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2445 a_83141_n19525# a_71281_n10073# a_82573_n19525# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2446 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2447 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2448 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2449 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2450 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2451 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2452 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2453 VDD a_83153_10448# a_83683_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2454 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2455 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2456 a_95105_n14095# a_71281_n10073# a_94537_n14095# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2457 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2458 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2459 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2460 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2461 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X2462 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2463 a_63683_n16906# a_50751_n19729# a_63161_n17803# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2464 a_90245_n15000# a_71281_n10073# a_89407_n14095# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2465 a_88839_n6960# a_71281_n10073# a_88271_n6960# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2466 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2467 a_53675_7563# a_47819_11614# a_55601_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2468 a_90969_10448# a_89163_10388# a_89009_7563# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2469 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2470 VDD a_31699_20742# a_31699_20742# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2471 a_95943_n8770# a_71281_n10073# a_95105_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2472 a_112559_4481# a_100992_4421# a_114516_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2473 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2474 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2475 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2476 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2477 VSS a_36162_n36382# a_36562_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2478 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2479 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2480 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2481 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2482 a_89407_n1530# a_71281_n10073# a_88839_n1530# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2483 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2484 a_67422_n35156# a_65486_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2485 a_83725_6405# a_83325_4421# a_83153_10448# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2486 VSS a_59558_n29181# a_60080_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2487 a_81735_n19525# a_71281_n10073# a_81205_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2488 a_51151_n8932# a_50751_n19729# a_50629_n8932# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2489 a_40053_n8033# a_31953_n19727# a_39531_n8033# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2490 VDD a_83153_10448# a_83683_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2491 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2492 a_93969_n9675# a_71281_n10073# a_93131_n9675# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2493 a_53145_n8932# a_50751_n19729# a_52585_n8932# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2494 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2495 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2496 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X2497 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2498 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2499 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2500 a_112559_4481# a_100992_4421# a_114516_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2501 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2502 a_94537_n4245# a_71281_n10073# a_93969_n4245# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2503 a_30682_n36322# a_30152_n35156# a_30152_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2504 a_88839_n14095# a_71281_n10073# a_88271_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2505 a_35781_n19595# a_31953_n19727# a_35221_n19595# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2506 a_41487_n8033# a_31953_n19727# a_40965_n8033# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2507 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2508 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2509 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2510 a_35221_n7136# a_31953_n19727# a_34699_n8033# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2511 a_67422_n33224# a_65486_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2512 a_89407_n15905# a_71281_n10073# a_88839_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2513 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2514 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2515 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2516 a_112507_n17715# a_71281_n8397# a_112199_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2517 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2518 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2519 a_100803_n15905# a_71281_n8397# a_100235_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2520 a_36562_13546# a_36162_10388# a_36032_13546# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2521 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2522 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2523 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2524 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2525 a_55635_n36322# a_53829_n36382# a_53675_n27257# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2526 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2527 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2528 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2529 a_41660_19698# a_35502_24538# a_41100_20251# VSS nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X2530 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2531 a_65117_n17803# a_50751_n19729# a_64595_n18700# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2532 a_55601_4481# a_47819_11614# a_47991_4421# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2533 a_35502_24538# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2534 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2535 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2536 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2537 a_53829_n36382# a_59558_n29181# a_61484_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2538 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2539 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2540 a_60109_n36322# a_53699_n35156# a_53829_n36382# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2541 a_59411_n17803# a_50751_n19729# a_58851_n17803# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2542 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2543 a_83141_n6960# a_71281_n10073# a_82573_n6960# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2544 a_36562_11614# a_36162_10388# a_36032_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2545 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2546 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2547 a_33379_34007# IN_POS cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
X2548 a_59558_4481# a_59558_4481# a_61484_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2549 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2550 a_33249_35053# a_35502_24538# OUT VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2551 VDD a_65486_11614# a_73268_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2552 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2553 a_100235_n6960# a_71281_n8397# a_99667_n6960# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2554 a_83709_n13190# a_71281_n10073# a_83141_n13190# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2555 a_46319_n1754# a_31953_n19727# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2556 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2557 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2558 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2559 a_47753_n6239# a_31953_n19727# a_47231_n6239# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2560 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2561 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2562 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2563 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2564 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2565 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2566 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2567 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2568 a_81735_n3340# a_71281_n10073# a_81205_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2569 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2570 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2571 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2572 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2573 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2574 a_94892_4481# a_83325_4421# a_96849_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2575 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2576 a_99667_n15000# a_71281_n8397# a_98829_n15000# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2577 a_59411_n17803# a_50751_n19729# a_60285_n16009# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2578 a_60677_10448# a_47991_4421# a_60109_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2579 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2580 a_98829_n3340# a_71281_n8397# a_98299_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2581 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2582 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2583 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2584 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2585 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2586 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X2587 a_48313_n2651# a_31953_n19727# a_47753_n2651# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2588 a_111063_n15000# a_71281_n8397# a_110225_n15000# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2589 a_33787_n14213# a_31953_n19727# a_33265_n14213# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2590 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2591 a_59411_n2653# a_50751_n19729# a_58851_n1756# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2592 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2593 a_113037_n6960# a_71281_n8397# a_112199_n6960# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2594 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2595 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2596 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2597 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2598 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2599 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2600 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2601 a_45445_n5342# a_31953_n19727# a_44885_n5342# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2602 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2603 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2604 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2605 a_30152_10448# a_30324_4421# a_32128_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2606 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2607 a_94892_4481# a_83325_4421# a_96849_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2608 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2609 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2610 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2611 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2612 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2613 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2614 a_87433_n4245# a_71281_n10073# a_86903_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2615 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2616 a_43010_n36322# a_36032_n35156# a_42442_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2617 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2618 a_64243_n5344# a_50751_n19729# a_63683_n5344# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2619 a_71864_6405# a_65486_11614# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2620 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2621 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2622 a_93131_n13190# a_71281_n10073# a_92601_n16810# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2623 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2624 a_101641_n8770# a_71281_n8397# a_100803_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2625 a_88271_n13190# a_71281_n10073# a_87433_n13190# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2626 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2627 a_53145_n17803# a_50751_n19729# a_54019_n16009# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2628 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2629 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2630 a_71342_n30339# a_65486_n36322# a_73268_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2631 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2632 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2633 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2634 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2635 a_64243_n16009# a_50751_n19729# a_63683_n16009# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2636 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2637 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2638 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2639 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2640 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2641 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2642 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2643 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2644 a_45138_22884# a_35922_19591# a_44608_22884# VDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X2645 a_100820_10448# a_100820_10448# a_102756_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2646 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2647 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2648 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2649 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2650 a_31831_n5342# a_83325_n29313# a_83725_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2651 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2652 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2653 a_32128_n27257# a_30324_n30399# a_31284_n30339# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2654 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2655 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2656 a_40053_n3548# a_31953_n19727# a_39531_n3548# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2657 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2658 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2659 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2660 a_99667_n20430# a_71281_n8397# a_98829_n20430# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2661 a_102796_7563# a_100992_4421# a_56895_n16009# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2662 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2663 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2664 a_61515_n36322# a_47991_n29313# a_60677_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2665 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2666 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2667 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2668 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2669 a_93131_n3340# a_71281_n10073# a_92601_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2670 a_73302_12380# a_71496_10388# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2671 a_57977_n16009# a_50751_n19729# a_57417_n16009# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2672 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2673 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2674 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2675 a_111063_n20430# a_71281_n8397# a_110225_n20430# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2676 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2677 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2678 a_42047_n13316# a_31953_n19727# a_41487_n12419# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2679 a_100820_10448# a_100820_10448# a_102756_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2680 a_41487_n3548# a_31953_n19727# a_40965_n3548# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2681 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2682 a_31699_20742# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2683 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2684 a_37968_n34390# a_36162_n36382# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2685 a_52585_n13318# a_50751_n19729# a_52063_n14215# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2686 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2687 VDD a_31699_20742# a_35502_25545# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2688 a_65486_n35156# a_65658_n29313# a_67462_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2689 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2690 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2691 a_36530_n27257# a_30152_n36322# a_36008_n27257# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2692 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2693 a_106501_n21335# a_71281_n8397# a_105933_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2694 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2695 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2696 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2697 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2698 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2699 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2700 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2701 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2702 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2703 a_44363_n16007# a_45445_n19595# a_66058_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2704 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2705 a_85089_13546# a_83153_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2706 a_41100_20251# a_35502_24538# a_35502_24538# VSS nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X2707 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2708 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2709 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2710 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2711 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2712 a_105933_n6960# a_71281_n8397# a_105365_n6960# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2713 a_32913_n1754# a_31953_n19727# a_32353_n1754# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2714 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2715 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2716 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2717 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2718 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2719 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2720 a_106501_n1530# a_71281_n8397# a_105933_n1530# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2721 a_113081_n28415# a_112559_n29181# a_106830_n36382# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2722 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2723 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2724 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2725 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2726 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2727 a_85089_11614# a_83153_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2728 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2729 a_52635_34067# a_35502_24538# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2730 a_111063_n9675# a_71281_n8397# a_110225_n9675# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2731 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2732 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2733 a_89563_n35156# a_89163_n36382# a_89033_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2734 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2735 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2736 a_104527_n3340# a_71281_n8397# a_103997_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2737 a_77225_n29181# a_65658_n29313# a_79182_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2738 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2739 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2740 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2741 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2742 a_111631_n4245# a_71281_n8397# a_111063_n4245# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2743 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2744 a_52635_34067# a_35502_24538# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2745 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2746 a_79182_n36322# a_65658_n29313# a_78344_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2747 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2748 a_67111_n8932# a_50751_n19729# a_66551_n8932# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2749 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2750 a_54019_n14215# a_50751_n19729# a_53497_n14215# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2751 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2752 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2753 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2754 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2755 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2756 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2757 a_39179_n12419# a_31953_n19727# a_38619_n12419# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2758 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2759 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2760 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2761 a_89563_n33224# a_89163_n36382# a_71366_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2762 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2763 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2764 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2765 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2766 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2767 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2768 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2769 a_81735_n2435# a_71281_n10073# a_36032_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2770 a_99667_n15905# a_71281_n8397# a_98829_n15905# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2771 a_107198_6405# a_100820_11614# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2772 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2773 a_47819_10448# a_47991_4421# a_49795_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2774 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2775 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2776 VSS a_77225_n29181# a_77747_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2777 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2778 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2779 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2780 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2781 a_98829_n2435# a_71281_n8397# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2782 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2783 a_89563_12380# a_89163_10388# a_81205_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2784 a_67422_12380# a_65486_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2785 a_111063_n15905# a_71281_n8397# a_110225_n15905# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2786 a_71266_n4019# a_71266_n4019# a_75602_n4019# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X2787 a_77776_n36322# a_71366_n35156# a_71496_n36382# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2788 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2789 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2790 a_43010_10448# a_30324_4421# a_42442_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2791 a_61515_13546# a_47991_4421# a_60677_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2792 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2793 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2794 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2795 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2796 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2797 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2798 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2799 a_35781_n2651# a_31953_n19727# a_35221_n1754# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2800 a_32913_n18698# a_31953_n19727# a_32353_n17801# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2801 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2802 a_84017_n5150# a_71281_n10073# a_83709_n1530# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2803 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2804 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2805 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2806 I1N I1N a_75585_n8397# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X2807 a_85129_7563# a_83325_4421# a_50629_n16009# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2808 VSS a_106830_n36382# a_107230_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2809 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2810 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2811 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2812 a_110225_n17715# a_71281_n8397# a_109695_n16810# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2813 a_61515_11614# a_47991_4421# a_60677_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2814 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2815 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2816 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2817 a_43848_n34390# a_30324_n29313# a_43010_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2818 a_30152_10448# a_30152_10448# a_32088_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2819 a_110225_n15000# a_71281_n8397# a_109695_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2820 a_53675_7563# a_53829_10388# a_54229_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2821 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2822 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2823 a_35502_24538# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2824 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2825 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2826 a_89009_7563# a_83153_11614# a_90935_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2827 a_93969_n13190# a_71281_n10073# a_93131_n13190# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2828 a_78344_10448# a_65658_4421# a_77776_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2829 a_53699_13546# a_53829_10388# a_55635_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2830 a_36008_n30339# a_36162_n36382# a_36562_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2831 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2832 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2833 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2834 a_48391_5639# a_47991_5507# a_47819_11614# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2835 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2836 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2837 a_106676_n27257# a_106830_n36382# a_107230_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2838 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2839 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2840 a_41487_n13316# a_31953_n19727# a_40965_n14213# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2841 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2842 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2843 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2844 a_38619_n6239# a_31953_n19727# a_38097_n7136# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2845 VSS a_112559_4481# a_113081_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2846 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2847 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2848 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2849 a_89407_n14095# a_71281_n10073# a_88839_n14095# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2850 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2851 VSS a_53829_10388# a_54229_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2852 a_30152_10448# a_30152_10448# a_32088_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2853 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2854 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X2855 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2856 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2857 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2858 a_47753_n5342# a_31953_n19727# a_46879_n7136# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2859 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2860 a_100803_n14095# a_71281_n8397# a_100235_n14095# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2861 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2862 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2863 a_48313_n19595# a_31953_n19727# a_47753_n19595# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2864 a_35502_24538# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2865 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2866 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2867 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2868 a_71496_10388# a_77225_4481# a_79151_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2869 a_71496_n36382# a_77225_n29181# a_79151_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2870 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2871 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2872 a_93131_n2435# a_71281_n10073# a_71366_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2873 a_89009_n30339# a_83153_n36322# a_90935_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2874 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2875 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2876 VDD a_31699_20742# a_31699_20742# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2877 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2878 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2879 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2880 a_95443_n35156# a_83325_n29313# a_94892_n29181# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2881 a_60845_n15112# a_50751_n19729# a_60285_n15112# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2882 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2883 a_63683_n8035# a_50751_n19729# a_63161_n8932# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2884 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2885 a_106676_n27257# a_100820_n36322# a_108602_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2886 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2887 a_51711_n16906# a_50751_n19729# a_51151_n16906# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2888 a_44885_n13316# a_31953_n19727# a_44363_n13316# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2889 a_65677_n8932# a_50751_n19729# a_65117_n8035# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2890 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2891 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2892 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2893 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2894 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2895 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2896 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2897 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2898 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2899 VSS VSS VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X2900 a_95413_n5150# a_71281_n10073# a_95105_n1530# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2901 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2902 a_39179_n8930# a_100820_n36322# a_107198_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2903 a_110225_n20430# a_71281_n8397# a_71366_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2904 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2905 a_95443_n33224# a_83325_n29313# a_94892_n29181# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2906 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2907 a_60845_n7138# a_50751_n19729# a_60285_n7138# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2908 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2909 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2910 a_71366_13546# a_71496_10388# a_73302_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2911 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2912 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2913 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2914 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2915 a_54579_n15112# a_50751_n19729# a_54019_n15112# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2916 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2917 a_106830_n36382# a_103997_n8770# a_114516_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2918 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2919 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2920 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2921 a_93969_n3340# a_71281_n10073# a_93131_n3340# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2922 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2923 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2924 a_64243_n16906# a_50751_n19729# a_63683_n15112# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2925 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2926 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2927 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2928 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2929 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2930 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2931 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2932 a_37934_n28415# a_30152_n36322# a_30324_n30399# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2933 a_104527_n2435# a_71281_n8397# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2934 a_82573_n4245# a_71281_n10073# a_81735_n4245# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2935 a_35221_n15110# a_31953_n19727# a_34699_n16904# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2936 a_106830_n36382# a_103997_n8770# a_114516_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2937 VSS a_94892_4481# a_95414_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2938 a_111631_n15000# a_71281_n8397# a_111063_n15000# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2939 a_73268_7563# a_65486_11614# a_65658_4421# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2940 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2941 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2942 a_40053_n2651# a_31953_n19727# a_39531_n3548# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2943 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2944 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2945 a_67111_n19597# a_50751_n19729# a_66551_n18700# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2946 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2947 a_106809_n5150# a_100992_n29313# a_113110_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2948 a_99667_n4245# a_71281_n8397# a_98829_n4245# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2949 VDD a_31699_20742# a_35502_25545# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2950 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2951 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X2952 a_46319_n14213# a_31953_n19727# a_45797_n14213# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2953 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2954 a_57977_n16906# a_50751_n19729# a_57417_n15112# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2955 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2956 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2957 a_41487_n2651# a_31953_n19727# a_40965_n3548# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2958 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2959 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2960 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2961 VDD a_71281_n10073# a_89407_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2962 a_35221_n1754# a_31953_n19727# a_32913_n1754# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2963 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2964 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2965 a_43010_n36322# a_36032_n35156# a_42442_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2966 a_108636_12380# a_106830_10388# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2967 a_52585_n12421# a_50751_n19729# a_51711_n16009# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2968 a_57977_n5344# a_50751_n19729# a_57417_n5344# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2969 a_107230_10448# a_106830_10388# a_89033_13546# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2970 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2971 a_106809_n5150# a_100992_n29313# a_113110_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2972 a_38619_n18698# a_31953_n19727# a_38097_n19595# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2973 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2974 a_37934_5639# a_30152_11614# a_30324_5507# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2975 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2976 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2977 a_30152_n36322# a_30324_n30399# a_32128_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2978 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2979 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2980 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2981 a_51151_n4447# a_50751_n19729# a_50629_n4447# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2982 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2983 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2984 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2985 a_49755_n35156# a_47819_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2986 VSS a_41891_n29181# a_42413_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2987 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2988 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2989 a_44885_n8930# a_31953_n19727# a_44363_n8930# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2990 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2991 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2992 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2993 VSS a_112559_n29181# a_113081_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2994 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2995 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2996 a_88271_n6960# a_71281_n10073# a_87433_n6960# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2997 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2998 a_84547_n20430# a_71281_n10073# a_83709_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2999 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3000 a_46879_n8930# a_31953_n19727# a_46319_n8930# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3001 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3002 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3003 a_87433_n13190# a_71281_n10073# a_86903_n16810# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3004 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3005 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3006 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3007 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3008 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3009 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3010 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3011 a_95414_6405# a_94892_4481# a_94892_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3012 a_110225_n15905# a_71281_n8397# a_109695_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3013 a_107230_n34390# a_106830_n36382# a_103997_n8770# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3014 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3015 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3016 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3017 VSS a_94892_n29181# a_95414_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3018 a_49755_n33224# a_47819_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3019 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3020 a_111631_n20430# a_71281_n8397# a_111063_n20430# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3021 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3022 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3023 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3024 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3025 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3026 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3027 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3028 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3029 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3030 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3031 a_36032_n35156# a_36162_n36382# a_37968_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3032 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3033 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3034 VSS VSS VSS VSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X3035 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3036 a_43848_12380# a_36032_11614# a_43010_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3037 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3038 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3039 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3040 a_37968_n36322# a_36162_n36382# a_36008_n27257# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3041 VDD a_31699_20742# a_35502_24538# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3042 a_65117_n13318# a_50751_n19729# a_64595_n14215# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3043 VSS VSS VSS VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X3044 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3045 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3046 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3047 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3048 a_63683_n3550# a_50751_n19729# a_63161_n4447# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3049 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3050 VDD a_71281_n8397# a_100803_n1530# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3051 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3052 a_40053_n17801# a_31953_n19727# a_39531_n18698# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3053 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3054 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3055 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3056 a_59411_n13318# a_50751_n19729# a_58851_n13318# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3057 a_65117_n8035# a_50751_n19729# a_64595_n8035# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3058 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3059 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3060 a_36162_n36382# a_41891_n29181# a_43817_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3061 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3062 a_65677_n3550# a_50751_n19729# a_65117_n3550# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3063 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3064 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3065 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3066 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3067 a_47819_10448# a_47819_10448# a_49755_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3068 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3069 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3070 a_50751_n19729# a_71266_n4019# a_75602_n4978# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3071 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3072 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3073 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3074 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3075 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3076 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3077 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3078 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3079 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3080 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3081 a_83153_11614# a_83153_10448# a_85089_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3082 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3083 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3084 VDD a_83153_10448# a_83683_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3085 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3086 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3087 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3088 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3089 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3090 a_47819_10448# a_47819_10448# a_49755_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3091 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3092 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3093 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3094 a_107339_n8770# a_71281_n8397# a_106501_n8770# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3095 a_77225_n29181# a_65658_n29313# a_79182_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3096 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3097 a_45445_n19595# a_31953_n19727# a_44885_n19595# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3098 a_106830_10388# a_86903_n14095# a_114516_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3099 a_30682_n35156# a_30152_n35156# a_30152_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3100 a_34347_n14213# a_31953_n19727# a_35221_n16007# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3101 VDD a_83153_n35156# a_83683_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3102 a_58851_n8932# a_50751_n19729# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3103 VSS a_35502_25545# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3104 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3105 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3106 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3107 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3108 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3109 a_93969_n2435# a_71281_n10073# a_93131_n2435# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3110 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3111 a_99667_n14095# a_71281_n8397# a_98829_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3112 a_66551_n19597# a_50751_n19729# a_64243_n19597# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3113 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3114 a_55601_n27257# a_47819_n36322# a_47991_n29313# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3115 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3116 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3117 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3118 a_111063_n14095# a_71281_n8397# a_110225_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3119 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3120 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3121 a_30682_n33224# a_30152_n35156# a_30152_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3122 a_113037_n6055# a_71281_n8397# a_112507_n6055# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3123 a_55635_n35156# a_53829_n36382# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3124 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3125 VSS a_59558_4481# a_60080_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3126 a_111631_n15905# a_71281_n8397# a_111063_n15905# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3127 a_31699_17542# I1U a_30377_18342# VSS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X3128 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3129 a_38619_n5342# a_31953_n19727# a_38097_n5342# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3130 a_64243_n1756# a_65486_11614# a_71864_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3131 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3132 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3133 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3134 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3135 a_83153_10448# a_83325_4421# a_85129_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3136 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3137 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3138 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3139 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3140 a_95413_n16810# a_71281_n10073# a_95105_n13190# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3141 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3142 VCM a_33379_34007# cap_mim_2f0_m4m5_noshield c_width=9.8u c_length=9.8u
X3143 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3144 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3145 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3146 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3147 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3148 a_65486_10448# a_65486_10448# a_67422_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3149 a_60109_n35156# a_47991_n29313# a_59558_n29181# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3150 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3151 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3152 a_35502_24538# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3153 a_113110_n34390# a_103997_n8770# a_106830_n36382# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3154 a_36562_10448# a_36162_10388# a_33379_34917# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3155 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3156 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3157 a_55635_n33224# a_53829_n36382# a_53675_n30339# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3158 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3159 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3160 a_35502_25545# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3161 a_82573_n18620# a_71281_n10073# a_81735_n18620# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3162 a_111063_n3340# a_71281_n8397# a_110225_n3340# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3163 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3164 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3165 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3166 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3167 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3168 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3169 a_41891_n29181# a_30324_n29313# a_43848_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3170 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3171 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3172 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3173 a_46319_n8930# a_31953_n19727# a_45445_n5342# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3174 a_65486_10448# a_65486_10448# a_67422_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3175 a_60109_n33224# a_47991_n29313# a_59558_n29181# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3176 a_94537_n13190# a_71281_n10073# a_93969_n13190# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3177 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3178 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3179 a_43848_n36322# a_30324_n29313# a_43010_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3180 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3181 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3182 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3183 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3184 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3185 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3186 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3187 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3188 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3189 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3190 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3191 a_114485_7563# a_112559_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3192 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3193 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3194 a_60845_n7138# a_50751_n19729# a_60285_n6241# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3195 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3196 a_47819_n35156# a_47991_n29313# a_49795_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3197 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3198 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3199 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3200 a_65677_n14215# a_50751_n19729# a_65117_n14215# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3201 a_51151_n19597# a_50751_n19729# a_50629_n19597# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3202 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3203 a_51711_n8035# a_50751_n19729# a_51151_n8035# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3204 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3205 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3206 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3207 a_89163_10388# a_81205_n14095# a_96849_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3208 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3209 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3210 a_54229_12380# a_53829_10388# a_53699_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3211 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3212 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3213 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3214 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3215 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3216 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X3217 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3218 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3219 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3220 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3221 a_60285_n5344# a_50751_n19729# a_59411_n3550# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3222 VDD VDD VDD VDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X3223 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3224 a_65117_n3550# a_50751_n19729# a_64595_n3550# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3225 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3226 a_35221_n14213# a_31953_n19727# a_34699_n14213# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3227 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3228 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3229 a_34347_n19595# a_31953_n19727# a_33787_n18698# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3230 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3231 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X3232 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3233 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3234 a_101392_n30339# a_39179_n8930# a_100820_n36322# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3235 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3236 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3237 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3238 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3239 VSS a_35502_25545# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3240 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3241 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3242 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3243 VDD a_31699_20742# a_35502_24538# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3244 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3245 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3246 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3247 a_67462_7563# a_65658_4421# a_63161_n5344# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3248 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3249 a_52585_n7138# a_50751_n19729# a_52063_n8035# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3250 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3251 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3252 a_67111_n4447# a_50751_n19729# a_66551_n4447# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3253 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3254 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3255 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3256 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3257 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3258 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3259 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3260 a_54579_n7138# a_50751_n19729# a_54019_n7138# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3261 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3262 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3263 a_61515_n35156# a_53699_n35156# a_60677_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3264 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3265 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3266 a_94892_4481# a_94892_4481# a_96818_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3267 VSS a_35502_25545# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3268 a_71864_n28415# a_65486_n36322# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3269 a_100820_11614# a_100820_10448# a_102756_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3270 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3271 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3272 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3273 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3274 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3275 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3276 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3277 VSS a_35502_25545# a_35922_19591# VSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X3278 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3279 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3280 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3281 a_31284_n30339# a_30324_n30399# a_30724_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3282 a_107339_n8770# a_71281_n8397# a_106501_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3283 a_57977_n12421# a_100820_11614# a_107198_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3284 a_71896_12380# a_71496_10388# a_71366_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3285 a_47753_n16904# a_31953_n19727# a_47231_n16904# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3286 a_114485_n30339# a_112559_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3287 a_61515_n33224# a_53699_n35156# a_60677_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3288 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3289 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3290 a_95414_n29181# a_94892_n29181# a_94892_n29181# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3291 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3292 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3293 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3294 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3295 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3296 a_32913_n14213# a_31953_n19727# a_32353_n13316# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3297 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3298 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3299 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3300 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3301 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3302 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3303 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3304 a_85089_n34390# a_83153_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3305 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3306 a_50629_n16009# a_51711_n12421# a_83725_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3307 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3308 a_32913_n8930# a_31953_n19727# a_32353_n8930# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3309 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3310 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3311 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3312 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3313 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3314 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3315 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3316 a_65117_n12421# a_50751_n19729# a_64243_n16009# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3317 a_45138_24920# a_35922_19591# a_44608_24195# VDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X3318 a_110225_n6055# a_71281_n8397# a_109695_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3319 a_85089_10448# a_83153_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3320 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3321 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3322 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3323 a_63683_n2653# a_50751_n19729# a_63161_n2653# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3324 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3325 a_96818_7563# a_94892_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3326 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3327 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3328 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3329 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3330 a_59411_n13318# a_50751_n19729# a_58851_n12421# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3331 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3332 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3333 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3334 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3335 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3336 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X3337 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3338 a_65677_n2653# a_50751_n19729# a_65117_n2653# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3339 VDD VDD VDD VDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X3340 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3341 a_48951_4481# a_47991_5507# a_48391_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3342 a_110225_n14095# a_71281_n8397# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3343 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3344 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3345 a_79182_n35156# a_71366_n35156# a_78344_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3346 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3347 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3348 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3349 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3350 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3351 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3352 a_111063_n2435# a_71281_n8397# a_110225_n2435# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3353 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3354 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3355 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3356 a_79182_12380# a_71366_11614# a_78344_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3357 a_112199_n8770# a_71281_n8397# a_111631_n8770# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3358 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3359 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3360 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3361 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3362 a_60080_5639# a_59558_4481# a_53829_10388# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3363 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3364 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3365 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3366 a_60845_n2653# a_50751_n19729# a_60285_n1756# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3367 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3368 a_107230_n36322# a_106830_n36382# VCM VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3369 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3370 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3371 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3372 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3373 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3374 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3375 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3376 a_79182_n33224# a_71366_n35156# a_78344_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3377 a_51711_n3550# a_50751_n19729# a_51151_n3550# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3378 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3379 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3380 a_83725_7563# a_51711_n12421# a_83153_11614# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3381 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3382 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3383 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3384 a_33379_34007# a_36162_n36382# a_37968_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3385 a_77776_n35156# a_65658_n29313# a_77225_n29181# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3386 a_32353_n16904# a_31953_n19727# a_31831_n17801# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3387 VDD a_35922_19591# a_45706_22884# VDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X3388 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3389 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3390 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3391 a_90245_n3340# a_71281_n10073# a_89407_n3340# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3392 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3393 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3394 a_44363_n16007# a_65658_n29313# a_66058_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3395 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3396 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3397 a_33787_n19595# a_31953_n19727# a_32913_n16007# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3398 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3399 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3400 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3401 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3402 a_35781_n8930# a_31953_n19727# a_35221_n8930# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3403 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3404 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3405 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3406 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3407 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3408 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3409 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3410 a_77776_n33224# a_65658_n29313# a_77225_n29181# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3411 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3412 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3413 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3414 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3415 a_61515_10448# a_53699_11614# a_60677_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3416 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3417 a_113081_n27257# a_112559_n29181# a_112559_n29181# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3418 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3419 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3420 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3421 a_30152_11614# a_30324_5507# a_32128_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3422 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3423 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3424 a_59558_n29181# a_59558_n29181# a_61484_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3425 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3426 a_39179_n6239# a_31953_n19727# a_38619_n6239# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3427 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3428 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3429 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3430 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3431 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3432 VSS a_36162_n36382# a_36562_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3433 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3434 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3435 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3436 a_54019_n7138# a_50751_n19729# a_53497_n8035# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3437 VSS a_77225_4481# a_77747_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3438 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3439 a_82573_n21335# a_71281_n10073# a_81735_n21335# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3440 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3441 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3442 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3443 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3444 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3445 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3446 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3447 a_57417_n17803# a_50751_n19729# a_56895_n17803# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3448 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3449 a_53675_4481# a_53829_10388# a_54229_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3450 a_30152_11614# a_30152_10448# a_32088_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3451 a_90969_n34390# a_89163_n36382# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3452 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X3453 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3454 a_45138_24195# a_35922_19591# a_44608_24195# VDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X3455 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3456 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3457 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3458 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3459 a_100235_n19525# a_71281_n8397# a_99667_n19525# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3460 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3461 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3462 a_36008_n27257# a_36162_n36382# a_36562_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3463 VDD a_83153_n35156# a_83683_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3464 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3465 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3466 a_46879_n14213# a_31953_n19727# a_47753_n16007# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3467 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3468 a_75585_n10073# I1N VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X3469 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3470 a_71342_4481# a_65486_11614# a_73268_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3471 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3472 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3473 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3474 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3475 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3476 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3477 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3478 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3479 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3480 a_111631_n14095# a_71281_n8397# a_111063_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3481 VSS a_77225_n29181# a_77747_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3482 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3483 a_102796_4481# a_57977_n12421# a_56895_n16009# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3484 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3485 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3486 VDD a_100820_11614# a_108602_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3487 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3488 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3489 a_30324_5507# a_30152_11614# a_36530_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3490 a_52635_34067# a_35502_24538# a_33249_34067# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3491 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3492 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3493 a_52585_n18700# a_50751_n19729# a_52063_n18700# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3494 a_98829_n19525# a_71281_n8397# a_98299_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3495 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3496 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3497 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3498 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3499 VDD a_31699_20742# a_35502_25545# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3500 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3501 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3502 a_105365_n19525# a_71281_n8397# a_104527_n19525# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3503 a_113110_n36322# a_103997_n8770# a_106830_n36382# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3504 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3505 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3506 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3507 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3508 a_53829_10388# a_59558_4481# a_61484_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3509 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3510 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3511 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3512 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3513 a_65117_n2653# a_50751_n19729# a_64595_n3550# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3514 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3515 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3516 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3517 a_95105_n18620# a_71281_n10073# a_94537_n18620# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3518 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3519 a_71864_7563# a_65486_11614# a_71342_7563# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3520 a_66551_n7138# a_50751_n19729# a_66029_n8035# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3521 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3522 a_90245_n18620# a_71281_n10073# a_89407_n18620# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3523 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3524 a_41891_n29181# a_30324_n29313# a_43848_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3525 a_110225_n4245# a_71281_n8397# a_109695_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3526 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3527 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3528 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3529 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3530 a_31831_n5342# a_32913_n8930# a_83725_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3531 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3532 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3533 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3534 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3535 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3536 VDD a_71281_n8397# a_100803_n13190# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3537 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3538 VSS a_35502_25545# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3539 VDD a_71266_n4019# a_72596_n4019# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3540 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3541 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3542 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3543 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3544 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3545 a_45445_n19595# a_65486_n36322# a_71864_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3546 a_40613_n13316# a_31953_n19727# a_40053_n12419# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3547 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3548 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3549 VSS VSS VSS VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X3550 a_54579_n7138# a_50751_n19729# a_54019_n6241# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3551 a_108602_5639# a_100820_11614# a_57977_n12421# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3552 a_36530_5639# a_30152_11614# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3553 a_112199_n7865# a_71281_n8397# a_111631_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3554 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3555 a_88839_n18620# a_71281_n10073# a_88271_n18620# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3556 a_54019_n19597# a_50751_n19729# a_51711_n19597# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3557 a_40053_n13316# a_31953_n19727# a_39531_n14213# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3558 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3559 a_94537_n6960# a_71281_n10073# a_93969_n6960# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3560 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3561 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3562 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3563 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3564 a_108636_n34390# a_106830_n36382# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3565 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3566 a_43010_n36322# a_30324_n29313# a_42442_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3567 VSS a_35502_25545# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3568 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3569 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3570 a_30724_n29181# a_30324_n29313# a_30152_n35156# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3571 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3572 a_60109_13546# a_53699_11614# a_53829_10388# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3573 VDD a_31699_20742# a_35502_24538# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3574 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3575 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3576 a_35221_n8930# a_31953_n19727# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3577 a_38619_n15110# a_31953_n19727# a_38097_n15110# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3578 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3579 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3580 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3581 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3582 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3583 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3584 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3585 VDD a_71281_n8397# a_106501_n13190# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3586 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3587 a_90245_n3340# a_71281_n10073# a_89407_n2435# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3588 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3589 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3590 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3591 a_100992_n29313# a_100820_n36322# a_107198_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3592 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3593 a_102796_n28415# a_100992_n29313# a_38097_n5342# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3594 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3595 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3596 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3597 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3598 a_43010_n36322# a_30324_n29313# a_42442_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3599 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3600 a_60109_11614# a_53699_11614# a_53829_10388# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3601 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3602 a_83709_n8770# a_71281_n10073# a_83141_n8770# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3603 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3604 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3605 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3606 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3607 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3608 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3609 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3610 a_44885_n8033# a_31953_n19727# a_44363_n8930# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3611 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3612 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3613 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3614 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3615 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3616 a_46879_n8930# a_31953_n19727# a_46319_n8033# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3617 a_85129_4481# a_51711_n12421# a_50629_n16009# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3618 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3619 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3620 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3621 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3622 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3623 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3624 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3625 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3626 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3627 a_32913_n8930# a_83153_n36322# a_89531_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3628 a_37934_n27257# a_30152_n36322# a_30324_n29313# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3629 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3630 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3631 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3632 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3633 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3634 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3635 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3636 a_37968_n35156# a_36162_n36382# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3637 a_89407_n9675# a_71281_n10073# a_88839_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3638 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3639 a_41487_n18698# a_31953_n19727# a_40965_n18698# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3640 a_42047_n7136# a_31953_n19727# a_41487_n7136# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3641 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3642 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3643 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3644 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3645 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3646 VSS a_36162_10388# a_36562_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3647 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3648 a_77776_13546# a_71366_11614# a_71496_10388# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3649 a_55635_13546# a_53829_10388# a_53675_4481# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3650 a_48391_n29181# a_47991_n29313# a_47819_n35156# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3651 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3652 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3653 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3654 a_83153_n35156# a_83153_n35156# a_85089_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3655 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3656 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3657 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3658 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3659 a_33249_35053# a_35502_24538# OUT VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3660 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3661 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3662 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3663 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3664 a_37968_n33224# a_36162_n36382# a_36008_n30339# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3665 a_51711_n3550# a_50751_n19729# a_51151_n2653# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3666 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3667 a_85089_n36322# a_83153_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3668 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3669 VDD a_31699_20742# a_31699_20742# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3670 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3671 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3672 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3673 a_87433_n6960# a_71281_n10073# a_86903_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3674 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3675 a_107198_7563# a_100820_11614# a_106676_7563# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3676 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3677 a_77776_11614# a_71366_11614# a_71496_10388# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3678 a_55635_11614# a_53829_10388# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3679 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3680 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3681 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3682 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3683 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3684 a_44885_n18698# a_31953_n19727# a_44363_n19595# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3685 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3686 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3687 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3688 a_47819_11614# a_47819_10448# a_49755_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3689 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3690 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3691 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3692 a_71496_n36382# a_71366_n35156# a_79182_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3693 a_45445_n16007# a_31953_n19727# a_44885_n16007# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3694 a_95105_n8770# a_71281_n10073# a_94537_n8770# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3695 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3696 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3697 a_90935_n28415# a_83153_n36322# a_32913_n8930# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3698 a_53145_n17803# a_50751_n19729# a_52585_n17803# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3699 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3700 a_114516_n34390# a_100992_n29313# a_106809_n5150# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3701 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3702 VSS a_94892_n29181# a_95414_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3703 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3704 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3705 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3706 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3707 a_66551_n16009# a_50751_n19729# a_65677_n14215# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3708 a_39179_n5342# a_31953_n19727# a_38619_n5342# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3709 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3710 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3711 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3712 a_90245_n17715# a_71281_n10073# a_89715_n17715# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3713 a_52585_n1756# a_50751_n19729# a_51711_n5344# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3714 VDD a_71281_n8397# a_106501_n1530# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3715 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3716 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3717 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3718 a_54019_n6241# a_50751_n19729# a_53497_n6241# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3719 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3720 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3721 a_71496_n36382# a_71366_n35156# a_79182_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3722 a_32353_n4445# a_31953_n19727# a_31831_n4445# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3723 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3724 a_54579_n2653# a_50751_n19729# a_54019_n1756# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3725 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3726 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3727 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3728 a_47819_11614# a_47991_5507# a_49795_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3729 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3730 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3731 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3732 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3733 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3734 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3735 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3736 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3737 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3738 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3739 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3740 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3741 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3742 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3743 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3744 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3745 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3746 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3747 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3748 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3749 a_46319_n19595# a_31953_n19727# a_45445_n16007# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3750 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3751 a_73268_4481# a_65486_11614# a_65658_4421# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3752 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3753 VSS VSS VSS VSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X3754 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3755 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3756 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3757 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3758 a_33249_34067# a_35502_24538# a_52635_34067# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3759 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3760 a_31953_n19727# a_71266_n4019# a_75602_n3060# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3761 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3762 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3763 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3764 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3765 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3766 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3767 a_65486_11614# a_65486_10448# a_67422_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3768 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3769 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3770 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3771 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3772 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3773 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3774 a_43848_n35156# a_36032_n35156# a_43010_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3775 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3776 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3777 a_54197_n28415# a_47819_n36322# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3778 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3779 a_44885_n3548# a_31953_n19727# a_44363_n4445# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3780 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3781 a_48391_6405# a_47991_4421# a_47819_10448# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3782 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3783 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3784 VSS VSS VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X3785 a_46319_n8033# a_31953_n19727# a_45797_n8033# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3786 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3787 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3788 a_95105_n21335# a_71281_n10073# a_94537_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3789 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3790 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3791 a_89033_n35156# a_89163_n36382# a_90969_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3792 a_57417_n7138# a_50751_n19729# a_56895_n7138# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3793 a_46879_n3548# a_31953_n19727# a_46319_n3548# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3794 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3795 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3796 a_47753_n12419# a_31953_n19727# a_45445_n12419# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3797 VDD a_71281_n10073# a_89407_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3798 a_83709_n7865# a_71281_n10073# a_83141_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3799 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3800 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3801 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3802 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3803 a_51151_n16009# a_50751_n19729# a_50629_n16009# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3804 a_43848_n33224# a_36032_n35156# a_43010_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3805 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3806 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3807 a_77747_n29181# a_77225_n29181# a_77225_n29181# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3808 a_90969_n36322# a_89163_n36382# a_89009_n27257# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3809 a_111631_n6960# a_71281_n8397# a_111063_n6960# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3810 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3811 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3812 a_66551_n6241# a_50751_n19729# a_66029_n6241# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3813 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3814 VDD a_31699_20742# a_35502_25545# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3815 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3816 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3817 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3818 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3819 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3820 a_108602_n28415# a_100820_n36322# a_39179_n8930# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3821 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3822 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3823 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3824 a_83709_n15000# a_71281_n10073# a_83141_n15000# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3825 VDD a_71266_n4019# a_72596_n4978# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3826 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3827 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3828 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3829 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3830 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3831 a_59411_n8932# a_50751_n19729# a_58851_n8035# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3832 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3833 a_66016_13546# a_65486_10448# a_65486_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3834 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3835 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3836 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3837 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3838 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3839 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3840 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3841 a_67111_n15112# a_50751_n19729# a_66551_n14215# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3842 a_88839_n21335# a_71281_n10073# a_88271_n21335# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3843 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3844 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3845 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3846 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3847 a_65117_n18700# a_50751_n19729# a_64595_n18700# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3848 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3849 VSS a_94892_4481# a_95414_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3850 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3851 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3852 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3853 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3854 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3855 a_100803_n8770# a_71281_n8397# a_100235_n8770# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3856 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3857 a_105933_n19525# a_71281_n8397# a_105365_n19525# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3858 a_105365_n4245# a_71281_n8397# a_104527_n4245# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3859 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3860 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3861 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3862 a_66016_11614# a_65486_10448# a_65486_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3863 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3864 a_59411_n19597# a_50751_n19729# a_58851_n18700# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3865 a_42047_n17801# a_31953_n19727# a_41487_n17801# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3866 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3867 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3868 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3869 a_30152_n35156# a_30324_n29313# a_32128_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3870 a_38619_n14213# a_31953_n19727# a_38097_n15110# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3871 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3872 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3873 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3874 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3875 a_35922_19591# a_35502_25545# VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X3876 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3877 a_93131_n17715# a_71281_n10073# a_92601_n16810# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3878 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X3879 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X3880 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3881 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3882 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3883 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3884 VSS a_112559_n29181# a_113081_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3885 a_93131_n15000# a_71281_n10073# a_92601_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3886 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3887 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3888 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3889 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3890 a_88271_n15000# a_71281_n10073# a_87433_n15000# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3891 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3892 a_31699_19142# I1U a_30377_19942# VSS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X3893 a_106501_n9675# a_71281_n8397# a_105933_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3894 a_83153_n35156# a_83325_n29313# a_85129_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3895 a_104527_n19525# a_71281_n8397# a_103997_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3896 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3897 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3898 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3899 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3900 a_32353_n12419# a_31953_n19727# a_31831_n13316# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3901 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3902 a_95105_n7865# a_71281_n10073# a_94537_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3903 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3904 a_54019_n1756# a_50751_n19729# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3905 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3906 a_83709_n20430# a_71281_n10073# a_83141_n20430# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3907 a_37968_12380# a_36162_10388# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3908 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3909 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3910 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3911 a_89407_n18620# a_71281_n10073# a_88839_n18620# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3912 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3913 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X3914 a_83683_13546# a_83153_10448# a_83153_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3915 a_95414_7563# a_94892_4481# a_89163_10388# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3916 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3917 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3918 a_100803_n18620# a_71281_n8397# a_100235_n18620# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3919 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3920 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3921 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3922 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3923 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3924 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3925 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3926 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3927 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3928 a_108636_n36322# a_106830_n36382# a_106676_n27257# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3929 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3930 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3931 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3932 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3933 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3934 a_72596_n4019# a_71266_n4019# a_71266_n4019# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X3935 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3936 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3937 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3938 a_42413_n28415# a_41891_n29181# a_36162_n36382# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3939 a_41891_n29181# a_41891_n29181# a_43817_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3940 a_37934_6405# a_30152_11614# a_30324_5507# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3941 a_83683_11614# a_83153_10448# a_83153_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3942 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3943 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3944 a_106830_n36382# a_112559_n29181# a_114485_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3945 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3946 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3947 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3948 a_39179_n18698# a_31953_n19727# a_38619_n17801# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3949 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3950 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3951 a_60845_n17803# a_50751_n19729# a_60285_n16906# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3952 a_32913_n8033# a_31953_n19727# a_32353_n8033# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3953 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3954 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3955 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3956 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3957 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3958 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3959 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3960 a_57417_n13318# a_50751_n19729# a_56895_n13318# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3961 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3962 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3963 a_93131_n20430# a_71281_n10073# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3964 VSS VSS VSS VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X3965 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3966 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3967 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3968 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3969 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3970 a_88271_n20430# a_71281_n10073# a_87433_n20430# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3971 a_60285_n17803# a_50751_n19729# a_59763_n18700# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3972 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3973 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3974 VDD a_30152_n36322# a_37934_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3975 a_94892_n29181# a_94892_n29181# a_96818_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3976 a_71864_n27257# a_65486_n36322# a_71342_n27257# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3977 VDD a_71281_n10073# a_83709_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3978 a_46319_n3548# a_31953_n19727# a_45797_n3548# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3979 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3980 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3981 a_107230_n35156# a_106830_n36382# a_103997_n8770# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3982 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3983 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3984 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3985 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3986 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3987 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3988 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3989 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3990 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3991 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3992 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3993 a_66551_n1756# a_50751_n19729# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3994 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3995 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3996 a_112199_n1530# a_71281_n8397# a_111631_n1530# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3997 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3998 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3999 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4000 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4001 a_54579_n17803# a_50751_n19729# a_54019_n16906# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4002 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4003 a_31284_n30339# a_30324_n29313# a_30724_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4004 a_36032_n35156# a_36162_n36382# a_37968_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4005 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4006 VDD a_31699_20742# a_35502_24538# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4007 a_64243_n16906# a_50751_n19729# a_63683_n16906# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4008 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4009 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4010 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4011 a_33787_n7136# a_31953_n19727# a_33265_n8033# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4012 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4013 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4014 a_107230_n33224# a_106830_n36382# a_89033_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4015 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4016 a_48313_n4445# a_31953_n19727# a_47753_n4445# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4017 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4018 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4019 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4020 a_66551_n15112# a_50751_n19729# a_66029_n16906# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4021 a_59411_n3550# a_50751_n19729# a_58851_n3550# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4022 a_82573_n6960# a_71281_n10073# a_81735_n6960# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4023 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4024 VSS I1N a_72603_n8397# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X4025 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4026 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4027 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4028 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4029 a_65677_n19597# a_50751_n19729# a_65117_n19597# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4030 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4031 a_45445_n8033# a_31953_n19727# a_44885_n7136# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4032 a_114485_4481# a_112559_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4033 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4034 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4035 a_83709_n15905# a_71281_n10073# a_83141_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4036 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4037 a_99667_n6960# a_71281_n8397# a_98829_n6960# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4038 a_36032_n36322# a_36162_n36382# a_37968_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4039 a_83153_n35156# a_83153_n35156# a_85089_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4040 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4041 a_64243_n8035# a_50751_n19729# a_63683_n7138# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4042 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4043 a_60080_n28415# a_59558_n29181# a_53829_n36382# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4044 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4045 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4046 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4047 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4048 a_113037_n20430# a_71281_n8397# a_112199_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4049 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4050 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4051 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4052 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4053 a_35781_n8930# a_31953_n19727# a_35221_n8033# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4054 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X4055 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4056 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4057 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4058 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4059 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4060 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4061 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4062 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4063 a_57977_n16906# a_50751_n19729# a_57417_n16906# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4064 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4065 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4066 a_35221_n19595# a_31953_n19727# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4067 a_65658_4421# a_65486_11614# a_71864_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4068 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4069 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4070 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4071 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4072 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4073 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4074 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4075 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4076 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4077 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4078 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4079 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4080 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4081 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4082 a_100803_n7865# a_71281_n8397# a_100235_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4083 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4084 OUT a_35502_24538# a_33249_35053# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4085 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4086 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4087 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4088 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4089 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4090 a_39179_n19595# a_47819_n36322# a_54197_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4091 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4092 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4093 a_88839_n8770# a_71281_n10073# a_88271_n8770# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4094 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4095 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4096 VDD a_83153_n35156# a_83683_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4097 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4098 VDD a_71281_n10073# a_95105_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4099 a_114516_n36322# a_100992_n29313# a_106809_n5150# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4100 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4101 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4102 a_93131_n15905# a_71281_n10073# a_92601_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4103 a_113110_12380# a_100992_4421# a_112559_4481# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4104 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4105 a_89407_n3340# a_71281_n10073# a_88839_n3340# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4106 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4107 a_67462_4481# a_64243_n1756# a_63161_n5344# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4108 a_88271_n15905# a_71281_n10073# a_87433_n15905# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4109 a_46274_24920# a_35922_19591# a_45706_24920# VDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X4110 a_48349_12380# a_47819_10448# a_47819_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4111 a_44885_n2651# a_31953_n19727# a_44363_n2651# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4112 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4113 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4114 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4115 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4116 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4117 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4118 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4119 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4120 a_57417_n6241# a_50751_n19729# a_56895_n7138# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4121 a_46879_n2651# a_31953_n19727# a_46319_n2651# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4122 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4123 a_93969_n15000# a_71281_n10073# a_93131_n15000# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4124 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4125 a_89163_10388# a_94892_4481# a_96818_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4126 VSS a_59558_4481# a_60080_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4127 VDD a_83153_n35156# a_83683_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4128 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4129 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4130 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4131 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4132 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4133 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4134 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4135 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4136 a_83153_11614# a_51711_n12421# a_85129_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4137 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4138 a_51151_n15112# a_50751_n19729# a_50629_n15112# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4139 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4140 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4141 a_33249_35053# a_35502_24538# OUT VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4142 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4143 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4144 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4145 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4146 a_102756_13546# a_100820_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4147 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4148 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4149 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4150 a_32913_n18698# a_31953_n19727# a_32353_n18698# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4151 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4152 a_42047_n2651# a_31953_n19727# a_41487_n1754# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4153 a_113110_n35156# a_100992_n29313# a_112559_n29181# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4154 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4155 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4156 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4157 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4158 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4159 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4160 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4161 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4162 a_32913_n3548# a_31953_n19727# a_32353_n3548# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4163 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4164 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4165 a_34347_n14213# a_31953_n19727# a_33787_n14213# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4166 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4167 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4168 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4169 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4170 a_36162_n36382# a_36032_n35156# a_43848_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4171 a_102756_11614# a_100820_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4172 a_50629_n16009# a_83325_4421# a_83725_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4173 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4174 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4175 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4176 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4177 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4178 a_113110_n33224# a_100992_n29313# a_112559_n29181# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4179 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4180 a_35502_25545# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4181 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4182 a_83141_n8770# a_71281_n10073# a_82573_n8770# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4183 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4184 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4185 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4186 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4187 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4188 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4189 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4190 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4191 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4192 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4193 VSS a_35502_25545# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4194 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4195 a_100235_n8770# a_71281_n8397# a_99667_n8770# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4196 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4197 a_36162_n36382# a_36032_n35156# a_43848_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4198 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4199 a_71366_n36322# a_89163_n36382# a_90969_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4200 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4201 a_96818_4481# a_94892_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4202 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4203 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4204 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4205 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4206 a_54019_n16009# a_50751_n19729# a_53145_n14215# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4207 a_63683_n17803# a_50751_n19729# a_63161_n17803# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4208 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4209 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4210 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4211 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4212 a_93969_n20430# a_71281_n10073# a_93131_n20430# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4213 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4214 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4215 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4216 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4217 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4218 a_81735_n6055# a_71281_n10073# a_81205_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4219 a_99667_n18620# a_71281_n8397# a_98829_n18620# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4220 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4221 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4222 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4223 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4224 a_95414_n30339# a_94892_n29181# a_89163_n36382# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4225 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4226 a_38097_n5342# a_39179_n8930# a_101392_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4227 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4228 a_72603_n9297# I1N a_71281_n10073# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X4229 a_111063_n18620# a_71281_n8397# a_110225_n18620# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4230 a_98829_n6055# a_71281_n8397# a_98299_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4231 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4232 a_89407_n21335# a_71281_n10073# a_88839_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4233 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4234 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4235 VSS a_35502_25545# a_35502_25545# VSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X4236 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4237 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4238 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4239 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4240 a_113037_n8770# a_71281_n8397# a_112199_n8770# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4241 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4242 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4243 a_100803_n21335# a_71281_n8397# a_100235_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4244 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4245 a_46274_23609# a_35922_19591# a_45706_24195# VDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X4246 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4247 a_100992_4421# a_100820_11614# a_107198_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4248 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4249 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4250 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4251 a_35221_n8033# a_31953_n19727# a_34699_n8033# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4252 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4253 a_83725_4481# a_83325_4421# a_83153_10448# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4254 a_106501_n19525# a_71281_n8397# a_105933_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4255 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4256 a_35781_n4445# a_31953_n19727# a_35221_n3548# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4257 a_60109_10448# a_47991_4421# a_59558_4481# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4258 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4259 a_87433_n6055# a_71281_n10073# a_86903_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4260 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4261 a_53145_n13318# a_50751_n19729# a_52585_n13318# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4262 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4263 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4264 a_101111_n6055# a_71281_n8397# a_100803_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4265 a_72596_n4978# a_71266_n4019# a_31953_n19727# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X4266 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4267 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4268 a_73268_n28415# a_65486_n36322# a_45445_n19595# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4269 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4270 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4271 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4272 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4273 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4274 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4275 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4276 a_33249_35053# a_35502_24538# OUT VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4277 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4278 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4279 a_52635_34067# a_35502_24538# a_33249_34067# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4280 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4281 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4282 a_83709_n1530# a_71281_n10073# a_83141_n1530# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4283 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4284 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4285 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4286 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4287 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4288 a_63683_n8932# a_50751_n19729# a_63161_n8932# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4289 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4290 a_96818_n29181# a_94892_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4291 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4292 a_57417_n12421# a_50751_n19729# a_56895_n13318# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4293 a_42442_12380# a_30324_4421# a_41891_4481# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4294 a_41487_n15110# a_31953_n19727# a_40965_n16904# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4295 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4296 a_65677_n8932# a_50751_n19729# a_65117_n8932# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4297 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4298 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4299 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4300 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4301 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4302 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4303 a_35502_24538# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4304 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4305 a_88839_n7865# a_71281_n10073# a_88271_n7865# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4306 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4307 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4308 a_87433_n17715# a_71281_n10073# a_86903_n16810# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4309 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4310 a_46319_n2651# a_31953_n19727# a_45797_n3548# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4311 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4312 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4313 a_47753_n7136# a_31953_n19727# a_47231_n8033# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4314 a_57417_n1756# a_50751_n19729# a_56895_n2653# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4315 a_93131_n6055# a_71281_n10073# a_92601_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4316 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4317 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4318 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4319 a_87433_n15000# a_71281_n10073# a_86903_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4320 a_89407_n2435# a_71281_n10073# a_88839_n2435# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4321 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4322 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4323 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4324 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4325 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4326 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4327 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4328 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4329 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4330 a_30324_n30399# a_30152_n36322# a_36530_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4331 a_85089_n35156# a_83153_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4332 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4333 a_93969_n15905# a_71281_n10073# a_93131_n15905# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4334 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4335 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4336 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4337 a_71342_7563# a_65486_11614# a_73268_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4338 a_55635_10448# a_53829_10388# a_53675_7563# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4339 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4340 a_77776_10448# a_65658_4421# a_77225_4481# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4341 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4342 a_44885_n15110# a_31953_n19727# a_44363_n15110# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4343 a_102796_n27257# a_39179_n8930# a_38097_n5342# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4344 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4345 a_59411_n2653# a_50751_n19729# a_58851_n2653# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4346 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4347 a_61484_5639# a_59558_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4348 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4349 a_85089_n33224# a_83153_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4350 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4351 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4352 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4353 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4354 a_105933_n8770# a_71281_n8397# a_105365_n8770# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4355 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4356 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4357 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4358 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4359 a_64243_n6241# a_50751_n19729# a_63683_n6241# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4360 a_48951_4481# a_47991_4421# a_48391_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4361 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4362 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4363 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4364 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4365 VDD a_31699_20742# a_35502_24538# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4366 a_106501_n3340# a_71281_n8397# a_105933_n3340# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4367 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4368 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4369 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4370 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4371 a_60080_6405# a_59558_4481# a_59558_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4372 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4373 a_95105_n1530# a_71281_n10073# a_94537_n1530# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4374 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4375 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4376 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4377 a_104527_n6055# a_71281_n8397# a_103997_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4378 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4379 a_112199_n13190# a_71281_n8397# a_111631_n13190# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4380 a_71864_4481# a_65486_11614# a_71342_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4381 a_83141_n7865# a_71281_n10073# a_82573_n7865# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4382 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4383 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4384 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4385 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4386 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4387 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4388 a_87433_n20430# a_71281_n10073# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4389 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4390 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4391 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4392 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4393 a_100235_n7865# a_71281_n8397# a_99667_n7865# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4394 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4395 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4396 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4397 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4398 a_83709_n14095# a_71281_n10073# a_83141_n14095# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4399 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4400 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4401 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4402 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4403 a_40053_n18698# a_31953_n19727# a_39531_n18698# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4404 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4405 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4406 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4407 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4408 a_81735_n4245# a_71281_n10073# a_81205_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4409 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4410 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4411 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4412 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4413 a_42047_n13316# a_31953_n19727# a_41487_n13316# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4414 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4415 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4416 a_41487_n4445# a_31953_n19727# a_40965_n6239# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4417 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4418 a_35221_n3548# a_31953_n19727# a_34699_n3548# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4419 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4420 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4421 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4422 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4423 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4424 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4425 a_98829_n4245# a_71281_n8397# a_98299_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4426 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4427 a_52585_n14215# a_50751_n19729# a_52063_n14215# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4428 a_57977_n8035# a_50751_n19729# a_57417_n7138# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4429 a_67462_n28415# a_65658_n29313# a_44363_n16007# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4430 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4431 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4432 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4433 a_113037_n8770# a_71281_n8397# a_112199_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4434 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4435 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4436 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4437 VSS a_77225_4481# a_77747_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4438 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4439 a_95943_n17715# a_71281_n10073# a_95413_n16810# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4440 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4441 a_84547_n3340# a_71281_n10073# a_83709_n3340# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4442 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4443 a_33249_34067# a_35502_24538# a_52635_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4444 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4445 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4446 a_90935_n27257# a_83153_n36322# a_83325_n29313# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4447 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4448 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4449 a_95943_n15000# a_71281_n10073# a_95105_n15000# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4450 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4451 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4452 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4453 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4454 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4455 a_93131_n14095# a_71281_n10073# IBPOUT VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4456 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4457 a_110225_n18620# a_71281_n8397# a_109695_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4458 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4459 a_32913_n3548# a_31953_n19727# a_32353_n2651# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4460 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4461 a_90969_n35156# a_89163_n36382# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4462 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4463 a_88271_n14095# a_71281_n10073# a_87433_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4464 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4465 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4466 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4467 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4468 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4469 a_65117_n8932# a_50751_n19729# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4470 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4471 a_59558_4481# a_59558_4481# a_61484_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4472 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4473 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4474 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4475 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4476 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4477 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4478 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4479 a_90969_12380# a_89163_10388# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4480 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4481 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4482 a_65658_n29313# a_65486_n36322# a_71864_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4483 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4484 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4485 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4486 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4487 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4488 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4489 a_94537_n15000# a_71281_n10073# a_93969_n15000# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4490 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4491 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4492 a_90969_n33224# a_89163_n36382# a_89009_n30339# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4493 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4494 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4495 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4496 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4497 VDD a_100820_11614# a_108602_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4498 a_30324_5507# a_30152_11614# a_36530_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4499 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4500 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4501 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4502 a_54019_n15112# a_50751_n19729# a_53497_n16906# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4503 a_99667_n21335# a_71281_n8397# a_98829_n21335# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4504 a_30724_n30339# a_30324_n30399# a_30152_n36322# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4505 a_39179_n14213# a_31953_n19727# a_38619_n13316# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4506 a_79151_n28415# a_77225_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4507 a_87433_n15905# a_71281_n10073# a_86903_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4508 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4509 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4510 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4511 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4512 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4513 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4514 a_93131_n4245# a_71281_n10073# a_92601_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4515 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4516 a_33787_n1754# a_31953_n19727# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4517 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4518 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4519 a_66016_10448# a_65486_10448# a_65486_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4520 a_111063_n21335# a_71281_n8397# a_110225_n21335# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4521 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4522 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4523 a_35781_n17801# a_31953_n19727# a_35221_n16904# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4524 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4525 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4526 a_60285_n13318# a_50751_n19729# a_59763_n14215# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4527 VSS VSS VSS VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X4528 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4529 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4530 a_45445_n1754# a_31953_n19727# a_44885_n1754# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4531 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4532 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4533 a_83141_n13190# a_71281_n10073# a_82573_n13190# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4534 a_100803_n1530# a_71281_n8397# a_100235_n1530# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4535 a_83725_n28415# a_32913_n8930# a_83153_n36322# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4536 a_95943_n20430# a_71281_n10073# a_95105_n20430# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4537 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4538 a_54197_n27257# a_47819_n36322# a_53675_n27257# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4539 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4540 a_64243_n1756# a_50751_n19729# a_63683_n1756# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4541 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4542 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4543 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4544 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4545 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4546 VDD a_65486_n36322# a_73268_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4547 a_95943_n3340# a_71281_n10073# a_95105_n3340# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4548 a_35781_n2651# a_31953_n19727# a_35221_n2651# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4549 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4550 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4551 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4552 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4553 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4554 a_107198_4481# a_100820_11614# a_106676_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4555 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4556 a_105933_n7865# a_71281_n8397# a_105365_n7865# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4557 a_53145_n13318# a_50751_n19729# a_52585_n12421# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4558 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4559 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4560 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4561 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4562 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4563 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4564 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4565 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4566 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4567 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4568 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4569 a_81735_n13190# a_71281_n10073# a_81205_n16810# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4570 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4571 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4572 a_35502_25545# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4573 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4574 a_83325_n29313# a_83153_n36322# a_89531_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4575 a_106501_n2435# a_71281_n8397# a_105933_n2435# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4576 a_94537_n20430# a_71281_n10073# a_93969_n20430# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4577 a_108602_6405# a_100820_11614# a_57977_n12421# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4578 a_36530_6405# a_30152_11614# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4579 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4580 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4581 a_49795_5639# a_47991_4421# a_48951_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4582 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4583 a_32128_n29181# a_30324_n30399# a_31284_n30339# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4584 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4585 a_108602_n27257# a_100820_n36322# a_100992_n29313# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4586 a_49755_13546# a_47819_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4587 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4588 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4589 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4590 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4591 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4592 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4593 VDD a_71266_n4019# a_72596_n3060# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X4594 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4595 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4596 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4597 a_108636_n35156# a_106830_n36382# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4598 a_111631_n18620# a_71281_n8397# a_111063_n18620# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4599 a_104527_n4245# a_71281_n8397# a_103997_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4600 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4601 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4602 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4603 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4604 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4605 a_41487_n14213# a_31953_n19727# a_40965_n14213# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4606 a_48391_n30339# a_39179_n19595# a_47819_n36322# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4607 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4608 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4609 a_38619_n7136# a_31953_n19727# a_38097_n7136# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4610 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4611 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4612 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4613 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4614 a_84017_n17715# a_81205_n14095# a_95443_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4615 a_83683_10448# a_83153_10448# a_83153_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4616 a_60677_10448# a_47991_4421# a_60109_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4617 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4618 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4619 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4620 a_49755_11614# a_47819_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4621 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4622 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4623 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4624 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4625 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4626 a_36530_n29181# a_30152_n36322# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4627 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4628 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4629 a_108636_n33224# a_106830_n36382# a_106676_n30339# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4630 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4631 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4632 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4633 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4634 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4635 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4636 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4637 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4638 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4639 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4640 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4641 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4642 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4643 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4644 a_84017_n17715# a_81205_n14095# a_95443_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4645 a_51711_n8932# a_50751_n19729# a_51151_n8932# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4646 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4647 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4648 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4649 a_51711_n18700# a_50751_n19729# a_51151_n17803# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4650 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4651 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4652 a_44885_n14213# a_31953_n19727# a_44363_n15110# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4653 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4654 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4655 a_83153_n36322# a_32913_n8930# a_85129_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4656 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4657 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4658 a_95943_n18620# a_71281_n10073# a_95105_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4659 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4660 a_110225_n6960# a_71281_n8397# a_109695_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4661 a_84547_n3340# a_71281_n10073# a_83709_n2435# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4662 a_88271_n8770# a_71281_n10073# a_87433_n8770# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4663 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4664 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4665 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4666 a_60845_n8932# a_50751_n19729# a_60285_n8035# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4667 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4668 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4669 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4670 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4671 VSS I1N a_72603_n10073# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X4672 a_110225_n17715# a_71281_n8397# a_109695_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4673 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4674 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4675 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4676 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4677 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4678 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4679 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4680 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4681 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4682 a_93969_n14095# a_71281_n10073# a_93131_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4683 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4684 a_83153_n36322# a_83153_n35156# a_85089_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4685 a_90935_5639# a_83153_11614# a_51711_n12421# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4686 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4687 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4688 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4689 a_94537_n15905# a_71281_n10073# a_93969_n15905# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4690 a_71266_n4019# I1N a_75585_n9297# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X4691 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4692 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X4693 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4694 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4695 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4696 a_60285_n7138# a_50751_n19729# a_59763_n8035# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4697 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4698 a_42413_n27257# a_41891_n29181# a_41891_n29181# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4699 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4700 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4701 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4702 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4703 a_35221_n16007# a_31953_n19727# a_34347_n17801# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4704 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4705 a_47819_10448# a_47991_4421# a_49795_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4706 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4707 a_67111_n19597# a_50751_n19729# a_66551_n19597# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4708 a_101641_n3340# a_71281_n8397# a_100803_n3340# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4709 a_66058_5639# a_64243_n1756# a_65486_11614# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4710 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4711 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4712 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4713 OUT a_35502_24538# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4714 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4715 a_83153_n36322# a_83153_n35156# a_85089_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4716 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4717 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4718 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4719 a_89163_n36382# a_94892_n29181# a_96818_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4720 a_31699_20742# I1U a_30377_19942# VSS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X4721 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4722 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4723 a_35221_n2651# a_31953_n19727# a_34699_n3548# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4724 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4725 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4726 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4727 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4728 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4729 VSS a_94892_4481# a_95414_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4730 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4731 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4732 a_114516_n35156# a_103997_n8770# a_106809_n5150# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4733 a_63683_n13318# a_50751_n19729# a_63161_n13318# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4734 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4735 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4736 a_57977_n6241# a_50751_n19729# a_57417_n6241# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4737 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4738 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4739 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4740 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4741 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4742 a_38619_n19595# a_31953_n19727# a_38097_n19595# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4743 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4744 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4745 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4746 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4747 a_31699_20742# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4748 a_51151_n5344# a_50751_n19729# a_31284_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4749 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4750 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4751 a_88839_n1530# a_71281_n10073# a_88271_n1530# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4752 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4753 a_95943_n3340# a_71281_n10073# a_95105_n2435# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4754 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4755 a_110225_n21335# a_71281_n8397# a_109695_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4756 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4757 a_77747_n30339# a_77225_n29181# a_71496_n36382# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4758 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4759 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4760 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4761 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4762 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4763 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4764 a_114516_n33224# a_103997_n8770# a_106809_n5150# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4765 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4766 a_46879_n13316# a_31953_n19727# a_46319_n12419# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4767 a_48391_7563# a_47991_5507# a_47819_11614# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4768 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4769 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4770 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4771 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4772 VDD a_47819_n36322# a_55601_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4773 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4774 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4775 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4776 a_93969_n4245# a_71281_n10073# a_93131_n4245# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4777 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4778 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4779 a_32913_n16904# a_31953_n19727# a_32353_n15110# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4780 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4781 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4782 a_60080_n27257# a_59558_n29181# a_59558_n29181# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4783 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4784 a_42047_n8930# a_31953_n19727# a_41487_n8930# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4785 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4786 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4787 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4788 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4789 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4790 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4791 a_47753_n1754# a_31953_n19727# a_45445_n1754# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4792 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4793 a_71496_n36382# a_77225_n29181# a_79151_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4794 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4795 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4796 VDD a_83153_n36322# a_90935_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4797 a_102756_10448# a_100820_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4798 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4799 a_95414_4481# a_94892_4481# a_94892_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4800 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4801 a_40613_n17801# a_31953_n19727# a_40053_n17801# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4802 VDD a_31699_20742# a_31699_20742# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4803 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4804 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4805 a_65117_n14215# a_50751_n19729# a_64595_n14215# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4806 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4807 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4808 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4809 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4810 a_63683_n4447# a_50751_n19729# a_63161_n4447# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4811 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4812 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4813 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4814 a_59411_n14215# a_50751_n19729# a_58851_n14215# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4815 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4816 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4817 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4818 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4819 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4820 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4821 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4822 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4823 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4824 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4825 a_60285_n12421# a_50751_n19729# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4826 a_89033_n35156# a_89163_n36382# a_90969_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4827 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4828 a_57417_n18700# a_50751_n19729# a_56895_n19597# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4829 VSS VSS VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X4830 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4831 a_83141_n1530# a_71281_n10073# a_82573_n1530# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4832 a_35502_25545# a_35502_25545# VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X4833 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4834 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4835 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4836 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4837 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4838 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4839 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4840 a_60845_n4447# a_50751_n19729# a_60285_n3550# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4841 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4842 a_100235_n1530# a_71281_n8397# a_99667_n1530# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4843 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4844 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4845 a_54197_5639# a_47819_11614# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4846 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4847 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4848 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4849 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4850 VDD a_30152_10448# a_30682_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4851 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4852 a_89033_n36322# a_89163_n36382# a_90969_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4853 a_78344_10448# a_65658_4421# a_77776_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4854 a_53699_11614# a_53829_10388# a_55635_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4855 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4856 a_96849_13546# a_83325_4421# a_84017_n17715# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4857 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4858 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4859 a_88271_n7865# a_71281_n10073# a_87433_n7865# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4860 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4861 a_101641_n17715# a_71281_n8397# a_43010_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4862 a_87433_n14095# a_71281_n10073# a_86903_n14095# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4863 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4864 a_101641_n15000# a_71281_n8397# a_100803_n15000# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4865 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4866 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4867 a_111631_n21335# a_71281_n8397# a_111063_n21335# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4868 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4869 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4870 VDD a_30152_10448# a_30682_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4871 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4872 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4873 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4874 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4875 a_96849_11614# a_83325_4421# a_84017_n17715# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4876 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4877 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4878 VDD a_71281_n8397# a_112199_n1530# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4879 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4880 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4881 a_33249_34067# a_35502_24538# a_52635_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4882 a_48313_n17801# a_31953_n19727# a_47753_n16904# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4883 a_112559_n29181# a_112559_n29181# a_114485_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4884 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4885 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4886 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4887 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4888 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4889 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4890 a_58851_n17803# a_50751_n19729# a_58329_n18700# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4891 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4892 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4893 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4894 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4895 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4896 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4897 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4898 a_101641_n3340# a_71281_n8397# a_100803_n2435# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4899 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4900 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4901 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4902 a_36008_n27257# a_30152_n36322# a_37934_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4903 a_107339_n17715# a_71281_n8397# a_60677_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4904 a_47991_5507# a_50751_n19729# a_57417_n1756# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4905 a_37934_7563# a_30152_11614# a_30324_4421# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4906 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4907 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4908 a_107339_n15000# a_71281_n8397# a_106501_n15000# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4909 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4910 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4911 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4912 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4913 a_65658_4421# a_65486_11614# a_71864_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4914 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4915 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4916 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4917 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4918 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4919 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4920 a_71366_11614# a_71496_10388# a_73302_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4921 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4922 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4923 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4924 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4925 a_38097_n5342# a_100992_n29313# a_101392_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4926 a_101641_n20430# a_71281_n8397# a_100803_n20430# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4927 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4928 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4929 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4930 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4931 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4932 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4933 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4934 a_43817_n28415# a_41891_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4935 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4936 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4937 VDD a_31699_20742# a_31699_20742# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4938 a_106809_n6055# a_71281_n8397# a_106501_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4939 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4940 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4941 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4942 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4943 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4944 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4945 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4946 a_49795_n28415# a_47991_n29313# a_38097_n16007# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4947 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4948 a_100820_n35156# a_100820_n35156# a_102756_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4949 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4950 a_41891_4481# a_30324_4421# a_43848_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4951 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4952 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4953 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4954 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4955 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4956 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4957 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4958 a_73268_n27257# a_65486_n36322# a_65658_n29313# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4959 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4960 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4961 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4962 a_72596_n3060# a_71266_n4019# a_50751_n19729# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X4963 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4964 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4965 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4966 a_105365_n6960# a_71281_n8397# a_104527_n6960# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4967 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4968 a_60285_n6241# a_50751_n19729# a_59763_n6241# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4969 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4970 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4971 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4972 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4973 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4974 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4975 a_107339_n20430# a_71281_n8397# a_106501_n20430# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4976 a_95943_n15000# a_71281_n10073# a_95105_n14095# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4977 a_105933_n1530# a_71281_n8397# a_105365_n1530# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4978 a_34347_n19595# a_31953_n19727# a_33787_n19595# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4979 VDD a_100820_n35156# a_101350_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4980 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4981 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4982 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4983 a_41891_4481# a_30324_4421# a_43848_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4984 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4985 a_107230_12380# a_106830_10388# a_86903_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4986 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4987 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4988 a_47991_n29313# a_47819_n36322# a_54197_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4989 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4990 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4991 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4992 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4993 a_75585_n10973# I1N VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X4994 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X4995 a_82573_n19525# a_71281_n10073# a_81735_n19525# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4996 a_111063_n4245# a_71281_n8397# a_110225_n4245# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4997 a_52585_n8035# a_50751_n19729# a_52063_n8035# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4998 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4999 a_65677_n7138# a_50751_n19729# a_66551_n5344# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5000 a_63683_n12421# a_50751_n19729# a_63161_n13318# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5001 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5002 a_54579_n8932# a_50751_n19729# a_54019_n8035# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5003 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5004 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5005 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5006 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5007 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5008 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5009 a_94537_n14095# a_71281_n10073# a_93969_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5010 a_30324_n29313# a_30152_n36322# a_36530_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5011 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5012 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5013 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5014 a_35781_n13316# a_31953_n19727# a_35221_n12419# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5015 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5016 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5017 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5018 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5019 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5020 a_36562_n34390# a_36162_n36382# a_36032_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5021 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5022 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5023 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5024 a_55601_n29181# a_47819_n36322# a_39179_n19595# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5025 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5026 a_101641_n18620# a_71281_n8397# a_100803_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5027 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5028 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5029 a_90245_n6055# a_71281_n10073# a_89715_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5030 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5031 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5032 a_47753_n17801# a_31953_n19727# a_47231_n18698# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5033 a_66058_n28415# a_45445_n19595# a_65486_n36322# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5034 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5035 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5036 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5037 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5038 VSS a_59558_4481# a_60080_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5039 VSS a_35502_25545# a_35502_25545# VSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X5040 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5041 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5042 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5043 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5044 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5045 a_32913_n14213# a_31953_n19727# a_32353_n14213# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5046 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5047 a_83153_10448# a_83325_4421# a_85129_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5048 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5049 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5050 a_38619_n1754# a_31953_n19727# a_38097_n2651# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5051 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5052 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5053 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5054 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5055 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5056 a_100992_4421# a_100820_11614# a_107198_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5057 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5058 a_53145_n19597# a_50751_n19729# a_52585_n18700# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5059 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X5060 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5061 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5062 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5063 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5064 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5065 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5066 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5067 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5068 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5069 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5070 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5071 a_32088_13546# a_30152_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5072 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5073 a_84017_n16810# a_71281_n10073# a_83709_n13190# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5074 VDD a_31699_20742# a_35502_24538# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5075 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5076 a_107339_n18620# a_71281_n8397# a_106501_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5077 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5078 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5079 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5080 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5081 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5082 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5083 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5084 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5085 VDD a_83153_10448# a_83683_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5086 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5087 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5088 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5089 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5090 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5091 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5092 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5093 a_106830_10388# a_86903_n14095# a_114516_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5094 a_32088_11614# a_30152_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5095 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5096 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5097 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5098 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5099 a_45445_n16904# a_31953_n19727# a_44885_n16904# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5100 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5101 a_60845_n2653# a_50751_n19729# a_60285_n2653# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5102 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5103 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5104 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5105 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5106 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5107 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5108 a_33787_n8930# a_31953_n19727# a_32913_n5342# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5109 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5110 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5111 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5112 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5113 a_51711_n6241# a_50751_n19729# a_51151_n4447# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5114 a_67462_n27257# a_45445_n19595# a_44363_n16007# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5115 a_66551_n16906# a_50751_n19729# a_66029_n16906# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5116 a_31699_20742# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5117 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5118 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5119 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5120 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5121 a_32353_n17801# a_31953_n19727# a_31831_n17801# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5122 VSS a_31953_n19727# a_44885_n8930# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5123 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5124 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5125 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5126 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5127 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5128 a_51711_n14215# a_50751_n19729# a_51151_n13318# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5129 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5130 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5131 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5132 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5133 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5134 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5135 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5136 a_60285_n1756# a_50751_n19729# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5137 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5138 a_33249_35053# a_35502_24538# OUT VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5139 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5140 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5141 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5142 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5143 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5144 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5145 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5146 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5147 a_36562_12380# a_36162_10388# a_36032_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5148 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5149 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5150 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5151 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5152 a_33379_34917# IN_NEG cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
X5153 a_42442_n34390# a_36032_n35156# a_36162_n36382# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5154 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5155 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5156 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5157 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5158 a_61484_n28415# a_59558_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5159 a_110225_n6055# a_71281_n8397# a_109695_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5160 a_39179_n8033# a_31953_n19727# a_38619_n7136# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5161 a_96818_n30339# a_94892_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5162 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5163 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5164 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5165 a_100820_n35156# a_100992_n29313# a_102796_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5166 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5167 a_52585_n3550# a_50751_n19729# a_52063_n3550# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5168 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5169 a_54019_n8035# a_50751_n19729# a_53497_n8035# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5170 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5171 a_32353_n6239# a_31953_n19727# a_31831_n7136# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5172 a_54579_n4447# a_50751_n19729# a_54019_n3550# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5173 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5174 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5175 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5176 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5177 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5178 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5179 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5180 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5181 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5182 a_79151_n27257# a_77225_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5183 OUT a_33379_34917# cap_mim_2f0_m4m5_noshield c_width=9.8u c_length=9.8u
X5184 a_112199_n9675# a_71281_n8397# a_111631_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5185 a_49755_10448# a_47819_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5186 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5187 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5188 VSS VSS VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X5189 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5190 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5191 a_94537_n8770# a_71281_n10073# a_93969_n8770# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5192 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5193 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5194 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5195 a_63161_n5344# a_64243_n1756# a_66058_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5196 a_71342_7563# a_71496_10388# a_71896_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5197 a_89163_10388# a_81205_n14095# a_96849_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5198 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5199 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5200 a_51151_n16906# a_50751_n19729# a_50629_n17803# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5201 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5202 a_84017_n17715# a_83325_4421# a_95443_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5203 VDD a_30152_11614# a_37934_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5204 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5205 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5206 a_42047_n19595# a_31953_n19727# a_41487_n18698# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5207 a_83725_n27257# a_83325_n29313# a_83153_n35156# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5208 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5209 a_77747_5639# a_77225_4481# a_71496_10388# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5210 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5211 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5212 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5213 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5214 a_90245_n6960# a_71281_n10073# a_89407_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5215 a_52585_n19597# a_50751_n19729# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5216 a_107198_n28415# a_100820_n36322# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5217 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5218 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5219 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5220 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5221 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5222 VSS a_71496_10388# a_71896_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5223 a_59411_n8932# a_50751_n19729# a_58851_n8932# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5224 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5225 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5226 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5227 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X5228 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5229 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5230 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5231 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5232 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5233 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5234 a_48951_4481# a_47991_5507# a_48391_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5235 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5236 a_66551_n8035# a_50751_n19729# a_66029_n8035# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5237 a_32128_5639# a_30324_4421# a_31284_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5238 a_88271_n1530# a_71281_n10073# a_87433_n1530# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5239 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5240 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5241 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5242 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5243 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X5244 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5245 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5246 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5247 a_60080_7563# a_59558_4481# a_53829_10388# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5248 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5249 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5250 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5251 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5252 a_77225_4481# a_65658_4421# a_79182_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5253 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5254 a_100820_11614# a_100820_10448# a_102756_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5255 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5256 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5257 a_53829_10388# a_59558_4481# a_61484_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5258 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5259 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5260 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5261 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5262 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5263 a_35502_24538# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5264 a_40613_n13316# a_31953_n19727# a_40053_n13316# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5265 a_65677_n17803# a_50751_n19729# a_66551_n16009# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5266 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5267 a_35502_24538# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5268 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5269 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5270 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5271 a_100820_n35156# a_100820_n35156# a_102756_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5272 a_35502_25545# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5273 a_40053_n14213# a_31953_n19727# a_39531_n14213# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5274 a_61484_6405# a_59558_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5275 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5276 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5277 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5278 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5279 a_77225_4481# a_65658_4421# a_79182_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5280 a_39179_n18698# a_31953_n19727# a_38619_n18698# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5281 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5282 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5283 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5284 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5285 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5286 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5287 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5288 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5289 a_44363_n16007# a_65658_n29313# a_66058_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5290 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5291 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5292 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5293 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5294 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5295 a_87433_n8770# a_71281_n10073# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5296 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5297 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5298 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5299 a_60285_n18700# a_50751_n19729# a_59763_n18700# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5300 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5301 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5302 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5303 a_38619_n16007# a_31953_n19727# a_38097_n16007# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5304 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5305 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5306 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5307 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5308 a_113081_n29181# a_112559_n29181# a_112559_n29181# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5309 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X5310 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5311 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5312 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5313 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5314 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5315 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5316 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5317 VDD a_100820_n35156# a_101350_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5318 a_85089_12380# a_83153_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5319 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5320 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5321 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5322 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5323 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5324 VSS a_77225_4481# a_77747_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5325 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5326 a_47991_5507# a_47819_11614# a_54197_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5327 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5328 a_54019_n3550# a_50751_n19729# a_53497_n3550# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5329 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5330 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5331 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5332 a_95105_n19525# a_71281_n10073# a_94537_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5333 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5334 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5335 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5336 a_41660_19698# a_35502_24538# a_41100_19698# VSS nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X5337 a_90245_n20430# a_71281_n10073# a_89407_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5338 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5339 a_107339_n3340# a_71281_n8397# a_106501_n3340# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5340 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5341 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5342 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5343 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5344 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5345 a_101641_n15000# a_71281_n8397# a_100803_n14095# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5346 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5347 a_45706_23609# a_35922_19591# a_45138_23609# VDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X5348 a_48313_n13316# a_31953_n19727# a_47753_n12419# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5349 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5350 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5351 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5352 a_36562_n36322# a_36162_n36382# a_36032_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5353 a_47753_n8930# a_31953_n19727# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5354 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5355 VSS a_77225_n29181# a_77747_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5356 a_41487_n19595# a_31953_n19727# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5357 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5358 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5359 a_58851_n13318# a_50751_n19729# a_58329_n14215# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5360 a_42047_n8930# a_31953_n19727# a_41487_n8033# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5361 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5362 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5363 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5364 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5365 a_88839_n19525# a_71281_n10073# a_88271_n19525# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5366 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5367 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5368 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5369 a_106676_4481# a_100820_11614# a_108602_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5370 a_30324_4421# a_30152_11614# a_36530_7563# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5371 a_94537_n7865# a_71281_n10073# a_93969_n7865# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5372 a_89715_n17715# a_86903_n14095# a_113110_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5373 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5374 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5375 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5376 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5377 VDD a_31699_20742# a_35502_24538# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5378 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5379 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5380 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5381 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5382 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5383 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5384 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5385 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5386 VDD a_31699_20742# a_35502_25545# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5387 a_66016_n34390# a_65486_n35156# a_65486_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5388 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5389 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5390 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5391 a_71342_n27257# a_65486_n36322# a_73268_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5392 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5393 a_51711_n12421# a_50751_n19729# a_51151_n12421# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5394 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5395 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5396 a_61515_12380# a_53699_11614# a_60677_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5397 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5398 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5399 a_107339_n15000# a_71281_n8397# a_106501_n14095# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5400 a_89715_n17715# a_86903_n14095# a_113110_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5401 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5402 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5403 a_52635_34067# a_35502_24538# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5404 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X5405 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5406 a_44885_n19595# a_31953_n19727# a_44363_n19595# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5407 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5408 a_66551_n3550# a_50751_n19729# a_66029_n3550# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5409 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5410 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5411 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5412 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5413 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5414 a_83709_n9675# a_71281_n10073# a_83141_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5415 a_32128_n30339# a_30324_n29313# a_31284_n30339# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5416 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5417 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5418 a_53675_n30339# a_47819_n36322# a_55601_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5419 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5420 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5421 a_111631_n8770# a_71281_n8397# a_111063_n8770# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5422 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5423 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5424 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5425 a_48313_n7136# a_31953_n19727# a_47753_n6239# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5426 a_89009_7563# a_89163_10388# a_89563_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5427 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5428 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5429 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5430 VSS a_53829_10388# a_54229_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5431 a_30152_11614# a_30152_10448# a_32088_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5432 a_83709_n18620# a_71281_n10073# a_83141_n18620# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5433 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5434 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5435 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5436 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5437 VDD a_30152_10448# a_30682_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5438 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5439 a_52585_n2653# a_50751_n19729# a_52063_n3550# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5440 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5441 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5442 a_96849_10448# a_81205_n14095# a_84017_n17715# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5443 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5444 a_108602_7563# a_100820_11614# a_100992_4421# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5445 a_36530_7563# a_30152_11614# a_36008_7563# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5446 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5447 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5448 a_85129_n28415# a_83325_n29313# a_31831_n5342# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5449 a_54579_n2653# a_50751_n19729# a_54019_n2653# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5450 a_32353_n5342# a_31953_n19727# a_31831_n5342# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5451 a_31699_20742# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5452 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5453 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5454 a_33249_34067# a_35502_24538# a_52635_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5455 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5456 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5457 a_81735_n6960# a_71281_n10073# a_81205_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5458 a_36530_n30339# a_30152_n36322# a_36008_n30339# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5459 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5460 VSS a_89163_10388# a_89563_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5461 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5462 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5463 a_75602_n4019# a_71266_n4019# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X5464 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5465 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5466 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5467 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5468 a_98829_n6960# a_71281_n8397# a_98299_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5469 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5470 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5471 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5472 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5473 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5474 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5475 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5476 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5477 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5478 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5479 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5480 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5481 a_47819_11614# a_47991_5507# a_49795_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5482 a_89531_n28415# a_83153_n36322# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5483 a_39179_n8930# a_100820_n36322# a_107198_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5484 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5485 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5486 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5487 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5488 a_93131_n18620# a_71281_n10073# a_92601_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5489 a_87433_n7865# a_71281_n10073# a_86903_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5490 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5491 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5492 a_88271_n18620# a_71281_n10073# a_87433_n18620# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5493 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5494 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5495 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5496 a_63683_n18700# a_50751_n19729# a_63161_n19597# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5497 a_42442_n36322# a_36032_n35156# a_36162_n36382# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5498 a_73302_n34390# a_71496_n36382# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5499 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5500 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5501 a_49795_6405# a_47991_5507# a_48951_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5502 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5503 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5504 a_38097_n16007# a_39179_n19595# a_48391_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5505 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5506 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5507 a_41100_19698# a_35502_24538# a_40578_19075# VSS nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X5508 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5509 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5510 a_44885_n4445# a_31953_n19727# a_44363_n4445# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5511 a_100235_n13190# a_71281_n8397# a_99667_n13190# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5512 a_95105_n9675# a_71281_n10073# a_94537_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5513 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5514 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5515 VSS VSS VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X5516 a_57417_n8035# a_50751_n19729# a_56895_n8932# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5517 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5518 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5519 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5520 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5521 a_37934_n29181# a_30152_n36322# a_30324_n30399# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5522 a_47753_n13316# a_31953_n19727# a_47231_n14213# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5523 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5524 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5525 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5526 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5527 a_107339_n3340# a_71281_n8397# a_106501_n2435# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5528 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5529 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5530 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5531 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5532 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5533 a_48391_4481# a_47991_4421# a_47819_10448# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5534 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5535 a_42047_n4445# a_31953_n19727# a_41487_n3548# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5536 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5537 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5538 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5539 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5540 a_98829_n13190# a_71281_n8397# a_98299_n16810# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5541 a_54019_n16906# a_50751_n19729# a_53497_n16906# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5542 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5543 a_93131_n6960# a_71281_n10073# a_92601_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5544 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5545 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5546 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5547 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5548 VDD a_100820_10448# a_101350_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5549 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5550 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5551 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5552 a_67111_n15112# a_50751_n19729# a_66551_n15112# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5553 a_36162_10388# a_36032_11614# a_43848_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5554 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5555 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5556 a_105365_n13190# a_71281_n8397# a_104527_n13190# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5557 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5558 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5559 a_65117_n19597# a_50751_n19729# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5560 a_35502_25545# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5561 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5562 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5563 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5564 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5565 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5566 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5567 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5568 a_59411_n19597# a_50751_n19729# a_58851_n19597# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5569 VDD a_100820_10448# a_101350_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5570 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5571 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5572 a_33249_35053# a_35502_24538# OUT VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5573 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5574 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5575 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5576 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5577 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5578 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5579 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5580 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5581 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5582 a_35502_24538# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5583 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5584 a_75585_n8397# I1N VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X5585 a_45445_n12419# a_31953_n19727# a_44885_n12419# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5586 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5587 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5588 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5589 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5590 VSS a_94892_n29181# a_95414_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5591 a_43817_n27257# a_41891_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5592 a_112199_n3340# a_71281_n8397# a_111631_n3340# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5593 a_90935_6405# a_83153_11614# a_51711_n12421# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5594 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5595 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5596 a_39179_n1754# a_31953_n19727# a_38619_n1754# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5597 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5598 a_49795_n27257# a_39179_n19595# a_38097_n16007# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5599 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5600 a_32353_n13316# a_31953_n19727# a_31831_n13316# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5601 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5602 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5603 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5604 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5605 a_54019_n2653# a_50751_n19729# a_53497_n3550# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5606 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5607 a_104527_n6960# a_71281_n8397# a_103997_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5608 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5609 a_89033_13546# a_106830_10388# a_108636_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5610 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5611 a_112199_n15000# a_71281_n8397# a_111631_n15000# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5612 a_82573_n8770# a_71281_n10073# a_81735_n8770# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5613 a_111631_n7865# a_71281_n8397# a_111063_n7865# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5614 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5615 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5616 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5617 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5618 a_66058_6405# a_65658_4421# a_65486_10448# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5619 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5620 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5621 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5622 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5623 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5624 a_83683_n34390# a_83153_n35156# a_83153_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5625 a_77225_n29181# a_77225_n29181# a_79151_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5626 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5627 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5628 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5629 a_99667_n8770# a_71281_n8397# a_98829_n8770# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5630 a_89009_n27257# a_83153_n36322# a_90935_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5631 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5632 a_38619_n8930# a_31953_n19727# a_38097_n8930# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5633 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5634 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5635 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5636 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5637 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5638 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5639 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5640 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5641 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5642 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5643 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5644 a_86903_n14095# a_106830_10388# a_108636_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5645 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5646 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5647 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5648 a_58851_n12421# a_50751_n19729# a_57977_n16009# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5649 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5650 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5651 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5652 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5653 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5654 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5655 a_100803_n9675# a_71281_n8397# a_100235_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5656 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5657 a_60845_n17803# a_50751_n19729# a_60285_n17803# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5658 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5659 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5660 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5661 a_57417_n14215# a_50751_n19729# a_56895_n15112# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5662 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5663 a_47819_11614# a_47819_10448# a_49755_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5664 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5665 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5666 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5667 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5668 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5669 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5670 a_32088_10448# a_30152_10448# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5671 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5672 a_37934_4481# a_30152_11614# a_30324_4421# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5673 a_93131_n17715# a_71281_n10073# a_92601_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5674 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5675 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5676 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5677 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5678 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5679 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5680 a_57417_n3550# a_50751_n19729# a_56895_n4447# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5681 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5682 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5683 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5684 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5685 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5686 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5687 a_112199_n20430# a_71281_n8397# a_111631_n20430# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5688 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5689 a_93969_n18620# a_71281_n10073# a_93131_n18620# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5690 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5691 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5692 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5693 a_66551_n2653# a_50751_n19729# a_66029_n3550# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5694 a_41891_4481# a_41891_4481# a_43817_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5695 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5696 a_54579_n17803# a_50751_n19729# a_54019_n17803# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5697 a_66058_n27257# a_65658_n29313# a_65486_n35156# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5698 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5699 a_83709_n21335# a_71281_n10073# a_83141_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5700 a_64243_n18700# a_50751_n19729# a_63683_n17803# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5701 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5702 a_33787_n8033# a_31953_n19727# a_33265_n8033# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5703 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5704 a_89407_n19525# a_71281_n10073# a_88839_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5705 a_46879_n3548# a_31953_n19727# a_47753_n5342# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5706 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5707 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5708 VSS a_59558_n29181# a_60080_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5709 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5710 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5711 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X5712 a_100803_n19525# a_71281_n8397# a_100235_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5713 a_45445_n8033# a_31953_n19727# a_44885_n8033# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5714 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5715 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5716 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5717 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5718 a_31699_20742# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5719 a_64243_n8035# a_50751_n19729# a_63683_n8035# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5720 a_75602_n4978# a_71266_n4019# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X5721 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5722 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5723 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5724 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5725 a_100820_10448# a_100992_4421# a_102796_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5726 a_31284_4481# a_30324_5507# a_30724_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5727 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5728 a_66016_n36322# a_65486_n35156# a_65486_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5729 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5730 a_40613_n7136# a_31953_n19727# a_40053_n7136# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5731 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5732 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5733 a_57977_n18700# a_50751_n19729# a_57417_n17803# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5734 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5735 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5736 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5737 a_65486_11614# a_65486_10448# a_67422_12380# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5738 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5739 a_83141_n15000# a_71281_n10073# a_82573_n15000# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5740 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5741 VSS VSS VSS VSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X5742 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5743 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5744 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5745 a_54197_6405# a_47819_11614# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5746 a_59558_4481# a_47991_4421# a_61515_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5747 a_93131_n21335# a_71281_n10073# a_92601_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5748 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5749 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5750 a_43817_5639# a_41891_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5751 a_88271_n21335# a_71281_n10073# a_87433_n21335# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5752 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5753 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5754 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5755 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5756 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5757 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5758 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5759 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5760 a_81735_n17715# a_71281_n10073# a_81205_n16810# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5761 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5762 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5763 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5764 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5765 a_59558_4481# a_47991_4421# a_61515_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5766 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5767 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5768 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5769 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5770 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5771 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5772 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5773 a_81735_n15000# a_71281_n10073# a_81205_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5774 a_93969_n6960# a_71281_n10073# a_93131_n6960# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5775 a_33379_34917# a_36162_10388# a_37968_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5776 a_112199_n2435# a_71281_n8397# a_111631_n2435# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5777 a_42047_n15110# a_31953_n19727# a_41487_n15110# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5778 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5779 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5780 a_41487_n6239# a_31953_n19727# a_40965_n6239# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5781 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5782 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5783 a_101392_5639# a_57977_n12421# a_100820_11614# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5784 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5785 a_94537_n1530# a_71281_n10073# a_93969_n1530# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5786 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5787 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5788 a_112199_n15905# a_71281_n8397# a_111631_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5789 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5790 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5791 a_30724_5639# a_30324_5507# a_30152_11614# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5792 a_82573_n7865# a_71281_n10073# a_81735_n7865# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5793 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5794 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5795 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5796 a_71342_4481# a_71496_10388# a_71896_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5797 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5798 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5799 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5800 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5801 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5802 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5803 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5804 a_36032_11614# a_36162_10388# a_37968_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5805 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5806 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5807 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5808 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5809 a_30324_n30399# a_31953_n19727# a_32353_n19595# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5810 a_99667_n7865# a_71281_n8397# a_98829_n7865# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5811 a_42047_n2651# a_31953_n19727# a_41487_n2651# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5812 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5813 VSS a_59558_4481# a_60080_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5814 a_83141_n20430# a_71281_n10073# a_82573_n20430# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5815 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5816 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5817 a_61484_n27257# a_59558_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5818 a_32913_n6239# a_31953_n19727# a_32353_n4445# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5819 a_83153_11614# a_51711_n12421# a_85129_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5820 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5821 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5822 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5823 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5824 a_100820_n36322# a_39179_n8930# a_102796_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5825 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5826 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5827 VSS I1N a_72603_n9297# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X5828 a_83709_n3340# a_71281_n10073# a_83141_n3340# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5829 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5830 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5831 a_73302_n36322# a_71496_n36382# a_71342_n27257# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5832 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5833 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5834 a_71864_n29181# a_65486_n36322# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5835 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5836 a_52635_34067# a_35502_24538# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5837 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5838 a_81735_n20430# a_71281_n10073# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5839 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5840 a_88839_n9675# a_71281_n10073# a_88271_n9675# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5841 a_31284_n30339# a_30324_n29313# a_30724_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5842 a_87433_n18620# a_71281_n10073# a_86903_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5843 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5844 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5845 a_100820_n36322# a_100820_n35156# a_102756_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5846 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5847 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5848 a_89407_n4245# a_71281_n10073# a_88839_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5849 a_39179_n16904# a_31953_n19727# a_38619_n15110# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5850 a_71496_10388# a_71366_11614# a_79182_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5851 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5852 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5853 a_55601_n30339# a_47819_n36322# a_47991_n29313# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5854 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5855 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5856 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5857 a_33787_n3548# a_31953_n19727# a_33265_n3548# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5858 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5859 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5860 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5861 a_33787_n12419# a_31953_n19727# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5862 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5863 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5864 a_45445_n3548# a_31953_n19727# a_44885_n3548# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5865 a_107198_n27257# a_100820_n36322# a_106676_n27257# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5866 a_51711_n12421# a_83153_11614# a_89531_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5867 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5868 a_48349_n34390# a_47819_n35156# a_47819_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5869 a_100820_n36322# a_100820_n35156# a_102756_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5870 a_105933_n13190# a_71281_n8397# a_105365_n13190# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5871 a_46879_n17801# a_31953_n19727# a_46319_n17801# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5872 VSS VSS VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X5873 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5874 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5875 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5876 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5877 VDD a_100820_n35156# a_101350_n35156# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5878 a_64243_n3550# a_50751_n19729# a_63683_n3550# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5879 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5880 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5881 a_51711_n18700# a_50751_n19729# a_51151_n18700# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5882 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5883 VSS a_35502_25545# a_35922_19591# VSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X5884 a_87433_n1530# a_71281_n10073# a_86903_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5885 a_31699_20742# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5886 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5887 a_35781_n4445# a_31953_n19727# a_35221_n4445# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5888 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5889 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5890 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5891 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5892 a_53145_n14215# a_50751_n19729# a_52585_n14215# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5893 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5894 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5895 a_65486_n35156# a_65658_n29313# a_67462_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5896 a_71281_n8397# a_71281_n8397# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5897 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5898 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5899 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5900 VDD a_100820_n35156# a_101350_n33224# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5901 a_104527_n13190# a_71281_n8397# a_103997_n16810# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5902 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5903 a_95105_n3340# a_71281_n10073# a_94537_n3340# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5904 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5905 a_31699_17542# I1U VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=6u
X5906 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5907 a_83141_n15905# a_71281_n10073# a_82573_n15905# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5908 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5909 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5910 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5911 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5912 a_83141_n9675# a_71281_n10073# a_82573_n9675# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5913 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5914 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5915 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X5916 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5917 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5918 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5919 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5920 a_36562_n35156# a_36162_n36382# a_36032_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5921 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5922 VSS a_89163_n36382# a_89563_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5923 a_41487_n16007# a_31953_n19727# a_40613_n17801# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5924 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5925 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5926 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5927 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5928 VSS a_35502_25545# a_33249_34067# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5929 a_100235_n9675# a_71281_n8397# a_99667_n9675# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5930 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5931 VDD a_47819_10448# a_48349_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5932 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5933 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5934 a_89531_5639# a_83153_11614# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5935 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5936 a_93969_n21335# a_71281_n10073# a_93131_n21335# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5937 a_47753_n8033# a_31953_n19727# a_47231_n8033# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5938 a_57417_n2653# a_50751_n19729# a_56895_n2653# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5939 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5940 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5941 a_81735_n15905# a_71281_n10073# a_81205_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5942 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5943 a_81735_n6055# a_71281_n10073# a_81205_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5944 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5945 a_99667_n19525# a_71281_n8397# a_98829_n19525# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5946 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5947 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5948 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5949 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5950 a_36562_n33224# a_36162_n36382# a_33379_34007# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5951 a_60845_n8932# a_50751_n19729# a_60285_n8932# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5952 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5953 a_83683_n36322# a_83153_n35156# a_83153_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5954 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5955 VDD a_31699_20742# a_35502_25545# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5956 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5957 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5958 VSS VSS VSS VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X5959 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5960 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5961 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5962 a_111063_n19525# a_71281_n8397# a_110225_n19525# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5963 a_98829_n6055# a_71281_n8397# a_98299_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5964 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5965 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5966 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5967 VDD a_47819_10448# a_48349_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5968 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5969 VSS a_35502_25545# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5970 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5971 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5972 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5973 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5974 a_112507_n6055# a_71281_n8397# a_112199_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5975 a_89715_n17715# a_100992_4421# a_113110_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5976 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5977 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5978 a_44885_n16007# a_31953_n19727# a_44363_n16007# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5979 a_95943_n18620# a_71281_n10073# a_95105_n18620# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5980 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5981 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5982 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5983 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5984 a_84547_n6055# a_71281_n10073# a_84017_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5985 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5986 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5987 a_95443_13546# a_81205_n14095# a_89163_10388# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5988 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5989 a_35221_n16904# a_31953_n19727# a_34699_n16904# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5990 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5991 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5992 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5993 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5994 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5995 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5996 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5997 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5998 a_111063_n6960# a_71281_n8397# a_110225_n6960# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5999 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6000 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6001 a_54229_n34390# a_53829_n36382# a_53699_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6002 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6003 a_83709_n2435# a_71281_n10073# a_83141_n2435# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6004 a_94537_n18620# a_71281_n10073# a_93969_n18620# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6005 a_95443_11614# a_81205_n14095# a_89163_10388# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6006 a_111631_n1530# a_71281_n8397# a_111063_n1530# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6007 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6008 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6009 VDD a_65486_10448# a_66016_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6010 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6011 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6012 a_48951_4481# a_47991_4421# a_48391_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6013 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6014 a_89009_4481# a_89163_10388# a_89563_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6015 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X6016 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6017 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6018 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6019 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6020 a_60080_4481# a_59558_4481# a_59558_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6021 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6022 a_40613_n19595# a_31953_n19727# a_40053_n18698# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6023 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6024 a_87433_n17715# a_71281_n10073# a_86903_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6025 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6026 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6027 a_93131_n6055# a_71281_n10073# a_92601_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6028 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6029 VDD a_71281_n8397# a_112199_n13190# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6030 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6031 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6032 VDD a_65486_10448# a_66016_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6033 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6034 a_40053_n19595# a_31953_n19727# a_39179_n16007# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6035 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6036 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6037 a_101350_13546# a_100820_10448# a_100820_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6038 a_42047_n15110# a_31953_n19727# a_41487_n14213# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6039 a_41487_n5342# a_31953_n19727# a_40613_n7136# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6040 a_35221_n4445# a_31953_n19727# a_34699_n6239# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6041 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6042 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6043 a_100803_n3340# a_71281_n8397# a_100235_n3340# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6044 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6045 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6046 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6047 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6048 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6049 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6050 a_42442_n35156# a_30324_n29313# a_41891_n29181# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6051 a_57977_n8035# a_50751_n19729# a_57417_n8035# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6052 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6053 a_96011_n36322# a_89033_n35156# a_95443_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6054 VSS VSS VSS VSS nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X6055 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6056 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6057 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6058 a_95943_n6055# a_71281_n10073# a_95413_n5150# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6059 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6060 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6061 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6062 a_51151_n7138# a_50751_n19729# a_50629_n7138# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6063 VSS I1N a_72603_n10973# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X6064 a_101350_11614# a_100820_10448# a_100820_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6065 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6066 a_105933_n9675# a_71281_n8397# a_105365_n9675# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6067 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6068 a_53145_n7138# a_50751_n19729# a_52585_n7138# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6069 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X6070 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6071 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6072 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6073 a_42442_n33224# a_30324_n29313# a_41891_n29181# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6074 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6075 VDD a_100820_n36322# a_108602_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6076 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6077 a_106501_n4245# a_71281_n8397# a_105933_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6078 VSS a_35502_25545# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X6079 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6080 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6081 a_52635_49681# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6082 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6083 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6084 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6085 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6086 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6087 a_95105_n2435# a_71281_n10073# a_94537_n2435# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6088 VSS a_77225_4481# a_77747_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6089 OUT a_33379_34917# cap_mim_2f0_m4m5_noshield c_width=9.8u c_length=9.8u
X6090 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6091 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6092 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6093 a_85129_n27257# a_32913_n8930# a_31831_n5342# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6094 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6095 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6096 a_63161_n5344# a_65658_4421# a_66058_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6097 a_104527_n6055# a_71281_n8397# a_103997_n9675# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6098 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6099 a_112199_n14095# a_71281_n8397# a_111631_n14095# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6100 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6101 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6102 VDD a_30152_11614# a_37934_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6103 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6104 a_47753_n3548# a_31953_n19727# a_47231_n3548# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6105 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6106 a_87433_n21335# a_71281_n10073# a_86903_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6107 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6108 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X6109 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6110 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6111 a_77747_6405# a_77225_4481# a_77225_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6112 VDD a_31699_20742# a_31699_20742# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6113 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X6114 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6115 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6116 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6117 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6118 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6119 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6120 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6121 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6122 a_44363_n16007# a_45445_n19595# a_66058_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6123 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6124 a_58851_n18700# a_50751_n19729# a_58329_n18700# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6125 a_39179_n14213# a_31953_n19727# a_38619_n14213# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6126 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6127 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6128 a_60845_n13318# a_50751_n19729# a_60285_n13318# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6129 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6130 a_89531_n27257# a_83153_n36322# a_89009_n27257# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6131 a_102796_n29181# a_39179_n8930# a_38097_n5342# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6132 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6133 a_33787_n2651# a_31953_n19727# a_33265_n3548# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6134 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6135 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6136 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6137 VDD a_100820_10448# a_101350_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6138 a_61484_7563# a_59558_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6139 a_60109_12380# a_47991_4421# a_59558_4481# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6140 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6141 a_35781_n17801# a_31953_n19727# a_35221_n17801# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6142 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6143 a_60285_n14215# a_50751_n19729# a_59763_n14215# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6144 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6145 OUT a_35502_24538# a_33249_35053# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6146 a_113081_n30339# a_112559_n29181# a_106830_n36382# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6147 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6148 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6149 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6150 a_106676_7563# a_100820_11614# a_108602_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6151 a_45445_n3548# a_31953_n19727# a_44885_n2651# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6152 a_30324_4421# a_30152_11614# a_36530_4481# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6153 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6154 a_38097_n16007# a_47991_n29313# a_48391_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6155 a_32128_6405# a_30324_5507# a_31284_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6156 VDD VDD VDD VDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X6157 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6158 a_64243_n3550# a_50751_n19729# a_63683_n2653# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6159 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6160 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6161 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6162 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6163 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6164 a_95943_n17715# a_71281_n10073# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6165 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6166 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6167 a_114516_13546# a_100992_4421# a_89715_n17715# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6168 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6169 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6170 a_110225_n8770# a_71281_n8397# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6171 a_84547_n6960# a_71281_n10073# a_83709_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6172 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6173 a_54579_n13318# a_50751_n19729# a_54019_n13318# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6174 a_40613_n2651# a_31953_n19727# a_40053_n1754# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6175 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6176 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6177 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6178 a_47819_n35156# a_47819_n35156# a_49755_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6179 a_39179_n8930# a_31953_n19727# a_38619_n8930# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6180 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6181 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6182 a_64243_n14215# a_50751_n19729# a_63683_n13318# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6183 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6184 a_110225_n19525# a_71281_n8397# a_109695_n19525# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6185 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6186 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6187 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6188 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6189 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6190 a_114516_11614# a_100992_4421# a_89715_n17715# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6191 VSS a_41891_n29181# a_42413_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6192 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X6193 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6194 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6195 VSS a_77225_n29181# a_77747_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6196 VDD a_71281_n10073# a_71281_n10073# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6197 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6198 a_106676_7563# a_106830_10388# a_107230_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6199 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6200 a_82573_n1530# a_71281_n10073# a_81735_n1530# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6201 OUT a_106830_10388# a_108636_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6202 VDD a_47819_n35156# a_48349_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6203 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6204 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6205 a_46319_n12419# a_31953_n19727# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6206 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6207 a_106501_n13190# a_71281_n8397# a_105933_n13190# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6208 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6209 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6210 a_99667_n1530# a_71281_n8397# a_98829_n1530# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6211 a_108602_4481# a_100820_11614# a_100992_4421# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6212 a_57977_n14215# a_50751_n19729# a_57417_n13318# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6213 a_38619_n8033# a_31953_n19727# a_38097_n8930# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6214 a_36530_4481# a_30152_11614# a_36008_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6215 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6216 a_48349_n36322# a_47819_n35156# a_47819_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6217 a_101641_n6055# a_71281_n8397# a_96011_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6218 a_30682_13546# a_30152_10448# a_30152_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6219 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6220 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6221 a_77776_12380# a_65658_4421# a_77225_4481# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6222 a_55635_12380# a_53829_10388# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6223 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6224 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6225 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6226 VSS a_106830_10388# a_107230_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6227 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6228 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6229 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6230 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6231 VSS VSS VSS VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X6232 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6233 a_57977_n3550# a_50751_n19729# a_57417_n3550# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6234 a_90245_n6960# a_71281_n10073# a_89407_n6960# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6235 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6236 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6237 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6238 a_112559_4481# a_112559_4481# a_114485_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6239 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6240 VSS a_41891_4481# a_42413_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6241 a_33249_34067# a_35502_24538# a_52635_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6242 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6243 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6244 a_47991_5507# a_47819_11614# a_54197_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6245 a_71896_n34390# a_71496_n36382# a_71366_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6246 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6247 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6248 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6249 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6250 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6251 a_83141_n14095# a_71281_n10073# a_82573_n14095# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6252 a_90935_n29181# a_83153_n36322# a_32913_n8930# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6253 a_100803_n2435# a_71281_n8397# a_100235_n2435# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6254 a_30682_11614# a_30152_10448# a_30152_11614# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6255 VDD a_71281_n10073# a_95105_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6256 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6257 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6258 a_33249_34067# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6259 a_88839_n3340# a_71281_n10073# a_88271_n3340# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6260 a_33379_34917# IN_NEG cap_mim_2f0_m4m5_noshield c_width=100u c_length=100u
X6261 a_95943_n6960# a_71281_n10073# a_95105_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6262 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6263 VSS a_35502_25545# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X6264 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6265 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6266 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6267 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6268 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6269 a_84547_n17715# a_71281_n10073# a_84017_n16810# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6270 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6271 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6272 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6273 a_96849_n34390# a_83325_n29313# a_96011_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6274 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6275 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6276 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6277 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6278 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6279 a_84547_n15000# a_71281_n10073# a_83709_n15000# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6280 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6281 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6282 a_89009_n30339# a_89163_n36382# a_89563_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6283 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6284 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6285 a_71366_13546# a_89163_10388# a_90969_13546# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6286 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6287 a_81735_n14095# a_71281_n10073# a_81205_n14095# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6288 a_71281_n10073# a_71281_n10073# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6289 a_56895_n16009# a_57977_n12421# a_101392_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6290 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6291 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6292 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6293 VDD VDD VDD VDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X6294 a_94537_n21335# a_71281_n10073# a_93969_n21335# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6295 a_47753_n18698# a_31953_n19727# a_47231_n18698# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6296 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6297 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6298 VDD a_30152_n35156# a_30682_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6299 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6300 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6301 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6302 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6303 a_113081_5639# a_112559_4481# a_106830_10388# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6304 a_52585_n8932# a_50751_n19729# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6305 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6306 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6307 a_65486_10448# a_65658_4421# a_67462_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6308 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6309 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6310 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6311 a_111631_n19525# a_71281_n8397# a_111063_n19525# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6312 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6313 a_54579_n8932# a_50751_n19729# a_54019_n8932# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6314 a_42413_5639# a_41891_4481# a_36162_10388# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6315 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6316 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6317 a_81205_n14095# a_89163_10388# a_90969_11614# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6318 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6319 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6320 a_60285_n8035# a_50751_n19729# a_59763_n8035# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6321 a_66016_n35156# a_65486_n35156# a_65486_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6322 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6323 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6324 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6325 a_79151_5639# a_77225_4481# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6326 VSS VSS VSS VSS nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X6327 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6328 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6329 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6330 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6331 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6332 a_53699_n35156# a_53829_n36382# a_55635_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6333 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6334 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6335 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6336 a_100992_n29313# a_100820_n36322# a_107198_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6337 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6338 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6339 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6340 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6341 a_54197_n29181# a_47819_n36322# VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6342 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6343 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6344 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6345 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6346 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6347 a_66016_n33224# a_65486_n35156# a_65486_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6348 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6349 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6350 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6351 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6352 a_83141_n3340# a_71281_n10073# a_82573_n3340# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6353 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6354 a_67111_n7138# a_50751_n19729# a_66551_n7138# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6355 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6356 a_63683_n14215# a_50751_n19729# a_63161_n15112# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6357 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6358 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6359 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6360 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6361 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6362 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6363 a_84547_n20430# a_71281_n10073# a_83709_n20430# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6364 a_33249_35053# a_33379_34917# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6365 a_53829_10388# a_53699_11614# a_61515_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6366 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6367 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6368 a_100235_n3340# a_71281_n8397# a_99667_n3340# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6369 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6370 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6371 a_35502_25545# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6372 a_37934_n30339# a_30152_n36322# a_30324_n29313# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6373 a_54229_n36322# a_53829_n36382# a_53699_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6374 a_51151_n6241# a_50751_n19729# a_50629_n7138# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6375 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6376 a_49795_7563# a_47991_4421# a_48951_4481# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6377 a_110225_n7865# a_71281_n8397# a_109695_n7865# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6378 a_108602_n29181# a_100820_n36322# a_39179_n8930# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6379 a_88271_n9675# a_71281_n10073# a_87433_n9675# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6380 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6381 a_101641_n18620# a_71281_n8397# a_100803_n18620# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6382 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6383 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6384 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6385 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6386 a_46879_n13316# a_31953_n19727# a_46319_n13316# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6387 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6388 a_32353_n18698# a_31953_n19727# a_31831_n19595# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6389 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6390 VSS a_59558_n29181# a_60080_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6391 a_36032_13546# a_36162_10388# a_37968_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6392 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6393 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6394 a_32913_n16007# a_31953_n19727# a_32353_n16007# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6395 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6396 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6397 a_38619_n3548# a_31953_n19727# a_38097_n4445# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6398 a_113037_n3340# a_71281_n8397# a_112199_n3340# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6399 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6400 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6401 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6402 a_66016_12380# a_65486_10448# a_65486_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6403 a_47753_n2651# a_31953_n19727# a_47231_n3548# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6404 a_47819_n35156# a_47991_n29313# a_49795_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6405 a_75602_n3060# a_71266_n4019# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X6406 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6407 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6408 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6409 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6410 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6411 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6412 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6413 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6414 a_73302_n35156# a_71496_n36382# VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6415 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6416 a_65486_n35156# a_65486_n35156# a_67422_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6417 a_101641_n6960# a_71281_n8397# a_100803_n4245# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6418 a_96011_n36322# a_89033_n35156# a_95443_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6419 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6420 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X6421 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6422 a_107339_n18620# a_71281_n8397# a_106501_n18620# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6423 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6424 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6425 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6426 a_60845_n13318# a_50751_n19729# a_60285_n12421# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6427 a_63683_n5344# a_50751_n19729# a_63161_n5344# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6428 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6429 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6430 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6431 a_83153_n36322# a_32913_n8930# a_85129_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6432 a_50751_n19729# a_50751_n19729# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6433 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6434 VDD a_47819_11614# a_55601_5639# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6435 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6436 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6437 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6438 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6439 a_57417_n19597# a_50751_n19729# a_56895_n19597# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6440 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6441 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6442 VSS a_94892_n29181# a_95414_n30339# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6443 a_73302_n33224# a_71496_n36382# a_71342_n30339# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6444 VDD a_31699_20742# a_35502_24538# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6445 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6446 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6447 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6448 a_101392_n28415# a_39179_n8930# a_100820_n36322# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6449 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6450 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6451 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6452 VSS VSS VSS VSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X6453 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6454 VDD a_65486_n35156# a_66016_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6455 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6456 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6457 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6458 a_60845_n4447# a_50751_n19729# a_60285_n4447# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6459 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6460 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6461 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6462 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6463 a_88839_n2435# a_71281_n10073# a_88271_n2435# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6464 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6465 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6466 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6467 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6468 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6469 a_54579_n13318# a_50751_n19729# a_54019_n12421# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6470 a_84547_n18620# a_71281_n10073# a_83709_n15905# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6471 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6472 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6473 IBNOUT a_50751_n19729# a_63683_n12421# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6474 a_90935_7563# a_83153_11614# a_83325_4421# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6475 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6476 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6477 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6478 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6479 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6480 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6481 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6482 a_54019_n8932# a_50751_n19729# a_51711_n8932# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6483 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6484 a_42413_n29181# a_41891_n29181# a_41891_n29181# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6485 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6486 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6487 VSS VSS VSS VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X6488 a_60285_n3550# a_50751_n19729# a_59763_n3550# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6489 a_83683_12380# a_83153_10448# a_83153_10448# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6490 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6491 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6492 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6493 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6494 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6495 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6496 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6497 a_52635_48695# a_35922_19591# a_52635_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6498 a_35221_n12419# a_31953_n19727# a_32913_n12419# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6499 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6500 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6501 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6502 a_66058_7563# a_64243_n1756# a_65486_11614# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6503 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6504 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6505 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6506 a_32088_n34390# a_30152_n35156# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6507 a_105365_n8770# a_71281_n8397# a_104527_n8770# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6508 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6509 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6510 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6511 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6512 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6513 a_48313_n17801# a_31953_n19727# a_47753_n17801# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6514 a_114485_n28415# a_112559_n29181# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6515 a_55601_5639# a_47819_11614# a_47991_5507# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6516 VDD a_31699_20742# a_33249_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6517 a_33249_34067# a_33379_34007# a_33249_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6518 a_89163_n36382# a_94892_n29181# a_96818_n29181# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6519 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6520 a_105933_n3340# a_71281_n8397# a_105365_n3340# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6521 a_57977_n12421# a_50751_n19729# a_57417_n12421# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6522 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X6523 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6524 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6525 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6526 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6527 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6528 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6529 VDD a_31699_20742# a_31699_20742# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6530 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6531 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6532 a_57977_n3550# a_50751_n19729# a_57417_n2653# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6533 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6534 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6535 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6536 VDD a_71281_n8397# a_71281_n8397# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6537 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6538 OUT a_35922_19591# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6539 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6540 a_47819_n35156# a_47819_n35156# a_49755_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6541 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6542 a_51151_n1756# a_50751_n19729# a_50629_n2653# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6543 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6544 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6545 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6546 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6547 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6548 a_83141_n2435# a_71281_n10073# a_82573_n2435# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6549 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6550 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6551 a_53145_n2653# a_50751_n19729# a_52585_n1756# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6552 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6553 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6554 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6555 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6556 a_83683_n35156# a_83153_n35156# a_83153_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6557 a_100235_n2435# a_71281_n8397# a_99667_n2435# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6558 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6559 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6560 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6561 a_71366_n35156# a_71496_n36382# a_73302_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6562 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6563 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6564 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6565 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6566 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6567 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6568 a_52635_48695# a_52635_34067# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6569 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6570 VDD a_47819_10448# a_48349_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6571 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6572 a_66551_n8932# a_50751_n19729# a_64243_n8932# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6573 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6574 VSS a_35502_25545# a_33249_34067# VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X6575 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6576 a_60080_n29181# a_59558_n29181# a_59558_n29181# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6577 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6578 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6579 a_101641_n17715# a_71281_n8397# a_101111_n17715# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6580 VDD a_47819_n35156# a_48349_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6581 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6582 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6583 a_33249_35053# a_35502_24538# OUT VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6584 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6585 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6586 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6587 a_78344_n36322# a_71366_n35156# a_77776_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6588 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6589 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6590 a_83683_n33224# a_83153_n35156# a_83153_n35156# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6591 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6592 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6593 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6594 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6595 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X6596 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6597 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6598 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6599 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6600 a_65486_n36322# a_45445_n19595# a_67462_n27257# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6601 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6602 a_67111_n17803# a_50751_n19729# a_66551_n16906# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6603 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6604 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6605 VSS a_71496_n36382# a_71896_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6606 a_113037_n3340# a_71281_n8397# a_112199_n2435# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6607 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6608 a_33249_48695# a_33379_34917# a_33249_35053# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6609 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6610 a_52635_34067# a_35922_19591# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6611 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6612 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6613 a_71896_n36322# a_71496_n36382# a_71366_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6614 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6615 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6616 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6617 VDD a_52635_34067# a_52635_49681# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6618 VSS a_50751_n19729# a_50751_n19729# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6619 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6620 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6621 a_33249_48695# a_31699_20742# VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6622 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6623 a_95443_10448# a_83325_4421# a_94892_4481# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6624 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6625 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6626 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6627 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6628 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6629 a_107339_n17715# a_71281_n8397# a_106809_n17715# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6630 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6631 a_94892_n29181# a_83325_n29313# a_96849_n34390# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6632 a_38619_n16904# a_31953_n19727# a_38097_n17801# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6633 a_31699_20742# a_31699_20742# VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6634 a_36162_10388# a_41891_4481# a_43817_6405# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6635 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6636 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6637 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6638 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6639 a_96849_n36322# a_83325_n29313# a_96011_n36322# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6640 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6641 a_54197_7563# a_47819_11614# a_53675_7563# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6642 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6643 a_71266_n4019# I1N a_75585_n10073# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X6644 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6645 a_31953_n19727# a_31953_n19727# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6646 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6647 a_59558_n29181# a_59558_n29181# a_61484_n28415# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6648 VSS a_35502_25545# a_33249_35053# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6649 a_33249_48695# a_33379_34007# a_33249_34067# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6650 a_67111_n7138# a_50751_n19729# a_66551_n6241# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6651 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6652 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6653 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6654 a_33249_35053# a_35502_25545# VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6655 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6656 a_52635_49681# a_35922_19591# OUT VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6657 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6658 VDD a_65486_10448# a_66016_10448# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6659 VDD a_30152_n35156# a_30682_n36322# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6660 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6661 VSS a_31953_n19727# a_31953_n19727# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6662 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6663 VDD VDD VDD VDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X6664 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6665 a_101111_n17715# a_71281_n8397# a_100803_n21335# VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6666 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6667 VDD a_52635_34067# a_52635_48695# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6668 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6669 a_35781_n13316# a_31953_n19727# a_35221_n13316# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6670 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6671 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
.ends

