* NGSPICE file created from clockGeneratorLayout.ext - technology: gf180mcuD

.subckt clockGeneratorLayout GND IBIAS VDD OUT
X0 a_16964_8348.t0 GND.t30 cap_mim_2f0_m4m5_noshield c_width=42u c_length=10u
X1 GND.t335 GND.t334 GND.t335 GND.t17 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X2 a_21743_6100.t13 a_21743_6748.t14 GND.t8 GND.t7 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X3 a_21743_6100.t3 a_16964_8348.t3 a_21659_3242.t7 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X4 a_21659_3242.t23 a_11345_12294.t2 VDD.t37 VDD.t10 pfet_03v3 ad=0.52p pd=2.52u as=1.3p ps=5.3u w=2u l=2u
X5 GND.t333 GND.t332 GND.t333 GND.t135 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X6 VDD.t262 VDD.t261 VDD.t262 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X7 a_11300_8092.t7 a_11300_8092.t6 a_16434_7468.t1 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X8 VDD.t260 VDD.t259 VDD.t260 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X9 a_19582_6043.t2 a_25891_6334.t4 a_28935_6098# w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X10 a_25891_n1726.t1 a_25891_n1726.t0 a_28583_n2146# w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X11 GND.t331 GND.t330 GND.t331 GND.t102 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X12 VDD.t36 a_11345_12294.t2 a_21659_3242.t15 VDD.t8 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=2u
X13 a_21743_n1960.t8 a_9120_14251.t2 a_21659_n106.t11 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X14 VDD.t258 VDD.t257 VDD.t258 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X15 VDD.t256 VDD.t255 VDD.t256 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X16 a_21743_n2608.t11 a_16964_8348.t4 a_21659_n106.t7 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X17 VDD.t254 VDD.t253 VDD.t254 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X18 a_16434_7468.t21 a_16434_7468.t20 VDD.t279 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X19 a_9120_14251.t1 a_28848_14251# GND.t0 ppolyf_u_1k r_width=1u r_length=98u
X20 a_9938_8092.t55 a_10060_n1528.t13 GND.t411 GND.t70 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X21 a_9938_8092.t54 a_10060_n1528.t14 GND.t375 GND.t204 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X22 a_21743_n2608.t10 a_16964_8348.t5 a_21659_n106.t1 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X23 GND.t329 GND.t328 GND.t329 GND.t89 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X24 a_9938_8092.t53 a_10060_n1528.t15 GND.t406 GND.t13 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X25 a_21743_6748.t5 a_21743_6100.t14 GND.t357 GND.t7 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X26 a_11618_8092.t6 a_10060_n1528.t16 GND.t416 GND.t175 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X27 VDD.t252 VDD.t251 VDD.t252 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X28 GND.t327 GND.t326 GND.t327 GND.t152 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X29 a_19718_7047# OUT.t0 a_19582_6479.t0 VDD.t271 pfet_03v3 ad=0.39p pd=2.5u as=0.39p ps=2.5u w=0.6u l=0.6u
X30 OUT.t0 a_19582_6043.t3 GND.t368 GND.t367 nfet_03v3 ad=0.366p pd=2.42u as=0.366p ps=2.42u w=0.6u l=0.6u
X31 VDD.t250 VDD.t249 VDD.t250 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X32 a_25891_6334.t1 a_21743_6748.t15 GND.t10 GND.t9 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X33 GND.t325 GND.t324 GND.t325 GND.t144 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X34 a_10778_8092.t27 a_10060_n1528.t17 GND.t354 GND.t13 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X35 a_11345_12294.t1 a_11345_12294.t0 VDD.t35 VDD.t34 pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X36 a_21743_n1960.t7 a_9120_14251.t3 a_21659_n106.t10 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X37 a_21743_6748.t4 a_21743_6100.t15 GND.t342 GND.t79 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X38 GND.t323 GND.t322 GND.t323 GND.t50 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X39 a_21743_n2608.t13 a_21743_n1960.t14 GND.t372 GND.t76 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X40 VDD.t248 VDD.t247 VDD.t248 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X41 VDD.t246 VDD.t245 VDD.t246 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X42 a_11345_12294.t0 a_10060_n1528.t18 GND.t346 GND.t345 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X43 VDD.t244 VDD.t243 VDD.t244 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X44 a_10778_8092.t26 a_10060_n1528.t19 GND.t419 GND.t175 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X45 GND.t321 GND.t320 GND.t321 GND.t204 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X46 a_21743_n1960.t9 a_21743_n2608.t14 GND.t446 GND.t76 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X47 VDD.t242 VDD.t241 VDD.t242 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X48 VDD.t240 VDD.t239 VDD.t240 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X49 VDD.t238 VDD.t237 VDD.t238 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X50 a_21659_3242.t13 a_11345_12294.t2 VDD.t33 VDD.t6 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=2u
X51 a_16964_8348.t2 a_11300_8092.t8 a_16434_8348.t1 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X52 VDD.t236 VDD.t235 VDD.t236 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X53 GND.t319 GND.t318 GND.t319 GND.t175 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X54 a_9938_8092.t52 a_10060_n1528.t20 GND.t426 GND.t172 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X55 a_25891_n1726.t2 a_21743_n2608.t15 GND.t16 GND.t15 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X56 GND.t317 GND.t316 GND.t317 GND.t50 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X57 VDD.t32 a_11345_12294.t2 a_21659_3242.t12 VDD.t4 pfet_03v3 ad=1.3p pd=5.3u as=0.52p ps=2.52u w=2u l=2u
X58 VDD.t234 VDD.t233 VDD.t234 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X59 GND.t315 GND.t314 GND.t315 GND.t172 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X60 a_9938_8092.t51 a_10060_n1528.t21 GND.t24 GND.t13 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X61 a_11618_8092.t5 a_10060_n1528.t22 GND.t6 GND.t5 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X62 a_19582_7363.t2 a_21743_n1960.t15 GND.t421 GND.t15 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X63 a_16434_8348.t11 a_16434_7468.t22 VDD.t280 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X64 a_21743_n2608.t9 a_16964_8348.t6 a_21659_n106.t5 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X65 VDD.t232 VDD.t231 VDD.t232 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X66 a_9938_8092.t50 a_10060_n1528.t23 GND.t14 GND.t13 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X67 a_19582_6043.t1 a_21743_6100.t16 GND.t343 GND.t9 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X68 VDD.t230 VDD.t229 VDD.t230 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X69 VDD.t228 VDD.t227 VDD.t228 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X70 VDD.t226 VDD.t225 VDD.t226 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X71 a_21743_6100.t12 a_21743_6748.t16 GND.t428 GND.t79 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X72 a_16964_8348.t0 GND.t29 cap_mim_2f0_m4m5_noshield c_width=42u c_length=10u
X73 GND.t313 GND.t312 GND.t313 GND.t86 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X74 GND.t311 GND.t310 GND.t311 GND.t3 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X75 a_21659_n106.t27 a_11345_12294.t3 VDD.t31 VDD.t26 pfet_03v3 ad=0.52p pd=2.52u as=1.3p ps=5.3u w=2u l=2u
X76 VDD.t224 VDD.t223 VDD.t224 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X77 GND.t309 GND.t308 GND.t309 GND.t105 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X78 VDD.t222 VDD.t221 VDD.t222 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X79 a_19582_7363.t0 a_25891_n1726.t4 a_28935_n1490# w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X80 GND.t307 GND.t306 GND.t307 GND.t58 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X81 GND.t305 GND.t304 GND.t305 GND.t99 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X82 a_16964_8348.t0 GND.t28 cap_mim_2f0_m4m5_noshield c_width=42u c_length=10u
X83 a_10460_8092.t9 IBIAS.t2 a_9938_8092.t7 GND.t276 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X84 VDD.t220 VDD.t219 VDD.t220 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X85 a_10778_8092.t25 a_10060_n1528.t24 GND.t371 GND.t5 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X86 a_9938_8092.t49 a_10060_n1528.t25 GND.t384 GND.t22 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X87 VDD.t218 VDD.t217 VDD.t218 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X88 GND.t303 GND.t302 GND.t303 GND.t163 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X89 a_10778_8092.t24 a_10060_n1528.t26 GND.t390 GND.t13 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X90 a_21743_n1960.t13 a_21743_n1960.t12 GND.t382 GND.t41 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X91 VDD.t216 VDD.t215 VDD.t216 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X92 a_11618_8092.t4 a_10060_n1528.t27 GND.t362 GND.t5 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X93 VDD.t214 VDD.t213 VDD.t214 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X94 VDD.t212 VDD.t211 VDD.t212 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X95 GND.t301 GND.t300 GND.t301 GND.t204 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X96 VDD.t210 VDD.t209 VDD.t210 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X97 VDD.t208 VDD.t207 VDD.t208 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X98 a_21743_n2608.t3 a_21743_n2608.t2 GND.t361 GND.t41 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X99 GND.t299 GND.t298 GND.t299 GND.t112 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X100 a_21743_6100.t11 a_21743_6100.t10 GND.t356 GND.t35 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X101 a_10778_8092.t23 a_10060_n1528.t28 GND.t23 GND.t22 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X102 VDD.t270 OUT.t0 a_10460_8092.t1 GND.t394 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X103 a_9938_8092.t48 a_10060_n1528.t29 GND.t369 GND.t13 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X104 a_9938_8092.t47 a_10060_n1528.t30 GND.t427 GND.t70 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X105 a_9938_8092.t46 a_10060_n1528.t31 GND.t388 GND.t11 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X106 a_28935_n1490# a_25891_n1726.t5 VDD.t267 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X107 a_10060_n1528.t12 a_10060_n1528.t11 GND.t364 GND.t5 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X108 a_16434_7468.t19 a_16434_7468.t18 VDD.t269 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X109 GND.t297 GND.t296 GND.t297 GND.t38 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X110 a_21743_6748.t3 a_9248_11691.t2 a_21659_3242.t11 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X111 a_21659_n106.t26 a_11345_12294.t3 VDD.t30 VDD.t26 pfet_03v3 ad=0.52p pd=2.52u as=1.3p ps=5.3u w=2u l=2u
X112 a_9938_8092.t45 a_10060_n1528.t32 GND.t398 GND.t22 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X113 GND.t295 GND.t294 GND.t295 GND.t112 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X114 VDD.t206 VDD.t205 VDD.t206 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X115 a_19582_6479.t1 OUT.t0 GND.t393 GND.t392 nfet_03v3 ad=0.366p pd=2.42u as=0.366p ps=2.42u w=0.6u l=0.6u
X116 VDD.t204 VDD.t203 VDD.t204 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X117 a_21743_6100.t4 a_16964_8348.t7 a_21659_3242.t6 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X118 a_9938_8092.t44 a_10060_n1528.t33 GND.t355 GND.t70 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X119 VDD.t202 VDD.t201 VDD.t202 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X120 a_11345_12294.t0 a_10060_n1528.t34 GND.t450 GND.t449 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X121 GND.t293 GND.t292 GND.t293 GND.t276 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X122 a_10778_8092.t22 a_10060_n1528.t35 GND.t381 GND.t5 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X123 a_10778_8092.t21 a_10060_n1528.t36 GND.t433 GND.t11 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X124 a_10778_8092.t20 a_10060_n1528.t37 GND.t435 GND.t22 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X125 a_21743_n1960.t6 a_9120_14251.t4 a_21659_n106.t15 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X126 VDD.t29 a_11345_12294.t4 a_21659_n106.t25 VDD.t23 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=2u
X127 VDD.t200 VDD.t199 VDD.t200 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X128 a_10060_n1528.t10 a_10060_n1528.t9 GND.t420 GND.t5 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X129 a_9938_8092.t43 a_10060_n1528.t38 GND.t452 GND.t22 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X130 a_21743_6748.t13 a_21743_6748.t12 GND.t445 GND.t35 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X131 a_28583_6754# a_25891_6334.t5 VDD.t0 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X132 GND.t291 GND.t290 GND.t291 GND.t13 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X133 GND.t289 GND.t288 GND.t289 GND.t63 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X134 a_16434_8348.t10 a_16434_7468.t23 VDD.t276 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X135 GND.t287 GND.t286 GND.t287 GND.t7 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X136 VDD.t264 a_19582_7363.t3 a_19718_7047# VDD.t263 pfet_03v3 ad=0.39p pd=2.5u as=0.39p ps=2.5u w=0.6u l=0.6u
X137 a_9938_8092.t42 a_10060_n1528.t39 GND.t431 GND.t86 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X138 a_21659_n106.t24 a_11345_12294.t3 VDD.t28 VDD.t19 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=2u
X139 a_21659_n106.t23 a_11345_12294.t3 VDD.t27 VDD.t26 pfet_03v3 ad=0.52p pd=2.52u as=1.3p ps=5.3u w=2u l=2u
X140 GND.t285 GND.t284 GND.t285 GND.t112 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X141 VDD.t198 VDD.t197 VDD.t198 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X142 VDD.t196 VDD.t195 VDD.t196 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X143 GND.t283 GND.t282 GND.t283 GND.t86 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X144 GND.t281 GND.t280 GND.t281 GND.t112 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X145 GND.t279 GND.t278 GND.t279 GND.t152 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X146 a_9938_8092.t41 a_10060_n1528.t40 GND.t444 GND.t70 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X147 a_21743_6748.t0 a_9248_11691.t3 a_21659_3242.t8 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X148 GND.t277 GND.t275 GND.t277 GND.t276 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X149 GND.t274 GND.t273 GND.t274 GND.t112 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X150 a_10778_8092.t19 a_10060_n1528.t41 GND.t21 GND.t11 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X151 GND.t272 GND.t271 GND.t272 GND.t144 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X152 VDD.t25 a_11345_12294.t3 a_21659_n106.t22 VDD.t23 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=2u
X153 a_21743_6100.t7 a_16964_8348.t8 a_21659_3242.t5 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X154 VDD.t194 VDD.t193 VDD.t194 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X155 a_10778_8092.t18 a_10060_n1528.t42 GND.t399 GND.t175 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X156 GND.t270 GND.t269 GND.t270 GND.t70 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X157 GND.t268 GND.t267 GND.t268 GND.t55 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X158 VDD.t192 VDD.t191 VDD.t192 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X159 a_9938_8092.t40 a_10060_n1528.t43 GND.t415 GND.t172 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X160 VDD.t24 a_11345_12294.t4 a_21659_n106.t21 VDD.t23 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=2u
X161 a_25891_6334.t3 a_25891_6334.t2 a_28583_6754# w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X162 a_9938_8092.t39 a_10060_n1528.t44 GND.t12 GND.t11 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X163 a_21743_6748.t1 a_9248_11691.t4 a_21659_3242.t9 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X164 VDD.t190 VDD.t189 VDD.t190 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X165 a_9938_8092.t38 a_10060_n1528.t45 GND.t397 GND.t204 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X166 GND.t19 GND.t20 GND.t0 ppolyf_u_1k r_width=1u r_length=98u
X167 VDD.t188 VDD.t187 VDD.t188 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X168 GND.t266 GND.t265 GND.t266 GND.t144 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X169 a_21743_n2608.t8 a_16964_8348.t9 a_21659_n106.t2 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X170 VDD.t186 VDD.t185 VDD.t186 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X171 GND.t264 GND.t263 GND.t264 GND.t50 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X172 a_21743_n1960.t5 a_9120_14251.t5 a_21659_n106.t14 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X173 VDD.t184 VDD.t183 VDD.t184 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X174 a_11618_8092.t3 a_10060_n1528.t46 GND.t348 GND.t175 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X175 a_9938_8092.t37 a_10060_n1528.t47 GND.t377 GND.t172 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X176 VDD.t182 VDD.t181 VDD.t182 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X177 a_16434_7468.t17 a_16434_7468.t16 VDD.t275 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X178 a_21743_n1960.t4 a_9120_14251.t6 a_21659_n106.t9 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X179 VDD.t180 VDD.t179 VDD.t180 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X180 a_10778_8092.t17 a_10060_n1528.t48 GND.t402 GND.t5 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X181 VDD.t178 VDD.t177 VDD.t178 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X182 a_11300_8092.t3 IBIAS.t3 a_10778_8092.t3 GND.t223 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X183 VDD.t176 VDD.t175 VDD.t176 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X184 a_21659_n106.t20 a_11345_12294.t3 VDD.t22 VDD.t19 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=2u
X185 a_21743_6748.t2 a_9248_11691.t5 a_21659_3242.t10 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X186 a_10778_8092.t16 a_10060_n1528.t49 GND.t359 GND.t22 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X187 GND.t262 GND.t261 GND.t262 GND.t152 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X188 VDD.t174 VDD.t173 VDD.t174 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X189 a_10778_8092.t15 a_10060_n1528.t50 GND.t387 GND.t5 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X190 a_10778_8092.t14 a_10060_n1528.t51 GND.t404 GND.t96 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X191 a_10460_8092.t8 IBIAS.t4 a_9938_8092.t5 GND.t276 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X192 a_9938_8092.t36 a_10060_n1528.t52 GND.t448 GND.t149 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X193 a_21743_6100.t5 a_16964_8348.t10 a_21659_3242.t4 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X194 VDD.t172 VDD.t171 VDD.t172 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X195 GND.t260 GND.t259 GND.t260 GND.t9 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X196 GND.t258 GND.t257 GND.t258 GND.t5 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X197 a_9938_8092.t35 a_10060_n1528.t53 GND.t396 GND.t22 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X198 GND.t256 GND.t255 GND.t256 GND.t32 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X199 VDD.t21 a_11345_12294.t5 a_21659_n106.t19 VDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0.52p ps=2.52u w=2u l=2u
X200 GND.t254 GND.t253 GND.t254 GND.t79 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X201 VDD.t170 VDD.t169 VDD.t170 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X202 GND.t252 GND.t251 GND.t252 GND.t76 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X203 GND.t250 GND.t249 GND.t250 GND.t17 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X204 a_16434_7468.t15 a_16434_7468.t14 VDD.t274 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X205 VDD.t168 VDD.t167 VDD.t168 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X206 GND.t248 GND.t247 GND.t248 GND.t135 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X207 GND.t246 GND.t245 GND.t246 GND.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X208 a_28583_n2146# a_25891_n1726.t6 VDD.t268 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X209 GND.t244 GND.t243 GND.t244 GND.t112 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X210 a_21743_n2608.t7 a_16964_8348.t11 a_21659_n106.t4 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X211 a_10778_8092.t13 a_10060_n1528.t54 GND.t409 GND.t175 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X212 a_11618_8092.t2 a_10060_n1528.t55 GND.t423 GND.t96 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X213 GND.t242 GND.t241 GND.t242 GND.t105 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X214 GND.t240 GND.t239 GND.t240 GND.t13 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X215 a_9938_8092.t34 a_10060_n1528.t56 GND.t391 GND.t172 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X216 a_10778_8092.t12 a_10060_n1528.t57 GND.t424 GND.t149 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X217 a_21743_n1960.t3 a_9120_14251.t7 a_21659_n106.t8 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X218 a_9938_8092.t33 a_10060_n1528.t58 GND.t400 GND.t70 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X219 GND.t238 GND.t237 GND.t238 GND.t102 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X220 a_10060_n1528.t8 a_10060_n1528.t7 GND.t434 GND.t96 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X221 a_10778_8092.t11 a_10060_n1528.t59 GND.t410 GND.t11 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X222 a_10060_n1528.t6 a_10060_n1528.t5 GND.t339 GND.t175 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X223 a_21659_n106.t18 a_11345_12294.t3 VDD.t20 VDD.t19 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=2u
X224 GND.t236 GND.t235 GND.t236 GND.t99 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X225 a_21743_n2608.t6 a_16964_8348.t12 a_21659_n106.t0 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X226 GND.t234 GND.t233 GND.t234 GND.t105 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X227 GND.t232 GND.t231 GND.t232 GND.t15 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X228 a_9938_8092.t32 a_10060_n1528.t60 GND.t373 GND.t172 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X229 a_21743_n2608.t5 a_16964_8348.t13 a_21659_n106.t3 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X230 GND.t230 GND.t229 GND.t230 GND.t5 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X231 GND.t1 GND.t2 GND.t0 ppolyf_u_1k r_width=1u r_length=98u
X232 a_21743_6748.t7 a_9248_11691.t6 a_21659_3242.t25 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X233 a_9938_8092.t31 a_10060_n1528.t61 GND.t376 GND.t149 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X234 GND.t228 GND.t227 GND.t228 GND.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X235 a_16434_7468.t13 a_16434_7468.t12 VDD.t282 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X236 VDD.t18 a_11345_12294.t3 a_21659_n106.t17 VDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0.52p ps=2.52u w=2u l=2u
X237 a_9120_15571# a_28848_15131# GND.t0 ppolyf_u_1k r_width=1u r_length=98u
X238 a_16964_8348.t1 a_19582_6479.t3 a_10460_8092.t0 GND.t379 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X239 VDD.t166 VDD.t165 VDD.t166 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X240 GND.t226 GND.t225 GND.t226 GND.t112 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X241 GND.t224 GND.t222 GND.t224 GND.t223 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X242 a_11618_8092.t1 a_10060_n1528.t62 GND.t414 GND.t96 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X243 GND.t221 GND.t220 GND.t221 GND.t89 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X244 a_10778_8092.t10 a_10060_n1528.t63 GND.t413 GND.t96 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X245 VDD.t164 VDD.t163 VDD.t164 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X246 GND.t219 GND.t218 GND.t219 GND.t112 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X247 a_9938_8092.t30 a_10060_n1528.t64 GND.t425 GND.t149 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X248 a_16434_7468.t11 a_16434_7468.t10 VDD.t273 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X249 VDD.t17 a_11345_12294.t3 a_21659_n106.t16 VDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0.52p ps=2.52u w=2u l=2u
X250 GND.t217 GND.t216 GND.t217 GND.t112 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X251 a_9938_8092.t29 a_10060_n1528.t65 GND.t389 GND.t204 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X252 GND.t215 GND.t214 GND.t215 GND.t73 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X253 GND.t213 GND.t212 GND.t213 GND.t73 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X254 a_10060_n1528.t4 a_10060_n1528.t3 GND.t401 GND.t96 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X255 a_16434_8348.t9 a_16434_7468.t24 VDD.t277 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X256 a_16434_8348.t8 a_16434_7468.t25 VDD.t278 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X257 a_9938_8092.t28 a_10060_n1528.t66 GND.t451 GND.t149 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X258 GND.t211 GND.t210 GND.t211 GND.t70 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X259 a_11345_12294.t0 a_10060_n1528.t67 GND.t408 GND.t407 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X260 a_21659_3242.t18 a_11345_12294.t2 VDD.t15 VDD.t10 pfet_03v3 ad=0.52p pd=2.52u as=1.3p ps=5.3u w=2u l=2u
X261 VDD.t162 VDD.t161 VDD.t162 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X262 VDD.t160 VDD.t159 VDD.t160 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X263 GND.t209 GND.t208 GND.t209 GND.t11 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X264 GND.t207 GND.t206 GND.t207 GND.t99 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X265 GND.t350 a_19582_7363.t4 a_19582_6479.t2 GND.t349 nfet_03v3 ad=0.366p pd=2.42u as=0.366p ps=2.42u w=0.6u l=0.6u
X266 VDD.t158 VDD.t157 VDD.t158 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X267 GND.t205 GND.t203 GND.t205 GND.t204 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X268 VDD.t156 VDD.t155 VDD.t156 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X269 VDD.t154 VDD.t153 VDD.t154 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X270 VDD.t14 a_11345_12294.t2 a_21659_3242.t21 VDD.t8 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=2u
X271 GND.t418 a_10060_n1528.t68 a_11345_12294.t0 GND.t417 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X272 a_16434_8348.t7 a_16434_7468.t26 VDD.t288 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X273 GND.t202 GND.t201 GND.t202 GND.t73 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X274 a_10460_8092.t7 IBIAS.t5 a_9938_8092.t6 GND.t223 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X275 a_10778_8092.t9 a_10060_n1528.t69 GND.t370 GND.t175 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X276 GND.t200 GND.t199 GND.t200 GND.t58 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X277 a_9938_8092.t27 a_10060_n1528.t70 GND.t340 GND.t172 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X278 GND.t198 GND.t197 GND.t198 GND.t41 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X279 a_9938_8092.t26 a_10060_n1528.t71 GND.t353 GND.t13 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X280 VDD.t152 VDD.t151 VDD.t152 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X281 a_9938_8092.t25 a_10060_n1528.t72 GND.t386 GND.t86 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X282 a_10778_8092.t8 a_10060_n1528.t73 GND.t395 GND.t11 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X283 VDD.t150 VDD.t149 VDD.t150 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X284 IBIAS.t1 IBIAS.t0 a_10060_n1528.t0 GND.t276 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X285 GND.t196 GND.t195 GND.t196 GND.t35 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X286 GND.t194 GND.t193 GND.t194 GND.t63 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X287 VDD.t148 VDD.t147 VDD.t148 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X288 VDD.t146 VDD.t145 VDD.t146 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X289 VDD.t144 VDD.t143 VDD.t144 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X290 a_9938_8092.t24 a_10060_n1528.t74 GND.t403 GND.t172 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X291 VDD.t142 VDD.t141 VDD.t142 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X292 GND.t192 GND.t191 GND.t192 GND.t38 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X293 a_16434_8348.t6 a_16434_7468.t27 VDD.t289 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X294 GND.t190 GND.t189 GND.t190 GND.t63 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X295 GND.t188 GND.t187 GND.t188 GND.t5 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X296 GND.t186 GND.t185 GND.t186 GND.t73 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X297 a_9120_14691# a_28848_14251# GND.t0 ppolyf_u_1k r_width=1u r_length=98u
X298 a_9938_8092.t23 a_10060_n1528.t75 GND.t405 GND.t86 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X299 VDD.t140 VDD.t139 VDD.t140 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X300 VDD.t138 VDD.t137 VDD.t138 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X301 a_10778_8092.t7 a_10060_n1528.t76 GND.t338 GND.t96 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X302 GND.t184 GND.t183 GND.t184 GND.t47 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X303 a_10778_8092.t6 a_10060_n1528.t77 GND.t447 GND.t96 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X304 VDD.t136 VDD.t135 VDD.t136 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X305 a_11300_8092.t2 IBIAS.t6 a_10778_8092.t2 GND.t276 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X306 a_10460_8092.t6 IBIAS.t7 a_9938_8092.t3 GND.t44 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X307 VDD.t134 VDD.t133 VDD.t134 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X308 a_9938_8092.t22 a_10060_n1528.t78 GND.t440 GND.t149 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X309 GND.t182 GND.t181 GND.t182 GND.t73 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X310 GND.t180 GND.t179 GND.t180 GND.t3 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X311 a_11300_8092.t1 IBIAS.t8 a_10778_8092.t1 GND.t223 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X312 GND.t178 GND.t177 GND.t178 GND.t96 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X313 a_9938_8092.t21 a_10060_n1528.t79 GND.t360 GND.t149 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X314 GND.t176 GND.t174 GND.t176 GND.t175 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X315 VDD.t132 VDD.t131 VDD.t132 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X316 VDD.t130 VDD.t129 VDD.t130 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X317 a_21743_6748.t11 a_21743_6748.t10 GND.t443 GND.t55 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X318 GND.t173 GND.t171 GND.t173 GND.t172 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X319 a_16434_8348.t5 a_16434_7468.t28 VDD.t290 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X320 a_16964_8348.t0 GND.t27 cap_mim_2f0_m4m5_noshield c_width=42u c_length=10u
X321 a_16434_7468.t9 a_16434_7468.t8 VDD.t272 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X322 GND.t170 GND.t169 GND.t170 GND.t149 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X323 a_9248_11691.t0 a_9248_11691.t0 VDD.t2 VDD.t1 pfet_03v3 ad=3.25p pd=11.299999u as=3.25p ps=11.299999u w=5u l=4u
X324 GND.t168 GND.t167 GND.t168 GND.t112 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X325 VDD.t128 VDD.t127 VDD.t128 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X326 a_21659_3242.t20 a_11345_12294.t2 VDD.t13 VDD.t6 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=2u
X327 a_16434_7468.t7 a_16434_7468.t6 VDD.t281 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X328 GND.t166 GND.t165 GND.t166 GND.t70 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X329 GND.t164 GND.t162 GND.t164 GND.t163 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X330 VDD.t126 VDD.t125 VDD.t126 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X331 GND.t161 GND.t160 GND.t161 GND.t11 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X332 VDD.t124 VDD.t123 VDD.t124 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X333 a_9938_8092.t20 a_10060_n1528.t80 GND.t337 GND.t86 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X334 VDD.t122 VDD.t121 VDD.t122 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X335 a_28935_6098# a_25891_6334.t6 VDD.t38 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X336 a_16434_7468.t5 a_16434_7468.t4 VDD.t287 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X337 VDD.t12 a_11345_12294.t2 a_21659_3242.t16 VDD.t4 pfet_03v3 ad=1.3p pd=5.3u as=0.52p ps=2.52u w=2u l=2u
X338 GND.t159 GND.t158 GND.t159 GND.t86 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X339 GND.t157 GND.t156 GND.t157 GND.t47 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X340 VDD.t120 VDD.t119 VDD.t120 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X341 a_10778_8092.t5 a_10060_n1528.t81 GND.t347 GND.t22 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X342 GND.t155 GND.t154 GND.t155 GND.t96 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X343 GND.t153 GND.t151 GND.t153 GND.t152 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X344 a_21743_n1960.t2 a_9120_14251.t8 a_21659_n106.t13 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X345 VDD.t118 VDD.t117 VDD.t118 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X346 VDD.t116 VDD.t115 VDD.t116 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X347 GND.t150 GND.t148 GND.t150 GND.t149 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X348 GND.t147 GND.t146 GND.t147 GND.t44 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X349 GND.t145 GND.t143 GND.t145 GND.t144 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X350 VDD.t114 VDD.t113 VDD.t114 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X351 a_21743_6100.t9 a_21743_6100.t8 GND.t358 GND.t55 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X352 a_19582_7363.t1 a_21743_n1960.t16 GND.t422 GND.t32 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X353 a_21743_n1960.t0 a_21743_n2608.t16 GND.t18 GND.t17 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X354 VDD.t112 VDD.t111 VDD.t112 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X355 GND.t142 GND.t141 GND.t142 GND.t135 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X356 GND.t140 GND.t139 GND.t140 GND.t58 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X357 a_25891_n1726.t3 a_21743_n2608.t17 GND.t363 GND.t32 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X358 a_9938_8092.t19 a_10060_n1528.t82 GND.t352 GND.t13 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X359 GND.t138 GND.t137 GND.t138 GND.t73 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X360 a_11345_12294.t0 a_10060_n1528.t83 GND.t26 GND.t25 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X361 a_21743_n2608.t12 a_21743_n1960.t17 GND.t385 GND.t17 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X362 VDD.t110 VDD.t109 VDD.t110 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X363 GND.t136 GND.t134 GND.t136 GND.t135 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X364 GND.t133 GND.t132 GND.t133 GND.t102 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X365 GND.t131 GND.t130 GND.t131 GND.t13 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X366 GND.t129 GND.t128 GND.t129 GND.t73 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X367 VDD.t108 VDD.t107 VDD.t108 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X368 VDD.t106 VDD.t105 VDD.t106 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X369 GND.t437 a_10060_n1528.t84 a_11345_12294.t0 GND.t436 nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X370 GND.t127 GND.t126 GND.t127 GND.t70 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X371 GND.t125 GND.t124 GND.t125 GND.t38 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X372 VDD.t104 VDD.t103 VDD.t104 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X373 a_21743_6100.t0 a_16964_8348.t14 a_21659_3242.t3 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X374 GND.t123 GND.t122 GND.t123 GND.t47 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X375 VDD.t102 VDD.t101 VDD.t102 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X376 a_9938_8092.t18 a_10060_n1528.t85 GND.t432 GND.t11 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X377 GND.t121 GND.t120 GND.t121 GND.t89 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X378 GND.t119 GND.t118 GND.t119 GND.t44 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X379 VDD.t100 VDD.t99 VDD.t100 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X380 GND.t117 GND.t116 GND.t117 GND.t50 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X381 GND.t115 GND.t114 GND.t115 GND.t7 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X382 a_16434_8348.t4 a_16434_7468.t29 VDD.t283 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X383 VDD.t98 VDD.t97 VDD.t98 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X384 VDD.t96 VDD.t95 VDD.t96 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X385 GND.t113 GND.t111 GND.t113 GND.t112 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X386 a_9938_8092.t17 a_10060_n1528.t86 GND.t439 GND.t86 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X387 GND.t110 GND.t109 GND.t110 GND.t58 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X388 a_21743_6748.t8 a_9248_11691.t7 a_21659_3242.t26 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X389 a_21743_n2608.t4 a_16964_8348.t15 a_21659_n106.t6 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X390 VDD.t94 VDD.t93 VDD.t94 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X391 VDD.t92 VDD.t91 VDD.t92 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X392 GND.t108 GND.t107 GND.t108 GND.t73 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X393 GND.t106 GND.t104 GND.t106 GND.t105 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X394 a_10460_8092.t5 IBIAS.t9 a_9938_8092.t4 GND.t223 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X395 VDD.t90 VDD.t89 VDD.t90 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X396 GND.t103 GND.t101 GND.t103 GND.t102 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X397 VDD.t88 VDD.t87 VDD.t88 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X398 VDD.t86 VDD.t85 VDD.t86 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X399 GND.t100 GND.t98 GND.t100 GND.t99 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X400 OUT.t0 a_19582_6479.t4 a_19718_6163# VDD.t3 pfet_03v3 ad=0.39p pd=2.5u as=0.39p ps=2.5u w=0.6u l=0.6u
X401 VDD.t84 VDD.t83 VDD.t84 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X402 VDD.t82 VDD.t81 VDD.t82 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X403 VDD.t80 VDD.t79 VDD.t80 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X404 VDD.t78 VDD.t77 VDD.t78 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X405 GND.t97 GND.t95 GND.t97 GND.t96 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X406 GND.t94 GND.t93 GND.t94 GND.t38 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X407 a_9120_14251.t0 IBIAS.t10 a_11618_8092.t0 GND.t223 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X408 GND.t92 GND.t91 GND.t92 GND.t47 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X409 VDD.t76 VDD.t75 VDD.t76 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X410 a_10460_8092.t4 IBIAS.t11 a_9938_8092.t1 GND.t44 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X411 VDD.t74 VDD.t73 VDD.t74 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X412 a_21743_6100.t6 a_16964_8348.t16 a_21659_3242.t2 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X413 GND.t90 GND.t88 GND.t90 GND.t89 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X414 VDD.t72 VDD.t71 VDD.t72 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X415 GND.t87 GND.t85 GND.t87 GND.t86 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X416 a_21743_6748.t9 a_9248_11691.t8 a_21659_3242.t27 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X417 VDD.t70 VDD.t69 VDD.t70 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X418 a_21743_n1960.t1 a_9120_14251.t9 a_21659_n106.t12 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X419 a_21743_6100.t1 a_16964_8348.t17 a_21659_3242.t1 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X420 VDD.t68 VDD.t67 VDD.t68 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X421 a_9120_15571# a_9248_11691.t1 GND.t0 ppolyf_u_1k r_width=1u r_length=98u
X422 GND.t84 GND.t83 GND.t84 GND.t9 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X423 a_21659_3242.t19 a_11345_12294.t2 VDD.t11 VDD.t10 pfet_03v3 ad=0.52p pd=2.52u as=1.3p ps=5.3u w=2u l=2u
X424 GND.t82 GND.t81 GND.t82 GND.t73 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X425 GND.t80 GND.t78 GND.t80 GND.t79 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X426 GND.t77 GND.t75 GND.t77 GND.t76 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X427 a_16434_7468.t3 a_16434_7468.t2 VDD.t286 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X428 a_19582_6043.t0 a_21743_6100.t17 GND.t4 GND.t3 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X429 VDD.t66 VDD.t65 VDD.t66 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X430 GND.t74 GND.t72 GND.t74 GND.t73 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X431 a_9938_8092.t16 a_10060_n1528.t87 GND.t351 GND.t204 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X432 VDD.t9 a_11345_12294.t2 a_21659_3242.t17 VDD.t8 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=2u
X433 a_9938_8092.t15 a_10060_n1528.t88 GND.t336 GND.t70 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X434 VDD.t64 VDD.t63 VDD.t64 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X435 VDD.t62 VDD.t61 VDD.t62 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X436 GND.t71 GND.t69 GND.t71 GND.t70 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X437 a_9938_8092.t14 a_10060_n1528.t89 GND.t442 GND.t11 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X438 a_16964_8348.t0 a_11300_8092.t9 a_16434_8348.t0 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X439 VDD.t60 VDD.t59 VDD.t60 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X440 GND.t68 GND.t67 GND.t68 GND.t15 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X441 VDD.t58 VDD.t57 VDD.t58 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X442 GND.t66 GND.t65 GND.t66 GND.t50 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X443 GND.t64 GND.t62 GND.t64 GND.t63 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X444 GND.t61 GND.t60 GND.t61 GND.t11 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X445 a_9938_8092.t13 a_10060_n1528.t90 GND.t344 GND.t204 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X446 a_19718_6163# a_19582_6043.t4 VDD.t266 VDD.t265 pfet_03v3 ad=0.39p pd=2.5u as=0.39p ps=2.5u w=0.6u l=0.6u
X447 a_21743_n2608.t1 a_21743_n2608.t0 GND.t380 GND.t163 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X448 VDD.t56 VDD.t55 VDD.t56 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X449 a_9938_8092.t12 a_10060_n1528.t91 GND.t430 GND.t204 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X450 VDD.t54 VDD.t53 VDD.t54 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X451 VDD.t52 VDD.t51 VDD.t52 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X452 GND.t59 GND.t57 GND.t59 GND.t58 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X453 a_21743_n1960.t11 a_21743_n1960.t10 GND.t383 GND.t163 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X454 a_9938_8092.t11 a_10060_n1528.t92 GND.t441 GND.t86 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X455 VDD.t50 VDD.t49 VDD.t50 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X456 a_25891_6334.t0 a_21743_6748.t17 GND.t429 GND.t3 nfet_03v3 ad=0.672p pd=3.44u as=0.672p ps=3.44u w=0.6u l=0.6u
X457 GND.t56 GND.t54 GND.t56 GND.t55 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X458 a_16434_8348.t3 a_16434_7468.t30 VDD.t284 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X459 a_9120_14691# a_28848_15131# GND.t0 ppolyf_u_1k r_width=1u r_length=98u
X460 a_21743_6100.t2 a_16964_8348.t18 a_21659_3242.t0 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X461 a_10460_8092.t3 IBIAS.t12 a_9938_8092.t2 GND.t58 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X462 VDD.t48 VDD.t47 VDD.t48 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X463 GND.t53 GND.t52 GND.t53 GND.t38 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X464 VDD.t46 VDD.t45 VDD.t46 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X465 VDD.t44 VDD.t43 VDD.t44 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X466 GND.t51 GND.t49 GND.t51 GND.t50 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X467 a_21743_6748.t6 a_9248_11691.t9 a_21659_3242.t24 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0.696p ps=3.52u w=0.6u l=0.6u
X468 a_9938_8092.t10 a_10060_n1528.t93 GND.t374 GND.t204 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X469 GND.t48 GND.t46 GND.t48 GND.t47 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X470 GND.t45 GND.t43 GND.t45 GND.t44 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X471 a_9938_8092.t9 a_10060_n1528.t94 GND.t378 GND.t204 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X472 a_21659_3242.t22 a_11345_12294.t2 VDD.t7 VDD.t6 pfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=2u
X473 a_16434_8348.t2 a_16434_7468.t31 VDD.t285 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X474 VDD.t42 VDD.t41 VDD.t42 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X475 GND.t42 GND.t40 GND.t42 GND.t41 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X476 GND.t366 a_19582_6479.t5 OUT.t0 GND.t365 nfet_03v3 ad=0.366p pd=2.42u as=0.366p ps=2.42u w=0.6u l=0.6u
X477 a_10060_n1528.t2 a_10060_n1528.t1 GND.t341 GND.t175 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X478 VDD.t40 VDD.t39 VDD.t40 w_23841_n458# pfet_03v3 ad=0.696p pd=3.52u as=0 ps=0 w=0.6u l=0.6u
X479 GND.t39 GND.t37 GND.t39 GND.t38 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X480 VDD.t5 a_11345_12294.t2 a_21659_3242.t14 VDD.t4 pfet_03v3 ad=1.3p pd=5.3u as=0.52p ps=2.52u w=2u l=2u
X481 a_10778_8092.t4 a_10060_n1528.t95 GND.t438 GND.t149 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X482 GND.t36 GND.t34 GND.t36 GND.t35 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
X483 a_10460_8092.t2 IBIAS.t13 a_9938_8092.t0 GND.t47 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X484 a_9938_8092.t8 a_10060_n1528.t96 GND.t412 GND.t172 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X485 a_11300_8092.t5 a_11300_8092.t4 a_16434_7468.t0 w_15348_6286# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X486 a_11300_8092.t0 IBIAS.t14 a_10778_8092.t0 GND.t44 nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=2u
X487 GND.t33 GND.t31 GND.t33 GND.t32 nfet_03v3 ad=0.672p pd=3.44u as=0 ps=0 w=0.6u l=0.6u
R0 a_16964_8348.n2 a_16964_8348.t13 20.1527
R1 a_16964_8348.n3 a_16964_8348.t12 19.2698
R2 a_16964_8348.n3 a_16964_8348.t6 19.2698
R3 a_16964_8348.n2 a_16964_8348.t11 19.2698
R4 a_16964_8348.n1 a_16964_8348.t7 19.2698
R5 a_16964_8348.n0 a_16964_8348.t8 19.2698
R6 a_16964_8348.n0 a_16964_8348.t14 19.2698
R7 a_16964_8348.n1 a_16964_8348.t10 19.2698
R8 a_16964_8348.n0 a_16964_8348.t3 17.8802
R9 a_16964_8348.n3 a_16964_8348.t15 16.9973
R10 a_16964_8348.n3 a_16964_8348.t4 16.9973
R11 a_16964_8348.n2 a_16964_8348.t5 16.9973
R12 a_16964_8348.n2 a_16964_8348.t9 16.9973
R13 a_16964_8348.n1 a_16964_8348.t17 16.9973
R14 a_16964_8348.n1 a_16964_8348.t18 16.9973
R15 a_16964_8348.n0 a_16964_8348.t16 16.9973
R16 a_16964_8348.t0 a_16964_8348.n1 13.7866
R17 a_16964_8348.n1 a_16964_8348.n0 13.0644
R18 a_16964_8348.t0 a_16964_8348.t2 11.5231
R19 a_16964_8348.n3 a_16964_8348.n2 11.4691
R20 a_16964_8348.n1 a_16964_8348.n3 11.078
R21 a_16964_8348.t0 a_16964_8348.t1 7.91829
R22 GND.n358 GND.n324 1.93097e+06
R23 GND.t38 GND.n358 1.13917e+06
R24 GND.n328 GND.n327 656338
R25 GND.n330 GND.n329 371800
R26 GND.n329 GND.n328 354412
R27 GND.t135 GND.n326 23177.7
R28 GND.n328 GND.t73 12601.6
R29 GND.n361 GND.n360 9225.03
R30 GND.n340 GND.n333 3687.83
R31 GND.t417 GND.t407 3018.24
R32 GND.n376 GND.n375 2831.47
R33 GND.n357 GND.n331 2687.63
R34 GND.t345 GND.n324 2409.2
R35 GND.t0 GND.n330 2340.02
R36 GND.n331 GND.t345 2161.28
R37 GND.t392 GND.t365 1630.46
R38 GND.t436 GND.t25 1619.22
R39 GND.t349 GND.t392 1586.79
R40 GND.t365 GND.t367 1586.79
R41 GND.n365 GND.t379 1580.25
R42 GND.n376 GND.t73 1411.95
R43 GND.n375 GND.n317 1295.63
R44 GND.n376 GND.n316 1245.9
R45 GND.n331 GND.t449 1159.48
R46 GND.n376 GND.t349 1026.32
R47 GND.t367 GND.n316 1026.32
R48 GND.n331 GND.t0 913.669
R49 GND.n331 GND.t417 856.966
R50 GND.t394 GND.n361 765.518
R51 GND.t144 GND.t105 591.636
R52 GND.t58 GND.t50 527.13
R53 GND.t44 GND.t223 527.13
R54 GND.t276 GND.t47 527.13
R55 GND.t47 GND.t38 527.13
R56 GND.n359 GND.t223 509.558
R57 GND.n331 GND.t436 459.743
R58 GND.n324 GND.t58 456.217
R59 GND.t3 GND.t102 445.05
R60 GND.t89 GND.t35 445.05
R61 GND.t35 GND.t7 445.05
R62 GND.t7 GND.t79 445.05
R63 GND.t79 GND.t55 445.05
R64 GND.t55 GND.t99 445.05
R65 GND.t15 GND.t135 418.409
R66 GND.t32 GND.t15 418.409
R67 GND.t105 GND.t41 418.409
R68 GND.t41 GND.t17 418.409
R69 GND.t17 GND.t76 418.409
R70 GND.t76 GND.t163 418.409
R71 GND.t163 GND.t63 418.409
R72 GND.t394 GND.n317 389.656
R73 GND.n326 GND.t152 367.813
R74 GND.t102 GND.n329 353.632
R75 GND.n327 GND.t144 286.49
R76 GND.t379 GND.n317 283.875
R77 GND.n329 GND.t89 275.676
R78 GND.t63 GND.t73 245.894
R79 GND.t86 GND.t172 234.697
R80 GND.t172 GND.t149 234.697
R81 GND.t149 GND.t22 234.697
R82 GND.t22 GND.t175 234.697
R83 GND.t175 GND.t96 234.697
R84 GND.t96 GND.t5 234.697
R85 GND.t5 GND.t11 234.697
R86 GND.t11 GND.t13 234.697
R87 GND.t204 GND.t70 234.697
R88 GND.t70 GND.t112 234.697
R89 GND.t13 GND.n359 226.875
R90 GND.n330 GND.n325 202.703
R91 GND.n360 GND.t86 180.494
R92 GND.n325 GND.t9 177.601
R93 GND.n376 GND.n312 176.462
R94 GND.n327 GND.t32 131.919
R95 GND.n326 GND.n325 105.168
R96 GND.n369 GND.n323 78.4742
R97 GND.n370 GND.n323 78.4742
R98 GND.n374 GND.n318 78.4742
R99 GND.n365 GND.n318 78.4742
R100 GND.n324 GND.t44 70.9119
R101 GND.n3029 GND.n1 68.0662
R102 GND.n360 GND.t73 54.2044
R103 GND.n374 GND.n319 42.0005
R104 GND.n370 GND.n319 42.0005
R105 GND.n365 GND.n362 42.0005
R106 GND.n369 GND.n362 42.0005
R107 GND.t99 GND.n312 40.3952
R108 GND.n355 GND.n336 36.6672
R109 GND.n351 GND.n335 36.6672
R110 GND.n349 GND.n333 36.6672
R111 GND.n364 GND.n362 36.4742
R112 GND.n364 GND.n319 36.4742
R113 GND.n361 GND.n323 21.5568
R114 GND.n343 GND.n342 21.1987
R115 GND.n359 GND.t276 17.5715
R116 GND.n499 GND.n449 16.0495
R117 GND.n316 GND.n315 15.0643
R118 GND.n311 GND.t350 15.0005
R119 GND.n313 GND.t393 15.0005
R120 GND.n314 GND.t366 15.0005
R121 GND.n315 GND.t368 15.0005
R122 GND.n345 GND.n344 14.9575
R123 GND.n377 GND.n376 14.9005
R124 GND.n389 GND.t98 14.6214
R125 GND.n215 GND.t151 14.6214
R126 GND.t62 GND.n809 14.6204
R127 GND.t332 GND.n573 14.6204
R128 GND.t143 GND.n99 14.6096
R129 GND.n222 GND.t330 14.6096
R130 GND.t104 GND.n99 14.6087
R131 GND.n222 GND.t328 14.6087
R132 GND.n100 GND.t143 14.6073
R133 GND.n102 GND.t265 14.6073
R134 GND.t265 GND.n101 14.6073
R135 GND.n104 GND.t271 14.6073
R136 GND.t271 GND.n103 14.6073
R137 GND.n113 GND.t324 14.6073
R138 GND.t324 GND.n105 14.6073
R139 GND.t237 GND.n197 14.6073
R140 GND.n198 GND.t237 14.6073
R141 GND.n202 GND.t132 14.6073
R142 GND.t132 GND.n201 14.6073
R143 GND.n204 GND.t101 14.6073
R144 GND.t101 GND.n203 14.6073
R145 GND.t330 GND.n205 14.6073
R146 GND.n810 GND.t62 14.606
R147 GND.n812 GND.t189 14.606
R148 GND.t189 GND.n811 14.606
R149 GND.n814 GND.t193 14.606
R150 GND.t193 GND.n813 14.606
R151 GND.t288 GND.n87 14.606
R152 GND.n815 GND.t288 14.606
R153 GND.n574 GND.t332 14.606
R154 GND.n576 GND.t134 14.606
R155 GND.t134 GND.n575 14.606
R156 GND.n578 GND.t141 14.606
R157 GND.t141 GND.n577 14.606
R158 GND.n580 GND.t247 14.606
R159 GND.t247 GND.n579 14.606
R160 GND.n383 GND.t304 14.606
R161 GND.t304 GND.n382 14.606
R162 GND.n385 GND.t235 14.606
R163 GND.t235 GND.n384 14.606
R164 GND.n387 GND.t206 14.606
R165 GND.t206 GND.n386 14.606
R166 GND.t98 GND.n388 14.606
R167 GND.n209 GND.t326 14.606
R168 GND.n448 GND.t326 14.606
R169 GND.n211 GND.t278 14.606
R170 GND.t278 GND.n210 14.606
R171 GND.n213 GND.t261 14.606
R172 GND.t261 GND.n212 14.606
R173 GND.t151 GND.n214 14.606
R174 GND.n793 GND.n792 14.2055
R175 GND.n786 GND.n785 14.2055
R176 GND.n791 GND.n790 14.2055
R177 GND.n779 GND.n778 14.2055
R178 GND.n784 GND.n783 14.2055
R179 GND.n115 GND.n114 14.2055
R180 GND.n777 GND.n776 14.2055
R181 GND.n418 GND.n417 14.2055
R182 GND.n200 GND.n199 14.2055
R183 GND.n411 GND.n410 14.2055
R184 GND.n416 GND.n415 14.2055
R185 GND.n404 GND.n403 14.2055
R186 GND.n409 GND.n408 14.2055
R187 GND.n402 GND.n401 14.2055
R188 GND.n347 GND.t2 11.69
R189 GND.n343 GND.t19 11.6812
R190 GND.n344 GND.t1 11.6779
R191 GND.n342 GND.t20 11.6773
R192 GND.n703 GND.n94 11.6555
R193 GND.n702 GND.n696 11.6555
R194 GND.n695 GND.n694 11.6555
R195 GND.n693 GND.n680 11.6555
R196 GND.n679 GND.n678 11.6555
R197 GND.n677 GND.n664 11.6555
R198 GND.n662 GND.n108 11.6555
R199 GND.n616 GND.n615 11.6555
R200 GND.n614 GND.n133 11.6555
R201 GND.n593 GND.n141 11.6555
R202 GND.n592 GND.n147 11.6555
R203 GND.n428 GND.n189 11.6555
R204 GND.n429 GND.n187 11.6555
R205 GND.n437 GND.n436 11.6555
R206 GND.n445 GND.n444 11.6555
R207 GND.n306 GND.n232 11.6555
R208 GND.n305 GND.n236 11.6555
R209 GND.n297 GND.n296 11.6555
R210 GND.n286 GND.n285 11.6555
R211 GND.n278 GND.n277 11.6555
R212 GND.n276 GND.n248 11.6555
R213 GND.n258 GND.n257 11.6555
R214 GND.n1078 GND.n1077 10.2176
R215 GND.n793 GND.t104 9.4905
R216 GND.n786 GND.t233 9.4905
R217 GND.n790 GND.t233 9.4905
R218 GND.n779 GND.t241 9.4905
R219 GND.n783 GND.t241 9.4905
R220 GND.n114 GND.t308 9.4905
R221 GND.n776 GND.t308 9.4905
R222 GND.n418 GND.t220 9.4905
R223 GND.t220 GND.n200 9.4905
R224 GND.n411 GND.t120 9.4905
R225 GND.n415 GND.t120 9.4905
R226 GND.n404 GND.t88 9.4905
R227 GND.n408 GND.t88 9.4905
R228 GND.n401 GND.t328 9.4905
R229 GND.n1978 GND.n1445 9.2465
R230 GND.n2953 GND.n1445 9.2465
R231 GND.n1684 GND.n1683 9.2465
R232 GND.n1684 GND.n1446 9.2465
R233 GND.n1107 GND.t386 8.844
R234 GND.n1100 GND.t373 8.844
R235 GND.n1093 GND.t451 8.844
R236 GND.n1086 GND.t452 8.844
R237 GND.n1116 GND.t401 8.844
R238 GND.n1123 GND.t420 8.844
R239 GND.n1130 GND.t12 8.844
R240 GND.n1137 GND.t14 8.844
R241 GND.n1144 GND.t378 8.844
R242 GND.n1151 GND.t427 8.844
R243 GND.n290 GND.t428 8.61761
R244 GND.n245 GND.t357 8.61761
R245 GND.n264 GND.t445 8.61761
R246 GND.n659 GND.t361 8.61761
R247 GND.n673 GND.t385 8.61761
R248 GND.n689 GND.t446 8.61761
R249 GND.n233 GND.t358 8.61578
R250 GND.n705 GND.t383 8.61578
R251 GND.n184 GND.t343 8.60755
R252 GND.n142 GND.t421 8.60755
R253 GND.n193 GND.t429 8.60204
R254 GND.n130 GND.t363 8.60204
R255 GND.n193 GND.t4 8.30644
R256 GND.n130 GND.t422 8.30644
R257 GND.n184 GND.t10 8.30099
R258 GND.n142 GND.t16 8.30099
R259 GND.n233 GND.t443 8.28997
R260 GND.n290 GND.t342 8.28997
R261 GND.n245 GND.t8 8.28997
R262 GND.n264 GND.t356 8.28997
R263 GND.n659 GND.t382 8.28997
R264 GND.n673 GND.t18 8.28997
R265 GND.n689 GND.t372 8.28997
R266 GND.n705 GND.t380 8.28997
R267 GND.n663 GND.t42 8.28759
R268 GND.t33 GND.n98 8.28759
R269 GND.n570 GND.t33 8.28759
R270 GND.t232 GND.n571 8.28759
R271 GND.n572 GND.t232 8.28759
R272 GND.n808 GND.t303 8.28759
R273 GND.n806 GND.t303 8.28759
R274 GND.n805 GND.t252 8.28759
R275 GND.n803 GND.t252 8.28759
R276 GND.n802 GND.t335 8.28759
R277 GND.n800 GND.t335 8.28759
R278 GND.n799 GND.t198 8.28759
R279 GND.n797 GND.t198 8.28759
R280 GND.t56 GND.n390 8.28759
R281 GND.n391 GND.t56 8.28759
R282 GND.t254 GND.n392 8.28759
R283 GND.n393 GND.t254 8.28759
R284 GND.t287 GND.n394 8.28759
R285 GND.n395 GND.t287 8.28759
R286 GND.t196 GND.n396 8.28759
R287 GND.n397 GND.t196 8.28759
R288 GND.n221 GND.t311 8.28759
R289 GND.n219 GND.t311 8.28759
R290 GND.n218 GND.t260 8.28759
R291 GND.n216 GND.t260 8.28759
R292 GND.n268 GND.t36 8.28759
R293 GND.t306 GND.n46 8.06917
R294 GND.n339 GND.t306 8.06917
R295 GND.t263 GND.n46 8.06917
R296 GND.n339 GND.t263 8.06917
R297 GND.t57 GND.n1328 8.06917
R298 GND.n1329 GND.t57 8.06917
R299 GND.n1328 GND.t322 8.06917
R300 GND.n1329 GND.t322 8.06917
R301 GND.t109 GND.n1326 8.06917
R302 GND.n1327 GND.t109 8.06917
R303 GND.n1326 GND.t49 8.06917
R304 GND.n1327 GND.t49 8.06917
R305 GND.t316 GND.n1324 8.06917
R306 GND.n1325 GND.t316 8.06917
R307 GND.n1301 GND.t85 8.06917
R308 GND.t85 GND.n55 8.06917
R309 GND.n1301 GND.t107 8.06917
R310 GND.t107 GND.n55 8.06917
R311 GND.t158 GND.n1299 8.06917
R312 GND.n1300 GND.t158 8.06917
R313 GND.n1299 GND.t181 8.06917
R314 GND.n1300 GND.t181 8.06917
R315 GND.t212 GND.n1297 8.06917
R316 GND.n1298 GND.t212 8.06917
R317 GND.t137 GND.n1295 8.06917
R318 GND.n1296 GND.t137 8.06917
R319 GND.t201 GND.n1293 8.06917
R320 GND.n1294 GND.t201 8.06917
R321 GND.t214 GND.n1291 8.06917
R322 GND.n1292 GND.t214 8.06917
R323 GND.t185 GND.n1289 8.06917
R324 GND.n1290 GND.t185 8.06917
R325 GND.t81 GND.n1287 8.06917
R326 GND.n1288 GND.t81 8.06917
R327 GND.t312 GND.n1285 8.06917
R328 GND.n1286 GND.t312 8.06917
R329 GND.n1285 GND.t128 8.06917
R330 GND.n1286 GND.t128 8.06917
R331 GND.t282 GND.n1283 8.06917
R332 GND.n1284 GND.t282 8.06917
R333 GND.n1283 GND.t72 8.06917
R334 GND.n1284 GND.t72 8.06917
R335 GND.n1374 GND.t280 8.06917
R336 GND.t280 GND.n1373 8.06917
R337 GND.n1374 GND.t126 8.06917
R338 GND.n1373 GND.t126 8.06917
R339 GND.t218 GND.n5 8.06917
R340 GND.n1375 GND.t218 8.06917
R341 GND.t69 GND.n5 8.06917
R342 GND.n1375 GND.t69 8.06917
R343 GND.n1362 GND.t298 8.06917
R344 GND.t298 GND.n1361 8.06917
R345 GND.n1364 GND.t243 8.06917
R346 GND.t243 GND.n1363 8.06917
R347 GND.n1366 GND.t294 8.06917
R348 GND.t294 GND.n1365 8.06917
R349 GND.n1368 GND.t111 8.06917
R350 GND.t111 GND.n1367 8.06917
R351 GND.n1370 GND.t284 8.06917
R352 GND.t284 GND.n1369 8.06917
R353 GND.n1372 GND.t225 8.06917
R354 GND.t225 GND.n1371 8.06917
R355 GND.n1351 GND.t124 8.06917
R356 GND.t124 GND.n1350 8.06917
R357 GND.n1351 GND.t122 8.06917
R358 GND.n1350 GND.t122 8.06917
R359 GND.n1351 GND.t275 8.06917
R360 GND.n1350 GND.t275 8.06917
R361 GND.n1353 GND.t167 8.06917
R362 GND.t167 GND.n1352 8.06917
R363 GND.n1353 GND.t165 8.06917
R364 GND.n1352 GND.t165 8.06917
R365 GND.n1353 GND.t300 8.06917
R366 GND.n1352 GND.t300 8.06917
R367 GND.n1356 GND.t216 8.06917
R368 GND.t216 GND.n1355 8.06917
R369 GND.n1356 GND.t210 8.06917
R370 GND.n1355 GND.t210 8.06917
R371 GND.n1356 GND.t320 8.06917
R372 GND.n1355 GND.t320 8.06917
R373 GND.n1346 GND.t37 8.06917
R374 GND.t37 GND.n1345 8.06917
R375 GND.n1340 GND.t296 8.06917
R376 GND.t296 GND.n1339 8.06917
R377 GND.n1340 GND.t156 8.06917
R378 GND.n1339 GND.t156 8.06917
R379 GND.n1342 GND.t52 8.06917
R380 GND.t52 GND.n1341 8.06917
R381 GND.n1342 GND.t46 8.06917
R382 GND.n1341 GND.t46 8.06917
R383 GND.n1344 GND.t93 8.06917
R384 GND.t93 GND.n1343 8.06917
R385 GND.n1344 GND.t91 8.06917
R386 GND.n1343 GND.t91 8.06917
R387 GND.n1331 GND.t146 8.06917
R388 GND.t146 GND.n44 8.06917
R389 GND.n776 GND.n775 8.0005
R390 GND.n114 GND.n107 8.0005
R391 GND.n783 GND.n782 8.0005
R392 GND.n780 GND.n779 8.0005
R393 GND.n790 GND.n789 8.0005
R394 GND.n787 GND.n786 8.0005
R395 GND.n794 GND.n793 8.0005
R396 GND.n401 GND.n400 8.0005
R397 GND.n408 GND.n407 8.0005
R398 GND.n405 GND.n404 8.0005
R399 GND.n415 GND.n414 8.0005
R400 GND.n412 GND.n411 8.0005
R401 GND.n200 GND.n196 8.0005
R402 GND.n419 GND.n418 8.0005
R403 GND.n1107 GND.t439 7.91829
R404 GND.n1108 GND.t405 7.91829
R405 GND.n1109 GND.t441 7.91829
R406 GND.n1110 GND.t337 7.91829
R407 GND.n1111 GND.t431 7.91829
R408 GND.n1100 GND.t415 7.91829
R409 GND.n1101 GND.t340 7.91829
R410 GND.n1102 GND.t377 7.91829
R411 GND.n1103 GND.t403 7.91829
R412 GND.n1104 GND.t391 7.91829
R413 GND.n1105 GND.t426 7.91829
R414 GND.n1106 GND.t412 7.91829
R415 GND.n1093 GND.t448 7.91829
R416 GND.n1094 GND.t440 7.91829
R417 GND.n1095 GND.t424 7.91829
R418 GND.n1096 GND.t438 7.91829
R419 GND.n1097 GND.t425 7.91829
R420 GND.n1098 GND.t360 7.91829
R421 GND.n1099 GND.t376 7.91829
R422 GND.n1086 GND.t384 7.91829
R423 GND.n1087 GND.t359 7.91829
R424 GND.n1088 GND.t23 7.91829
R425 GND.n1089 GND.t347 7.91829
R426 GND.n1090 GND.t435 7.91829
R427 GND.n1091 GND.t396 7.91829
R428 GND.n1092 GND.t398 7.91829
R429 GND.n1078 GND.t339 7.91829
R430 GND.n1079 GND.t399 7.91829
R431 GND.n1080 GND.t370 7.91829
R432 GND.n1081 GND.t348 7.91829
R433 GND.n1082 GND.t416 7.91829
R434 GND.n1083 GND.t409 7.91829
R435 GND.n1084 GND.t419 7.91829
R436 GND.n1085 GND.t341 7.91829
R437 GND.n1076 GND.t450 7.91829
R438 GND.n1077 GND.t346 7.91829
R439 GND.n1116 GND.t404 7.91829
R440 GND.n1117 GND.t447 7.91829
R441 GND.n1118 GND.t423 7.91829
R442 GND.n1119 GND.t414 7.91829
R443 GND.n1120 GND.t413 7.91829
R444 GND.n1121 GND.t338 7.91829
R445 GND.n1122 GND.t434 7.91829
R446 GND.n1123 GND.t371 7.91829
R447 GND.n1124 GND.t402 7.91829
R448 GND.n1125 GND.t362 7.91829
R449 GND.n1126 GND.t6 7.91829
R450 GND.n1127 GND.t381 7.91829
R451 GND.n1128 GND.t387 7.91829
R452 GND.n1129 GND.t364 7.91829
R453 GND.n1130 GND.t388 7.91829
R454 GND.n1131 GND.t410 7.91829
R455 GND.n1132 GND.t433 7.91829
R456 GND.n1133 GND.t395 7.91829
R457 GND.n1134 GND.t21 7.91829
R458 GND.n1135 GND.t442 7.91829
R459 GND.n1136 GND.t432 7.91829
R460 GND.n1137 GND.t406 7.91829
R461 GND.n1138 GND.t369 7.91829
R462 GND.n1139 GND.t354 7.91829
R463 GND.n1140 GND.t390 7.91829
R464 GND.n1141 GND.t24 7.91829
R465 GND.n1142 GND.t352 7.91829
R466 GND.n1143 GND.t353 7.91829
R467 GND.n1144 GND.t351 7.91829
R468 GND.n1145 GND.t375 7.91829
R469 GND.n1146 GND.t430 7.91829
R470 GND.n1147 GND.t344 7.91829
R471 GND.n1148 GND.t374 7.91829
R472 GND.n1149 GND.t389 7.91829
R473 GND.n1150 GND.t397 7.91829
R474 GND.n1151 GND.t400 7.91829
R475 GND.n1152 GND.t355 7.91829
R476 GND.n1153 GND.t411 7.91829
R477 GND.n1154 GND.t444 7.91829
R478 GND.n1155 GND.t336 7.91829
R479 GND.n359 GND.t204 7.82375
R480 GND.n330 GND.t3 7.53391
R481 GND.n2954 GND.n2953 7.35912
R482 GND.n149 GND.t67 7.30624
R483 GND.n135 GND.t255 7.30624
R484 GND.n798 GND.t197 7.30624
R485 GND.n801 GND.t334 7.30624
R486 GND.n804 GND.t251 7.30624
R487 GND.n807 GND.t302 7.30624
R488 GND.n568 GND.t231 7.30624
R489 GND.n569 GND.t31 7.30624
R490 GND.n764 GND.t40 7.30624
R491 GND.n747 GND.t249 7.30624
R492 GND.n730 GND.t75 7.30624
R493 GND.n713 GND.t162 7.30624
R494 GND.n217 GND.t259 7.30624
R495 GND.n220 GND.t310 7.30624
R496 GND.n260 GND.t34 7.30624
R497 GND.n251 GND.t114 7.30624
R498 GND.n241 GND.t78 7.30624
R499 GND.n238 GND.t267 7.30624
R500 GND.n179 GND.t83 7.30624
R501 GND.n190 GND.t179 7.30624
R502 GND.n223 GND.t195 7.30624
R503 GND.n224 GND.t286 7.30624
R504 GND.n225 GND.t253 7.30624
R505 GND.n226 GND.t54 7.30624
R506 GND.n592 GND.n591 6.3005
R507 GND.n594 GND.n593 6.3005
R508 GND.n614 GND.n613 6.3005
R509 GND.n615 GND.n132 6.3005
R510 GND.n662 GND.n655 6.3005
R511 GND.n677 GND.n669 6.3005
R512 GND.n678 GND.n670 6.3005
R513 GND.n693 GND.n685 6.3005
R514 GND.n694 GND.n686 6.3005
R515 GND.n702 GND.n701 6.3005
R516 GND.n704 GND.n703 6.3005
R517 GND.n259 GND.n258 6.3005
R518 GND.n276 GND.n275 6.3005
R519 GND.n277 GND.n247 6.3005
R520 GND.n287 GND.n286 6.3005
R521 GND.n296 GND.n295 6.3005
R522 GND.n305 GND.n304 6.3005
R523 GND.n307 GND.n306 6.3005
R524 GND.n444 GND.n443 6.3005
R525 GND.n438 GND.n437 6.3005
R526 GND.n430 GND.n429 6.3005
R527 GND.n428 GND.n427 6.3005
R528 GND.n1686 GND.n1685 6.16867
R529 GND.n1685 GND.n1444 6.16866
R530 GND.n1978 GND.n1977 5.79988
R531 GND.n337 GND.n336 5.2005
R532 GND.n355 GND.n354 5.2005
R533 GND.n353 GND.n335 5.2005
R534 GND.n352 GND.n351 5.2005
R535 GND.n350 GND.n349 5.2005
R536 GND.n348 GND.n333 5.2005
R537 GND.n357 GND.n333 5.2005
R538 GND.n341 GND.n340 5.2005
R539 GND.n1075 GND.n1073 4.98524
R540 GND.n494 GND.n493 4.5005
R541 GND.n493 GND.n453 4.5005
R542 GND.n496 GND.n453 4.5005
R543 GND.n380 GND.n379 4.5005
R544 GND.n309 GND.n308 4.5005
R545 GND.n235 GND.n234 4.5005
R546 GND.n303 GND.n302 4.5005
R547 GND.n301 GND.n237 4.5005
R548 GND.n300 GND.n299 4.5005
R549 GND.n298 GND.n239 4.5005
R550 GND.n292 GND.n240 4.5005
R551 GND.n294 GND.n293 4.5005
R552 GND.n289 GND.n288 4.5005
R553 GND.n243 GND.n242 4.5005
R554 GND.n284 GND.n283 4.5005
R555 GND.n282 GND.n244 4.5005
R556 GND.n280 GND.n279 4.5005
R557 GND.n250 GND.n246 4.5005
R558 GND.n274 GND.n273 4.5005
R559 GND.n272 GND.n249 4.5005
R560 GND.n271 GND.n270 4.5005
R561 GND.n269 GND.n252 4.5005
R562 GND.n267 GND.n266 4.5005
R563 GND.n263 GND.n253 4.5005
R564 GND.n262 GND.n261 4.5005
R565 GND.n256 GND.n255 4.5005
R566 GND.n254 GND.n195 4.5005
R567 GND.n423 GND.n422 4.5005
R568 GND.n426 GND.n425 4.5005
R569 GND.n192 GND.n191 4.5005
R570 GND.n188 GND.n186 4.5005
R571 GND.n432 GND.n431 4.5005
R572 GND.n433 GND.n183 4.5005
R573 GND.n435 GND.n434 4.5005
R574 GND.n182 GND.n181 4.5005
R575 GND.n440 GND.n439 4.5005
R576 GND.n442 GND.n441 4.5005
R577 GND.n180 GND.n178 4.5005
R578 GND.n446 GND.n176 4.5005
R579 GND.n831 GND.n84 4.5005
R580 GND.n832 GND.n831 4.5005
R581 GND.n831 GND.n830 4.5005
R582 GND.n831 GND.n91 4.5005
R583 GND.n831 GND.n90 4.5005
R584 GND.n831 GND.n89 4.5005
R585 GND.n831 GND.n88 4.5005
R586 GND.n819 GND.n818 4.5005
R587 GND.n708 GND.n707 4.5005
R588 GND.n712 GND.n711 4.5005
R589 GND.n715 GND.n714 4.5005
R590 GND.n700 GND.n697 4.5005
R591 GND.n721 GND.n720 4.5005
R592 GND.n723 GND.n722 4.5005
R593 GND.n692 GND.n687 4.5005
R594 GND.n729 GND.n728 4.5005
R595 GND.n732 GND.n731 4.5005
R596 GND.n684 GND.n681 4.5005
R597 GND.n738 GND.n737 4.5005
R598 GND.n740 GND.n739 4.5005
R599 GND.n676 GND.n671 4.5005
R600 GND.n746 GND.n745 4.5005
R601 GND.n749 GND.n748 4.5005
R602 GND.n668 GND.n665 4.5005
R603 GND.n755 GND.n754 4.5005
R604 GND.n757 GND.n756 4.5005
R605 GND.n657 GND.n656 4.5005
R606 GND.n763 GND.n762 4.5005
R607 GND.n766 GND.n765 4.5005
R608 GND.n654 GND.n110 4.5005
R609 GND.n772 GND.n771 4.5005
R610 GND.n648 GND.n647 4.5005
R611 GND.n647 GND.n112 4.5005
R612 GND.n647 GND.n122 4.5005
R613 GND.n647 GND.n123 4.5005
R614 GND.n647 GND.n120 4.5005
R615 GND.n647 GND.n124 4.5005
R616 GND.n647 GND.n119 4.5005
R617 GND.n647 GND.n125 4.5005
R618 GND.n647 GND.n118 4.5005
R619 GND.n647 GND.n126 4.5005
R620 GND.n647 GND.n117 4.5005
R621 GND.n647 GND.n127 4.5005
R622 GND.n647 GND.n116 4.5005
R623 GND.n647 GND.n646 4.5005
R624 GND.n620 GND.n106 4.5005
R625 GND.n618 GND.n617 4.5005
R626 GND.n138 GND.n137 4.5005
R627 GND.n612 GND.n611 4.5005
R628 GND.n605 GND.n134 4.5005
R629 GND.n604 GND.n603 4.5005
R630 GND.n602 GND.n601 4.5005
R631 GND.n596 GND.n595 4.5005
R632 GND.n146 GND.n145 4.5005
R633 GND.n590 GND.n589 4.5005
R634 GND.n150 GND.n148 4.5005
R635 GND.n583 GND.n582 4.5005
R636 GND.n564 GND.n157 4.5005
R637 GND.n564 GND.n156 4.5005
R638 GND.n564 GND.n158 4.5005
R639 GND.n564 GND.n155 4.5005
R640 GND.n564 GND.n159 4.5005
R641 GND.n564 GND.n154 4.5005
R642 GND.n564 GND.n563 4.5005
R643 GND.n1408 GND.n2 4.5005
R644 GND.n1409 GND.n1408 4.5005
R645 GND.n1408 GND.n12 4.5005
R646 GND.n1408 GND.n11 4.5005
R647 GND.n1408 GND.n13 4.5005
R648 GND.n1408 GND.n10 4.5005
R649 GND.n1408 GND.n14 4.5005
R650 GND.n1408 GND.n9 4.5005
R651 GND.n1408 GND.n15 4.5005
R652 GND.n1408 GND.n8 4.5005
R653 GND.n1408 GND.n16 4.5005
R654 GND.n1408 GND.n7 4.5005
R655 GND.n1408 GND.n17 4.5005
R656 GND.n1408 GND.n6 4.5005
R657 GND.n1408 GND.n1407 4.5005
R658 GND.n1379 GND.n1378 4.5005
R659 GND.n21 GND.n20 4.5005
R660 GND.n1005 GND.n1004 4.5005
R661 GND.n984 GND.n983 4.5005
R662 GND.n998 GND.n997 4.5005
R663 GND.n995 GND.n994 4.5005
R664 GND.n988 GND.n987 4.5005
R665 GND.n989 GND.n982 4.5005
R666 GND.n1009 GND.n1008 4.5005
R667 GND.n979 GND.n978 4.5005
R668 GND.n1015 GND.n1014 4.5005
R669 GND.n1018 GND.n1017 4.5005
R670 GND.n977 GND.n974 4.5005
R671 GND.n1024 GND.n1023 4.5005
R672 GND.n1026 GND.n1025 4.5005
R673 GND.n972 GND.n969 4.5005
R674 GND.n1032 GND.n1031 4.5005
R675 GND.n1034 GND.n1033 4.5005
R676 GND.n967 GND.n964 4.5005
R677 GND.n1040 GND.n1039 4.5005
R678 GND.n1042 GND.n1041 4.5005
R679 GND.n959 GND.n958 4.5005
R680 GND.n1048 GND.n1047 4.5005
R681 GND.n1050 GND.n1049 4.5005
R682 GND.n932 GND.n930 4.5005
R683 GND.n1056 GND.n1055 4.5005
R684 GND.n951 GND.n929 4.5005
R685 GND.n950 GND.n949 4.5005
R686 GND.n948 GND.n947 4.5005
R687 GND.n940 GND.n936 4.5005
R688 GND.n942 GND.n941 4.5005
R689 GND.n938 GND.n928 4.5005
R690 GND.n1060 GND.n1059 4.5005
R691 GND.n927 GND.n924 4.5005
R692 GND.n1066 GND.n1065 4.5005
R693 GND.n1068 GND.n1067 4.5005
R694 GND.n922 GND.n919 4.5005
R695 GND.n1164 GND.n1163 4.5005
R696 GND.n1166 GND.n1165 4.5005
R697 GND.n917 GND.n914 4.5005
R698 GND.n1172 GND.n1171 4.5005
R699 GND.n1174 GND.n1173 4.5005
R700 GND.n909 GND.n908 4.5005
R701 GND.n1180 GND.n1179 4.5005
R702 GND.n1182 GND.n1181 4.5005
R703 GND.n904 GND.n903 4.5005
R704 GND.n1188 GND.n1187 4.5005
R705 GND.n1190 GND.n1189 4.5005
R706 GND.n881 GND.n879 4.5005
R707 GND.n1196 GND.n1195 4.5005
R708 GND.n896 GND.n878 4.5005
R709 GND.n895 GND.n894 4.5005
R710 GND.n893 GND.n892 4.5005
R711 GND.n886 GND.n885 4.5005
R712 GND.n887 GND.n877 4.5005
R713 GND.n1200 GND.n1199 4.5005
R714 GND.n874 GND.n873 4.5005
R715 GND.n1206 GND.n1205 4.5005
R716 GND.n1209 GND.n1208 4.5005
R717 GND.n870 GND.n869 4.5005
R718 GND.n1215 GND.n1214 4.5005
R719 GND.n1218 GND.n1217 4.5005
R720 GND.n868 GND.n865 4.5005
R721 GND.n1224 GND.n1223 4.5005
R722 GND.n1226 GND.n1225 4.5005
R723 GND.n863 GND.n860 4.5005
R724 GND.n1232 GND.n1231 4.5005
R725 GND.n1234 GND.n1233 4.5005
R726 GND.n858 GND.n855 4.5005
R727 GND.n1240 GND.n1239 4.5005
R728 GND.n1242 GND.n1241 4.5005
R729 GND.n850 GND.n849 4.5005
R730 GND.n1248 GND.n1247 4.5005
R731 GND.n1250 GND.n1249 4.5005
R732 GND.n1282 GND.n73 4.5005
R733 GND.n1282 GND.n72 4.5005
R734 GND.n1282 GND.n74 4.5005
R735 GND.n1282 GND.n71 4.5005
R736 GND.n1282 GND.n75 4.5005
R737 GND.n1282 GND.n70 4.5005
R738 GND.n1282 GND.n76 4.5005
R739 GND.n1282 GND.n69 4.5005
R740 GND.n1282 GND.n77 4.5005
R741 GND.n1282 GND.n68 4.5005
R742 GND.n1282 GND.n78 4.5005
R743 GND.n1282 GND.n67 4.5005
R744 GND.n1282 GND.n79 4.5005
R745 GND.n1282 GND.n66 4.5005
R746 GND.n1282 GND.n1281 4.5005
R747 GND.n3025 GND.n1419 4.5005
R748 GND.n3025 GND.n3024 4.5005
R749 GND.n3029 GND.n3028 4.5005
R750 GND.n1414 GND.n0 4.5005
R751 GND.n1413 GND.n1412 4.5005
R752 GND.n1411 GND.n1410 4.5005
R753 GND.n4 GND.n3 4.5005
R754 GND.n1384 GND.n1383 4.5005
R755 GND.n1386 GND.n1385 4.5005
R756 GND.n1388 GND.n1387 4.5005
R757 GND.n1390 GND.n1389 4.5005
R758 GND.n1392 GND.n1391 4.5005
R759 GND.n1394 GND.n1393 4.5005
R760 GND.n1396 GND.n1395 4.5005
R761 GND.n1398 GND.n1397 4.5005
R762 GND.n1400 GND.n1399 4.5005
R763 GND.n1402 GND.n1401 4.5005
R764 GND.n1404 GND.n1403 4.5005
R765 GND.n1406 GND.n1405 4.5005
R766 GND.n1382 GND.n18 4.5005
R767 GND.n1381 GND.n1380 4.5005
R768 GND.n1003 GND.n19 4.5005
R769 GND.n1002 GND.n1001 4.5005
R770 GND.n1000 GND.n999 4.5005
R771 GND.n986 GND.n985 4.5005
R772 GND.n993 GND.n992 4.5005
R773 GND.n991 GND.n990 4.5005
R774 GND.n981 GND.n980 4.5005
R775 GND.n1011 GND.n1010 4.5005
R776 GND.n1013 GND.n1012 4.5005
R777 GND.n976 GND.n975 4.5005
R778 GND.n1020 GND.n1019 4.5005
R779 GND.n1022 GND.n1021 4.5005
R780 GND.n971 GND.n970 4.5005
R781 GND.n1028 GND.n1027 4.5005
R782 GND.n1030 GND.n1029 4.5005
R783 GND.n966 GND.n965 4.5005
R784 GND.n1036 GND.n1035 4.5005
R785 GND.n1038 GND.n1037 4.5005
R786 GND.n961 GND.n960 4.5005
R787 GND.n1044 GND.n1043 4.5005
R788 GND.n1046 GND.n1045 4.5005
R789 GND.n956 GND.n955 4.5005
R790 GND.n1052 GND.n1051 4.5005
R791 GND.n1054 GND.n1053 4.5005
R792 GND.n954 GND.n931 4.5005
R793 GND.n953 GND.n952 4.5005
R794 GND.n934 GND.n933 4.5005
R795 GND.n946 GND.n945 4.5005
R796 GND.n944 GND.n943 4.5005
R797 GND.n939 GND.n937 4.5005
R798 GND.n926 GND.n925 4.5005
R799 GND.n1062 GND.n1061 4.5005
R800 GND.n1064 GND.n1063 4.5005
R801 GND.n921 GND.n920 4.5005
R802 GND.n1070 GND.n1069 4.5005
R803 GND.n1072 GND.n1071 4.5005
R804 GND.n916 GND.n915 4.5005
R805 GND.n1168 GND.n1167 4.5005
R806 GND.n1170 GND.n1169 4.5005
R807 GND.n911 GND.n910 4.5005
R808 GND.n1176 GND.n1175 4.5005
R809 GND.n1178 GND.n1177 4.5005
R810 GND.n906 GND.n905 4.5005
R811 GND.n1184 GND.n1183 4.5005
R812 GND.n1186 GND.n1185 4.5005
R813 GND.n901 GND.n900 4.5005
R814 GND.n1192 GND.n1191 4.5005
R815 GND.n1194 GND.n1193 4.5005
R816 GND.n899 GND.n880 4.5005
R817 GND.n898 GND.n897 4.5005
R818 GND.n883 GND.n882 4.5005
R819 GND.n891 GND.n890 4.5005
R820 GND.n889 GND.n888 4.5005
R821 GND.n876 GND.n875 4.5005
R822 GND.n1202 GND.n1201 4.5005
R823 GND.n1204 GND.n1203 4.5005
R824 GND.n872 GND.n871 4.5005
R825 GND.n1211 GND.n1210 4.5005
R826 GND.n1213 GND.n1212 4.5005
R827 GND.n867 GND.n866 4.5005
R828 GND.n1220 GND.n1219 4.5005
R829 GND.n1222 GND.n1221 4.5005
R830 GND.n862 GND.n861 4.5005
R831 GND.n1228 GND.n1227 4.5005
R832 GND.n1230 GND.n1229 4.5005
R833 GND.n857 GND.n856 4.5005
R834 GND.n1236 GND.n1235 4.5005
R835 GND.n1238 GND.n1237 4.5005
R836 GND.n852 GND.n851 4.5005
R837 GND.n1244 GND.n1243 4.5005
R838 GND.n1246 GND.n1245 4.5005
R839 GND.n848 GND.n847 4.5005
R840 GND.n1252 GND.n1251 4.5005
R841 GND.n1254 GND.n1253 4.5005
R842 GND.n1256 GND.n1255 4.5005
R843 GND.n1258 GND.n1257 4.5005
R844 GND.n1260 GND.n1259 4.5005
R845 GND.n1262 GND.n1261 4.5005
R846 GND.n1264 GND.n1263 4.5005
R847 GND.n1266 GND.n1265 4.5005
R848 GND.n1268 GND.n1267 4.5005
R849 GND.n1270 GND.n1269 4.5005
R850 GND.n1272 GND.n1271 4.5005
R851 GND.n1274 GND.n1273 4.5005
R852 GND.n1276 GND.n1275 4.5005
R853 GND.n1278 GND.n1277 4.5005
R854 GND.n1280 GND.n1279 4.5005
R855 GND.n846 GND.n80 4.5005
R856 GND.n845 GND.n844 4.5005
R857 GND.n843 GND.n81 4.5005
R858 GND.n842 GND.n841 4.5005
R859 GND.n840 GND.n82 4.5005
R860 GND.n839 GND.n838 4.5005
R861 GND.n837 GND.n83 4.5005
R862 GND.n836 GND.n835 4.5005
R863 GND.n834 GND.n833 4.5005
R864 GND.n86 GND.n85 4.5005
R865 GND.n829 GND.n828 4.5005
R866 GND.n827 GND.n826 4.5005
R867 GND.n825 GND.n824 4.5005
R868 GND.n823 GND.n822 4.5005
R869 GND.n821 GND.n820 4.5005
R870 GND.n93 GND.n92 4.5005
R871 GND.n710 GND.n709 4.5005
R872 GND.n699 GND.n698 4.5005
R873 GND.n717 GND.n716 4.5005
R874 GND.n719 GND.n718 4.5005
R875 GND.n691 GND.n688 4.5005
R876 GND.n725 GND.n724 4.5005
R877 GND.n727 GND.n726 4.5005
R878 GND.n683 GND.n682 4.5005
R879 GND.n734 GND.n733 4.5005
R880 GND.n736 GND.n735 4.5005
R881 GND.n675 GND.n672 4.5005
R882 GND.n742 GND.n741 4.5005
R883 GND.n744 GND.n743 4.5005
R884 GND.n667 GND.n666 4.5005
R885 GND.n751 GND.n750 4.5005
R886 GND.n753 GND.n752 4.5005
R887 GND.n661 GND.n658 4.5005
R888 GND.n759 GND.n758 4.5005
R889 GND.n761 GND.n760 4.5005
R890 GND.n653 GND.n652 4.5005
R891 GND.n768 GND.n767 4.5005
R892 GND.n770 GND.n769 4.5005
R893 GND.n651 GND.n109 4.5005
R894 GND.n650 GND.n649 4.5005
R895 GND.n121 GND.n111 4.5005
R896 GND.n625 GND.n624 4.5005
R897 GND.n627 GND.n626 4.5005
R898 GND.n629 GND.n628 4.5005
R899 GND.n631 GND.n630 4.5005
R900 GND.n633 GND.n632 4.5005
R901 GND.n635 GND.n634 4.5005
R902 GND.n637 GND.n636 4.5005
R903 GND.n639 GND.n638 4.5005
R904 GND.n641 GND.n640 4.5005
R905 GND.n643 GND.n642 4.5005
R906 GND.n645 GND.n644 4.5005
R907 GND.n623 GND.n128 4.5005
R908 GND.n622 GND.n621 4.5005
R909 GND.n131 GND.n129 4.5005
R910 GND.n610 GND.n609 4.5005
R911 GND.n608 GND.n136 4.5005
R912 GND.n607 GND.n606 4.5005
R913 GND.n140 GND.n139 4.5005
R914 GND.n600 GND.n599 4.5005
R915 GND.n598 GND.n597 4.5005
R916 GND.n588 GND.n144 4.5005
R917 GND.n587 GND.n586 4.5005
R918 GND.n585 GND.n584 4.5005
R919 GND.n152 GND.n151 4.5005
R920 GND.n552 GND.n551 4.5005
R921 GND.n554 GND.n553 4.5005
R922 GND.n556 GND.n555 4.5005
R923 GND.n558 GND.n557 4.5005
R924 GND.n560 GND.n559 4.5005
R925 GND.n562 GND.n561 4.5005
R926 GND.n550 GND.n160 4.5005
R927 GND.n549 GND.n548 4.5005
R928 GND.n547 GND.n161 4.5005
R929 GND.n546 GND.n545 4.5005
R930 GND.n544 GND.n162 4.5005
R931 GND.n543 GND.n542 4.5005
R932 GND.n541 GND.n163 4.5005
R933 GND.n540 GND.n539 4.5005
R934 GND.n538 GND.n164 4.5005
R935 GND.n537 GND.n536 4.5005
R936 GND.n535 GND.n165 4.5005
R937 GND.n534 GND.n533 4.5005
R938 GND.n532 GND.n166 4.5005
R939 GND.n531 GND.n530 4.5005
R940 GND.n529 GND.n167 4.5005
R941 GND.n528 GND.n527 4.5005
R942 GND.n526 GND.n168 4.5005
R943 GND.n525 GND.n524 4.5005
R944 GND.n523 GND.n169 4.5005
R945 GND.n522 GND.n521 4.5005
R946 GND.n520 GND.n170 4.5005
R947 GND.n519 GND.n518 4.5005
R948 GND.n517 GND.n171 4.5005
R949 GND.n516 GND.n515 4.5005
R950 GND.n514 GND.n172 4.5005
R951 GND.n513 GND.n512 4.5005
R952 GND.n511 GND.n173 4.5005
R953 GND.n510 GND.n509 4.5005
R954 GND.n508 GND.n174 4.5005
R955 GND.n507 GND.n506 4.5005
R956 GND.n505 GND.n175 4.5005
R957 GND.n504 GND.n503 4.5005
R958 GND.n502 GND.n501 4.5005
R959 GND.n500 GND.n1 4.5005
R960 GND.n1075 GND.n1074 4.35135
R961 GND.n1076 GND.n1075 4.31387
R962 GND.n703 GND.t164 4.2005
R963 GND.t164 GND.n702 4.2005
R964 GND.n694 GND.t77 4.2005
R965 GND.t77 GND.n693 4.2005
R966 GND.n678 GND.t250 4.2005
R967 GND.t250 GND.n677 4.2005
R968 GND.t42 GND.n662 4.2005
R969 GND.n615 GND.t256 4.2005
R970 GND.t256 GND.n614 4.2005
R971 GND.n593 GND.t68 4.2005
R972 GND.t68 GND.n592 4.2005
R973 GND.t180 GND.n428 4.2005
R974 GND.n429 GND.t180 4.2005
R975 GND.n437 GND.t84 4.2005
R976 GND.n444 GND.t84 4.2005
R977 GND.n306 GND.t268 4.2005
R978 GND.t268 GND.n305 4.2005
R979 GND.n296 GND.t80 4.2005
R980 GND.n286 GND.t80 4.2005
R981 GND.n277 GND.t115 4.2005
R982 GND.t115 GND.n276 4.2005
R983 GND.n258 GND.t36 4.2005
R984 GND.n97 GND.t64 4.14649
R985 GND.n96 GND.t190 4.14649
R986 GND.n95 GND.t194 4.14649
R987 GND.n816 GND.t289 4.14649
R988 GND.n795 GND.t106 4.14649
R989 GND.n788 GND.t234 4.14649
R990 GND.n781 GND.t242 4.14649
R991 GND.n774 GND.t309 4.14649
R992 GND.n567 GND.t333 4.14649
R993 GND.n566 GND.t136 4.14649
R994 GND.n565 GND.t142 4.14649
R995 GND.n153 GND.t248 4.14649
R996 GND.n230 GND.t305 4.14649
R997 GND.n229 GND.t236 4.14649
R998 GND.n228 GND.t207 4.14649
R999 GND.n227 GND.t100 4.14649
R1000 GND.n420 GND.t221 4.14649
R1001 GND.n413 GND.t121 4.14649
R1002 GND.n406 GND.t90 4.14649
R1003 GND.n399 GND.t329 4.14649
R1004 GND.n177 GND.t327 4.14649
R1005 GND.n208 GND.t279 4.14649
R1006 GND.n207 GND.t262 4.14649
R1007 GND.n206 GND.t153 4.14649
R1008 GND.n774 GND.t325 4.14549
R1009 GND.n781 GND.t272 4.14549
R1010 GND.n788 GND.t266 4.14549
R1011 GND.n795 GND.t145 4.14549
R1012 GND.n399 GND.t331 4.14549
R1013 GND.n406 GND.t103 4.14549
R1014 GND.n413 GND.t133 4.14549
R1015 GND.n420 GND.t238 4.14549
R1016 GND.n336 GND.n332 4.05199
R1017 GND.n356 GND.n355 4.05199
R1018 GND.n351 GND.n334 4.05199
R1019 GND.n356 GND.n335 4.05199
R1020 GND.n349 GND.n334 4.05199
R1021 GND.n340 GND.n332 4.05199
R1022 GND.n1357 GND.t269 4.05092
R1023 GND.n36 GND.t183 4.0509
R1024 GND.n1319 GND.t199 4.0509
R1025 GND.n43 GND.t222 4.03583
R1026 GND.n42 GND.t292 4.03583
R1027 GND.n37 GND.t191 4.03583
R1028 GND.n29 GND.t273 4.03583
R1029 GND.n854 GND.t314 4.03583
R1030 GND.n1216 GND.t169 4.03583
R1031 GND.n884 GND.t245 4.03583
R1032 GND.n907 GND.t318 4.03583
R1033 GND.n918 GND.t177 4.03583
R1034 GND.n935 GND.t257 4.03583
R1035 GND.n962 GND.t60 4.03583
R1036 GND.n973 GND.t130 4.03583
R1037 GND.n996 GND.t203 4.03583
R1038 GND.n54 GND.t171 4.03583
R1039 GND.n53 GND.t148 4.03583
R1040 GND.n52 GND.t227 4.03583
R1041 GND.n51 GND.t174 4.03583
R1042 GND.n50 GND.t154 4.03583
R1043 GND.n1314 GND.t229 4.03583
R1044 GND.n1315 GND.t208 4.03583
R1045 GND.n50 GND.t95 4.03583
R1046 GND.n1314 GND.t187 4.03583
R1047 GND.n1315 GND.t160 4.03583
R1048 GND.n50 GND.t65 4.03583
R1049 GND.n1314 GND.t139 4.03583
R1050 GND.n1315 GND.t118 4.03583
R1051 GND.n1322 GND.t116 4.03583
R1052 GND.n45 GND.t43 4.03533
R1053 GND.n31 GND.t239 4.03533
R1054 GND.n33 GND.t290 4.03533
R1055 GND.n344 GND.n343 3.92729
R1056 GND.n347 GND.n346 3.92607
R1057 GND.n358 GND.n357 3.91751
R1058 GND.n1360 GND.t274 3.37894
R1059 GND.n1323 GND.t117 3.37892
R1060 GND.t192 GND.n1347 3.37892
R1061 GND.n1321 GND.t117 3.3605
R1062 GND.t119 GND.n32 3.3605
R1063 GND.n1316 GND.t119 3.3605
R1064 GND.t140 GND.n1317 3.3605
R1065 GND.n1318 GND.t140 3.3605
R1066 GND.n1313 GND.t66 3.3605
R1067 GND.t66 GND.n1312 3.3605
R1068 GND.t161 GND.n32 3.3605
R1069 GND.n1316 GND.t161 3.3605
R1070 GND.n1317 GND.t188 3.3605
R1071 GND.n1318 GND.t188 3.3605
R1072 GND.n1313 GND.t97 3.3605
R1073 GND.n1312 GND.t97 3.3605
R1074 GND.t209 GND.n32 3.3605
R1075 GND.n1316 GND.t209 3.3605
R1076 GND.n1317 GND.t230 3.3605
R1077 GND.n1318 GND.t230 3.3605
R1078 GND.n1313 GND.t155 3.3605
R1079 GND.n1312 GND.t155 3.3605
R1080 GND.n1311 GND.t176 3.3605
R1081 GND.t176 GND.n1310 3.3605
R1082 GND.n1309 GND.t228 3.3605
R1083 GND.t228 GND.n1308 3.3605
R1084 GND.n1307 GND.t150 3.3605
R1085 GND.t150 GND.n1306 3.3605
R1086 GND.n1305 GND.t173 3.3605
R1087 GND.t173 GND.n1304 3.3605
R1088 GND.t205 GND.n1006 3.3605
R1089 GND.n1007 GND.t205 3.3605
R1090 GND.n1016 GND.t131 3.3605
R1091 GND.t131 GND.n968 3.3605
R1092 GND.n963 GND.t61 3.3605
R1093 GND.t61 GND.n957 3.3605
R1094 GND.t258 GND.n1057 3.3605
R1095 GND.n1058 GND.t258 3.3605
R1096 GND.n923 GND.t178 3.3605
R1097 GND.t178 GND.n913 3.3605
R1098 GND.n912 GND.t319 3.3605
R1099 GND.t319 GND.n902 3.3605
R1100 GND.t246 GND.n1197 3.3605
R1101 GND.n1198 GND.t246 3.3605
R1102 GND.n1207 GND.t170 3.3605
R1103 GND.t170 GND.n864 3.3605
R1104 GND.n859 GND.t315 3.3605
R1105 GND.t315 GND.n853 3.3605
R1106 GND.t274 GND.n1359 3.3605
R1107 GND.n1348 GND.t192 3.3605
R1108 GND.n1337 GND.t293 3.3605
R1109 GND.t293 GND.n1336 3.3605
R1110 GND.n1335 GND.t224 3.3605
R1111 GND.t224 GND.n1334 3.3605
R1112 GND.n424 GND.n193 3.2947
R1113 GND.n185 GND.n184 3.27989
R1114 GND.n281 GND.n245 3.24384
R1115 GND.n291 GND.n290 3.24341
R1116 GND.n265 GND.n264 3.24341
R1117 GND.n310 GND.n233 3.24335
R1118 GND.n619 GND.n130 3.20256
R1119 GND.n143 GND.n142 3.18774
R1120 GND.n1112 GND.n1111 3.16121
R1121 GND.n1156 GND.n1155 3.16121
R1122 GND.n674 GND.n673 3.15269
R1123 GND.n660 GND.n659 3.15227
R1124 GND.n706 GND.n705 3.1522
R1125 GND.n690 GND.n689 3.15127
R1126 GND.n488 GND.t28 3.15121
R1127 GND.t28 GND.n487 3.15121
R1128 GND.n2954 GND.n1444 2.96543
R1129 GND.n1687 GND.n1686 2.65676
R1130 GND.n2956 GND.n1443 2.46014
R1131 GND.n490 GND.n489 2.4452
R1132 GND.n2768 GND.n2740 2.29025
R1133 GND.n2160 GND.n1621 2.288
R1134 GND.n2499 GND.n1508 2.288
R1135 GND.n1940 GND.n1939 2.2505
R1136 GND.n1938 GND.n1700 2.2505
R1137 GND.n1937 GND.n1936 2.2505
R1138 GND.n1935 GND.n1701 2.2505
R1139 GND.n1934 GND.n1933 2.2505
R1140 GND.n1932 GND.n1702 2.2505
R1141 GND.n1931 GND.n1930 2.2505
R1142 GND.n1929 GND.n1703 2.2505
R1143 GND.n1928 GND.n1927 2.2505
R1144 GND.n1926 GND.n1704 2.2505
R1145 GND.n1925 GND.n1924 2.2505
R1146 GND.n1923 GND.n1705 2.2505
R1147 GND.n1922 GND.n1921 2.2505
R1148 GND.n1920 GND.n1706 2.2505
R1149 GND.n1919 GND.n1918 2.2505
R1150 GND.n1917 GND.n1707 2.2505
R1151 GND.n1916 GND.n1915 2.2505
R1152 GND.n1914 GND.n1708 2.2505
R1153 GND.n1913 GND.n1912 2.2505
R1154 GND.n1911 GND.n1709 2.2505
R1155 GND.n1910 GND.n1909 2.2505
R1156 GND.n1908 GND.n1710 2.2505
R1157 GND.n1907 GND.n1906 2.2505
R1158 GND.n1905 GND.n1711 2.2505
R1159 GND.n1904 GND.n1903 2.2505
R1160 GND.n1902 GND.n1712 2.2505
R1161 GND.n1901 GND.n1900 2.2505
R1162 GND.n1899 GND.n1713 2.2505
R1163 GND.n1898 GND.n1897 2.2505
R1164 GND.n1896 GND.n1714 2.2505
R1165 GND.n1895 GND.n1894 2.2505
R1166 GND.n1893 GND.n1715 2.2505
R1167 GND.n1892 GND.n1891 2.2505
R1168 GND.n1890 GND.n1716 2.2505
R1169 GND.n1889 GND.n1888 2.2505
R1170 GND.n1887 GND.n1717 2.2505
R1171 GND.n1886 GND.n1885 2.2505
R1172 GND.n1884 GND.n1718 2.2505
R1173 GND.n1883 GND.n1882 2.2505
R1174 GND.n1881 GND.n1719 2.2505
R1175 GND.n1880 GND.n1879 2.2505
R1176 GND.n1878 GND.n1720 2.2505
R1177 GND.n1877 GND.n1876 2.2505
R1178 GND.n1875 GND.n1721 2.2505
R1179 GND.n1874 GND.n1873 2.2505
R1180 GND.n1872 GND.n1722 2.2505
R1181 GND.n1871 GND.n1870 2.2505
R1182 GND.n1869 GND.n1723 2.2505
R1183 GND.n1868 GND.n1867 2.2505
R1184 GND.n1866 GND.n1724 2.2505
R1185 GND.n1865 GND.n1864 2.2505
R1186 GND.n1863 GND.n1725 2.2505
R1187 GND.n1862 GND.n1861 2.2505
R1188 GND.n1860 GND.n1726 2.2505
R1189 GND.n1859 GND.n1858 2.2505
R1190 GND.n1857 GND.n1727 2.2505
R1191 GND.n1856 GND.n1855 2.2505
R1192 GND.n1854 GND.n1728 2.2505
R1193 GND.n1853 GND.n1852 2.2505
R1194 GND.n1851 GND.n1729 2.2505
R1195 GND.n1850 GND.n1849 2.2505
R1196 GND.n1848 GND.n1730 2.2505
R1197 GND.n1847 GND.n1846 2.2505
R1198 GND.n1845 GND.n1731 2.2505
R1199 GND.n1844 GND.n1843 2.2505
R1200 GND.n1842 GND.n1732 2.2505
R1201 GND.n1841 GND.n1840 2.2505
R1202 GND.n1839 GND.n1733 2.2505
R1203 GND.n1838 GND.n1837 2.2505
R1204 GND.n1836 GND.n1734 2.2505
R1205 GND.n1835 GND.n1834 2.2505
R1206 GND.n1833 GND.n1735 2.2505
R1207 GND.n1832 GND.n1831 2.2505
R1208 GND.n1830 GND.n1736 2.2505
R1209 GND.n1829 GND.n1828 2.2505
R1210 GND.n1827 GND.n1737 2.2505
R1211 GND.n1826 GND.n1825 2.2505
R1212 GND.n1824 GND.n1738 2.2505
R1213 GND.n1823 GND.n1822 2.2505
R1214 GND.n1821 GND.n1739 2.2505
R1215 GND.n1820 GND.n1819 2.2505
R1216 GND.n1818 GND.n1740 2.2505
R1217 GND.n1817 GND.n1816 2.2505
R1218 GND.n1815 GND.n1741 2.2505
R1219 GND.n1814 GND.n1813 2.2505
R1220 GND.n1812 GND.n1742 2.2505
R1221 GND.n1811 GND.n1810 2.2505
R1222 GND.n1809 GND.n1743 2.2505
R1223 GND.n1808 GND.n1807 2.2505
R1224 GND.n1806 GND.n1744 2.2505
R1225 GND.n1805 GND.n1804 2.2505
R1226 GND.n1803 GND.n1745 2.2505
R1227 GND.n1802 GND.n1801 2.2505
R1228 GND.n1800 GND.n1746 2.2505
R1229 GND.n1799 GND.n1798 2.2505
R1230 GND.n1797 GND.n1747 2.2505
R1231 GND.n1796 GND.n1795 2.2505
R1232 GND.n1794 GND.n1748 2.2505
R1233 GND.n1793 GND.n1792 2.2505
R1234 GND.n1791 GND.n1749 2.2505
R1235 GND.n1790 GND.n1789 2.2505
R1236 GND.n1788 GND.n1750 2.2505
R1237 GND.n1787 GND.n1786 2.2505
R1238 GND.n1785 GND.n1751 2.2505
R1239 GND.n1784 GND.n1783 2.2505
R1240 GND.n1782 GND.n1752 2.2505
R1241 GND.n1781 GND.n1780 2.2505
R1242 GND.n1779 GND.n1753 2.2505
R1243 GND.n1778 GND.n1777 2.2505
R1244 GND.n1776 GND.n1754 2.2505
R1245 GND.n1775 GND.n1774 2.2505
R1246 GND.n1773 GND.n1755 2.2505
R1247 GND.n1772 GND.n1771 2.2505
R1248 GND.n1770 GND.n1756 2.2505
R1249 GND.n1769 GND.n1768 2.2505
R1250 GND.n1767 GND.n1757 2.2505
R1251 GND.n1766 GND.n1765 2.2505
R1252 GND.n1764 GND.n1758 2.2505
R1253 GND.n1763 GND.n1762 2.2505
R1254 GND.n1761 GND.n1760 2.2505
R1255 GND.n1759 GND.n1682 2.2505
R1256 GND.n1980 GND.n1681 2.2505
R1257 GND.n1982 GND.n1981 2.2505
R1258 GND.n1983 GND.n1680 2.2505
R1259 GND.n1985 GND.n1984 2.2505
R1260 GND.n1986 GND.n1679 2.2505
R1261 GND.n1988 GND.n1987 2.2505
R1262 GND.n1989 GND.n1678 2.2505
R1263 GND.n1991 GND.n1990 2.2505
R1264 GND.n1992 GND.n1677 2.2505
R1265 GND.n1994 GND.n1993 2.2505
R1266 GND.n1995 GND.n1676 2.2505
R1267 GND.n1997 GND.n1996 2.2505
R1268 GND.n1998 GND.n1675 2.2505
R1269 GND.n2000 GND.n1999 2.2505
R1270 GND.n2001 GND.n1674 2.2505
R1271 GND.n2003 GND.n2002 2.2505
R1272 GND.n2004 GND.n1673 2.2505
R1273 GND.n2006 GND.n2005 2.2505
R1274 GND.n2007 GND.n1672 2.2505
R1275 GND.n2009 GND.n2008 2.2505
R1276 GND.n2010 GND.n1671 2.2505
R1277 GND.n2012 GND.n2011 2.2505
R1278 GND.n2013 GND.n1670 2.2505
R1279 GND.n2015 GND.n2014 2.2505
R1280 GND.n2016 GND.n1669 2.2505
R1281 GND.n2018 GND.n2017 2.2505
R1282 GND.n2019 GND.n1668 2.2505
R1283 GND.n2021 GND.n2020 2.2505
R1284 GND.n2022 GND.n1667 2.2505
R1285 GND.n2024 GND.n2023 2.2505
R1286 GND.n2025 GND.n1666 2.2505
R1287 GND.n2027 GND.n2026 2.2505
R1288 GND.n2028 GND.n1665 2.2505
R1289 GND.n2030 GND.n2029 2.2505
R1290 GND.n2031 GND.n1664 2.2505
R1291 GND.n2033 GND.n2032 2.2505
R1292 GND.n2034 GND.n1663 2.2505
R1293 GND.n2036 GND.n2035 2.2505
R1294 GND.n2037 GND.n1662 2.2505
R1295 GND.n2039 GND.n2038 2.2505
R1296 GND.n2040 GND.n1661 2.2505
R1297 GND.n2042 GND.n2041 2.2505
R1298 GND.n2043 GND.n1660 2.2505
R1299 GND.n2045 GND.n2044 2.2505
R1300 GND.n2046 GND.n1659 2.2505
R1301 GND.n2048 GND.n2047 2.2505
R1302 GND.n2049 GND.n1658 2.2505
R1303 GND.n2051 GND.n2050 2.2505
R1304 GND.n2052 GND.n1657 2.2505
R1305 GND.n2054 GND.n2053 2.2505
R1306 GND.n2055 GND.n1656 2.2505
R1307 GND.n2057 GND.n2056 2.2505
R1308 GND.n2058 GND.n1655 2.2505
R1309 GND.n2060 GND.n2059 2.2505
R1310 GND.n2061 GND.n1654 2.2505
R1311 GND.n2063 GND.n2062 2.2505
R1312 GND.n2064 GND.n1653 2.2505
R1313 GND.n2066 GND.n2065 2.2505
R1314 GND.n2067 GND.n1652 2.2505
R1315 GND.n2069 GND.n2068 2.2505
R1316 GND.n2070 GND.n1651 2.2505
R1317 GND.n2072 GND.n2071 2.2505
R1318 GND.n2073 GND.n1650 2.2505
R1319 GND.n2075 GND.n2074 2.2505
R1320 GND.n2076 GND.n1649 2.2505
R1321 GND.n2078 GND.n2077 2.2505
R1322 GND.n2079 GND.n1648 2.2505
R1323 GND.n2081 GND.n2080 2.2505
R1324 GND.n2082 GND.n1647 2.2505
R1325 GND.n2084 GND.n2083 2.2505
R1326 GND.n2085 GND.n1646 2.2505
R1327 GND.n2087 GND.n2086 2.2505
R1328 GND.n2088 GND.n1645 2.2505
R1329 GND.n2090 GND.n2089 2.2505
R1330 GND.n2091 GND.n1644 2.2505
R1331 GND.n2093 GND.n2092 2.2505
R1332 GND.n2094 GND.n1643 2.2505
R1333 GND.n2096 GND.n2095 2.2505
R1334 GND.n2097 GND.n1642 2.2505
R1335 GND.n2099 GND.n2098 2.2505
R1336 GND.n2100 GND.n1641 2.2505
R1337 GND.n2102 GND.n2101 2.2505
R1338 GND.n2103 GND.n1640 2.2505
R1339 GND.n2105 GND.n2104 2.2505
R1340 GND.n2106 GND.n1639 2.2505
R1341 GND.n2108 GND.n2107 2.2505
R1342 GND.n2109 GND.n1638 2.2505
R1343 GND.n2111 GND.n2110 2.2505
R1344 GND.n2112 GND.n1637 2.2505
R1345 GND.n2114 GND.n2113 2.2505
R1346 GND.n2115 GND.n1636 2.2505
R1347 GND.n2117 GND.n2116 2.2505
R1348 GND.n2118 GND.n1635 2.2505
R1349 GND.n2120 GND.n2119 2.2505
R1350 GND.n2121 GND.n1634 2.2505
R1351 GND.n2123 GND.n2122 2.2505
R1352 GND.n2124 GND.n1633 2.2505
R1353 GND.n2126 GND.n2125 2.2505
R1354 GND.n2127 GND.n1632 2.2505
R1355 GND.n2129 GND.n2128 2.2505
R1356 GND.n2130 GND.n1631 2.2505
R1357 GND.n2132 GND.n2131 2.2505
R1358 GND.n2133 GND.n1630 2.2505
R1359 GND.n2135 GND.n2134 2.2505
R1360 GND.n2136 GND.n1629 2.2505
R1361 GND.n2138 GND.n2137 2.2505
R1362 GND.n2139 GND.n1628 2.2505
R1363 GND.n2141 GND.n2140 2.2505
R1364 GND.n2142 GND.n1627 2.2505
R1365 GND.n2144 GND.n2143 2.2505
R1366 GND.n2145 GND.n1626 2.2505
R1367 GND.n2147 GND.n2146 2.2505
R1368 GND.n2148 GND.n1625 2.2505
R1369 GND.n2150 GND.n2149 2.2505
R1370 GND.n2151 GND.n1624 2.2505
R1371 GND.n2153 GND.n2152 2.2505
R1372 GND.n2154 GND.n1623 2.2505
R1373 GND.n2156 GND.n2155 2.2505
R1374 GND.n2157 GND.n1622 2.2505
R1375 GND.n2159 GND.n2158 2.2505
R1376 GND.n2162 GND.n2161 2.2505
R1377 GND.n2163 GND.n1620 2.2505
R1378 GND.n2165 GND.n2164 2.2505
R1379 GND.n2166 GND.n1619 2.2505
R1380 GND.n2168 GND.n2167 2.2505
R1381 GND.n2169 GND.n1618 2.2505
R1382 GND.n2171 GND.n2170 2.2505
R1383 GND.n2172 GND.n1617 2.2505
R1384 GND.n2174 GND.n2173 2.2505
R1385 GND.n2175 GND.n1616 2.2505
R1386 GND.n2177 GND.n2176 2.2505
R1387 GND.n2178 GND.n1615 2.2505
R1388 GND.n2180 GND.n2179 2.2505
R1389 GND.n2181 GND.n1614 2.2505
R1390 GND.n2183 GND.n2182 2.2505
R1391 GND.n2184 GND.n1613 2.2505
R1392 GND.n2186 GND.n2185 2.2505
R1393 GND.n2187 GND.n1612 2.2505
R1394 GND.n2189 GND.n2188 2.2505
R1395 GND.n2190 GND.n1611 2.2505
R1396 GND.n2192 GND.n2191 2.2505
R1397 GND.n2193 GND.n1610 2.2505
R1398 GND.n2195 GND.n2194 2.2505
R1399 GND.n2196 GND.n1609 2.2505
R1400 GND.n2198 GND.n2197 2.2505
R1401 GND.n2199 GND.n1608 2.2505
R1402 GND.n2201 GND.n2200 2.2505
R1403 GND.n2202 GND.n1607 2.2505
R1404 GND.n2204 GND.n2203 2.2505
R1405 GND.n2205 GND.n1606 2.2505
R1406 GND.n2207 GND.n2206 2.2505
R1407 GND.n2208 GND.n1605 2.2505
R1408 GND.n2210 GND.n2209 2.2505
R1409 GND.n2211 GND.n1604 2.2505
R1410 GND.n2213 GND.n2212 2.2505
R1411 GND.n2214 GND.n1603 2.2505
R1412 GND.n2216 GND.n2215 2.2505
R1413 GND.n2217 GND.n1602 2.2505
R1414 GND.n2219 GND.n2218 2.2505
R1415 GND.n2220 GND.n1601 2.2505
R1416 GND.n2222 GND.n2221 2.2505
R1417 GND.n2223 GND.n1600 2.2505
R1418 GND.n2225 GND.n2224 2.2505
R1419 GND.n2226 GND.n1599 2.2505
R1420 GND.n2228 GND.n2227 2.2505
R1421 GND.n2229 GND.n1598 2.2505
R1422 GND.n2231 GND.n2230 2.2505
R1423 GND.n2232 GND.n1597 2.2505
R1424 GND.n2234 GND.n2233 2.2505
R1425 GND.n2235 GND.n1596 2.2505
R1426 GND.n2237 GND.n2236 2.2505
R1427 GND.n2238 GND.n1595 2.2505
R1428 GND.n2240 GND.n2239 2.2505
R1429 GND.n2241 GND.n1594 2.2505
R1430 GND.n2243 GND.n2242 2.2505
R1431 GND.n2244 GND.n1593 2.2505
R1432 GND.n2246 GND.n2245 2.2505
R1433 GND.n2247 GND.n1592 2.2505
R1434 GND.n2249 GND.n2248 2.2505
R1435 GND.n2250 GND.n1591 2.2505
R1436 GND.n2252 GND.n2251 2.2505
R1437 GND.n2253 GND.n1590 2.2505
R1438 GND.n2255 GND.n2254 2.2505
R1439 GND.n2256 GND.n1589 2.2505
R1440 GND.n2258 GND.n2257 2.2505
R1441 GND.n2259 GND.n1588 2.2505
R1442 GND.n2261 GND.n2260 2.2505
R1443 GND.n2262 GND.n1587 2.2505
R1444 GND.n2264 GND.n2263 2.2505
R1445 GND.n2265 GND.n1586 2.2505
R1446 GND.n2267 GND.n2266 2.2505
R1447 GND.n2268 GND.n1585 2.2505
R1448 GND.n2270 GND.n2269 2.2505
R1449 GND.n2271 GND.n1584 2.2505
R1450 GND.n2273 GND.n2272 2.2505
R1451 GND.n2274 GND.n1583 2.2505
R1452 GND.n2276 GND.n2275 2.2505
R1453 GND.n2277 GND.n1582 2.2505
R1454 GND.n2279 GND.n2278 2.2505
R1455 GND.n2280 GND.n1581 2.2505
R1456 GND.n2282 GND.n2281 2.2505
R1457 GND.n2283 GND.n1580 2.2505
R1458 GND.n2285 GND.n2284 2.2505
R1459 GND.n2286 GND.n1579 2.2505
R1460 GND.n2288 GND.n2287 2.2505
R1461 GND.n2289 GND.n1578 2.2505
R1462 GND.n2291 GND.n2290 2.2505
R1463 GND.n2292 GND.n1577 2.2505
R1464 GND.n2294 GND.n2293 2.2505
R1465 GND.n2295 GND.n1576 2.2505
R1466 GND.n2297 GND.n2296 2.2505
R1467 GND.n2298 GND.n1575 2.2505
R1468 GND.n2300 GND.n2299 2.2505
R1469 GND.n2301 GND.n1574 2.2505
R1470 GND.n2303 GND.n2302 2.2505
R1471 GND.n2304 GND.n1573 2.2505
R1472 GND.n2306 GND.n2305 2.2505
R1473 GND.n2307 GND.n1572 2.2505
R1474 GND.n2309 GND.n2308 2.2505
R1475 GND.n2310 GND.n1571 2.2505
R1476 GND.n2312 GND.n2311 2.2505
R1477 GND.n2313 GND.n1570 2.2505
R1478 GND.n2315 GND.n2314 2.2505
R1479 GND.n2316 GND.n1569 2.2505
R1480 GND.n2318 GND.n2317 2.2505
R1481 GND.n2319 GND.n1568 2.2505
R1482 GND.n2321 GND.n2320 2.2505
R1483 GND.n2322 GND.n1567 2.2505
R1484 GND.n2324 GND.n2323 2.2505
R1485 GND.n2325 GND.n1566 2.2505
R1486 GND.n2327 GND.n2326 2.2505
R1487 GND.n2328 GND.n1565 2.2505
R1488 GND.n2330 GND.n2329 2.2505
R1489 GND.n2331 GND.n1564 2.2505
R1490 GND.n2333 GND.n2332 2.2505
R1491 GND.n2334 GND.n1563 2.2505
R1492 GND.n2336 GND.n2335 2.2505
R1493 GND.n2337 GND.n1562 2.2505
R1494 GND.n2339 GND.n2338 2.2505
R1495 GND.n2340 GND.n1561 2.2505
R1496 GND.n2342 GND.n2341 2.2505
R1497 GND.n2343 GND.n1560 2.2505
R1498 GND.n2345 GND.n2344 2.2505
R1499 GND.n2346 GND.n1559 2.2505
R1500 GND.n2348 GND.n2347 2.2505
R1501 GND.n2349 GND.n1558 2.2505
R1502 GND.n2351 GND.n2350 2.2505
R1503 GND.n2352 GND.n1557 2.2505
R1504 GND.n2354 GND.n2353 2.2505
R1505 GND.n2355 GND.n1556 2.2505
R1506 GND.n2357 GND.n2356 2.2505
R1507 GND.n2358 GND.n1555 2.2505
R1508 GND.n2360 GND.n2359 2.2505
R1509 GND.n2361 GND.n1554 2.2505
R1510 GND.n2363 GND.n2362 2.2505
R1511 GND.n2364 GND.n1553 2.2505
R1512 GND.n2366 GND.n2365 2.2505
R1513 GND.n2367 GND.n1552 2.2505
R1514 GND.n2369 GND.n2368 2.2505
R1515 GND.n2370 GND.n1551 2.2505
R1516 GND.n2372 GND.n2371 2.2505
R1517 GND.n2373 GND.n1550 2.2505
R1518 GND.n2375 GND.n2374 2.2505
R1519 GND.n2376 GND.n1549 2.2505
R1520 GND.n2378 GND.n2377 2.2505
R1521 GND.n2379 GND.n1548 2.2505
R1522 GND.n2381 GND.n2380 2.2505
R1523 GND.n2382 GND.n1547 2.2505
R1524 GND.n2384 GND.n2383 2.2505
R1525 GND.n2385 GND.n1546 2.2505
R1526 GND.n2387 GND.n2386 2.2505
R1527 GND.n2388 GND.n1545 2.2505
R1528 GND.n2390 GND.n2389 2.2505
R1529 GND.n2391 GND.n1544 2.2505
R1530 GND.n2393 GND.n2392 2.2505
R1531 GND.n2394 GND.n1543 2.2505
R1532 GND.n2396 GND.n2395 2.2505
R1533 GND.n2397 GND.n1542 2.2505
R1534 GND.n2399 GND.n2398 2.2505
R1535 GND.n2400 GND.n1541 2.2505
R1536 GND.n2402 GND.n2401 2.2505
R1537 GND.n2403 GND.n1540 2.2505
R1538 GND.n2405 GND.n2404 2.2505
R1539 GND.n2406 GND.n1539 2.2505
R1540 GND.n2408 GND.n2407 2.2505
R1541 GND.n2409 GND.n1538 2.2505
R1542 GND.n2411 GND.n2410 2.2505
R1543 GND.n2412 GND.n1537 2.2505
R1544 GND.n2414 GND.n2413 2.2505
R1545 GND.n2415 GND.n1536 2.2505
R1546 GND.n2417 GND.n2416 2.2505
R1547 GND.n2418 GND.n1535 2.2505
R1548 GND.n2420 GND.n2419 2.2505
R1549 GND.n2421 GND.n1534 2.2505
R1550 GND.n2423 GND.n2422 2.2505
R1551 GND.n2424 GND.n1533 2.2505
R1552 GND.n2426 GND.n2425 2.2505
R1553 GND.n2427 GND.n1532 2.2505
R1554 GND.n2429 GND.n2428 2.2505
R1555 GND.n2430 GND.n1531 2.2505
R1556 GND.n2432 GND.n2431 2.2505
R1557 GND.n2433 GND.n1530 2.2505
R1558 GND.n2435 GND.n2434 2.2505
R1559 GND.n2436 GND.n1529 2.2505
R1560 GND.n2438 GND.n2437 2.2505
R1561 GND.n2439 GND.n1528 2.2505
R1562 GND.n2441 GND.n2440 2.2505
R1563 GND.n2442 GND.n1527 2.2505
R1564 GND.n2444 GND.n2443 2.2505
R1565 GND.n2445 GND.n1526 2.2505
R1566 GND.n2447 GND.n2446 2.2505
R1567 GND.n2448 GND.n1525 2.2505
R1568 GND.n2450 GND.n2449 2.2505
R1569 GND.n2451 GND.n1524 2.2505
R1570 GND.n2453 GND.n2452 2.2505
R1571 GND.n2454 GND.n1523 2.2505
R1572 GND.n2456 GND.n2455 2.2505
R1573 GND.n2457 GND.n1522 2.2505
R1574 GND.n2459 GND.n2458 2.2505
R1575 GND.n2460 GND.n1521 2.2505
R1576 GND.n2462 GND.n2461 2.2505
R1577 GND.n2463 GND.n1520 2.2505
R1578 GND.n2465 GND.n2464 2.2505
R1579 GND.n2466 GND.n1519 2.2505
R1580 GND.n2468 GND.n2467 2.2505
R1581 GND.n2469 GND.n1518 2.2505
R1582 GND.n2471 GND.n2470 2.2505
R1583 GND.n2472 GND.n1517 2.2505
R1584 GND.n2474 GND.n2473 2.2505
R1585 GND.n2475 GND.n1516 2.2505
R1586 GND.n2477 GND.n2476 2.2505
R1587 GND.n2478 GND.n1515 2.2505
R1588 GND.n2480 GND.n2479 2.2505
R1589 GND.n2481 GND.n1514 2.2505
R1590 GND.n2483 GND.n2482 2.2505
R1591 GND.n2484 GND.n1513 2.2505
R1592 GND.n2486 GND.n2485 2.2505
R1593 GND.n2487 GND.n1512 2.2505
R1594 GND.n2489 GND.n2488 2.2505
R1595 GND.n2490 GND.n1511 2.2505
R1596 GND.n2492 GND.n2491 2.2505
R1597 GND.n2493 GND.n1510 2.2505
R1598 GND.n2495 GND.n2494 2.2505
R1599 GND.n2496 GND.n1509 2.2505
R1600 GND.n2498 GND.n2497 2.2505
R1601 GND.n2771 GND.n2770 2.2505
R1602 GND.n2772 GND.n2738 2.2505
R1603 GND.n2774 GND.n2773 2.2505
R1604 GND.n2775 GND.n2737 2.2505
R1605 GND.n2777 GND.n2776 2.2505
R1606 GND.n2778 GND.n2736 2.2505
R1607 GND.n2780 GND.n2779 2.2505
R1608 GND.n2781 GND.n2735 2.2505
R1609 GND.n2783 GND.n2782 2.2505
R1610 GND.n2784 GND.n2734 2.2505
R1611 GND.n2786 GND.n2785 2.2505
R1612 GND.n2787 GND.n2733 2.2505
R1613 GND.n2789 GND.n2788 2.2505
R1614 GND.n2790 GND.n2732 2.2505
R1615 GND.n2792 GND.n2791 2.2505
R1616 GND.n2793 GND.n2731 2.2505
R1617 GND.n2795 GND.n2794 2.2505
R1618 GND.n2796 GND.n2730 2.2505
R1619 GND.n2798 GND.n2797 2.2505
R1620 GND.n2799 GND.n2729 2.2505
R1621 GND.n2801 GND.n2800 2.2505
R1622 GND.n2802 GND.n2728 2.2505
R1623 GND.n2804 GND.n2803 2.2505
R1624 GND.n2805 GND.n2727 2.2505
R1625 GND.n2807 GND.n2806 2.2505
R1626 GND.n2808 GND.n2726 2.2505
R1627 GND.n2810 GND.n2809 2.2505
R1628 GND.n2811 GND.n2725 2.2505
R1629 GND.n2813 GND.n2812 2.2505
R1630 GND.n2814 GND.n2724 2.2505
R1631 GND.n2816 GND.n2815 2.2505
R1632 GND.n2817 GND.n2723 2.2505
R1633 GND.n2819 GND.n2818 2.2505
R1634 GND.n2820 GND.n2722 2.2505
R1635 GND.n2822 GND.n2821 2.2505
R1636 GND.n2823 GND.n2721 2.2505
R1637 GND.n2825 GND.n2824 2.2505
R1638 GND.n2826 GND.n2720 2.2505
R1639 GND.n2828 GND.n2827 2.2505
R1640 GND.n2829 GND.n2719 2.2505
R1641 GND.n2831 GND.n2830 2.2505
R1642 GND.n2832 GND.n2718 2.2505
R1643 GND.n2834 GND.n2833 2.2505
R1644 GND.n2835 GND.n2717 2.2505
R1645 GND.n2837 GND.n2836 2.2505
R1646 GND.n2838 GND.n2716 2.2505
R1647 GND.n2840 GND.n2839 2.2505
R1648 GND.n2841 GND.n2715 2.2505
R1649 GND.n2843 GND.n2842 2.2505
R1650 GND.n2844 GND.n2714 2.2505
R1651 GND.n2846 GND.n2845 2.2505
R1652 GND.n2847 GND.n2713 2.2505
R1653 GND.n2849 GND.n2848 2.2505
R1654 GND.n2850 GND.n2712 2.2505
R1655 GND.n2852 GND.n2851 2.2505
R1656 GND.n2853 GND.n2711 2.2505
R1657 GND.n2855 GND.n2854 2.2505
R1658 GND.n2856 GND.n2710 2.2505
R1659 GND.n2858 GND.n2857 2.2505
R1660 GND.n2859 GND.n2709 2.2505
R1661 GND.n2861 GND.n2860 2.2505
R1662 GND.n2862 GND.n2708 2.2505
R1663 GND.n2864 GND.n2863 2.2505
R1664 GND.n2865 GND.n2707 2.2505
R1665 GND.n2867 GND.n2866 2.2505
R1666 GND.n2868 GND.n2706 2.2505
R1667 GND.n2870 GND.n2869 2.2505
R1668 GND.n2871 GND.n2705 2.2505
R1669 GND.n2873 GND.n2872 2.2505
R1670 GND.n2874 GND.n2704 2.2505
R1671 GND.n2876 GND.n2875 2.2505
R1672 GND.n2877 GND.n2703 2.2505
R1673 GND.n2879 GND.n2878 2.2505
R1674 GND.n2880 GND.n2702 2.2505
R1675 GND.n2882 GND.n2881 2.2505
R1676 GND.n2883 GND.n2701 2.2505
R1677 GND.n2885 GND.n2884 2.2505
R1678 GND.n2886 GND.n2700 2.2505
R1679 GND.n2888 GND.n2887 2.2505
R1680 GND.n2889 GND.n2699 2.2505
R1681 GND.n2891 GND.n2890 2.2505
R1682 GND.n2892 GND.n2698 2.2505
R1683 GND.n2894 GND.n2893 2.2505
R1684 GND.n2895 GND.n2697 2.2505
R1685 GND.n2897 GND.n2896 2.2505
R1686 GND.n2898 GND.n2696 2.2505
R1687 GND.n2900 GND.n2899 2.2505
R1688 GND.n2901 GND.n2695 2.2505
R1689 GND.n2903 GND.n2902 2.2505
R1690 GND.n2904 GND.n2694 2.2505
R1691 GND.n2906 GND.n2905 2.2505
R1692 GND.n2907 GND.n2693 2.2505
R1693 GND.n2909 GND.n2908 2.2505
R1694 GND.n2910 GND.n2692 2.2505
R1695 GND.n2912 GND.n2911 2.2505
R1696 GND.n2913 GND.n2691 2.2505
R1697 GND.n2915 GND.n2914 2.2505
R1698 GND.n2916 GND.n2690 2.2505
R1699 GND.n2918 GND.n2917 2.2505
R1700 GND.n2919 GND.n2689 2.2505
R1701 GND.n2921 GND.n2920 2.2505
R1702 GND.n2922 GND.n2688 2.2505
R1703 GND.n2924 GND.n2923 2.2505
R1704 GND.n2925 GND.n2687 2.2505
R1705 GND.n2927 GND.n2926 2.2505
R1706 GND.n2928 GND.n2686 2.2505
R1707 GND.n2930 GND.n2929 2.2505
R1708 GND.n2931 GND.n2685 2.2505
R1709 GND.n2933 GND.n2932 2.2505
R1710 GND.n2934 GND.n2684 2.2505
R1711 GND.n2936 GND.n2935 2.2505
R1712 GND.n2937 GND.n2683 2.2505
R1713 GND.n2939 GND.n2938 2.2505
R1714 GND.n2940 GND.n2682 2.2505
R1715 GND.n2942 GND.n2941 2.2505
R1716 GND.n2943 GND.n2681 2.2505
R1717 GND.n2945 GND.n2944 2.2505
R1718 GND.n2946 GND.n2680 2.2505
R1719 GND.n2948 GND.n2947 2.2505
R1720 GND.n2949 GND.n1448 2.2505
R1721 GND.n2951 GND.n2950 2.2505
R1722 GND.n2679 GND.n1447 2.2505
R1723 GND.n2678 GND.n2677 2.2505
R1724 GND.n2676 GND.n1449 2.2505
R1725 GND.n2675 GND.n2674 2.2505
R1726 GND.n2673 GND.n1450 2.2505
R1727 GND.n2672 GND.n2671 2.2505
R1728 GND.n2670 GND.n1451 2.2505
R1729 GND.n2669 GND.n2668 2.2505
R1730 GND.n2667 GND.n1452 2.2505
R1731 GND.n2666 GND.n2665 2.2505
R1732 GND.n2664 GND.n1453 2.2505
R1733 GND.n2663 GND.n2662 2.2505
R1734 GND.n2661 GND.n1454 2.2505
R1735 GND.n2660 GND.n2659 2.2505
R1736 GND.n2658 GND.n1455 2.2505
R1737 GND.n2657 GND.n2656 2.2505
R1738 GND.n2655 GND.n1456 2.2505
R1739 GND.n2654 GND.n2653 2.2505
R1740 GND.n2652 GND.n1457 2.2505
R1741 GND.n2651 GND.n2650 2.2505
R1742 GND.n2649 GND.n1458 2.2505
R1743 GND.n2648 GND.n2647 2.2505
R1744 GND.n2646 GND.n1459 2.2505
R1745 GND.n2645 GND.n2644 2.2505
R1746 GND.n2643 GND.n1460 2.2505
R1747 GND.n2642 GND.n2641 2.2505
R1748 GND.n2640 GND.n1461 2.2505
R1749 GND.n2639 GND.n2638 2.2505
R1750 GND.n2637 GND.n1462 2.2505
R1751 GND.n2636 GND.n2635 2.2505
R1752 GND.n2634 GND.n1463 2.2505
R1753 GND.n2633 GND.n2632 2.2505
R1754 GND.n2631 GND.n1464 2.2505
R1755 GND.n2630 GND.n2629 2.2505
R1756 GND.n2628 GND.n1465 2.2505
R1757 GND.n2627 GND.n2626 2.2505
R1758 GND.n2625 GND.n1466 2.2505
R1759 GND.n2624 GND.n2623 2.2505
R1760 GND.n2622 GND.n1467 2.2505
R1761 GND.n2621 GND.n2620 2.2505
R1762 GND.n2619 GND.n1468 2.2505
R1763 GND.n2618 GND.n2617 2.2505
R1764 GND.n2616 GND.n1469 2.2505
R1765 GND.n2615 GND.n2614 2.2505
R1766 GND.n2613 GND.n1470 2.2505
R1767 GND.n2612 GND.n2611 2.2505
R1768 GND.n2610 GND.n1471 2.2505
R1769 GND.n2609 GND.n2608 2.2505
R1770 GND.n2607 GND.n1472 2.2505
R1771 GND.n2606 GND.n2605 2.2505
R1772 GND.n2604 GND.n1473 2.2505
R1773 GND.n2603 GND.n2602 2.2505
R1774 GND.n2601 GND.n1474 2.2505
R1775 GND.n2600 GND.n2599 2.2505
R1776 GND.n2598 GND.n1475 2.2505
R1777 GND.n2597 GND.n2596 2.2505
R1778 GND.n2595 GND.n1476 2.2505
R1779 GND.n2594 GND.n2593 2.2505
R1780 GND.n2592 GND.n1477 2.2505
R1781 GND.n2591 GND.n2590 2.2505
R1782 GND.n2589 GND.n1478 2.2505
R1783 GND.n2588 GND.n2587 2.2505
R1784 GND.n2586 GND.n1479 2.2505
R1785 GND.n2585 GND.n2584 2.2505
R1786 GND.n2583 GND.n1480 2.2505
R1787 GND.n2582 GND.n2581 2.2505
R1788 GND.n2580 GND.n1481 2.2505
R1789 GND.n2579 GND.n2578 2.2505
R1790 GND.n2577 GND.n1482 2.2505
R1791 GND.n2576 GND.n2575 2.2505
R1792 GND.n2574 GND.n1483 2.2505
R1793 GND.n2573 GND.n2572 2.2505
R1794 GND.n2571 GND.n1484 2.2505
R1795 GND.n2570 GND.n2569 2.2505
R1796 GND.n2568 GND.n1485 2.2505
R1797 GND.n2567 GND.n2566 2.2505
R1798 GND.n2565 GND.n1486 2.2505
R1799 GND.n2564 GND.n2563 2.2505
R1800 GND.n2562 GND.n1487 2.2505
R1801 GND.n2561 GND.n2560 2.2505
R1802 GND.n2559 GND.n1488 2.2505
R1803 GND.n2558 GND.n2557 2.2505
R1804 GND.n2556 GND.n1489 2.2505
R1805 GND.n2555 GND.n2554 2.2505
R1806 GND.n2553 GND.n1490 2.2505
R1807 GND.n2552 GND.n2551 2.2505
R1808 GND.n2550 GND.n1491 2.2505
R1809 GND.n2549 GND.n2548 2.2505
R1810 GND.n2547 GND.n1492 2.2505
R1811 GND.n2546 GND.n2545 2.2505
R1812 GND.n2544 GND.n1493 2.2505
R1813 GND.n2543 GND.n2542 2.2505
R1814 GND.n2541 GND.n1494 2.2505
R1815 GND.n2540 GND.n2539 2.2505
R1816 GND.n2538 GND.n1495 2.2505
R1817 GND.n2537 GND.n2536 2.2505
R1818 GND.n2535 GND.n1496 2.2505
R1819 GND.n2534 GND.n2533 2.2505
R1820 GND.n2532 GND.n1497 2.2505
R1821 GND.n2531 GND.n2530 2.2505
R1822 GND.n2529 GND.n1498 2.2505
R1823 GND.n2528 GND.n2527 2.2505
R1824 GND.n2526 GND.n1499 2.2505
R1825 GND.n2525 GND.n2524 2.2505
R1826 GND.n2523 GND.n1500 2.2505
R1827 GND.n2522 GND.n2521 2.2505
R1828 GND.n2520 GND.n1501 2.2505
R1829 GND.n2519 GND.n2518 2.2505
R1830 GND.n2517 GND.n1502 2.2505
R1831 GND.n2516 GND.n2515 2.2505
R1832 GND.n2514 GND.n1503 2.2505
R1833 GND.n2513 GND.n2512 2.2505
R1834 GND.n2511 GND.n1504 2.2505
R1835 GND.n2510 GND.n2509 2.2505
R1836 GND.n2508 GND.n1505 2.2505
R1837 GND.n2507 GND.n2506 2.2505
R1838 GND.n2505 GND.n1506 2.2505
R1839 GND.n2504 GND.n2503 2.2505
R1840 GND.n2502 GND.n1507 2.2505
R1841 GND.n2501 GND.n2500 2.2505
R1842 GND.n2769 GND.n2739 2.2505
R1843 GND.n1974 GND.n1688 2.2505
R1844 GND.n1973 GND.n1972 2.2505
R1845 GND.n1971 GND.n1689 2.2505
R1846 GND.n1970 GND.n1969 2.2505
R1847 GND.n1968 GND.n1690 2.2505
R1848 GND.n1967 GND.n1966 2.2505
R1849 GND.n1965 GND.n1691 2.2505
R1850 GND.n1964 GND.n1963 2.2505
R1851 GND.n1962 GND.n1692 2.2505
R1852 GND.n1961 GND.n1960 2.2505
R1853 GND.n1959 GND.n1693 2.2505
R1854 GND.n1958 GND.n1957 2.2505
R1855 GND.n1956 GND.n1694 2.2505
R1856 GND.n1955 GND.n1954 2.2505
R1857 GND.n1953 GND.n1695 2.2505
R1858 GND.n1952 GND.n1951 2.2505
R1859 GND.n1950 GND.n1696 2.2505
R1860 GND.n1949 GND.n1948 2.2505
R1861 GND.n1947 GND.n1697 2.2505
R1862 GND.n1946 GND.n1945 2.2505
R1863 GND.n1944 GND.n1698 2.2505
R1864 GND.n1943 GND.n1942 2.2505
R1865 GND.n1941 GND.n1699 2.2505
R1866 GND.n3023 GND.n1417 2.2505
R1867 GND.n3022 GND.n3021 2.2505
R1868 GND.n3020 GND.n1421 2.2505
R1869 GND.n3019 GND.n3018 2.2505
R1870 GND.n3017 GND.n1422 2.2505
R1871 GND.n3016 GND.n3015 2.2505
R1872 GND.n3014 GND.n1423 2.2505
R1873 GND.n3013 GND.n3012 2.2505
R1874 GND.n3011 GND.n1424 2.2505
R1875 GND.n3010 GND.n3009 2.2505
R1876 GND.n3008 GND.n1425 2.2505
R1877 GND.n3007 GND.n3006 2.2505
R1878 GND.n3005 GND.n1426 2.2505
R1879 GND.n3004 GND.n3003 2.2505
R1880 GND.n3002 GND.n1427 2.2505
R1881 GND.n3001 GND.n3000 2.2505
R1882 GND.n2999 GND.n1428 2.2505
R1883 GND.n2998 GND.n2997 2.2505
R1884 GND.n2996 GND.n1429 2.2505
R1885 GND.n2995 GND.n2994 2.2505
R1886 GND.n2993 GND.n1430 2.2505
R1887 GND.n2992 GND.n2991 2.2505
R1888 GND.n2990 GND.n1431 2.2505
R1889 GND.n2989 GND.n2988 2.2505
R1890 GND.n2987 GND.n1432 2.2505
R1891 GND.n2986 GND.n2985 2.2505
R1892 GND.n2984 GND.n1433 2.2505
R1893 GND.n2983 GND.n2982 2.2505
R1894 GND.n2981 GND.n1434 2.2505
R1895 GND.n2980 GND.n2979 2.2505
R1896 GND.n2978 GND.n1435 2.2505
R1897 GND.n2977 GND.n2976 2.2505
R1898 GND.n2975 GND.n1436 2.2505
R1899 GND.n2974 GND.n2973 2.2505
R1900 GND.n2972 GND.n1437 2.2505
R1901 GND.n2971 GND.n2970 2.2505
R1902 GND.n2969 GND.n1438 2.2505
R1903 GND.n2968 GND.n2967 2.2505
R1904 GND.n2966 GND.n1439 2.2505
R1905 GND.n2965 GND.n2964 2.2505
R1906 GND.n2963 GND.n1440 2.2505
R1907 GND.n2962 GND.n2961 2.2505
R1908 GND.n2960 GND.n1441 2.2505
R1909 GND.n2959 GND.n2958 2.2505
R1910 GND.n2957 GND.n1442 2.2505
R1911 GND.n2767 GND.n2766 2.2505
R1912 GND.n2765 GND.n2741 2.2505
R1913 GND.n2764 GND.n2763 2.2505
R1914 GND.n2762 GND.n2742 2.2505
R1915 GND.n2761 GND.n2760 2.2505
R1916 GND.n2759 GND.n2743 2.2505
R1917 GND.n2758 GND.n2757 2.2505
R1918 GND.n2756 GND.n2744 2.2505
R1919 GND.n2755 GND.n2754 2.2505
R1920 GND.n2753 GND.n2745 2.2505
R1921 GND.n2752 GND.n2751 2.2505
R1922 GND.n2750 GND.n2746 2.2505
R1923 GND.n2749 GND.n2748 2.2505
R1924 GND.n2747 GND.n1418 2.2505
R1925 GND.n496 GND.n495 2.24636
R1926 GND.n491 GND.n452 2.24636
R1927 GND.n492 GND.n490 2.24405
R1928 GND.n3027 GND.n1416 2.24111
R1929 GND.n3025 GND.n1420 2.24111
R1930 GND.n3027 GND.n1415 2.24111
R1931 GND.n45 GND.t45 1.69686
R1932 GND.n31 GND.t240 1.69376
R1933 GND.n33 GND.t291 1.69376
R1934 GND.n1319 GND.t200 1.681
R1935 GND.n1357 GND.t270 1.681
R1936 GND.n36 GND.t184 1.681
R1937 GND.n338 GND.t307 1.6805
R1938 GND.n338 GND.t264 1.6805
R1939 GND.n47 GND.t59 1.6805
R1940 GND.n47 GND.t323 1.6805
R1941 GND.n48 GND.t110 1.6805
R1942 GND.n48 GND.t51 1.6805
R1943 GND.n49 GND.t317 1.6805
R1944 GND.n1302 GND.t87 1.6805
R1945 GND.n1302 GND.t108 1.6805
R1946 GND.n56 GND.t159 1.6805
R1947 GND.n56 GND.t182 1.6805
R1948 GND.n57 GND.t213 1.6805
R1949 GND.n58 GND.t138 1.6805
R1950 GND.n59 GND.t202 1.6805
R1951 GND.n60 GND.t215 1.6805
R1952 GND.n61 GND.t186 1.6805
R1953 GND.n62 GND.t82 1.6805
R1954 GND.n63 GND.t313 1.6805
R1955 GND.n63 GND.t129 1.6805
R1956 GND.n64 GND.t283 1.6805
R1957 GND.n64 GND.t74 1.6805
R1958 GND.n22 GND.t281 1.6805
R1959 GND.n22 GND.t127 1.6805
R1960 GND.n1376 GND.t219 1.6805
R1961 GND.n1376 GND.t71 1.6805
R1962 GND.n28 GND.t299 1.6805
R1963 GND.n27 GND.t244 1.6805
R1964 GND.n26 GND.t295 1.6805
R1965 GND.n25 GND.t113 1.6805
R1966 GND.n24 GND.t285 1.6805
R1967 GND.n23 GND.t226 1.6805
R1968 GND.n35 GND.t125 1.6805
R1969 GND.n35 GND.t123 1.6805
R1970 GND.n35 GND.t277 1.6805
R1971 GND.n34 GND.t168 1.6805
R1972 GND.n34 GND.t166 1.6805
R1973 GND.n34 GND.t301 1.6805
R1974 GND.n30 GND.t217 1.6805
R1975 GND.n30 GND.t211 1.6805
R1976 GND.n30 GND.t321 1.6805
R1977 GND.n38 GND.t39 1.6805
R1978 GND.n41 GND.t297 1.6805
R1979 GND.n41 GND.t157 1.6805
R1980 GND.n40 GND.t53 1.6805
R1981 GND.n40 GND.t48 1.6805
R1982 GND.n39 GND.t94 1.6805
R1983 GND.n39 GND.t92 1.6805
R1984 GND.n1332 GND.t147 1.6805
R1985 GND.n493 GND.n450 1.51495
R1986 GND.n487 GND.n486 1.5005
R1987 GND.n485 GND.n458 1.5005
R1988 GND.n484 GND.n483 1.5005
R1989 GND.n482 GND.n459 1.5005
R1990 GND.n481 GND.n480 1.5005
R1991 GND.n479 GND.n460 1.5005
R1992 GND.n478 GND.n477 1.5005
R1993 GND.n476 GND.n475 1.5005
R1994 GND.n474 GND.n457 1.5005
R1995 GND.n473 GND.n456 1.5005
R1996 GND.n472 GND.n471 1.5005
R1997 GND.n470 GND.n461 1.5005
R1998 GND.n469 GND.n468 1.5005
R1999 GND.n467 GND.n462 1.5005
R2000 GND.n466 GND.n465 1.5005
R2001 GND.n464 GND.n463 1.5005
R2002 GND.n455 GND.n454 1.5005
R2003 GND.n489 GND.n488 1.5005
R2004 GND.n452 GND.n451 1.5005
R2005 GND.n497 GND.n496 1.5005
R2006 GND.n498 GND.n497 1.5005
R2007 GND.n346 GND.n44 1.47371
R2008 GND.n345 GND.n339 1.4646
R2009 GND.n1112 GND.n1106 1.3355
R2010 GND.n1113 GND.n1099 1.3355
R2011 GND.n1114 GND.n1092 1.3355
R2012 GND.n1115 GND.n1085 1.3355
R2013 GND.n1160 GND.n1122 1.3355
R2014 GND.n1159 GND.n1129 1.3355
R2015 GND.n1158 GND.n1136 1.3355
R2016 GND.n1157 GND.n1143 1.3355
R2017 GND.n1156 GND.n1150 1.3355
R2018 GND.n1074 GND.t26 1.2605
R2019 GND.n1074 GND.t437 1.2605
R2020 GND.n1073 GND.t408 1.2605
R2021 GND.n1073 GND.t418 1.2605
R2022 GND.n1975 GND.n1443 1.19266
R2023 GND.n1687 GND.n1443 1.17423
R2024 GND.n378 GND.n377 1.15205
R2025 GND.n368 GND.n322 1.00945
R2026 GND.n371 GND.n322 1.00945
R2027 GND.n366 GND.n363 1.00945
R2028 GND.n1108 GND.n1107 0.926214
R2029 GND.n1109 GND.n1108 0.926214
R2030 GND.n1110 GND.n1109 0.926214
R2031 GND.n1111 GND.n1110 0.926214
R2032 GND.n1101 GND.n1100 0.926214
R2033 GND.n1102 GND.n1101 0.926214
R2034 GND.n1103 GND.n1102 0.926214
R2035 GND.n1104 GND.n1103 0.926214
R2036 GND.n1105 GND.n1104 0.926214
R2037 GND.n1106 GND.n1105 0.926214
R2038 GND.n1094 GND.n1093 0.926214
R2039 GND.n1095 GND.n1094 0.926214
R2040 GND.n1096 GND.n1095 0.926214
R2041 GND.n1097 GND.n1096 0.926214
R2042 GND.n1098 GND.n1097 0.926214
R2043 GND.n1099 GND.n1098 0.926214
R2044 GND.n1087 GND.n1086 0.926214
R2045 GND.n1088 GND.n1087 0.926214
R2046 GND.n1089 GND.n1088 0.926214
R2047 GND.n1090 GND.n1089 0.926214
R2048 GND.n1091 GND.n1090 0.926214
R2049 GND.n1092 GND.n1091 0.926214
R2050 GND.n1079 GND.n1078 0.926214
R2051 GND.n1080 GND.n1079 0.926214
R2052 GND.n1081 GND.n1080 0.926214
R2053 GND.n1082 GND.n1081 0.926214
R2054 GND.n1083 GND.n1082 0.926214
R2055 GND.n1084 GND.n1083 0.926214
R2056 GND.n1085 GND.n1084 0.926214
R2057 GND.n1117 GND.n1116 0.926214
R2058 GND.n1118 GND.n1117 0.926214
R2059 GND.n1119 GND.n1118 0.926214
R2060 GND.n1120 GND.n1119 0.926214
R2061 GND.n1121 GND.n1120 0.926214
R2062 GND.n1122 GND.n1121 0.926214
R2063 GND.n1124 GND.n1123 0.926214
R2064 GND.n1125 GND.n1124 0.926214
R2065 GND.n1126 GND.n1125 0.926214
R2066 GND.n1127 GND.n1126 0.926214
R2067 GND.n1128 GND.n1127 0.926214
R2068 GND.n1129 GND.n1128 0.926214
R2069 GND.n1131 GND.n1130 0.926214
R2070 GND.n1132 GND.n1131 0.926214
R2071 GND.n1133 GND.n1132 0.926214
R2072 GND.n1134 GND.n1133 0.926214
R2073 GND.n1135 GND.n1134 0.926214
R2074 GND.n1136 GND.n1135 0.926214
R2075 GND.n1138 GND.n1137 0.926214
R2076 GND.n1139 GND.n1138 0.926214
R2077 GND.n1140 GND.n1139 0.926214
R2078 GND.n1141 GND.n1140 0.926214
R2079 GND.n1142 GND.n1141 0.926214
R2080 GND.n1143 GND.n1142 0.926214
R2081 GND.n1145 GND.n1144 0.926214
R2082 GND.n1146 GND.n1145 0.926214
R2083 GND.n1147 GND.n1146 0.926214
R2084 GND.n1148 GND.n1147 0.926214
R2085 GND.n1149 GND.n1148 0.926214
R2086 GND.n1150 GND.n1149 0.926214
R2087 GND.n1152 GND.n1151 0.926214
R2088 GND.n1153 GND.n1152 0.926214
R2089 GND.n1154 GND.n1153 0.926214
R2090 GND.n1155 GND.n1154 0.926214
R2091 GND.n1113 GND.n1112 0.9005
R2092 GND.n1114 GND.n1113 0.9005
R2093 GND.n1115 GND.n1114 0.9005
R2094 GND.n1160 GND.n1159 0.9005
R2095 GND.n1159 GND.n1158 0.9005
R2096 GND.n1158 GND.n1157 0.9005
R2097 GND.n1157 GND.n1156 0.9005
R2098 GND.n323 GND.n322 0.867167
R2099 GND.n363 GND.n318 0.867167
R2100 GND.n318 GND.n312 0.867167
R2101 GND.n364 GND.n321 0.867167
R2102 GND.t379 GND.n364 0.867167
R2103 GND.n313 GND.n311 0.826654
R2104 GND.n315 GND.n314 0.826654
R2105 GND.n498 GND.n450 0.7789
R2106 GND.n1977 GND.n1687 0.755
R2107 GND.n369 GND.n368 0.743357
R2108 GND.t394 GND.n369 0.743357
R2109 GND.n371 GND.n370 0.743357
R2110 GND.n370 GND.t394 0.743357
R2111 GND.n366 GND.n365 0.743357
R2112 GND.n374 GND.n373 0.743357
R2113 GND.n375 GND.n374 0.743357
R2114 GND.n1077 GND.n1076 0.634786
R2115 GND.n449 GND.n448 0.600741
R2116 GND.n1161 GND.n1115 0.6005
R2117 GND.n378 GND.n231 0.57754
R2118 GND.n357 GND.n332 0.575504
R2119 GND.n357 GND.n356 0.575504
R2120 GND.n357 GND.n334 0.575504
R2121 GND.n342 GND.n341 0.548
R2122 GND.n348 GND.n347 0.545857
R2123 GND.n373 GND.n372 0.5405
R2124 GND.n372 GND.n371 0.5405
R2125 GND.n367 GND.n366 0.5405
R2126 GND.n368 GND.n367 0.5405
R2127 GND.n363 GND.n320 0.513219
R2128 GND.n341 GND.n337 0.471929
R2129 GND.n354 GND.n337 0.471929
R2130 GND.n354 GND.n353 0.471929
R2131 GND.n353 GND.n352 0.471929
R2132 GND.n352 GND.n350 0.471929
R2133 GND.n350 GND.n348 0.471929
R2134 GND.n367 GND.n321 0.469447
R2135 GND.n372 GND.n321 0.469447
R2136 GND.n254 GND.n194 0.399459
R2137 GND.n423 GND.n194 0.396656
R2138 GND.n3028 GND.n3027 0.363875
R2139 GND.n1161 GND.n1160 0.3005
R2140 GND.n486 GND.t30 0.25547
R2141 GND.n449 GND.n176 0.243441
R2142 GND.n379 GND.n378 0.242328
R2143 GND.n2957 GND.n2956 0.234366
R2144 GND.n1975 GND.n1974 0.229823
R2145 GND.n199 GND.n194 0.220722
R2146 GND.n499 GND.n498 0.2183
R2147 GND.n2956 GND.n2955 0.214495
R2148 GND.n346 GND.n345 0.206158
R2149 GND.n1976 GND.n1975 0.199263
R2150 GND.n314 GND.n313 0.194346
R2151 GND.n377 GND.n311 0.164346
R2152 GND.n502 GND.n1 0.114071
R2153 GND.n503 GND.n502 0.114071
R2154 GND.n503 GND.n175 0.114071
R2155 GND.n507 GND.n175 0.114071
R2156 GND.n508 GND.n507 0.114071
R2157 GND.n509 GND.n508 0.114071
R2158 GND.n509 GND.n173 0.114071
R2159 GND.n513 GND.n173 0.114071
R2160 GND.n514 GND.n513 0.114071
R2161 GND.n515 GND.n514 0.114071
R2162 GND.n515 GND.n171 0.114071
R2163 GND.n519 GND.n171 0.114071
R2164 GND.n520 GND.n519 0.114071
R2165 GND.n521 GND.n520 0.114071
R2166 GND.n521 GND.n169 0.114071
R2167 GND.n525 GND.n169 0.114071
R2168 GND.n526 GND.n525 0.114071
R2169 GND.n527 GND.n526 0.114071
R2170 GND.n527 GND.n167 0.114071
R2171 GND.n531 GND.n167 0.114071
R2172 GND.n532 GND.n531 0.114071
R2173 GND.n533 GND.n532 0.114071
R2174 GND.n533 GND.n165 0.114071
R2175 GND.n537 GND.n165 0.114071
R2176 GND.n538 GND.n537 0.114071
R2177 GND.n539 GND.n538 0.114071
R2178 GND.n539 GND.n163 0.114071
R2179 GND.n543 GND.n163 0.114071
R2180 GND.n544 GND.n543 0.114071
R2181 GND.n545 GND.n544 0.114071
R2182 GND.n545 GND.n161 0.114071
R2183 GND.n549 GND.n161 0.114071
R2184 GND.n550 GND.n549 0.114071
R2185 GND.n561 GND.n550 0.114071
R2186 GND.n561 GND.n560 0.114071
R2187 GND.n560 GND.n558 0.114071
R2188 GND.n558 GND.n556 0.114071
R2189 GND.n556 GND.n554 0.114071
R2190 GND.n554 GND.n552 0.114071
R2191 GND.n552 GND.n151 0.114071
R2192 GND.n585 GND.n151 0.114071
R2193 GND.n586 GND.n585 0.114071
R2194 GND.n586 GND.n144 0.114071
R2195 GND.n598 GND.n144 0.114071
R2196 GND.n599 GND.n598 0.114071
R2197 GND.n599 GND.n139 0.114071
R2198 GND.n607 GND.n139 0.114071
R2199 GND.n608 GND.n607 0.114071
R2200 GND.n609 GND.n608 0.114071
R2201 GND.n609 GND.n129 0.114071
R2202 GND.n622 GND.n129 0.114071
R2203 GND.n623 GND.n622 0.114071
R2204 GND.n644 GND.n623 0.114071
R2205 GND.n644 GND.n643 0.114071
R2206 GND.n643 GND.n641 0.114071
R2207 GND.n641 GND.n639 0.114071
R2208 GND.n639 GND.n637 0.114071
R2209 GND.n637 GND.n635 0.114071
R2210 GND.n635 GND.n633 0.114071
R2211 GND.n633 GND.n631 0.114071
R2212 GND.n631 GND.n629 0.114071
R2213 GND.n629 GND.n627 0.114071
R2214 GND.n627 GND.n625 0.114071
R2215 GND.n625 GND.n111 0.114071
R2216 GND.n650 GND.n111 0.114071
R2217 GND.n651 GND.n650 0.114071
R2218 GND.n769 GND.n651 0.114071
R2219 GND.n769 GND.n768 0.114071
R2220 GND.n768 GND.n652 0.114071
R2221 GND.n760 GND.n652 0.114071
R2222 GND.n760 GND.n759 0.114071
R2223 GND.n759 GND.n658 0.114071
R2224 GND.n752 GND.n658 0.114071
R2225 GND.n752 GND.n751 0.114071
R2226 GND.n751 GND.n666 0.114071
R2227 GND.n743 GND.n666 0.114071
R2228 GND.n743 GND.n742 0.114071
R2229 GND.n742 GND.n672 0.114071
R2230 GND.n735 GND.n672 0.114071
R2231 GND.n735 GND.n734 0.114071
R2232 GND.n734 GND.n682 0.114071
R2233 GND.n726 GND.n682 0.114071
R2234 GND.n726 GND.n725 0.114071
R2235 GND.n725 GND.n688 0.114071
R2236 GND.n718 GND.n688 0.114071
R2237 GND.n718 GND.n717 0.114071
R2238 GND.n717 GND.n698 0.114071
R2239 GND.n709 GND.n698 0.114071
R2240 GND.n709 GND.n92 0.114071
R2241 GND.n821 GND.n92 0.114071
R2242 GND.n823 GND.n821 0.114071
R2243 GND.n825 GND.n823 0.114071
R2244 GND.n827 GND.n825 0.114071
R2245 GND.n828 GND.n827 0.114071
R2246 GND.n828 GND.n85 0.114071
R2247 GND.n834 GND.n85 0.114071
R2248 GND.n835 GND.n834 0.114071
R2249 GND.n835 GND.n83 0.114071
R2250 GND.n839 GND.n83 0.114071
R2251 GND.n840 GND.n839 0.114071
R2252 GND.n841 GND.n840 0.114071
R2253 GND.n841 GND.n81 0.114071
R2254 GND.n845 GND.n81 0.114071
R2255 GND.n846 GND.n845 0.114071
R2256 GND.n1279 GND.n846 0.114071
R2257 GND.n1279 GND.n1278 0.114071
R2258 GND.n1278 GND.n1276 0.114071
R2259 GND.n1276 GND.n1274 0.114071
R2260 GND.n1274 GND.n1272 0.114071
R2261 GND.n1272 GND.n1270 0.114071
R2262 GND.n1270 GND.n1268 0.114071
R2263 GND.n1268 GND.n1266 0.114071
R2264 GND.n1266 GND.n1264 0.114071
R2265 GND.n1264 GND.n1262 0.114071
R2266 GND.n1262 GND.n1260 0.114071
R2267 GND.n1260 GND.n1258 0.114071
R2268 GND.n1258 GND.n1256 0.114071
R2269 GND.n1256 GND.n1254 0.114071
R2270 GND.n1254 GND.n1252 0.114071
R2271 GND.n1252 GND.n847 0.114071
R2272 GND.n1245 GND.n847 0.114071
R2273 GND.n1245 GND.n1244 0.114071
R2274 GND.n1244 GND.n851 0.114071
R2275 GND.n1237 GND.n851 0.114071
R2276 GND.n1237 GND.n1236 0.114071
R2277 GND.n1236 GND.n856 0.114071
R2278 GND.n1229 GND.n856 0.114071
R2279 GND.n1229 GND.n1228 0.114071
R2280 GND.n1228 GND.n861 0.114071
R2281 GND.n1221 GND.n861 0.114071
R2282 GND.n1221 GND.n1220 0.114071
R2283 GND.n1220 GND.n866 0.114071
R2284 GND.n1212 GND.n866 0.114071
R2285 GND.n1212 GND.n1211 0.114071
R2286 GND.n1211 GND.n871 0.114071
R2287 GND.n1203 GND.n871 0.114071
R2288 GND.n1203 GND.n1202 0.114071
R2289 GND.n1202 GND.n875 0.114071
R2290 GND.n889 GND.n875 0.114071
R2291 GND.n890 GND.n889 0.114071
R2292 GND.n890 GND.n882 0.114071
R2293 GND.n898 GND.n882 0.114071
R2294 GND.n899 GND.n898 0.114071
R2295 GND.n1193 GND.n899 0.114071
R2296 GND.n1193 GND.n1192 0.114071
R2297 GND.n1192 GND.n900 0.114071
R2298 GND.n1185 GND.n900 0.114071
R2299 GND.n1185 GND.n1184 0.114071
R2300 GND.n1184 GND.n905 0.114071
R2301 GND.n1177 GND.n905 0.114071
R2302 GND.n1177 GND.n1176 0.114071
R2303 GND.n1176 GND.n910 0.114071
R2304 GND.n1169 GND.n910 0.114071
R2305 GND.n1169 GND.n1168 0.114071
R2306 GND.n1168 GND.n915 0.114071
R2307 GND.n1071 GND.n915 0.114071
R2308 GND.n1071 GND.n1070 0.114071
R2309 GND.n1070 GND.n920 0.114071
R2310 GND.n1063 GND.n920 0.114071
R2311 GND.n1063 GND.n1062 0.114071
R2312 GND.n1062 GND.n925 0.114071
R2313 GND.n937 GND.n925 0.114071
R2314 GND.n944 GND.n937 0.114071
R2315 GND.n945 GND.n944 0.114071
R2316 GND.n945 GND.n933 0.114071
R2317 GND.n953 GND.n933 0.114071
R2318 GND.n954 GND.n953 0.114071
R2319 GND.n1053 GND.n954 0.114071
R2320 GND.n1053 GND.n1052 0.114071
R2321 GND.n1052 GND.n955 0.114071
R2322 GND.n1045 GND.n955 0.114071
R2323 GND.n1045 GND.n1044 0.114071
R2324 GND.n1044 GND.n960 0.114071
R2325 GND.n1037 GND.n960 0.114071
R2326 GND.n1037 GND.n1036 0.114071
R2327 GND.n1036 GND.n965 0.114071
R2328 GND.n1029 GND.n965 0.114071
R2329 GND.n1029 GND.n1028 0.114071
R2330 GND.n1028 GND.n970 0.114071
R2331 GND.n1021 GND.n970 0.114071
R2332 GND.n1021 GND.n1020 0.114071
R2333 GND.n1020 GND.n975 0.114071
R2334 GND.n1012 GND.n975 0.114071
R2335 GND.n1012 GND.n1011 0.114071
R2336 GND.n1011 GND.n980 0.114071
R2337 GND.n991 GND.n980 0.114071
R2338 GND.n992 GND.n991 0.114071
R2339 GND.n992 GND.n985 0.114071
R2340 GND.n1000 GND.n985 0.114071
R2341 GND.n1001 GND.n1000 0.114071
R2342 GND.n1001 GND.n19 0.114071
R2343 GND.n1381 GND.n19 0.114071
R2344 GND.n1382 GND.n1381 0.114071
R2345 GND.n1405 GND.n1382 0.114071
R2346 GND.n1405 GND.n1404 0.114071
R2347 GND.n1404 GND.n1402 0.114071
R2348 GND.n1402 GND.n1400 0.114071
R2349 GND.n1400 GND.n1398 0.114071
R2350 GND.n1398 GND.n1396 0.114071
R2351 GND.n1396 GND.n1394 0.114071
R2352 GND.n1394 GND.n1392 0.114071
R2353 GND.n1392 GND.n1390 0.114071
R2354 GND.n1390 GND.n1388 0.114071
R2355 GND.n1388 GND.n1386 0.114071
R2356 GND.n1386 GND.n1384 0.114071
R2357 GND.n1384 GND.n3 0.114071
R2358 GND.n1411 GND.n3 0.114071
R2359 GND.n1412 GND.n1411 0.114071
R2360 GND.n1412 GND.n0 0.114071
R2361 GND.n1941 GND.n1940 0.09575
R2362 GND.n1939 GND.n1699 0.09575
R2363 GND.n373 GND.n320 0.0845084
R2364 GND.n180 GND.n176 0.0632632
R2365 GND.n441 GND.n180 0.0632632
R2366 GND.n441 GND.n440 0.0632632
R2367 GND.n440 GND.n181 0.0632632
R2368 GND.n434 GND.n433 0.0632632
R2369 GND.n433 GND.n432 0.0632632
R2370 GND.n432 GND.n186 0.0632632
R2371 GND.n192 GND.n186 0.0632632
R2372 GND.n425 GND.n192 0.0632632
R2373 GND.n255 GND.n254 0.0632632
R2374 GND.n262 GND.n255 0.0632632
R2375 GND.n263 GND.n262 0.0632632
R2376 GND.n266 GND.n263 0.0632632
R2377 GND.n271 GND.n252 0.0632632
R2378 GND.n272 GND.n271 0.0632632
R2379 GND.n273 GND.n272 0.0632632
R2380 GND.n273 GND.n246 0.0632632
R2381 GND.n280 GND.n246 0.0632632
R2382 GND.n283 GND.n282 0.0632632
R2383 GND.n283 GND.n242 0.0632632
R2384 GND.n289 GND.n242 0.0632632
R2385 GND.n293 GND.n289 0.0632632
R2386 GND.n293 GND.n292 0.0632632
R2387 GND.n300 GND.n239 0.0632632
R2388 GND.n301 GND.n300 0.0632632
R2389 GND.n302 GND.n301 0.0632632
R2390 GND.n302 GND.n234 0.0632632
R2391 GND.n309 GND.n234 0.0632632
R2392 GND GND.n0 0.0572857
R2393 GND GND.n3029 0.0572857
R2394 GND.n424 GND.n423 0.0520132
R2395 GND.n2771 GND.n2739 0.051875
R2396 GND.n2770 GND.n2769 0.051875
R2397 GND.n1977 GND.n1976 0.0483723
R2398 GND.n434 GND.n185 0.0472763
R2399 GND.n379 GND.n310 0.0455
R2400 GND.n291 GND.n239 0.0449079
R2401 GND.n1162 GND.n1161 0.0433571
R2402 GND.t28 GND.t27 0.0414821
R2403 GND.t30 GND.t29 0.041442
R2404 GND.n1420 GND.n1415 0.0410752
R2405 GND.n1420 GND.n1416 0.0410752
R2406 GND.n1358 GND.n1357 0.0407703
R2407 GND.n1349 GND.n36 0.0407245
R2408 GND.n1320 GND.n1319 0.0407245
R2409 GND.n1942 GND.n1941 0.04025
R2410 GND.n1942 GND.n1698 0.04025
R2411 GND.n1946 GND.n1698 0.04025
R2412 GND.n1947 GND.n1946 0.04025
R2413 GND.n1948 GND.n1947 0.04025
R2414 GND.n1948 GND.n1696 0.04025
R2415 GND.n1952 GND.n1696 0.04025
R2416 GND.n1953 GND.n1952 0.04025
R2417 GND.n1954 GND.n1953 0.04025
R2418 GND.n1954 GND.n1694 0.04025
R2419 GND.n1958 GND.n1694 0.04025
R2420 GND.n1959 GND.n1958 0.04025
R2421 GND.n1960 GND.n1959 0.04025
R2422 GND.n1960 GND.n1692 0.04025
R2423 GND.n1964 GND.n1692 0.04025
R2424 GND.n1965 GND.n1964 0.04025
R2425 GND.n1966 GND.n1965 0.04025
R2426 GND.n1966 GND.n1690 0.04025
R2427 GND.n1970 GND.n1690 0.04025
R2428 GND.n1971 GND.n1970 0.04025
R2429 GND.n1972 GND.n1971 0.04025
R2430 GND.n1972 GND.n1688 0.04025
R2431 GND.n1976 GND.n1688 0.04025
R2432 GND.n2502 GND.n2501 0.04025
R2433 GND.n2503 GND.n2502 0.04025
R2434 GND.n2503 GND.n1506 0.04025
R2435 GND.n2507 GND.n1506 0.04025
R2436 GND.n2508 GND.n2507 0.04025
R2437 GND.n2509 GND.n2508 0.04025
R2438 GND.n2509 GND.n1504 0.04025
R2439 GND.n2513 GND.n1504 0.04025
R2440 GND.n2514 GND.n2513 0.04025
R2441 GND.n2515 GND.n2514 0.04025
R2442 GND.n2515 GND.n1502 0.04025
R2443 GND.n2519 GND.n1502 0.04025
R2444 GND.n2520 GND.n2519 0.04025
R2445 GND.n2521 GND.n2520 0.04025
R2446 GND.n2521 GND.n1500 0.04025
R2447 GND.n2525 GND.n1500 0.04025
R2448 GND.n2526 GND.n2525 0.04025
R2449 GND.n2527 GND.n2526 0.04025
R2450 GND.n2527 GND.n1498 0.04025
R2451 GND.n2531 GND.n1498 0.04025
R2452 GND.n2532 GND.n2531 0.04025
R2453 GND.n2533 GND.n2532 0.04025
R2454 GND.n2533 GND.n1496 0.04025
R2455 GND.n2537 GND.n1496 0.04025
R2456 GND.n2538 GND.n2537 0.04025
R2457 GND.n2539 GND.n2538 0.04025
R2458 GND.n2539 GND.n1494 0.04025
R2459 GND.n2543 GND.n1494 0.04025
R2460 GND.n2544 GND.n2543 0.04025
R2461 GND.n2545 GND.n2544 0.04025
R2462 GND.n2545 GND.n1492 0.04025
R2463 GND.n2549 GND.n1492 0.04025
R2464 GND.n2550 GND.n2549 0.04025
R2465 GND.n2551 GND.n2550 0.04025
R2466 GND.n2551 GND.n1490 0.04025
R2467 GND.n2555 GND.n1490 0.04025
R2468 GND.n2556 GND.n2555 0.04025
R2469 GND.n2557 GND.n2556 0.04025
R2470 GND.n2557 GND.n1488 0.04025
R2471 GND.n2561 GND.n1488 0.04025
R2472 GND.n2562 GND.n2561 0.04025
R2473 GND.n2563 GND.n2562 0.04025
R2474 GND.n2563 GND.n1486 0.04025
R2475 GND.n2567 GND.n1486 0.04025
R2476 GND.n2568 GND.n2567 0.04025
R2477 GND.n2569 GND.n2568 0.04025
R2478 GND.n2569 GND.n1484 0.04025
R2479 GND.n2573 GND.n1484 0.04025
R2480 GND.n2574 GND.n2573 0.04025
R2481 GND.n2575 GND.n2574 0.04025
R2482 GND.n2575 GND.n1482 0.04025
R2483 GND.n2579 GND.n1482 0.04025
R2484 GND.n2580 GND.n2579 0.04025
R2485 GND.n2581 GND.n2580 0.04025
R2486 GND.n2581 GND.n1480 0.04025
R2487 GND.n2585 GND.n1480 0.04025
R2488 GND.n2586 GND.n2585 0.04025
R2489 GND.n2587 GND.n2586 0.04025
R2490 GND.n2587 GND.n1478 0.04025
R2491 GND.n2591 GND.n1478 0.04025
R2492 GND.n2592 GND.n2591 0.04025
R2493 GND.n2593 GND.n2592 0.04025
R2494 GND.n2593 GND.n1476 0.04025
R2495 GND.n2597 GND.n1476 0.04025
R2496 GND.n2598 GND.n2597 0.04025
R2497 GND.n2599 GND.n2598 0.04025
R2498 GND.n2599 GND.n1474 0.04025
R2499 GND.n2603 GND.n1474 0.04025
R2500 GND.n2604 GND.n2603 0.04025
R2501 GND.n2605 GND.n2604 0.04025
R2502 GND.n2605 GND.n1472 0.04025
R2503 GND.n2609 GND.n1472 0.04025
R2504 GND.n2610 GND.n2609 0.04025
R2505 GND.n2611 GND.n2610 0.04025
R2506 GND.n2611 GND.n1470 0.04025
R2507 GND.n2615 GND.n1470 0.04025
R2508 GND.n2616 GND.n2615 0.04025
R2509 GND.n2617 GND.n2616 0.04025
R2510 GND.n2617 GND.n1468 0.04025
R2511 GND.n2621 GND.n1468 0.04025
R2512 GND.n2622 GND.n2621 0.04025
R2513 GND.n2623 GND.n2622 0.04025
R2514 GND.n2623 GND.n1466 0.04025
R2515 GND.n2627 GND.n1466 0.04025
R2516 GND.n2628 GND.n2627 0.04025
R2517 GND.n2629 GND.n2628 0.04025
R2518 GND.n2629 GND.n1464 0.04025
R2519 GND.n2633 GND.n1464 0.04025
R2520 GND.n2634 GND.n2633 0.04025
R2521 GND.n2635 GND.n2634 0.04025
R2522 GND.n2635 GND.n1462 0.04025
R2523 GND.n2639 GND.n1462 0.04025
R2524 GND.n2640 GND.n2639 0.04025
R2525 GND.n2641 GND.n2640 0.04025
R2526 GND.n2641 GND.n1460 0.04025
R2527 GND.n2645 GND.n1460 0.04025
R2528 GND.n2646 GND.n2645 0.04025
R2529 GND.n2647 GND.n2646 0.04025
R2530 GND.n2647 GND.n1458 0.04025
R2531 GND.n2651 GND.n1458 0.04025
R2532 GND.n2652 GND.n2651 0.04025
R2533 GND.n2653 GND.n2652 0.04025
R2534 GND.n2653 GND.n1456 0.04025
R2535 GND.n2657 GND.n1456 0.04025
R2536 GND.n2658 GND.n2657 0.04025
R2537 GND.n2659 GND.n2658 0.04025
R2538 GND.n2659 GND.n1454 0.04025
R2539 GND.n2663 GND.n1454 0.04025
R2540 GND.n2664 GND.n2663 0.04025
R2541 GND.n2665 GND.n2664 0.04025
R2542 GND.n2665 GND.n1452 0.04025
R2543 GND.n2669 GND.n1452 0.04025
R2544 GND.n2670 GND.n2669 0.04025
R2545 GND.n2671 GND.n2670 0.04025
R2546 GND.n2671 GND.n1450 0.04025
R2547 GND.n2675 GND.n1450 0.04025
R2548 GND.n2676 GND.n2675 0.04025
R2549 GND.n2677 GND.n2676 0.04025
R2550 GND.n2677 GND.n1447 0.04025
R2551 GND.n2951 GND.n1448 0.04025
R2552 GND.n2947 GND.n1448 0.04025
R2553 GND.n2947 GND.n2946 0.04025
R2554 GND.n2946 GND.n2945 0.04025
R2555 GND.n2945 GND.n2681 0.04025
R2556 GND.n2941 GND.n2681 0.04025
R2557 GND.n2941 GND.n2940 0.04025
R2558 GND.n2940 GND.n2939 0.04025
R2559 GND.n2939 GND.n2683 0.04025
R2560 GND.n2935 GND.n2683 0.04025
R2561 GND.n2935 GND.n2934 0.04025
R2562 GND.n2934 GND.n2933 0.04025
R2563 GND.n2933 GND.n2685 0.04025
R2564 GND.n2929 GND.n2685 0.04025
R2565 GND.n2929 GND.n2928 0.04025
R2566 GND.n2928 GND.n2927 0.04025
R2567 GND.n2927 GND.n2687 0.04025
R2568 GND.n2923 GND.n2687 0.04025
R2569 GND.n2923 GND.n2922 0.04025
R2570 GND.n2922 GND.n2921 0.04025
R2571 GND.n2921 GND.n2689 0.04025
R2572 GND.n2917 GND.n2689 0.04025
R2573 GND.n2917 GND.n2916 0.04025
R2574 GND.n2916 GND.n2915 0.04025
R2575 GND.n2915 GND.n2691 0.04025
R2576 GND.n2911 GND.n2691 0.04025
R2577 GND.n2911 GND.n2910 0.04025
R2578 GND.n2910 GND.n2909 0.04025
R2579 GND.n2909 GND.n2693 0.04025
R2580 GND.n2905 GND.n2693 0.04025
R2581 GND.n2905 GND.n2904 0.04025
R2582 GND.n2904 GND.n2903 0.04025
R2583 GND.n2903 GND.n2695 0.04025
R2584 GND.n2899 GND.n2695 0.04025
R2585 GND.n2899 GND.n2898 0.04025
R2586 GND.n2898 GND.n2897 0.04025
R2587 GND.n2897 GND.n2697 0.04025
R2588 GND.n2893 GND.n2697 0.04025
R2589 GND.n2893 GND.n2892 0.04025
R2590 GND.n2892 GND.n2891 0.04025
R2591 GND.n2891 GND.n2699 0.04025
R2592 GND.n2887 GND.n2699 0.04025
R2593 GND.n2887 GND.n2886 0.04025
R2594 GND.n2886 GND.n2885 0.04025
R2595 GND.n2885 GND.n2701 0.04025
R2596 GND.n2881 GND.n2701 0.04025
R2597 GND.n2881 GND.n2880 0.04025
R2598 GND.n2880 GND.n2879 0.04025
R2599 GND.n2879 GND.n2703 0.04025
R2600 GND.n2875 GND.n2703 0.04025
R2601 GND.n2875 GND.n2874 0.04025
R2602 GND.n2874 GND.n2873 0.04025
R2603 GND.n2873 GND.n2705 0.04025
R2604 GND.n2869 GND.n2705 0.04025
R2605 GND.n2869 GND.n2868 0.04025
R2606 GND.n2868 GND.n2867 0.04025
R2607 GND.n2867 GND.n2707 0.04025
R2608 GND.n2863 GND.n2707 0.04025
R2609 GND.n2863 GND.n2862 0.04025
R2610 GND.n2862 GND.n2861 0.04025
R2611 GND.n2861 GND.n2709 0.04025
R2612 GND.n2857 GND.n2709 0.04025
R2613 GND.n2857 GND.n2856 0.04025
R2614 GND.n2856 GND.n2855 0.04025
R2615 GND.n2855 GND.n2711 0.04025
R2616 GND.n2851 GND.n2711 0.04025
R2617 GND.n2851 GND.n2850 0.04025
R2618 GND.n2850 GND.n2849 0.04025
R2619 GND.n2849 GND.n2713 0.04025
R2620 GND.n2845 GND.n2713 0.04025
R2621 GND.n2845 GND.n2844 0.04025
R2622 GND.n2844 GND.n2843 0.04025
R2623 GND.n2843 GND.n2715 0.04025
R2624 GND.n2839 GND.n2715 0.04025
R2625 GND.n2839 GND.n2838 0.04025
R2626 GND.n2838 GND.n2837 0.04025
R2627 GND.n2837 GND.n2717 0.04025
R2628 GND.n2833 GND.n2717 0.04025
R2629 GND.n2833 GND.n2832 0.04025
R2630 GND.n2832 GND.n2831 0.04025
R2631 GND.n2831 GND.n2719 0.04025
R2632 GND.n2827 GND.n2719 0.04025
R2633 GND.n2827 GND.n2826 0.04025
R2634 GND.n2826 GND.n2825 0.04025
R2635 GND.n2825 GND.n2721 0.04025
R2636 GND.n2821 GND.n2721 0.04025
R2637 GND.n2821 GND.n2820 0.04025
R2638 GND.n2820 GND.n2819 0.04025
R2639 GND.n2819 GND.n2723 0.04025
R2640 GND.n2815 GND.n2723 0.04025
R2641 GND.n2815 GND.n2814 0.04025
R2642 GND.n2814 GND.n2813 0.04025
R2643 GND.n2813 GND.n2725 0.04025
R2644 GND.n2809 GND.n2725 0.04025
R2645 GND.n2809 GND.n2808 0.04025
R2646 GND.n2808 GND.n2807 0.04025
R2647 GND.n2807 GND.n2727 0.04025
R2648 GND.n2803 GND.n2727 0.04025
R2649 GND.n2803 GND.n2802 0.04025
R2650 GND.n2802 GND.n2801 0.04025
R2651 GND.n2801 GND.n2729 0.04025
R2652 GND.n2797 GND.n2729 0.04025
R2653 GND.n2797 GND.n2796 0.04025
R2654 GND.n2796 GND.n2795 0.04025
R2655 GND.n2795 GND.n2731 0.04025
R2656 GND.n2791 GND.n2731 0.04025
R2657 GND.n2791 GND.n2790 0.04025
R2658 GND.n2790 GND.n2789 0.04025
R2659 GND.n2789 GND.n2733 0.04025
R2660 GND.n2785 GND.n2733 0.04025
R2661 GND.n2785 GND.n2784 0.04025
R2662 GND.n2784 GND.n2783 0.04025
R2663 GND.n2783 GND.n2735 0.04025
R2664 GND.n2779 GND.n2735 0.04025
R2665 GND.n2779 GND.n2778 0.04025
R2666 GND.n2778 GND.n2777 0.04025
R2667 GND.n2777 GND.n2737 0.04025
R2668 GND.n2773 GND.n2737 0.04025
R2669 GND.n2773 GND.n2772 0.04025
R2670 GND.n2772 GND.n2771 0.04025
R2671 GND.n2161 GND.n1620 0.04025
R2672 GND.n2165 GND.n1620 0.04025
R2673 GND.n2166 GND.n2165 0.04025
R2674 GND.n2167 GND.n2166 0.04025
R2675 GND.n2167 GND.n1618 0.04025
R2676 GND.n2171 GND.n1618 0.04025
R2677 GND.n2172 GND.n2171 0.04025
R2678 GND.n2173 GND.n2172 0.04025
R2679 GND.n2173 GND.n1616 0.04025
R2680 GND.n2177 GND.n1616 0.04025
R2681 GND.n2178 GND.n2177 0.04025
R2682 GND.n2179 GND.n2178 0.04025
R2683 GND.n2179 GND.n1614 0.04025
R2684 GND.n2183 GND.n1614 0.04025
R2685 GND.n2184 GND.n2183 0.04025
R2686 GND.n2185 GND.n2184 0.04025
R2687 GND.n2185 GND.n1612 0.04025
R2688 GND.n2189 GND.n1612 0.04025
R2689 GND.n2190 GND.n2189 0.04025
R2690 GND.n2191 GND.n2190 0.04025
R2691 GND.n2191 GND.n1610 0.04025
R2692 GND.n2195 GND.n1610 0.04025
R2693 GND.n2196 GND.n2195 0.04025
R2694 GND.n2197 GND.n2196 0.04025
R2695 GND.n2197 GND.n1608 0.04025
R2696 GND.n2201 GND.n1608 0.04025
R2697 GND.n2202 GND.n2201 0.04025
R2698 GND.n2203 GND.n2202 0.04025
R2699 GND.n2203 GND.n1606 0.04025
R2700 GND.n2207 GND.n1606 0.04025
R2701 GND.n2208 GND.n2207 0.04025
R2702 GND.n2209 GND.n2208 0.04025
R2703 GND.n2209 GND.n1604 0.04025
R2704 GND.n2213 GND.n1604 0.04025
R2705 GND.n2214 GND.n2213 0.04025
R2706 GND.n2215 GND.n2214 0.04025
R2707 GND.n2215 GND.n1602 0.04025
R2708 GND.n2219 GND.n1602 0.04025
R2709 GND.n2220 GND.n2219 0.04025
R2710 GND.n2221 GND.n2220 0.04025
R2711 GND.n2221 GND.n1600 0.04025
R2712 GND.n2225 GND.n1600 0.04025
R2713 GND.n2226 GND.n2225 0.04025
R2714 GND.n2227 GND.n2226 0.04025
R2715 GND.n2227 GND.n1598 0.04025
R2716 GND.n2231 GND.n1598 0.04025
R2717 GND.n2232 GND.n2231 0.04025
R2718 GND.n2233 GND.n2232 0.04025
R2719 GND.n2233 GND.n1596 0.04025
R2720 GND.n2237 GND.n1596 0.04025
R2721 GND.n2238 GND.n2237 0.04025
R2722 GND.n2239 GND.n2238 0.04025
R2723 GND.n2239 GND.n1594 0.04025
R2724 GND.n2243 GND.n1594 0.04025
R2725 GND.n2244 GND.n2243 0.04025
R2726 GND.n2245 GND.n2244 0.04025
R2727 GND.n2245 GND.n1592 0.04025
R2728 GND.n2249 GND.n1592 0.04025
R2729 GND.n2250 GND.n2249 0.04025
R2730 GND.n2251 GND.n2250 0.04025
R2731 GND.n2251 GND.n1590 0.04025
R2732 GND.n2255 GND.n1590 0.04025
R2733 GND.n2256 GND.n2255 0.04025
R2734 GND.n2257 GND.n2256 0.04025
R2735 GND.n2257 GND.n1588 0.04025
R2736 GND.n2261 GND.n1588 0.04025
R2737 GND.n2262 GND.n2261 0.04025
R2738 GND.n2263 GND.n2262 0.04025
R2739 GND.n2263 GND.n1586 0.04025
R2740 GND.n2267 GND.n1586 0.04025
R2741 GND.n2268 GND.n2267 0.04025
R2742 GND.n2269 GND.n2268 0.04025
R2743 GND.n2269 GND.n1584 0.04025
R2744 GND.n2273 GND.n1584 0.04025
R2745 GND.n2274 GND.n2273 0.04025
R2746 GND.n2275 GND.n2274 0.04025
R2747 GND.n2275 GND.n1582 0.04025
R2748 GND.n2279 GND.n1582 0.04025
R2749 GND.n2280 GND.n2279 0.04025
R2750 GND.n2281 GND.n2280 0.04025
R2751 GND.n2281 GND.n1580 0.04025
R2752 GND.n2285 GND.n1580 0.04025
R2753 GND.n2286 GND.n2285 0.04025
R2754 GND.n2287 GND.n2286 0.04025
R2755 GND.n2287 GND.n1578 0.04025
R2756 GND.n2291 GND.n1578 0.04025
R2757 GND.n2292 GND.n2291 0.04025
R2758 GND.n2293 GND.n2292 0.04025
R2759 GND.n2293 GND.n1576 0.04025
R2760 GND.n2297 GND.n1576 0.04025
R2761 GND.n2298 GND.n2297 0.04025
R2762 GND.n2299 GND.n2298 0.04025
R2763 GND.n2299 GND.n1574 0.04025
R2764 GND.n2303 GND.n1574 0.04025
R2765 GND.n2304 GND.n2303 0.04025
R2766 GND.n2305 GND.n2304 0.04025
R2767 GND.n2305 GND.n1572 0.04025
R2768 GND.n2309 GND.n1572 0.04025
R2769 GND.n2310 GND.n2309 0.04025
R2770 GND.n2311 GND.n2310 0.04025
R2771 GND.n2311 GND.n1570 0.04025
R2772 GND.n2315 GND.n1570 0.04025
R2773 GND.n2316 GND.n2315 0.04025
R2774 GND.n2317 GND.n2316 0.04025
R2775 GND.n2317 GND.n1568 0.04025
R2776 GND.n2321 GND.n1568 0.04025
R2777 GND.n2322 GND.n2321 0.04025
R2778 GND.n2323 GND.n2322 0.04025
R2779 GND.n2323 GND.n1566 0.04025
R2780 GND.n2327 GND.n1566 0.04025
R2781 GND.n2328 GND.n2327 0.04025
R2782 GND.n2329 GND.n2328 0.04025
R2783 GND.n2329 GND.n1564 0.04025
R2784 GND.n2333 GND.n1564 0.04025
R2785 GND.n2334 GND.n2333 0.04025
R2786 GND.n2335 GND.n2334 0.04025
R2787 GND.n2335 GND.n1562 0.04025
R2788 GND.n2339 GND.n1562 0.04025
R2789 GND.n2340 GND.n2339 0.04025
R2790 GND.n2341 GND.n2340 0.04025
R2791 GND.n2341 GND.n1560 0.04025
R2792 GND.n2345 GND.n1560 0.04025
R2793 GND.n2346 GND.n2345 0.04025
R2794 GND.n2347 GND.n2346 0.04025
R2795 GND.n2347 GND.n1558 0.04025
R2796 GND.n2351 GND.n1558 0.04025
R2797 GND.n2352 GND.n2351 0.04025
R2798 GND.n2353 GND.n2352 0.04025
R2799 GND.n2353 GND.n1556 0.04025
R2800 GND.n2357 GND.n1556 0.04025
R2801 GND.n2358 GND.n2357 0.04025
R2802 GND.n2359 GND.n2358 0.04025
R2803 GND.n2359 GND.n1554 0.04025
R2804 GND.n2363 GND.n1554 0.04025
R2805 GND.n2364 GND.n2363 0.04025
R2806 GND.n2365 GND.n2364 0.04025
R2807 GND.n2365 GND.n1552 0.04025
R2808 GND.n2369 GND.n1552 0.04025
R2809 GND.n2370 GND.n2369 0.04025
R2810 GND.n2371 GND.n2370 0.04025
R2811 GND.n2371 GND.n1550 0.04025
R2812 GND.n2375 GND.n1550 0.04025
R2813 GND.n2376 GND.n2375 0.04025
R2814 GND.n2377 GND.n2376 0.04025
R2815 GND.n2377 GND.n1548 0.04025
R2816 GND.n2381 GND.n1548 0.04025
R2817 GND.n2382 GND.n2381 0.04025
R2818 GND.n2383 GND.n2382 0.04025
R2819 GND.n2383 GND.n1546 0.04025
R2820 GND.n2387 GND.n1546 0.04025
R2821 GND.n2388 GND.n2387 0.04025
R2822 GND.n2389 GND.n2388 0.04025
R2823 GND.n2389 GND.n1544 0.04025
R2824 GND.n2393 GND.n1544 0.04025
R2825 GND.n2394 GND.n2393 0.04025
R2826 GND.n2395 GND.n2394 0.04025
R2827 GND.n2395 GND.n1542 0.04025
R2828 GND.n2399 GND.n1542 0.04025
R2829 GND.n2400 GND.n2399 0.04025
R2830 GND.n2401 GND.n2400 0.04025
R2831 GND.n2401 GND.n1540 0.04025
R2832 GND.n2405 GND.n1540 0.04025
R2833 GND.n2406 GND.n2405 0.04025
R2834 GND.n2407 GND.n2406 0.04025
R2835 GND.n2407 GND.n1538 0.04025
R2836 GND.n2411 GND.n1538 0.04025
R2837 GND.n2412 GND.n2411 0.04025
R2838 GND.n2413 GND.n2412 0.04025
R2839 GND.n2413 GND.n1536 0.04025
R2840 GND.n2417 GND.n1536 0.04025
R2841 GND.n2418 GND.n2417 0.04025
R2842 GND.n2419 GND.n2418 0.04025
R2843 GND.n2419 GND.n1534 0.04025
R2844 GND.n2423 GND.n1534 0.04025
R2845 GND.n2424 GND.n2423 0.04025
R2846 GND.n2425 GND.n2424 0.04025
R2847 GND.n2425 GND.n1532 0.04025
R2848 GND.n2429 GND.n1532 0.04025
R2849 GND.n2430 GND.n2429 0.04025
R2850 GND.n2431 GND.n2430 0.04025
R2851 GND.n2431 GND.n1530 0.04025
R2852 GND.n2435 GND.n1530 0.04025
R2853 GND.n2436 GND.n2435 0.04025
R2854 GND.n2437 GND.n2436 0.04025
R2855 GND.n2437 GND.n1528 0.04025
R2856 GND.n2441 GND.n1528 0.04025
R2857 GND.n2442 GND.n2441 0.04025
R2858 GND.n2443 GND.n2442 0.04025
R2859 GND.n2443 GND.n1526 0.04025
R2860 GND.n2447 GND.n1526 0.04025
R2861 GND.n2448 GND.n2447 0.04025
R2862 GND.n2449 GND.n2448 0.04025
R2863 GND.n2449 GND.n1524 0.04025
R2864 GND.n2453 GND.n1524 0.04025
R2865 GND.n2454 GND.n2453 0.04025
R2866 GND.n2455 GND.n2454 0.04025
R2867 GND.n2455 GND.n1522 0.04025
R2868 GND.n2459 GND.n1522 0.04025
R2869 GND.n2460 GND.n2459 0.04025
R2870 GND.n2461 GND.n2460 0.04025
R2871 GND.n2461 GND.n1520 0.04025
R2872 GND.n2465 GND.n1520 0.04025
R2873 GND.n2466 GND.n2465 0.04025
R2874 GND.n2467 GND.n2466 0.04025
R2875 GND.n2467 GND.n1518 0.04025
R2876 GND.n2471 GND.n1518 0.04025
R2877 GND.n2472 GND.n2471 0.04025
R2878 GND.n2473 GND.n2472 0.04025
R2879 GND.n2473 GND.n1516 0.04025
R2880 GND.n2477 GND.n1516 0.04025
R2881 GND.n2478 GND.n2477 0.04025
R2882 GND.n2479 GND.n2478 0.04025
R2883 GND.n2479 GND.n1514 0.04025
R2884 GND.n2483 GND.n1514 0.04025
R2885 GND.n2484 GND.n2483 0.04025
R2886 GND.n2485 GND.n2484 0.04025
R2887 GND.n2485 GND.n1512 0.04025
R2888 GND.n2489 GND.n1512 0.04025
R2889 GND.n2490 GND.n2489 0.04025
R2890 GND.n2491 GND.n2490 0.04025
R2891 GND.n2491 GND.n1510 0.04025
R2892 GND.n2495 GND.n1510 0.04025
R2893 GND.n2496 GND.n2495 0.04025
R2894 GND.n2497 GND.n2496 0.04025
R2895 GND.n2159 GND.n1622 0.04025
R2896 GND.n2155 GND.n1622 0.04025
R2897 GND.n2155 GND.n2154 0.04025
R2898 GND.n2154 GND.n2153 0.04025
R2899 GND.n2153 GND.n1624 0.04025
R2900 GND.n2149 GND.n1624 0.04025
R2901 GND.n2149 GND.n2148 0.04025
R2902 GND.n2148 GND.n2147 0.04025
R2903 GND.n2147 GND.n1626 0.04025
R2904 GND.n2143 GND.n1626 0.04025
R2905 GND.n2143 GND.n2142 0.04025
R2906 GND.n2142 GND.n2141 0.04025
R2907 GND.n2141 GND.n1628 0.04025
R2908 GND.n2137 GND.n1628 0.04025
R2909 GND.n2137 GND.n2136 0.04025
R2910 GND.n2136 GND.n2135 0.04025
R2911 GND.n2135 GND.n1630 0.04025
R2912 GND.n2131 GND.n1630 0.04025
R2913 GND.n2131 GND.n2130 0.04025
R2914 GND.n2130 GND.n2129 0.04025
R2915 GND.n2129 GND.n1632 0.04025
R2916 GND.n2125 GND.n1632 0.04025
R2917 GND.n2125 GND.n2124 0.04025
R2918 GND.n2124 GND.n2123 0.04025
R2919 GND.n2123 GND.n1634 0.04025
R2920 GND.n2119 GND.n1634 0.04025
R2921 GND.n2119 GND.n2118 0.04025
R2922 GND.n2118 GND.n2117 0.04025
R2923 GND.n2117 GND.n1636 0.04025
R2924 GND.n2113 GND.n1636 0.04025
R2925 GND.n2113 GND.n2112 0.04025
R2926 GND.n2112 GND.n2111 0.04025
R2927 GND.n2111 GND.n1638 0.04025
R2928 GND.n2107 GND.n1638 0.04025
R2929 GND.n2107 GND.n2106 0.04025
R2930 GND.n2106 GND.n2105 0.04025
R2931 GND.n2105 GND.n1640 0.04025
R2932 GND.n2101 GND.n1640 0.04025
R2933 GND.n2101 GND.n2100 0.04025
R2934 GND.n2100 GND.n2099 0.04025
R2935 GND.n2099 GND.n1642 0.04025
R2936 GND.n2095 GND.n1642 0.04025
R2937 GND.n2095 GND.n2094 0.04025
R2938 GND.n2094 GND.n2093 0.04025
R2939 GND.n2093 GND.n1644 0.04025
R2940 GND.n2089 GND.n1644 0.04025
R2941 GND.n2089 GND.n2088 0.04025
R2942 GND.n2088 GND.n2087 0.04025
R2943 GND.n2087 GND.n1646 0.04025
R2944 GND.n2083 GND.n1646 0.04025
R2945 GND.n2083 GND.n2082 0.04025
R2946 GND.n2082 GND.n2081 0.04025
R2947 GND.n2081 GND.n1648 0.04025
R2948 GND.n2077 GND.n1648 0.04025
R2949 GND.n2077 GND.n2076 0.04025
R2950 GND.n2076 GND.n2075 0.04025
R2951 GND.n2075 GND.n1650 0.04025
R2952 GND.n2071 GND.n1650 0.04025
R2953 GND.n2071 GND.n2070 0.04025
R2954 GND.n2070 GND.n2069 0.04025
R2955 GND.n2069 GND.n1652 0.04025
R2956 GND.n2065 GND.n1652 0.04025
R2957 GND.n2065 GND.n2064 0.04025
R2958 GND.n2064 GND.n2063 0.04025
R2959 GND.n2063 GND.n1654 0.04025
R2960 GND.n2059 GND.n1654 0.04025
R2961 GND.n2059 GND.n2058 0.04025
R2962 GND.n2058 GND.n2057 0.04025
R2963 GND.n2057 GND.n1656 0.04025
R2964 GND.n2053 GND.n1656 0.04025
R2965 GND.n2053 GND.n2052 0.04025
R2966 GND.n2052 GND.n2051 0.04025
R2967 GND.n2051 GND.n1658 0.04025
R2968 GND.n2047 GND.n1658 0.04025
R2969 GND.n2047 GND.n2046 0.04025
R2970 GND.n2046 GND.n2045 0.04025
R2971 GND.n2045 GND.n1660 0.04025
R2972 GND.n2041 GND.n1660 0.04025
R2973 GND.n2041 GND.n2040 0.04025
R2974 GND.n2040 GND.n2039 0.04025
R2975 GND.n2039 GND.n1662 0.04025
R2976 GND.n2035 GND.n1662 0.04025
R2977 GND.n2035 GND.n2034 0.04025
R2978 GND.n2034 GND.n2033 0.04025
R2979 GND.n2033 GND.n1664 0.04025
R2980 GND.n2029 GND.n1664 0.04025
R2981 GND.n2029 GND.n2028 0.04025
R2982 GND.n2028 GND.n2027 0.04025
R2983 GND.n2027 GND.n1666 0.04025
R2984 GND.n2023 GND.n1666 0.04025
R2985 GND.n2023 GND.n2022 0.04025
R2986 GND.n2022 GND.n2021 0.04025
R2987 GND.n2021 GND.n1668 0.04025
R2988 GND.n2017 GND.n1668 0.04025
R2989 GND.n2017 GND.n2016 0.04025
R2990 GND.n2016 GND.n2015 0.04025
R2991 GND.n2015 GND.n1670 0.04025
R2992 GND.n2011 GND.n1670 0.04025
R2993 GND.n2011 GND.n2010 0.04025
R2994 GND.n2010 GND.n2009 0.04025
R2995 GND.n2009 GND.n1672 0.04025
R2996 GND.n2005 GND.n1672 0.04025
R2997 GND.n2005 GND.n2004 0.04025
R2998 GND.n2004 GND.n2003 0.04025
R2999 GND.n2003 GND.n1674 0.04025
R3000 GND.n1999 GND.n1674 0.04025
R3001 GND.n1999 GND.n1998 0.04025
R3002 GND.n1998 GND.n1997 0.04025
R3003 GND.n1997 GND.n1676 0.04025
R3004 GND.n1993 GND.n1676 0.04025
R3005 GND.n1993 GND.n1992 0.04025
R3006 GND.n1992 GND.n1991 0.04025
R3007 GND.n1991 GND.n1678 0.04025
R3008 GND.n1987 GND.n1678 0.04025
R3009 GND.n1987 GND.n1986 0.04025
R3010 GND.n1986 GND.n1985 0.04025
R3011 GND.n1985 GND.n1680 0.04025
R3012 GND.n1981 GND.n1680 0.04025
R3013 GND.n1981 GND.n1980 0.04025
R3014 GND.n1761 GND.n1682 0.04025
R3015 GND.n1762 GND.n1761 0.04025
R3016 GND.n1762 GND.n1758 0.04025
R3017 GND.n1766 GND.n1758 0.04025
R3018 GND.n1767 GND.n1766 0.04025
R3019 GND.n1768 GND.n1767 0.04025
R3020 GND.n1768 GND.n1756 0.04025
R3021 GND.n1772 GND.n1756 0.04025
R3022 GND.n1773 GND.n1772 0.04025
R3023 GND.n1774 GND.n1773 0.04025
R3024 GND.n1774 GND.n1754 0.04025
R3025 GND.n1778 GND.n1754 0.04025
R3026 GND.n1779 GND.n1778 0.04025
R3027 GND.n1780 GND.n1779 0.04025
R3028 GND.n1780 GND.n1752 0.04025
R3029 GND.n1784 GND.n1752 0.04025
R3030 GND.n1785 GND.n1784 0.04025
R3031 GND.n1786 GND.n1785 0.04025
R3032 GND.n1786 GND.n1750 0.04025
R3033 GND.n1790 GND.n1750 0.04025
R3034 GND.n1791 GND.n1790 0.04025
R3035 GND.n1792 GND.n1791 0.04025
R3036 GND.n1792 GND.n1748 0.04025
R3037 GND.n1796 GND.n1748 0.04025
R3038 GND.n1797 GND.n1796 0.04025
R3039 GND.n1798 GND.n1797 0.04025
R3040 GND.n1798 GND.n1746 0.04025
R3041 GND.n1802 GND.n1746 0.04025
R3042 GND.n1803 GND.n1802 0.04025
R3043 GND.n1804 GND.n1803 0.04025
R3044 GND.n1804 GND.n1744 0.04025
R3045 GND.n1808 GND.n1744 0.04025
R3046 GND.n1809 GND.n1808 0.04025
R3047 GND.n1810 GND.n1809 0.04025
R3048 GND.n1810 GND.n1742 0.04025
R3049 GND.n1814 GND.n1742 0.04025
R3050 GND.n1815 GND.n1814 0.04025
R3051 GND.n1816 GND.n1815 0.04025
R3052 GND.n1816 GND.n1740 0.04025
R3053 GND.n1820 GND.n1740 0.04025
R3054 GND.n1821 GND.n1820 0.04025
R3055 GND.n1822 GND.n1821 0.04025
R3056 GND.n1822 GND.n1738 0.04025
R3057 GND.n1826 GND.n1738 0.04025
R3058 GND.n1827 GND.n1826 0.04025
R3059 GND.n1828 GND.n1827 0.04025
R3060 GND.n1828 GND.n1736 0.04025
R3061 GND.n1832 GND.n1736 0.04025
R3062 GND.n1833 GND.n1832 0.04025
R3063 GND.n1834 GND.n1833 0.04025
R3064 GND.n1834 GND.n1734 0.04025
R3065 GND.n1838 GND.n1734 0.04025
R3066 GND.n1839 GND.n1838 0.04025
R3067 GND.n1840 GND.n1839 0.04025
R3068 GND.n1840 GND.n1732 0.04025
R3069 GND.n1844 GND.n1732 0.04025
R3070 GND.n1845 GND.n1844 0.04025
R3071 GND.n1846 GND.n1845 0.04025
R3072 GND.n1846 GND.n1730 0.04025
R3073 GND.n1850 GND.n1730 0.04025
R3074 GND.n1851 GND.n1850 0.04025
R3075 GND.n1852 GND.n1851 0.04025
R3076 GND.n1852 GND.n1728 0.04025
R3077 GND.n1856 GND.n1728 0.04025
R3078 GND.n1857 GND.n1856 0.04025
R3079 GND.n1858 GND.n1857 0.04025
R3080 GND.n1858 GND.n1726 0.04025
R3081 GND.n1862 GND.n1726 0.04025
R3082 GND.n1863 GND.n1862 0.04025
R3083 GND.n1864 GND.n1863 0.04025
R3084 GND.n1864 GND.n1724 0.04025
R3085 GND.n1868 GND.n1724 0.04025
R3086 GND.n1869 GND.n1868 0.04025
R3087 GND.n1870 GND.n1869 0.04025
R3088 GND.n1870 GND.n1722 0.04025
R3089 GND.n1874 GND.n1722 0.04025
R3090 GND.n1875 GND.n1874 0.04025
R3091 GND.n1876 GND.n1875 0.04025
R3092 GND.n1876 GND.n1720 0.04025
R3093 GND.n1880 GND.n1720 0.04025
R3094 GND.n1881 GND.n1880 0.04025
R3095 GND.n1882 GND.n1881 0.04025
R3096 GND.n1882 GND.n1718 0.04025
R3097 GND.n1886 GND.n1718 0.04025
R3098 GND.n1887 GND.n1886 0.04025
R3099 GND.n1888 GND.n1887 0.04025
R3100 GND.n1888 GND.n1716 0.04025
R3101 GND.n1892 GND.n1716 0.04025
R3102 GND.n1893 GND.n1892 0.04025
R3103 GND.n1894 GND.n1893 0.04025
R3104 GND.n1894 GND.n1714 0.04025
R3105 GND.n1898 GND.n1714 0.04025
R3106 GND.n1899 GND.n1898 0.04025
R3107 GND.n1900 GND.n1899 0.04025
R3108 GND.n1900 GND.n1712 0.04025
R3109 GND.n1904 GND.n1712 0.04025
R3110 GND.n1905 GND.n1904 0.04025
R3111 GND.n1906 GND.n1905 0.04025
R3112 GND.n1906 GND.n1710 0.04025
R3113 GND.n1910 GND.n1710 0.04025
R3114 GND.n1911 GND.n1910 0.04025
R3115 GND.n1912 GND.n1911 0.04025
R3116 GND.n1912 GND.n1708 0.04025
R3117 GND.n1916 GND.n1708 0.04025
R3118 GND.n1917 GND.n1916 0.04025
R3119 GND.n1918 GND.n1917 0.04025
R3120 GND.n1918 GND.n1706 0.04025
R3121 GND.n1922 GND.n1706 0.04025
R3122 GND.n1923 GND.n1922 0.04025
R3123 GND.n1924 GND.n1923 0.04025
R3124 GND.n1924 GND.n1704 0.04025
R3125 GND.n1928 GND.n1704 0.04025
R3126 GND.n1929 GND.n1928 0.04025
R3127 GND.n1930 GND.n1929 0.04025
R3128 GND.n1930 GND.n1702 0.04025
R3129 GND.n1934 GND.n1702 0.04025
R3130 GND.n1935 GND.n1934 0.04025
R3131 GND.n1936 GND.n1935 0.04025
R3132 GND.n1936 GND.n1700 0.04025
R3133 GND.n1940 GND.n1700 0.04025
R3134 GND.n2158 GND.n2157 0.04025
R3135 GND.n2157 GND.n2156 0.04025
R3136 GND.n2156 GND.n1623 0.04025
R3137 GND.n2152 GND.n1623 0.04025
R3138 GND.n2152 GND.n2151 0.04025
R3139 GND.n2151 GND.n2150 0.04025
R3140 GND.n2150 GND.n1625 0.04025
R3141 GND.n2146 GND.n1625 0.04025
R3142 GND.n2146 GND.n2145 0.04025
R3143 GND.n2145 GND.n2144 0.04025
R3144 GND.n2144 GND.n1627 0.04025
R3145 GND.n2140 GND.n1627 0.04025
R3146 GND.n2140 GND.n2139 0.04025
R3147 GND.n2139 GND.n2138 0.04025
R3148 GND.n2138 GND.n1629 0.04025
R3149 GND.n2134 GND.n1629 0.04025
R3150 GND.n2134 GND.n2133 0.04025
R3151 GND.n2133 GND.n2132 0.04025
R3152 GND.n2132 GND.n1631 0.04025
R3153 GND.n2128 GND.n1631 0.04025
R3154 GND.n2128 GND.n2127 0.04025
R3155 GND.n2127 GND.n2126 0.04025
R3156 GND.n2126 GND.n1633 0.04025
R3157 GND.n2122 GND.n1633 0.04025
R3158 GND.n2122 GND.n2121 0.04025
R3159 GND.n2121 GND.n2120 0.04025
R3160 GND.n2120 GND.n1635 0.04025
R3161 GND.n2116 GND.n1635 0.04025
R3162 GND.n2116 GND.n2115 0.04025
R3163 GND.n2115 GND.n2114 0.04025
R3164 GND.n2114 GND.n1637 0.04025
R3165 GND.n2110 GND.n1637 0.04025
R3166 GND.n2110 GND.n2109 0.04025
R3167 GND.n2109 GND.n2108 0.04025
R3168 GND.n2108 GND.n1639 0.04025
R3169 GND.n2104 GND.n1639 0.04025
R3170 GND.n2104 GND.n2103 0.04025
R3171 GND.n2103 GND.n2102 0.04025
R3172 GND.n2102 GND.n1641 0.04025
R3173 GND.n2098 GND.n1641 0.04025
R3174 GND.n2098 GND.n2097 0.04025
R3175 GND.n2097 GND.n2096 0.04025
R3176 GND.n2096 GND.n1643 0.04025
R3177 GND.n2092 GND.n1643 0.04025
R3178 GND.n2092 GND.n2091 0.04025
R3179 GND.n2091 GND.n2090 0.04025
R3180 GND.n2090 GND.n1645 0.04025
R3181 GND.n2086 GND.n1645 0.04025
R3182 GND.n2086 GND.n2085 0.04025
R3183 GND.n2085 GND.n2084 0.04025
R3184 GND.n2084 GND.n1647 0.04025
R3185 GND.n2080 GND.n1647 0.04025
R3186 GND.n2080 GND.n2079 0.04025
R3187 GND.n2079 GND.n2078 0.04025
R3188 GND.n2078 GND.n1649 0.04025
R3189 GND.n2074 GND.n1649 0.04025
R3190 GND.n2074 GND.n2073 0.04025
R3191 GND.n2073 GND.n2072 0.04025
R3192 GND.n2072 GND.n1651 0.04025
R3193 GND.n2068 GND.n1651 0.04025
R3194 GND.n2068 GND.n2067 0.04025
R3195 GND.n2067 GND.n2066 0.04025
R3196 GND.n2066 GND.n1653 0.04025
R3197 GND.n2062 GND.n1653 0.04025
R3198 GND.n2062 GND.n2061 0.04025
R3199 GND.n2061 GND.n2060 0.04025
R3200 GND.n2060 GND.n1655 0.04025
R3201 GND.n2056 GND.n1655 0.04025
R3202 GND.n2056 GND.n2055 0.04025
R3203 GND.n2055 GND.n2054 0.04025
R3204 GND.n2054 GND.n1657 0.04025
R3205 GND.n2050 GND.n1657 0.04025
R3206 GND.n2050 GND.n2049 0.04025
R3207 GND.n2049 GND.n2048 0.04025
R3208 GND.n2048 GND.n1659 0.04025
R3209 GND.n2044 GND.n1659 0.04025
R3210 GND.n2044 GND.n2043 0.04025
R3211 GND.n2043 GND.n2042 0.04025
R3212 GND.n2042 GND.n1661 0.04025
R3213 GND.n2038 GND.n1661 0.04025
R3214 GND.n2038 GND.n2037 0.04025
R3215 GND.n2037 GND.n2036 0.04025
R3216 GND.n2036 GND.n1663 0.04025
R3217 GND.n2032 GND.n1663 0.04025
R3218 GND.n2032 GND.n2031 0.04025
R3219 GND.n2031 GND.n2030 0.04025
R3220 GND.n2030 GND.n1665 0.04025
R3221 GND.n2026 GND.n1665 0.04025
R3222 GND.n2026 GND.n2025 0.04025
R3223 GND.n2025 GND.n2024 0.04025
R3224 GND.n2024 GND.n1667 0.04025
R3225 GND.n2020 GND.n1667 0.04025
R3226 GND.n2020 GND.n2019 0.04025
R3227 GND.n2019 GND.n2018 0.04025
R3228 GND.n2018 GND.n1669 0.04025
R3229 GND.n2014 GND.n1669 0.04025
R3230 GND.n2014 GND.n2013 0.04025
R3231 GND.n2013 GND.n2012 0.04025
R3232 GND.n2012 GND.n1671 0.04025
R3233 GND.n2008 GND.n1671 0.04025
R3234 GND.n2008 GND.n2007 0.04025
R3235 GND.n2007 GND.n2006 0.04025
R3236 GND.n2006 GND.n1673 0.04025
R3237 GND.n2002 GND.n1673 0.04025
R3238 GND.n2002 GND.n2001 0.04025
R3239 GND.n2001 GND.n2000 0.04025
R3240 GND.n2000 GND.n1675 0.04025
R3241 GND.n1996 GND.n1675 0.04025
R3242 GND.n1996 GND.n1995 0.04025
R3243 GND.n1995 GND.n1994 0.04025
R3244 GND.n1994 GND.n1677 0.04025
R3245 GND.n1990 GND.n1677 0.04025
R3246 GND.n1990 GND.n1989 0.04025
R3247 GND.n1989 GND.n1988 0.04025
R3248 GND.n1988 GND.n1679 0.04025
R3249 GND.n1984 GND.n1679 0.04025
R3250 GND.n1984 GND.n1983 0.04025
R3251 GND.n1983 GND.n1982 0.04025
R3252 GND.n1982 GND.n1681 0.04025
R3253 GND.n1759 GND.n1681 0.04025
R3254 GND.n1760 GND.n1759 0.04025
R3255 GND.n1763 GND.n1760 0.04025
R3256 GND.n1764 GND.n1763 0.04025
R3257 GND.n1765 GND.n1764 0.04025
R3258 GND.n1765 GND.n1757 0.04025
R3259 GND.n1769 GND.n1757 0.04025
R3260 GND.n1770 GND.n1769 0.04025
R3261 GND.n1771 GND.n1770 0.04025
R3262 GND.n1771 GND.n1755 0.04025
R3263 GND.n1775 GND.n1755 0.04025
R3264 GND.n1776 GND.n1775 0.04025
R3265 GND.n1777 GND.n1776 0.04025
R3266 GND.n1777 GND.n1753 0.04025
R3267 GND.n1781 GND.n1753 0.04025
R3268 GND.n1782 GND.n1781 0.04025
R3269 GND.n1783 GND.n1782 0.04025
R3270 GND.n1783 GND.n1751 0.04025
R3271 GND.n1787 GND.n1751 0.04025
R3272 GND.n1788 GND.n1787 0.04025
R3273 GND.n1789 GND.n1788 0.04025
R3274 GND.n1789 GND.n1749 0.04025
R3275 GND.n1793 GND.n1749 0.04025
R3276 GND.n1794 GND.n1793 0.04025
R3277 GND.n1795 GND.n1794 0.04025
R3278 GND.n1795 GND.n1747 0.04025
R3279 GND.n1799 GND.n1747 0.04025
R3280 GND.n1800 GND.n1799 0.04025
R3281 GND.n1801 GND.n1800 0.04025
R3282 GND.n1801 GND.n1745 0.04025
R3283 GND.n1805 GND.n1745 0.04025
R3284 GND.n1806 GND.n1805 0.04025
R3285 GND.n1807 GND.n1806 0.04025
R3286 GND.n1807 GND.n1743 0.04025
R3287 GND.n1811 GND.n1743 0.04025
R3288 GND.n1812 GND.n1811 0.04025
R3289 GND.n1813 GND.n1812 0.04025
R3290 GND.n1813 GND.n1741 0.04025
R3291 GND.n1817 GND.n1741 0.04025
R3292 GND.n1818 GND.n1817 0.04025
R3293 GND.n1819 GND.n1818 0.04025
R3294 GND.n1819 GND.n1739 0.04025
R3295 GND.n1823 GND.n1739 0.04025
R3296 GND.n1824 GND.n1823 0.04025
R3297 GND.n1825 GND.n1824 0.04025
R3298 GND.n1825 GND.n1737 0.04025
R3299 GND.n1829 GND.n1737 0.04025
R3300 GND.n1830 GND.n1829 0.04025
R3301 GND.n1831 GND.n1830 0.04025
R3302 GND.n1831 GND.n1735 0.04025
R3303 GND.n1835 GND.n1735 0.04025
R3304 GND.n1836 GND.n1835 0.04025
R3305 GND.n1837 GND.n1836 0.04025
R3306 GND.n1837 GND.n1733 0.04025
R3307 GND.n1841 GND.n1733 0.04025
R3308 GND.n1842 GND.n1841 0.04025
R3309 GND.n1843 GND.n1842 0.04025
R3310 GND.n1843 GND.n1731 0.04025
R3311 GND.n1847 GND.n1731 0.04025
R3312 GND.n1848 GND.n1847 0.04025
R3313 GND.n1849 GND.n1848 0.04025
R3314 GND.n1849 GND.n1729 0.04025
R3315 GND.n1853 GND.n1729 0.04025
R3316 GND.n1854 GND.n1853 0.04025
R3317 GND.n1855 GND.n1854 0.04025
R3318 GND.n1855 GND.n1727 0.04025
R3319 GND.n1859 GND.n1727 0.04025
R3320 GND.n1860 GND.n1859 0.04025
R3321 GND.n1861 GND.n1860 0.04025
R3322 GND.n1861 GND.n1725 0.04025
R3323 GND.n1865 GND.n1725 0.04025
R3324 GND.n1866 GND.n1865 0.04025
R3325 GND.n1867 GND.n1866 0.04025
R3326 GND.n1867 GND.n1723 0.04025
R3327 GND.n1871 GND.n1723 0.04025
R3328 GND.n1872 GND.n1871 0.04025
R3329 GND.n1873 GND.n1872 0.04025
R3330 GND.n1873 GND.n1721 0.04025
R3331 GND.n1877 GND.n1721 0.04025
R3332 GND.n1878 GND.n1877 0.04025
R3333 GND.n1879 GND.n1878 0.04025
R3334 GND.n1879 GND.n1719 0.04025
R3335 GND.n1883 GND.n1719 0.04025
R3336 GND.n1884 GND.n1883 0.04025
R3337 GND.n1885 GND.n1884 0.04025
R3338 GND.n1885 GND.n1717 0.04025
R3339 GND.n1889 GND.n1717 0.04025
R3340 GND.n1890 GND.n1889 0.04025
R3341 GND.n1891 GND.n1890 0.04025
R3342 GND.n1891 GND.n1715 0.04025
R3343 GND.n1895 GND.n1715 0.04025
R3344 GND.n1896 GND.n1895 0.04025
R3345 GND.n1897 GND.n1896 0.04025
R3346 GND.n1897 GND.n1713 0.04025
R3347 GND.n1901 GND.n1713 0.04025
R3348 GND.n1902 GND.n1901 0.04025
R3349 GND.n1903 GND.n1902 0.04025
R3350 GND.n1903 GND.n1711 0.04025
R3351 GND.n1907 GND.n1711 0.04025
R3352 GND.n1908 GND.n1907 0.04025
R3353 GND.n1909 GND.n1908 0.04025
R3354 GND.n1909 GND.n1709 0.04025
R3355 GND.n1913 GND.n1709 0.04025
R3356 GND.n1914 GND.n1913 0.04025
R3357 GND.n1915 GND.n1914 0.04025
R3358 GND.n1915 GND.n1707 0.04025
R3359 GND.n1919 GND.n1707 0.04025
R3360 GND.n1920 GND.n1919 0.04025
R3361 GND.n1921 GND.n1920 0.04025
R3362 GND.n1921 GND.n1705 0.04025
R3363 GND.n1925 GND.n1705 0.04025
R3364 GND.n1926 GND.n1925 0.04025
R3365 GND.n1927 GND.n1926 0.04025
R3366 GND.n1927 GND.n1703 0.04025
R3367 GND.n1931 GND.n1703 0.04025
R3368 GND.n1932 GND.n1931 0.04025
R3369 GND.n1933 GND.n1932 0.04025
R3370 GND.n1933 GND.n1701 0.04025
R3371 GND.n1937 GND.n1701 0.04025
R3372 GND.n1938 GND.n1937 0.04025
R3373 GND.n1939 GND.n1938 0.04025
R3374 GND.n2163 GND.n2162 0.04025
R3375 GND.n2164 GND.n2163 0.04025
R3376 GND.n2164 GND.n1619 0.04025
R3377 GND.n2168 GND.n1619 0.04025
R3378 GND.n2169 GND.n2168 0.04025
R3379 GND.n2170 GND.n2169 0.04025
R3380 GND.n2170 GND.n1617 0.04025
R3381 GND.n2174 GND.n1617 0.04025
R3382 GND.n2175 GND.n2174 0.04025
R3383 GND.n2176 GND.n2175 0.04025
R3384 GND.n2176 GND.n1615 0.04025
R3385 GND.n2180 GND.n1615 0.04025
R3386 GND.n2181 GND.n2180 0.04025
R3387 GND.n2182 GND.n2181 0.04025
R3388 GND.n2182 GND.n1613 0.04025
R3389 GND.n2186 GND.n1613 0.04025
R3390 GND.n2187 GND.n2186 0.04025
R3391 GND.n2188 GND.n2187 0.04025
R3392 GND.n2188 GND.n1611 0.04025
R3393 GND.n2192 GND.n1611 0.04025
R3394 GND.n2193 GND.n2192 0.04025
R3395 GND.n2194 GND.n2193 0.04025
R3396 GND.n2194 GND.n1609 0.04025
R3397 GND.n2198 GND.n1609 0.04025
R3398 GND.n2199 GND.n2198 0.04025
R3399 GND.n2200 GND.n2199 0.04025
R3400 GND.n2200 GND.n1607 0.04025
R3401 GND.n2204 GND.n1607 0.04025
R3402 GND.n2205 GND.n2204 0.04025
R3403 GND.n2206 GND.n2205 0.04025
R3404 GND.n2206 GND.n1605 0.04025
R3405 GND.n2210 GND.n1605 0.04025
R3406 GND.n2211 GND.n2210 0.04025
R3407 GND.n2212 GND.n2211 0.04025
R3408 GND.n2212 GND.n1603 0.04025
R3409 GND.n2216 GND.n1603 0.04025
R3410 GND.n2217 GND.n2216 0.04025
R3411 GND.n2218 GND.n2217 0.04025
R3412 GND.n2218 GND.n1601 0.04025
R3413 GND.n2222 GND.n1601 0.04025
R3414 GND.n2223 GND.n2222 0.04025
R3415 GND.n2224 GND.n2223 0.04025
R3416 GND.n2224 GND.n1599 0.04025
R3417 GND.n2228 GND.n1599 0.04025
R3418 GND.n2229 GND.n2228 0.04025
R3419 GND.n2230 GND.n2229 0.04025
R3420 GND.n2230 GND.n1597 0.04025
R3421 GND.n2234 GND.n1597 0.04025
R3422 GND.n2235 GND.n2234 0.04025
R3423 GND.n2236 GND.n2235 0.04025
R3424 GND.n2236 GND.n1595 0.04025
R3425 GND.n2240 GND.n1595 0.04025
R3426 GND.n2241 GND.n2240 0.04025
R3427 GND.n2242 GND.n2241 0.04025
R3428 GND.n2242 GND.n1593 0.04025
R3429 GND.n2246 GND.n1593 0.04025
R3430 GND.n2247 GND.n2246 0.04025
R3431 GND.n2248 GND.n2247 0.04025
R3432 GND.n2248 GND.n1591 0.04025
R3433 GND.n2252 GND.n1591 0.04025
R3434 GND.n2253 GND.n2252 0.04025
R3435 GND.n2254 GND.n2253 0.04025
R3436 GND.n2254 GND.n1589 0.04025
R3437 GND.n2258 GND.n1589 0.04025
R3438 GND.n2259 GND.n2258 0.04025
R3439 GND.n2260 GND.n2259 0.04025
R3440 GND.n2260 GND.n1587 0.04025
R3441 GND.n2264 GND.n1587 0.04025
R3442 GND.n2265 GND.n2264 0.04025
R3443 GND.n2266 GND.n2265 0.04025
R3444 GND.n2266 GND.n1585 0.04025
R3445 GND.n2270 GND.n1585 0.04025
R3446 GND.n2271 GND.n2270 0.04025
R3447 GND.n2272 GND.n2271 0.04025
R3448 GND.n2272 GND.n1583 0.04025
R3449 GND.n2276 GND.n1583 0.04025
R3450 GND.n2277 GND.n2276 0.04025
R3451 GND.n2278 GND.n2277 0.04025
R3452 GND.n2278 GND.n1581 0.04025
R3453 GND.n2282 GND.n1581 0.04025
R3454 GND.n2283 GND.n2282 0.04025
R3455 GND.n2284 GND.n2283 0.04025
R3456 GND.n2284 GND.n1579 0.04025
R3457 GND.n2288 GND.n1579 0.04025
R3458 GND.n2289 GND.n2288 0.04025
R3459 GND.n2290 GND.n2289 0.04025
R3460 GND.n2290 GND.n1577 0.04025
R3461 GND.n2294 GND.n1577 0.04025
R3462 GND.n2295 GND.n2294 0.04025
R3463 GND.n2296 GND.n2295 0.04025
R3464 GND.n2296 GND.n1575 0.04025
R3465 GND.n2300 GND.n1575 0.04025
R3466 GND.n2301 GND.n2300 0.04025
R3467 GND.n2302 GND.n2301 0.04025
R3468 GND.n2302 GND.n1573 0.04025
R3469 GND.n2306 GND.n1573 0.04025
R3470 GND.n2307 GND.n2306 0.04025
R3471 GND.n2308 GND.n2307 0.04025
R3472 GND.n2308 GND.n1571 0.04025
R3473 GND.n2312 GND.n1571 0.04025
R3474 GND.n2313 GND.n2312 0.04025
R3475 GND.n2314 GND.n2313 0.04025
R3476 GND.n2314 GND.n1569 0.04025
R3477 GND.n2318 GND.n1569 0.04025
R3478 GND.n2319 GND.n2318 0.04025
R3479 GND.n2320 GND.n2319 0.04025
R3480 GND.n2320 GND.n1567 0.04025
R3481 GND.n2324 GND.n1567 0.04025
R3482 GND.n2325 GND.n2324 0.04025
R3483 GND.n2326 GND.n2325 0.04025
R3484 GND.n2326 GND.n1565 0.04025
R3485 GND.n2330 GND.n1565 0.04025
R3486 GND.n2331 GND.n2330 0.04025
R3487 GND.n2332 GND.n2331 0.04025
R3488 GND.n2332 GND.n1563 0.04025
R3489 GND.n2336 GND.n1563 0.04025
R3490 GND.n2337 GND.n2336 0.04025
R3491 GND.n2338 GND.n2337 0.04025
R3492 GND.n2338 GND.n1561 0.04025
R3493 GND.n2342 GND.n1561 0.04025
R3494 GND.n2343 GND.n2342 0.04025
R3495 GND.n2344 GND.n2343 0.04025
R3496 GND.n2344 GND.n1559 0.04025
R3497 GND.n2348 GND.n1559 0.04025
R3498 GND.n2349 GND.n2348 0.04025
R3499 GND.n2350 GND.n2349 0.04025
R3500 GND.n2350 GND.n1557 0.04025
R3501 GND.n2354 GND.n1557 0.04025
R3502 GND.n2355 GND.n2354 0.04025
R3503 GND.n2356 GND.n2355 0.04025
R3504 GND.n2356 GND.n1555 0.04025
R3505 GND.n2360 GND.n1555 0.04025
R3506 GND.n2361 GND.n2360 0.04025
R3507 GND.n2362 GND.n2361 0.04025
R3508 GND.n2362 GND.n1553 0.04025
R3509 GND.n2366 GND.n1553 0.04025
R3510 GND.n2367 GND.n2366 0.04025
R3511 GND.n2368 GND.n2367 0.04025
R3512 GND.n2368 GND.n1551 0.04025
R3513 GND.n2372 GND.n1551 0.04025
R3514 GND.n2373 GND.n2372 0.04025
R3515 GND.n2374 GND.n2373 0.04025
R3516 GND.n2374 GND.n1549 0.04025
R3517 GND.n2378 GND.n1549 0.04025
R3518 GND.n2379 GND.n2378 0.04025
R3519 GND.n2380 GND.n2379 0.04025
R3520 GND.n2380 GND.n1547 0.04025
R3521 GND.n2384 GND.n1547 0.04025
R3522 GND.n2385 GND.n2384 0.04025
R3523 GND.n2386 GND.n2385 0.04025
R3524 GND.n2386 GND.n1545 0.04025
R3525 GND.n2390 GND.n1545 0.04025
R3526 GND.n2391 GND.n2390 0.04025
R3527 GND.n2392 GND.n2391 0.04025
R3528 GND.n2392 GND.n1543 0.04025
R3529 GND.n2396 GND.n1543 0.04025
R3530 GND.n2397 GND.n2396 0.04025
R3531 GND.n2398 GND.n2397 0.04025
R3532 GND.n2398 GND.n1541 0.04025
R3533 GND.n2402 GND.n1541 0.04025
R3534 GND.n2403 GND.n2402 0.04025
R3535 GND.n2404 GND.n2403 0.04025
R3536 GND.n2404 GND.n1539 0.04025
R3537 GND.n2408 GND.n1539 0.04025
R3538 GND.n2409 GND.n2408 0.04025
R3539 GND.n2410 GND.n2409 0.04025
R3540 GND.n2410 GND.n1537 0.04025
R3541 GND.n2414 GND.n1537 0.04025
R3542 GND.n2415 GND.n2414 0.04025
R3543 GND.n2416 GND.n2415 0.04025
R3544 GND.n2416 GND.n1535 0.04025
R3545 GND.n2420 GND.n1535 0.04025
R3546 GND.n2421 GND.n2420 0.04025
R3547 GND.n2422 GND.n2421 0.04025
R3548 GND.n2422 GND.n1533 0.04025
R3549 GND.n2426 GND.n1533 0.04025
R3550 GND.n2427 GND.n2426 0.04025
R3551 GND.n2428 GND.n2427 0.04025
R3552 GND.n2428 GND.n1531 0.04025
R3553 GND.n2432 GND.n1531 0.04025
R3554 GND.n2433 GND.n2432 0.04025
R3555 GND.n2434 GND.n2433 0.04025
R3556 GND.n2434 GND.n1529 0.04025
R3557 GND.n2438 GND.n1529 0.04025
R3558 GND.n2439 GND.n2438 0.04025
R3559 GND.n2440 GND.n2439 0.04025
R3560 GND.n2440 GND.n1527 0.04025
R3561 GND.n2444 GND.n1527 0.04025
R3562 GND.n2445 GND.n2444 0.04025
R3563 GND.n2446 GND.n2445 0.04025
R3564 GND.n2446 GND.n1525 0.04025
R3565 GND.n2450 GND.n1525 0.04025
R3566 GND.n2451 GND.n2450 0.04025
R3567 GND.n2452 GND.n2451 0.04025
R3568 GND.n2452 GND.n1523 0.04025
R3569 GND.n2456 GND.n1523 0.04025
R3570 GND.n2457 GND.n2456 0.04025
R3571 GND.n2458 GND.n2457 0.04025
R3572 GND.n2458 GND.n1521 0.04025
R3573 GND.n2462 GND.n1521 0.04025
R3574 GND.n2463 GND.n2462 0.04025
R3575 GND.n2464 GND.n2463 0.04025
R3576 GND.n2464 GND.n1519 0.04025
R3577 GND.n2468 GND.n1519 0.04025
R3578 GND.n2469 GND.n2468 0.04025
R3579 GND.n2470 GND.n2469 0.04025
R3580 GND.n2470 GND.n1517 0.04025
R3581 GND.n2474 GND.n1517 0.04025
R3582 GND.n2475 GND.n2474 0.04025
R3583 GND.n2476 GND.n2475 0.04025
R3584 GND.n2476 GND.n1515 0.04025
R3585 GND.n2480 GND.n1515 0.04025
R3586 GND.n2481 GND.n2480 0.04025
R3587 GND.n2482 GND.n2481 0.04025
R3588 GND.n2482 GND.n1513 0.04025
R3589 GND.n2486 GND.n1513 0.04025
R3590 GND.n2487 GND.n2486 0.04025
R3591 GND.n2488 GND.n2487 0.04025
R3592 GND.n2488 GND.n1511 0.04025
R3593 GND.n2492 GND.n1511 0.04025
R3594 GND.n2493 GND.n2492 0.04025
R3595 GND.n2494 GND.n2493 0.04025
R3596 GND.n2494 GND.n1509 0.04025
R3597 GND.n2498 GND.n1509 0.04025
R3598 GND.n2500 GND.n1507 0.04025
R3599 GND.n2504 GND.n1507 0.04025
R3600 GND.n2505 GND.n2504 0.04025
R3601 GND.n2506 GND.n2505 0.04025
R3602 GND.n2506 GND.n1505 0.04025
R3603 GND.n2510 GND.n1505 0.04025
R3604 GND.n2511 GND.n2510 0.04025
R3605 GND.n2512 GND.n2511 0.04025
R3606 GND.n2512 GND.n1503 0.04025
R3607 GND.n2516 GND.n1503 0.04025
R3608 GND.n2517 GND.n2516 0.04025
R3609 GND.n2518 GND.n2517 0.04025
R3610 GND.n2518 GND.n1501 0.04025
R3611 GND.n2522 GND.n1501 0.04025
R3612 GND.n2523 GND.n2522 0.04025
R3613 GND.n2524 GND.n2523 0.04025
R3614 GND.n2524 GND.n1499 0.04025
R3615 GND.n2528 GND.n1499 0.04025
R3616 GND.n2529 GND.n2528 0.04025
R3617 GND.n2530 GND.n2529 0.04025
R3618 GND.n2530 GND.n1497 0.04025
R3619 GND.n2534 GND.n1497 0.04025
R3620 GND.n2535 GND.n2534 0.04025
R3621 GND.n2536 GND.n2535 0.04025
R3622 GND.n2536 GND.n1495 0.04025
R3623 GND.n2540 GND.n1495 0.04025
R3624 GND.n2541 GND.n2540 0.04025
R3625 GND.n2542 GND.n2541 0.04025
R3626 GND.n2542 GND.n1493 0.04025
R3627 GND.n2546 GND.n1493 0.04025
R3628 GND.n2547 GND.n2546 0.04025
R3629 GND.n2548 GND.n2547 0.04025
R3630 GND.n2548 GND.n1491 0.04025
R3631 GND.n2552 GND.n1491 0.04025
R3632 GND.n2553 GND.n2552 0.04025
R3633 GND.n2554 GND.n2553 0.04025
R3634 GND.n2554 GND.n1489 0.04025
R3635 GND.n2558 GND.n1489 0.04025
R3636 GND.n2559 GND.n2558 0.04025
R3637 GND.n2560 GND.n2559 0.04025
R3638 GND.n2560 GND.n1487 0.04025
R3639 GND.n2564 GND.n1487 0.04025
R3640 GND.n2565 GND.n2564 0.04025
R3641 GND.n2566 GND.n2565 0.04025
R3642 GND.n2566 GND.n1485 0.04025
R3643 GND.n2570 GND.n1485 0.04025
R3644 GND.n2571 GND.n2570 0.04025
R3645 GND.n2572 GND.n2571 0.04025
R3646 GND.n2572 GND.n1483 0.04025
R3647 GND.n2576 GND.n1483 0.04025
R3648 GND.n2577 GND.n2576 0.04025
R3649 GND.n2578 GND.n2577 0.04025
R3650 GND.n2578 GND.n1481 0.04025
R3651 GND.n2582 GND.n1481 0.04025
R3652 GND.n2583 GND.n2582 0.04025
R3653 GND.n2584 GND.n2583 0.04025
R3654 GND.n2584 GND.n1479 0.04025
R3655 GND.n2588 GND.n1479 0.04025
R3656 GND.n2589 GND.n2588 0.04025
R3657 GND.n2590 GND.n2589 0.04025
R3658 GND.n2590 GND.n1477 0.04025
R3659 GND.n2594 GND.n1477 0.04025
R3660 GND.n2595 GND.n2594 0.04025
R3661 GND.n2596 GND.n2595 0.04025
R3662 GND.n2596 GND.n1475 0.04025
R3663 GND.n2600 GND.n1475 0.04025
R3664 GND.n2601 GND.n2600 0.04025
R3665 GND.n2602 GND.n2601 0.04025
R3666 GND.n2602 GND.n1473 0.04025
R3667 GND.n2606 GND.n1473 0.04025
R3668 GND.n2607 GND.n2606 0.04025
R3669 GND.n2608 GND.n2607 0.04025
R3670 GND.n2608 GND.n1471 0.04025
R3671 GND.n2612 GND.n1471 0.04025
R3672 GND.n2613 GND.n2612 0.04025
R3673 GND.n2614 GND.n2613 0.04025
R3674 GND.n2614 GND.n1469 0.04025
R3675 GND.n2618 GND.n1469 0.04025
R3676 GND.n2619 GND.n2618 0.04025
R3677 GND.n2620 GND.n2619 0.04025
R3678 GND.n2620 GND.n1467 0.04025
R3679 GND.n2624 GND.n1467 0.04025
R3680 GND.n2625 GND.n2624 0.04025
R3681 GND.n2626 GND.n2625 0.04025
R3682 GND.n2626 GND.n1465 0.04025
R3683 GND.n2630 GND.n1465 0.04025
R3684 GND.n2631 GND.n2630 0.04025
R3685 GND.n2632 GND.n2631 0.04025
R3686 GND.n2632 GND.n1463 0.04025
R3687 GND.n2636 GND.n1463 0.04025
R3688 GND.n2637 GND.n2636 0.04025
R3689 GND.n2638 GND.n2637 0.04025
R3690 GND.n2638 GND.n1461 0.04025
R3691 GND.n2642 GND.n1461 0.04025
R3692 GND.n2643 GND.n2642 0.04025
R3693 GND.n2644 GND.n2643 0.04025
R3694 GND.n2644 GND.n1459 0.04025
R3695 GND.n2648 GND.n1459 0.04025
R3696 GND.n2649 GND.n2648 0.04025
R3697 GND.n2650 GND.n2649 0.04025
R3698 GND.n2650 GND.n1457 0.04025
R3699 GND.n2654 GND.n1457 0.04025
R3700 GND.n2655 GND.n2654 0.04025
R3701 GND.n2656 GND.n2655 0.04025
R3702 GND.n2656 GND.n1455 0.04025
R3703 GND.n2660 GND.n1455 0.04025
R3704 GND.n2661 GND.n2660 0.04025
R3705 GND.n2662 GND.n2661 0.04025
R3706 GND.n2662 GND.n1453 0.04025
R3707 GND.n2666 GND.n1453 0.04025
R3708 GND.n2667 GND.n2666 0.04025
R3709 GND.n2668 GND.n2667 0.04025
R3710 GND.n2668 GND.n1451 0.04025
R3711 GND.n2672 GND.n1451 0.04025
R3712 GND.n2673 GND.n2672 0.04025
R3713 GND.n2674 GND.n2673 0.04025
R3714 GND.n2674 GND.n1449 0.04025
R3715 GND.n2678 GND.n1449 0.04025
R3716 GND.n2679 GND.n2678 0.04025
R3717 GND.n2950 GND.n2679 0.04025
R3718 GND.n2950 GND.n2949 0.04025
R3719 GND.n2949 GND.n2948 0.04025
R3720 GND.n2948 GND.n2680 0.04025
R3721 GND.n2944 GND.n2680 0.04025
R3722 GND.n2944 GND.n2943 0.04025
R3723 GND.n2943 GND.n2942 0.04025
R3724 GND.n2942 GND.n2682 0.04025
R3725 GND.n2938 GND.n2682 0.04025
R3726 GND.n2938 GND.n2937 0.04025
R3727 GND.n2937 GND.n2936 0.04025
R3728 GND.n2936 GND.n2684 0.04025
R3729 GND.n2932 GND.n2684 0.04025
R3730 GND.n2932 GND.n2931 0.04025
R3731 GND.n2931 GND.n2930 0.04025
R3732 GND.n2930 GND.n2686 0.04025
R3733 GND.n2926 GND.n2686 0.04025
R3734 GND.n2926 GND.n2925 0.04025
R3735 GND.n2925 GND.n2924 0.04025
R3736 GND.n2924 GND.n2688 0.04025
R3737 GND.n2920 GND.n2688 0.04025
R3738 GND.n2920 GND.n2919 0.04025
R3739 GND.n2919 GND.n2918 0.04025
R3740 GND.n2918 GND.n2690 0.04025
R3741 GND.n2914 GND.n2690 0.04025
R3742 GND.n2914 GND.n2913 0.04025
R3743 GND.n2913 GND.n2912 0.04025
R3744 GND.n2912 GND.n2692 0.04025
R3745 GND.n2908 GND.n2692 0.04025
R3746 GND.n2908 GND.n2907 0.04025
R3747 GND.n2907 GND.n2906 0.04025
R3748 GND.n2906 GND.n2694 0.04025
R3749 GND.n2902 GND.n2694 0.04025
R3750 GND.n2902 GND.n2901 0.04025
R3751 GND.n2901 GND.n2900 0.04025
R3752 GND.n2900 GND.n2696 0.04025
R3753 GND.n2896 GND.n2696 0.04025
R3754 GND.n2896 GND.n2895 0.04025
R3755 GND.n2895 GND.n2894 0.04025
R3756 GND.n2894 GND.n2698 0.04025
R3757 GND.n2890 GND.n2698 0.04025
R3758 GND.n2890 GND.n2889 0.04025
R3759 GND.n2889 GND.n2888 0.04025
R3760 GND.n2888 GND.n2700 0.04025
R3761 GND.n2884 GND.n2700 0.04025
R3762 GND.n2884 GND.n2883 0.04025
R3763 GND.n2883 GND.n2882 0.04025
R3764 GND.n2882 GND.n2702 0.04025
R3765 GND.n2878 GND.n2702 0.04025
R3766 GND.n2878 GND.n2877 0.04025
R3767 GND.n2877 GND.n2876 0.04025
R3768 GND.n2876 GND.n2704 0.04025
R3769 GND.n2872 GND.n2704 0.04025
R3770 GND.n2872 GND.n2871 0.04025
R3771 GND.n2871 GND.n2870 0.04025
R3772 GND.n2870 GND.n2706 0.04025
R3773 GND.n2866 GND.n2706 0.04025
R3774 GND.n2866 GND.n2865 0.04025
R3775 GND.n2865 GND.n2864 0.04025
R3776 GND.n2864 GND.n2708 0.04025
R3777 GND.n2860 GND.n2708 0.04025
R3778 GND.n2860 GND.n2859 0.04025
R3779 GND.n2859 GND.n2858 0.04025
R3780 GND.n2858 GND.n2710 0.04025
R3781 GND.n2854 GND.n2710 0.04025
R3782 GND.n2854 GND.n2853 0.04025
R3783 GND.n2853 GND.n2852 0.04025
R3784 GND.n2852 GND.n2712 0.04025
R3785 GND.n2848 GND.n2712 0.04025
R3786 GND.n2848 GND.n2847 0.04025
R3787 GND.n2847 GND.n2846 0.04025
R3788 GND.n2846 GND.n2714 0.04025
R3789 GND.n2842 GND.n2714 0.04025
R3790 GND.n2842 GND.n2841 0.04025
R3791 GND.n2841 GND.n2840 0.04025
R3792 GND.n2840 GND.n2716 0.04025
R3793 GND.n2836 GND.n2716 0.04025
R3794 GND.n2836 GND.n2835 0.04025
R3795 GND.n2835 GND.n2834 0.04025
R3796 GND.n2834 GND.n2718 0.04025
R3797 GND.n2830 GND.n2718 0.04025
R3798 GND.n2830 GND.n2829 0.04025
R3799 GND.n2829 GND.n2828 0.04025
R3800 GND.n2828 GND.n2720 0.04025
R3801 GND.n2824 GND.n2720 0.04025
R3802 GND.n2824 GND.n2823 0.04025
R3803 GND.n2823 GND.n2822 0.04025
R3804 GND.n2822 GND.n2722 0.04025
R3805 GND.n2818 GND.n2722 0.04025
R3806 GND.n2818 GND.n2817 0.04025
R3807 GND.n2817 GND.n2816 0.04025
R3808 GND.n2816 GND.n2724 0.04025
R3809 GND.n2812 GND.n2724 0.04025
R3810 GND.n2812 GND.n2811 0.04025
R3811 GND.n2811 GND.n2810 0.04025
R3812 GND.n2810 GND.n2726 0.04025
R3813 GND.n2806 GND.n2726 0.04025
R3814 GND.n2806 GND.n2805 0.04025
R3815 GND.n2805 GND.n2804 0.04025
R3816 GND.n2804 GND.n2728 0.04025
R3817 GND.n2800 GND.n2728 0.04025
R3818 GND.n2800 GND.n2799 0.04025
R3819 GND.n2799 GND.n2798 0.04025
R3820 GND.n2798 GND.n2730 0.04025
R3821 GND.n2794 GND.n2730 0.04025
R3822 GND.n2794 GND.n2793 0.04025
R3823 GND.n2793 GND.n2792 0.04025
R3824 GND.n2792 GND.n2732 0.04025
R3825 GND.n2788 GND.n2732 0.04025
R3826 GND.n2788 GND.n2787 0.04025
R3827 GND.n2787 GND.n2786 0.04025
R3828 GND.n2786 GND.n2734 0.04025
R3829 GND.n2782 GND.n2734 0.04025
R3830 GND.n2782 GND.n2781 0.04025
R3831 GND.n2781 GND.n2780 0.04025
R3832 GND.n2780 GND.n2736 0.04025
R3833 GND.n2776 GND.n2736 0.04025
R3834 GND.n2776 GND.n2775 0.04025
R3835 GND.n2775 GND.n2774 0.04025
R3836 GND.n2774 GND.n2738 0.04025
R3837 GND.n2770 GND.n2738 0.04025
R3838 GND.n1943 GND.n1699 0.04025
R3839 GND.n1944 GND.n1943 0.04025
R3840 GND.n1945 GND.n1944 0.04025
R3841 GND.n1945 GND.n1697 0.04025
R3842 GND.n1949 GND.n1697 0.04025
R3843 GND.n1950 GND.n1949 0.04025
R3844 GND.n1951 GND.n1950 0.04025
R3845 GND.n1951 GND.n1695 0.04025
R3846 GND.n1955 GND.n1695 0.04025
R3847 GND.n1956 GND.n1955 0.04025
R3848 GND.n1957 GND.n1956 0.04025
R3849 GND.n1957 GND.n1693 0.04025
R3850 GND.n1961 GND.n1693 0.04025
R3851 GND.n1962 GND.n1961 0.04025
R3852 GND.n1963 GND.n1962 0.04025
R3853 GND.n1963 GND.n1691 0.04025
R3854 GND.n1967 GND.n1691 0.04025
R3855 GND.n1968 GND.n1967 0.04025
R3856 GND.n1969 GND.n1968 0.04025
R3857 GND.n1969 GND.n1689 0.04025
R3858 GND.n1973 GND.n1689 0.04025
R3859 GND.n1974 GND.n1973 0.04025
R3860 GND.n2958 GND.n2957 0.04025
R3861 GND.n2958 GND.n1441 0.04025
R3862 GND.n2962 GND.n1441 0.04025
R3863 GND.n2963 GND.n2962 0.04025
R3864 GND.n2964 GND.n2963 0.04025
R3865 GND.n2964 GND.n1439 0.04025
R3866 GND.n2968 GND.n1439 0.04025
R3867 GND.n2969 GND.n2968 0.04025
R3868 GND.n2970 GND.n2969 0.04025
R3869 GND.n2970 GND.n1437 0.04025
R3870 GND.n2974 GND.n1437 0.04025
R3871 GND.n2975 GND.n2974 0.04025
R3872 GND.n2976 GND.n2975 0.04025
R3873 GND.n2976 GND.n1435 0.04025
R3874 GND.n2980 GND.n1435 0.04025
R3875 GND.n2981 GND.n2980 0.04025
R3876 GND.n2982 GND.n2981 0.04025
R3877 GND.n2982 GND.n1433 0.04025
R3878 GND.n2986 GND.n1433 0.04025
R3879 GND.n2987 GND.n2986 0.04025
R3880 GND.n2988 GND.n2987 0.04025
R3881 GND.n2988 GND.n1431 0.04025
R3882 GND.n2992 GND.n1431 0.04025
R3883 GND.n2993 GND.n2992 0.04025
R3884 GND.n2994 GND.n2993 0.04025
R3885 GND.n2994 GND.n1429 0.04025
R3886 GND.n2998 GND.n1429 0.04025
R3887 GND.n2999 GND.n2998 0.04025
R3888 GND.n3000 GND.n2999 0.04025
R3889 GND.n3000 GND.n1427 0.04025
R3890 GND.n3004 GND.n1427 0.04025
R3891 GND.n3005 GND.n3004 0.04025
R3892 GND.n3006 GND.n3005 0.04025
R3893 GND.n3006 GND.n1425 0.04025
R3894 GND.n3010 GND.n1425 0.04025
R3895 GND.n3011 GND.n3010 0.04025
R3896 GND.n3012 GND.n3011 0.04025
R3897 GND.n3012 GND.n1423 0.04025
R3898 GND.n3016 GND.n1423 0.04025
R3899 GND.n3017 GND.n3016 0.04025
R3900 GND.n3018 GND.n3017 0.04025
R3901 GND.n3018 GND.n1421 0.04025
R3902 GND.n3022 GND.n1421 0.04025
R3903 GND.n3023 GND.n3022 0.04025
R3904 GND.n3024 GND.n3023 0.04025
R3905 GND.n2747 GND.n1419 0.04025
R3906 GND.n2749 GND.n2747 0.04025
R3907 GND.n2750 GND.n2749 0.04025
R3908 GND.n2751 GND.n2750 0.04025
R3909 GND.n2751 GND.n2745 0.04025
R3910 GND.n2755 GND.n2745 0.04025
R3911 GND.n2756 GND.n2755 0.04025
R3912 GND.n2757 GND.n2756 0.04025
R3913 GND.n2757 GND.n2743 0.04025
R3914 GND.n2761 GND.n2743 0.04025
R3915 GND.n2762 GND.n2761 0.04025
R3916 GND.n2763 GND.n2762 0.04025
R3917 GND.n2763 GND.n2741 0.04025
R3918 GND.n2767 GND.n2741 0.04025
R3919 GND.n2959 GND.n1442 0.04025
R3920 GND.n2960 GND.n2959 0.04025
R3921 GND.n2961 GND.n2960 0.04025
R3922 GND.n2961 GND.n1440 0.04025
R3923 GND.n2965 GND.n1440 0.04025
R3924 GND.n2966 GND.n2965 0.04025
R3925 GND.n2967 GND.n2966 0.04025
R3926 GND.n2967 GND.n1438 0.04025
R3927 GND.n2971 GND.n1438 0.04025
R3928 GND.n2972 GND.n2971 0.04025
R3929 GND.n2973 GND.n2972 0.04025
R3930 GND.n2973 GND.n1436 0.04025
R3931 GND.n2977 GND.n1436 0.04025
R3932 GND.n2978 GND.n2977 0.04025
R3933 GND.n2979 GND.n2978 0.04025
R3934 GND.n2979 GND.n1434 0.04025
R3935 GND.n2983 GND.n1434 0.04025
R3936 GND.n2984 GND.n2983 0.04025
R3937 GND.n2985 GND.n2984 0.04025
R3938 GND.n2985 GND.n1432 0.04025
R3939 GND.n2989 GND.n1432 0.04025
R3940 GND.n2990 GND.n2989 0.04025
R3941 GND.n2991 GND.n2990 0.04025
R3942 GND.n2991 GND.n1430 0.04025
R3943 GND.n2995 GND.n1430 0.04025
R3944 GND.n2996 GND.n2995 0.04025
R3945 GND.n2997 GND.n2996 0.04025
R3946 GND.n2997 GND.n1428 0.04025
R3947 GND.n3001 GND.n1428 0.04025
R3948 GND.n3002 GND.n3001 0.04025
R3949 GND.n3003 GND.n3002 0.04025
R3950 GND.n3003 GND.n1426 0.04025
R3951 GND.n3007 GND.n1426 0.04025
R3952 GND.n3008 GND.n3007 0.04025
R3953 GND.n3009 GND.n3008 0.04025
R3954 GND.n3009 GND.n1424 0.04025
R3955 GND.n3013 GND.n1424 0.04025
R3956 GND.n3014 GND.n3013 0.04025
R3957 GND.n3015 GND.n3014 0.04025
R3958 GND.n3015 GND.n1422 0.04025
R3959 GND.n3019 GND.n1422 0.04025
R3960 GND.n3020 GND.n3019 0.04025
R3961 GND.n3021 GND.n3020 0.04025
R3962 GND.n3021 GND.n1417 0.04025
R3963 GND.n2748 GND.n1418 0.04025
R3964 GND.n2748 GND.n2746 0.04025
R3965 GND.n2752 GND.n2746 0.04025
R3966 GND.n2753 GND.n2752 0.04025
R3967 GND.n2754 GND.n2753 0.04025
R3968 GND.n2754 GND.n2744 0.04025
R3969 GND.n2758 GND.n2744 0.04025
R3970 GND.n2759 GND.n2758 0.04025
R3971 GND.n2760 GND.n2759 0.04025
R3972 GND.n2760 GND.n2742 0.04025
R3973 GND.n2764 GND.n2742 0.04025
R3974 GND.n2765 GND.n2764 0.04025
R3975 GND.n2766 GND.n2765 0.04025
R3976 GND.n1330 GND.n45 0.0381165
R3977 GND.n800 GND.n799 0.0358501
R3978 GND.n803 GND.n802 0.0358501
R3979 GND.n806 GND.n805 0.0358501
R3980 GND.n571 GND.n570 0.0358501
R3981 GND.n219 GND.n218 0.0358501
R3982 GND.n396 GND.n395 0.0358501
R3983 GND.n394 GND.n393 0.0358501
R3984 GND.n392 GND.n391 0.0358501
R3985 GND.n282 GND.n281 0.03425
R3986 GND.n266 GND.n265 0.0324737
R3987 GND.n575 GND.n574 0.0323341
R3988 GND.n577 GND.n576 0.0323341
R3989 GND.n579 GND.n578 0.0323341
R3990 GND.n811 GND.n810 0.0323341
R3991 GND.n813 GND.n812 0.0323341
R3992 GND.n815 GND.n814 0.0323341
R3993 GND.n210 GND.n209 0.0323341
R3994 GND.n212 GND.n211 0.0323341
R3995 GND.n214 GND.n213 0.0323341
R3996 GND.n384 GND.n383 0.0323341
R3997 GND.n386 GND.n385 0.0323341
R3998 GND.n388 GND.n387 0.0323341
R3999 GND.n1332 GND.n1331 0.0322143
R4000 GND.n1345 GND.n38 0.032139
R4001 GND.n1346 GND.n38 0.032139
R4002 GND.n1361 GND.n28 0.032139
R4003 GND.n1362 GND.n28 0.032139
R4004 GND.n1363 GND.n27 0.032139
R4005 GND.n1364 GND.n27 0.032139
R4006 GND.n1365 GND.n26 0.032139
R4007 GND.n1366 GND.n26 0.032139
R4008 GND.n1367 GND.n25 0.032139
R4009 GND.n1368 GND.n25 0.032139
R4010 GND.n1369 GND.n24 0.032139
R4011 GND.n1370 GND.n24 0.032139
R4012 GND.n1371 GND.n23 0.032139
R4013 GND.n1372 GND.n23 0.032139
R4014 GND.n1325 GND.n49 0.032139
R4015 GND.n1324 GND.n49 0.032139
R4016 GND.n1298 GND.n57 0.0320266
R4017 GND.n1297 GND.n57 0.0320266
R4018 GND.n1296 GND.n58 0.0320266
R4019 GND.n1295 GND.n58 0.0320266
R4020 GND.n1294 GND.n59 0.0320266
R4021 GND.n1293 GND.n59 0.0320266
R4022 GND.n1292 GND.n60 0.0320266
R4023 GND.n1291 GND.n60 0.0320266
R4024 GND.n1290 GND.n61 0.0320266
R4025 GND.n1289 GND.n61 0.0320266
R4026 GND.n1288 GND.n62 0.0320266
R4027 GND.n1287 GND.n62 0.0320266
R4028 GND.n1334 GND.n43 0.0318433
R4029 GND.n1335 GND.n43 0.0318433
R4030 GND.n1336 GND.n1335 0.0318433
R4031 GND.n1336 GND.n42 0.0318433
R4032 GND.n1337 GND.n42 0.0318433
R4033 GND.n1304 GND.n54 0.0318433
R4034 GND.n1305 GND.n54 0.0318433
R4035 GND.n1306 GND.n1305 0.0318433
R4036 GND.n1306 GND.n53 0.0318433
R4037 GND.n1307 GND.n53 0.0318433
R4038 GND.n1308 GND.n1307 0.0318433
R4039 GND.n1308 GND.n52 0.0318433
R4040 GND.n1309 GND.n52 0.0318433
R4041 GND.n1310 GND.n1309 0.0318433
R4042 GND.n1310 GND.n51 0.0318433
R4043 GND.n1311 GND.n51 0.0318433
R4044 GND.n265 GND.n252 0.0312895
R4045 GND.n1359 GND.n29 0.0296667
R4046 GND.n1348 GND.n37 0.0296329
R4047 GND.n1322 GND.n1321 0.0296329
R4048 GND.n1363 GND.n1362 0.0295736
R4049 GND.n1365 GND.n1364 0.0295736
R4050 GND.n1367 GND.n1366 0.0295736
R4051 GND.n1369 GND.n1368 0.0295736
R4052 GND.n1371 GND.n1370 0.0295736
R4053 GND.n281 GND.n280 0.0295132
R4054 GND.n1297 GND.n1296 0.0294704
R4055 GND.n1295 GND.n1294 0.0294704
R4056 GND.n1293 GND.n1292 0.0294704
R4057 GND.n1291 GND.n1290 0.0294704
R4058 GND.n1289 GND.n1288 0.0294704
R4059 GND.n496 GND.n452 0.0284
R4060 GND.n497 GND.n451 0.0284
R4061 GND.n3026 GND.n1418 0.027875
R4062 GND.n1334 GND.n1333 0.0275896
R4063 GND.n1338 GND.n1337 0.0274776
R4064 GND.n1304 GND.n1303 0.0274776
R4065 GND.n1373 GND.n1372 0.027385
R4066 GND.n1326 GND.n1325 0.0273316
R4067 GND.n1287 GND.n1286 0.0272974
R4068 GND.n1345 GND.n1344 0.0272769
R4069 GND.n1299 GND.n1298 0.027243
R4070 GND.n1333 GND.n44 0.0253571
R4071 GND.n1361 GND.n1360 0.0250843
R4072 GND.n1347 GND.n1346 0.0249774
R4073 GND.n1324 GND.n1323 0.0249774
R4074 GND.n1354 GND.n31 0.0247529
R4075 GND.n1354 GND.n33 0.0247529
R4076 GND.n501 GND.n500 0.02435
R4077 GND.n504 GND.n501 0.02435
R4078 GND.n505 GND.n504 0.02435
R4079 GND.n506 GND.n505 0.02435
R4080 GND.n506 GND.n174 0.02435
R4081 GND.n510 GND.n174 0.02435
R4082 GND.n511 GND.n510 0.02435
R4083 GND.n512 GND.n511 0.02435
R4084 GND.n512 GND.n172 0.02435
R4085 GND.n516 GND.n172 0.02435
R4086 GND.n517 GND.n516 0.02435
R4087 GND.n518 GND.n517 0.02435
R4088 GND.n518 GND.n170 0.02435
R4089 GND.n522 GND.n170 0.02435
R4090 GND.n523 GND.n522 0.02435
R4091 GND.n524 GND.n523 0.02435
R4092 GND.n524 GND.n168 0.02435
R4093 GND.n528 GND.n168 0.02435
R4094 GND.n529 GND.n528 0.02435
R4095 GND.n530 GND.n529 0.02435
R4096 GND.n530 GND.n166 0.02435
R4097 GND.n534 GND.n166 0.02435
R4098 GND.n535 GND.n534 0.02435
R4099 GND.n536 GND.n535 0.02435
R4100 GND.n536 GND.n164 0.02435
R4101 GND.n540 GND.n164 0.02435
R4102 GND.n541 GND.n540 0.02435
R4103 GND.n542 GND.n541 0.02435
R4104 GND.n542 GND.n162 0.02435
R4105 GND.n546 GND.n162 0.02435
R4106 GND.n547 GND.n546 0.02435
R4107 GND.n548 GND.n547 0.02435
R4108 GND.n548 GND.n160 0.02435
R4109 GND.n837 GND.n836 0.02435
R4110 GND.n838 GND.n837 0.02435
R4111 GND.n838 GND.n82 0.02435
R4112 GND.n842 GND.n82 0.02435
R4113 GND.n843 GND.n842 0.02435
R4114 GND.n844 GND.n843 0.02435
R4115 GND.n844 GND.n80 0.02435
R4116 GND.n1414 GND.n1413 0.02435
R4117 GND.n3028 GND.n1414 0.02435
R4118 GND.n580 GND.n564 0.0237017
R4119 GND.n831 GND.n87 0.0237017
R4120 GND.n382 GND.n231 0.0237017
R4121 GND.n574 GND.n567 0.0236444
R4122 GND.n575 GND.n566 0.0236444
R4123 GND.n576 GND.n566 0.0236444
R4124 GND.n577 GND.n565 0.0236444
R4125 GND.n578 GND.n565 0.0236444
R4126 GND.n579 GND.n153 0.0236444
R4127 GND.n810 GND.n97 0.0236444
R4128 GND.n811 GND.n96 0.0236444
R4129 GND.n812 GND.n96 0.0236444
R4130 GND.n813 GND.n95 0.0236444
R4131 GND.n814 GND.n95 0.0236444
R4132 GND.n816 GND.n815 0.0236444
R4133 GND.n209 GND.n177 0.0236444
R4134 GND.n210 GND.n208 0.0236444
R4135 GND.n211 GND.n208 0.0236444
R4136 GND.n212 GND.n207 0.0236444
R4137 GND.n213 GND.n207 0.0236444
R4138 GND.n214 GND.n206 0.0236444
R4139 GND.n383 GND.n230 0.0236444
R4140 GND.n384 GND.n229 0.0236444
R4141 GND.n385 GND.n229 0.0236444
R4142 GND.n386 GND.n228 0.0236444
R4143 GND.n387 GND.n228 0.0236444
R4144 GND.n388 GND.n227 0.0236444
R4145 GND.n2161 GND.n2160 0.023375
R4146 GND.n2497 GND.n1508 0.023375
R4147 GND.n2162 GND.n1621 0.023375
R4148 GND.n2499 GND.n2498 0.023375
R4149 GND.n798 GND.n797 0.0228491
R4150 GND.n799 GND.n798 0.0228491
R4151 GND.n801 GND.n800 0.0228491
R4152 GND.n802 GND.n801 0.0228491
R4153 GND.n804 GND.n803 0.0228491
R4154 GND.n805 GND.n804 0.0228491
R4155 GND.n807 GND.n806 0.0228491
R4156 GND.n808 GND.n807 0.0228491
R4157 GND.n572 GND.n568 0.0228491
R4158 GND.n571 GND.n568 0.0228491
R4159 GND.n570 GND.n569 0.0228491
R4160 GND.n569 GND.n98 0.0228491
R4161 GND.n217 GND.n216 0.0228491
R4162 GND.n218 GND.n217 0.0228491
R4163 GND.n220 GND.n219 0.0228491
R4164 GND.n221 GND.n220 0.0228491
R4165 GND.n397 GND.n223 0.0228491
R4166 GND.n396 GND.n223 0.0228491
R4167 GND.n395 GND.n224 0.0228491
R4168 GND.n394 GND.n224 0.0228491
R4169 GND.n393 GND.n225 0.0228491
R4170 GND.n392 GND.n225 0.0228491
R4171 GND.n391 GND.n226 0.0228491
R4172 GND.n390 GND.n226 0.0228491
R4173 GND.n797 GND.n796 0.0224016
R4174 GND.n809 GND.n808 0.0224016
R4175 GND.n573 GND.n572 0.0224016
R4176 GND.n796 GND.n98 0.0224016
R4177 GND.n216 GND.n215 0.0224016
R4178 GND.n398 GND.n221 0.0224016
R4179 GND.n398 GND.n397 0.0224016
R4180 GND.n390 GND.n389 0.0224016
R4181 GND.n3026 GND.n1417 0.021875
R4182 GND.n2501 GND.n1508 0.0215
R4183 GND.n2160 GND.n2159 0.0215
R4184 GND.n2158 GND.n1621 0.0215
R4185 GND.n2500 GND.n2499 0.0215
R4186 GND.n1419 GND.n1416 0.0207876
R4187 GND.n3024 GND.n1415 0.0207876
R4188 GND.n2952 GND.n1447 0.020375
R4189 GND.n2952 GND.n2951 0.020375
R4190 GND.n2740 GND.n2739 0.020375
R4191 GND.n1980 GND.n1979 0.020375
R4192 GND.n1979 GND.n1682 0.020375
R4193 GND.n2769 GND.n2768 0.020375
R4194 GND.n2955 GND.n1442 0.020375
R4195 GND.n563 GND.n562 0.01985
R4196 GND.n559 GND.n154 0.01985
R4197 GND.n557 GND.n159 0.01985
R4198 GND.n555 GND.n155 0.01985
R4199 GND.n553 GND.n158 0.01985
R4200 GND.n551 GND.n156 0.01985
R4201 GND.n157 GND.n152 0.01985
R4202 GND.n584 GND.n583 0.01985
R4203 GND.n587 GND.n150 0.01985
R4204 GND.n589 GND.n588 0.01985
R4205 GND.n597 GND.n145 0.01985
R4206 GND.n601 GND.n140 0.01985
R4207 GND.n606 GND.n604 0.01985
R4208 GND.n605 GND.n136 0.01985
R4209 GND.n611 GND.n610 0.01985
R4210 GND.n138 GND.n131 0.01985
R4211 GND.n620 GND.n128 0.01985
R4212 GND.n646 GND.n645 0.01985
R4213 GND.n642 GND.n116 0.01985
R4214 GND.n640 GND.n127 0.01985
R4215 GND.n638 GND.n117 0.01985
R4216 GND.n636 GND.n126 0.01985
R4217 GND.n634 GND.n118 0.01985
R4218 GND.n632 GND.n125 0.01985
R4219 GND.n630 GND.n119 0.01985
R4220 GND.n628 GND.n124 0.01985
R4221 GND.n626 GND.n120 0.01985
R4222 GND.n624 GND.n123 0.01985
R4223 GND.n122 GND.n121 0.01985
R4224 GND.n649 GND.n112 0.01985
R4225 GND.n648 GND.n109 0.01985
R4226 GND.n771 GND.n770 0.01985
R4227 GND.n767 GND.n110 0.01985
R4228 GND.n766 GND.n653 0.01985
R4229 GND.n762 GND.n761 0.01985
R4230 GND.n757 GND.n661 0.01985
R4231 GND.n754 GND.n753 0.01985
R4232 GND.n750 GND.n665 0.01985
R4233 GND.n749 GND.n667 0.01985
R4234 GND.n745 GND.n744 0.01985
R4235 GND.n740 GND.n675 0.01985
R4236 GND.n737 GND.n736 0.01985
R4237 GND.n733 GND.n681 0.01985
R4238 GND.n732 GND.n683 0.01985
R4239 GND.n728 GND.n727 0.01985
R4240 GND.n723 GND.n691 0.01985
R4241 GND.n720 GND.n719 0.01985
R4242 GND.n716 GND.n697 0.01985
R4243 GND.n715 GND.n699 0.01985
R4244 GND.n711 GND.n710 0.01985
R4245 GND.n820 GND.n819 0.01985
R4246 GND.n822 GND.n88 0.01985
R4247 GND.n824 GND.n89 0.01985
R4248 GND.n826 GND.n90 0.01985
R4249 GND.n829 GND.n91 0.01985
R4250 GND.n830 GND.n86 0.01985
R4251 GND.n833 GND.n832 0.01985
R4252 GND.n836 GND.n84 0.01985
R4253 GND.n486 GND.n485 0.0191
R4254 GND.n485 GND.n484 0.0191
R4255 GND.n484 GND.n459 0.0191
R4256 GND.n480 GND.n459 0.0191
R4257 GND.n480 GND.n479 0.0191
R4258 GND.n479 GND.n478 0.0191
R4259 GND.n478 GND.n475 0.0191
R4260 GND.n475 GND.n474 0.0191
R4261 GND.n474 GND.n473 0.0191
R4262 GND.n473 GND.n472 0.0191
R4263 GND.n472 GND.n461 0.0191
R4264 GND.n468 GND.n461 0.0191
R4265 GND.n468 GND.n467 0.0191
R4266 GND.n467 GND.n466 0.0191
R4267 GND.n466 GND.n463 0.0191
R4268 GND.n463 GND.n454 0.0191
R4269 GND.n489 GND.n454 0.0191
R4270 GND.n292 GND.n291 0.0188553
R4271 GND.n310 GND.n309 0.0182632
R4272 GND.n2955 GND.n2954 0.0175455
R4273 GND.n185 GND.n181 0.0164868
R4274 GND.n1373 GND.n22 0.0163383
R4275 GND.n1374 GND.n22 0.0163383
R4276 GND.n1376 GND.n1375 0.0163383
R4277 GND.n1286 GND.n63 0.0163383
R4278 GND.n1285 GND.n63 0.0163383
R4279 GND.n1284 GND.n64 0.0163383
R4280 GND.n339 GND.n338 0.0163383
R4281 GND.n338 GND.n46 0.0163383
R4282 GND.n1329 GND.n47 0.0163383
R4283 GND.n1328 GND.n47 0.0163383
R4284 GND.n1327 GND.n48 0.0163383
R4285 GND.n1326 GND.n48 0.0163383
R4286 GND.n1340 GND.n41 0.0163289
R4287 GND.n1341 GND.n40 0.0163289
R4288 GND.n1342 GND.n40 0.0163289
R4289 GND.n1343 GND.n39 0.0163289
R4290 GND.n1344 GND.n39 0.0163289
R4291 GND.n1302 GND.n1301 0.0163289
R4292 GND.n1300 GND.n56 0.0163289
R4293 GND.n1299 GND.n56 0.0163289
R4294 GND.n581 GND.n580 0.0158898
R4295 GND.n817 GND.n87 0.0158898
R4296 GND.n448 GND.n447 0.0158898
R4297 GND.n382 GND.n381 0.0158898
R4298 GND.n621 GND.n619 0.015575
R4299 GND.n487 GND.n458 0.0151842
R4300 GND.n483 GND.n458 0.0151842
R4301 GND.n483 GND.n482 0.0151842
R4302 GND.n482 GND.n481 0.0151842
R4303 GND.n481 GND.n460 0.0151842
R4304 GND.n477 GND.n460 0.0151842
R4305 GND.n477 GND.n476 0.0151842
R4306 GND.n476 GND.n457 0.0151842
R4307 GND.n471 GND.n456 0.0151842
R4308 GND.n471 GND.n470 0.0151842
R4309 GND.n470 GND.n469 0.0151842
R4310 GND.n469 GND.n462 0.0151842
R4311 GND.n465 GND.n462 0.0151842
R4312 GND.n465 GND.n464 0.0151842
R4313 GND.n464 GND.n455 0.0151842
R4314 GND.n488 GND.n455 0.0151842
R4315 GND.n1375 GND.n1374 0.0150541
R4316 GND.n1285 GND.n1284 0.0150541
R4317 GND.n1328 GND.n1327 0.0150541
R4318 GND.n1341 GND.n1340 0.0150455
R4319 GND.n1343 GND.n1342 0.0150455
R4320 GND.n1301 GND.n1300 0.0150455
R4321 GND.n492 GND.n452 0.0149069
R4322 GND.n493 GND.n492 0.0149069
R4323 GND.n451 GND.n450 0.0146953
R4324 GND.n1281 GND.n1280 0.014225
R4325 GND.n1277 GND.n66 0.014225
R4326 GND.n1275 GND.n79 0.014225
R4327 GND.n1273 GND.n67 0.014225
R4328 GND.n1271 GND.n78 0.014225
R4329 GND.n1269 GND.n68 0.014225
R4330 GND.n1267 GND.n77 0.014225
R4331 GND.n1265 GND.n69 0.014225
R4332 GND.n1263 GND.n76 0.014225
R4333 GND.n1261 GND.n70 0.014225
R4334 GND.n1259 GND.n75 0.014225
R4335 GND.n1257 GND.n71 0.014225
R4336 GND.n1255 GND.n74 0.014225
R4337 GND.n1253 GND.n72 0.014225
R4338 GND.n1251 GND.n73 0.014225
R4339 GND.n1250 GND.n848 0.014225
R4340 GND.n1247 GND.n1246 0.014225
R4341 GND.n1243 GND.n850 0.014225
R4342 GND.n1242 GND.n852 0.014225
R4343 GND.n1239 GND.n1238 0.014225
R4344 GND.n1235 GND.n855 0.014225
R4345 GND.n1234 GND.n857 0.014225
R4346 GND.n1231 GND.n1230 0.014225
R4347 GND.n1227 GND.n860 0.014225
R4348 GND.n1226 GND.n862 0.014225
R4349 GND.n1223 GND.n1222 0.014225
R4350 GND.n1219 GND.n865 0.014225
R4351 GND.n1218 GND.n867 0.014225
R4352 GND.n1214 GND.n1213 0.014225
R4353 GND.n1210 GND.n870 0.014225
R4354 GND.n1209 GND.n872 0.014225
R4355 GND.n1205 GND.n1204 0.014225
R4356 GND.n1201 GND.n874 0.014225
R4357 GND.n1200 GND.n876 0.014225
R4358 GND.n888 GND.n887 0.014225
R4359 GND.n891 GND.n886 0.014225
R4360 GND.n892 GND.n883 0.014225
R4361 GND.n897 GND.n895 0.014225
R4362 GND.n896 GND.n880 0.014225
R4363 GND.n1195 GND.n1194 0.014225
R4364 GND.n1191 GND.n881 0.014225
R4365 GND.n1190 GND.n901 0.014225
R4366 GND.n1187 GND.n1186 0.014225
R4367 GND.n1183 GND.n904 0.014225
R4368 GND.n1182 GND.n906 0.014225
R4369 GND.n1179 GND.n1178 0.014225
R4370 GND.n1175 GND.n909 0.014225
R4371 GND.n1174 GND.n911 0.014225
R4372 GND.n1171 GND.n1170 0.014225
R4373 GND.n1167 GND.n914 0.014225
R4374 GND.n1166 GND.n916 0.014225
R4375 GND.n1069 GND.n919 0.014225
R4376 GND.n1068 GND.n921 0.014225
R4377 GND.n1065 GND.n1064 0.014225
R4378 GND.n1061 GND.n924 0.014225
R4379 GND.n1060 GND.n926 0.014225
R4380 GND.n939 GND.n938 0.014225
R4381 GND.n943 GND.n942 0.014225
R4382 GND.n946 GND.n936 0.014225
R4383 GND.n947 GND.n934 0.014225
R4384 GND.n952 GND.n950 0.014225
R4385 GND.n951 GND.n931 0.014225
R4386 GND.n1055 GND.n1054 0.014225
R4387 GND.n1051 GND.n932 0.014225
R4388 GND.n1050 GND.n956 0.014225
R4389 GND.n1047 GND.n1046 0.014225
R4390 GND.n1043 GND.n959 0.014225
R4391 GND.n1042 GND.n961 0.014225
R4392 GND.n1039 GND.n1038 0.014225
R4393 GND.n1035 GND.n964 0.014225
R4394 GND.n1034 GND.n966 0.014225
R4395 GND.n1031 GND.n1030 0.014225
R4396 GND.n1027 GND.n969 0.014225
R4397 GND.n1026 GND.n971 0.014225
R4398 GND.n1023 GND.n1022 0.014225
R4399 GND.n1019 GND.n974 0.014225
R4400 GND.n1018 GND.n976 0.014225
R4401 GND.n1014 GND.n1013 0.014225
R4402 GND.n1010 GND.n979 0.014225
R4403 GND.n1009 GND.n981 0.014225
R4404 GND.n990 GND.n989 0.014225
R4405 GND.n993 GND.n988 0.014225
R4406 GND.n994 GND.n986 0.014225
R4407 GND.n999 GND.n998 0.014225
R4408 GND.n1002 GND.n984 0.014225
R4409 GND.n1004 GND.n1003 0.014225
R4410 GND.n1380 GND.n20 0.014225
R4411 GND.n1379 GND.n18 0.014225
R4412 GND.n1407 GND.n1406 0.014225
R4413 GND.n1403 GND.n6 0.014225
R4414 GND.n1401 GND.n17 0.014225
R4415 GND.n1399 GND.n7 0.014225
R4416 GND.n1397 GND.n16 0.014225
R4417 GND.n1395 GND.n8 0.014225
R4418 GND.n1393 GND.n15 0.014225
R4419 GND.n1391 GND.n9 0.014225
R4420 GND.n1389 GND.n14 0.014225
R4421 GND.n1387 GND.n10 0.014225
R4422 GND.n1385 GND.n13 0.014225
R4423 GND.n1383 GND.n11 0.014225
R4424 GND.n12 GND.n4 0.014225
R4425 GND.n1410 GND.n1409 0.014225
R4426 GND.n1413 GND.n2 0.014225
R4427 GND.n600 GND.n143 0.013775
R4428 GND.n1312 GND.n1311 0.0137258
R4429 GND.n603 GND.n602 0.0136768
R4430 GND.n763 GND.n656 0.0136768
R4431 GND.n756 GND.n755 0.0136768
R4432 GND.n739 GND.n738 0.0136768
R4433 GND.n722 GND.n721 0.0136768
R4434 GND.n267 GND.n253 0.0136768
R4435 GND.n270 GND.n269 0.0136768
R4436 GND.n284 GND.n244 0.0136768
R4437 GND.n299 GND.n298 0.0136768
R4438 GND.n435 GND.n183 0.0136768
R4439 GND.n2768 GND.n2767 0.013625
R4440 GND.n2766 GND.n2740 0.013625
R4441 GND.n706 GND.n93 0.0131
R4442 GND.n1377 GND.n5 0.0129138
R4443 GND.n1283 GND.n65 0.0129138
R4444 GND.n1339 GND.n1338 0.0129064
R4445 GND.n1303 GND.n55 0.0129064
R4446 GND.n724 GND.n690 0.012875
R4447 GND.n746 GND.n670 0.0128066
R4448 GND.n250 GND.n247 0.0128066
R4449 GND.n660 GND.n657 0.01265
R4450 GND.n1163 GND.n1162 0.012425
R4451 GND.n3027 GND.n3026 0.012425
R4452 GND.n3026 GND.n3025 0.012425
R4453 GND.n1249 GND.n1248 0.0123657
R4454 GND.n1248 GND.n849 0.0123657
R4455 GND.n1241 GND.n1240 0.0123657
R4456 GND.n1233 GND.n858 0.0123657
R4457 GND.n1233 GND.n1232 0.0123657
R4458 GND.n1225 GND.n863 0.0123657
R4459 GND.n1225 GND.n1224 0.0123657
R4460 GND.n1217 GND.n868 0.0123657
R4461 GND.n1215 GND.n869 0.0123657
R4462 GND.n1208 GND.n869 0.0123657
R4463 GND.n1206 GND.n873 0.0123657
R4464 GND.n1199 GND.n873 0.0123657
R4465 GND.n885 GND.n877 0.0123657
R4466 GND.n894 GND.n893 0.0123657
R4467 GND.n894 GND.n878 0.0123657
R4468 GND.n1196 GND.n879 0.0123657
R4469 GND.n1189 GND.n1188 0.0123657
R4470 GND.n1188 GND.n903 0.0123657
R4471 GND.n1181 GND.n1180 0.0123657
R4472 GND.n1180 GND.n908 0.0123657
R4473 GND.n1173 GND.n1172 0.0123657
R4474 GND.n1165 GND.n917 0.0123657
R4475 GND.n1165 GND.n1164 0.0123657
R4476 GND.n1067 GND.n922 0.0123657
R4477 GND.n1067 GND.n1066 0.0123657
R4478 GND.n1059 GND.n927 0.0123657
R4479 GND.n941 GND.n928 0.0123657
R4480 GND.n941 GND.n940 0.0123657
R4481 GND.n949 GND.n948 0.0123657
R4482 GND.n949 GND.n929 0.0123657
R4483 GND.n1056 GND.n930 0.0123657
R4484 GND.n1049 GND.n1048 0.0123657
R4485 GND.n1048 GND.n958 0.0123657
R4486 GND.n1041 GND.n1040 0.0123657
R4487 GND.n1033 GND.n967 0.0123657
R4488 GND.n1033 GND.n1032 0.0123657
R4489 GND.n1025 GND.n972 0.0123657
R4490 GND.n1025 GND.n1024 0.0123657
R4491 GND.n1017 GND.n977 0.0123657
R4492 GND.n1015 GND.n978 0.0123657
R4493 GND.n1008 GND.n978 0.0123657
R4494 GND.n987 GND.n982 0.0123657
R4495 GND.n995 GND.n987 0.0123657
R4496 GND.n997 GND.n983 0.0123657
R4497 GND.n1005 GND.n21 0.0123657
R4498 GND.n1378 GND.n21 0.0123657
R4499 GND.n679 GND.n676 0.0123094
R4500 GND.n279 GND.n278 0.0123094
R4501 GND.n1198 GND.n877 0.0122537
R4502 GND.n1040 GND.n963 0.0122537
R4503 GND.n594 GND.n146 0.0118122
R4504 GND.n613 GND.n612 0.0118122
R4505 GND.n729 GND.n686 0.0118122
R4506 GND.n714 GND.n701 0.0118122
R4507 GND.n295 GND.n294 0.0118122
R4508 GND.n304 GND.n303 0.0118122
R4509 GND.n439 GND.n438 0.0118122
R4510 GND.n430 GND.n188 0.0118122
R4511 GND.n425 GND.n424 0.01175
R4512 GND.n902 GND.n879 0.0115821
R4513 GND.n1057 GND.n1056 0.0115821
R4514 GND.n674 GND.n671 0.011525
R4515 GND.n868 GND.n864 0.0113582
R4516 GND.n1017 GND.n1016 0.0113582
R4517 GND.n595 GND.n141 0.0113149
R4518 GND.n134 GND.n133 0.0113149
R4519 GND.n695 GND.n692 0.0113149
R4520 GND.n700 GND.n696 0.0113149
R4521 GND.n297 GND.n240 0.0113149
R4522 GND.n237 GND.n236 0.0113149
R4523 GND.n436 GND.n182 0.0113149
R4524 GND.n431 GND.n187 0.0113149
R4525 GND.n1360 GND.n29 0.0112292
R4526 GND.n1347 GND.n37 0.0112168
R4527 GND.n1323 GND.n1322 0.0112168
R4528 GND.n1330 GND.n1329 0.011148
R4529 GND.n1350 GND.n35 0.011063
R4530 GND.n1351 GND.n35 0.011063
R4531 GND.n1352 GND.n34 0.011063
R4532 GND.n1353 GND.n34 0.011063
R4533 GND.n1355 GND.n30 0.011063
R4534 GND.n1356 GND.n30 0.011063
R4535 GND.n1312 GND.n50 0.0110528
R4536 GND.n1313 GND.n50 0.0110528
R4537 GND.n1318 GND.n1314 0.0110528
R4538 GND.n1317 GND.n1314 0.0110528
R4539 GND.n1317 GND.n1316 0.0110528
R4540 GND.n1316 GND.n1315 0.0110528
R4541 GND.n1315 GND.n32 0.0110528
R4542 GND.n591 GND.n590 0.0108177
R4543 GND.n137 GND.n132 0.0108177
R4544 GND.n731 GND.n685 0.0108177
R4545 GND.n712 GND.n704 0.0108177
R4546 GND.n288 GND.n287 0.0108177
R4547 GND.n307 GND.n235 0.0108177
R4548 GND.n443 GND.n442 0.0108177
R4549 GND.n427 GND.n191 0.0108177
R4550 GND.n1172 GND.n913 0.0106866
R4551 GND.n927 GND.n923 0.0106866
R4552 GND.n1281 GND.n80 0.010625
R4553 GND.n1280 GND.n66 0.010625
R4554 GND.n1277 GND.n79 0.010625
R4555 GND.n1275 GND.n67 0.010625
R4556 GND.n1273 GND.n78 0.010625
R4557 GND.n1271 GND.n68 0.010625
R4558 GND.n1269 GND.n77 0.010625
R4559 GND.n1267 GND.n69 0.010625
R4560 GND.n1265 GND.n76 0.010625
R4561 GND.n1263 GND.n70 0.010625
R4562 GND.n1261 GND.n75 0.010625
R4563 GND.n1259 GND.n71 0.010625
R4564 GND.n1257 GND.n74 0.010625
R4565 GND.n1255 GND.n72 0.010625
R4566 GND.n1253 GND.n73 0.010625
R4567 GND.n1251 GND.n1250 0.010625
R4568 GND.n1247 GND.n848 0.010625
R4569 GND.n1246 GND.n850 0.010625
R4570 GND.n1243 GND.n1242 0.010625
R4571 GND.n1239 GND.n852 0.010625
R4572 GND.n1238 GND.n855 0.010625
R4573 GND.n1235 GND.n1234 0.010625
R4574 GND.n1231 GND.n857 0.010625
R4575 GND.n1230 GND.n860 0.010625
R4576 GND.n1227 GND.n1226 0.010625
R4577 GND.n1223 GND.n862 0.010625
R4578 GND.n1222 GND.n865 0.010625
R4579 GND.n1219 GND.n1218 0.010625
R4580 GND.n1214 GND.n867 0.010625
R4581 GND.n1213 GND.n870 0.010625
R4582 GND.n1210 GND.n1209 0.010625
R4583 GND.n1205 GND.n872 0.010625
R4584 GND.n1204 GND.n874 0.010625
R4585 GND.n1201 GND.n1200 0.010625
R4586 GND.n887 GND.n876 0.010625
R4587 GND.n888 GND.n886 0.010625
R4588 GND.n892 GND.n891 0.010625
R4589 GND.n895 GND.n883 0.010625
R4590 GND.n897 GND.n896 0.010625
R4591 GND.n1195 GND.n880 0.010625
R4592 GND.n1194 GND.n881 0.010625
R4593 GND.n1191 GND.n1190 0.010625
R4594 GND.n1187 GND.n901 0.010625
R4595 GND.n1186 GND.n904 0.010625
R4596 GND.n1183 GND.n1182 0.010625
R4597 GND.n1179 GND.n906 0.010625
R4598 GND.n1178 GND.n909 0.010625
R4599 GND.n1175 GND.n1174 0.010625
R4600 GND.n1171 GND.n911 0.010625
R4601 GND.n1170 GND.n914 0.010625
R4602 GND.n1167 GND.n1166 0.010625
R4603 GND.n1163 GND.n916 0.010625
R4604 GND.n1072 GND.n919 0.010625
R4605 GND.n1069 GND.n1068 0.010625
R4606 GND.n1065 GND.n921 0.010625
R4607 GND.n1064 GND.n924 0.010625
R4608 GND.n1061 GND.n1060 0.010625
R4609 GND.n938 GND.n926 0.010625
R4610 GND.n942 GND.n939 0.010625
R4611 GND.n943 GND.n936 0.010625
R4612 GND.n947 GND.n946 0.010625
R4613 GND.n950 GND.n934 0.010625
R4614 GND.n952 GND.n951 0.010625
R4615 GND.n1055 GND.n931 0.010625
R4616 GND.n1054 GND.n932 0.010625
R4617 GND.n1051 GND.n1050 0.010625
R4618 GND.n1047 GND.n956 0.010625
R4619 GND.n1046 GND.n959 0.010625
R4620 GND.n1043 GND.n1042 0.010625
R4621 GND.n1039 GND.n961 0.010625
R4622 GND.n1038 GND.n964 0.010625
R4623 GND.n1035 GND.n1034 0.010625
R4624 GND.n1031 GND.n966 0.010625
R4625 GND.n1030 GND.n969 0.010625
R4626 GND.n1027 GND.n1026 0.010625
R4627 GND.n1023 GND.n971 0.010625
R4628 GND.n1022 GND.n974 0.010625
R4629 GND.n1019 GND.n1018 0.010625
R4630 GND.n1014 GND.n976 0.010625
R4631 GND.n1013 GND.n979 0.010625
R4632 GND.n1010 GND.n1009 0.010625
R4633 GND.n989 GND.n981 0.010625
R4634 GND.n990 GND.n988 0.010625
R4635 GND.n994 GND.n993 0.010625
R4636 GND.n998 GND.n986 0.010625
R4637 GND.n999 GND.n984 0.010625
R4638 GND.n1004 GND.n1002 0.010625
R4639 GND.n1003 GND.n20 0.010625
R4640 GND.n1380 GND.n1379 0.010625
R4641 GND.n1407 GND.n18 0.010625
R4642 GND.n1406 GND.n6 0.010625
R4643 GND.n1403 GND.n17 0.010625
R4644 GND.n1401 GND.n7 0.010625
R4645 GND.n1399 GND.n16 0.010625
R4646 GND.n1397 GND.n8 0.010625
R4647 GND.n1395 GND.n15 0.010625
R4648 GND.n1393 GND.n9 0.010625
R4649 GND.n1391 GND.n14 0.010625
R4650 GND.n1389 GND.n10 0.010625
R4651 GND.n1387 GND.n13 0.010625
R4652 GND.n1385 GND.n11 0.010625
R4653 GND.n1383 GND.n12 0.010625
R4654 GND.n1409 GND.n4 0.010625
R4655 GND.n1410 GND.n2 0.010625
R4656 GND.n1241 GND.n853 0.0104627
R4657 GND.n1006 GND.n983 0.0104627
R4658 GND.n1684 GND.n1445 0.0103253
R4659 GND.n1685 GND.n1684 0.0103253
R4660 GND.n2329 GND.n1445 0.0103253
R4661 GND.n582 GND.n581 0.0103204
R4662 GND.n148 GND.n147 0.0103204
R4663 GND.n617 GND.n616 0.0103204
R4664 GND.n773 GND.n106 0.0103204
R4665 GND.n684 GND.n680 0.0103204
R4666 GND.n707 GND.n94 0.0103204
R4667 GND.n818 GND.n817 0.0103204
R4668 GND.n285 GND.n243 0.0103204
R4669 GND.n308 GND.n232 0.0103204
R4670 GND.n381 GND.n380 0.0103204
R4671 GND.n447 GND.n446 0.0103204
R4672 GND.n445 GND.n178 0.0103204
R4673 GND.n426 GND.n189 0.0103204
R4674 GND.n422 GND.n421 0.0103204
R4675 GND.n495 GND.n494 0.0102808
R4676 GND.n491 GND.n453 0.0102808
R4677 GND.n494 GND.n491 0.0102808
R4678 GND.n495 GND.n490 0.0102808
R4679 GND.n1352 GND.n1351 0.0102066
R4680 GND.n795 GND.n794 0.0101961
R4681 GND.n789 GND.n788 0.0101961
R4682 GND.n788 GND.n787 0.0101961
R4683 GND.n782 GND.n781 0.0101961
R4684 GND.n781 GND.n780 0.0101961
R4685 GND.n775 GND.n774 0.0101961
R4686 GND.n420 GND.n419 0.0101961
R4687 GND.n414 GND.n413 0.0101961
R4688 GND.n413 GND.n412 0.0101961
R4689 GND.n407 GND.n406 0.0101961
R4690 GND.n406 GND.n405 0.0101961
R4691 GND.n400 GND.n399 0.0101961
R4692 GND.n1240 GND.n854 0.0100149
R4693 GND.n997 GND.n996 0.0100149
R4694 GND.n748 GND.n669 0.0098232
R4695 GND.n275 GND.n274 0.0098232
R4696 GND.n1173 GND.n912 0.00979105
R4697 GND.n1059 GND.n1058 0.00979105
R4698 GND.n1320 GND.n1318 0.00965829
R4699 GND.n1978 GND.n1683 0.00964634
R4700 GND.n2953 GND.n1446 0.00964634
R4701 GND.n2953 GND.n2952 0.00964634
R4702 GND.n1979 GND.n1978 0.00964634
R4703 GND.n756 GND.n663 0.00959771
R4704 GND.n269 GND.n268 0.00959771
R4705 GND.n765 GND.n764 0.00957459
R4706 GND.n261 GND.n260 0.00957459
R4707 GND.n668 GND.n664 0.00932597
R4708 GND.n249 GND.n248 0.00932597
R4709 GND.n1217 GND.n1216 0.0091194
R4710 GND.n977 GND.n973 0.0091194
R4711 GND.n1197 GND.n1196 0.00889552
R4712 GND.n957 GND.n930 0.00889552
R4713 GND.n765 GND.n655 0.00882873
R4714 GND.n261 GND.n259 0.00882873
R4715 GND.n741 GND.n674 0.008825
R4716 GND.n792 GND.n791 0.00870442
R4717 GND.n785 GND.n784 0.00870442
R4718 GND.n778 GND.n777 0.00870442
R4719 GND.n417 GND.n416 0.00870442
R4720 GND.n410 GND.n409 0.00870442
R4721 GND.n403 GND.n402 0.00870442
R4722 GND.n748 GND.n747 0.00858011
R4723 GND.n274 GND.n251 0.00858011
R4724 GND.n647 GND.n115 0.0084558
R4725 GND.n773 GND.n772 0.00833149
R4726 GND.n654 GND.n108 0.00833149
R4727 GND.n421 GND.n195 0.00833149
R4728 GND.n257 GND.n256 0.00833149
R4729 GND.n1331 GND.n1330 0.00832143
R4730 GND.n573 GND.n567 0.00825457
R4731 GND.n581 GND.n153 0.00825457
R4732 GND.n809 GND.n97 0.00825457
R4733 GND.n817 GND.n816 0.00825457
R4734 GND.n447 GND.n177 0.00825457
R4735 GND.n215 GND.n206 0.00825457
R4736 GND.n381 GND.n230 0.00825457
R4737 GND.n389 GND.n227 0.00825457
R4738 GND.n885 GND.n884 0.00822388
R4739 GND.n1041 GND.n962 0.00822388
R4740 GND.n1207 GND.n1206 0.008
R4741 GND.n1032 GND.n968 0.008
R4742 GND.t28 GND.n457 0.00784211
R4743 GND.t28 GND.n456 0.00784211
R4744 GND.n758 GND.n660 0.0077
R4745 GND.n796 GND.n99 0.00759641
R4746 GND.n398 GND.n222 0.00759641
R4747 GND.n590 GND.n149 0.00758564
R4748 GND.n137 GND.n135 0.00758564
R4749 GND.n731 GND.n730 0.00758564
R4750 GND.n713 GND.n712 0.00758564
R4751 GND.n288 GND.n241 0.00758564
R4752 GND.n238 GND.n235 0.00758564
R4753 GND.n442 GND.n179 0.00758564
R4754 GND.n191 GND.n190 0.00758564
R4755 GND.n690 GND.n687 0.007475
R4756 GND.n1333 GND.n1332 0.00735714
R4757 GND.n1408 GND.n5 0.00734899
R4758 GND.n1283 GND.n1282 0.00734899
R4759 GND.n907 GND.n903 0.00732836
R4760 GND.n948 GND.n935 0.00732836
R4761 GND.n708 GND.n706 0.00725
R4762 GND.n863 GND.n859 0.00710448
R4763 GND.n1008 GND.n1007 0.00710448
R4764 GND.n149 GND.n146 0.00659116
R4765 GND.n612 GND.n135 0.00659116
R4766 GND.n730 GND.n729 0.00659116
R4767 GND.n714 GND.n713 0.00659116
R4768 GND.n294 GND.n241 0.00659116
R4769 GND.n303 GND.n238 0.00659116
R4770 GND.n439 GND.n179 0.00659116
R4771 GND.n190 GND.n188 0.00659116
R4772 GND.n596 GND.n143 0.006575
R4773 GND.n1446 GND.n1444 0.00647611
R4774 GND.n1686 GND.n1683 0.00646981
R4775 GND.n1164 GND.n918 0.00643284
R4776 GND.n922 GND.n918 0.00643284
R4777 GND.n773 GND.n107 0.00609392
R4778 GND.n421 GND.n196 0.00609392
R4779 GND.n772 GND.n108 0.0058453
R4780 GND.n257 GND.n195 0.0058453
R4781 GND.n1232 GND.n859 0.00576119
R4782 GND.n1007 GND.n982 0.00576119
R4783 GND.n747 GND.n746 0.00559669
R4784 GND.n251 GND.n250 0.00559669
R4785 GND.n663 GND.n656 0.00557014
R4786 GND.n268 GND.n267 0.00557014
R4787 GND.n1181 GND.n907 0.00553731
R4788 GND.n940 GND.n935 0.00553731
R4789 GND.n320 GND.n231 0.00543473
R4790 GND.n655 GND.n654 0.00534807
R4791 GND.n259 GND.n256 0.00534807
R4792 GND.n1354 GND.n1353 0.0050678
R4793 GND.n1355 GND.n1354 0.0050678
R4794 GND.n792 GND.n100 0.00505453
R4795 GND.n791 GND.n101 0.00505453
R4796 GND.n785 GND.n102 0.00505453
R4797 GND.n784 GND.n103 0.00505453
R4798 GND.n778 GND.n104 0.00505453
R4799 GND.n777 GND.n105 0.00505453
R4800 GND.n115 GND.n113 0.00505453
R4801 GND.n199 GND.n198 0.00505453
R4802 GND.n417 GND.n197 0.00505453
R4803 GND.n416 GND.n201 0.00505453
R4804 GND.n410 GND.n202 0.00505453
R4805 GND.n409 GND.n203 0.00505453
R4806 GND.n403 GND.n204 0.00505453
R4807 GND.n402 GND.n205 0.00505453
R4808 GND.n563 GND.n160 0.005
R4809 GND.n562 GND.n154 0.005
R4810 GND.n559 GND.n159 0.005
R4811 GND.n557 GND.n155 0.005
R4812 GND.n555 GND.n158 0.005
R4813 GND.n553 GND.n156 0.005
R4814 GND.n551 GND.n157 0.005
R4815 GND.n583 GND.n152 0.005
R4816 GND.n584 GND.n150 0.005
R4817 GND.n589 GND.n587 0.005
R4818 GND.n588 GND.n145 0.005
R4819 GND.n597 GND.n596 0.005
R4820 GND.n601 GND.n600 0.005
R4821 GND.n604 GND.n140 0.005
R4822 GND.n606 GND.n605 0.005
R4823 GND.n611 GND.n136 0.005
R4824 GND.n610 GND.n138 0.005
R4825 GND.n618 GND.n131 0.005
R4826 GND.n621 GND.n620 0.005
R4827 GND.n646 GND.n128 0.005
R4828 GND.n645 GND.n116 0.005
R4829 GND.n642 GND.n127 0.005
R4830 GND.n640 GND.n117 0.005
R4831 GND.n638 GND.n126 0.005
R4832 GND.n636 GND.n118 0.005
R4833 GND.n634 GND.n125 0.005
R4834 GND.n632 GND.n119 0.005
R4835 GND.n630 GND.n124 0.005
R4836 GND.n628 GND.n120 0.005
R4837 GND.n626 GND.n123 0.005
R4838 GND.n624 GND.n122 0.005
R4839 GND.n121 GND.n112 0.005
R4840 GND.n649 GND.n648 0.005
R4841 GND.n771 GND.n109 0.005
R4842 GND.n770 GND.n110 0.005
R4843 GND.n767 GND.n766 0.005
R4844 GND.n762 GND.n653 0.005
R4845 GND.n761 GND.n657 0.005
R4846 GND.n758 GND.n757 0.005
R4847 GND.n754 GND.n661 0.005
R4848 GND.n753 GND.n665 0.005
R4849 GND.n750 GND.n749 0.005
R4850 GND.n745 GND.n667 0.005
R4851 GND.n744 GND.n671 0.005
R4852 GND.n741 GND.n740 0.005
R4853 GND.n737 GND.n675 0.005
R4854 GND.n736 GND.n681 0.005
R4855 GND.n733 GND.n732 0.005
R4856 GND.n728 GND.n683 0.005
R4857 GND.n727 GND.n687 0.005
R4858 GND.n724 GND.n723 0.005
R4859 GND.n720 GND.n691 0.005
R4860 GND.n719 GND.n697 0.005
R4861 GND.n716 GND.n715 0.005
R4862 GND.n711 GND.n699 0.005
R4863 GND.n710 GND.n708 0.005
R4864 GND.n819 GND.n93 0.005
R4865 GND.n820 GND.n88 0.005
R4866 GND.n822 GND.n89 0.005
R4867 GND.n824 GND.n90 0.005
R4868 GND.n826 GND.n91 0.005
R4869 GND.n830 GND.n829 0.005
R4870 GND.n832 GND.n86 0.005
R4871 GND.n833 GND.n84 0.005
R4872 GND.n1208 GND.n1207 0.00486567
R4873 GND.n972 GND.n968 0.00486567
R4874 GND.n755 GND.n664 0.00485083
R4875 GND.n270 GND.n248 0.00485083
R4876 GND.n619 GND.n618 0.004775
R4877 GND.n893 GND.n884 0.00464179
R4878 GND.n962 GND.n958 0.00464179
R4879 GND.n796 GND.n795 0.00460221
R4880 GND.n774 GND.n773 0.00460221
R4881 GND.n764 GND.n763 0.00460221
R4882 GND.n260 GND.n253 0.00460221
R4883 GND.n421 GND.n420 0.00460221
R4884 GND.n399 GND.n398 0.00460221
R4885 GND.n500 GND.n499 0.00455
R4886 GND.n1330 GND.n46 0.00440606
R4887 GND.n1359 GND.n1358 0.00435417
R4888 GND.n669 GND.n668 0.00435359
R4889 GND.n275 GND.n249 0.00435359
R4890 GND.n1349 GND.n1348 0.00434971
R4891 GND.n1321 GND.n1320 0.00434971
R4892 GND.n1197 GND.n878 0.00397015
R4893 GND.n1049 GND.n957 0.00397015
R4894 GND.n1377 GND.n1376 0.00392449
R4895 GND.n65 GND.n64 0.00392449
R4896 GND.n1338 GND.n41 0.00392246
R4897 GND.n1303 GND.n1302 0.00392246
R4898 GND.n582 GND.n147 0.00385635
R4899 GND.n616 GND.n106 0.00385635
R4900 GND.n738 GND.n680 0.00385635
R4901 GND.n818 GND.n94 0.00385635
R4902 GND.n285 GND.n284 0.00385635
R4903 GND.n380 GND.n232 0.00385635
R4904 GND.n446 GND.n445 0.00385635
R4905 GND.n422 GND.n189 0.00385635
R4906 GND.n1216 GND.n1215 0.00374627
R4907 GND.n1024 GND.n973 0.00374627
R4908 GND.n591 GND.n148 0.00335912
R4909 GND.n617 GND.n132 0.00335912
R4910 GND.n685 GND.n684 0.00335912
R4911 GND.n707 GND.n704 0.00335912
R4912 GND.n287 GND.n243 0.00335912
R4913 GND.n308 GND.n307 0.00335912
R4914 GND.n443 GND.n178 0.00335912
R4915 GND.n427 GND.n426 0.00335912
R4916 GND.n775 GND.n105 0.00328344
R4917 GND.n113 GND.n107 0.00328344
R4918 GND.n782 GND.n103 0.00328344
R4919 GND.n780 GND.n104 0.00328344
R4920 GND.n789 GND.n101 0.00328344
R4921 GND.n787 GND.n102 0.00328344
R4922 GND.n794 GND.n100 0.00328344
R4923 GND.n400 GND.n205 0.00328344
R4924 GND.n407 GND.n203 0.00328344
R4925 GND.n405 GND.n204 0.00328344
R4926 GND.n414 GND.n201 0.00328344
R4927 GND.n412 GND.n202 0.00328344
R4928 GND.n198 GND.n196 0.00328344
R4929 GND.n419 GND.n197 0.00328344
R4930 GND.n912 GND.n908 0.00307463
R4931 GND.n1058 GND.n928 0.00307463
R4932 GND.n602 GND.n141 0.00286188
R4933 GND.n603 GND.n133 0.00286188
R4934 GND.n722 GND.n695 0.00286188
R4935 GND.n721 GND.n696 0.00286188
R4936 GND.n298 GND.n297 0.00286188
R4937 GND.n299 GND.n236 0.00286188
R4938 GND.n436 GND.n435 0.00286188
R4939 GND.n187 GND.n183 0.00286188
R4940 GND.n858 GND.n854 0.00285075
R4941 GND.n996 GND.n995 0.00285075
R4942 GND.n853 GND.n849 0.00240299
R4943 GND.n1006 GND.n1005 0.00240299
R4944 GND.n595 GND.n594 0.00236464
R4945 GND.n613 GND.n134 0.00236464
R4946 GND.n692 GND.n686 0.00236464
R4947 GND.n701 GND.n700 0.00236464
R4948 GND.n295 GND.n240 0.00236464
R4949 GND.n304 GND.n237 0.00236464
R4950 GND.n438 GND.n182 0.00236464
R4951 GND.n431 GND.n430 0.00236464
R4952 GND.n1162 GND.n1072 0.0023
R4953 GND.n917 GND.n913 0.0021791
R4954 GND.n1066 GND.n923 0.0021791
R4955 GND.n1350 GND.n1349 0.00199881
R4956 GND.n1358 GND.n1356 0.00199881
R4957 GND.n1249 GND.n65 0.00195522
R4958 GND.n1378 GND.n1377 0.00195522
R4959 GND.n1354 GND.n32 0.00193216
R4960 GND.n1320 GND.n1313 0.00189447
R4961 GND.n739 GND.n679 0.0018674
R4962 GND.n278 GND.n244 0.0018674
R4963 GND.n1224 GND.n864 0.00150746
R4964 GND.n1016 GND.n1015 0.00150746
R4965 GND.n676 GND.n670 0.00137017
R4966 GND.n279 GND.n247 0.00137017
R4967 GND.n1189 GND.n902 0.00128358
R4968 GND.n1057 GND.n929 0.00128358
R4969 GND.n1199 GND.n1198 0.00061194
R4970 GND.n967 GND.n963 0.00061194
R4971 a_21743_6748.n1 a_21743_6748.n0 16.2768
R4972 a_21743_6748.t10 a_21743_6748.n2 8.42794
R4973 a_21743_6748.n1 a_21743_6748.t12 8.44632
R4974 a_21743_6748.n0 a_21743_6748.t6 14.0566
R4975 a_21743_6748.n1 a_21743_6748.t5 13.9025
R4976 a_21743_6748.n2 a_21743_6748.t4 13.5018
R4977 a_21743_6748.n0 a_21743_6748.t1 13.3613
R4978 a_21743_6748.n0 a_21743_6748.t3 13.3613
R4979 a_21743_6748.n0 a_21743_6748.t0 13.3606
R4980 a_21743_6748.n0 a_21743_6748.t7 13.3305
R4981 a_21743_6748.n0 a_21743_6748.t2 13.3292
R4982 a_21743_6748.n0 a_21743_6748.t9 13.3288
R4983 a_21743_6748.n0 a_21743_6748.t8 13.3182
R4984 a_21743_6748.n1 a_21743_6748.t15 10.7255
R4985 a_21743_6748.t13 a_21743_6748.n1 10.5667
R4986 a_21743_6748.n2 a_21743_6748.t11 10.5446
R4987 a_21743_6748.n1 a_21743_6748.t17 9.65646
R4988 a_21743_6748.n1 a_21743_6748.t16 8.61301
R4989 a_21743_6748.n1 a_21743_6748.t14 8.57431
R4990 a_21743_6748.n1 a_21743_6748.n2 7.8313
R4991 a_21743_6100.t10 a_21743_6100.n1 8.45596
R4992 a_21743_6100.n2 a_21743_6100.t4 15.2205
R4993 a_21743_6100.n1 a_21743_6100.t13 13.8811
R4994 a_21743_6100.n1 a_21743_6100.t12 13.5061
R4995 a_21743_6100.n2 a_21743_6100.t2 13.1505
R4996 a_21743_6100.n2 a_21743_6100.t0 13.1484
R4997 a_21743_6100.n2 a_21743_6100.t7 13.1469
R4998 a_21743_6100.n2 a_21743_6100.t1 13.1463
R4999 a_21743_6100.n2 a_21743_6100.t6 13.1463
R5000 a_21743_6100.n2 a_21743_6100.t3 13.1436
R5001 a_21743_6100.n0 a_21743_6100.n2 10.8237
R5002 a_21743_6100.n0 a_21743_6100.t5 10.7513
R5003 a_21743_6100.t11 a_21743_6100.n1 10.5704
R5004 a_21743_6100.n1 a_21743_6100.t9 10.5629
R5005 a_21743_6100.n1 a_21743_6100.t16 10.3448
R5006 a_21743_6100.n1 a_21743_6100.n0 9.61388
R5007 a_21743_6100.n1 a_21743_6100.t14 8.61428
R5008 a_21743_6100.n1 a_21743_6100.t15 8.57979
R5009 a_21743_6100.n1 a_21743_6100.t8 8.53382
R5010 a_21743_6100.n1 a_21743_6100.t17 8.51529
R5011 a_21659_3242.n0 a_21659_3242.t1 13.6222
R5012 a_21659_3242.n0 a_21659_3242.t10 13.5669
R5013 a_21659_3242.n3 a_21659_3242.t25 13.5669
R5014 a_21659_3242.n0 a_21659_3242.t4 13.5665
R5015 a_21659_3242.n4 a_21659_3242.t27 13.5665
R5016 a_21659_3242.n4 a_21659_3242.t3 13.5665
R5017 a_21659_3242.n3 a_21659_3242.t2 13.5665
R5018 a_21659_3242.n1 a_21659_3242.t9 13.5654
R5019 a_21659_3242.n2 a_21659_3242.t5 13.5643
R5020 a_21659_3242.n1 a_21659_3242.t24 13.5643
R5021 a_21659_3242.t7 a_21659_3242.n5 13.5643
R5022 a_21659_3242.n2 a_21659_3242.t11 13.5639
R5023 a_21659_3242.n1 a_21659_3242.t0 13.5635
R5024 a_21659_3242.n5 a_21659_3242.t8 13.5596
R5025 a_21659_3242.n15 a_21659_3242.t26 11.4211
R5026 a_21659_3242.n17 a_21659_3242.t6 11.2961
R5027 a_21659_3242.n6 a_21659_3242.n12 4.62286
R5028 a_21659_3242.n7 a_21659_3242.n9 4.62286
R5029 a_21659_3242.n5 a_21659_3242.n3 4.33657
R5030 a_21659_3242.n6 a_21659_3242.n14 3.98468
R5031 a_21659_3242.n6 a_21659_3242.n13 3.98468
R5032 a_21659_3242.n8 a_21659_3242.n11 3.98468
R5033 a_21659_3242.n7 a_21659_3242.n10 3.98468
R5034 a_21659_3242.n17 a_21659_3242.n16 2.97211
R5035 a_21659_3242.n1 a_21659_3242.n17 2.93779
R5036 a_21659_3242.n15 a_21659_3242.n0 2.92
R5037 a_21659_3242.n0 a_21659_3242.n4 2.75836
R5038 a_21659_3242.n8 a_21659_3242.n6 2.15026
R5039 a_21659_3242.n5 a_21659_3242.n2 2.0705
R5040 a_21659_3242.n2 a_21659_3242.n1 2.06773
R5041 a_21659_3242.n16 a_21659_3242.n8 1.57764
R5042 a_21659_3242.n4 a_21659_3242.n3 1.37836
R5043 a_21659_3242.n8 a_21659_3242.n7 1.07026
R5044 a_21659_3242.n16 a_21659_3242.n15 0.927751
R5045 a_21659_3242.n14 a_21659_3242.t17 0.9105
R5046 a_21659_3242.n14 a_21659_3242.t19 0.9105
R5047 a_21659_3242.n13 a_21659_3242.t15 0.9105
R5048 a_21659_3242.n13 a_21659_3242.t23 0.9105
R5049 a_21659_3242.n12 a_21659_3242.t21 0.9105
R5050 a_21659_3242.n12 a_21659_3242.t18 0.9105
R5051 a_21659_3242.n11 a_21659_3242.t14 0.9105
R5052 a_21659_3242.n11 a_21659_3242.t22 0.9105
R5053 a_21659_3242.n10 a_21659_3242.t12 0.9105
R5054 a_21659_3242.n10 a_21659_3242.t13 0.9105
R5055 a_21659_3242.n9 a_21659_3242.t16 0.9105
R5056 a_21659_3242.n9 a_21659_3242.t20 0.9105
R5057 a_11345_12294.t0 a_11345_12294.t3 23.7444
R5058 a_11345_12294.t1 a_11345_12294.t0 14.5807
R5059 a_11345_12294.t3 a_11345_12294.t4 7.58125
R5060 a_11345_12294.t5 a_11345_12294.t3 7.34053
R5061 a_11345_12294.t3 a_11345_12294.t2 7.26371
R5062 VDD.t3 VDD.t271 1513.51
R5063 VDD.t271 VDD.t263 1193.15
R5064 VDD.t265 VDD.t3 1193.15
R5065 VDD.t263 VDD.n1 749.592
R5066 VDD.n2 VDD.t265 749.423
R5067 VDD.t19 VDD.t16 204.879
R5068 VDD.t26 VDD.t23 204.879
R5069 VDD.t6 VDD.t4 204.879
R5070 VDD.t10 VDD.t8 204.879
R5071 VDD.n493 VDD.n39 195.466
R5072 VDD.n495 VDD.n39 195.466
R5073 VDD.n548 VDD.n8 195.466
R5074 VDD.n550 VDD.n8 195.466
R5075 VDD.t16 VDD.n493 188.95
R5076 VDD.n495 VDD.t26 188.95
R5077 VDD.t4 VDD.n548 188.95
R5078 VDD.n550 VDD.t10 188.95
R5079 VDD.n493 VDD.n40 183.53
R5080 VDD.n495 VDD.n40 183.53
R5081 VDD.n548 VDD.n7 183.53
R5082 VDD.n550 VDD.n7 183.53
R5083 VDD.n891 VDD.n568 112.903
R5084 VDD.n889 VDD.n888 112.903
R5085 VDD.n494 VDD.t19 102.439
R5086 VDD.t23 VDD.n494 102.439
R5087 VDD.n549 VDD.t6 102.439
R5088 VDD.t8 VDD.n549 102.439
R5089 VDD.n888 VDD.n887 87.2367
R5090 VDD.n891 VDD.n890 87.2367
R5091 VDD.n919 VDD.n562 71.4558
R5092 VDD.n917 VDD.n916 71.4558
R5093 VDD.n916 VDD.n915 60.8228
R5094 VDD.n919 VDD.n918 60.8228
R5095 VDD.n582 VDD.n575 17.0302
R5096 VDD.n169 VDD.t165 14.743
R5097 VDD.n147 VDD.t247 14.743
R5098 VDD.n140 VDD.t139 14.743
R5099 VDD.n260 VDD.t241 14.742
R5100 VDD.t253 VDD.n241 14.742
R5101 VDD.n234 VDD.t195 14.742
R5102 VDD.n165 VDD.t73 14.7277
R5103 VDD.t73 VDD.n164 14.7277
R5104 VDD.n167 VDD.t55 14.7277
R5105 VDD.t55 VDD.n166 14.7277
R5106 VDD.t165 VDD.n168 14.7277
R5107 VDD.n211 VDD.t119 14.7277
R5108 VDD.n213 VDD.t119 14.7277
R5109 VDD.n208 VDD.t117 14.7277
R5110 VDD.n210 VDD.t117 14.7277
R5111 VDD.n153 VDD.t125 14.7277
R5112 VDD.n155 VDD.t125 14.7277
R5113 VDD.n150 VDD.t179 14.7277
R5114 VDD.n152 VDD.t179 14.7277
R5115 VDD.n149 VDD.t247 14.7277
R5116 VDD.n136 VDD.t237 14.7277
R5117 VDD.t237 VDD.n125 14.7277
R5118 VDD.n138 VDD.t57 14.7277
R5119 VDD.t57 VDD.n137 14.7277
R5120 VDD.t139 VDD.n139 14.7277
R5121 VDD.n258 VDD.t241 14.7277
R5122 VDD.n255 VDD.t225 14.7277
R5123 VDD.n257 VDD.t225 14.7277
R5124 VDD.n252 VDD.t107 14.7277
R5125 VDD.n254 VDD.t107 14.7277
R5126 VDD.n300 VDD.t259 14.7277
R5127 VDD.t259 VDD.n299 14.7277
R5128 VDD.n302 VDD.t149 14.7277
R5129 VDD.t149 VDD.n301 14.7277
R5130 VDD.n242 VDD.t253 14.7277
R5131 VDD.n244 VDD.t203 14.7277
R5132 VDD.t203 VDD.n243 14.7277
R5133 VDD.n246 VDD.t143 14.7277
R5134 VDD.t143 VDD.n245 14.7277
R5135 VDD.n232 VDD.t195 14.7277
R5136 VDD.n229 VDD.t145 14.7277
R5137 VDD.n231 VDD.t145 14.7277
R5138 VDD.t63 VDD.n216 14.7277
R5139 VDD.n228 VDD.t63 14.7277
R5140 VDD.n1 VDD.t264 14.6005
R5141 VDD.n0 VDD.t266 14.6005
R5142 VDD.n1014 VDD.t270 12.6668
R5143 VDD.n441 VDD.n440 11.1505
R5144 VDD.n431 VDD.n430 11.1505
R5145 VDD.n423 VDD.n56 11.1505
R5146 VDD.n422 VDD.n60 11.1505
R5147 VDD.n413 VDD.n412 11.1505
R5148 VDD.n403 VDD.n402 11.1505
R5149 VDD.n396 VDD.n71 11.1505
R5150 VDD.n395 VDD.n75 11.1505
R5151 VDD.n385 VDD.n384 11.1505
R5152 VDD.n376 VDD.n375 11.1505
R5153 VDD.n369 VDD.n368 11.1505
R5154 VDD.n367 VDD.n90 11.1505
R5155 VDD.n359 VDD.n358 11.1505
R5156 VDD.n350 VDD.n349 11.1505
R5157 VDD.n343 VDD.n342 11.1505
R5158 VDD.n341 VDD.n106 11.1505
R5159 VDD.n333 VDD.n332 11.1505
R5160 VDD.n323 VDD.n322 11.1505
R5161 VDD.n315 VDD.n118 11.1505
R5162 VDD.n314 VDD.n122 11.1505
R5163 VDD.n441 VDD.n51 11.1505
R5164 VDD.n430 VDD.n55 11.1505
R5165 VDD.n59 VDD.n56 11.1505
R5166 VDD.n62 VDD.n60 11.1505
R5167 VDD.n413 VDD.n66 11.1505
R5168 VDD.n402 VDD.n70 11.1505
R5169 VDD.n74 VDD.n71 11.1505
R5170 VDD.n77 VDD.n75 11.1505
R5171 VDD.n385 VDD.n81 11.1505
R5172 VDD.n375 VDD.n85 11.1505
R5173 VDD.n369 VDD.n89 11.1505
R5174 VDD.n92 VDD.n90 11.1505
R5175 VDD.n359 VDD.n97 11.1505
R5176 VDD.n349 VDD.n101 11.1505
R5177 VDD.n343 VDD.n105 11.1505
R5178 VDD.n108 VDD.n106 11.1505
R5179 VDD.n333 VDD.n113 11.1505
R5180 VDD.n322 VDD.n117 11.1505
R5181 VDD.n121 VDD.n118 11.1505
R5182 VDD.n124 VDD.n122 11.1505
R5183 VDD.n182 VDD.n181 11.1505
R5184 VDD.n188 VDD.n187 11.1505
R5185 VDD.n190 VDD.n189 11.1505
R5186 VDD.n195 VDD.n194 11.1505
R5187 VDD.n197 VDD.n196 11.1505
R5188 VDD.n202 VDD.n201 11.1505
R5189 VDD.n204 VDD.n203 11.1505
R5190 VDD.n273 VDD.n272 11.1505
R5191 VDD.n279 VDD.n278 11.1505
R5192 VDD.n281 VDD.n280 11.1505
R5193 VDD.n286 VDD.n285 11.1505
R5194 VDD.n288 VDD.n287 11.1505
R5195 VDD.n293 VDD.n292 11.1505
R5196 VDD.n295 VDD.n294 11.1505
R5197 VDD.n304 VDD.t38 11.0944
R5198 VDD.n305 VDD.t267 11.0944
R5199 VDD.n304 VDD.t0 10.8102
R5200 VDD.n305 VDD.t268 10.8102
R5201 VDD.t66 VDD.n126 8.44802
R5202 VDD.t42 VDD.n217 8.44802
R5203 VDD.t208 VDD.n126 8.44712
R5204 VDD.t228 VDD.n217 8.44712
R5205 VDD.n156 VDD.t148 8.44573
R5206 VDD.t148 VDD.n132 8.44573
R5207 VDD.n131 VDD.t122 8.44573
R5208 VDD.t122 VDD.n130 8.44573
R5209 VDD.n129 VDD.t200 8.44573
R5210 VDD.t200 VDD.n128 8.44573
R5211 VDD.n127 VDD.t66 8.44573
R5212 VDD.n247 VDD.t112 8.44573
R5213 VDD.t112 VDD.n223 8.44573
R5214 VDD.n222 VDD.t94 8.44573
R5215 VDD.t94 VDD.n221 8.44573
R5216 VDD.n220 VDD.t172 8.44573
R5217 VDD.t172 VDD.n219 8.44573
R5218 VDD.n218 VDD.t42 8.44573
R5219 VDD.n180 VDD.t124 8.44566
R5220 VDD.n271 VDD.t90 8.44566
R5221 VDD.t198 VDD.n170 8.44445
R5222 VDD.n171 VDD.t198 8.44445
R5223 VDD.t40 VDD.n172 8.44445
R5224 VDD.n173 VDD.t40 8.44445
R5225 VDD.t60 VDD.n174 8.44445
R5226 VDD.n175 VDD.t60 8.44445
R5227 VDD.t102 VDD.n176 8.44445
R5228 VDD.n177 VDD.t102 8.44445
R5229 VDD.n178 VDD.t124 8.44445
R5230 VDD.n146 VDD.t104 8.44445
R5231 VDD.n144 VDD.t104 8.44445
R5232 VDD.n143 VDD.t52 8.44445
R5233 VDD.n141 VDD.t52 8.44445
R5234 VDD.t110 VDD.n261 8.44445
R5235 VDD.n262 VDD.t110 8.44445
R5236 VDD.t190 VDD.n263 8.44445
R5237 VDD.n264 VDD.t190 8.44445
R5238 VDD.t86 VDD.n265 8.44445
R5239 VDD.n266 VDD.t86 8.44445
R5240 VDD.t194 VDD.n267 8.44445
R5241 VDD.n268 VDD.t194 8.44445
R5242 VDD.n269 VDD.t90 8.44445
R5243 VDD.n240 VDD.t244 8.44445
R5244 VDD.n238 VDD.t244 8.44445
R5245 VDD.n237 VDD.t80 8.44445
R5246 VDD.n235 VDD.t80 8.44445
R5247 VDD.n936 VDD.n557 8.2871
R5248 VDD.t127 VDD.n1209 8.13022
R5249 VDD.n1204 VDD.t105 8.13022
R5250 VDD.t151 VDD.n1170 8.13014
R5251 VDD.n1177 VDD.t47 8.13014
R5252 VDD.n1230 VDD.t261 8.10567
R5253 VDD.t261 VDD.n1229 8.10567
R5254 VDD.t239 VDD.n1227 8.10567
R5255 VDD.n1228 VDD.t239 8.10567
R5256 VDD.t215 VDD.n1225 8.10567
R5257 VDD.n1226 VDD.t215 8.10567
R5258 VDD.n1171 VDD.t151 8.10567
R5259 VDD.n1173 VDD.t115 8.10567
R5260 VDD.t115 VDD.n1172 8.10567
R5261 VDD.n1175 VDD.t83 8.10567
R5262 VDD.t83 VDD.n1174 8.10567
R5263 VDD.t47 VDD.n1176 8.10567
R5264 VDD.t173 VDD.n1213 8.10567
R5265 VDD.n1214 VDD.t173 8.10567
R5266 VDD.t157 VDD.n1211 8.10567
R5267 VDD.n1212 VDD.t157 8.10567
R5268 VDD.n1210 VDD.t127 8.10567
R5269 VDD.n1200 VDD.t163 8.10567
R5270 VDD.t163 VDD.n942 8.10567
R5271 VDD.n1202 VDD.t131 8.10567
R5272 VDD.t131 VDD.n1201 8.10567
R5273 VDD.t105 VDD.n1203 8.10567
R5274 VDD.n142 VDD.t51 7.36707
R5275 VDD.n145 VDD.t103 7.36707
R5276 VDD.n206 VDD.t65 7.36707
R5277 VDD.n199 VDD.t199 7.36707
R5278 VDD.n192 VDD.t121 7.36707
R5279 VDD.n185 VDD.t147 7.36707
R5280 VDD.n206 VDD.t207 7.36707
R5281 VDD.n199 VDD.t255 7.36707
R5282 VDD.n192 VDD.t177 7.36707
R5283 VDD.n185 VDD.t209 7.36707
R5284 VDD.n179 VDD.t123 7.36707
R5285 VDD.n157 VDD.t101 7.36707
R5286 VDD.n158 VDD.t59 7.36707
R5287 VDD.n159 VDD.t39 7.36707
R5288 VDD.n160 VDD.t197 7.36707
R5289 VDD.n236 VDD.t79 7.36707
R5290 VDD.n239 VDD.t243 7.36707
R5291 VDD.n297 VDD.t41 7.36707
R5292 VDD.n290 VDD.t171 7.36707
R5293 VDD.n283 VDD.t93 7.36707
R5294 VDD.n276 VDD.t111 7.36707
R5295 VDD.n297 VDD.t227 7.36707
R5296 VDD.n290 VDD.t129 7.36707
R5297 VDD.n283 VDD.t43 7.36707
R5298 VDD.n276 VDD.t61 7.36707
R5299 VDD.n270 VDD.t89 7.36707
R5300 VDD.n248 VDD.t193 7.36707
R5301 VDD.n249 VDD.t85 7.36707
R5302 VDD.n250 VDD.t189 7.36707
R5303 VDD.n251 VDD.t109 7.36707
R5304 VDD.n308 VDD.t187 7.36707
R5305 VDD.n114 VDD.t71 7.36707
R5306 VDD.n110 VDD.t233 7.36707
R5307 VDD.n98 VDD.t251 7.36707
R5308 VDD.n94 VDD.t231 7.36707
R5309 VDD.n82 VDD.t95 7.36707
R5310 VDD.n78 VDD.t229 7.36707
R5311 VDD.n405 VDD.t91 7.36707
R5312 VDD.n63 VDD.t249 7.36707
R5313 VDD.n434 VDD.t159 7.36707
R5314 VDD.n308 VDD.t75 7.36707
R5315 VDD.n114 VDD.t213 7.36707
R5316 VDD.n110 VDD.t141 7.36707
R5317 VDD.n98 VDD.t161 7.36707
R5318 VDD.n94 VDD.t137 7.36707
R5319 VDD.n82 VDD.t223 7.36707
R5320 VDD.n78 VDD.t133 7.36707
R5321 VDD.n405 VDD.t221 7.36707
R5322 VDD.n63 VDD.t153 7.36707
R5323 VDD.n434 VDD.t45 7.36707
R5324 VDD.n1061 VDD.t289 6.39714
R5325 VDD.n1056 VDD.t269 6.39714
R5326 VDD.n1038 VDD.t290 6.39714
R5327 VDD.n1033 VDD.t279 6.39714
R5328 VDD.n1009 VDD.t272 6.39714
R5329 VDD.n991 VDD.t285 6.39714
R5330 VDD.n986 VDD.t287 6.39714
R5331 VDD.n969 VDD.t283 6.39714
R5332 VDD.n963 VDD.t274 6.39714
R5333 VDD.n42 VDD.t21 6.09286
R5334 VDD.n10 VDD.t5 6.09286
R5335 VDD.n924 VDD.t35 5.8777
R5336 VDD.n35 VDD.t30 5.74671
R5337 VDD.n1014 VDD.t278 5.48273
R5338 VDD.n556 VDD.t11 5.47086
R5339 VDD.n555 VDD.t37 5.47086
R5340 VDD.n554 VDD.t15 5.47086
R5341 VDD.n36 VDD.t27 5.47086
R5342 VDD.n35 VDD.t31 5.47086
R5343 VDD.n43 VDD.t18 5.45468
R5344 VDD.n42 VDD.t17 5.45468
R5345 VDD.n10 VDD.t32 5.45468
R5346 VDD.n11 VDD.t12 5.45468
R5347 VDD.n1061 VDD.t282 5.45468
R5348 VDD.n1056 VDD.t280 5.45468
R5349 VDD.n1038 VDD.t273 5.45468
R5350 VDD.n1033 VDD.t284 5.45468
R5351 VDD.n1015 VDD.t275 5.45468
R5352 VDD.n1009 VDD.t277 5.45468
R5353 VDD.n991 VDD.t286 5.45468
R5354 VDD.n986 VDD.t288 5.45468
R5355 VDD.n969 VDD.t281 5.45468
R5356 VDD.n963 VDD.t276 5.45468
R5357 VDD.n205 VDD.n204 5.2005
R5358 VDD.n201 VDD.n200 5.2005
R5359 VDD.n198 VDD.n197 5.2005
R5360 VDD.n194 VDD.n193 5.2005
R5361 VDD.n191 VDD.n190 5.2005
R5362 VDD.n187 VDD.n186 5.2005
R5363 VDD.n183 VDD.n182 5.2005
R5364 VDD.n296 VDD.n295 5.2005
R5365 VDD.n292 VDD.n291 5.2005
R5366 VDD.n289 VDD.n288 5.2005
R5367 VDD.n285 VDD.n284 5.2005
R5368 VDD.n282 VDD.n281 5.2005
R5369 VDD.n278 VDD.n277 5.2005
R5370 VDD.n274 VDD.n273 5.2005
R5371 VDD.n313 VDD.n124 5.2005
R5372 VDD.n316 VDD.n121 5.2005
R5373 VDD.n324 VDD.n117 5.2005
R5374 VDD.n331 VDD.n113 5.2005
R5375 VDD.n340 VDD.n108 5.2005
R5376 VDD.n105 VDD.n104 5.2005
R5377 VDD.n351 VDD.n101 5.2005
R5378 VDD.n357 VDD.n97 5.2005
R5379 VDD.n366 VDD.n92 5.2005
R5380 VDD.n89 VDD.n88 5.2005
R5381 VDD.n377 VDD.n85 5.2005
R5382 VDD.n383 VDD.n81 5.2005
R5383 VDD.n394 VDD.n77 5.2005
R5384 VDD.n397 VDD.n74 5.2005
R5385 VDD.n404 VDD.n70 5.2005
R5386 VDD.n411 VDD.n66 5.2005
R5387 VDD.n421 VDD.n62 5.2005
R5388 VDD.n424 VDD.n59 5.2005
R5389 VDD.n432 VDD.n55 5.2005
R5390 VDD.n439 VDD.n51 5.2005
R5391 VDD.n314 VDD.n313 5.2005
R5392 VDD.n316 VDD.n315 5.2005
R5393 VDD.n324 VDD.n323 5.2005
R5394 VDD.n332 VDD.n331 5.2005
R5395 VDD.n341 VDD.n340 5.2005
R5396 VDD.n342 VDD.n104 5.2005
R5397 VDD.n351 VDD.n350 5.2005
R5398 VDD.n358 VDD.n357 5.2005
R5399 VDD.n367 VDD.n366 5.2005
R5400 VDD.n368 VDD.n88 5.2005
R5401 VDD.n377 VDD.n376 5.2005
R5402 VDD.n384 VDD.n383 5.2005
R5403 VDD.n395 VDD.n394 5.2005
R5404 VDD.n397 VDD.n396 5.2005
R5405 VDD.n404 VDD.n403 5.2005
R5406 VDD.n412 VDD.n411 5.2005
R5407 VDD.n422 VDD.n421 5.2005
R5408 VDD.n424 VDD.n423 5.2005
R5409 VDD.n432 VDD.n431 5.2005
R5410 VDD.n440 VDD.n439 5.2005
R5411 VDD.n440 VDD.t46 4.9005
R5412 VDD.n431 VDD.t46 4.9005
R5413 VDD.n423 VDD.t154 4.9005
R5414 VDD.t154 VDD.n422 4.9005
R5415 VDD.n412 VDD.t222 4.9005
R5416 VDD.n403 VDD.t222 4.9005
R5417 VDD.n396 VDD.t134 4.9005
R5418 VDD.t134 VDD.n395 4.9005
R5419 VDD.n384 VDD.t224 4.9005
R5420 VDD.n376 VDD.t224 4.9005
R5421 VDD.n368 VDD.t138 4.9005
R5422 VDD.t138 VDD.n367 4.9005
R5423 VDD.n358 VDD.t162 4.9005
R5424 VDD.n350 VDD.t162 4.9005
R5425 VDD.n342 VDD.t142 4.9005
R5426 VDD.t142 VDD.n341 4.9005
R5427 VDD.n332 VDD.t214 4.9005
R5428 VDD.n323 VDD.t214 4.9005
R5429 VDD.n315 VDD.t76 4.9005
R5430 VDD.t76 VDD.n314 4.9005
R5431 VDD.t160 VDD.n51 4.9005
R5432 VDD.n55 VDD.t160 4.9005
R5433 VDD.t250 VDD.n59 4.9005
R5434 VDD.n62 VDD.t250 4.9005
R5435 VDD.t92 VDD.n66 4.9005
R5436 VDD.n70 VDD.t92 4.9005
R5437 VDD.t230 VDD.n74 4.9005
R5438 VDD.n77 VDD.t230 4.9005
R5439 VDD.t96 VDD.n81 4.9005
R5440 VDD.n85 VDD.t96 4.9005
R5441 VDD.t232 VDD.n89 4.9005
R5442 VDD.n92 VDD.t232 4.9005
R5443 VDD.t252 VDD.n97 4.9005
R5444 VDD.n101 VDD.t252 4.9005
R5445 VDD.t234 VDD.n105 4.9005
R5446 VDD.n108 VDD.t234 4.9005
R5447 VDD.t72 VDD.n113 4.9005
R5448 VDD.n117 VDD.t72 4.9005
R5449 VDD.t188 VDD.n121 4.9005
R5450 VDD.n124 VDD.t188 4.9005
R5451 VDD.n182 VDD.t210 4.9005
R5452 VDD.n187 VDD.t210 4.9005
R5453 VDD.n190 VDD.t178 4.9005
R5454 VDD.n194 VDD.t178 4.9005
R5455 VDD.n197 VDD.t256 4.9005
R5456 VDD.n201 VDD.t256 4.9005
R5457 VDD.n204 VDD.t208 4.9005
R5458 VDD.n273 VDD.t62 4.9005
R5459 VDD.n278 VDD.t62 4.9005
R5460 VDD.n281 VDD.t44 4.9005
R5461 VDD.n285 VDD.t44 4.9005
R5462 VDD.n288 VDD.t130 4.9005
R5463 VDD.n292 VDD.t130 4.9005
R5464 VDD.n295 VDD.t228 4.9005
R5465 VDD.n26 VDD.n24 4.62286
R5466 VDD.n19 VDD.n17 4.62286
R5467 VDD.n5 VDD.n3 4.5005
R5468 VDD.n519 VDD.n518 4.5005
R5469 VDD.n521 VDD.n520 4.5005
R5470 VDD.n522 VDD.n517 4.5005
R5471 VDD.n524 VDD.n523 4.5005
R5472 VDD.n525 VDD.n516 4.5005
R5473 VDD.n527 VDD.n526 4.5005
R5474 VDD.n528 VDD.n514 4.5005
R5475 VDD.n530 VDD.n529 4.5005
R5476 VDD.n532 VDD.n16 4.5005
R5477 VDD.n534 VDD.n533 4.5005
R5478 VDD.n535 VDD.n15 4.5005
R5479 VDD.n537 VDD.n536 4.5005
R5480 VDD.n538 VDD.n14 4.5005
R5481 VDD.n540 VDD.n539 4.5005
R5482 VDD.n541 VDD.n13 4.5005
R5483 VDD.n543 VDD.n542 4.5005
R5484 VDD.n544 VDD.n9 4.5005
R5485 VDD.n546 VDD.n545 4.5005
R5486 VDD.n457 VDD.n22 4.5005
R5487 VDD.n459 VDD.n458 4.5005
R5488 VDD.n460 VDD.n456 4.5005
R5489 VDD.n462 VDD.n461 4.5005
R5490 VDD.n463 VDD.n455 4.5005
R5491 VDD.n465 VDD.n464 4.5005
R5492 VDD.n466 VDD.n454 4.5005
R5493 VDD.n468 VDD.n467 4.5005
R5494 VDD.n469 VDD.n45 4.5005
R5495 VDD.n471 VDD.n470 4.5005
R5496 VDD.n453 VDD.n44 4.5005
R5497 VDD.n452 VDD.n451 4.5005
R5498 VDD.n450 VDD.n46 4.5005
R5499 VDD.n449 VDD.n448 4.5005
R5500 VDD.n447 VDD.n47 4.5005
R5501 VDD.n446 VDD.n445 4.5005
R5502 VDD.n444 VDD.n48 4.5005
R5503 VDD.n443 VDD.n442 4.5005
R5504 VDD.n50 VDD.n49 4.5005
R5505 VDD.n438 VDD.n437 4.5005
R5506 VDD.n436 VDD.n435 4.5005
R5507 VDD.n433 VDD.n53 4.5005
R5508 VDD.n427 VDD.n54 4.5005
R5509 VDD.n429 VDD.n428 4.5005
R5510 VDD.n426 VDD.n425 4.5005
R5511 VDD.n58 VDD.n57 4.5005
R5512 VDD.n418 VDD.n417 4.5005
R5513 VDD.n420 VDD.n419 4.5005
R5514 VDD.n416 VDD.n61 4.5005
R5515 VDD.n415 VDD.n414 4.5005
R5516 VDD.n65 VDD.n64 4.5005
R5517 VDD.n410 VDD.n409 4.5005
R5518 VDD.n408 VDD.n67 4.5005
R5519 VDD.n407 VDD.n406 4.5005
R5520 VDD.n69 VDD.n68 4.5005
R5521 VDD.n401 VDD.n400 4.5005
R5522 VDD.n399 VDD.n398 4.5005
R5523 VDD.n73 VDD.n72 4.5005
R5524 VDD.n391 VDD.n390 4.5005
R5525 VDD.n393 VDD.n392 4.5005
R5526 VDD.n389 VDD.n76 4.5005
R5527 VDD.n388 VDD.n387 4.5005
R5528 VDD.n386 VDD.n79 4.5005
R5529 VDD.n380 VDD.n80 4.5005
R5530 VDD.n382 VDD.n381 4.5005
R5531 VDD.n379 VDD.n378 4.5005
R5532 VDD.n84 VDD.n83 4.5005
R5533 VDD.n374 VDD.n373 4.5005
R5534 VDD.n372 VDD.n86 4.5005
R5535 VDD.n371 VDD.n370 4.5005
R5536 VDD.n93 VDD.n87 4.5005
R5537 VDD.n365 VDD.n364 4.5005
R5538 VDD.n363 VDD.n91 4.5005
R5539 VDD.n362 VDD.n361 4.5005
R5540 VDD.n360 VDD.n95 4.5005
R5541 VDD.n354 VDD.n96 4.5005
R5542 VDD.n356 VDD.n355 4.5005
R5543 VDD.n353 VDD.n352 4.5005
R5544 VDD.n100 VDD.n99 4.5005
R5545 VDD.n348 VDD.n347 4.5005
R5546 VDD.n346 VDD.n102 4.5005
R5547 VDD.n345 VDD.n344 4.5005
R5548 VDD.n109 VDD.n103 4.5005
R5549 VDD.n339 VDD.n338 4.5005
R5550 VDD.n337 VDD.n107 4.5005
R5551 VDD.n336 VDD.n335 4.5005
R5552 VDD.n334 VDD.n111 4.5005
R5553 VDD.n328 VDD.n112 4.5005
R5554 VDD.n330 VDD.n329 4.5005
R5555 VDD.n327 VDD.n326 4.5005
R5556 VDD.n325 VDD.n115 4.5005
R5557 VDD.n319 VDD.n116 4.5005
R5558 VDD.n321 VDD.n320 4.5005
R5559 VDD.n318 VDD.n317 4.5005
R5560 VDD.n120 VDD.n119 4.5005
R5561 VDD.n310 VDD.n309 4.5005
R5562 VDD.n312 VDD.n311 4.5005
R5563 VDD.n307 VDD.n123 4.5005
R5564 VDD.n499 VDD.n498 4.5005
R5565 VDD.n500 VDD.n34 4.5005
R5566 VDD.n502 VDD.n501 4.5005
R5567 VDD.n503 VDD.n33 4.5005
R5568 VDD.n505 VDD.n504 4.5005
R5569 VDD.n506 VDD.n32 4.5005
R5570 VDD.n508 VDD.n507 4.5005
R5571 VDD.n509 VDD.n30 4.5005
R5572 VDD.n511 VDD.n510 4.5005
R5573 VDD.n477 VDD.n29 4.5005
R5574 VDD.n479 VDD.n478 4.5005
R5575 VDD.n480 VDD.n476 4.5005
R5576 VDD.n482 VDD.n481 4.5005
R5577 VDD.n483 VDD.n475 4.5005
R5578 VDD.n485 VDD.n484 4.5005
R5579 VDD.n486 VDD.n474 4.5005
R5580 VDD.n488 VDD.n487 4.5005
R5581 VDD.n489 VDD.n41 4.5005
R5582 VDD.n491 VDD.n490 4.5005
R5583 VDD.n497 VDD.n37 4.5005
R5584 VDD.n553 VDD.n552 4.5005
R5585 VDD.n894 VDD.n893 4.5005
R5586 VDD.n895 VDD.n571 4.5005
R5587 VDD.n898 VDD.n897 4.5005
R5588 VDD.n899 VDD.n570 4.5005
R5589 VDD.n901 VDD.n900 4.5005
R5590 VDD.n902 VDD.n569 4.5005
R5591 VDD.n904 VDD.n903 4.5005
R5592 VDD.n905 VDD.n567 4.5005
R5593 VDD.n907 VDD.n906 4.5005
R5594 VDD.n908 VDD.n566 4.5005
R5595 VDD.n910 VDD.n909 4.5005
R5596 VDD.n911 VDD.n564 4.5005
R5597 VDD.n913 VDD.n912 4.5005
R5598 VDD.n883 VDD.n576 4.5005
R5599 VDD.n883 VDD.n882 4.5005
R5600 VDD.n922 VDD.n921 4.5005
R5601 VDD.n935 VDD.n934 4.5005
R5602 VDD.n933 VDD.n558 4.5005
R5603 VDD.n932 VDD.n931 4.5005
R5604 VDD.n930 VDD.n560 4.5005
R5605 VDD.n929 VDD.n928 4.5005
R5606 VDD.n927 VDD.n561 4.5005
R5607 VDD.n926 VDD.n925 4.5005
R5608 VDD.n923 VDD.n563 4.5005
R5609 VDD.n1074 VDD.n1060 4.5005
R5610 VDD.n1076 VDD.n1075 4.5005
R5611 VDD.n1072 VDD.n1059 4.5005
R5612 VDD.n1071 VDD.n1070 4.5005
R5613 VDD.n1069 VDD.n1062 4.5005
R5614 VDD.n1067 VDD.n1066 4.5005
R5615 VDD.n1065 VDD.n1063 4.5005
R5616 VDD.n1064 VDD.n1058 4.5005
R5617 VDD.n1079 VDD.n1057 4.5005
R5618 VDD.n1081 VDD.n1080 4.5005
R5619 VDD.n1084 VDD.n1083 4.5005
R5620 VDD.n1085 VDD.n1054 4.5005
R5621 VDD.n1087 VDD.n1086 4.5005
R5622 VDD.n1089 VDD.n1088 4.5005
R5623 VDD.n1090 VDD.n1051 4.5005
R5624 VDD.n1092 VDD.n1091 4.5005
R5625 VDD.n1093 VDD.n1037 4.5005
R5626 VDD.n1095 VDD.n1094 4.5005
R5627 VDD.n1049 VDD.n1036 4.5005
R5628 VDD.n1048 VDD.n1047 4.5005
R5629 VDD.n1046 VDD.n1039 4.5005
R5630 VDD.n1044 VDD.n1043 4.5005
R5631 VDD.n1042 VDD.n1040 4.5005
R5632 VDD.n1041 VDD.n1035 4.5005
R5633 VDD.n1098 VDD.n1034 4.5005
R5634 VDD.n1100 VDD.n1099 4.5005
R5635 VDD.n1103 VDD.n1102 4.5005
R5636 VDD.n1104 VDD.n1031 4.5005
R5637 VDD.n1106 VDD.n1105 4.5005
R5638 VDD.n1108 VDD.n1107 4.5005
R5639 VDD.n1109 VDD.n1028 4.5005
R5640 VDD.n1111 VDD.n1110 4.5005
R5641 VDD.n1112 VDD.n1013 4.5005
R5642 VDD.n1114 VDD.n1113 4.5005
R5643 VDD.n1026 VDD.n1012 4.5005
R5644 VDD.n1025 VDD.n1024 4.5005
R5645 VDD.n1023 VDD.n1016 4.5005
R5646 VDD.n1021 VDD.n1020 4.5005
R5647 VDD.n1019 VDD.n1017 4.5005
R5648 VDD.n1018 VDD.n1011 4.5005
R5649 VDD.n1117 VDD.n1010 4.5005
R5650 VDD.n1119 VDD.n1118 4.5005
R5651 VDD.n1122 VDD.n1121 4.5005
R5652 VDD.n1123 VDD.n1007 4.5005
R5653 VDD.n1125 VDD.n1124 4.5005
R5654 VDD.n1127 VDD.n1126 4.5005
R5655 VDD.n1128 VDD.n1004 4.5005
R5656 VDD.n1130 VDD.n1129 4.5005
R5657 VDD.n1131 VDD.n990 4.5005
R5658 VDD.n1133 VDD.n1132 4.5005
R5659 VDD.n1002 VDD.n989 4.5005
R5660 VDD.n1001 VDD.n1000 4.5005
R5661 VDD.n999 VDD.n992 4.5005
R5662 VDD.n997 VDD.n996 4.5005
R5663 VDD.n995 VDD.n993 4.5005
R5664 VDD.n994 VDD.n988 4.5005
R5665 VDD.n1136 VDD.n987 4.5005
R5666 VDD.n1138 VDD.n1137 4.5005
R5667 VDD.n1141 VDD.n1140 4.5005
R5668 VDD.n1142 VDD.n984 4.5005
R5669 VDD.n1144 VDD.n1143 4.5005
R5670 VDD.n1146 VDD.n1145 4.5005
R5671 VDD.n1147 VDD.n981 4.5005
R5672 VDD.n1149 VDD.n1148 4.5005
R5673 VDD.n1150 VDD.n968 4.5005
R5674 VDD.n1152 VDD.n1151 4.5005
R5675 VDD.n979 VDD.n967 4.5005
R5676 VDD.n978 VDD.n977 4.5005
R5677 VDD.n976 VDD.n970 4.5005
R5678 VDD.n974 VDD.n973 4.5005
R5679 VDD.n972 VDD.n971 4.5005
R5680 VDD.n966 VDD.n965 4.5005
R5681 VDD.n1156 VDD.n1155 4.5005
R5682 VDD.n1157 VDD.n962 4.5005
R5683 VDD.n1159 VDD.n1158 4.5005
R5684 VDD.n1161 VDD.n961 4.5005
R5685 VDD.n1163 VDD.n1162 4.5005
R5686 VDD.n1165 VDD.n1164 4.5005
R5687 VDD.n1166 VDD.n959 4.5005
R5688 VDD.n1168 VDD.n1167 4.5005
R5689 VDD.n163 VDD.t74 4.22484
R5690 VDD.n162 VDD.t56 4.22484
R5691 VDD.n161 VDD.t166 4.22484
R5692 VDD.n212 VDD.t120 4.22484
R5693 VDD.n209 VDD.t118 4.22484
R5694 VDD.n154 VDD.t126 4.22484
R5695 VDD.n151 VDD.t180 4.22484
R5696 VDD.n148 VDD.t248 4.22484
R5697 VDD.n135 VDD.t238 4.22484
R5698 VDD.n134 VDD.t58 4.22484
R5699 VDD.n133 VDD.t140 4.22484
R5700 VDD.n259 VDD.t242 4.22484
R5701 VDD.n256 VDD.t226 4.22484
R5702 VDD.n253 VDD.t108 4.22484
R5703 VDD.n215 VDD.t260 4.22484
R5704 VDD.n214 VDD.t150 4.22484
R5705 VDD.n226 VDD.t254 4.22484
R5706 VDD.n225 VDD.t204 4.22484
R5707 VDD.n224 VDD.t144 4.22484
R5708 VDD.n233 VDD.t196 4.22484
R5709 VDD.n230 VDD.t146 4.22484
R5710 VDD.n227 VDD.t64 4.22484
R5711 VDD.n960 VDD.t219 4.05408
R5712 VDD.n975 VDD.t155 4.05408
R5713 VDD.n983 VDD.t169 4.05408
R5714 VDD.n998 VDD.t99 4.05408
R5715 VDD.n1006 VDD.t181 4.05408
R5716 VDD.n1022 VDD.t205 4.05408
R5717 VDD.n1030 VDD.t67 4.05408
R5718 VDD.n1045 VDD.t183 4.05408
R5719 VDD.n1053 VDD.t257 4.05408
R5720 VDD.n1068 VDD.t191 4.05408
R5721 VDD.n953 VDD.t135 4.05408
R5722 VDD.n952 VDD.t49 4.05408
R5723 VDD.n951 VDD.t69 4.05408
R5724 VDD.n950 VDD.t235 4.05408
R5725 VDD.n949 VDD.t77 4.05408
R5726 VDD.n948 VDD.t113 4.05408
R5727 VDD.n947 VDD.t217 4.05408
R5728 VDD.n1195 VDD.t211 4.05408
R5729 VDD.n1196 VDD.t245 4.05408
R5730 VDD.n946 VDD.t201 4.05408
R5731 VDD.n945 VDD.t53 4.05408
R5732 VDD.n944 VDD.t87 4.05408
R5733 VDD.n943 VDD.t185 4.05408
R5734 VDD.n946 VDD.t81 4.05408
R5735 VDD.n945 VDD.t167 4.05408
R5736 VDD.n944 VDD.t97 4.05408
R5737 VDD.n943 VDD.t175 4.05408
R5738 VDD.n28 VDD.n27 3.98468
R5739 VDD.n26 VDD.n25 3.98468
R5740 VDD.n19 VDD.n18 3.98468
R5741 VDD.n21 VDD.n20 3.98468
R5742 VDD.n1223 VDD.t176 3.20383
R5743 VDD.t176 VDD.n1222 3.20383
R5744 VDD.n1221 VDD.t98 3.20383
R5745 VDD.t98 VDD.n1220 3.20383
R5746 VDD.n1219 VDD.t168 3.20383
R5747 VDD.t168 VDD.n1218 3.20383
R5748 VDD.n1217 VDD.t82 3.20383
R5749 VDD.t82 VDD.n1216 3.20383
R5750 VDD.n1223 VDD.t186 3.20383
R5751 VDD.n1222 VDD.t186 3.20383
R5752 VDD.n1221 VDD.t88 3.20383
R5753 VDD.n1220 VDD.t88 3.20383
R5754 VDD.n1219 VDD.t54 3.20383
R5755 VDD.n1218 VDD.t54 3.20383
R5756 VDD.n1217 VDD.t202 3.20383
R5757 VDD.n1216 VDD.t202 3.20383
R5758 VDD.n1191 VDD.t218 3.20383
R5759 VDD.t218 VDD.n1190 3.20383
R5760 VDD.n1189 VDD.t114 3.20383
R5761 VDD.t114 VDD.n1188 3.20383
R5762 VDD.n1187 VDD.t78 3.20383
R5763 VDD.t78 VDD.n1186 3.20383
R5764 VDD.n1185 VDD.t236 3.20383
R5765 VDD.t236 VDD.n1184 3.20383
R5766 VDD.n1183 VDD.t70 3.20383
R5767 VDD.t70 VDD.n1182 3.20383
R5768 VDD.n1181 VDD.t50 3.20383
R5769 VDD.t50 VDD.n1180 3.20383
R5770 VDD.n1179 VDD.t136 3.20383
R5771 VDD.t136 VDD.n1178 3.20383
R5772 VDD.t192 VDD.n1077 3.20383
R5773 VDD.n1078 VDD.t192 3.20383
R5774 VDD.n1055 VDD.t258 3.20383
R5775 VDD.t258 VDD.n1052 3.20383
R5776 VDD.t184 VDD.n1096 3.20383
R5777 VDD.n1097 VDD.t184 3.20383
R5778 VDD.n1032 VDD.t68 3.20383
R5779 VDD.t68 VDD.n1029 3.20383
R5780 VDD.t206 VDD.n1115 3.20383
R5781 VDD.n1116 VDD.t206 3.20383
R5782 VDD.n1008 VDD.t182 3.20383
R5783 VDD.t182 VDD.n1005 3.20383
R5784 VDD.t100 VDD.n1134 3.20383
R5785 VDD.n1135 VDD.t100 3.20383
R5786 VDD.n985 VDD.t170 3.20383
R5787 VDD.t170 VDD.n982 3.20383
R5788 VDD.t156 VDD.n1153 3.20383
R5789 VDD.n1154 VDD.t156 3.20383
R5790 VDD.n1160 VDD.t220 3.20383
R5791 VDD.t220 VDD.n958 3.20383
R5792 VDD.t246 VDD.n1205 3.20383
R5793 VDD.n1206 VDD.t246 3.20383
R5794 VDD.t212 VDD.n1207 3.20383
R5795 VDD.n1208 VDD.t212 3.20383
R5796 VDD.n496 VDD.n38 2.62234
R5797 VDD.n492 VDD.n38 2.62234
R5798 VDD.n551 VDD.n6 2.62234
R5799 VDD.n547 VDD.n6 2.62234
R5800 VDD.n896 VDD.t2 2.38623
R5801 VDD.n1169 VDD.n1168 2.27786
R5802 VDD.n306 VDD.n122 2.25958
R5803 VDD.n702 VDD.n639 2.2505
R5804 VDD.n703 VDD.n638 2.2505
R5805 VDD.n705 VDD.n704 2.2505
R5806 VDD.n706 VDD.n637 2.2505
R5807 VDD.n708 VDD.n707 2.2505
R5808 VDD.n709 VDD.n636 2.2505
R5809 VDD.n711 VDD.n710 2.2505
R5810 VDD.n712 VDD.n635 2.2505
R5811 VDD.n714 VDD.n713 2.2505
R5812 VDD.n715 VDD.n634 2.2505
R5813 VDD.n717 VDD.n716 2.2505
R5814 VDD.n718 VDD.n633 2.2505
R5815 VDD.n720 VDD.n719 2.2505
R5816 VDD.n721 VDD.n632 2.2505
R5817 VDD.n723 VDD.n722 2.2505
R5818 VDD.n724 VDD.n631 2.2505
R5819 VDD.n726 VDD.n725 2.2505
R5820 VDD.n727 VDD.n630 2.2505
R5821 VDD.n729 VDD.n728 2.2505
R5822 VDD.n730 VDD.n629 2.2505
R5823 VDD.n732 VDD.n731 2.2505
R5824 VDD.n733 VDD.n628 2.2505
R5825 VDD.n735 VDD.n734 2.2505
R5826 VDD.n736 VDD.n627 2.2505
R5827 VDD.n738 VDD.n737 2.2505
R5828 VDD.n739 VDD.n626 2.2505
R5829 VDD.n741 VDD.n740 2.2505
R5830 VDD.n742 VDD.n625 2.2505
R5831 VDD.n744 VDD.n743 2.2505
R5832 VDD.n745 VDD.n624 2.2505
R5833 VDD.n747 VDD.n746 2.2505
R5834 VDD.n748 VDD.n623 2.2505
R5835 VDD.n750 VDD.n749 2.2505
R5836 VDD.n751 VDD.n622 2.2505
R5837 VDD.n753 VDD.n752 2.2505
R5838 VDD.n754 VDD.n621 2.2505
R5839 VDD.n756 VDD.n755 2.2505
R5840 VDD.n757 VDD.n620 2.2505
R5841 VDD.n759 VDD.n758 2.2505
R5842 VDD.n760 VDD.n619 2.2505
R5843 VDD.n762 VDD.n761 2.2505
R5844 VDD.n763 VDD.n618 2.2505
R5845 VDD.n765 VDD.n764 2.2505
R5846 VDD.n766 VDD.n617 2.2505
R5847 VDD.n768 VDD.n767 2.2505
R5848 VDD.n769 VDD.n616 2.2505
R5849 VDD.n771 VDD.n770 2.2505
R5850 VDD.n772 VDD.n615 2.2505
R5851 VDD.n774 VDD.n773 2.2505
R5852 VDD.n775 VDD.n614 2.2505
R5853 VDD.n777 VDD.n776 2.2505
R5854 VDD.n778 VDD.n613 2.2505
R5855 VDD.n780 VDD.n779 2.2505
R5856 VDD.n781 VDD.n612 2.2505
R5857 VDD.n783 VDD.n782 2.2505
R5858 VDD.n784 VDD.n611 2.2505
R5859 VDD.n786 VDD.n785 2.2505
R5860 VDD.n787 VDD.n610 2.2505
R5861 VDD.n789 VDD.n788 2.2505
R5862 VDD.n790 VDD.n609 2.2505
R5863 VDD.n792 VDD.n791 2.2505
R5864 VDD.n793 VDD.n608 2.2505
R5865 VDD.n795 VDD.n794 2.2505
R5866 VDD.n796 VDD.n607 2.2505
R5867 VDD.n798 VDD.n797 2.2505
R5868 VDD.n799 VDD.n606 2.2505
R5869 VDD.n801 VDD.n800 2.2505
R5870 VDD.n802 VDD.n605 2.2505
R5871 VDD.n804 VDD.n803 2.2505
R5872 VDD.n805 VDD.n604 2.2505
R5873 VDD.n807 VDD.n806 2.2505
R5874 VDD.n808 VDD.n603 2.2505
R5875 VDD.n810 VDD.n809 2.2505
R5876 VDD.n811 VDD.n602 2.2505
R5877 VDD.n813 VDD.n812 2.2505
R5878 VDD.n814 VDD.n601 2.2505
R5879 VDD.n816 VDD.n815 2.2505
R5880 VDD.n817 VDD.n600 2.2505
R5881 VDD.n819 VDD.n818 2.2505
R5882 VDD.n820 VDD.n599 2.2505
R5883 VDD.n822 VDD.n821 2.2505
R5884 VDD.n823 VDD.n598 2.2505
R5885 VDD.n825 VDD.n824 2.2505
R5886 VDD.n826 VDD.n597 2.2505
R5887 VDD.n828 VDD.n827 2.2505
R5888 VDD.n829 VDD.n596 2.2505
R5889 VDD.n831 VDD.n830 2.2505
R5890 VDD.n832 VDD.n595 2.2505
R5891 VDD.n834 VDD.n833 2.2505
R5892 VDD.n835 VDD.n594 2.2505
R5893 VDD.n837 VDD.n836 2.2505
R5894 VDD.n838 VDD.n593 2.2505
R5895 VDD.n840 VDD.n839 2.2505
R5896 VDD.n841 VDD.n592 2.2505
R5897 VDD.n843 VDD.n842 2.2505
R5898 VDD.n844 VDD.n591 2.2505
R5899 VDD.n846 VDD.n845 2.2505
R5900 VDD.n847 VDD.n590 2.2505
R5901 VDD.n849 VDD.n848 2.2505
R5902 VDD.n850 VDD.n589 2.2505
R5903 VDD.n852 VDD.n851 2.2505
R5904 VDD.n853 VDD.n588 2.2505
R5905 VDD.n855 VDD.n854 2.2505
R5906 VDD.n856 VDD.n587 2.2505
R5907 VDD.n858 VDD.n857 2.2505
R5908 VDD.n859 VDD.n586 2.2505
R5909 VDD.n861 VDD.n860 2.2505
R5910 VDD.n862 VDD.n585 2.2505
R5911 VDD.n864 VDD.n863 2.2505
R5912 VDD.n865 VDD.n584 2.2505
R5913 VDD.n867 VDD.n866 2.2505
R5914 VDD.n868 VDD.n583 2.2505
R5915 VDD.n870 VDD.n869 2.2505
R5916 VDD.n881 VDD.n574 2.2505
R5917 VDD.n880 VDD.n879 2.2505
R5918 VDD.n878 VDD.n578 2.2505
R5919 VDD.n877 VDD.n876 2.2505
R5920 VDD.n875 VDD.n579 2.2505
R5921 VDD.n874 VDD.n873 2.2505
R5922 VDD.n581 VDD.n580 2.2505
R5923 VDD.n656 VDD.n655 2.2505
R5924 VDD.n657 VDD.n654 2.2505
R5925 VDD.n659 VDD.n658 2.2505
R5926 VDD.n660 VDD.n653 2.2505
R5927 VDD.n662 VDD.n661 2.2505
R5928 VDD.n663 VDD.n652 2.2505
R5929 VDD.n665 VDD.n664 2.2505
R5930 VDD.n666 VDD.n651 2.2505
R5931 VDD.n668 VDD.n667 2.2505
R5932 VDD.n669 VDD.n650 2.2505
R5933 VDD.n671 VDD.n670 2.2505
R5934 VDD.n672 VDD.n649 2.2505
R5935 VDD.n674 VDD.n673 2.2505
R5936 VDD.n675 VDD.n648 2.2505
R5937 VDD.n677 VDD.n676 2.2505
R5938 VDD.n678 VDD.n647 2.2505
R5939 VDD.n680 VDD.n679 2.2505
R5940 VDD.n681 VDD.n646 2.2505
R5941 VDD.n683 VDD.n682 2.2505
R5942 VDD.n684 VDD.n645 2.2505
R5943 VDD.n686 VDD.n685 2.2505
R5944 VDD.n687 VDD.n644 2.2505
R5945 VDD.n689 VDD.n688 2.2505
R5946 VDD.n690 VDD.n643 2.2505
R5947 VDD.n692 VDD.n691 2.2505
R5948 VDD.n693 VDD.n642 2.2505
R5949 VDD.n695 VDD.n694 2.2505
R5950 VDD.n696 VDD.n641 2.2505
R5951 VDD.n698 VDD.n697 2.2505
R5952 VDD.n699 VDD.n640 2.2505
R5953 VDD.n701 VDD.n700 2.2505
R5954 VDD.n885 VDD.n573 2.24111
R5955 VDD.n883 VDD.n577 2.24111
R5956 VDD.n885 VDD.n572 2.24111
R5957 VDD.n306 VDD.n304 2.17535
R5958 VDD.n306 VDD.n305 2.17535
R5959 VDD.n1 VDD.n0 1.85588
R5960 VDD.n872 VDD.n871 1.84648
R5961 VDD.n892 VDD.n886 1.61339
R5962 VDD.n886 VDD.n565 1.61339
R5963 VDD.n939 VDD.t262 1.60217
R5964 VDD.n940 VDD.t240 1.60217
R5965 VDD.n941 VDD.t216 1.60217
R5966 VDD.n957 VDD.t152 1.60217
R5967 VDD.n956 VDD.t116 1.60217
R5968 VDD.n955 VDD.t84 1.60217
R5969 VDD.n954 VDD.t48 1.60217
R5970 VDD.n1192 VDD.t174 1.60217
R5971 VDD.n1193 VDD.t158 1.60217
R5972 VDD.n1194 VDD.t128 1.60217
R5973 VDD.n1199 VDD.t164 1.60217
R5974 VDD.n1198 VDD.t132 1.60217
R5975 VDD.n1197 VDD.t106 1.60217
R5976 VDD.n497 VDD.n496 1.59191
R5977 VDD.n492 VDD.n491 1.59191
R5978 VDD.n552 VDD.n551 1.59191
R5979 VDD.n547 VDD.n546 1.59191
R5980 VDD.n1073 VDD.n1061 1.05137
R5981 VDD.n1082 VDD.n1056 1.05137
R5982 VDD.n1050 VDD.n1038 1.05137
R5983 VDD.n1101 VDD.n1033 1.05137
R5984 VDD.n1027 VDD.n1015 1.05137
R5985 VDD.n1120 VDD.n1009 1.05137
R5986 VDD.n1003 VDD.n991 1.05137
R5987 VDD.n1139 VDD.n986 1.05137
R5988 VDD.n980 VDD.n969 1.05137
R5989 VDD.n964 VDD.n963 1.05137
R5990 VDD.n920 VDD.n919 1.0505
R5991 VDD.n916 VDD.n559 1.0505
R5992 VDD.n920 VDD.n914 1.02129
R5993 VDD.n914 VDD.n559 1.02129
R5994 VDD.n557 VDD.n556 0.998076
R5995 VDD.n1015 VDD.n1014 0.914916
R5996 VDD.n27 VDD.t20 0.9105
R5997 VDD.n27 VDD.t25 0.9105
R5998 VDD.n25 VDD.t28 0.9105
R5999 VDD.n25 VDD.t24 0.9105
R6000 VDD.n24 VDD.t22 0.9105
R6001 VDD.n24 VDD.t29 0.9105
R6002 VDD.n17 VDD.t7 0.9105
R6003 VDD.n17 VDD.t9 0.9105
R6004 VDD.n18 VDD.t33 0.9105
R6005 VDD.n18 VDD.t36 0.9105
R6006 VDD.n20 VDD.t13 0.9105
R6007 VDD.n20 VDD.t14 0.9105
R6008 VDD.n917 VDD.n914 0.9005
R6009 VDD.n928 VDD.n562 0.9005
R6010 VDD.n893 VDD.n892 0.857079
R6011 VDD.n912 VDD.n565 0.857079
R6012 VDD.n918 VDD.t34 0.767069
R6013 VDD.n915 VDD.t34 0.767069
R6014 VDD.n936 VDD.n935 0.759875
R6015 VDD.n457 VDD.n23 0.653559
R6016 VDD.n43 VDD.n42 0.638674
R6017 VDD.n11 VDD.n10 0.638674
R6018 VDD.n21 VDD.n19 0.638674
R6019 VDD.n28 VDD.n26 0.638674
R6020 VDD.n473 VDD.n43 0.577801
R6021 VDD.n12 VDD.n11 0.577801
R6022 VDD.n531 VDD.n21 0.577801
R6023 VDD.n512 VDD.n28 0.577801
R6024 VDD.n889 VDD.n886 0.573227
R6025 VDD.n904 VDD.n568 0.573227
R6026 VDD VDD.n937 0.53378
R6027 VDD.n892 VDD.n891 0.5255
R6028 VDD.n888 VDD.n565 0.5255
R6029 VDD.n921 VDD.n920 0.51112
R6030 VDD.n934 VDD.n559 0.51112
R6031 VDD.n513 VDD.n23 0.464857
R6032 VDD.n890 VDD.t1 0.443525
R6033 VDD.n887 VDD.t1 0.443525
R6034 VDD.n531 VDD.n513 0.443
R6035 VDD.n472 VDD.n12 0.443
R6036 VDD.n473 VDD.n472 0.443
R6037 VDD.n513 VDD.n512 0.443
R6038 VDD.n23 VDD.n4 0.430752
R6039 VDD.n496 VDD.n495 0.332079
R6040 VDD.n493 VDD.n492 0.332079
R6041 VDD.n551 VDD.n550 0.332079
R6042 VDD.n548 VDD.n547 0.332079
R6043 VDD.n40 VDD.n38 0.274413
R6044 VDD.n494 VDD.n40 0.274413
R6045 VDD.n39 VDD.n31 0.274413
R6046 VDD.n494 VDD.n39 0.274413
R6047 VDD.n7 VDD.n6 0.274413
R6048 VDD.n549 VDD.n7 0.274413
R6049 VDD.n515 VDD.n8 0.274413
R6050 VDD.n549 VDD.n8 0.274413
R6051 VDD.n556 VDD.n555 0.269452
R6052 VDD.n555 VDD.n554 0.269452
R6053 VDD.n36 VDD.n35 0.269452
R6054 VDD.n554 VDD.n553 0.262326
R6055 VDD.n37 VDD.n36 0.262326
R6056 VDD.n700 VDD.n639 0.240125
R6057 VDD.n702 VDD.n701 0.240125
R6058 VDD.n869 VDD.n582 0.234368
R6059 VDD.n894 VDD.n885 0.233375
R6060 VDD.n576 VDD.n575 0.229823
R6061 VDD.n553 VDD.n4 0.22415
R6062 VDD.n37 VDD.n4 0.22415
R6063 VDD.n884 VDD.n575 0.216513
R6064 VDD.n871 VDD.n582 0.214494
R6065 VDD.n922 VDD.n913 0.188825
R6066 VDD.n2 VDD.n0 0.168962
R6067 VDD.n915 VDD.n562 0.133266
R6068 VDD.n918 VDD.n917 0.133266
R6069 VDD.n887 VDD.n568 0.130545
R6070 VDD.n890 VDD.n889 0.130545
R6071 VDD.n557 VDD.n2 0.118192
R6072 VDD.n934 VDD.n933 0.114071
R6073 VDD.n933 VDD.n932 0.114071
R6074 VDD.n932 VDD.n560 0.114071
R6075 VDD.n928 VDD.n560 0.114071
R6076 VDD.n928 VDD.n927 0.114071
R6077 VDD.n927 VDD.n926 0.114071
R6078 VDD.n926 VDD.n563 0.114071
R6079 VDD.n921 VDD.n563 0.114071
R6080 VDD.n912 VDD.n911 0.114071
R6081 VDD.n911 VDD.n910 0.114071
R6082 VDD.n910 VDD.n566 0.114071
R6083 VDD.n906 VDD.n566 0.114071
R6084 VDD.n906 VDD.n905 0.114071
R6085 VDD.n905 VDD.n904 0.114071
R6086 VDD.n904 VDD.n569 0.114071
R6087 VDD.n900 VDD.n569 0.114071
R6088 VDD.n900 VDD.n899 0.114071
R6089 VDD.n899 VDD.n898 0.114071
R6090 VDD.n898 VDD.n571 0.114071
R6091 VDD.n893 VDD.n571 0.114071
R6092 VDD.n491 VDD.n41 0.114071
R6093 VDD.n487 VDD.n41 0.114071
R6094 VDD.n487 VDD.n486 0.114071
R6095 VDD.n486 VDD.n485 0.114071
R6096 VDD.n485 VDD.n475 0.114071
R6097 VDD.n481 VDD.n475 0.114071
R6098 VDD.n481 VDD.n480 0.114071
R6099 VDD.n480 VDD.n479 0.114071
R6100 VDD.n479 VDD.n477 0.114071
R6101 VDD.n510 VDD.n509 0.114071
R6102 VDD.n509 VDD.n508 0.114071
R6103 VDD.n508 VDD.n32 0.114071
R6104 VDD.n504 VDD.n32 0.114071
R6105 VDD.n504 VDD.n503 0.114071
R6106 VDD.n503 VDD.n502 0.114071
R6107 VDD.n502 VDD.n34 0.114071
R6108 VDD.n498 VDD.n34 0.114071
R6109 VDD.n498 VDD.n497 0.114071
R6110 VDD.n447 VDD.n446 0.114071
R6111 VDD.n448 VDD.n447 0.114071
R6112 VDD.n448 VDD.n46 0.114071
R6113 VDD.n452 VDD.n46 0.114071
R6114 VDD.n453 VDD.n452 0.114071
R6115 VDD.n470 VDD.n453 0.114071
R6116 VDD.n470 VDD.n469 0.114071
R6117 VDD.n469 VDD.n468 0.114071
R6118 VDD.n468 VDD.n454 0.114071
R6119 VDD.n464 VDD.n454 0.114071
R6120 VDD.n464 VDD.n463 0.114071
R6121 VDD.n463 VDD.n462 0.114071
R6122 VDD.n462 VDD.n456 0.114071
R6123 VDD.n458 VDD.n456 0.114071
R6124 VDD.n458 VDD.n457 0.114071
R6125 VDD.n546 VDD.n9 0.114071
R6126 VDD.n542 VDD.n9 0.114071
R6127 VDD.n542 VDD.n541 0.114071
R6128 VDD.n541 VDD.n540 0.114071
R6129 VDD.n540 VDD.n14 0.114071
R6130 VDD.n536 VDD.n14 0.114071
R6131 VDD.n536 VDD.n535 0.114071
R6132 VDD.n535 VDD.n534 0.114071
R6133 VDD.n534 VDD.n16 0.114071
R6134 VDD.n529 VDD.n528 0.114071
R6135 VDD.n528 VDD.n527 0.114071
R6136 VDD.n527 VDD.n516 0.114071
R6137 VDD.n523 VDD.n516 0.114071
R6138 VDD.n523 VDD.n522 0.114071
R6139 VDD.n522 VDD.n521 0.114071
R6140 VDD.n521 VDD.n518 0.114071
R6141 VDD.n518 VDD.n5 0.114071
R6142 VDD.n552 VDD.n5 0.114071
R6143 VDD.n545 VDD.n544 0.114071
R6144 VDD.n544 VDD.n543 0.114071
R6145 VDD.n543 VDD.n13 0.114071
R6146 VDD.n539 VDD.n13 0.114071
R6147 VDD.n539 VDD.n538 0.114071
R6148 VDD.n538 VDD.n537 0.114071
R6149 VDD.n537 VDD.n15 0.114071
R6150 VDD.n533 VDD.n15 0.114071
R6151 VDD.n533 VDD.n532 0.114071
R6152 VDD.n530 VDD.n514 0.114071
R6153 VDD.n526 VDD.n514 0.114071
R6154 VDD.n526 VDD.n525 0.114071
R6155 VDD.n525 VDD.n524 0.114071
R6156 VDD.n524 VDD.n517 0.114071
R6157 VDD.n520 VDD.n517 0.114071
R6158 VDD.n520 VDD.n519 0.114071
R6159 VDD.n519 VDD.n3 0.114071
R6160 VDD.n311 VDD.n307 0.114071
R6161 VDD.n311 VDD.n310 0.114071
R6162 VDD.n310 VDD.n119 0.114071
R6163 VDD.n318 VDD.n119 0.114071
R6164 VDD.n320 VDD.n318 0.114071
R6165 VDD.n320 VDD.n319 0.114071
R6166 VDD.n319 VDD.n115 0.114071
R6167 VDD.n327 VDD.n115 0.114071
R6168 VDD.n329 VDD.n327 0.114071
R6169 VDD.n329 VDD.n328 0.114071
R6170 VDD.n328 VDD.n111 0.114071
R6171 VDD.n336 VDD.n111 0.114071
R6172 VDD.n337 VDD.n336 0.114071
R6173 VDD.n338 VDD.n337 0.114071
R6174 VDD.n338 VDD.n103 0.114071
R6175 VDD.n345 VDD.n103 0.114071
R6176 VDD.n346 VDD.n345 0.114071
R6177 VDD.n347 VDD.n346 0.114071
R6178 VDD.n347 VDD.n99 0.114071
R6179 VDD.n353 VDD.n99 0.114071
R6180 VDD.n355 VDD.n353 0.114071
R6181 VDD.n355 VDD.n354 0.114071
R6182 VDD.n354 VDD.n95 0.114071
R6183 VDD.n362 VDD.n95 0.114071
R6184 VDD.n363 VDD.n362 0.114071
R6185 VDD.n364 VDD.n363 0.114071
R6186 VDD.n364 VDD.n87 0.114071
R6187 VDD.n371 VDD.n87 0.114071
R6188 VDD.n372 VDD.n371 0.114071
R6189 VDD.n373 VDD.n372 0.114071
R6190 VDD.n373 VDD.n83 0.114071
R6191 VDD.n379 VDD.n83 0.114071
R6192 VDD.n381 VDD.n379 0.114071
R6193 VDD.n381 VDD.n380 0.114071
R6194 VDD.n380 VDD.n79 0.114071
R6195 VDD.n388 VDD.n79 0.114071
R6196 VDD.n389 VDD.n388 0.114071
R6197 VDD.n392 VDD.n389 0.114071
R6198 VDD.n392 VDD.n391 0.114071
R6199 VDD.n391 VDD.n72 0.114071
R6200 VDD.n399 VDD.n72 0.114071
R6201 VDD.n400 VDD.n399 0.114071
R6202 VDD.n400 VDD.n68 0.114071
R6203 VDD.n407 VDD.n68 0.114071
R6204 VDD.n408 VDD.n407 0.114071
R6205 VDD.n409 VDD.n408 0.114071
R6206 VDD.n409 VDD.n64 0.114071
R6207 VDD.n415 VDD.n64 0.114071
R6208 VDD.n416 VDD.n415 0.114071
R6209 VDD.n419 VDD.n416 0.114071
R6210 VDD.n419 VDD.n418 0.114071
R6211 VDD.n418 VDD.n57 0.114071
R6212 VDD.n426 VDD.n57 0.114071
R6213 VDD.n428 VDD.n426 0.114071
R6214 VDD.n428 VDD.n427 0.114071
R6215 VDD.n427 VDD.n53 0.114071
R6216 VDD.n436 VDD.n53 0.114071
R6217 VDD.n437 VDD.n436 0.114071
R6218 VDD.n437 VDD.n49 0.114071
R6219 VDD.n443 VDD.n49 0.114071
R6220 VDD.n444 VDD.n443 0.114071
R6221 VDD.n445 VDD.n444 0.114071
R6222 VDD.n445 VDD.n47 0.114071
R6223 VDD.n449 VDD.n47 0.114071
R6224 VDD.n450 VDD.n449 0.114071
R6225 VDD.n451 VDD.n450 0.114071
R6226 VDD.n451 VDD.n44 0.114071
R6227 VDD.n471 VDD.n45 0.114071
R6228 VDD.n467 VDD.n45 0.114071
R6229 VDD.n467 VDD.n466 0.114071
R6230 VDD.n466 VDD.n465 0.114071
R6231 VDD.n465 VDD.n455 0.114071
R6232 VDD.n461 VDD.n455 0.114071
R6233 VDD.n461 VDD.n460 0.114071
R6234 VDD.n460 VDD.n459 0.114071
R6235 VDD.n459 VDD.n22 0.114071
R6236 VDD.n490 VDD.n489 0.114071
R6237 VDD.n489 VDD.n488 0.114071
R6238 VDD.n488 VDD.n474 0.114071
R6239 VDD.n484 VDD.n474 0.114071
R6240 VDD.n484 VDD.n483 0.114071
R6241 VDD.n483 VDD.n482 0.114071
R6242 VDD.n482 VDD.n476 0.114071
R6243 VDD.n478 VDD.n476 0.114071
R6244 VDD.n478 VDD.n29 0.114071
R6245 VDD.n511 VDD.n30 0.114071
R6246 VDD.n507 VDD.n30 0.114071
R6247 VDD.n507 VDD.n506 0.114071
R6248 VDD.n506 VDD.n505 0.114071
R6249 VDD.n505 VDD.n33 0.114071
R6250 VDD.n501 VDD.n33 0.114071
R6251 VDD.n501 VDD.n500 0.114071
R6252 VDD.n500 VDD.n499 0.114071
R6253 VDD.n937 VDD.n936 0.11015
R6254 VDD.n1074 VDD.n937 0.10822
R6255 VDD.n553 VDD.n3 0.104429
R6256 VDD.n499 VDD.n37 0.104429
R6257 VDD.n307 VDD.n306 0.0926429
R6258 VDD.n472 VDD.n471 0.068
R6259 VDD.n477 VDD.n31 0.0572857
R6260 VDD.n510 VDD.n31 0.0572857
R6261 VDD.n515 VDD.n16 0.0572857
R6262 VDD.n529 VDD.n515 0.0572857
R6263 VDD.n532 VDD.n531 0.0572857
R6264 VDD.n531 VDD.n530 0.0572857
R6265 VDD.n512 VDD.n29 0.0572857
R6266 VDD.n512 VDD.n511 0.0572857
R6267 VDD.n446 VDD.n48 0.0527041
R6268 VDD.n472 VDD.n44 0.0465714
R6269 VDD.n577 VDD.n572 0.0410752
R6270 VDD.n577 VDD.n573 0.0410752
R6271 VDD.n700 VDD.n699 0.04025
R6272 VDD.n699 VDD.n698 0.04025
R6273 VDD.n698 VDD.n641 0.04025
R6274 VDD.n694 VDD.n641 0.04025
R6275 VDD.n694 VDD.n693 0.04025
R6276 VDD.n693 VDD.n692 0.04025
R6277 VDD.n692 VDD.n643 0.04025
R6278 VDD.n688 VDD.n643 0.04025
R6279 VDD.n688 VDD.n687 0.04025
R6280 VDD.n687 VDD.n686 0.04025
R6281 VDD.n686 VDD.n645 0.04025
R6282 VDD.n682 VDD.n645 0.04025
R6283 VDD.n682 VDD.n681 0.04025
R6284 VDD.n681 VDD.n680 0.04025
R6285 VDD.n680 VDD.n647 0.04025
R6286 VDD.n676 VDD.n647 0.04025
R6287 VDD.n676 VDD.n675 0.04025
R6288 VDD.n675 VDD.n674 0.04025
R6289 VDD.n674 VDD.n649 0.04025
R6290 VDD.n670 VDD.n649 0.04025
R6291 VDD.n670 VDD.n669 0.04025
R6292 VDD.n669 VDD.n668 0.04025
R6293 VDD.n668 VDD.n651 0.04025
R6294 VDD.n664 VDD.n651 0.04025
R6295 VDD.n664 VDD.n663 0.04025
R6296 VDD.n663 VDD.n662 0.04025
R6297 VDD.n662 VDD.n653 0.04025
R6298 VDD.n658 VDD.n653 0.04025
R6299 VDD.n658 VDD.n657 0.04025
R6300 VDD.n657 VDD.n656 0.04025
R6301 VDD.n656 VDD.n580 0.04025
R6302 VDD.n874 VDD.n580 0.04025
R6303 VDD.n875 VDD.n874 0.04025
R6304 VDD.n876 VDD.n875 0.04025
R6305 VDD.n876 VDD.n578 0.04025
R6306 VDD.n880 VDD.n578 0.04025
R6307 VDD.n881 VDD.n880 0.04025
R6308 VDD.n882 VDD.n881 0.04025
R6309 VDD.n869 VDD.n868 0.04025
R6310 VDD.n868 VDD.n867 0.04025
R6311 VDD.n867 VDD.n584 0.04025
R6312 VDD.n863 VDD.n584 0.04025
R6313 VDD.n863 VDD.n862 0.04025
R6314 VDD.n862 VDD.n861 0.04025
R6315 VDD.n861 VDD.n586 0.04025
R6316 VDD.n857 VDD.n586 0.04025
R6317 VDD.n857 VDD.n856 0.04025
R6318 VDD.n856 VDD.n855 0.04025
R6319 VDD.n855 VDD.n588 0.04025
R6320 VDD.n851 VDD.n588 0.04025
R6321 VDD.n851 VDD.n850 0.04025
R6322 VDD.n850 VDD.n849 0.04025
R6323 VDD.n849 VDD.n590 0.04025
R6324 VDD.n845 VDD.n590 0.04025
R6325 VDD.n845 VDD.n844 0.04025
R6326 VDD.n844 VDD.n843 0.04025
R6327 VDD.n843 VDD.n592 0.04025
R6328 VDD.n839 VDD.n592 0.04025
R6329 VDD.n839 VDD.n838 0.04025
R6330 VDD.n838 VDD.n837 0.04025
R6331 VDD.n837 VDD.n594 0.04025
R6332 VDD.n833 VDD.n594 0.04025
R6333 VDD.n833 VDD.n832 0.04025
R6334 VDD.n832 VDD.n831 0.04025
R6335 VDD.n831 VDD.n596 0.04025
R6336 VDD.n827 VDD.n596 0.04025
R6337 VDD.n827 VDD.n826 0.04025
R6338 VDD.n826 VDD.n825 0.04025
R6339 VDD.n825 VDD.n598 0.04025
R6340 VDD.n821 VDD.n598 0.04025
R6341 VDD.n821 VDD.n820 0.04025
R6342 VDD.n820 VDD.n819 0.04025
R6343 VDD.n819 VDD.n600 0.04025
R6344 VDD.n815 VDD.n600 0.04025
R6345 VDD.n815 VDD.n814 0.04025
R6346 VDD.n814 VDD.n813 0.04025
R6347 VDD.n813 VDD.n602 0.04025
R6348 VDD.n809 VDD.n602 0.04025
R6349 VDD.n809 VDD.n808 0.04025
R6350 VDD.n808 VDD.n807 0.04025
R6351 VDD.n807 VDD.n604 0.04025
R6352 VDD.n803 VDD.n604 0.04025
R6353 VDD.n803 VDD.n802 0.04025
R6354 VDD.n802 VDD.n801 0.04025
R6355 VDD.n801 VDD.n606 0.04025
R6356 VDD.n797 VDD.n606 0.04025
R6357 VDD.n797 VDD.n796 0.04025
R6358 VDD.n796 VDD.n795 0.04025
R6359 VDD.n795 VDD.n608 0.04025
R6360 VDD.n791 VDD.n608 0.04025
R6361 VDD.n791 VDD.n790 0.04025
R6362 VDD.n790 VDD.n789 0.04025
R6363 VDD.n789 VDD.n610 0.04025
R6364 VDD.n785 VDD.n610 0.04025
R6365 VDD.n785 VDD.n784 0.04025
R6366 VDD.n784 VDD.n783 0.04025
R6367 VDD.n783 VDD.n612 0.04025
R6368 VDD.n779 VDD.n612 0.04025
R6369 VDD.n779 VDD.n778 0.04025
R6370 VDD.n778 VDD.n777 0.04025
R6371 VDD.n777 VDD.n614 0.04025
R6372 VDD.n773 VDD.n614 0.04025
R6373 VDD.n773 VDD.n772 0.04025
R6374 VDD.n772 VDD.n771 0.04025
R6375 VDD.n771 VDD.n616 0.04025
R6376 VDD.n767 VDD.n616 0.04025
R6377 VDD.n767 VDD.n766 0.04025
R6378 VDD.n766 VDD.n765 0.04025
R6379 VDD.n765 VDD.n618 0.04025
R6380 VDD.n761 VDD.n618 0.04025
R6381 VDD.n761 VDD.n760 0.04025
R6382 VDD.n760 VDD.n759 0.04025
R6383 VDD.n759 VDD.n620 0.04025
R6384 VDD.n755 VDD.n620 0.04025
R6385 VDD.n755 VDD.n754 0.04025
R6386 VDD.n754 VDD.n753 0.04025
R6387 VDD.n753 VDD.n622 0.04025
R6388 VDD.n749 VDD.n622 0.04025
R6389 VDD.n749 VDD.n748 0.04025
R6390 VDD.n748 VDD.n747 0.04025
R6391 VDD.n747 VDD.n624 0.04025
R6392 VDD.n743 VDD.n624 0.04025
R6393 VDD.n743 VDD.n742 0.04025
R6394 VDD.n742 VDD.n741 0.04025
R6395 VDD.n741 VDD.n626 0.04025
R6396 VDD.n737 VDD.n626 0.04025
R6397 VDD.n737 VDD.n736 0.04025
R6398 VDD.n736 VDD.n735 0.04025
R6399 VDD.n735 VDD.n628 0.04025
R6400 VDD.n731 VDD.n628 0.04025
R6401 VDD.n731 VDD.n730 0.04025
R6402 VDD.n730 VDD.n729 0.04025
R6403 VDD.n729 VDD.n630 0.04025
R6404 VDD.n725 VDD.n630 0.04025
R6405 VDD.n725 VDD.n724 0.04025
R6406 VDD.n724 VDD.n723 0.04025
R6407 VDD.n723 VDD.n632 0.04025
R6408 VDD.n719 VDD.n632 0.04025
R6409 VDD.n719 VDD.n718 0.04025
R6410 VDD.n718 VDD.n717 0.04025
R6411 VDD.n717 VDD.n634 0.04025
R6412 VDD.n713 VDD.n634 0.04025
R6413 VDD.n713 VDD.n712 0.04025
R6414 VDD.n712 VDD.n711 0.04025
R6415 VDD.n711 VDD.n636 0.04025
R6416 VDD.n707 VDD.n636 0.04025
R6417 VDD.n707 VDD.n706 0.04025
R6418 VDD.n706 VDD.n705 0.04025
R6419 VDD.n705 VDD.n638 0.04025
R6420 VDD.n639 VDD.n638 0.04025
R6421 VDD.n870 VDD.n583 0.04025
R6422 VDD.n866 VDD.n583 0.04025
R6423 VDD.n866 VDD.n865 0.04025
R6424 VDD.n865 VDD.n864 0.04025
R6425 VDD.n864 VDD.n585 0.04025
R6426 VDD.n860 VDD.n585 0.04025
R6427 VDD.n860 VDD.n859 0.04025
R6428 VDD.n859 VDD.n858 0.04025
R6429 VDD.n858 VDD.n587 0.04025
R6430 VDD.n854 VDD.n587 0.04025
R6431 VDD.n854 VDD.n853 0.04025
R6432 VDD.n853 VDD.n852 0.04025
R6433 VDD.n852 VDD.n589 0.04025
R6434 VDD.n848 VDD.n589 0.04025
R6435 VDD.n848 VDD.n847 0.04025
R6436 VDD.n847 VDD.n846 0.04025
R6437 VDD.n846 VDD.n591 0.04025
R6438 VDD.n842 VDD.n591 0.04025
R6439 VDD.n842 VDD.n841 0.04025
R6440 VDD.n841 VDD.n840 0.04025
R6441 VDD.n840 VDD.n593 0.04025
R6442 VDD.n836 VDD.n593 0.04025
R6443 VDD.n836 VDD.n835 0.04025
R6444 VDD.n835 VDD.n834 0.04025
R6445 VDD.n834 VDD.n595 0.04025
R6446 VDD.n830 VDD.n595 0.04025
R6447 VDD.n830 VDD.n829 0.04025
R6448 VDD.n829 VDD.n828 0.04025
R6449 VDD.n828 VDD.n597 0.04025
R6450 VDD.n824 VDD.n597 0.04025
R6451 VDD.n824 VDD.n823 0.04025
R6452 VDD.n823 VDD.n822 0.04025
R6453 VDD.n822 VDD.n599 0.04025
R6454 VDD.n818 VDD.n599 0.04025
R6455 VDD.n818 VDD.n817 0.04025
R6456 VDD.n817 VDD.n816 0.04025
R6457 VDD.n816 VDD.n601 0.04025
R6458 VDD.n812 VDD.n601 0.04025
R6459 VDD.n812 VDD.n811 0.04025
R6460 VDD.n811 VDD.n810 0.04025
R6461 VDD.n810 VDD.n603 0.04025
R6462 VDD.n806 VDD.n603 0.04025
R6463 VDD.n806 VDD.n805 0.04025
R6464 VDD.n805 VDD.n804 0.04025
R6465 VDD.n804 VDD.n605 0.04025
R6466 VDD.n800 VDD.n605 0.04025
R6467 VDD.n800 VDD.n799 0.04025
R6468 VDD.n799 VDD.n798 0.04025
R6469 VDD.n798 VDD.n607 0.04025
R6470 VDD.n794 VDD.n607 0.04025
R6471 VDD.n794 VDD.n793 0.04025
R6472 VDD.n793 VDD.n792 0.04025
R6473 VDD.n792 VDD.n609 0.04025
R6474 VDD.n788 VDD.n609 0.04025
R6475 VDD.n788 VDD.n787 0.04025
R6476 VDD.n787 VDD.n786 0.04025
R6477 VDD.n786 VDD.n611 0.04025
R6478 VDD.n782 VDD.n611 0.04025
R6479 VDD.n782 VDD.n781 0.04025
R6480 VDD.n781 VDD.n780 0.04025
R6481 VDD.n780 VDD.n613 0.04025
R6482 VDD.n776 VDD.n613 0.04025
R6483 VDD.n776 VDD.n775 0.04025
R6484 VDD.n775 VDD.n774 0.04025
R6485 VDD.n774 VDD.n615 0.04025
R6486 VDD.n770 VDD.n615 0.04025
R6487 VDD.n770 VDD.n769 0.04025
R6488 VDD.n769 VDD.n768 0.04025
R6489 VDD.n768 VDD.n617 0.04025
R6490 VDD.n764 VDD.n617 0.04025
R6491 VDD.n764 VDD.n763 0.04025
R6492 VDD.n763 VDD.n762 0.04025
R6493 VDD.n762 VDD.n619 0.04025
R6494 VDD.n758 VDD.n619 0.04025
R6495 VDD.n758 VDD.n757 0.04025
R6496 VDD.n757 VDD.n756 0.04025
R6497 VDD.n756 VDD.n621 0.04025
R6498 VDD.n752 VDD.n621 0.04025
R6499 VDD.n752 VDD.n751 0.04025
R6500 VDD.n751 VDD.n750 0.04025
R6501 VDD.n750 VDD.n623 0.04025
R6502 VDD.n746 VDD.n623 0.04025
R6503 VDD.n746 VDD.n745 0.04025
R6504 VDD.n745 VDD.n744 0.04025
R6505 VDD.n744 VDD.n625 0.04025
R6506 VDD.n740 VDD.n625 0.04025
R6507 VDD.n740 VDD.n739 0.04025
R6508 VDD.n739 VDD.n738 0.04025
R6509 VDD.n738 VDD.n627 0.04025
R6510 VDD.n734 VDD.n627 0.04025
R6511 VDD.n734 VDD.n733 0.04025
R6512 VDD.n733 VDD.n732 0.04025
R6513 VDD.n732 VDD.n629 0.04025
R6514 VDD.n728 VDD.n629 0.04025
R6515 VDD.n728 VDD.n727 0.04025
R6516 VDD.n727 VDD.n726 0.04025
R6517 VDD.n726 VDD.n631 0.04025
R6518 VDD.n722 VDD.n631 0.04025
R6519 VDD.n722 VDD.n721 0.04025
R6520 VDD.n721 VDD.n720 0.04025
R6521 VDD.n720 VDD.n633 0.04025
R6522 VDD.n716 VDD.n633 0.04025
R6523 VDD.n716 VDD.n715 0.04025
R6524 VDD.n715 VDD.n714 0.04025
R6525 VDD.n714 VDD.n635 0.04025
R6526 VDD.n710 VDD.n635 0.04025
R6527 VDD.n710 VDD.n709 0.04025
R6528 VDD.n709 VDD.n708 0.04025
R6529 VDD.n708 VDD.n637 0.04025
R6530 VDD.n704 VDD.n637 0.04025
R6531 VDD.n704 VDD.n703 0.04025
R6532 VDD.n703 VDD.n702 0.04025
R6533 VDD.n701 VDD.n640 0.04025
R6534 VDD.n697 VDD.n640 0.04025
R6535 VDD.n697 VDD.n696 0.04025
R6536 VDD.n696 VDD.n695 0.04025
R6537 VDD.n695 VDD.n642 0.04025
R6538 VDD.n691 VDD.n642 0.04025
R6539 VDD.n691 VDD.n690 0.04025
R6540 VDD.n690 VDD.n689 0.04025
R6541 VDD.n689 VDD.n644 0.04025
R6542 VDD.n685 VDD.n644 0.04025
R6543 VDD.n685 VDD.n684 0.04025
R6544 VDD.n684 VDD.n683 0.04025
R6545 VDD.n683 VDD.n646 0.04025
R6546 VDD.n679 VDD.n646 0.04025
R6547 VDD.n679 VDD.n678 0.04025
R6548 VDD.n678 VDD.n677 0.04025
R6549 VDD.n677 VDD.n648 0.04025
R6550 VDD.n673 VDD.n648 0.04025
R6551 VDD.n673 VDD.n672 0.04025
R6552 VDD.n672 VDD.n671 0.04025
R6553 VDD.n671 VDD.n650 0.04025
R6554 VDD.n667 VDD.n650 0.04025
R6555 VDD.n667 VDD.n666 0.04025
R6556 VDD.n666 VDD.n665 0.04025
R6557 VDD.n665 VDD.n652 0.04025
R6558 VDD.n661 VDD.n652 0.04025
R6559 VDD.n661 VDD.n660 0.04025
R6560 VDD.n660 VDD.n659 0.04025
R6561 VDD.n659 VDD.n654 0.04025
R6562 VDD.n655 VDD.n654 0.04025
R6563 VDD.n655 VDD.n581 0.04025
R6564 VDD.n873 VDD.n581 0.04025
R6565 VDD.n877 VDD.n579 0.04025
R6566 VDD.n878 VDD.n877 0.04025
R6567 VDD.n879 VDD.n878 0.04025
R6568 VDD.n879 VDD.n574 0.04025
R6569 VDD.n144 VDD.n143 0.0373782
R6570 VDD.n178 VDD.n177 0.0373782
R6571 VDD.n176 VDD.n175 0.0373782
R6572 VDD.n174 VDD.n173 0.0373782
R6573 VDD.n172 VDD.n171 0.0373782
R6574 VDD.n238 VDD.n237 0.0373782
R6575 VDD.n269 VDD.n268 0.0373782
R6576 VDD.n267 VDD.n266 0.0373782
R6577 VDD.n265 VDD.n264 0.0373782
R6578 VDD.n263 VDD.n262 0.0373782
R6579 VDD.n545 VDD.n12 0.0358571
R6580 VDD.n490 VDD.n473 0.0358571
R6581 VDD.n211 VDD.n210 0.0323214
R6582 VDD.n137 VDD.n136 0.0323214
R6583 VDD.n139 VDD.n138 0.0323214
R6584 VDD.n153 VDD.n152 0.0323214
R6585 VDD.n150 VDD.n149 0.0323214
R6586 VDD.n301 VDD.n300 0.0323214
R6587 VDD.n232 VDD.n231 0.0323214
R6588 VDD.n229 VDD.n228 0.0323214
R6589 VDD.n243 VDD.n242 0.0323214
R6590 VDD.n245 VDD.n244 0.0323214
R6591 VDD.n258 VDD.n257 0.0323214
R6592 VDD.n255 VDD.n254 0.0323214
R6593 VDD.n166 VDD.n165 0.0323214
R6594 VDD.n168 VDD.n167 0.0323214
R6595 VDD.n1178 VDD.n953 0.0320556
R6596 VDD.n1179 VDD.n953 0.0320556
R6597 VDD.n1180 VDD.n1179 0.0320556
R6598 VDD.n1180 VDD.n952 0.0320556
R6599 VDD.n1181 VDD.n952 0.0320556
R6600 VDD.n1182 VDD.n1181 0.0320556
R6601 VDD.n1182 VDD.n951 0.0320556
R6602 VDD.n1183 VDD.n951 0.0320556
R6603 VDD.n1184 VDD.n1183 0.0320556
R6604 VDD.n1184 VDD.n950 0.0320556
R6605 VDD.n1185 VDD.n950 0.0320556
R6606 VDD.n1186 VDD.n1185 0.0320556
R6607 VDD.n1186 VDD.n949 0.0320556
R6608 VDD.n1187 VDD.n949 0.0320556
R6609 VDD.n1188 VDD.n1187 0.0320556
R6610 VDD.n1188 VDD.n948 0.0320556
R6611 VDD.n1189 VDD.n948 0.0320556
R6612 VDD.n1190 VDD.n1189 0.0320556
R6613 VDD.n1190 VDD.n947 0.0320556
R6614 VDD.n1191 VDD.n947 0.0320556
R6615 VDD.n1208 VDD.n1195 0.0320556
R6616 VDD.n1207 VDD.n1195 0.0320556
R6617 VDD.n1207 VDD.n1206 0.0320556
R6618 VDD.n1206 VDD.n1196 0.0320556
R6619 VDD.n1205 VDD.n1196 0.0320556
R6620 VDD.n884 VDD.n574 0.032
R6621 VDD.n1199 VDD.n942 0.0319052
R6622 VDD.n1200 VDD.n1199 0.0319052
R6623 VDD.n1201 VDD.n1198 0.0319052
R6624 VDD.n1202 VDD.n1198 0.0319052
R6625 VDD.n1203 VDD.n1197 0.0319052
R6626 VDD.n1214 VDD.n1192 0.0319052
R6627 VDD.n1213 VDD.n1192 0.0319052
R6628 VDD.n1212 VDD.n1193 0.0319052
R6629 VDD.n1211 VDD.n1193 0.0319052
R6630 VDD.n1210 VDD.n1194 0.0319052
R6631 VDD.n1229 VDD.n939 0.0319052
R6632 VDD.n1228 VDD.n940 0.0319052
R6633 VDD.n1227 VDD.n940 0.0319052
R6634 VDD.n1226 VDD.n941 0.0319052
R6635 VDD.n1225 VDD.n941 0.0319052
R6636 VDD.n1171 VDD.n957 0.0317952
R6637 VDD.n1172 VDD.n956 0.0317952
R6638 VDD.n1173 VDD.n956 0.0317952
R6639 VDD.n1174 VDD.n955 0.0317952
R6640 VDD.n1175 VDD.n955 0.0317952
R6641 VDD.n1176 VDD.n954 0.0317952
R6642 VDD.n1201 VDD.n1200 0.0304297
R6643 VDD.n1203 VDD.n1202 0.0304297
R6644 VDD.n1213 VDD.n1212 0.0304297
R6645 VDD.n1211 VDD.n1210 0.0304297
R6646 VDD.n1229 VDD.n1228 0.0304297
R6647 VDD.n1227 VDD.n1226 0.0304297
R6648 VDD.n1172 VDD.n1171 0.030325
R6649 VDD.n1174 VDD.n1173 0.030325
R6650 VDD.n1176 VDD.n1175 0.030325
R6651 VDD.n1209 VDD.n1208 0.0278333
R6652 VDD.n1205 VDD.n1204 0.0278333
R6653 VDD.n1178 VDD.n1177 0.0275
R6654 VDD.n1225 VDD.n1224 0.0260035
R6655 VDD.n1224 VDD.n942 0.0258981
R6656 VDD.n1215 VDD.n1214 0.0258981
R6657 VDD.n513 VDD.n22 0.0251429
R6658 VDD.n1230 VDD.n938 0.025055
R6659 VDD.n1168 VDD.n959 0.02435
R6660 VDD.n1164 VDD.n959 0.02435
R6661 VDD.n1164 VDD.n1163 0.02435
R6662 VDD.n1163 VDD.n961 0.02435
R6663 VDD.n1158 VDD.n1157 0.02435
R6664 VDD.n1157 VDD.n1156 0.02435
R6665 VDD.n1156 VDD.n965 0.02435
R6666 VDD.n972 VDD.n965 0.02435
R6667 VDD.n973 VDD.n972 0.02435
R6668 VDD.n973 VDD.n970 0.02435
R6669 VDD.n978 VDD.n970 0.02435
R6670 VDD.n979 VDD.n978 0.02435
R6671 VDD.n1151 VDD.n1150 0.02435
R6672 VDD.n1150 VDD.n1149 0.02435
R6673 VDD.n1149 VDD.n981 0.02435
R6674 VDD.n1145 VDD.n981 0.02435
R6675 VDD.n1145 VDD.n1144 0.02435
R6676 VDD.n1144 VDD.n984 0.02435
R6677 VDD.n1140 VDD.n984 0.02435
R6678 VDD.n1138 VDD.n987 0.02435
R6679 VDD.n994 VDD.n987 0.02435
R6680 VDD.n995 VDD.n994 0.02435
R6681 VDD.n996 VDD.n995 0.02435
R6682 VDD.n996 VDD.n992 0.02435
R6683 VDD.n1001 VDD.n992 0.02435
R6684 VDD.n1002 VDD.n1001 0.02435
R6685 VDD.n1132 VDD.n1131 0.02435
R6686 VDD.n1131 VDD.n1130 0.02435
R6687 VDD.n1130 VDD.n1004 0.02435
R6688 VDD.n1126 VDD.n1004 0.02435
R6689 VDD.n1126 VDD.n1125 0.02435
R6690 VDD.n1125 VDD.n1007 0.02435
R6691 VDD.n1121 VDD.n1007 0.02435
R6692 VDD.n1119 VDD.n1010 0.02435
R6693 VDD.n1018 VDD.n1010 0.02435
R6694 VDD.n1019 VDD.n1018 0.02435
R6695 VDD.n1020 VDD.n1019 0.02435
R6696 VDD.n1020 VDD.n1016 0.02435
R6697 VDD.n1025 VDD.n1016 0.02435
R6698 VDD.n1026 VDD.n1025 0.02435
R6699 VDD.n1113 VDD.n1112 0.02435
R6700 VDD.n1112 VDD.n1111 0.02435
R6701 VDD.n1111 VDD.n1028 0.02435
R6702 VDD.n1107 VDD.n1028 0.02435
R6703 VDD.n1107 VDD.n1106 0.02435
R6704 VDD.n1106 VDD.n1031 0.02435
R6705 VDD.n1102 VDD.n1031 0.02435
R6706 VDD.n1100 VDD.n1034 0.02435
R6707 VDD.n1041 VDD.n1034 0.02435
R6708 VDD.n1042 VDD.n1041 0.02435
R6709 VDD.n1043 VDD.n1042 0.02435
R6710 VDD.n1043 VDD.n1039 0.02435
R6711 VDD.n1048 VDD.n1039 0.02435
R6712 VDD.n1049 VDD.n1048 0.02435
R6713 VDD.n1094 VDD.n1093 0.02435
R6714 VDD.n1093 VDD.n1092 0.02435
R6715 VDD.n1092 VDD.n1051 0.02435
R6716 VDD.n1088 VDD.n1051 0.02435
R6717 VDD.n1088 VDD.n1087 0.02435
R6718 VDD.n1087 VDD.n1054 0.02435
R6719 VDD.n1083 VDD.n1054 0.02435
R6720 VDD.n1081 VDD.n1057 0.02435
R6721 VDD.n1064 VDD.n1057 0.02435
R6722 VDD.n1065 VDD.n1064 0.02435
R6723 VDD.n1066 VDD.n1065 0.02435
R6724 VDD.n1066 VDD.n1062 0.02435
R6725 VDD.n1071 VDD.n1062 0.02435
R6726 VDD.n1072 VDD.n1071 0.02435
R6727 VDD.n1075 VDD.n1074 0.02435
R6728 VDD.n935 VDD.n558 0.02435
R6729 VDD.n931 VDD.n558 0.02435
R6730 VDD.n931 VDD.n930 0.02435
R6731 VDD.n930 VDD.n929 0.02435
R6732 VDD.n929 VDD.n561 0.02435
R6733 VDD.n925 VDD.n561 0.02435
R6734 VDD.n923 VDD.n922 0.02435
R6735 VDD.n913 VDD.n564 0.02435
R6736 VDD.n909 VDD.n564 0.02435
R6737 VDD.n909 VDD.n908 0.02435
R6738 VDD.n908 VDD.n907 0.02435
R6739 VDD.n907 VDD.n567 0.02435
R6740 VDD.n903 VDD.n567 0.02435
R6741 VDD.n903 VDD.n902 0.02435
R6742 VDD.n902 VDD.n901 0.02435
R6743 VDD.n901 VDD.n570 0.02435
R6744 VDD.n897 VDD.n570 0.02435
R6745 VDD.n895 VDD.n894 0.02435
R6746 VDD.n964 VDD.n961 0.024125
R6747 VDD.n141 VDD.n140 0.023624
R6748 VDD.n147 VDD.n146 0.023624
R6749 VDD.n170 VDD.n169 0.023624
R6750 VDD.n235 VDD.n234 0.023624
R6751 VDD.n241 VDD.n240 0.023624
R6752 VDD.n261 VDD.n260 0.023624
R6753 VDD.n213 VDD.n212 0.0235265
R6754 VDD.n212 VDD.n211 0.0235265
R6755 VDD.n210 VDD.n209 0.0235265
R6756 VDD.n209 VDD.n208 0.0235265
R6757 VDD.n135 VDD.n125 0.0235265
R6758 VDD.n136 VDD.n135 0.0235265
R6759 VDD.n137 VDD.n134 0.0235265
R6760 VDD.n138 VDD.n134 0.0235265
R6761 VDD.n139 VDD.n133 0.0235265
R6762 VDD.n155 VDD.n154 0.0235265
R6763 VDD.n154 VDD.n153 0.0235265
R6764 VDD.n152 VDD.n151 0.0235265
R6765 VDD.n151 VDD.n150 0.0235265
R6766 VDD.n149 VDD.n148 0.0235265
R6767 VDD.n299 VDD.n215 0.0235265
R6768 VDD.n300 VDD.n215 0.0235265
R6769 VDD.n301 VDD.n214 0.0235265
R6770 VDD.n302 VDD.n214 0.0235265
R6771 VDD.n233 VDD.n232 0.0235265
R6772 VDD.n231 VDD.n230 0.0235265
R6773 VDD.n230 VDD.n229 0.0235265
R6774 VDD.n228 VDD.n227 0.0235265
R6775 VDD.n227 VDD.n216 0.0235265
R6776 VDD.n242 VDD.n226 0.0235265
R6777 VDD.n243 VDD.n225 0.0235265
R6778 VDD.n244 VDD.n225 0.0235265
R6779 VDD.n245 VDD.n224 0.0235265
R6780 VDD.n246 VDD.n224 0.0235265
R6781 VDD.n259 VDD.n258 0.0235265
R6782 VDD.n257 VDD.n256 0.0235265
R6783 VDD.n256 VDD.n255 0.0235265
R6784 VDD.n254 VDD.n253 0.0235265
R6785 VDD.n253 VDD.n252 0.0235265
R6786 VDD.n164 VDD.n163 0.0235265
R6787 VDD.n165 VDD.n163 0.0235265
R6788 VDD.n166 VDD.n162 0.0235265
R6789 VDD.n167 VDD.n162 0.0235265
R6790 VDD.n168 VDD.n161 0.0235265
R6791 VDD.n1151 VDD.n980 0.02345
R6792 VDD.n1139 VDD.n1138 0.022775
R6793 VDD.n142 VDD.n141 0.0227498
R6794 VDD.n143 VDD.n142 0.0227498
R6795 VDD.n145 VDD.n144 0.0227498
R6796 VDD.n146 VDD.n145 0.0227498
R6797 VDD.n179 VDD.n178 0.0227498
R6798 VDD.n177 VDD.n157 0.0227498
R6799 VDD.n176 VDD.n157 0.0227498
R6800 VDD.n175 VDD.n158 0.0227498
R6801 VDD.n174 VDD.n158 0.0227498
R6802 VDD.n173 VDD.n159 0.0227498
R6803 VDD.n172 VDD.n159 0.0227498
R6804 VDD.n171 VDD.n160 0.0227498
R6805 VDD.n170 VDD.n160 0.0227498
R6806 VDD.n236 VDD.n235 0.0227498
R6807 VDD.n237 VDD.n236 0.0227498
R6808 VDD.n239 VDD.n238 0.0227498
R6809 VDD.n240 VDD.n239 0.0227498
R6810 VDD.n270 VDD.n269 0.0227498
R6811 VDD.n268 VDD.n248 0.0227498
R6812 VDD.n267 VDD.n248 0.0227498
R6813 VDD.n266 VDD.n249 0.0227498
R6814 VDD.n265 VDD.n249 0.0227498
R6815 VDD.n264 VDD.n250 0.0227498
R6816 VDD.n263 VDD.n250 0.0227498
R6817 VDD.n262 VDD.n251 0.0227498
R6818 VDD.n261 VDD.n251 0.0227498
R6819 VDD.n1132 VDD.n1003 0.021875
R6820 VDD.n180 VDD.n179 0.0209847
R6821 VDD.n271 VDD.n270 0.0209847
R6822 VDD.n1120 VDD.n1119 0.020975
R6823 VDD.n576 VDD.n573 0.0207876
R6824 VDD.n882 VDD.n572 0.0207876
R6825 VDD.n871 VDD.n870 0.020375
R6826 VDD.n873 VDD.n872 0.020375
R6827 VDD.n872 VDD.n579 0.020375
R6828 VDD.n1113 VDD.n1027 0.020075
R6829 VDD.n303 VDD.n213 0.0198811
R6830 VDD.n208 VDD.n207 0.0198811
R6831 VDD.n207 VDD.n125 0.0198811
R6832 VDD.n184 VDD.n155 0.0198811
R6833 VDD.n299 VDD.n298 0.0198811
R6834 VDD.n303 VDD.n302 0.0198811
R6835 VDD.n298 VDD.n216 0.0198811
R6836 VDD.n275 VDD.n246 0.0198811
R6837 VDD.n252 VDD.n52 0.0198811
R6838 VDD.n164 VDD.n52 0.0198811
R6839 VDD.n1101 VDD.n1100 0.019175
R6840 VDD.n1216 VDD.n1191 0.0190218
R6841 VDD.n1094 VDD.n1050 0.018275
R6842 VDD.n1082 VDD.n1081 0.017375
R6843 VDD.n1217 VDD.n946 0.0171298
R6844 VDD.n1218 VDD.n1217 0.0171298
R6845 VDD.n1218 VDD.n945 0.0171298
R6846 VDD.n1219 VDD.n945 0.0171298
R6847 VDD.n1220 VDD.n1219 0.0171298
R6848 VDD.n1220 VDD.n944 0.0171298
R6849 VDD.n1221 VDD.n944 0.0171298
R6850 VDD.n1222 VDD.n1221 0.0171298
R6851 VDD.n1222 VDD.n943 0.0171298
R6852 VDD.n925 VDD.n924 0.0167
R6853 VDD.n1075 VDD.n1073 0.016475
R6854 VDD.n181 VDD.n180 0.0157263
R6855 VDD.n272 VDD.n271 0.0157263
R6856 VDD.n1170 VDD.n1169 0.0146745
R6857 VDD.n1169 VDD.n958 0.0143101
R6858 VDD.n897 VDD.n896 0.014
R6859 VDD VDD.n1230 0.0135679
R6860 VDD.n885 VDD.n884 0.012425
R6861 VDD.n884 VDD.n883 0.012425
R6862 VDD.n1167 VDD.n1166 0.0122778
R6863 VDD.n1166 VDD.n1165 0.0122778
R6864 VDD.n1162 VDD.n1161 0.0122778
R6865 VDD.n1159 VDD.n962 0.0122778
R6866 VDD.n1155 VDD.n962 0.0122778
R6867 VDD.n971 VDD.n966 0.0122778
R6868 VDD.n974 VDD.n971 0.0122778
R6869 VDD.n977 VDD.n976 0.0122778
R6870 VDD.n977 VDD.n967 0.0122778
R6871 VDD.n1152 VDD.n968 0.0122778
R6872 VDD.n1148 VDD.n1147 0.0122778
R6873 VDD.n1147 VDD.n1146 0.0122778
R6874 VDD.n1143 VDD.n1142 0.0122778
R6875 VDD.n1142 VDD.n1141 0.0122778
R6876 VDD.n1137 VDD.n1136 0.0122778
R6877 VDD.n993 VDD.n988 0.0122778
R6878 VDD.n997 VDD.n993 0.0122778
R6879 VDD.n1000 VDD.n999 0.0122778
R6880 VDD.n1000 VDD.n989 0.0122778
R6881 VDD.n1133 VDD.n990 0.0122778
R6882 VDD.n1129 VDD.n1128 0.0122778
R6883 VDD.n1128 VDD.n1127 0.0122778
R6884 VDD.n1124 VDD.n1123 0.0122778
R6885 VDD.n1123 VDD.n1122 0.0122778
R6886 VDD.n1118 VDD.n1117 0.0122778
R6887 VDD.n1017 VDD.n1011 0.0122778
R6888 VDD.n1021 VDD.n1017 0.0122778
R6889 VDD.n1024 VDD.n1023 0.0122778
R6890 VDD.n1024 VDD.n1012 0.0122778
R6891 VDD.n1114 VDD.n1013 0.0122778
R6892 VDD.n1110 VDD.n1109 0.0122778
R6893 VDD.n1109 VDD.n1108 0.0122778
R6894 VDD.n1105 VDD.n1104 0.0122778
R6895 VDD.n1104 VDD.n1103 0.0122778
R6896 VDD.n1099 VDD.n1098 0.0122778
R6897 VDD.n1040 VDD.n1035 0.0122778
R6898 VDD.n1044 VDD.n1040 0.0122778
R6899 VDD.n1047 VDD.n1046 0.0122778
R6900 VDD.n1047 VDD.n1036 0.0122778
R6901 VDD.n1095 VDD.n1037 0.0122778
R6902 VDD.n1091 VDD.n1090 0.0122778
R6903 VDD.n1090 VDD.n1089 0.0122778
R6904 VDD.n1086 VDD.n1085 0.0122778
R6905 VDD.n1085 VDD.n1084 0.0122778
R6906 VDD.n1080 VDD.n1079 0.0122778
R6907 VDD.n1063 VDD.n1058 0.0122778
R6908 VDD.n1067 VDD.n1063 0.0122778
R6909 VDD.n1070 VDD.n1069 0.0122778
R6910 VDD.n1070 VDD.n1059 0.0122778
R6911 VDD.n1076 VDD.n1060 0.0122778
R6912 VDD.n1161 VDD.n1160 0.0121667
R6913 VDD.n1153 VDD.n1152 0.0119444
R6914 VDD.n1079 VDD.n1078 0.0119444
R6915 VDD.n1137 VDD.n985 0.0115
R6916 VDD.n1052 VDD.n1037 0.0115
R6917 VDD.n1134 VDD.n1133 0.0110556
R6918 VDD.n1098 VDD.n1097 0.0110556
R6919 VDD.n1216 VDD.n1215 0.0109815
R6920 VDD.n1224 VDD.n1223 0.0109815
R6921 VDD.n896 VDD.n895 0.01085
R6922 VDD.n1118 VDD.n1008 0.0106111
R6923 VDD.n1029 VDD.n1013 0.0106111
R6924 VDD.n203 VDD.n202 0.0104419
R6925 VDD.n196 VDD.n195 0.0104419
R6926 VDD.n189 VDD.n188 0.0104419
R6927 VDD.n294 VDD.n293 0.0104419
R6928 VDD.n287 VDD.n286 0.0104419
R6929 VDD.n280 VDD.n279 0.0104419
R6930 VDD.n1117 VDD.n1116 0.0101667
R6931 VDD.n1115 VDD.n1114 0.0101667
R6932 VDD.n206 VDD.n205 0.0099186
R6933 VDD.n200 VDD.n199 0.0099186
R6934 VDD.n199 VDD.n198 0.0099186
R6935 VDD.n193 VDD.n192 0.0099186
R6936 VDD.n192 VDD.n191 0.0099186
R6937 VDD.n186 VDD.n185 0.0099186
R6938 VDD.n297 VDD.n296 0.0099186
R6939 VDD.n291 VDD.n290 0.0099186
R6940 VDD.n290 VDD.n289 0.0099186
R6941 VDD.n284 VDD.n283 0.0099186
R6942 VDD.n283 VDD.n282 0.0099186
R6943 VDD.n277 VDD.n276 0.0099186
R6944 VDD.n1005 VDD.n990 0.00972222
R6945 VDD.n1099 VDD.n1032 0.00972222
R6946 VDD.n1136 VDD.n1135 0.00927778
R6947 VDD.n1096 VDD.n1095 0.00927778
R6948 VDD.n982 VDD.n968 0.00883333
R6949 VDD.n1080 VDD.n1055 0.00883333
R6950 VDD.n1162 VDD.n960 0.00861111
R6951 VDD.n1155 VDD.n1154 0.00838889
R6952 VDD.n1077 VDD.n1076 0.00838889
R6953 VDD.n1073 VDD.n1072 0.008375
R6954 VDD.n140 VDD.n133 0.00825064
R6955 VDD.n148 VDD.n147 0.00825064
R6956 VDD.n234 VDD.n233 0.00825064
R6957 VDD.n241 VDD.n226 0.00825064
R6958 VDD.n260 VDD.n259 0.00825064
R6959 VDD.n169 VDD.n161 0.00825064
R6960 VDD.n976 VDD.n975 0.00816667
R6961 VDD.n1068 VDD.n1067 0.00816667
R6962 VDD.n1060 VDD.n938 0.00816667
R6963 VDD.n924 VDD.n923 0.00815
R6964 VDD.n1143 VDD.n983 0.00772222
R6965 VDD.n1089 VDD.n1053 0.00772222
R6966 VDD.n1083 VDD.n1082 0.007475
R6967 VDD.n326 VDD.n325 0.00743314
R6968 VDD.n335 VDD.n334 0.00743314
R6969 VDD.n348 VDD.n102 0.00743314
R6970 VDD.n361 VDD.n360 0.00743314
R6971 VDD.n374 VDD.n86 0.00743314
R6972 VDD.n387 VDD.n386 0.00743314
R6973 VDD.n390 VDD.n73 0.00743314
R6974 VDD.n410 VDD.n67 0.00743314
R6975 VDD.n417 VDD.n58 0.00743314
R6976 VDD.n442 VDD.n48 0.00743314
R6977 VDD.n207 VDD.n206 0.00736773
R6978 VDD.n185 VDD.n184 0.00736773
R6979 VDD.n298 VDD.n297 0.00736773
R6980 VDD.n276 VDD.n275 0.00736773
R6981 VDD.n322 VDD.n321 0.00736773
R6982 VDD.n401 VDD.n71 0.00736773
R6983 VDD.n1204 VDD.n1197 0.00735012
R6984 VDD.n1209 VDD.n1194 0.00735012
R6985 VDD.n939 VDD.n938 0.00735012
R6986 VDD.n1170 VDD.n957 0.00732614
R6987 VDD.n1177 VDD.n954 0.00732614
R6988 VDD.n999 VDD.n998 0.00727778
R6989 VDD.n1045 VDD.n1044 0.00727778
R6990 VDD.n340 VDD.n339 0.00723692
R6991 VDD.n383 VDD.n382 0.00723692
R6992 VDD.n324 VDD.n116 0.0071061
R6993 VDD.n398 VDD.n397 0.0071061
R6994 VDD.n107 VDD.n106 0.00697529
R6995 VDD.n385 VDD.n80 0.00697529
R6996 VDD.n414 VDD.n413 0.00684448
R6997 VDD.n434 VDD.n433 0.00684448
R6998 VDD.n1124 VDD.n1006 0.00683333
R6999 VDD.n1108 VDD.n1030 0.00683333
R7000 VDD.n435 VDD.n52 0.00677907
R7001 VDD.n352 VDD.n351 0.00671366
R7002 VDD.n93 VDD.n88 0.00671366
R7003 VDD.n1215 VDD.n946 0.00664834
R7004 VDD.n1224 VDD.n943 0.00664834
R7005 VDD.n313 VDD.n123 0.00658285
R7006 VDD.n411 VDD.n65 0.00658285
R7007 VDD.n1050 VDD.n1049 0.006575
R7008 VDD.n349 VDD.n100 0.00645204
R7009 VDD.n370 VDD.n369 0.00645204
R7010 VDD.n1022 VDD.n1021 0.00638889
R7011 VDD.n1023 VDD.n1022 0.00638889
R7012 VDD.n420 VDD.n63 0.00632122
R7013 VDD.n429 VDD.n56 0.00632122
R7014 VDD.n357 VDD.n356 0.00619041
R7015 VDD.n366 VDD.n365 0.00619041
R7016 VDD.n425 VDD.n424 0.00605959
R7017 VDD.n1127 VDD.n1006 0.00594444
R7018 VDD.n1105 VDD.n1030 0.00594444
R7019 VDD.n359 VDD.n96 0.00592878
R7020 VDD.n91 VDD.n90 0.00592878
R7021 VDD.n308 VDD.n120 0.00579796
R7022 VDD.n406 VDD.n405 0.00579796
R7023 VDD.n442 VDD.n441 0.00579796
R7024 VDD.n309 VDD.n303 0.00573256
R7025 VDD.n1102 VDD.n1101 0.005675
R7026 VDD.n109 VDD.n104 0.00566715
R7027 VDD.n378 VDD.n377 0.00566715
R7028 VDD.n203 VDD.n127 0.00554783
R7029 VDD.n202 VDD.n128 0.00554783
R7030 VDD.n196 VDD.n129 0.00554783
R7031 VDD.n195 VDD.n130 0.00554783
R7032 VDD.n189 VDD.n131 0.00554783
R7033 VDD.n188 VDD.n132 0.00554783
R7034 VDD.n181 VDD.n156 0.00554783
R7035 VDD.n294 VDD.n218 0.00554783
R7036 VDD.n293 VDD.n219 0.00554783
R7037 VDD.n287 VDD.n220 0.00554783
R7038 VDD.n286 VDD.n221 0.00554783
R7039 VDD.n280 VDD.n222 0.00554783
R7040 VDD.n279 VDD.n223 0.00554783
R7041 VDD.n272 VDD.n247 0.00554783
R7042 VDD.n439 VDD.n50 0.00553634
R7043 VDD.n998 VDD.n997 0.0055
R7044 VDD.n1046 VDD.n1045 0.0055
R7045 VDD.n344 VDD.n343 0.00540552
R7046 VDD.n375 VDD.n84 0.00540552
R7047 VDD.n330 VDD.n114 0.00527471
R7048 VDD.n393 VDD.n78 0.00527471
R7049 VDD.n331 VDD.n330 0.0051439
R7050 VDD.n394 VDD.n393 0.0051439
R7051 VDD.n1146 VDD.n983 0.00505556
R7052 VDD.n1086 VDD.n1053 0.00505556
R7053 VDD.n333 VDD.n112 0.00488227
R7054 VDD.n76 VDD.n75 0.00488227
R7055 VDD.n1167 VDD.n958 0.00483333
R7056 VDD.n1027 VDD.n1026 0.004775
R7057 VDD.n110 VDD.n109 0.00475145
R7058 VDD.n378 VDD.n82 0.00475145
R7059 VDD.n316 VDD.n120 0.00462064
R7060 VDD.n406 VDD.n404 0.00462064
R7061 VDD.n430 VDD.n429 0.00462064
R7062 VDD.n975 VDD.n974 0.00461111
R7063 VDD.n1069 VDD.n1068 0.00461111
R7064 VDD.n1154 VDD.n966 0.00438889
R7065 VDD.n1077 VDD.n1059 0.00438889
R7066 VDD.n207 VDD.n126 0.00438406
R7067 VDD.n298 VDD.n217 0.00438406
R7068 VDD.n317 VDD.n118 0.00435901
R7069 VDD.n402 VDD.n69 0.00435901
R7070 VDD.n432 VDD.n54 0.00435901
R7071 VDD.n356 VDD.n98 0.0042282
R7072 VDD.n365 VDD.n94 0.0042282
R7073 VDD.n1165 VDD.n960 0.00416667
R7074 VDD.n414 VDD.n60 0.00409738
R7075 VDD.n421 VDD.n420 0.00409738
R7076 VDD.n1148 VDD.n982 0.00394444
R7077 VDD.n1084 VDD.n1055 0.00394444
R7078 VDD.n1121 VDD.n1120 0.003875
R7079 VDD.n61 VDD.n60 0.00383576
R7080 VDD.n421 VDD.n61 0.00383576
R7081 VDD.n352 VDD.n98 0.00370494
R7082 VDD.n94 VDD.n93 0.00370494
R7083 VDD.n321 VDD.n118 0.00357413
R7084 VDD.n402 VDD.n401 0.00357413
R7085 VDD.n433 VDD.n432 0.00357413
R7086 VDD.n1135 VDD.n988 0.0035
R7087 VDD.n1096 VDD.n1036 0.0035
R7088 VDD.n317 VDD.n316 0.0033125
R7089 VDD.n404 VDD.n69 0.0033125
R7090 VDD.n430 VDD.n54 0.0033125
R7091 VDD.n339 VDD.n110 0.00318169
R7092 VDD.n382 VDD.n82 0.00318169
R7093 VDD.n205 VDD.n127 0.00312096
R7094 VDD.n200 VDD.n128 0.00312096
R7095 VDD.n198 VDD.n129 0.00312096
R7096 VDD.n193 VDD.n130 0.00312096
R7097 VDD.n191 VDD.n131 0.00312096
R7098 VDD.n186 VDD.n132 0.00312096
R7099 VDD.n183 VDD.n156 0.00312096
R7100 VDD.n296 VDD.n218 0.00312096
R7101 VDD.n291 VDD.n219 0.00312096
R7102 VDD.n289 VDD.n220 0.00312096
R7103 VDD.n284 VDD.n221 0.00312096
R7104 VDD.n282 VDD.n222 0.00312096
R7105 VDD.n277 VDD.n223 0.00312096
R7106 VDD.n274 VDD.n247 0.00312096
R7107 VDD.n1129 VDD.n1005 0.00305556
R7108 VDD.n1103 VDD.n1032 0.00305556
R7109 VDD.n184 VDD.n183 0.00305087
R7110 VDD.n275 VDD.n274 0.00305087
R7111 VDD.n334 VDD.n333 0.00305087
R7112 VDD.n387 VDD.n75 0.00305087
R7113 VDD.n1003 VDD.n1002 0.002975
R7114 VDD.n331 VDD.n112 0.00278924
R7115 VDD.n394 VDD.n76 0.00278924
R7116 VDD.n326 VDD.n114 0.00265843
R7117 VDD.n390 VDD.n78 0.00265843
R7118 VDD.n1116 VDD.n1011 0.00261111
R7119 VDD.n1115 VDD.n1012 0.00261111
R7120 VDD.n343 VDD.n102 0.00252762
R7121 VDD.n375 VDD.n374 0.00252762
R7122 VDD.n439 VDD.n438 0.0023968
R7123 VDD.n344 VDD.n104 0.00226599
R7124 VDD.n377 VDD.n84 0.00226599
R7125 VDD.n312 VDD.n303 0.00220058
R7126 VDD.n1122 VDD.n1008 0.00216667
R7127 VDD.n1110 VDD.n1029 0.00216667
R7128 VDD.n309 VDD.n308 0.00213517
R7129 VDD.n405 VDD.n67 0.00213517
R7130 VDD.n441 VDD.n50 0.00213517
R7131 VDD.n1140 VDD.n1139 0.002075
R7132 VDD.n360 VDD.n359 0.00200436
R7133 VDD.n361 VDD.n90 0.00200436
R7134 VDD.n424 VDD.n58 0.00187355
R7135 VDD.n357 VDD.n96 0.00174273
R7136 VDD.n366 VDD.n91 0.00174273
R7137 VDD.n1134 VDD.n989 0.00172222
R7138 VDD.n1097 VDD.n1035 0.00172222
R7139 VDD.n417 VDD.n63 0.00161192
R7140 VDD.n425 VDD.n56 0.00161192
R7141 VDD.n349 VDD.n348 0.0014811
R7142 VDD.n369 VDD.n86 0.0014811
R7143 VDD.n980 VDD.n979 0.0014
R7144 VDD.n313 VDD.n312 0.00135029
R7145 VDD.n411 VDD.n410 0.00135029
R7146 VDD.n1141 VDD.n985 0.00127778
R7147 VDD.n1091 VDD.n1052 0.00127778
R7148 VDD.n351 VDD.n100 0.00121948
R7149 VDD.n370 VDD.n88 0.00121948
R7150 VDD.n438 VDD.n52 0.00115407
R7151 VDD.n123 VDD.n122 0.00108866
R7152 VDD.n413 VDD.n65 0.00108866
R7153 VDD.n435 VDD.n434 0.00108866
R7154 VDD.n335 VDD.n106 0.000957849
R7155 VDD.n386 VDD.n385 0.000957849
R7156 VDD.n1153 VDD.n967 0.000833333
R7157 VDD.n1078 VDD.n1058 0.000833333
R7158 VDD.n325 VDD.n324 0.000827035
R7159 VDD.n397 VDD.n73 0.000827035
R7160 VDD.n1158 VDD.n964 0.000725
R7161 VDD.n340 VDD.n107 0.000696221
R7162 VDD.n383 VDD.n80 0.000696221
R7163 VDD.n1160 VDD.n1159 0.000611111
R7164 VDD.n322 VDD.n116 0.000565407
R7165 VDD.n398 VDD.n71 0.000565407
R7166 a_11300_8092.n0 a_11300_8092.t0 7.34559
R7167 a_11300_8092.t9 a_11300_8092.t5 4.26279
R7168 a_11300_8092.t4 a_11300_8092.t5 3.86838
R7169 a_11300_8092.t5 a_11300_8092.t6 4.06156
R7170 a_11300_8092.t5 a_11300_8092.t8 4.06783
R7171 a_11300_8092.n0 a_11300_8092.t3 6.78329
R7172 a_11300_8092.n0 a_11300_8092.t2 6.78222
R7173 a_11300_8092.t5 a_11300_8092.n0 6.48046
R7174 a_11300_8092.n0 a_11300_8092.t1 6.17579
R7175 a_11300_8092.t7 a_11300_8092.t5 4.65501
R7176 a_16434_7468.n20 a_16434_7468.t0 11.8062
R7177 a_16434_7468.n14 a_16434_7468.t27 8.87887
R7178 a_16434_7468.t23 a_16434_7468.n15 4.06758
R7179 a_16434_7468.t27 a_16434_7468.n2 8.10567
R7180 a_16434_7468.t18 a_16434_7468.n0 3.82054
R7181 a_16434_7468.t28 a_16434_7468.n14 8.10567
R7182 a_16434_7468.n2 a_16434_7468.t28 8.10567
R7183 a_16434_7468.t20 a_16434_7468.n2 3.85103
R7184 a_16434_7468.n5 a_16434_7468.n13 0.478235
R7185 a_16434_7468.n5 a_16434_7468.t25 3.81497
R7186 a_16434_7468.n11 a_16434_7468.t8 3.85103
R7187 a_16434_7468.t31 a_16434_7468.n12 8.10567
R7188 a_16434_7468.n2 a_16434_7468.t31 8.10567
R7189 a_16434_7468.t4 a_16434_7468.n17 3.85103
R7190 a_16434_7468.t29 a_16434_7468.n10 8.10567
R7191 a_16434_7468.n2 a_16434_7468.t29 8.10567
R7192 a_16434_7468.t14 a_16434_7468.n18 3.91392
R7193 a_16434_7468.n19 a_16434_7468.t12 3.94737
R7194 a_16434_7468.n2 a_16434_7468.t22 8.10567
R7195 a_16434_7468.t22 a_16434_7468.n9 8.10567
R7196 a_16434_7468.t10 a_16434_7468.n2 3.85103
R7197 a_16434_7468.n3 a_16434_7468.t30 3.81497
R7198 a_16434_7468.n3 a_16434_7468.n8 0.478235
R7199 a_16434_7468.t16 a_16434_7468.n1 3.85103
R7200 a_16434_7468.n2 a_16434_7468.t24 8.10567
R7201 a_16434_7468.t24 a_16434_7468.n7 8.10567
R7202 a_16434_7468.t2 a_16434_7468.n4 3.85103
R7203 a_16434_7468.n2 a_16434_7468.t26 8.10567
R7204 a_16434_7468.t26 a_16434_7468.n6 8.10567
R7205 a_16434_7468.t6 a_16434_7468.n16 3.77854
R7206 a_16434_7468.n15 a_16434_7468.n16 0.551084
R7207 a_16434_7468.n20 a_16434_7468.t1 5.48273
R7208 a_16434_7468.n14 a_16434_7468.n20 3.97956
R7209 a_16434_7468.n14 a_16434_7468.t19 3.20383
R7210 a_16434_7468.n9 a_16434_7468.t13 3.20383
R7211 a_16434_7468.n2 a_16434_7468.t11 3.20383
R7212 a_16434_7468.n2 a_16434_7468.t17 3.20383
R7213 a_16434_7468.n2 a_16434_7468.t3 3.20383
R7214 a_16434_7468.n2 a_16434_7468.t7 3.20383
R7215 a_16434_7468.n12 a_16434_7468.t9 3.20383
R7216 a_16434_7468.n10 a_16434_7468.t5 3.20383
R7217 a_16434_7468.n2 a_16434_7468.t15 3.20383
R7218 a_16434_7468.t21 a_16434_7468.n13 3.20383
R7219 a_16434_7468.n6 a_16434_7468.n15 0.913357
R7220 a_16434_7468.n7 a_16434_7468.n6 0.913357
R7221 a_16434_7468.n8 a_16434_7468.n7 0.913357
R7222 a_16434_7468.n8 a_16434_7468.n9 0.913357
R7223 a_16434_7468.n10 a_16434_7468.n18 1.19317
R7224 a_16434_7468.n14 a_16434_7468.n0 1.07565
R7225 a_16434_7468.n5 a_16434_7468.n2 0.478235
R7226 a_16434_7468.n12 a_16434_7468.n11 1.01469
R7227 a_16434_7468.n10 a_16434_7468.n17 1.01469
R7228 a_16434_7468.n3 a_16434_7468.n2 0.478235
R7229 a_16434_7468.n7 a_16434_7468.n1 1.01469
R7230 a_16434_7468.n6 a_16434_7468.n4 1.01469
R7231 a_16434_7468.n19 a_16434_7468.n9 0.978123
R7232 a_16434_7468.n2 a_16434_7468.n16 0.551084
R7233 a_16434_7468.n2 a_16434_7468.n0 0.467078
R7234 a_16434_7468.n12 a_16434_7468.n10 0.913357
R7235 a_16434_7468.n12 a_16434_7468.n13 0.913357
R7236 a_16434_7468.n13 a_16434_7468.n14 0.913357
R7237 a_16434_7468.n11 a_16434_7468.n2 0.822854
R7238 a_16434_7468.n2 a_16434_7468.n17 0.822854
R7239 a_16434_7468.n2 a_16434_7468.n4 0.811729
R7240 a_16434_7468.n2 a_16434_7468.n1 0.811729
R7241 a_16434_7468.n19 a_16434_7468.n2 0.772955
R7242 a_16434_7468.n18 a_16434_7468.n2 0.697056
R7243 a_25891_6334.n6 a_25891_6334.t6 19.7931
R7244 a_25891_6334.t5 a_25891_6334.n6 19.4417
R7245 a_25891_6334.n10 a_25891_6334.t0 18.1584
R7246 a_25891_6334.n8 a_25891_6334.t4 17.4851
R7247 a_25891_6334.n9 a_25891_6334.t2 16.998
R7248 a_25891_6334.t4 a_25891_6334.n7 14.8382
R7249 a_25891_6334.n7 a_25891_6334.t5 14.8163
R7250 a_25891_6334.t1 a_25891_6334.n10 11.4638
R7251 a_25891_6334.n0 a_25891_6334.t3 10.7336
R7252 a_25891_6334.n5 a_25891_6334.n4 2.25359
R7253 a_25891_6334.n2 a_25891_6334.n1 2.2435
R7254 a_25891_6334.n7 a_25891_6334.n3 3.51079
R7255 a_25891_6334.n4 a_25891_6334.n3 2.783
R7256 a_25891_6334.n10 a_25891_6334.n9 1.43621
R7257 a_25891_6334.n6 a_25891_6334.n3 0.404429
R7258 a_25891_6334.n1 a_25891_6334.n0 0.281214
R7259 a_25891_6334.n9 a_25891_6334.n8 0.204071
R7260 a_25891_6334.n8 a_25891_6334.n0 0.154786
R7261 a_25891_6334.n2 a_25891_6334.n5 0.19972
R7262 a_25891_6334.t6 a_25891_6334.n5 14.7562
R7263 a_25891_6334.n4 a_25891_6334.n1 0.249071
R7264 a_25891_6334.n2 a_25891_6334.t2 14.7419
R7265 a_19582_6043.n0 a_19582_6043.t3 30.2519
R7266 a_19582_6043.t3 a_19582_6043.t4 27.8013
R7267 a_19582_6043.n0 a_19582_6043.t2 16.4135
R7268 a_19582_6043.t1 a_19582_6043.n0 14.3567
R7269 a_19582_6043.n0 a_19582_6043.t0 14.3488
R7270 a_25891_n1726.n6 a_25891_n1726.t5 19.7931
R7271 a_25891_n1726.n6 a_25891_n1726.t6 19.4417
R7272 a_25891_n1726.n7 a_25891_n1726.t3 18.1574
R7273 a_25891_n1726.n9 a_25891_n1726.t4 17.4851
R7274 a_25891_n1726.n8 a_25891_n1726.t0 16.998
R7275 a_25891_n1726.n5 a_25891_n1726.t4 14.8382
R7276 a_25891_n1726.t6 a_25891_n1726.n5 14.8163
R7277 a_25891_n1726.n7 a_25891_n1726.t2 11.4638
R7278 a_25891_n1726.t1 a_25891_n1726.n10 10.7346
R7279 a_25891_n1726.n0 a_25891_n1726.n4 2.25359
R7280 a_25891_n1726.n2 a_25891_n1726.n1 2.2435
R7281 a_25891_n1726.n3 a_25891_n1726.n5 3.51079
R7282 a_25891_n1726.n0 a_25891_n1726.n3 2.783
R7283 a_25891_n1726.n8 a_25891_n1726.n7 1.43621
R7284 a_25891_n1726.n3 a_25891_n1726.n6 0.404429
R7285 a_25891_n1726.n10 a_25891_n1726.n1 0.281214
R7286 a_25891_n1726.n9 a_25891_n1726.n8 0.204071
R7287 a_25891_n1726.n10 a_25891_n1726.n9 0.154786
R7288 a_25891_n1726.n2 a_25891_n1726.n4 0.19972
R7289 a_25891_n1726.t5 a_25891_n1726.n4 14.7562
R7290 a_25891_n1726.n1 a_25891_n1726.n0 0.249071
R7291 a_25891_n1726.t0 a_25891_n1726.n2 14.7419
R7292 a_9120_14251.n1 a_9120_14251.n0 32.8505
R7293 a_9120_14251.n0 a_9120_14251.t4 28.4659
R7294 a_9120_14251.n0 a_9120_14251.t5 19.2698
R7295 a_9120_14251.n0 a_9120_14251.t6 19.2698
R7296 a_9120_14251.n0 a_9120_14251.t7 19.2698
R7297 a_9120_14251.n0 a_9120_14251.t8 19.2698
R7298 a_9120_14251.n1 a_9120_14251.t1 18.2981
R7299 a_9120_14251.n0 a_9120_14251.t3 17.8802
R7300 a_9120_14251.n0 a_9120_14251.t2 16.9973
R7301 a_9120_14251.n0 a_9120_14251.t9 16.9973
R7302 a_9120_14251.t0 a_9120_14251.n1 15.1831
R7303 a_21659_n106.n21 a_21659_n106.t15 13.6232
R7304 a_21659_n106.n20 a_21659_n106.t5 13.5679
R7305 a_21659_n106.n16 a_21659_n106.t3 13.5679
R7306 a_21659_n106.n22 a_21659_n106.t9 13.5675
R7307 a_21659_n106.n19 a_21659_n106.t1 13.5675
R7308 a_21659_n106.n18 a_21659_n106.t13 13.5675
R7309 a_21659_n106.n17 a_21659_n106.t12 13.5675
R7310 a_21659_n106.n10 a_21659_n106.t0 13.5644
R7311 a_21659_n106.n12 a_21659_n106.t8 13.5633
R7312 a_21659_n106.n15 a_21659_n106.t10 13.5633
R7313 a_21659_n106.n9 a_21659_n106.t7 13.5633
R7314 a_21659_n106.n13 a_21659_n106.t2 13.5629
R7315 a_21659_n106.n11 a_21659_n106.t11 13.5625
R7316 a_21659_n106.n14 a_21659_n106.t4 13.5596
R7317 a_21659_n106.n23 a_21659_n106.t6 11.4221
R7318 a_21659_n106.n8 a_21659_n106.t14 11.2951
R7319 a_21659_n106.n6 a_21659_n106.n4 4.62286
R7320 a_21659_n106.n3 a_21659_n106.n1 4.62286
R7321 a_21659_n106.n16 a_21659_n106.n15 4.33657
R7322 a_21659_n106.n3 a_21659_n106.n2 3.98468
R7323 a_21659_n106.n6 a_21659_n106.n5 3.98468
R7324 a_21659_n106.n0 a_21659_n106.n7 3.98468
R7325 a_21659_n106.n26 a_21659_n106.n25 3.98468
R7326 a_21659_n106.n24 a_21659_n106.n8 2.97211
R7327 a_21659_n106.n9 a_21659_n106.n8 2.93779
R7328 a_21659_n106.n23 a_21659_n106.n22 2.92
R7329 a_21659_n106.n0 a_21659_n106.n24 1.57764
R7330 a_21659_n106.n25 a_21659_n106.n0 1.51209
R7331 a_21659_n106.n0 a_21659_n106.n6 1.07026
R7332 a_21659_n106.n24 a_21659_n106.n23 0.927751
R7333 a_21659_n106.n1 a_21659_n106.t22 0.9105
R7334 a_21659_n106.n1 a_21659_n106.t23 0.9105
R7335 a_21659_n106.n2 a_21659_n106.t21 0.9105
R7336 a_21659_n106.n2 a_21659_n106.t27 0.9105
R7337 a_21659_n106.n4 a_21659_n106.t17 0.9105
R7338 a_21659_n106.n4 a_21659_n106.t18 0.9105
R7339 a_21659_n106.n5 a_21659_n106.t16 0.9105
R7340 a_21659_n106.n5 a_21659_n106.t24 0.9105
R7341 a_21659_n106.n7 a_21659_n106.t19 0.9105
R7342 a_21659_n106.n7 a_21659_n106.t20 0.9105
R7343 a_21659_n106.n26 a_21659_n106.t25 0.9105
R7344 a_21659_n106.t26 a_21659_n106.n26 0.9105
R7345 a_21659_n106.n22 a_21659_n106.n21 0.763357
R7346 a_21659_n106.n20 a_21659_n106.n19 0.700143
R7347 a_21659_n106.n14 a_21659_n106.n13 0.699071
R7348 a_21659_n106.n13 a_21659_n106.n12 0.692643
R7349 a_21659_n106.n18 a_21659_n106.n17 0.692643
R7350 a_21659_n106.n10 a_21659_n106.n9 0.692328
R7351 a_21659_n106.n12 a_21659_n106.n11 0.689429
R7352 a_21659_n106.n19 a_21659_n106.n18 0.688357
R7353 a_21659_n106.n11 a_21659_n106.n10 0.686971
R7354 a_21659_n106.n17 a_21659_n106.n16 0.686214
R7355 a_21659_n106.n15 a_21659_n106.n14 0.679786
R7356 a_21659_n106.n25 a_21659_n106.n3 0.638674
R7357 a_21659_n106.n21 a_21659_n106.n20 0.608
R7358 a_21743_n1960.n3 a_21743_n1960.t12 8.45596
R7359 a_21743_n1960.n2 a_21743_n1960.t5 15.2205
R7360 a_21743_n1960.n5 a_21743_n1960.t0 13.8811
R7361 a_21743_n1960.n8 a_21743_n1960.t9 13.5061
R7362 a_21743_n1960.t8 a_21743_n1960.n2 13.1505
R7363 a_21743_n1960.n1 a_21743_n1960.t2 13.1484
R7364 a_21743_n1960.n1 a_21743_n1960.t1 13.1473
R7365 a_21743_n1960.n11 a_21743_n1960.t6 13.1473
R7366 a_21743_n1960.n2 a_21743_n1960.t3 13.1459
R7367 a_21743_n1960.n12 a_21743_n1960.t7 13.1426
R7368 a_21743_n1960.n10 a_21743_n1960.t4 10.7513
R7369 a_21743_n1960.n0 a_21743_n1960.t13 10.5704
R7370 a_21743_n1960.n4 a_21743_n1960.t11 10.5629
R7371 a_21743_n1960.n6 a_21743_n1960.t15 10.3448
R7372 a_21743_n1960.n0 a_21743_n1960.t17 8.61428
R7373 a_21743_n1960.n7 a_21743_n1960.t14 8.57979
R7374 a_21743_n1960.n4 a_21743_n1960.t10 8.53382
R7375 a_21743_n1960.n6 a_21743_n1960.t16 8.51529
R7376 a_21743_n1960.n9 a_21743_n1960.n5 4.42661
R7377 a_21743_n1960.n7 a_21743_n1960.n0 4.2562
R7378 a_21743_n1960.n9 a_21743_n1960.n8 3.833
R7379 a_21743_n1960.n8 a_21743_n1960.n4 3.62733
R7380 a_21743_n1960.n3 a_21743_n1960.n6 4.58528
R7381 a_21743_n1960.n10 a_21743_n1960.n9 3.30586
R7382 a_21743_n1960.n11 a_21743_n1960.n10 3.08583
R7383 a_21743_n1960.n1 a_21743_n1960.n11 2.7605
R7384 a_21743_n1960.n2 a_21743_n1960.n12 2.74014
R7385 a_21743_n1960.n0 a_21743_n1960.n5 2.64801
R7386 a_21743_n1960.n12 a_21743_n1960.n1 2.23871
R7387 a_21743_n1960.n4 a_21743_n1960.n7 1.76955
R7388 a_21743_n1960.n0 a_21743_n1960.n3 0.986849
R7389 a_21743_n2608.t0 a_21743_n2608.n5 8.42794
R7390 a_21743_n2608.n4 a_21743_n2608.n5 0.109799
R7391 a_21743_n2608.n3 a_21743_n2608.t2 8.44633
R7392 a_21743_n2608.t11 a_21743_n2608.n13 14.0556
R7393 a_21743_n2608.n2 a_21743_n2608.t12 13.9025
R7394 a_21743_n2608.n10 a_21743_n2608.t13 13.5018
R7395 a_21743_n2608.n13 a_21743_n2608.t6 13.3613
R7396 a_21743_n2608.n0 a_21743_n2608.t8 13.3603
R7397 a_21743_n2608.n0 a_21743_n2608.t7 13.3596
R7398 a_21743_n2608.n12 a_21743_n2608.t5 13.3305
R7399 a_21743_n2608.n1 a_21743_n2608.t9 13.3302
R7400 a_21743_n2608.n1 a_21743_n2608.t10 13.3298
R7401 a_21743_n2608.n11 a_21743_n2608.t4 13.3182
R7402 a_21743_n2608.n6 a_21743_n2608.t15 10.7255
R7403 a_21743_n2608.n3 a_21743_n2608.t3 10.5667
R7404 a_21743_n2608.n4 a_21743_n2608.t1 10.5446
R7405 a_21743_n2608.n6 a_21743_n2608.t17 9.65646
R7406 a_21743_n2608.n9 a_21743_n2608.t14 8.61301
R7407 a_21743_n2608.n8 a_21743_n2608.t16 8.57431
R7408 a_21743_n2608.n2 a_21743_n2608.n10 8.43907
R7409 a_21743_n2608.n10 a_21743_n2608.n4 3.63275
R7410 a_21743_n2608.n0 a_21743_n2608.n12 3.16014
R7411 a_21743_n2608.n5 a_21743_n2608.n9 4.39668
R7412 a_21743_n2608.n11 a_21743_n2608.n2 2.88157
R7413 a_21743_n2608.n13 a_21743_n2608.n0 2.75376
R7414 a_21743_n2608.n1 a_21743_n2608.n11 2.75086
R7415 a_21743_n2608.n3 a_21743_n2608.n2 2.65709
R7416 a_21743_n2608.n7 a_21743_n2608.n3 2.49995
R7417 a_21743_n2608.n7 a_21743_n2608.n6 2.17989
R7418 a_21743_n2608.n12 a_21743_n2608.n1 2.07586
R7419 a_21743_n2608.n8 a_21743_n2608.n7 1.97873
R7420 a_21743_n2608.n9 a_21743_n2608.n8 1.83916
R7421 a_10060_n1528.n12 a_10060_n1528.t34 8.61238
R7422 a_10060_n1528.t83 a_10060_n1528.n13 8.66897
R7423 a_10060_n1528.n14 a_10060_n1528.t18 8.60673
R7424 a_10060_n1528.t67 a_10060_n1528.n15 8.66202
R7425 a_10060_n1528.n6 a_10060_n1528.t45 4.02487
R7426 a_10060_n1528.n4 a_10060_n1528.t71 4.33277
R7427 a_10060_n1528.t11 a_10060_n1528.n6 4.02653
R7428 a_10060_n1528.n6 a_10060_n1528.t7 4.07081
R7429 a_10060_n1528.n6 a_10060_n1528.t1 4.02308
R7430 a_10060_n1528.t96 a_10060_n1528.n6 4.02396
R7431 a_10060_n1528.n6 a_10060_n1528.t65 4.21719
R7432 a_10060_n1528.n6 a_10060_n1528.t82 4.00119
R7433 a_10060_n1528.n6 a_10060_n1528.t89 4.02086
R7434 a_10060_n1528.t76 a_10060_n1528.n6 3.99212
R7435 a_10060_n1528.t19 a_10060_n1528.n6 3.9037
R7436 a_10060_n1528.t53 a_10060_n1528.n6 4.01604
R7437 a_10060_n1528.n6 a_10060_n1528.t20 4.00273
R7438 a_10060_n1528.n6 a_10060_n1528.t39 4.01944
R7439 a_10060_n1528.t40 a_10060_n1528.n6 3.90521
R7440 a_10060_n1528.t93 a_10060_n1528.n6 3.90521
R7441 a_10060_n1528.t21 a_10060_n1528.n6 3.95908
R7442 a_10060_n1528.t41 a_10060_n1528.n6 4.09206
R7443 a_10060_n1528.n6 a_10060_n1528.t63 4.00218
R7444 a_10060_n1528.n6 a_10060_n1528.t54 4.0029
R7445 a_10060_n1528.n6 a_10060_n1528.t37 3.99183
R7446 a_10060_n1528.n6 a_10060_n1528.t64 3.95427
R7447 a_10060_n1528.n6 a_10060_n1528.t56 4.06931
R7448 a_10060_n1528.t80 a_10060_n1528.n6 4.05576
R7449 a_10060_n1528.t13 a_10060_n1528.n6 3.97871
R7450 a_10060_n1528.n6 a_10060_n1528.t90 3.99598
R7451 a_10060_n1528.t26 a_10060_n1528.n6 3.99538
R7452 a_10060_n1528.n2 a_10060_n1528.t73 3.93188
R7453 a_10060_n1528.n9 a_10060_n1528.t22 3.9037
R7454 a_10060_n1528.t62 a_10060_n1528.n6 3.9037
R7455 a_10060_n1528.n3 a_10060_n1528.t16 4.05025
R7456 a_10060_n1528.t81 a_10060_n1528.n6 8.06917
R7457 a_10060_n1528.n2 a_10060_n1528.t81 8.06917
R7458 a_10060_n1528.t95 a_10060_n1528.n2 4.03115
R7459 a_10060_n1528.n5 a_10060_n1528.t74 3.92429
R7460 a_10060_n1528.n5 a_10060_n1528.n8 0.223084
R7461 a_10060_n1528.t92 a_10060_n1528.n8 3.98326
R7462 a_10060_n1528.n6 a_10060_n1528.t33 3.97614
R7463 a_10060_n1528.n0 a_10060_n1528.t91 4.1682
R7464 a_10060_n1528.t17 a_10060_n1528.n6 3.90323
R7465 a_10060_n1528.n0 a_10060_n1528.t36 3.97045
R7466 a_10060_n1528.n1 a_10060_n1528.t27 4.03608
R7467 a_10060_n1528.t55 a_10060_n1528.n2 3.98164
R7468 a_10060_n1528.n0 a_10060_n1528.t46 3.9037
R7469 a_10060_n1528.t28 a_10060_n1528.n2 3.85016
R7470 a_10060_n1528.n1 a_10060_n1528.n0 0.157031
R7471 a_10060_n1528.t57 a_10060_n1528.n0 3.87955
R7472 a_10060_n1528.n7 a_10060_n1528.t47 3.89343
R7473 a_10060_n1528.n7 a_10060_n1528.n0 0.284815
R7474 a_10060_n1528.t75 a_10060_n1528.n0 3.96911
R7475 a_10060_n1528.t58 a_10060_n1528.n0 4.00942
R7476 a_10060_n1528.t14 a_10060_n1528.n0 3.9761
R7477 a_10060_n1528.n0 a_10060_n1528.t29 4.00545
R7478 a_10060_n1528.n0 a_10060_n1528.t59 3.95578
R7479 a_10060_n1528.n0 a_10060_n1528.t48 3.95443
R7480 a_10060_n1528.n0 a_10060_n1528.t77 4.0138
R7481 a_10060_n1528.n0 a_10060_n1528.t69 4.24121
R7482 a_10060_n1528.t49 a_10060_n1528.n0 3.9791
R7483 a_10060_n1528.t78 a_10060_n1528.n0 3.93908
R7484 a_10060_n1528.n0 a_10060_n1528.t70 3.9037
R7485 a_10060_n1528.t86 a_10060_n1528.n0 4.26514
R7486 a_10060_n1528.t30 a_10060_n1528.n0 4.03998
R7487 a_10060_n1528.n0 a_10060_n1528.t87 3.9881
R7488 a_10060_n1528.n0 a_10060_n1528.t15 4.00952
R7489 a_10060_n1528.n0 a_10060_n1528.t31 4.01485
R7490 a_10060_n1528.t24 a_10060_n1528.n0 4.06522
R7491 a_10060_n1528.n0 a_10060_n1528.t51 4.07654
R7492 a_10060_n1528.n0 a_10060_n1528.t42 3.99982
R7493 a_10060_n1528.t25 a_10060_n1528.n0 3.99229
R7494 a_10060_n1528.t52 a_10060_n1528.n0 4.01575
R7495 a_10060_n1528.t43 a_10060_n1528.n0 4.00307
R7496 a_10060_n1528.t72 a_10060_n1528.n0 4.01945
R7497 a_10060_n1528.t94 a_10060_n1528.n0 4.32229
R7498 a_10060_n1528.n0 a_10060_n1528.t23 4.04959
R7499 a_10060_n1528.n0 a_10060_n1528.t9 4.02528
R7500 a_10060_n1528.t3 a_10060_n1528.n0 4.02638
R7501 a_10060_n1528.n0 a_10060_n1528.t5 4.03071
R7502 a_10060_n1528.t38 a_10060_n1528.n0 4.04387
R7503 a_10060_n1528.t66 a_10060_n1528.n0 4.33661
R7504 a_10060_n1528.t60 a_10060_n1528.n0 4.02396
R7505 a_10060_n1528.n12 a_10060_n1528.t84 8.06917
R7506 a_10060_n1528.t68 a_10060_n1528.n14 8.06917
R7507 a_10060_n1528.t84 a_10060_n1528.n18 5.4025
R7508 a_10060_n1528.n18 a_10060_n1528.t68 5.4025
R7509 a_10060_n1528.n22 a_10060_n1528.t34 5.4025
R7510 a_10060_n1528.t18 a_10060_n1528.n22 5.4025
R7511 a_10060_n1528.n20 a_10060_n1528.t67 5.4025
R7512 a_10060_n1528.n20 a_10060_n1528.t83 5.4025
R7513 a_10060_n1528.n23 a_10060_n1528.n15 4.50199
R7514 a_10060_n1528.n15 a_10060_n1528.n14 0.0557981
R7515 a_10060_n1528.n21 a_10060_n1528.n11 4.50135
R7516 a_10060_n1528.n10 a_10060_n1528.n11 0.0570868
R7517 a_10060_n1528.n13 a_10060_n1528.n19 4.50135
R7518 a_10060_n1528.n13 a_10060_n1528.n12 0.0570868
R7519 a_10060_n1528.n0 a_10060_n1528.n24 13.1977
R7520 a_10060_n1528.n0 a_10060_n1528.t0 17.6996
R7521 a_10060_n1528.n6 a_10060_n1528.t2 3.3605
R7522 a_10060_n1528.n6 a_10060_n1528.t8 3.3605
R7523 a_10060_n1528.n0 a_10060_n1528.t10 3.3605
R7524 a_10060_n1528.n0 a_10060_n1528.t4 3.3605
R7525 a_10060_n1528.n0 a_10060_n1528.t6 3.3605
R7526 a_10060_n1528.t12 a_10060_n1528.n6 3.3605
R7527 a_10060_n1528.n11 a_10060_n1528.n20 3.26697
R7528 a_10060_n1528.n22 a_10060_n1528.n10 3.21038
R7529 a_10060_n1528.n18 a_10060_n1528.n10 2.66717
R7530 a_10060_n1528.n19 a_10060_n1528.n17 0.844786
R7531 a_10060_n1528.n19 a_10060_n1528.n16 0.844786
R7532 a_10060_n1528.n23 a_10060_n1528.n17 0.838357
R7533 a_10060_n1528.t61 a_10060_n1528.n6 4.04879
R7534 a_10060_n1528.n3 a_10060_n1528.n6 0.0627636
R7535 a_10060_n1528.n9 a_10060_n1528.n6 0.264263
R7536 a_10060_n1528.n1 a_10060_n1528.n2 0.0724718
R7537 a_10060_n1528.n6 a_10060_n1528.t79 4.00266
R7538 a_10060_n1528.n24 a_10060_n1528.n16 0.538357
R7539 a_10060_n1528.n4 a_10060_n1528.t85 4.04767
R7540 a_10060_n1528.t44 a_10060_n1528.n0 4.02649
R7541 a_10060_n1528.t88 a_10060_n1528.n6 4.04662
R7542 a_10060_n1528.n21 a_10060_n1528.n16 0.3005
R7543 a_10060_n1528.n21 a_10060_n1528.n17 0.3005
R7544 a_10060_n1528.n24 a_10060_n1528.n23 0.3005
R7545 a_10060_n1528.n6 a_10060_n1528.n0 0.490269
R7546 a_10060_n1528.t35 a_10060_n1528.n6 4.03551
R7547 a_10060_n1528.n9 a_10060_n1528.n2 0.684037
R7548 a_10060_n1528.n6 a_10060_n1528.n5 0.640764
R7549 a_10060_n1528.n8 a_10060_n1528.n2 0.637579
R7550 a_10060_n1528.n7 a_10060_n1528.n8 0.284815
R7551 a_10060_n1528.n6 a_10060_n1528.t50 4.05843
R7552 a_10060_n1528.n2 a_10060_n1528.n3 0.162217
R7553 a_10060_n1528.n6 a_10060_n1528.n4 0.577923
R7554 a_10060_n1528.t32 a_10060_n1528.n6 4.32986
R7555 a_9938_8092.n44 a_9938_8092.t0 13.9633
R7556 a_9938_8092.n33 a_9938_8092.t2 13.3633
R7557 a_9938_8092.n0 a_9938_8092.t4 11.6211
R7558 a_9938_8092.n6 a_9938_8092.t1 9.76971
R7559 a_9938_8092.n38 a_9938_8092.t5 9.76971
R7560 a_9938_8092.n49 a_9938_8092.t38 8.844
R7561 a_9938_8092.n39 a_9938_8092.t15 8.844
R7562 a_9938_8092.n1 a_9938_8092.t26 8.844
R7563 a_9938_8092.n7 a_9938_8092.t18 8.844
R7564 a_9938_8092.n10 a_9938_8092.t45 8.844
R7565 a_9938_8092.n13 a_9938_8092.t31 8.844
R7566 a_9938_8092.n18 a_9938_8092.t8 8.844
R7567 a_9938_8092.n25 a_9938_8092.t42 8.844
R7568 a_9938_8092.n47 a_9938_8092.t9 7.91829
R7569 a_9938_8092.n48 a_9938_8092.t16 7.91829
R7570 a_9938_8092.n52 a_9938_8092.t12 7.91829
R7571 a_9938_8092.n51 a_9938_8092.t13 7.91829
R7572 a_9938_8092.n50 a_9938_8092.t10 7.91829
R7573 a_9938_8092.n49 a_9938_8092.t29 7.91829
R7574 a_9938_8092.n6 a_9938_8092.t3 7.91829
R7575 a_9938_8092.n0 a_9938_8092.t6 7.91829
R7576 a_9938_8092.n38 a_9938_8092.t7 7.91829
R7577 a_9938_8092.n43 a_9938_8092.t47 7.91829
R7578 a_9938_8092.n42 a_9938_8092.t33 7.91829
R7579 a_9938_8092.n41 a_9938_8092.t44 7.91829
R7580 a_9938_8092.n40 a_9938_8092.t55 7.91829
R7581 a_9938_8092.n39 a_9938_8092.t41 7.91829
R7582 a_9938_8092.n5 a_9938_8092.t50 7.91829
R7583 a_9938_8092.n4 a_9938_8092.t53 7.91829
R7584 a_9938_8092.n3 a_9938_8092.t48 7.91829
R7585 a_9938_8092.n2 a_9938_8092.t51 7.91829
R7586 a_9938_8092.n1 a_9938_8092.t19 7.91829
R7587 a_9938_8092.n9 a_9938_8092.t39 7.91829
R7588 a_9938_8092.n8 a_9938_8092.t46 7.91829
R7589 a_9938_8092.n7 a_9938_8092.t14 7.91829
R7590 a_9938_8092.n12 a_9938_8092.t43 7.91829
R7591 a_9938_8092.n11 a_9938_8092.t49 7.91829
R7592 a_9938_8092.n10 a_9938_8092.t35 7.91829
R7593 a_9938_8092.n17 a_9938_8092.t28 7.91829
R7594 a_9938_8092.n16 a_9938_8092.t36 7.91829
R7595 a_9938_8092.n15 a_9938_8092.t22 7.91829
R7596 a_9938_8092.n14 a_9938_8092.t30 7.91829
R7597 a_9938_8092.n13 a_9938_8092.t21 7.91829
R7598 a_9938_8092.n24 a_9938_8092.t32 7.91829
R7599 a_9938_8092.n23 a_9938_8092.t40 7.91829
R7600 a_9938_8092.n22 a_9938_8092.t27 7.91829
R7601 a_9938_8092.n21 a_9938_8092.t37 7.91829
R7602 a_9938_8092.n20 a_9938_8092.t24 7.91829
R7603 a_9938_8092.n19 a_9938_8092.t34 7.91829
R7604 a_9938_8092.n18 a_9938_8092.t52 7.91829
R7605 a_9938_8092.n29 a_9938_8092.t25 7.91829
R7606 a_9938_8092.n28 a_9938_8092.t17 7.91829
R7607 a_9938_8092.n27 a_9938_8092.t23 7.91829
R7608 a_9938_8092.n26 a_9938_8092.t11 7.91829
R7609 a_9938_8092.n25 a_9938_8092.t20 7.91829
R7610 a_9938_8092.t54 a_9938_8092.n53 7.91829
R7611 a_9938_8092.n30 a_9938_8092.n29 5.40264
R7612 a_9938_8092.n8 a_9938_8092.n7 4.62907
R7613 a_9938_8092.n11 a_9938_8092.n10 4.62907
R7614 a_9938_8092.n35 a_9938_8092.n6 4.51979
R7615 a_9938_8092.n45 a_9938_8092.n38 4.51802
R7616 a_9938_8092.n44 a_9938_8092.n43 4.50264
R7617 a_9938_8092.n37 a_9938_8092.n0 3.59407
R7618 a_9938_8092.n36 a_9938_8092.n5 3.57693
R7619 a_9938_8092.n34 a_9938_8092.n9 3.57693
R7620 a_9938_8092.n32 a_9938_8092.n12 3.57693
R7621 a_9938_8092.n31 a_9938_8092.n17 3.57693
R7622 a_9938_8092.n30 a_9938_8092.n24 3.57693
R7623 a_9938_8092.n47 a_9938_8092.n46 3.57693
R7624 a_9938_8092.n33 a_9938_8092.n32 3.3005
R7625 a_9938_8092.n3 a_9938_8092.n2 2.77764
R7626 a_9938_8092.n15 a_9938_8092.n14 2.77764
R7627 a_9938_8092.n43 a_9938_8092.n42 0.926214
R7628 a_9938_8092.n42 a_9938_8092.n41 0.926214
R7629 a_9938_8092.n41 a_9938_8092.n40 0.926214
R7630 a_9938_8092.n40 a_9938_8092.n39 0.926214
R7631 a_9938_8092.n5 a_9938_8092.n4 0.926214
R7632 a_9938_8092.n4 a_9938_8092.n3 0.926214
R7633 a_9938_8092.n2 a_9938_8092.n1 0.926214
R7634 a_9938_8092.n9 a_9938_8092.n8 0.926214
R7635 a_9938_8092.n12 a_9938_8092.n11 0.926214
R7636 a_9938_8092.n17 a_9938_8092.n16 0.926214
R7637 a_9938_8092.n16 a_9938_8092.n15 0.926214
R7638 a_9938_8092.n14 a_9938_8092.n13 0.926214
R7639 a_9938_8092.n24 a_9938_8092.n23 0.926214
R7640 a_9938_8092.n23 a_9938_8092.n22 0.926214
R7641 a_9938_8092.n22 a_9938_8092.n21 0.926214
R7642 a_9938_8092.n21 a_9938_8092.n20 0.926214
R7643 a_9938_8092.n20 a_9938_8092.n19 0.926214
R7644 a_9938_8092.n19 a_9938_8092.n18 0.926214
R7645 a_9938_8092.n29 a_9938_8092.n28 0.926214
R7646 a_9938_8092.n28 a_9938_8092.n27 0.926214
R7647 a_9938_8092.n27 a_9938_8092.n26 0.926214
R7648 a_9938_8092.n26 a_9938_8092.n25 0.926214
R7649 a_9938_8092.n48 a_9938_8092.n47 0.926214
R7650 a_9938_8092.n53 a_9938_8092.n48 0.926214
R7651 a_9938_8092.n53 a_9938_8092.n52 0.926214
R7652 a_9938_8092.n52 a_9938_8092.n51 0.926214
R7653 a_9938_8092.n51 a_9938_8092.n50 0.926214
R7654 a_9938_8092.n50 a_9938_8092.n49 0.926214
R7655 a_9938_8092.n31 a_9938_8092.n30 0.9005
R7656 a_9938_8092.n32 a_9938_8092.n31 0.9005
R7657 a_9938_8092.n35 a_9938_8092.n34 0.6005
R7658 a_9938_8092.n37 a_9938_8092.n36 0.6005
R7659 a_9938_8092.n46 a_9938_8092.n45 0.599429
R7660 a_9938_8092.n45 a_9938_8092.n44 0.301571
R7661 a_9938_8092.n34 a_9938_8092.n33 0.3005
R7662 a_9938_8092.n36 a_9938_8092.n35 0.3005
R7663 a_9938_8092.n46 a_9938_8092.n37 0.3005
R7664 a_11618_8092.n1 a_11618_8092.t0 24.1799
R7665 a_11618_8092.n0 a_11618_8092.t1 6.53667
R7666 a_11618_8092.n0 a_11618_8092.t6 6.53667
R7667 a_11618_8092.t5 a_11618_8092.n1 6.53667
R7668 a_11618_8092.n1 a_11618_8092.t4 5.61135
R7669 a_11618_8092.n0 a_11618_8092.t2 5.61135
R7670 a_11618_8092.n0 a_11618_8092.t3 5.61135
R7671 a_11618_8092.n1 a_11618_8092.n0 3.04062
R7672 OUT OUT.t0 1.5334
R7673 a_19582_6479.t4 a_19582_6479.t5 27.8013
R7674 a_19582_6479.n0 a_19582_6479.t4 17.911
R7675 a_19582_6479.n0 a_19582_6479.t3 13.7109
R7676 a_19582_6479.t0 a_19582_6479.n0 11.1076
R7677 a_19582_6479.n0 a_19582_6479.t2 10.5905
R7678 a_19582_6479.n0 a_19582_6479.t1 10.5905
R7679 a_10778_8092.n9 a_10778_8092.t15 8.844
R7680 a_10778_8092.n6 a_10778_8092.t7 8.844
R7681 a_10778_8092.t26 a_10778_8092.n24 8.844
R7682 a_10778_8092.n0 a_10778_8092.n17 8.48173
R7683 a_10778_8092.n22 a_10778_8092.t18 7.91829
R7684 a_10778_8092.n23 a_10778_8092.t9 7.91829
R7685 a_10778_8092.n11 a_10778_8092.t25 7.91829
R7686 a_10778_8092.n10 a_10778_8092.t17 7.91829
R7687 a_10778_8092.n9 a_10778_8092.t22 7.91829
R7688 a_10778_8092.n8 a_10778_8092.t14 7.91829
R7689 a_10778_8092.n7 a_10778_8092.t6 7.91829
R7690 a_10778_8092.n6 a_10778_8092.t10 7.91829
R7691 a_10778_8092.n24 a_10778_8092.t13 7.91829
R7692 a_10778_8092.n15 a_10778_8092.t1 7.34667
R7693 a_10778_8092.n16 a_10778_8092.t0 6.78437
R7694 a_10778_8092.n18 a_10778_8092.t24 6.55326
R7695 a_10778_8092.n12 a_10778_8092.t19 6.55326
R7696 a_10778_8092.n1 a_10778_8092.t20 6.55326
R7697 a_10778_8092.n4 a_10778_8092.t4 6.55326
R7698 a_10778_8092.n18 a_10778_8092.t27 5.62796
R7699 a_10778_8092.n13 a_10778_8092.t21 5.62796
R7700 a_10778_8092.n12 a_10778_8092.t8 5.62796
R7701 a_10778_8092.n14 a_10778_8092.t11 5.62796
R7702 a_10778_8092.n1 a_10778_8092.t5 5.62796
R7703 a_10778_8092.n2 a_10778_8092.t23 5.62796
R7704 a_10778_8092.n3 a_10778_8092.t16 5.62796
R7705 a_10778_8092.n4 a_10778_8092.t12 5.62796
R7706 a_10778_8092.n17 a_10778_8092.t3 5.61135
R7707 a_10778_8092.n15 a_10778_8092.t2 5.61135
R7708 a_10778_8092.n5 a_10778_8092.n4 4.40815
R7709 a_10778_8092.n0 a_10778_8092.n18 3.96458
R7710 a_10778_8092.n19 a_10778_8092.n11 3.90693
R7711 a_10778_8092.n20 a_10778_8092.n8 3.90693
R7712 a_10778_8092.n22 a_10778_8092.n21 3.90693
R7713 a_10778_8092.n10 a_10778_8092.n9 2.77764
R7714 a_10778_8092.n7 a_10778_8092.n6 2.77764
R7715 a_10778_8092.n24 a_10778_8092.n23 2.77764
R7716 a_10778_8092.n0 a_10778_8092.n14 2.58244
R7717 a_10778_8092.n5 a_10778_8092.n3 2.58244
R7718 a_10778_8092.n19 a_10778_8092.n0 1.19407
R7719 a_10778_8092.n16 a_10778_8092.n15 1.17352
R7720 a_10778_8092.n21 a_10778_8092.n5 1.0505
R7721 a_10778_8092.n11 a_10778_8092.n10 0.926214
R7722 a_10778_8092.n8 a_10778_8092.n7 0.926214
R7723 a_10778_8092.n23 a_10778_8092.n22 0.926214
R7724 a_10778_8092.n14 a_10778_8092.n13 0.925799
R7725 a_10778_8092.n13 a_10778_8092.n12 0.925799
R7726 a_10778_8092.n3 a_10778_8092.n2 0.925799
R7727 a_10778_8092.n2 a_10778_8092.n1 0.925799
R7728 a_10778_8092.n21 a_10778_8092.n20 0.9005
R7729 a_10778_8092.n20 a_10778_8092.n19 0.9005
R7730 a_10778_8092.n17 a_10778_8092.n16 0.562801
R7731 a_16434_8348.t10 a_16434_8348.n9 9.12983
R7732 a_16434_8348.n8 a_16434_8348.t7 8.2159
R7733 a_16434_8348.n6 a_16434_8348.t9 8.2159
R7734 a_16434_8348.n4 a_16434_8348.t3 8.2159
R7735 a_16434_8348.n2 a_16434_8348.t11 8.2159
R7736 a_16434_8348.n3 a_16434_8348.t5 8.16019
R7737 a_16434_8348.n5 a_16434_8348.t8 8.16019
R7738 a_16434_8348.n7 a_16434_8348.t2 8.16019
R7739 a_16434_8348.n9 a_16434_8348.t4 8.16019
R7740 a_16434_8348.n0 a_16434_8348.t1 7.22
R7741 a_16434_8348.n1 a_16434_8348.t6 5.48273
R7742 a_16434_8348.n0 a_16434_8348.t0 5.45468
R7743 a_16434_8348.n2 a_16434_8348.n1 3.59082
R7744 a_16434_8348.n1 a_16434_8348.n0 3.29349
R7745 a_16434_8348.n8 a_16434_8348.n7 0.913357
R7746 a_16434_8348.n7 a_16434_8348.n6 0.913357
R7747 a_16434_8348.n6 a_16434_8348.n5 0.913357
R7748 a_16434_8348.n5 a_16434_8348.n4 0.913357
R7749 a_16434_8348.n4 a_16434_8348.n3 0.913357
R7750 a_16434_8348.n3 a_16434_8348.n2 0.913357
R7751 a_16434_8348.n9 a_16434_8348.n8 0.912286
R7752 a_19582_7363.n0 a_19582_7363.t4 45.8134
R7753 a_19582_7363.t4 a_19582_7363.t3 27.8013
R7754 a_19582_7363.n0 a_19582_7363.t0 16.4111
R7755 a_19582_7363.t2 a_19582_7363.n0 14.3567
R7756 a_19582_7363.n0 a_19582_7363.t1 14.3498
R7757 IBIAS.t0 IBIAS.n45 8.06917
R7758 IBIAS.n46 IBIAS.t0 8.06917
R7759 IBIAS.t9 IBIAS.n31 8.06917
R7760 IBIAS.n32 IBIAS.t9 8.06917
R7761 IBIAS.n46 IBIAS.t4 8.06917
R7762 IBIAS.n28 IBIAS.t4 8.06917
R7763 IBIAS.n31 IBIAS.t8 8.06917
R7764 IBIAS.n8 IBIAS.t8 8.06917
R7765 IBIAS.n18 IBIAS.t11 8.06917
R7766 IBIAS.t11 IBIAS.n17 8.06917
R7767 IBIAS.n28 IBIAS.t6 8.06917
R7768 IBIAS.t6 IBIAS.n27 8.06917
R7769 IBIAS.t10 IBIAS.n8 8.06917
R7770 IBIAS.n21 IBIAS.t10 8.06917
R7771 IBIAS.t14 IBIAS.n18 8.06917
R7772 IBIAS.n19 IBIAS.t14 8.06917
R7773 IBIAS.t3 IBIAS.n21 8.06917
R7774 IBIAS.n22 IBIAS.t3 8.06917
R7775 IBIAS.n27 IBIAS.t2 8.06917
R7776 IBIAS.n24 IBIAS.t2 8.06917
R7777 IBIAS.n19 IBIAS.t7 8.06917
R7778 IBIAS.t7 IBIAS.n13 8.06917
R7779 IBIAS.n22 IBIAS.t5 8.06917
R7780 IBIAS.t5 IBIAS.n10 8.06917
R7781 IBIAS.n38 IBIAS.n4 4.5005
R7782 IBIAS.n37 IBIAS.n36 4.5005
R7783 IBIAS.n35 IBIAS.n5 4.5005
R7784 IBIAS.n34 IBIAS.n33 4.5005
R7785 IBIAS.n44 IBIAS.n43 4.5005
R7786 IBIAS.n42 IBIAS.n3 4.5005
R7787 IBIAS.n25 IBIAS.t13 4.13523
R7788 IBIAS.n14 IBIAS.t12 4.13523
R7789 IBIAS.n39 IBIAS.t1 3.3605
R7790 IBIAS.n41 IBIAS.n40 2.22296
R7791 IBIAS.n34 IBIAS.n6 1.26744
R7792 IBIAS.n43 IBIAS.n0 1.26744
R7793 IBIAS.n17 IBIAS.n15 0.994786
R7794 IBIAS.n26 IBIAS.n24 0.994786
R7795 IBIAS.n13 IBIAS.n12 0.994786
R7796 IBIAS.n23 IBIAS.n10 0.994786
R7797 IBIAS.n11 IBIAS.n10 0.993714
R7798 IBIAS.n7 IBIAS.n6 0.765244
R7799 IBIAS IBIAS.n47 0.558714
R7800 IBIAS.n16 IBIAS.n7 0.544786
R7801 IBIAS.n23 IBIAS.n9 0.544786
R7802 IBIAS.n20 IBIAS.n11 0.544786
R7803 IBIAS.n47 IBIAS.n1 0.544786
R7804 IBIAS.n30 IBIAS.n29 0.544786
R7805 IBIAS.n13 IBIAS.n11 0.417189
R7806 IBIAS.n17 IBIAS.n7 0.416118
R7807 IBIAS.n24 IBIAS.n23 0.416118
R7808 IBIAS.n32 IBIAS.n6 0.219765
R7809 IBIAS.n45 IBIAS.n0 0.219765
R7810 IBIAS.n26 IBIAS.n25 0.218332
R7811 IBIAS.n14 IBIAS.n12 0.218332
R7812 IBIAS.n15 IBIAS.n14 0.21832
R7813 IBIAS.n25 IBIAS.n1 0.21832
R7814 IBIAS IBIAS.n0 0.207029
R7815 IBIAS.n41 IBIAS.n4 0.170649
R7816 IBIAS.n42 IBIAS.n41 0.170649
R7817 IBIAS.n40 IBIAS.n39 0.119429
R7818 IBIAS.n33 IBIAS.n5 0.114071
R7819 IBIAS.n37 IBIAS.n5 0.114071
R7820 IBIAS.n38 IBIAS.n37 0.114071
R7821 IBIAS.n35 IBIAS.n34 0.114071
R7822 IBIAS.n36 IBIAS.n35 0.114071
R7823 IBIAS.n36 IBIAS.n4 0.114071
R7824 IBIAS.n43 IBIAS.n42 0.114071
R7825 IBIAS.n44 IBIAS.n3 0.114071
R7826 IBIAS.n20 IBIAS.n19 0.107232
R7827 IBIAS.n19 IBIAS.n12 0.106979
R7828 IBIAS.n21 IBIAS.n9 0.106979
R7829 IBIAS.n27 IBIAS.n9 0.106979
R7830 IBIAS.n27 IBIAS.n26 0.106979
R7831 IBIAS.n21 IBIAS.n20 0.106725
R7832 IBIAS.n23 IBIAS.n22 0.10668
R7833 IBIAS.n31 IBIAS.n7 0.10668
R7834 IBIAS.n31 IBIAS.n30 0.10668
R7835 IBIAS.n47 IBIAS.n46 0.10668
R7836 IBIAS.n22 IBIAS.n11 0.106427
R7837 IBIAS.n18 IBIAS.n15 0.106382
R7838 IBIAS.n18 IBIAS.n16 0.106382
R7839 IBIAS.n16 IBIAS.n8 0.106382
R7840 IBIAS.n29 IBIAS.n8 0.106382
R7841 IBIAS.n29 IBIAS.n28 0.106382
R7842 IBIAS.n28 IBIAS.n1 0.106382
R7843 IBIAS.n39 IBIAS.n2 0.102554
R7844 IBIAS.n40 IBIAS.n3 0.0894286
R7845 IBIAS.n46 IBIAS.n2 0.0889831
R7846 IBIAS.n33 IBIAS.n32 0.053
R7847 IBIAS.n45 IBIAS.n44 0.053
R7848 IBIAS.n30 IBIAS.n2 0.0181966
R7849 IBIAS.n40 IBIAS.n38 0.0122857
R7850 a_10460_8092.n1 a_10460_8092.t7 13.9
R7851 a_10460_8092.n1 a_10460_8092.t2 12.4044
R7852 a_10460_8092.n2 a_10460_8092.n4 10.9246
R7853 a_10460_8092.n1 a_10460_8092.t9 10.9095
R7854 a_10460_8092.n3 a_10460_8092.t6 10.9296
R7855 a_10460_8092.n4 a_10460_8092.t0 7.68524
R7856 a_10460_8092.n2 a_10460_8092.t3 6.73722
R7857 a_10460_8092.t8 a_10460_8092.n1 5.78102
R7858 a_10460_8092.n1 a_10460_8092.t5 5.63939
R7859 a_10460_8092.n4 a_10460_8092.t1 5.61135
R7860 a_10460_8092.n0 a_10460_8092.n3 0.119086
R7861 a_10460_8092.n0 a_10460_8092.n2 0.9005
R7862 a_10460_8092.t4 a_10460_8092.n3 5.74338
R7863 a_10460_8092.n1 a_10460_8092.n0 2.47915
R7864 a_9248_11691.t0 a_9248_11691.t1 39.5206
R7865 a_9248_11691.t0 a_9248_11691.n1 36.848
R7866 a_9248_11691.n0 a_9248_11691.t6 20.1527
R7867 a_9248_11691.n1 a_9248_11691.t4 19.2698
R7868 a_9248_11691.n0 a_9248_11691.t3 19.2698
R7869 a_9248_11691.n1 a_9248_11691.t5 19.2698
R7870 a_9248_11691.n1 a_9248_11691.t7 16.9973
R7871 a_9248_11691.n1 a_9248_11691.t9 16.9973
R7872 a_9248_11691.n0 a_9248_11691.t8 16.9973
R7873 a_9248_11691.n0 a_9248_11691.t2 16.9973
R7874 a_9248_11691.n1 a_9248_11691.n0 11.4691
C0 VDD OUT 1.85953f
C1 w_23841_n458# VDD 53.0454f
C2 w_15348_6286# VDD 37.9712f
C3 dw_7680_n4606# VDD 16.9601f
C4 OUT GND 3.54746f
C5 IBIAS GND 25.426878f
C6 VDD GND 0.231527p
C7 w_23841_n458# GND 0.165642p
C8 w_15348_6286# GND 0.153798p
C9 a_9248_11691.t0 GND 21.0358f
C10 a_9248_11691.n0 GND 1.61236f
C11 a_9248_11691.n1 GND 6.73324f
C12 a_9248_11691.t1 GND 3.97576f
C13 a_10460_8092.n1 GND 3.21967f
C14 a_10460_8092.n2 GND 1.58139f
C15 a_10460_8092.n4 GND 1.69928f
C16 a_19582_7363.n0 GND 4.51519f
C17 a_19582_7363.t4 GND 1.24671f
C18 a_10778_8092.n0 GND 1.83283f
C19 a_10778_8092.n4 GND 1.2861f
C20 a_10778_8092.n5 GND 1.22638f
C21 a_10778_8092.n18 GND 1.21782f
C22 OUT.t0 GND 5.3846f
C23 a_11618_8092.n0 GND 1.52895f
C24 a_11618_8092.n1 GND 2.81759f
C25 a_11618_8092.t0 GND 1.58708f
C26 a_9938_8092.n0 GND 1.35804f
C27 a_9938_8092.n6 GND 1.15116f
C28 a_9938_8092.n7 GND 1.10136f
C29 a_9938_8092.n10 GND 1.10136f
C30 a_9938_8092.n33 GND 1.25963f
C31 a_9938_8092.n38 GND 1.13846f
C32 a_9938_8092.n44 GND 1.17122f
C33 a_10060_n1528.n0 GND 16.8616f
C34 a_10060_n1528.n2 GND 2.51493f
C35 a_10060_n1528.n6 GND 16.712f
C36 a_21743_n2608.n0 GND 1.69696f
C37 a_21743_n2608.n1 GND 1.4942f
C38 a_21743_n2608.n2 GND 1.84456f
C39 a_21743_n2608.n3 GND 1.03842f
C40 a_21743_n2608.n6 GND 1.61068f
C41 a_21743_n2608.n9 GND 1.09151f
C42 a_21743_n2608.n10 GND 1.69126f
C43 a_21743_n2608.n11 GND 1.01041f
C44 a_21743_n2608.n12 GND 1.16017f
C45 a_21743_n2608.n13 GND 1.17717f
C46 a_21743_n1960.n0 GND 1.11113f
C47 a_21743_n1960.n2 GND 1.26257f
C48 a_21743_n1960.n6 GND 1.0284f
C49 a_21659_n106.n0 GND 1.01769f
C50 a_21659_n106.n8 GND 1.2138f
C51 a_21659_n106.n15 GND 1.5121f
C52 a_21659_n106.n16 GND 1.51445f
C53 a_21659_n106.n24 GND 1.17766f
C54 a_9120_14251.n0 GND 12.1644f
C55 a_9120_14251.n1 GND 11.8027f
C56 a_9120_14251.t0 GND 1.6182f
C57 a_25891_n1726.n7 GND 1.34194f
C58 a_19582_6043.n0 GND 2.34752f
C59 a_25891_6334.n10 GND 1.34195f
C60 a_16434_7468.n2 GND 12.7474f
C61 a_16434_7468.n14 GND 1.36177f
C62 a_11300_8092.n0 GND 1.41472f
C63 a_11300_8092.t5 GND 2.7079f
C64 VDD.n493 GND 1.03229f
C65 VDD.t16 GND 1.16547f
C66 VDD.t26 GND 1.16547f
C67 VDD.n495 GND 1.03229f
C68 VDD.n548 GND 1.03229f
C69 VDD.t4 GND 1.16547f
C70 VDD.t10 GND 1.16547f
C71 VDD.n550 GND 1.03229f
C72 VDD.n557 GND 1.61472f
C73 VDD.n575 GND 37.7025f
C74 VDD.n582 GND 17.0505f
C75 VDD.n871 GND 14.6204f
C76 VDD.n872 GND 8.29386f
C77 VDD.t1 GND 1.12118f
C78 VDD.n936 GND 1.99441f
C79 a_11345_12294.t0 GND 5.66055f
C80 a_11345_12294.t3 GND 14.368199f
C81 a_11345_12294.t2 GND 14.1238f
C82 a_11345_12294.t4 GND 1.16198f
C83 a_21659_3242.n0 GND 2.34034f
C84 a_21659_3242.n1 GND 2.34458f
C85 a_21659_3242.n2 GND 1.47921f
C86 a_21659_3242.n3 GND 2.25342f
C87 a_21659_3242.n4 GND 1.48038f
C88 a_21659_3242.n5 GND 2.23095f
C89 a_21659_3242.n6 GND 1.04999f
C90 a_21659_3242.n8 GND 1.01769f
C91 a_21659_3242.n16 GND 1.17766f
C92 a_21659_3242.n17 GND 1.21379f
C93 a_21743_6100.n0 GND 1.35102f
C94 a_21743_6100.n1 GND 5.4767f
C95 a_21743_6100.n2 GND 3.40422f
C96 a_21743_6748.n0 GND 6.50468f
C97 a_21743_6748.n1 GND 6.76473f
C98 a_21743_6748.n2 GND 2.76095f
C99 a_16964_8348.t0 GND 41.9053f
.ends

