** sch_path: /home/gmaranhao/Desktop/Bracolin/Voltage_Reference/LDO/Pass_tran.sch
.subckt Pass_tran VDD D G
*.PININFO VDD:B D:B G:B
M1[1] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[2] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[3] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[4] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[5] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[6] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[7] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[8] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[9] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[10] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[11] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[12] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[13] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[14] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[15] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[16] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[17] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[18] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[19] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[20] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[21] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[22] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[23] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[24] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[25] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[26] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[27] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[28] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[29] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[30] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[31] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[32] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[33] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[34] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[35] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[36] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[37] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[38] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[39] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[40] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[41] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[42] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[43] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[44] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[45] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[46] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[47] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[48] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[49] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[50] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[51] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[52] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[53] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[54] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[55] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[56] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[57] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[58] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[59] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[60] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[61] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[62] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[63] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[64] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[65] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[66] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[67] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[68] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[69] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[70] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[71] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[72] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[73] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[74] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[75] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[76] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[77] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[78] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[79] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[80] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[81] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[82] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[83] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[84] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[85] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[86] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[87] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[88] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[89] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[90] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[91] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[92] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[93] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[94] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[95] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[96] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[97] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[98] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[99] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[100] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[101] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[102] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[103] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[104] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[105] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[106] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[107] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[108] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[109] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[110] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[111] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[112] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[113] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[114] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[115] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[116] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[117] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[118] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[119] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[120] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[121] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[122] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[123] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[124] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[125] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[126] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[127] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[128] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[129] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[130] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[131] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[132] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[133] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[134] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[135] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[136] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[137] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[138] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[139] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[140] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[141] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[142] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[143] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[144] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[145] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[146] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[147] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[148] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[149] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[150] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[151] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[152] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[153] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[154] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[155] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[156] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[157] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[158] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[159] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[160] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[161] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[162] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[163] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[164] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[165] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[166] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[167] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[168] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[169] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[170] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[171] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[172] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[173] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[174] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[175] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[176] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[177] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[178] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[179] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[180] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[181] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[182] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[183] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[184] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[185] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[186] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[187] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[188] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[189] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[190] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[191] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[192] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[193] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[194] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[195] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[196] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[197] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[198] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[199] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
M1[200] D G VDD VDD pfet_03v3 L=1u W=16u nf=1 m=1
.ends
.end
