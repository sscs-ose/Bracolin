* Extracted by KLayout with GF180MCU LVS runset on : 15/03/2024 18:23

.SUBCKT CM_input VSS ISBCS IP IP2 VDD IN IN2

M1[1] ISBCS ISBCS net1[1] VSS nfet_03v3 L=6u W=2u nf=1 m=1
M1[2] ISBCS ISBCS net1[0] VSS nfet_03v3 L=6u W=2u nf=1 m=1
M2[1] vgp vgp net5[1] VDD pfet_03v3 L=6u W=2u nf=1 m=1
M2[2] vgp vgp net5[0] VDD pfet_03v3 L=6u W=2u nf=1 m=1
M3[1] net1[1] ISBCS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M3[2] net1[0] ISBCS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M4[1] IP ISBCS net2[1] VSS nfet_03v3 L=6u W=2u nf=1 m=1
M4[2] IP ISBCS net2[0] VSS nfet_03v3 L=6u W=2u nf=1 m=1
M5[1] net2[1] ISBCS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M5[2] net2[0] ISBCS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M6[1] IP2 ISBCS net3[1] VSS nfet_03v3 L=6u W=2u nf=1 m=1
M6[2] IP2 ISBCS net3[0] VSS nfet_03v3 L=6u W=2u nf=1 m=1
M7[1] net3[1] ISBCS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M7[2] net3[0] ISBCS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M8[1] vgp ISBCS net4[1] VSS nfet_03v3 L=6u W=2u nf=1 m=1
M8[2] vgp ISBCS net4[0] VSS nfet_03v3 L=6u W=2u nf=1 m=1
M9[1] net4[1] ISBCS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M9[2] net4[0] ISBCS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M10[1] net5[1] vgp VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M10[2] net5[0] vgp VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M11[1] IN vgp net6[1] VDD pfet_03v3 L=6u W=2u nf=1 m=1
M11[2] IN vgp net6[0] VDD pfet_03v3 L=6u W=2u nf=1 m=1
M12[1] net6[1] vgp VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M12[2] net6[0] vgp VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M13[1] IN2 vgp net7[1] VDD pfet_03v3 L=6u W=2u nf=1 m=1
M13[2] IN2 vgp net7[0] VDD pfet_03v3 L=6u W=2u nf=1 m=1
M16[1] net7[1] vgp VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M16[2] net7[0] vgp VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M14[1] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[2] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[3] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[4] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[5] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[6] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[7] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[8] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[9] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[10] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[11] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[12] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[13] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[14] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[15] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[16] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[17] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[18] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[19] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M14[20] VSS VSS VSS VSS nfet_03v3 L=6u W=2u nf=1 m=1
M15[1] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[2] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[3] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[4] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[5] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[6] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[7] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[8] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[9] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[10] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[11] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[12] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[13] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[14] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[15] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[16] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[17] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
M15[18] VDD VDD VDD VDD pfet_03v3 L=6u W=2u nf=1 m=1
.ENDS CM_input
