* NGSPICE file created from Filter_TOP.ext - technology: gf180mcuD

.subckt Filter_TOP
X0 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1 a_43695_n39042# PRbiased_net_x5_0.IBP1 PRbiased_net_x5_0.ITP1 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2 a_30415_n5302# CM_n_net_1.IN a_29855_n4405# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3 a_94739_n33067# a_83172_n33199# a_96696_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4 a_72648_n11674# a_71318_n10715# CM_input_0.IN CM_input_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X5 a_35879_13393# a_36009_10235# a_37815_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6 a_89378_n34225# a_83000_n40208# a_88856_n34225# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X7 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X8 a_48196_12227# a_47666_10295# a_47666_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X9 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X10 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X11 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X12 a_84976_7410# a_83172_4268# PRbiased_net_x5_1.ITN4 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X13 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X14 a_65360_n16095# CM_n_net_0.IN a_64838_n16095# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X15 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X16 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X17 a_n7828_n20082# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X18 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X19 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X20 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X21 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X22 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X23 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X24 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X25 a_84952_n9617# CM_p_net_0.IN a_84384_n9617# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X26 a_29999_n40208# PRbiased_net_x5_0.IBN1 a_31975_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X27 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X28 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X29 CM_n_net_1.VSS a_71343_10235# a_71743_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X30 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X31 a_29855_n3508# CM_n_net_1.IN a_29333_n4405# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X32 a_100929_n16633# CM_p_net_1.IN a_100399_n17538# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X33 a_84952_n17657# CM_p_net_0.IN a_84384_n17657# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X34 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X35 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X36 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X37 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X38 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X39 PRbiased_net_x5_0.ITP4 PRbiased_net_x5_0.IBP4 a_95290_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X40 a_45255_n20452# CM_n_net_1.IN a_44733_n20452# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X41 a_45255_n17761# CM_n_net_1.IN a_44381_n15967# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X42 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X43 PRbiased_net_x5_1.VDD a_29999_11461# a_37781_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X44 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X45 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X46 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X47 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X48 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X49 a_94942_n22182# CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X50 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X51 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X52 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X53 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X54 a_90082_n22182# CM_p_net_0.IN a_89244_n22182# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X55 a_59094_n16095# CM_n_net_0.IN a_58572_n16095# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X56 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X57 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X58 a_49960_n20580# CM_n_net_0.IN a_49438_n21477# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X59 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X60 a_83546_n4187# CM_p_net_0.IN CM_p_net_0.OUT1 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X61 a_115137_n19348# CM_p_net_1.IN CM_p_net_1.OUT12 CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X62 a_49960_n17889# CM_n_net_0.IN CM_n_net_0.OUT8 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X63 a_n2230_n26552# a_n7828_n21089# a_n2752_n26552# CM_n_net_1.VSS nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X64 a_90650_n5092# CM_p_net_0.IN a_90082_n5092# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X65 a_59094_n9915# CM_n_net_0.IN a_58572_n9915# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X66 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X67 a_83546_n17657# CM_p_net_0.IN a_83016_n17657# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X68 a_112928_n33067# a_112406_n33067# a_112406_n33067# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X69 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X70 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X71 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X72 CM_n_net_1.VSS a_94739_4328# a_95261_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X73 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X74 a_83530_n37110# a_83000_n39042# a_83000_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X75 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X76 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X77 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X78 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X79 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X80 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X81 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X82 a_38989_n20452# CM_n_net_1.IN a_38467_n20452# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X83 a_102335_n20253# CM_p_net_1.IN a_101767_n20253# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X84 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X85 a_38989_n17761# CM_n_net_1.IN a_38115_n15967# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X86 a_37815_n40208# a_36009_n40268# a_35855_n31143# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X87 a_63052_n16095# CM_n_net_0.IN a_62492_n15198# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X88 a_83000_n40208# a_83000_n39042# a_84936_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X89 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X90 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X91 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X92 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X93 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X94 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X95 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X96 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X97 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X98 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X99 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X100 a_36009_n40268# a_41738_n33067# a_43664_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X101 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X102 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X103 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X104 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X105 a_92056_n8712# CM_p_net_0.IN a_91218_n8712# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X106 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X107 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X108 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X109 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X110 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X111 a_100929_n5878# CM_p_net_1.IN a_100399_n5878# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X112 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X113 a_100929_n20253# CM_p_net_1.IN a_100399_n21158# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X114 a_42947_n18658# CM_n_net_1.IN a_42387_n16864# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X115 a_100667_n40208# a_100667_n39042# a_102603_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X116 a_84952_n21277# CM_p_net_0.IN a_84384_n21277# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X117 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X118 a_36409_n40208# a_36009_n40268# a_35879_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X119 a_107465_n9498# CM_p_net_1.IN a_106627_n9498# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X120 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X121 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X122 a_106627_n19348# CM_p_net_1.IN a_106097_n18443# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X123 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X124 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X125 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X126 a_56786_n16095# CM_n_net_0.IN a_56226_n15198# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X127 a_89378_n32301# a_83000_n40208# PRbiased_net_x5_0.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X128 a_61331_6252# a_59405_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X129 a_108601_n4973# CM_p_net_1.IN a_108033_n4973# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X130 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X131 a_114299_n3163# CM_p_net_1.IN a_113731_n3163# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X132 a_53388_n10812# CM_n_net_0.IN a_52828_n10812# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X133 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X134 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X135 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X136 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X137 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X138 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X139 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X140 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X141 a_31935_13393# a_29999_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X142 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X143 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X144 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X145 a_54076_13393# a_53676_10235# a_53546_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X146 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X147 PRbiased_net_x5_1.VDD a_65333_10295# a_65863_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X148 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X149 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X150 a_29999_n40208# PRbiased_net_x5_0.IBN1 a_31975_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X151 a_106627_n7688# CM_p_net_1.IN a_106097_n6783# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X152 a_102903_n17538# CM_p_net_1.IN a_102335_n17538# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X153 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X154 a_83546_n21277# CM_p_net_0.IN a_83016_n21277# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X155 PRbiased_net_x5_0.VDD a_100667_n39042# a_101197_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X156 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X157 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X158 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X159 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X160 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X161 a_94942_n4187# CM_p_net_0.IN CM_p_net_0.OUT5 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X162 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X163 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X164 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X165 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X166 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X167 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X168 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X169 a_51954_n9018# CM_n_net_0.IN a_51394_n9018# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X170 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X171 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X172 a_31935_11461# a_29999_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X173 a_54076_11461# a_53676_10235# PRbiased_net_x5_1.IBP2 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X174 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X175 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X176 a_47666_10295# a_47838_4268# a_49642_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X177 a_108033_n22063# CM_p_net_1.IN a_107465_n22063# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X178 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X179 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X180 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X181 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X182 a_71318_n10715# CM_input_0.ISBCS a_75637_n16769# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X183 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X184 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X185 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X186 a_109439_n8593# CM_p_net_1.IN a_108601_n5878# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X187 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X188 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X189 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X190 CM_n_net_1.VSS a_71343_n40268# a_71743_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X191 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X192 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X193 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X194 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X195 a_112928_n31143# a_112406_n33067# a_112406_n33067# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X196 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X197 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X198 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X199 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X200 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X201 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X202 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X203 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X204 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X205 a_49960_n10812# CM_n_net_0.IN a_49438_n10812# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X206 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X207 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X208 CM_p_net_1.VDD CM_p_net_1.IN a_108601_n22968# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X209 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X210 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X211 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X212 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X213 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X214 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X215 a_92056_n20372# CM_p_net_0.IN a_91218_n17657# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X216 a_96348_n5997# CM_p_net_0.IN a_95780_n5997# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X217 a_106627_n22063# CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X218 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X219 CM_n_net_1.VSS a_59405_4328# a_59927_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X220 a_112325_n5878# CM_p_net_1.IN a_111795_n5878# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X221 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X222 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X223 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X224 a_65360_n5430# CM_n_net_0.IN a_64838_n5430# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X225 a_1808_n21432# a_n7408_n26036# a_1278_n21432# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X226 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X227 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X228 a_84952_n8712# CM_p_net_0.IN a_84384_n8712# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X229 a_36009_n40268# a_41738_n33067# a_43664_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X230 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X231 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X232 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X233 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X234 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X235 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X236 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X237 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X238 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X239 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X240 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X241 a_84952_n16752# CM_p_net_0.IN a_84384_n16752# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X242 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X243 a_37555_n5302# CM_n_net_1.IN a_37033_n5302# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X244 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X245 a_95290_10295# a_83172_4268# a_94739_4328# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X246 a_33283_n8890# CM_n_net_1.IN a_32723_n7993# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X247 a_102903_n21158# CM_p_net_1.IN a_102335_n21158# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X248 FC_top_0.AVDD FC_top_0.IREF a_n7828_n20082# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X249 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X250 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X251 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X252 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X253 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X254 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X255 a_51394_n4533# CM_n_net_0.IN a_50872_n5430# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X256 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X257 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X258 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X259 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X260 a_39549_n6199# CM_n_net_1.IN a_38989_n5302# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X261 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X262 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X263 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X264 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X265 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X266 a_53388_n4533# CM_n_net_0.IN a_52828_n4533# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X267 a_63052_n5430# CM_n_net_0.IN a_62492_n4533# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X268 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X269 a_67269_n39042# a_65333_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X270 a_9305_n11560# a_n7828_n21089# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X271 a_32723_n4405# CM_n_net_1.IN a_32201_n5302# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X272 a_62492_n16095# CM_n_net_0.IN a_61970_n16992# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X273 a_58220_n19683# CM_n_net_0.IN a_57660_n19683# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X274 a_83546_n3282# CM_p_net_0.IN a_83016_n6902# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X275 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X276 a_115137_n19348# CM_p_net_1.IN a_114607_n18443# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X277 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X278 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X279 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X280 a_49602_10295# a_47666_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X281 a_83546_n16752# CM_p_net_0.IN a_83016_n17657# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X282 a_103741_n8593# CM_p_net_1.IN a_102903_n5878# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X283 PRbiased_net_x5_0.VDD a_29999_n39042# a_30529_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X284 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X285 a_71343_n40268# a_77072_n33067# a_78998_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X286 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X287 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X288 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X289 a_83000_10295# a_83172_4268# a_84976_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X290 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X291 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X292 a_n10081_n11560# a_n7828_n21089# a_9305_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X293 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X294 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X295 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X296 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X297 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X298 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X299 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X300 a_73149_12227# a_71343_10235# CM_n_net_1.VSS PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X301 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X302 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X303 a_101239_4328# a_100839_4268# a_100667_10295# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X304 a_91218_n5092# CM_p_net_0.IN a_90650_n5092# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X305 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X306 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X307 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X308 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X309 a_96665_5486# a_94739_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X310 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X311 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X312 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X313 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X314 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X315 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X316 a_92056_n22182# CM_p_net_0.IN a_91218_n21277# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X317 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X318 a_53388_n16992# CM_n_net_0.IN a_52828_n16992# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X319 a_n7828_n21089# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X320 a_97754_n19467# CM_p_net_0.IN CM_p_net_0.OUT12 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X321 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X322 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X323 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X324 a_67309_4328# PRbiased_net_x5_1.IBN3 PRbiased_net_x5_1.ITN3 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X325 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X326 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X327 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X328 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X329 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X330 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X331 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X332 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X333 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X334 a_52828_n14301# CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X335 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X336 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X337 a_36681_n9787# CM_n_net_1.IN a_36121_n8890# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X338 a_35855_4328# a_29999_11461# a_37781_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X339 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X340 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X341 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X342 a_100929_n4973# CM_p_net_1.IN a_100399_n5878# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X343 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X344 a_89244_n7807# CM_p_net_0.IN a_88714_n11427# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X345 a_84952_n20372# CM_p_net_0.IN a_84384_n20372# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X346 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X347 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X348 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X349 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X350 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X351 a_107465_n8593# CM_p_net_1.IN a_106627_n8593# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X352 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X353 a_89244_n5997# CM_p_net_0.IN a_88714_n5997# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X354 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X355 a_56786_n5430# CM_n_net_0.IN a_56226_n5430# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X356 a_55482_n40208# a_53676_n40268# a_53522_n31143# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X357 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X358 a_83572_5486# PRbiased_net_x5_1.IBN4 a_83000_11461# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X359 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X360 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X361 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X362 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X363 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X364 CM_n_net_1.VSS a_106677_10235# a_107077_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X365 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X366 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X367 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X368 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X369 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X370 a_32723_n19555# CM_n_net_1.IN a_32201_n20452# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X371 a_53676_n40268# a_59405_n33067# a_61331_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X372 a_115137_n22063# CM_p_net_1.IN a_114299_n22063# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X373 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X374 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X375 a_59956_n40208# PRbiased_net_x5_0.IBP2 a_53676_n40268# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X376 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X377 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X378 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X379 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X380 a_102903_n16633# CM_p_net_1.IN a_102335_n16633# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X381 a_83546_n20372# CM_p_net_0.IN a_83016_n21277# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X382 a_56226_n14301# CM_n_net_0.IN a_55704_n15198# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X383 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X384 a_94942_n3282# CM_p_net_0.IN a_94412_n6902# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X385 a_49960_n16992# CM_n_net_0.IN a_49438_n16992# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X386 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X387 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X388 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X389 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X390 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X391 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X392 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X393 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X394 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X395 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X396 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X397 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X398 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X399 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X400 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X401 CM_p_net_0.VDD CM_p_net_0.IN a_96916_n23087# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X402 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X403 a_109439_n4973# CM_p_net_1.IN a_108601_n4973# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X404 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X405 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X406 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X407 a_85520_n17657# CM_p_net_0.IN a_84952_n17657# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X408 a_83172_4268# a_83000_11461# a_89378_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X409 CM_n_net_1.VSS a_n7828_n20082# a_n7408_n26036# CM_n_net_1.VSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X410 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X411 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X412 a_36121_n19555# CM_n_net_1.IN a_35599_n19555# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X413 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X414 a_71343_n40268# a_77072_n33067# a_78998_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X415 a_71343_10235# PRbiased_net_x5_1.IBP3 a_79029_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X416 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X417 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X418 a_51394_n15198# CM_n_net_0.IN a_50872_n16095# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X419 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X420 a_73149_n39042# a_71343_n40268# CM_n_net_1.VSS PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X421 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X422 PRbiased_net_x5_1.ITP1 a_30171_4268# a_42289_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X423 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X424 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X425 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X426 a_92056_n16752# CM_p_net_0.IN a_91218_n16752# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X427 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X428 a_112325_n4973# CM_p_net_1.IN a_111795_n5878# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X429 PRbiased_net_x5_1.VDD a_65333_11461# a_73115_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X430 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X431 a_47838_n33199# a_47666_n40208# a_54044_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X432 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X433 a_30415_n21349# CM_n_net_1.IN a_29855_n21349# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X434 a_30415_n18658# CM_n_net_1.IN a_29855_n18658# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X435 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X436 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X437 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X438 a_113163_n17538# CM_p_net_1.IN a_112325_n17538# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X439 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X440 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X441 a_102335_n9498# CM_p_net_1.IN a_101767_n9498# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X442 a_114363_10295# PRbiased_net_x5_1.IBP5 PRbiased_net_x5_1.ITP5 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X443 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X444 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X445 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X446 a_42387_n4405# CM_n_net_1.IN a_41865_n4405# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X447 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X448 a_29855_n19555# CM_n_net_1.IN a_29333_n19555# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X449 PRbiased_net_x5_1.IBN5 a_100667_11461# a_107045_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X450 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X451 PRbiased_net_x5_1.ITN2 PRbiased_net_x5_1.IBN2 a_48238_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X452 a_102903_n20253# CM_p_net_1.IN a_102335_n20253# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X453 a_102903_n4068# CM_p_net_1.IN a_102335_n4068# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X454 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X455 a_65920_n9018# CM_n_net_0.IN a_65360_n9018# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X456 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X457 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X458 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X459 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X460 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X461 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X462 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X463 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X464 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X465 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X466 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X467 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X468 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X469 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X470 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X471 CM_n_net_1.VSS CM_input_0.ISBCS a_72655_n15993# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X472 a_109439_n19348# CM_p_net_1.IN CM_p_net_1.OUT10 CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X473 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X474 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X475 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X476 a_30415_n10684# CM_n_net_1.IN a_29855_n10684# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X477 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X478 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X479 a_44381_n5302# CM_n_net_1.IN a_43821_n5302# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X480 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X481 a_53676_10235# a_59405_4328# a_61331_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X482 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X483 a_103741_n4973# CM_p_net_1.IN a_102903_n4973# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X484 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X485 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X486 a_53676_n40268# a_59405_n33067# a_61331_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X487 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X488 a_85520_n21277# CM_p_net_0.IN a_84952_n21277# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X489 PRbiased_net_x5_1.ITP5 PRbiased_net_x5_1.IBP5 a_112957_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X490 CM_n_net_1.VSS a_59405_4328# a_59927_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X491 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X492 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X493 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X494 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X495 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X496 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X497 a_36121_n8890# CM_n_net_1.IN a_35599_n8890# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X498 a_90082_n9617# CM_p_net_0.IN a_89244_n9617# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X499 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X500 a_92056_n20372# CM_p_net_0.IN a_91218_n20372# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X501 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X502 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X503 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X504 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X505 a_38115_n8890# CM_n_net_1.IN a_37555_n8890# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X506 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X507 a_97754_n19467# CM_p_net_0.IN a_97224_n18562# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X508 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X509 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X510 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X511 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X512 a_56226_n5430# CM_n_net_0.IN a_55704_n6327# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X513 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X514 PRbiased_net_x5_1.ITP5 PRbiased_net_x5_1.IBP5 a_112957_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X515 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X516 a_65920_n21477# CM_n_net_0.IN a_65360_n21477# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X517 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X518 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X519 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X520 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X521 a_65920_n19683# CM_n_net_0.IN a_65360_n18786# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X522 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X523 a_113163_n21158# CM_p_net_1.IN a_112325_n21158# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X524 a_65360_n4533# CM_n_net_0.IN a_64838_n5430# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X525 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X526 a_89244_n7807# CM_p_net_0.IN a_88714_n6902# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X527 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X528 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X529 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X530 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X531 a_62492_n7224# CM_n_net_0.IN CM_n_net_0.OUT6 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X532 a_95780_n5092# CM_p_net_0.IN a_94942_n5092# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X533 a_108601_n22063# CM_p_net_1.IN a_108033_n22063# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X534 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X535 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X536 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X537 a_55448_n33067# a_47666_n40208# PRbiased_net_x5_0.IBN2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X538 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X539 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X540 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X541 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X542 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X543 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X544 PRbiased_net_x5_0.IBN2 a_47666_n40208# a_54044_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X545 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X546 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X547 a_83000_10295# a_83172_4268# a_84976_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X548 a_88880_13393# a_89010_10235# a_90816_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X549 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X550 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X551 a_59654_n21477# CM_n_net_0.IN a_59094_n21477# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X552 a_108483_10295# a_106677_10235# a_106523_7410# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X553 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X554 a_59654_n19683# CM_n_net_0.IN a_59094_n18786# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X555 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X556 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X557 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X558 FC_top_0.AVDD FC_top_0.IREF a_n7828_n21089# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X559 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X560 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X561 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X562 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X563 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X564 a_96665_7410# a_94739_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X565 a_42947_n7096# CM_n_net_1.IN a_42387_n7096# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X566 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X567 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X568 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X569 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X570 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X571 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X572 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X573 a_65333_11461# a_65333_10295# a_67269_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X574 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X575 a_88856_4328# a_89010_10235# a_89410_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X576 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X577 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X578 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X579 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X580 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X581 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X582 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X583 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X584 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X585 a_97754_n22182# CM_p_net_0.IN a_96916_n22182# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X586 a_59094_n5430# CM_n_net_0.IN a_58572_n5430# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X587 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X588 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X589 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X590 a_85520_n16752# CM_p_net_0.IN a_84952_n16752# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X591 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X592 a_n7828_n21089# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X593 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X594 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X595 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X596 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X597 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X598 a_83572_7410# PRbiased_net_x5_1.IBN4 a_83000_11461# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X599 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X600 a_65863_n37110# a_65333_n39042# a_65333_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X601 a_101197_13393# a_100667_10295# a_100667_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X602 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X603 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X604 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X605 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X606 a_43695_10295# PRbiased_net_x5_1.IBP1 PRbiased_net_x5_1.ITP1 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X607 a_36681_n7993# CM_n_net_1.IN a_36121_n7993# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X608 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X609 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X610 a_65333_n40208# a_65333_n39042# a_67269_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X611 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X612 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X613 a_n10081_n10574# a_n7828_n21089# FC_top_0.VOUT CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X614 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X615 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X616 a_n10081_n10574# a_n7828_n21089# FC_top_0.VOUT CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X617 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X618 a_56786_n5430# CM_n_net_0.IN a_56226_n4533# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X619 a_113163_n16633# CM_p_net_1.IN a_112325_n16633# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X620 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X621 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X622 a_102335_n8593# CM_p_net_1.IN a_101767_n8593# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X623 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X624 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X625 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X626 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X627 a_101197_11461# a_100667_10295# a_100667_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X628 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X629 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X630 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X631 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X632 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X633 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X634 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X635 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X636 a_102903_n3163# CM_p_net_1.IN a_102335_n3163# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X637 a_43821_n21349# CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X638 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X639 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X640 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X641 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X642 a_51954_n4533# CM_n_net_0.IN a_51394_n3636# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X643 a_108449_5486# a_100667_11461# PRbiased_net_x5_1.IBN5 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X644 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X645 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X646 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X647 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X648 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X649 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X650 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X651 a_55448_n31143# a_47666_n40208# a_47838_n33199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X652 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X653 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X654 a_109439_n19348# CM_p_net_1.IN a_108909_n18443# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X655 a_95780_n17657# CM_p_net_0.IN a_94942_n17657# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X656 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X657 a_84384_n5997# CM_p_net_0.IN a_83546_n5997# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X658 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X659 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X660 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X661 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X662 a_101767_n11308# CM_p_net_1.IN a_100929_n11308# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X663 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X664 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X665 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X666 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X667 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X668 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X669 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X670 a_85520_n20372# CM_p_net_0.IN a_84952_n20372# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X671 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X672 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X673 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X674 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X675 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X676 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X677 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X678 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X679 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X680 a_37555_n21349# CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X681 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X682 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X683 a_43821_n10684# CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X684 a_71189_4328# a_65333_11461# a_73115_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X685 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X686 a_59927_n34225# a_59405_n33067# a_53676_n40268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X687 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X688 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X689 a_30571_n34225# PRbiased_net_x5_0.IBN1 a_29999_n40208# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X690 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X691 a_50520_n16095# CM_n_net_0.IN a_49960_n16095# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X692 a_90082_n8712# CM_p_net_0.IN a_89244_n8712# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X693 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X694 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X695 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X696 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X697 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X698 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X699 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X700 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X701 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X702 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X703 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X704 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X705 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X706 a_1808_n22743# a_n7408_n26036# a_1278_n22743# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X707 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X708 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X709 PRbiased_net_x5_1.ITN2 PRbiased_net_x5_1.IBN2 a_48238_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X710 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X711 a_113163_n20253# CM_p_net_1.IN a_112325_n20253# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X712 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X713 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X714 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X715 a_30415_n20452# CM_n_net_1.IN a_29855_n20452# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X716 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X717 a_30415_n17761# CM_n_net_1.IN a_29855_n17761# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X718 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X719 a_89378_n33067# a_83000_n40208# PRbiased_net_x5_0.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X720 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X721 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X722 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X723 a_42387_n15967# CM_n_net_1.IN a_41865_n16864# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X724 a_37555_n10684# CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X725 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X726 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X727 a_84976_6252# PRbiased_net_x5_1.IBN4 PRbiased_net_x5_1.ITN4 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X728 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X729 a_101767_n15728# CM_p_net_1.IN a_100929_n15728# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X730 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X731 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X732 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X733 a_84936_n40208# a_83000_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X734 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X735 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X736 a_89244_n11427# CM_p_net_0.IN a_88714_n11427# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X737 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X738 a_36681_n15967# CM_n_net_1.IN a_36121_n15967# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X739 a_n2230_n25929# a_n7828_n21089# a_n2752_n26552# CM_n_net_1.VSS nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X740 PRbiased_net_x5_1.ITP3 a_65505_4268# a_77623_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X741 PRbiased_net_x5_1.IBP2 a_53676_10235# a_55482_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X742 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X743 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X744 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X745 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X746 a_65920_n9018# CM_n_net_0.IN a_65360_n8121# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X747 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X748 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X749 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X750 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X751 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X752 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X753 a_71743_n37110# a_71343_n40268# a_53546_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X754 a_109439_n22063# CM_p_net_1.IN a_108601_n22063# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X755 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X756 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X757 a_95780_n21277# CM_p_net_0.IN a_94942_n21277# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X758 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X759 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X760 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X761 a_96348_n5092# CM_p_net_0.IN a_95780_n5092# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X762 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X763 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X764 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X765 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X766 PRbiased_net_x5_0.IBP3 a_71343_n40268# a_73149_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X767 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X768 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X769 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X770 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X771 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X772 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X773 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X774 a_49642_4328# PRbiased_net_x5_1.IBN2 PRbiased_net_x5_1.ITN2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X775 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X776 a_42260_n34225# a_41738_n33067# a_36009_n40268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X777 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X778 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X779 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X780 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X781 a_108483_n39042# a_106677_n40268# CM_n_net_1.VSS PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X782 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X783 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X784 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X785 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X786 a_64486_n15198# CM_n_net_0.IN a_63926_n14301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X787 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X788 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X789 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X790 a_58220_n15198# CM_n_net_0.IN a_57660_n15198# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X791 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X792 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X793 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X794 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X795 a_113731_n17538# CM_p_net_1.IN a_113163_n17538# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X796 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X797 a_36121_n7993# CM_n_net_1.IN a_35599_n8890# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X798 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X799 a_89378_5486# a_83000_11461# PRbiased_net_x5_1.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X800 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X801 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X802 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X803 a_115137_n4973# CM_p_net_1.IN a_114299_n4068# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X804 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X805 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X806 a_31935_10295# a_29999_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X807 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X808 a_54076_10295# a_53676_10235# a_35879_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X809 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X810 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X811 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X812 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X813 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X814 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X815 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X816 a_56226_n4533# CM_n_net_0.IN a_55704_n4533# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X817 a_88856_7410# a_83000_11461# a_90782_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X818 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X819 a_57660_n9018# CM_n_net_0.IN a_57138_n9915# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X820 a_89244_n15847# CM_p_net_0.IN CM_p_net_0.OUT9 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X821 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X822 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X823 a_59927_n32301# a_59405_n33067# a_53676_n40268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X824 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X825 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X826 a_59654_n9018# CM_n_net_0.IN a_59094_n9018# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X827 a_30571_n32301# PRbiased_net_x5_0.IBN1 a_29999_n40208# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X828 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X829 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X830 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X831 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X832 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X833 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X834 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X835 a_45255_n7096# CM_n_net_1.IN a_44381_n5302# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X836 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X837 a_101197_n38276# a_100667_n39042# a_100667_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X838 a_107465_n17538# CM_p_net_1.IN a_106627_n17538# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X839 a_31289_n3508# CM_n_net_1.IN a_30415_n7096# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X840 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X841 a_30415_n9787# CM_n_net_1.IN a_29855_n9787# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X842 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X843 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X844 a_112928_4328# a_112406_4328# a_112406_4328# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X845 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X846 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X847 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X848 CM_n_net_1.OUT5 CM_n_net_1.IN a_42387_n3508# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X849 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X850 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X851 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X852 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X853 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X854 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X855 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X856 a_89378_n31143# a_83000_n40208# a_88856_n31143# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X857 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X858 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X859 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X860 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X861 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X862 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X863 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X864 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X865 a_33283_n4405# CM_n_net_1.IN a_32723_n4405# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X866 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X867 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X868 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X869 a_29855_n8890# CM_n_net_1.IN a_29333_n8890# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X870 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X871 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X872 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X873 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X874 a_90650_n11427# CM_p_net_0.IN a_90082_n11427# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X875 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X876 a_95780_n16752# CM_p_net_0.IN a_94942_n16752# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X877 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X878 a_50520_n7224# CM_n_net_0.IN a_49960_n7224# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X879 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X880 a_101767_n10403# CM_p_net_1.IN a_100929_n10403# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X881 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X882 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X883 a_113731_n21158# CM_p_net_1.IN a_113163_n21158# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X884 a_32723_n15070# CM_n_net_1.IN a_32201_n15967# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X885 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X886 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X887 a_89244_n5092# CM_p_net_0.IN a_88714_n5997# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X888 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X889 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X890 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X891 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X892 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X893 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X894 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X895 a_59405_4328# a_47838_4268# a_61362_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X896 a_90816_n40208# a_89010_n40268# a_88856_n31143# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X897 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X898 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X899 CM_n_net_1.VSS a_89010_n40268# a_89410_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X900 a_72655_n16769# CM_input_0.ISBCS CM_input_0.IP2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X901 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X902 a_59094_n4533# CM_n_net_0.IN a_58572_n5430# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X903 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X904 a_42260_n32301# a_41738_n33067# a_36009_n40268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X905 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X906 a_47666_11461# PRbiased_net_x5_1.IBN2 a_49642_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X907 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X908 a_51954_n21477# CM_n_net_0.IN a_51394_n20580# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X909 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X910 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X911 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X912 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X913 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X914 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X915 a_49960_n6327# CM_n_net_0.IN a_49438_n6327# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X916 a_65905_4328# a_65505_4268# a_65333_10295# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X917 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X918 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X919 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X920 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X921 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X922 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X923 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X924 a_59405_4328# a_47838_4268# a_61362_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X925 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X926 a_37781_4328# a_29999_11461# a_30171_4268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X927 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X928 a_108033_n4068# CM_p_net_1.IN a_107465_n4068# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X929 a_107465_n21158# CM_p_net_1.IN a_106627_n21158# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X930 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X931 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X932 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X933 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X934 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X935 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X936 a_96348_n11427# CM_p_net_0.IN a_95780_n11427# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X937 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X938 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X939 a_36121_n15070# CM_n_net_1.IN a_35599_n15070# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X940 a_108449_7410# a_100667_11461# a_100839_4268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X941 a_65920_n4533# CM_n_net_0.IN a_65360_n3636# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X942 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X943 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X944 a_90650_n15847# CM_p_net_0.IN a_90082_n15847# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X945 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X946 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X947 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X948 a_101767_n14823# CM_p_net_1.IN a_100929_n14823# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X949 a_77594_n34225# a_77072_n33067# a_71343_n40268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X950 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X951 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X952 a_43821_n20452# CM_n_net_1.IN a_43299_n20452# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X953 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X954 a_89244_n10522# CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X955 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X956 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X957 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X958 a_30171_n33199# a_29999_n40208# a_36377_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X959 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X960 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X961 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X962 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X963 a_33283_n21349# CM_n_net_1.IN a_32723_n21349# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X964 a_33283_n19555# CM_n_net_1.IN a_32723_n18658# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X965 FC_top_0.AVDD FC_top_0.IREF a_n7828_n21089# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X966 a_95780_n20372# CM_p_net_0.IN a_94942_n20372# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X967 a_57660_n16095# CM_n_net_0.IN a_57138_n16095# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X968 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X969 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X970 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X971 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X972 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X973 a_29855_n15070# CM_n_net_1.IN a_29333_n15070# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X974 a_9305_n11560# a_n7828_n21089# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X975 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X976 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X977 PRbiased_net_x5_0.VDD a_65333_n39042# a_65863_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X978 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X979 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X980 a_9305_n11560# a_n7828_n21089# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X981 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X982 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X983 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X984 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X985 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X986 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X987 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X988 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X989 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X990 a_95290_n37110# a_83172_n33199# a_94739_n33067# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X991 a_53522_7410# a_47666_11461# a_55448_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X992 a_37555_n20452# CM_n_net_1.IN a_37033_n20452# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X993 a_96348_n15847# CM_p_net_0.IN a_95780_n15847# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X994 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X995 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X996 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X997 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X998 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X999 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1000 a_113731_n16633# CM_p_net_1.IN a_113163_n16633# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1001 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1002 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1003 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1004 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1005 CM_p_net_1.VDD CM_p_net_1.IN a_102903_n11308# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1006 a_89010_n40268# PRbiased_net_x5_0.IBP4 a_96696_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1007 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1008 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1009 a_114607_n6783# CM_p_net_1.IN a_114299_n3163# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1010 a_33283_n10684# CM_n_net_1.IN a_32723_n10684# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1011 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1012 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1013 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1014 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1015 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1016 a_43695_n40208# a_30171_n33199# PRbiased_net_x5_0.ITP1 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1017 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1018 a_89410_12227# a_89010_10235# PRbiased_net_x5_1.IBP4 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1019 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1020 a_89244_n14942# CM_p_net_0.IN a_88714_n18562# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1021 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1022 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1023 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1024 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1025 a_31935_n37110# a_29999_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1026 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1027 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1028 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1029 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1030 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1031 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1032 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1033 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1034 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1035 PRbiased_net_x5_0.ITP4 a_83172_n33199# a_95290_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1036 a_107465_n16633# CM_p_net_1.IN a_106627_n16633# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1037 PRbiased_net_x5_1.VDD a_29999_11461# a_37781_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1038 a_51954_n10812# CM_n_net_0.IN a_51394_n10812# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1039 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1040 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1041 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1042 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1043 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1044 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1045 a_48196_13393# a_47666_10295# a_47666_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1046 a_54044_4328# a_47666_11461# a_53522_4328# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1047 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1048 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1049 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1050 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1051 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1052 a_30529_n37110# a_29999_n39042# a_29999_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1053 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1054 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1055 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1056 a_103741_n16633# CM_p_net_1.IN a_102903_n15728# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1057 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1058 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1059 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1060 a_89378_7410# a_83000_11461# a_88856_7410# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1061 a_71189_7410# a_71343_10235# a_71743_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1062 a_77594_n32301# a_77072_n33067# a_71343_n40268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1063 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1064 a_45815_n16864# CM_n_net_1.IN a_45255_n15967# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1065 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1066 a_90650_n10522# CM_p_net_0.IN a_90082_n10522# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1067 a_48196_11461# a_47666_10295# a_47666_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1068 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1069 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1070 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1071 a_n7828_n21089# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1072 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X1073 PRbiased_net_x5_0.IBN1 a_29999_n40208# a_36377_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1074 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1075 a_113731_n20253# CM_p_net_1.IN a_113163_n20253# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1076 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1077 a_112406_n33067# a_112406_n33067# a_114332_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1078 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1079 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1080 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1081 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1082 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1083 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1084 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1085 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1086 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1087 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1088 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1089 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1090 CM_n_net_1.VSS a_71343_10235# a_71743_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1091 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1092 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1093 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1094 a_32723_n9787# CM_n_net_1.IN a_32201_n9787# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1095 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1096 a_83000_n39042# a_83000_n39042# a_84936_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1097 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1098 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1099 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1100 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1101 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1102 a_45255_n3508# CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1103 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1104 a_39549_n16864# CM_n_net_1.IN a_38989_n15967# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1105 a_52828_n6327# CM_n_net_0.IN a_52306_n8121# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1106 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1107 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1108 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1109 a_83530_n38276# a_83000_n39042# a_83000_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1110 a_108033_n3163# CM_p_net_1.IN a_107465_n3163# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1111 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1112 a_107465_n20253# CM_p_net_1.IN a_106627_n20253# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1113 a_59654_n9018# CM_n_net_0.IN a_59094_n8121# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1114 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1115 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1116 a_65360_n20580# CM_n_net_0.IN a_64838_n20580# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1117 a_96348_n10522# CM_p_net_0.IN a_95780_n10522# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1118 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1119 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1120 a_65360_n17889# CM_n_net_0.IN a_64486_n16095# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1121 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1122 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1123 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1124 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1125 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1126 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1127 PRbiased_net_x5_1.ITP5 a_100839_4268# a_112957_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1128 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1129 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1130 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1131 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1132 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1133 a_90650_n14942# CM_p_net_0.IN a_90082_n14942# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1134 a_48196_n37110# a_47666_n39042# a_47666_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1135 PRbiased_net_x5_0.IBN2 a_47666_n40208# a_54044_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1136 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1137 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1138 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1139 a_52828_n19683# CM_n_net_0.IN a_52306_n20580# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1140 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1141 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1142 a_n7828_n20082# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1143 a_100667_n39042# a_100667_n39042# a_102603_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1144 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1145 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1146 a_90650_n9617# CM_p_net_0.IN a_90082_n9617# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1147 a_59094_n20580# CM_n_net_0.IN a_58572_n20580# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1148 a_29855_n7993# CM_n_net_1.IN a_29333_n8890# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1149 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1150 a_59094_n17889# CM_n_net_0.IN a_58220_n16095# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1151 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1152 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1153 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1154 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1155 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1156 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1157 a_32723_n14173# CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1158 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1159 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1160 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1161 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1162 a_67269_12227# a_65333_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1163 PRbiased_net_x5_1.VDD a_65333_10295# a_65863_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1164 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1165 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1166 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1167 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1168 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1169 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1170 a_102335_n22968# CM_p_net_1.IN a_101767_n22968# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1171 PRbiased_net_x5_0.VDD a_100667_n39042# a_101197_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1172 a_96348_n14942# CM_p_net_0.IN a_95780_n14942# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1173 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1174 a_56226_n19683# CM_n_net_0.IN a_55704_n19683# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1175 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1176 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1177 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1178 a_71189_n34225# a_71343_n40268# a_71743_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1179 a_103741_n10403# CM_p_net_1.IN a_102903_n10403# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1180 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1181 a_38989_n7096# CM_n_net_1.IN a_38115_n5302# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1182 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1183 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1184 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1185 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1186 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1187 a_112406_n33067# a_112406_n33067# a_114332_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1188 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1189 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1190 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1191 CM_n_net_1.VSS a_59405_4328# a_59927_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1192 a_100667_11461# a_100667_10295# a_102603_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1193 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1194 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1195 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1196 PRbiased_net_x5_1.VDD a_65333_10295# a_65863_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1197 a_84384_n5092# CM_p_net_0.IN a_83546_n5092# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1198 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1199 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1200 a_61331_n34225# a_59405_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1201 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1202 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1203 a_36121_n14173# CM_n_net_1.IN a_35599_n15070# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1204 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1205 a_100929_n22968# CM_p_net_1.IN a_100399_n22968# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1206 a_n1670_n25929# a_n7828_n21089# a_n2230_n25376# CM_n_net_1.VSS nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X1207 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1208 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1209 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1210 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1211 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1212 a_101239_5486# PRbiased_net_x5_1.IBN5 a_100667_11461# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1213 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1214 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1215 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1216 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1217 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1218 a_45815_n6199# CM_n_net_1.IN a_45255_n6199# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1219 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1220 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1221 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1222 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1223 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1224 a_114299_n5878# CM_p_net_1.IN a_113731_n5878# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1225 a_36681_n5302# CM_n_net_1.IN a_36121_n4405# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1226 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1227 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1228 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1229 a_67309_5486# a_65505_4268# PRbiased_net_x5_1.ITN3 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1230 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1231 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1232 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1233 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1234 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1235 a_33283_n21349# CM_n_net_1.IN a_32723_n20452# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1236 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1237 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1238 a_31849_n19555# CM_n_net_1.IN a_32723_n17761# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1239 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1240 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1241 a_101197_10295# a_100667_10295# a_100667_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1242 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1243 a_29855_n14173# CM_n_net_1.IN a_29333_n15070# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1244 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1245 a_103211_n18443# CM_p_net_1.IN a_102903_n14823# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1246 a_65360_n10812# CM_n_net_0.IN a_63052_n10812# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1247 PRbiased_net_x5_0.VDD a_29999_n39042# a_30529_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1248 a_108449_n34225# a_100667_n40208# a_100839_n33199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1249 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1250 a_47838_n33199# a_47666_n40208# a_54044_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1251 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1252 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1253 a_42387_n9787# CM_n_net_1.IN a_41865_n10684# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1254 a_67269_n40208# a_65333_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1255 a_83000_11461# PRbiased_net_x5_1.IBN4 a_84976_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1256 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1257 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1258 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1259 a_31849_n19555# CM_n_net_1.IN a_31289_n19555# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1260 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1261 a_96916_n11427# CM_p_net_0.IN a_96348_n11427# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1262 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1263 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1264 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1265 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1266 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1267 a_96665_6252# a_94739_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1268 a_54076_n37110# a_53676_n40268# a_35879_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1269 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1270 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1271 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1272 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1273 a_57660_n3636# CM_n_net_0.IN a_56786_n7224# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1274 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1275 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1276 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1277 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1278 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1279 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1280 a_59654_n4533# CM_n_net_0.IN a_59094_n3636# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1281 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1282 CM_n_net_1.VSS a_36009_10235# a_36409_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1283 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1284 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1285 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1286 a_59094_n10812# CM_n_net_0.IN a_56786_n10812# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1287 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1288 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1289 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1290 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1291 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1292 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1293 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1294 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1295 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1296 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1297 a_79029_n37110# PRbiased_net_x5_0.IBP3 PRbiased_net_x5_0.ITP3 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1298 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1299 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1300 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1301 a_73149_13393# a_71343_10235# a_71189_4328# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1302 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1303 a_83000_11461# a_83000_10295# a_84936_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1304 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1305 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1306 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1307 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1308 a_83572_6252# a_83172_4268# a_83000_10295# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1309 PRbiased_net_x5_1.IBN4 a_83000_11461# a_89378_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1310 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1311 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1312 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1313 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1314 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1315 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1316 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1317 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1318 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1319 a_61331_n32301# a_59405_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1320 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1321 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1322 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1323 a_96916_n15847# CM_p_net_0.IN a_96348_n15847# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1324 a_73149_11461# a_71343_10235# CM_n_net_1.VSS PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1325 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1326 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1327 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1328 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1329 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1330 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1331 a_83546_n7807# CM_p_net_0.IN a_83016_n11427# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1332 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1333 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1334 a_90650_n8712# CM_p_net_0.IN a_90082_n8712# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1335 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1336 a_n10081_n10574# a_n7828_n21089# FC_top_0.VOUT CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1337 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1338 a_83546_n5997# CM_p_net_0.IN a_83016_n5997# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1339 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1340 a_62492_n20580# CM_n_net_0.IN a_61970_n21477# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1341 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1342 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1343 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1344 a_62492_n17889# CM_n_net_0.IN CM_n_net_0.OUT12 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1345 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1346 a_29999_n40208# a_29999_n39042# a_31935_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1347 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1348 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1349 a_106523_7410# a_106677_10235# a_107077_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1350 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1351 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1352 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1353 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1354 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1355 CM_n_net_1.VSS a_77072_4328# a_77594_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1356 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1357 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1358 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1359 a_91218_n9617# CM_p_net_0.IN a_90650_n9617# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1360 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1361 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1362 a_96665_n34225# a_94739_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1363 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1364 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1365 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1366 a_108449_n32301# a_100667_n40208# PRbiased_net_x5_0.IBN5 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1367 a_61362_n37110# PRbiased_net_x5_0.IBP2 PRbiased_net_x5_0.ITP2 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1368 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1369 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1370 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1371 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1372 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1373 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1374 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1375 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1376 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1377 a_53522_n31143# a_47666_n40208# a_55448_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1378 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1379 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1380 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1381 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1382 CM_n_net_1.VSS a_106677_10235# a_107077_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1383 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1384 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1385 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1386 a_59405_4328# a_59405_4328# a_61331_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1387 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1388 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1389 a_84384_n23087# CM_p_net_0.IN a_83546_n23087# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1390 PRbiased_net_x5_1.VDD a_65333_11461# a_73115_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1391 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1392 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1393 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1394 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1395 a_59927_n33067# a_59405_n33067# a_59405_n33067# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1396 a_73149_n40208# a_71343_n40268# a_71189_n31143# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1397 a_36121_n4405# CM_n_net_1.IN a_35599_n4405# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1398 a_30571_n33067# a_30171_n33199# a_29999_n39042# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1399 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1400 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1401 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1402 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1403 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1404 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1405 a_65360_n16992# CM_n_net_0.IN a_64838_n18786# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1406 a_38115_n4405# CM_n_net_1.IN a_37555_n4405# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1407 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1408 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1409 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1410 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1411 a_65920_n15198# CM_n_net_0.IN a_65360_n14301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1412 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X1413 PRbiased_net_x5_1.ITN2 a_47838_4268# a_48238_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1414 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1415 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1416 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1417 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1418 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1419 a_114299_n4973# CM_p_net_1.IN a_113731_n4973# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1420 PRbiased_net_x5_1.ITP1 PRbiased_net_x5_1.IBP1 a_42289_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1421 a_63926_n21477# CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1422 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1423 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1424 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1425 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1426 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1427 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1428 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1429 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1430 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1431 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1432 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1433 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1434 a_94942_n7807# CM_p_net_0.IN a_94412_n11427# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1435 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1436 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1437 a_47666_n40208# a_47666_n39042# a_49602_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1438 a_94942_n5997# CM_p_net_0.IN a_94412_n5997# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1439 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1440 a_59094_n16992# CM_n_net_0.IN a_58572_n18786# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1441 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1442 CM_n_net_1.VSS a_n7828_n20082# a_n7408_n26036# CM_n_net_1.VSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X1443 PRbiased_net_x5_1.ITP1 PRbiased_net_x5_1.IBP1 a_42289_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1444 a_38989_n3508# CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1445 a_59654_n15198# CM_n_net_0.IN a_59094_n14301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1446 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1447 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1448 a_100929_n19348# CM_p_net_1.IN a_100399_n22968# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1449 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1450 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1451 a_96916_n10522# CM_p_net_0.IN a_96348_n10522# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1452 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1453 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1454 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1455 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1456 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1457 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1458 a_42260_n33067# a_41738_n33067# a_41738_n33067# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1459 FC_top_0.VOUT a_n7828_n21089# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1460 a_101239_7410# PRbiased_net_x5_1.IBN5 a_100667_11461# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1461 FC_top_0.VOUT a_n7828_n21089# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1462 PRbiased_net_x5_0.VDD a_47666_n39042# a_48196_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1463 a_45255_n19555# CM_n_net_1.IN a_44733_n20452# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1464 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1465 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1466 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1467 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1468 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1469 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1470 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1471 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1472 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1473 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1474 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1475 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1476 a_62492_n10812# CM_n_net_0.IN a_61970_n10812# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1477 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1478 a_96665_n32301# a_94739_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1479 a_67309_7410# a_65505_4268# PRbiased_net_x5_1.ITN3 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1480 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1481 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1482 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1483 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1484 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1485 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1486 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1487 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1488 PRbiased_net_x5_0.VDD a_47666_n40208# a_55448_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1489 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1490 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1491 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1492 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1493 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1494 a_53676_10235# PRbiased_net_x5_1.IBP2 a_61362_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1495 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1496 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1497 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1498 a_71743_12227# a_71343_10235# PRbiased_net_x5_1.IBP3 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1499 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1500 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1501 a_59927_n31143# a_59405_n33067# a_59405_n33067# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1502 a_38989_n19555# CM_n_net_1.IN a_38467_n20452# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1503 a_30571_n31143# a_30171_n33199# a_29999_n39042# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1504 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1505 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1506 a_102903_n22968# CM_p_net_1.IN a_102335_n22968# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1507 a_96916_n14942# CM_p_net_0.IN a_96348_n14942# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1508 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1509 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1510 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1511 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1512 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1513 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1514 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1515 a_96696_n37110# PRbiased_net_x5_0.IBP4 PRbiased_net_x5_0.ITP4 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1516 a_83546_n7807# CM_p_net_0.IN a_83016_n6902# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1517 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1518 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1519 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1520 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1521 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1522 a_42947_n21349# CM_n_net_1.IN a_42387_n21349# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1523 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1524 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1525 a_42947_n18658# CM_n_net_1.IN a_42387_n18658# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1526 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1527 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1528 a_47838_4268# a_47666_11461# a_54044_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1529 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1530 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1531 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1532 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1533 a_51954_n10812# CM_n_net_0.IN a_51394_n9915# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1534 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1535 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1536 a_91218_n8712# CM_p_net_0.IN a_90650_n8712# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1537 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1538 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1539 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1540 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1541 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1542 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1543 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1544 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1545 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1546 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1547 a_106627_n9498# CM_p_net_1.IN a_106097_n9498# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1548 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1549 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1550 a_83172_4268# a_83000_11461# a_89378_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1551 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1552 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1553 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1554 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1555 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1556 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1557 a_39549_n6199# CM_n_net_1.IN a_38989_n6199# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1558 a_53546_n40208# a_53676_n40268# a_55482_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1559 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1560 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1561 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1562 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1563 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1564 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1565 a_64486_n19683# CM_n_net_0.IN a_63926_n19683# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1566 a_84384_n22182# CM_p_net_0.IN a_83546_n22182# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1567 a_42947_n10684# CM_n_net_1.IN a_42387_n10684# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1568 a_42260_n31143# a_41738_n33067# a_41738_n33067# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1569 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1570 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1571 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1572 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1573 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1574 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1575 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1576 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1577 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1578 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1579 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1580 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1581 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1582 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1583 a_95780_n9617# CM_p_net_0.IN a_94942_n9617# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1584 a_65333_n39042# a_65333_n39042# a_67269_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1585 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1586 PRbiased_net_x5_0.ITN5 PRbiased_net_x5_0.IBN5 a_101239_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1587 a_n7828_n20082# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1588 a_47666_11461# a_47666_10295# a_49602_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1589 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1590 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1591 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1592 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1593 a_53522_n31143# a_53676_n40268# a_54076_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1594 a_65863_n38276# a_65333_n39042# a_65333_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1595 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1596 a_108449_6252# a_100667_11461# PRbiased_net_x5_1.IBN5 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1597 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1598 a_71189_n31143# a_65333_n40208# a_73115_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1599 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1600 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1601 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1602 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1603 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1604 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1605 a_94942_n7807# CM_p_net_0.IN a_94412_n6902# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1606 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1607 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1608 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1609 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1610 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1611 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1612 a_77594_n33067# a_77072_n33067# a_77072_n33067# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1613 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1614 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1615 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1616 a_31289_n8890# CM_n_net_1.IN a_30767_n9787# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1617 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1618 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1619 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1620 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1621 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1622 a_62492_n16992# CM_n_net_0.IN a_61970_n16992# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1623 a_52828_n15198# CM_n_net_0.IN a_52306_n16095# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1624 PRbiased_net_x5_0.IBN1 a_29999_n40208# a_36377_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1625 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1626 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1627 a_31975_n34225# a_30171_n33199# PRbiased_net_x5_0.ITN1 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1628 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X1629 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1630 a_42947_n9787# CM_n_net_1.IN a_42387_n8890# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1631 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1632 a_59405_4328# a_59405_4328# a_61331_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1633 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1634 a_100929_n19348# CM_p_net_1.IN a_100399_n18443# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1635 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1636 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1637 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1638 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1639 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1640 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1641 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1642 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1643 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1644 a_85520_n4187# CM_p_net_0.IN a_84952_n4187# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1645 a_48196_10295# a_47666_10295# a_47666_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1646 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1647 a_33283_n10684# CM_n_net_1.IN a_32723_n9787# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1648 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1649 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1650 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1651 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1652 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1653 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1654 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1655 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1656 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1657 a_49642_5486# a_47838_4268# PRbiased_net_x5_1.ITN2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1658 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1659 a_n10081_n11560# a_n7828_n21089# a_9305_n11560# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1660 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1661 a_53388_n6327# CM_n_net_0.IN a_52828_n6327# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1662 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1663 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1664 a_n10081_n11560# a_n7828_n21089# a_9305_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1665 a_63052_n8121# CM_n_net_0.IN a_62492_n6327# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1666 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1667 a_71189_4328# a_71343_10235# a_71743_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1668 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1669 a_56226_n15198# CM_n_net_0.IN a_55704_n15198# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1670 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1671 a_83546_n19467# CM_p_net_0.IN a_83016_n23087# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1672 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1673 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1674 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1675 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1676 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1677 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1678 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1679 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1680 a_112957_12227# a_100839_4268# a_112406_4328# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1681 a_102335_n22063# CM_p_net_1.IN a_101767_n22063# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1682 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1683 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1684 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1685 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1686 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1687 PRbiased_net_x5_1.VDD a_83000_11461# a_90782_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1688 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1689 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1690 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1691 a_102903_n5878# CM_p_net_1.IN a_102335_n5878# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1692 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1693 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1694 a_53388_n21477# CM_n_net_0.IN a_52828_n21477# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1695 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1696 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1697 a_53676_n40268# PRbiased_net_x5_0.IBP2 a_61362_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1698 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1699 a_53388_n19683# CM_n_net_0.IN a_52828_n18786# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1700 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1701 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1702 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1703 a_30415_n5302# CM_n_net_1.IN a_29855_n5302# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1704 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1705 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1706 PRbiased_net_x5_0.ITN5 PRbiased_net_x5_0.IBN5 a_101239_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1707 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1708 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1709 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X1710 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1711 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1712 a_100929_n7688# CM_p_net_1.IN a_100399_n11308# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1713 a_100929_n22063# CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1714 a_84952_n23087# CM_p_net_0.IN a_84384_n23087# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1715 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1716 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1717 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1718 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1719 PRbiased_net_x5_0.VDD a_65333_n40208# a_73115_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1720 a_53546_n40208# a_71343_n40268# a_73149_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1721 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1722 a_112928_5486# a_112406_4328# a_106677_10235# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1723 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1724 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1725 PRbiased_net_x5_1.ITP3 PRbiased_net_x5_1.IBP3 a_77623_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1726 a_35879_13393# a_53676_10235# a_55482_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1727 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1728 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1729 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1730 a_108483_n40208# a_106677_n40268# a_106523_n31143# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1731 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1732 a_89378_6252# a_83000_11461# PRbiased_net_x5_1.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1733 a_77594_n31143# a_77072_n33067# a_77072_n33067# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1734 PRbiased_net_x5_0.ITP2 a_47838_n33199# a_59956_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1735 a_71743_n38276# a_71343_n40268# PRbiased_net_x5_0.IBP3 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1736 a_29855_n4405# CM_n_net_1.IN a_29333_n4405# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1737 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1738 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1739 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1740 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1741 a_30171_n33199# a_29999_n40208# a_36377_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1742 a_31975_n32301# a_30171_n33199# PRbiased_net_x5_0.ITN1 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1743 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1744 a_106677_n40268# a_112406_n33067# a_114332_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1745 a_31849_n15070# CM_n_net_1.IN a_31289_n15070# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1746 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1747 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1748 a_106627_n8593# CM_p_net_1.IN a_106097_n9498# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1749 a_50520_n20580# CM_n_net_0.IN a_49960_n20580# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1750 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1751 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1752 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1753 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1754 a_83546_n23087# CM_p_net_0.IN a_83016_n23087# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1755 a_50520_n17889# CM_n_net_0.IN a_49960_n17889# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1756 PRbiased_net_x5_1.ITP3 PRbiased_net_x5_1.IBP3 a_77623_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1757 PRbiased_net_x5_1.IBP2 a_53676_10235# a_55482_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1758 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1759 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1760 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1761 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1762 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1763 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1764 a_49960_n21477# CM_n_net_0.IN a_49438_n21477# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1765 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1766 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1767 CM_input_0.ISBCS CM_input_0.ISBCS a_75637_n15093# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X1768 a_49960_n18786# CM_n_net_0.IN a_49438_n19683# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1769 a_114299_n11308# CM_p_net_1.IN a_113731_n11308# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1770 a_113163_n22968# CM_p_net_1.IN a_112325_n22968# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1771 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1772 a_101197_n39042# a_100667_n39042# a_100667_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1773 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1774 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1775 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1776 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1777 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1778 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X1779 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1780 a_95780_n8712# CM_p_net_0.IN a_94942_n8712# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1781 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1782 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1783 PRbiased_net_x5_1.VDD a_65333_10295# a_65863_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1784 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1785 a_109439_n7688# CM_p_net_1.IN CM_p_net_1.OUT4 CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1786 a_65905_5486# PRbiased_net_x5_1.IBN3 a_65333_11461# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1787 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1788 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1789 a_63052_n16095# CM_n_net_0.IN a_62492_n16095# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1790 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1791 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1792 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1793 a_37781_5486# a_29999_11461# PRbiased_net_x5_1.IBN1 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1794 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1795 a_96348_n9617# CM_p_net_0.IN a_95780_n9617# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1796 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1797 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1798 a_65920_n10812# CM_n_net_0.IN a_65360_n9915# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1799 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1800 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1801 a_92056_n19467# CM_p_net_0.IN CM_p_net_0.OUT10 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1802 a_9305_n11560# a_n7828_n21089# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1803 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1804 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1805 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1806 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1807 a_112325_n7688# CM_p_net_1.IN a_111795_n11308# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1808 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1809 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1810 a_100839_n33199# a_100667_n40208# a_107045_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1811 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1812 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1813 a_42947_n20452# CM_n_net_1.IN a_42387_n20452# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1814 PRbiased_net_x5_0.ITP3 a_65505_n33199# a_77623_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1815 a_42947_n17761# CM_n_net_1.IN a_42387_n17761# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1816 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1817 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1818 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1819 a_71318_n10715# a_71318_n10715# a_75654_n10715# CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X1820 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1821 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1822 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1823 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1824 a_56786_n16095# CM_n_net_0.IN a_56226_n16095# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1825 a_31289_n21349# CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1826 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1827 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1828 a_114299_n15728# CM_p_net_1.IN a_113731_n15728# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1829 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1830 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1831 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1832 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1833 a_85520_n3282# CM_p_net_0.IN a_84952_n3282# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1834 a_88856_n34225# a_89010_n40268# a_89410_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1835 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1836 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1837 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1838 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1839 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1840 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1841 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1842 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1843 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1844 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1845 a_83546_n5092# CM_p_net_0.IN a_83016_n5997# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1846 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1847 a_89010_10235# PRbiased_net_x5_1.IBP4 a_96696_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1848 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1849 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1850 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1851 a_78998_n34225# a_77072_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1852 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1853 a_83546_n19467# CM_p_net_0.IN a_83016_n18562# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1854 a_103741_n7688# CM_p_net_1.IN CM_p_net_1.OUT2 CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1855 PRbiased_net_x5_1.VDD a_47666_11461# a_55448_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1856 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1857 a_106677_n40268# a_112406_n33067# a_114332_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1858 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1859 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1860 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1861 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1862 a_31289_n10684# CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1863 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1864 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1865 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1866 a_102603_n37110# a_100667_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1867 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1868 a_45255_n8890# CM_n_net_1.IN a_44733_n9787# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1869 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1870 a_61331_n33067# a_59405_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1871 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1872 a_101767_n9498# CM_p_net_1.IN a_100929_n9498# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1873 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1874 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1875 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1876 a_50520_n10812# CM_n_net_0.IN a_49960_n10812# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1877 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1878 CM_p_net_0.VDD CM_p_net_0.IN a_91218_n23087# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1879 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1880 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1881 a_102903_n4973# CM_p_net_1.IN a_102335_n4973# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1882 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1883 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1884 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1885 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1886 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1887 a_42289_n37110# a_30171_n33199# a_41738_n33067# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1888 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1889 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1890 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1891 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1892 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1893 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1894 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1895 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1896 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1897 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1898 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1899 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1900 a_100929_n7688# CM_p_net_1.IN a_100399_n6783# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1901 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1902 a_73149_10295# a_71343_10235# a_71189_7410# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1903 a_89244_n9617# CM_p_net_0.IN a_88714_n9617# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1904 a_84952_n22182# CM_p_net_0.IN a_84384_n22182# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1905 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1906 a_36009_10235# a_41738_4328# a_43664_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1907 a_65360_n6327# CM_n_net_0.IN a_64838_n8121# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1908 a_42947_n7993# CM_n_net_1.IN a_42387_n7993# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1909 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1910 a_49642_7410# a_47838_4268# PRbiased_net_x5_1.ITN2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1911 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1912 a_54044_5486# a_47666_11461# PRbiased_net_x5_1.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1913 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1914 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1915 a_n7408_n26036# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X1916 a_62492_n9018# CM_n_net_0.IN a_61970_n9018# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1917 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1918 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1919 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1920 a_108449_n33067# a_100667_n40208# PRbiased_net_x5_0.IBN5 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1921 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1922 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1923 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1924 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1925 CM_n_net_1.VSS a_94739_n33067# a_95261_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1926 a_64486_n9018# CM_n_net_0.IN a_63926_n9018# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1927 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1928 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1929 PRbiased_net_x5_0.IBN5 a_100667_n40208# a_107045_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1930 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1931 FC_top_0.AVDD FC_top_0.IREF a_n7828_n20082# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1932 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1933 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1934 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1935 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1936 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1937 PRbiased_net_x5_0.VDD a_65333_n39042# a_65863_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1938 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1939 a_94739_n33067# a_83172_n33199# a_96696_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1940 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1941 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1942 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1943 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1944 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1945 a_83546_n22182# CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1946 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1947 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1948 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1949 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1950 a_94942_n5092# CM_p_net_0.IN a_94412_n5997# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1951 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1952 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X1953 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1954 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1955 a_32723_n5302# CM_n_net_1.IN a_32201_n5302# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1956 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1957 a_88856_4328# a_83000_11461# a_90782_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1958 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1959 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1960 a_95290_n38276# PRbiased_net_x5_0.IBP4 a_89010_n40268# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1961 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1962 a_100667_11461# PRbiased_net_x5_1.IBN5 a_102643_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1963 PRbiased_net_x5_1.ITN1 a_30171_4268# a_30571_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X1964 a_114299_n10403# CM_p_net_1.IN a_113731_n10403# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1965 a_45255_n15070# CM_n_net_1.IN a_44733_n15967# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1966 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1967 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1968 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1969 a_106523_4328# a_106677_10235# a_107077_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1970 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1971 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1972 a_114332_4328# a_112406_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1973 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1974 a_42260_4328# a_41738_4328# a_41738_4328# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1975 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1976 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1977 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X1978 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1979 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1980 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1981 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1982 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1983 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X1984 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1985 a_113163_n9498# CM_p_net_1.IN a_112325_n9498# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1986 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1987 a_109439_n7688# CM_p_net_1.IN a_108909_n6783# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1988 PRbiased_net_x5_0.ITP4 PRbiased_net_x5_0.IBP4 a_95290_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1989 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X1990 a_78998_n32301# a_77072_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1991 a_97754_n5092# CM_p_net_0.IN a_96916_n4187# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X1992 a_89410_13393# a_89010_10235# a_88880_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1993 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1994 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1995 a_112928_7410# a_112406_4328# a_106677_10235# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1996 a_113731_n4068# CM_p_net_1.IN a_113163_n4068# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X1997 a_31935_n38276# a_29999_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X1998 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X1999 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2000 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2001 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2002 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2003 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2004 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2005 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2006 a_96348_n8712# CM_p_net_0.IN a_95780_n8712# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2007 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2008 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2009 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2010 CM_input_0.IP CM_input_0.ISBCS a_75637_n17669# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X2011 a_92056_n19467# CM_p_net_0.IN a_91526_n18562# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2012 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2013 a_61331_n31143# a_59405_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2014 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X2015 a_38989_n15070# CM_n_net_1.IN a_38467_n15967# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2016 a_112325_n7688# CM_p_net_1.IN a_111795_n6783# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2017 a_57660_n20580# CM_n_net_0.IN a_57138_n20580# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2018 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2019 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2020 a_36681_n9787# CM_n_net_1.IN a_36121_n9787# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2021 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2022 a_89410_11461# a_89010_10235# PRbiased_net_x5_1.IBP4 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2023 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2024 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2025 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2026 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2027 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2028 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2029 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2030 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2031 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2032 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2033 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2034 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2035 a_30529_n38276# a_29999_n39042# a_29999_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2036 a_56786_n8121# CM_n_net_0.IN a_56226_n6327# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2037 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2038 a_114299_n14823# CM_p_net_1.IN a_113731_n14823# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2039 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2040 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2041 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2042 PRbiased_net_x5_1.ITP1 a_30171_4268# a_42289_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2043 a_102903_n22063# CM_p_net_1.IN a_102335_n22063# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2044 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2045 a_30529_12227# a_29999_10295# a_29999_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2046 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2047 a_115137_n8593# CM_p_net_1.IN a_114299_n5878# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2048 a_31849_n15070# CM_n_net_1.IN a_31289_n14173# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2049 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2050 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X2051 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2052 a_83530_n39042# a_83000_n39042# a_83000_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2053 a_50520_n18786# CM_n_net_0.IN a_49960_n16992# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2054 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2055 a_51954_n5430# CM_n_net_0.IN a_51394_n5430# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2056 a_96665_n33067# a_94739_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2057 a_65905_7410# PRbiased_net_x5_1.IBN3 a_65333_11461# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2058 a_108449_n31143# a_100667_n40208# a_100839_n33199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2059 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2060 CM_n_net_1.VSS a_94739_n33067# a_95261_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2061 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2062 a_37781_7410# a_29999_11461# a_30171_4268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2063 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2064 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2065 PRbiased_net_x5_0.VDD a_47666_n40208# a_55448_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2066 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2067 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2068 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2069 a_103741_n7688# CM_p_net_1.IN a_103211_n6783# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2070 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2071 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2072 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2073 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2074 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2075 a_85520_n23087# CM_p_net_0.IN a_84952_n23087# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2076 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2077 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2078 a_61362_12227# PRbiased_net_x5_1.IBP2 PRbiased_net_x5_1.ITP2 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2079 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2080 a_64486_n15198# CM_n_net_0.IN a_63926_n15198# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2081 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2082 a_35879_n40208# a_36009_n40268# a_37815_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2083 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2084 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2085 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2086 a_101767_n8593# CM_p_net_1.IN a_100929_n8593# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2087 a_100667_n40208# a_100667_n39042# a_102603_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2088 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2089 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2090 a_92056_n22182# CM_p_net_0.IN a_91218_n22182# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2091 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2092 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2093 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2094 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2095 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2096 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2097 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2098 a_51394_n16095# CM_n_net_0.IN a_50872_n16095# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2099 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2100 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2101 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2102 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2103 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2104 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2105 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2106 a_37815_12227# a_36009_10235# CM_n_net_1.VSS PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2107 a_59956_12227# a_47838_4268# a_59405_4328# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2108 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2109 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2110 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2111 a_63926_n9018# CM_n_net_0.IN a_63404_n9915# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2112 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2113 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2114 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2115 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2116 a_35855_n31143# a_36009_n40268# a_36409_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2117 a_48196_n38276# a_47666_n39042# a_47666_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2118 a_89244_n8712# CM_p_net_0.IN a_88714_n9617# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2119 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2120 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2121 a_113731_n22968# CM_p_net_1.IN a_113163_n22968# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2122 a_30415_n20452# CM_n_net_1.IN a_29855_n19555# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2123 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2124 PRbiased_net_x5_0.VDD a_100667_n39042# a_101197_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2125 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2126 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2127 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2128 a_31289_n20452# CM_n_net_1.IN a_30767_n20452# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2129 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2130 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2131 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2132 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2133 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2134 a_42387_n5302# CM_n_net_1.IN a_41865_n6199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2135 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2136 a_53522_4328# a_47666_11461# a_55448_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2137 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2138 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2139 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2140 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2141 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2142 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2143 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2144 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2145 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2146 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2147 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2148 a_57660_n10812# CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2149 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2150 a_67269_13393# a_65333_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2151 a_108033_n5878# CM_p_net_1.IN a_107465_n5878# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2152 a_101239_6252# a_100839_4268# a_100667_10295# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2153 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2154 a_57660_n9915# CM_n_net_0.IN a_57138_n9915# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2155 a_107465_n22968# CM_p_net_1.IN a_106627_n22968# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2156 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2157 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2158 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2159 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2160 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2161 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2162 a_59654_n10812# CM_n_net_0.IN a_59094_n9915# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2163 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2164 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2165 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2166 a_96665_n31143# a_94739_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2167 a_45255_n7993# CM_n_net_1.IN a_44733_n7993# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2168 a_67309_6252# PRbiased_net_x5_1.IBN3 PRbiased_net_x5_1.ITN3 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2169 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2170 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2171 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2172 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2173 a_113163_n8593# CM_p_net_1.IN a_112325_n8593# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2174 a_100667_10295# a_100667_10295# a_102603_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2175 a_67269_11461# a_65333_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2176 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2177 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2178 a_53522_n34225# a_47666_n40208# a_55448_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2179 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2180 a_97224_n6902# CM_p_net_0.IN a_96916_n3282# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2181 a_36121_n9787# CM_n_net_1.IN a_35599_n10684# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2182 a_113731_n3163# CM_p_net_1.IN a_113163_n3163# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2183 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2184 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2185 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2186 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2187 a_55482_12227# a_53676_10235# CM_n_net_1.VSS PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2188 a_n10081_n11560# a_n7828_n21089# a_9305_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2189 a_54044_7410# a_47666_11461# a_53522_7410# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2190 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2191 a_71711_n34225# a_65333_n40208# a_71189_n34225# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2192 a_38115_n10684# CM_n_net_1.IN a_37555_n9787# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2193 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2194 a_56226_n6327# CM_n_net_0.IN a_55704_n6327# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2195 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2196 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2197 a_65920_n19683# CM_n_net_0.IN a_65360_n19683# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2198 a_100667_10295# a_100667_10295# a_102603_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2199 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2200 a_38115_n21349# CM_n_net_1.IN a_37555_n21349# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2201 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2202 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2203 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2204 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2205 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2206 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2207 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2208 PRbiased_net_x5_0.VDD a_29999_n39042# a_30529_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2209 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2210 PRbiased_net_x5_0.ITN1 PRbiased_net_x5_0.IBN1 a_30571_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2211 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2212 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2213 a_36009_n40268# PRbiased_net_x5_0.IBP1 a_43695_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2214 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2215 a_62492_n8121# CM_n_net_0.IN a_61970_n9018# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2216 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2217 a_32723_n15967# CM_n_net_1.IN a_32201_n15967# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2218 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2219 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2220 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2221 FC_top_0.AVDD FC_top_0.IREF a_n7828_n20082# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2222 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2223 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2224 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2225 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2226 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2227 a_n10081_n10574# a_n7828_n21089# FC_top_0.VOUT CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2228 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2229 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2230 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X2231 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2232 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2233 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2234 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2235 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2236 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2237 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2238 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2239 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2240 a_115137_n4973# CM_p_net_1.IN a_114299_n4973# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2241 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2242 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2243 a_38989_n8890# CM_n_net_1.IN a_38467_n9787# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2244 a_59654_n19683# CM_n_net_0.IN a_59094_n19683# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2245 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2246 a_84384_n9617# CM_p_net_0.IN a_83546_n9617# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2247 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2248 a_38115_n10684# CM_n_net_1.IN a_37555_n10684# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2249 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2250 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2251 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2252 PRbiased_net_x5_0.ITP1 a_30171_n33199# a_42289_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2253 a_54076_n38276# a_53676_n40268# PRbiased_net_x5_0.IBP2 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2254 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2255 CM_n_net_1.VSS a_77072_4328# a_77594_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2256 PRbiased_net_x5_1.IBN4 a_83000_11461# a_89378_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2257 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2258 a_45255_n14173# CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2259 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2260 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2261 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2262 a_50520_n9915# CM_n_net_0.IN a_49960_n9018# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2263 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2264 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2265 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2266 a_85520_n22182# CM_p_net_0.IN a_84952_n22182# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2267 a_36121_n15967# CM_n_net_1.IN a_35599_n16864# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2268 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2269 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2270 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2271 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2272 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2273 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2274 a_35855_7410# a_36009_10235# a_36409_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2275 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2276 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2277 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2278 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2279 a_59094_n6327# CM_n_net_0.IN a_58572_n8121# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2280 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2281 a_79029_n38276# a_65505_n33199# PRbiased_net_x5_0.ITP3 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2282 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2283 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2284 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2285 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2286 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2287 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2288 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2289 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2290 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2291 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2292 a_83000_10295# a_83000_10295# a_84936_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2293 PRbiased_net_x5_0.ITN5 a_100839_n33199# a_101239_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2294 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2295 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2296 a_38989_n14173# CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2297 CM_n_net_1.VSS a_36009_10235# a_36409_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2298 a_63926_n14301# CM_n_net_0.IN a_63052_n17889# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2299 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2300 a_113163_n22063# CM_p_net_1.IN a_112325_n22063# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2301 PRbiased_net_x5_0.VDD a_65333_n40208# a_73115_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2302 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2303 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2304 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2305 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2306 a_n7828_n21089# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2307 a_29855_n15967# CM_n_net_1.IN a_29333_n16864# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2308 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2309 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2310 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2311 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2312 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2313 a_71711_n32301# a_65333_n40208# PRbiased_net_x5_0.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2314 a_65920_n6327# CM_n_net_0.IN a_65360_n5430# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2315 a_83000_10295# a_83000_10295# a_84936_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2316 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2317 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2318 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2319 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2320 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2321 a_101767_n17538# CM_p_net_1.IN a_100929_n17538# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2322 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2323 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2324 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2325 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2326 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2327 a_31975_n33067# PRbiased_net_x5_0.IBN1 PRbiased_net_x5_0.ITN1 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2328 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2329 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2330 a_53676_10235# a_59405_4328# a_61331_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2331 PRbiased_net_x5_0.ITN1 PRbiased_net_x5_0.IBN1 a_30571_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2332 a_95780_n23087# CM_p_net_0.IN a_94942_n23087# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2333 a_43821_n19555# CM_n_net_1.IN a_43299_n20452# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2334 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2335 a_51954_n4533# CM_n_net_0.IN a_51394_n4533# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2336 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2337 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2338 a_29999_n39042# a_29999_n39042# a_31935_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2339 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2340 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2341 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2342 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2343 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2344 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2345 a_108033_n4973# CM_p_net_1.IN a_107465_n4973# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2346 a_107465_n4068# CM_p_net_1.IN a_106627_n4068# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2347 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2348 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2349 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2350 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2351 a_61362_n38276# a_47838_n33199# PRbiased_net_x5_0.ITP2 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2352 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2353 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2354 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2355 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2356 a_53546_13393# a_53676_10235# a_55482_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2357 PRbiased_net_x5_1.ITP3 a_65505_4268# a_77623_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2358 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2359 a_65863_12227# a_65333_10295# a_65333_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2360 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2361 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2362 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2363 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2364 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2365 a_37555_n19555# CM_n_net_1.IN a_37033_n20452# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2366 PRbiased_net_x5_0.ITN3 PRbiased_net_x5_0.IBN3 a_65905_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2367 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2368 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2369 a_71343_n40268# PRbiased_net_x5_0.IBP3 a_79029_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2370 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2371 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2372 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2373 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2374 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2375 a_89244_n17657# CM_p_net_0.IN a_88714_n17657# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2376 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2377 a_62492_n3636# CM_n_net_0.IN a_61970_n4533# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2378 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2379 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2380 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2381 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2382 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2383 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2384 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2385 a_64486_n4533# CM_n_net_0.IN a_63926_n3636# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2386 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2387 CM_input_0.IN a_71318_n10715# a_75654_n9756# CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X2388 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2389 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2390 a_101767_n21158# CM_p_net_1.IN a_100929_n21158# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2391 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2392 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2393 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2394 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2395 PRbiased_net_x5_0.ITN5 a_100839_n33199# a_101239_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2396 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2397 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2398 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2399 a_42387_n16864# CM_n_net_1.IN a_41865_n16864# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2400 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2401 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2402 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2403 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2404 a_71189_n34225# a_65333_n40208# a_73115_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2405 a_47666_n39042# a_47666_n39042# a_49602_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2406 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2407 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2408 a_36681_n18658# CM_n_net_1.IN a_36121_n16864# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2409 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2410 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2411 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2412 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2413 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2414 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2415 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2416 a_84384_n8712# CM_p_net_0.IN a_83546_n8712# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2417 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2418 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2419 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2420 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2421 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2422 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2423 PRbiased_net_x5_1.IBN2 a_47666_11461# a_54044_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2424 CM_input_0.IN2 a_71318_n10715# a_75654_n11674# CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X2425 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2426 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2427 a_31975_n31143# PRbiased_net_x5_0.IBN1 PRbiased_net_x5_0.ITN1 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2428 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2429 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2430 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2431 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2432 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2433 CM_n_net_1.VSS a_77072_n33067# a_77594_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2434 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2435 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2436 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2437 a_72655_n15093# CM_input_0.ISBCS CM_input_0.IP CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X2438 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2439 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2440 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2441 PRbiased_net_x5_0.VDD a_47666_n39042# a_48196_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2442 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2443 a_58220_n16095# CM_n_net_0.IN a_57660_n16095# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2444 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2445 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2446 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2447 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2448 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2449 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2450 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2451 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2452 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2453 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2454 a_89244_n21277# CM_p_net_0.IN a_88714_n21277# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2455 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2456 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2457 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2458 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2459 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2460 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2461 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2462 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2463 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2464 PRbiased_net_x5_1.ITN5 a_100839_4268# a_101239_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2465 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2466 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2467 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2468 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2469 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2470 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2471 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2472 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2473 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2474 a_38115_n21349# CM_n_net_1.IN a_37555_n20452# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2475 CM_n_net_1.VSS a_41738_4328# a_42260_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2476 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2477 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2478 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2479 a_71743_13393# a_71343_10235# a_71213_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2480 PRbiased_net_x5_0.ITN3 PRbiased_net_x5_0.IBN3 a_65905_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2481 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2482 a_65333_11461# PRbiased_net_x5_1.IBN3 a_67309_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2483 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2484 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2485 a_90650_n17657# CM_p_net_0.IN a_90082_n17657# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2486 a_31289_n4405# CM_n_net_1.IN a_30767_n5302# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2487 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2488 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2489 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2490 a_78998_4328# a_77072_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2491 PRbiased_net_x5_0.IBN5 a_100667_n40208# a_107045_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2492 a_101767_n16633# CM_p_net_1.IN a_100929_n16633# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2493 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2494 CM_n_net_1.VSS a_77072_4328# a_77594_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2495 a_102643_n34225# a_100839_n33199# PRbiased_net_x5_0.ITN5 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2496 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2497 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2498 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2499 a_96696_n38276# a_83172_n33199# PRbiased_net_x5_0.ITP4 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2500 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2501 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2502 a_42947_n5302# CM_n_net_1.IN a_42387_n4405# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2503 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2504 a_71743_11461# a_71343_10235# PRbiased_net_x5_1.IBP3 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2505 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2506 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2507 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2508 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2509 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2510 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2511 a_95780_n22182# CM_p_net_0.IN a_94942_n22182# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2512 a_38989_n7993# CM_n_net_1.IN a_38467_n7993# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2513 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2514 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2515 a_90782_4328# a_83000_11461# a_83172_4268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2516 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2517 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2518 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2519 a_33283_n6199# CM_n_net_1.IN a_32723_n5302# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2520 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2521 a_29855_n9787# CM_n_net_1.IN a_29333_n10684# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2522 a_107465_n3163# CM_p_net_1.IN a_106627_n3163# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2523 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2524 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2525 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2526 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2527 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2528 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X2529 a_50520_n8121# CM_n_net_0.IN a_49960_n8121# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2530 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2531 a_107077_12227# a_106677_10235# PRbiased_net_x5_1.IBP5 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2532 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2533 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2534 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2535 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2536 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2537 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2538 a_65863_n39042# a_65333_n39042# a_65333_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2539 a_96348_n17657# CM_p_net_0.IN a_95780_n17657# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2540 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2541 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2542 a_78998_n33067# a_77072_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2543 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2544 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2545 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2546 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2547 PRbiased_net_x5_0.IBP2 a_53676_n40268# a_55482_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2548 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2549 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2550 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2551 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2552 a_9305_n11560# a_n7828_n21089# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2553 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2554 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2555 CM_n_net_1.VSS a_77072_n33067# a_77594_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2556 a_63926_n3636# CM_n_net_0.IN a_63052_n7224# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2557 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2558 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2559 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2560 a_51954_n21477# CM_n_net_0.IN a_51394_n21477# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2561 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2562 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2563 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2564 a_49960_n7224# CM_n_net_0.IN CM_n_net_0.OUT2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2565 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2566 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2567 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2568 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2569 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2570 a_89244_n16752# CM_p_net_0.IN a_88714_n17657# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2571 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2572 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2573 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2574 a_114332_n34225# a_112406_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2575 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2576 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2577 a_n7828_n20082# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X2578 a_90650_n21277# CM_p_net_0.IN a_90082_n21277# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2579 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2580 a_47666_10295# a_47666_10295# a_49602_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2581 a_53388_n15198# CM_n_net_0.IN a_52828_n14301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2582 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2583 a_101767_n20253# CM_p_net_1.IN a_100929_n20253# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2584 CM_n_net_1.VSS a_53676_n40268# a_54076_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2585 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2586 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2587 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2588 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2589 a_65920_n4533# CM_n_net_0.IN a_65360_n4533# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2590 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2591 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2592 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2593 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2594 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2595 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2596 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2597 a_37781_n34225# a_29999_n40208# a_30171_n33199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2598 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2599 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2600 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2601 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2602 a_42289_12227# a_30171_4268# a_41738_4328# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2603 a_n7828_n21089# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2604 a_89410_10295# a_89010_10235# a_71213_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2605 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2606 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2607 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2608 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2609 a_49642_6252# PRbiased_net_x5_1.IBN2 PRbiased_net_x5_1.ITN2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2610 a_47666_10295# a_47666_10295# a_49602_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2611 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2612 a_30415_n15967# CM_n_net_1.IN a_29855_n15070# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2613 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2614 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2615 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X2616 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2617 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2618 a_90816_12227# a_89010_10235# CM_n_net_1.VSS PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2619 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2620 a_103741_n20253# CM_p_net_1.IN a_102903_n17538# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2621 a_33283_n19555# CM_n_net_1.IN a_32723_n19555# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2622 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2623 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2624 CM_n_net_1.VSS a_94739_n33067# a_95261_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2625 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2626 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2627 a_100839_n33199# a_100667_n40208# a_107045_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2628 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2629 a_102643_n32301# a_100839_n33199# PRbiased_net_x5_0.ITN5 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2630 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2631 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2632 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2633 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2634 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2635 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2636 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2637 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2638 a_96348_n21277# CM_p_net_0.IN a_95780_n21277# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2639 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2640 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2641 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2642 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2643 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2644 a_86358_n5092# CM_p_net_0.IN a_85520_n4187# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2645 a_113731_n22063# CM_p_net_1.IN a_113163_n22063# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2646 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2647 a_102335_n4068# CM_p_net_1.IN a_101767_n4068# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2648 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2649 a_n7828_n20082# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2650 a_107077_n37110# a_106677_n40268# a_88880_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2651 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2652 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2653 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2654 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2655 PRbiased_net_x5_1.VDD a_83000_11461# a_90782_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2656 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2657 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2658 a_49960_n14301# CM_n_net_0.IN a_49438_n15198# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2659 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2660 PRbiased_net_x5_1.VDD a_83000_10295# a_83530_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2661 a_57660_n5430# CM_n_net_0.IN a_57138_n5430# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2662 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2663 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2664 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2665 a_89244_n20372# CM_p_net_0.IN a_88714_n21277# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2666 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2667 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2668 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2669 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2670 a_59654_n6327# CM_n_net_0.IN a_59094_n5430# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2671 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2672 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2673 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2674 a_75654_n10715# a_71318_n10715# CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X2675 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2676 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2677 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2678 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2679 a_78998_n31143# a_77072_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2680 a_112957_13393# PRbiased_net_x5_1.IBP5 a_106677_10235# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2681 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2682 a_112928_6252# a_112406_4328# a_112406_4328# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2683 a_107465_n22063# CM_p_net_1.IN a_106627_n22063# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2684 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2685 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2686 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2687 a_72655_n17669# CM_input_0.ISBCS CM_input_0.ISBCS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X2688 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2689 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2690 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2691 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2692 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2693 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2694 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2695 a_71743_n39042# a_71343_n40268# PRbiased_net_x5_0.IBP3 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2696 FC_top_0.VOUT a_n7828_n21089# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2697 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2698 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2699 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2700 a_59405_n33067# a_47838_n33199# a_61362_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2701 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2702 a_55448_4328# a_47666_11461# a_47838_4268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2703 a_90650_n16752# CM_p_net_0.IN a_90082_n16752# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2704 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2705 a_54044_n34225# a_47666_n40208# a_53522_n34225# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2706 a_47838_4268# a_47666_11461# a_54044_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2707 a_114332_n32301# a_112406_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2708 a_65920_n15198# CM_n_net_0.IN a_65360_n15198# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2709 a_112957_11461# PRbiased_net_x5_1.IBP5 a_106677_10235# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2710 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2711 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2712 a_103741_n22063# CM_p_net_1.IN a_102903_n21158# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2713 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2714 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2715 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2716 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2717 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2718 a_n7408_n26036# a_n7408_n26036# a_2944_n20707# FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0.78p ps=3.7u w=1.2u l=2u
X2719 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2720 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2721 a_n2230_n25376# a_n7828_n21089# a_n7828_n21089# CM_n_net_1.VSS nfet_03v3 ad=0.48p pd=2u as=0.732p ps=3.62u w=1.2u l=2u
X2722 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2723 CM_n_net_0.OUT1 CM_n_net_0.IN a_49960_n3636# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2724 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2725 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2726 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2727 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2728 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2729 a_37781_n32301# a_29999_n40208# PRbiased_net_x5_0.IBN1 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2730 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2731 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2732 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2733 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2734 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2735 PRbiased_net_x5_0.ITP2 PRbiased_net_x5_0.IBP2 a_59956_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2736 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2737 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2738 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2739 a_45815_n16864# CM_n_net_1.IN a_45255_n16864# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2740 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2741 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2742 PRbiased_net_x5_0.VDD a_83000_n39042# a_83530_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2743 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2744 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2745 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2746 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2747 a_65905_6252# a_65505_4268# a_65333_10295# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2748 PRbiased_net_x5_1.ITP2 a_47838_4268# a_59956_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2749 a_101197_n40208# a_100667_n39042# a_100667_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2750 a_59654_n15198# CM_n_net_0.IN a_59094_n15198# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2751 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2752 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2753 a_91218_n11427# CM_p_net_0.IN a_90650_n11427# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2754 CM_n_net_1.VSS a_94739_n33067# a_95261_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2755 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2756 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2757 a_96348_n16752# CM_p_net_0.IN a_95780_n16752# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2758 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2759 a_37781_6252# a_29999_11461# PRbiased_net_x5_1.IBN1 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2760 a_114363_n37110# PRbiased_net_x5_0.IBP5 PRbiased_net_x5_0.ITP5 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2761 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2762 CM_p_net_0.VDD CM_p_net_0.IN a_85520_n11427# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2763 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2764 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2765 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2766 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2767 a_106523_n31143# a_100667_n40208# a_108449_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2768 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2769 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2770 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2771 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2772 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2773 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2774 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2775 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2776 a_45255_n4405# CM_n_net_1.IN a_44733_n5302# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2777 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2778 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2779 a_52828_n7224# CM_n_net_0.IN a_51954_n5430# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2780 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2781 a_39549_n16864# CM_n_net_1.IN a_38989_n16864# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2782 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2783 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2784 a_67269_10295# a_65333_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2785 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2786 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2787 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2788 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2789 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2790 a_90650_n20372# CM_p_net_0.IN a_90082_n20372# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2791 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2792 a_112957_n37110# a_100839_n33199# a_112406_n33067# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2793 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X2794 a_65360_n21477# CM_n_net_0.IN a_63052_n21477# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2795 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2796 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2797 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2798 a_75654_n9756# a_71318_n10715# CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X2799 a_65360_n18786# CM_n_net_0.IN a_64838_n18786# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2800 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2801 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2802 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2803 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2804 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X2805 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2806 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2807 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2808 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2809 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X2810 a_100667_11461# a_100667_10295# a_102603_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2811 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2812 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2813 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2814 a_83000_n39042# a_83172_n33199# a_84976_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2815 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2816 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2817 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2818 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2819 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2820 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2821 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2822 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2823 a_91218_n15847# CM_p_net_0.IN a_90650_n15847# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2824 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2825 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2826 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2827 PRbiased_net_x5_0.ITP3 PRbiased_net_x5_0.IBP3 a_77623_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2828 a_86358_n16752# CM_p_net_0.IN a_85520_n15847# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2829 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X2830 a_n7828_n20082# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2831 a_41738_4328# a_41738_4328# a_43664_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2832 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2833 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2834 a_54044_n32301# a_47666_n40208# PRbiased_net_x5_0.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2835 a_103741_n16633# CM_p_net_1.IN a_102903_n16633# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2836 PRbiased_net_x5_1.VDD a_47666_11461# a_55448_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2837 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2838 a_59094_n21477# CM_n_net_0.IN a_56786_n21477# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2839 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2840 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2841 a_59094_n18786# CM_n_net_0.IN a_58572_n18786# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2842 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2843 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2844 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2845 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X2846 a_96348_n20372# CM_p_net_0.IN a_95780_n20372# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2847 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2848 a_85828_n6902# CM_p_net_0.IN a_85520_n3282# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2849 a_43821_n15070# CM_n_net_1.IN a_43299_n15967# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2850 a_102335_n3163# CM_p_net_1.IN a_101767_n3163# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2851 a_88880_n40208# a_89010_n40268# a_90816_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2852 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2853 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2854 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2855 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2856 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2857 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2858 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2859 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2860 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X2861 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2862 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2863 FC_top_0.VOUT a_n7828_n21089# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2864 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2865 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2866 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2867 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2868 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2869 a_94739_4328# a_83172_4268# a_96696_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2870 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2871 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2872 a_63052_n20580# CM_n_net_0.IN a_62492_n20580# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2873 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2874 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2875 a_63052_n17889# CM_n_net_0.IN a_62492_n17889# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2876 a_100667_10295# a_100839_4268# a_102643_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2877 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2878 PRbiased_net_x5_1.ITN1 PRbiased_net_x5_1.IBN1 a_30571_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2879 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2880 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2881 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2882 a_102603_n38276# a_100667_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2883 a_114332_5486# a_112406_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2884 a_37555_n15070# CM_n_net_1.IN a_37033_n15967# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2885 a_42260_5486# a_41738_4328# a_36009_10235# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2886 a_94739_n33067# a_94739_n33067# a_96665_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2887 a_54044_6252# a_47666_11461# PRbiased_net_x5_1.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2888 PRbiased_net_x5_0.VDD a_100667_n40208# a_108449_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2889 PRbiased_net_x5_0.ITN2 PRbiased_net_x5_0.IBN2 a_48238_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2890 a_71711_n33067# a_65333_n40208# PRbiased_net_x5_0.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2891 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2892 a_94739_4328# a_83172_4268# a_96696_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2893 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2894 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2895 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2896 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2897 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2898 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2899 a_44381_n8890# CM_n_net_1.IN a_45255_n7096# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2900 a_35855_4328# a_36009_10235# a_36409_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2901 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2902 a_42289_n38276# PRbiased_net_x5_0.IBP1 a_36009_n40268# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2903 a_31849_n4405# CM_n_net_1.IN a_31289_n3508# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2904 a_56786_n20580# CM_n_net_0.IN a_56226_n20580# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2905 a_36681_n5302# CM_n_net_1.IN a_36121_n5302# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2906 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2907 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2908 PRbiased_net_x5_0.VDD a_65333_n39042# a_65863_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2909 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2910 a_56786_n17889# CM_n_net_0.IN a_56226_n17889# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2911 a_96916_n17657# CM_p_net_0.IN a_96348_n17657# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2912 a_85520_n5997# CM_p_net_0.IN a_84952_n5997# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2913 PRbiased_net_x5_0.ITN1 a_30171_n33199# a_30571_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2914 a_103741_n20253# CM_p_net_1.IN a_102903_n20253# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2915 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2916 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2917 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2918 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2919 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2920 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2921 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2922 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2923 a_75637_n16769# CM_input_0.ISBCS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X2924 CM_n_net_1.OUT7 CM_n_net_1.IN a_29855_n14173# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2925 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2926 a_83000_11461# a_83000_10295# a_84936_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2927 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2928 a_44381_n21349# CM_n_net_1.IN a_43821_n21349# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2929 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2930 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2931 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2932 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2933 a_83546_n9617# CM_p_net_0.IN a_83016_n9617# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2934 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2935 a_95290_n39042# a_83172_n33199# a_94739_n33067# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2936 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2937 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2938 a_89410_n37110# a_89010_n40268# a_71213_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2939 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2940 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2941 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2942 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2943 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2944 a_83000_n39042# a_83172_n33199# a_84976_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2945 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2946 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2947 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2948 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2949 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2950 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2951 a_91218_n10522# CM_p_net_0.IN a_90650_n10522# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2952 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2953 a_31935_n39042# a_29999_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2954 a_57660_n4533# CM_n_net_0.IN a_57138_n5430# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2955 a_86358_n10522# CM_p_net_0.IN a_85520_n10522# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2956 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2957 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2958 a_44381_n10684# CM_n_net_1.IN a_43821_n10684# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2959 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2960 a_59654_n4533# CM_n_net_0.IN a_59094_n4533# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2961 FC_top_0.AVDD FC_top_0.IREF a_n7828_n21089# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2962 PRbiased_net_x5_0.VB a_106677_n40268# a_108483_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2963 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2964 a_112325_n11308# CM_p_net_1.IN a_111795_n11308# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X2965 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2966 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2967 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2968 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2969 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2970 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2971 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2972 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2973 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2974 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2975 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2976 a_30529_n39042# a_29999_n39042# a_29999_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2977 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2978 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X2979 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2980 a_96916_n21277# CM_p_net_0.IN a_96348_n21277# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2981 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2982 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X2983 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2984 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2985 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2986 FC_top_0.AVDD FC_top_0.IREF a_n7828_n20082# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X2987 a_106523_n31143# a_106677_n40268# a_107077_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X2988 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X2989 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2990 a_63052_n10812# CM_n_net_0.IN a_62492_n10812# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2991 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2992 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2993 a_94739_n33067# a_94739_n33067# a_96665_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2994 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2995 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2996 PRbiased_net_x5_0.ITN2 PRbiased_net_x5_0.IBN2 a_48238_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X2997 a_71711_n31143# a_65333_n40208# a_71189_n31143# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X2998 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X2999 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3000 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3001 a_91218_n14942# CM_p_net_0.IN a_90650_n14942# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3002 a_94942_n9617# CM_p_net_0.IN a_94412_n9617# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3003 CM_n_net_1.VSS a_112406_4328# a_112928_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3004 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3005 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3006 a_85828_n18562# CM_p_net_0.IN a_85520_n14942# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3007 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3008 a_83530_n40208# a_83000_n39042# a_83000_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3009 a_30415_n7993# CM_n_net_1.IN a_29855_n6199# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3010 PRbiased_net_x5_0.ITN1 a_30171_n33199# a_30571_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3011 a_112325_n15728# CM_p_net_1.IN CM_p_net_1.OUT11 CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3012 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3013 a_62492_n21477# CM_n_net_0.IN a_61970_n21477# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3014 a_71343_10235# a_77072_4328# a_78998_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3015 a_62492_n18786# CM_n_net_0.IN a_61970_n19683# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3016 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3017 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3018 a_30529_13393# a_29999_10295# a_29999_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3019 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3020 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3021 a_56786_n10812# CM_n_net_0.IN a_56226_n10812# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3022 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3023 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3024 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3025 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3026 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3027 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3028 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3029 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3030 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3031 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3032 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3033 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3034 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3035 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3036 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3037 a_100667_n39042# a_100667_n39042# a_102603_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3038 a_30529_11461# a_29999_10295# a_29999_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3039 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3040 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3041 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3042 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3043 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3044 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3045 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3046 a_48196_n39042# a_47666_n39042# a_47666_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3047 a_61362_13393# a_47838_4268# PRbiased_net_x5_1.ITP2 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3048 PRbiased_net_x5_0.ITN3 a_65505_n33199# a_65905_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3049 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3050 a_36121_n5302# CM_n_net_1.IN a_35599_n6199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3051 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3052 PRbiased_net_x5_1.ITN3 a_65505_4268# a_65905_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3053 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3054 PRbiased_net_x5_0.IBP1 a_36009_n40268# a_37815_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3055 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3056 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3057 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3058 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3059 a_38115_n5302# CM_n_net_1.IN a_37555_n5302# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3060 a_41738_4328# a_41738_4328# a_43664_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3061 a_77594_4328# a_77072_4328# a_77072_4328# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3062 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3063 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3064 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3065 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3066 PRbiased_net_x5_0.VDD a_100667_n39042# a_101197_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3067 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3068 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3069 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3070 a_61362_11461# a_47838_4268# PRbiased_net_x5_1.ITP2 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3071 a_106677_n40268# PRbiased_net_x5_0.IBP5 a_114363_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3072 a_96916_n16752# CM_p_net_0.IN a_96348_n16752# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3073 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X3074 a_37815_13393# a_36009_10235# a_35855_4328# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3075 a_63926_n19683# CM_n_net_0.IN a_63404_n20580# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3076 a_59956_13393# PRbiased_net_x5_1.IBP2 a_53676_10235# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3077 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3078 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3079 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3080 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3081 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3082 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3083 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3084 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3085 CM_n_net_1.VSS a_36009_n40268# a_36409_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3086 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3087 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3088 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3089 a_83546_n8712# CM_p_net_0.IN a_83016_n9617# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3090 a_31849_n15967# CM_n_net_1.IN a_31289_n15967# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3091 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3092 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3093 CM_n_net_1.VSS a_59405_n33067# a_59927_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3094 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3095 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3096 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3097 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3098 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3099 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3100 a_101239_n34225# PRbiased_net_x5_0.IBN5 a_100667_n40208# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3101 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3102 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3103 a_71743_10295# a_71343_10235# a_53546_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3104 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3105 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3106 a_31975_4328# PRbiased_net_x5_1.IBN1 PRbiased_net_x5_1.ITN1 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3107 a_37815_11461# a_36009_10235# CM_n_net_1.VSS PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3108 a_43821_n14173# CM_n_net_1.IN a_42947_n17761# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3109 a_100667_10295# a_100839_4268# a_102643_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3110 a_59956_11461# PRbiased_net_x5_1.IBP2 a_53676_10235# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3111 PRbiased_net_x5_1.ITN1 PRbiased_net_x5_1.IBN1 a_30571_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3112 a_38989_n4405# CM_n_net_1.IN a_38467_n5302# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3113 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3114 a_108601_n9498# CM_p_net_1.IN a_108033_n9498# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3115 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3116 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3117 PRbiased_net_x5_0.ITP5 a_100839_n33199# a_112957_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3118 a_73115_n34225# a_65333_n40208# a_65505_n33199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3119 a_33283_n15070# CM_n_net_1.IN a_32723_n15070# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3120 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3121 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3122 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3123 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3124 a_114332_7410# a_112406_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3125 a_42260_7410# a_41738_4328# a_36009_10235# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3126 CM_n_net_1.VSS a_77072_n33067# a_77594_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3127 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3128 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3129 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3130 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3131 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3132 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3133 a_63052_n18786# CM_n_net_0.IN a_62492_n16992# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3134 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3135 CM_input_0.VDD a_71318_n10715# a_72648_n9756# CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3136 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3137 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X3138 a_43821_n3508# CM_n_net_1.IN a_42947_n7096# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3139 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3140 a_112325_n10403# CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3141 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3142 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3143 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3144 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3145 a_51394_n20580# CM_n_net_0.IN a_50872_n20580# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3146 a_45815_n4405# CM_n_net_1.IN a_45255_n3508# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3147 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3148 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3149 a_37555_n14173# CM_n_net_1.IN a_36681_n17761# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3150 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3151 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3152 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3153 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3154 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3155 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3156 a_49602_n37110# a_47666_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3157 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3158 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3159 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3160 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3161 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3162 a_96916_n20372# CM_p_net_0.IN a_96348_n20372# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3163 a_55482_13393# a_53676_10235# a_53522_4328# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3164 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3165 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3166 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3167 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3168 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3169 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3170 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3171 PRbiased_net_x5_0.ITN3 a_65505_n33199# a_65905_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3172 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3173 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3174 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3175 a_94942_n11427# CM_p_net_0.IN a_94412_n11427# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3176 a_56786_n18786# CM_n_net_0.IN a_56226_n16992# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3177 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3178 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3179 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3180 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3181 a_90082_n11427# CM_p_net_0.IN a_89244_n11427# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3182 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3183 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3184 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3185 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3186 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3187 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3188 a_44381_n21349# CM_n_net_1.IN a_43821_n20452# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3189 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3190 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3191 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X3192 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3193 a_94942_n8712# CM_p_net_0.IN a_94412_n9617# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3194 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3195 a_54076_n39042# a_53676_n40268# PRbiased_net_x5_0.IBP2 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3196 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3197 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3198 CM_n_net_1.VSS a_77072_4328# a_77594_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3199 a_102643_n33067# PRbiased_net_x5_0.IBN5 PRbiased_net_x5_0.ITN5 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3200 a_55482_11461# a_53676_10235# CM_n_net_1.VSS PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3201 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3202 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3203 a_41738_n33067# a_30171_n33199# a_43695_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3204 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3205 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3206 a_36377_n34225# a_29999_n40208# a_35855_n34225# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3207 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3208 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3209 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3210 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3211 a_47666_11461# a_47666_10295# a_49602_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3212 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3213 a_112325_n14823# CM_p_net_1.IN a_111795_n18443# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3214 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3215 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3216 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3217 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3218 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3219 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3220 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3221 a_42947_n20452# CM_n_net_1.IN a_42387_n19555# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3222 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3223 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X3224 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3225 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3226 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3227 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3228 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3229 a_79029_12227# PRbiased_net_x5_1.IBP3 PRbiased_net_x5_1.ITP3 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3230 CM_n_net_1.VSS a_59405_n33067# a_59927_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3231 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3232 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3233 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3234 a_79029_n39042# PRbiased_net_x5_0.IBP3 PRbiased_net_x5_0.ITP3 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3235 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3236 a_97754_n7807# CM_p_net_0.IN CM_p_net_0.OUT6 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3237 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X3238 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3239 FC_top_0.AVDD FC_top_0.IREF a_n7828_n20082# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3240 a_101239_n32301# PRbiased_net_x5_0.IBN5 a_100667_n40208# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3241 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3242 a_97754_n8712# CM_p_net_0.IN a_96916_n5997# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3243 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3244 PRbiased_net_x5_0.ITP1 PRbiased_net_x5_0.IBP1 a_42289_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3245 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3246 a_113731_n5878# CM_p_net_1.IN a_113163_n5878# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3247 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3248 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3249 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3250 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3251 a_71318_n10715# CM_input_0.ISBCS a_75637_n15993# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X3252 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3253 a_73115_n32301# a_65333_n40208# PRbiased_net_x5_0.IBN3 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3254 a_38115_n8890# CM_n_net_1.IN a_38989_n7096# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3255 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3256 a_94942_n15847# CM_p_net_0.IN CM_p_net_0.OUT11 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3257 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3258 a_106677_10235# PRbiased_net_x5_1.IBP5 a_114363_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3259 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3260 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3261 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3262 a_90082_n15847# CM_p_net_0.IN a_89244_n15847# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3263 CM_n_net_1.VSS a_77072_n33067# a_77594_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3264 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3265 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3266 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3267 a_32723_n6199# CM_n_net_1.IN a_32201_n7993# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3268 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3269 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3270 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3271 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3272 a_n10081_n11560# a_n7828_n21089# a_9305_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3273 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3274 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3275 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3276 a_n7828_n20082# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3277 a_114332_n33067# a_112406_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3278 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3279 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3280 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3281 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3282 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3283 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3284 a_62492_n9915# CM_n_net_0.IN a_61970_n10812# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3285 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3286 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3287 a_75654_n11674# a_71318_n10715# CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X3288 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3289 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3290 a_29999_n40208# a_29999_n39042# a_31935_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3291 a_64486_n10812# CM_n_net_0.IN a_63926_n9915# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3292 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3293 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3294 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3295 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3296 a_37781_n33067# a_29999_n40208# PRbiased_net_x5_0.IBN1 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3297 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3298 a_51394_n10812# CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3299 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3300 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3301 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3302 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3303 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3304 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3305 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3306 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3307 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3308 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X3309 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3310 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3311 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3312 a_100929_n9498# CM_p_net_1.IN a_100399_n9498# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3313 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3314 a_61362_n39042# PRbiased_net_x5_0.IBP2 PRbiased_net_x5_0.ITP2 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3315 a_112957_10295# a_100839_4268# a_112406_4328# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3316 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3317 a_31289_n9787# CM_n_net_1.IN a_30767_n9787# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3318 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3319 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3320 a_108033_n11308# CM_p_net_1.IN a_107465_n11308# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3321 a_96696_12227# PRbiased_net_x5_1.IBP4 PRbiased_net_x5_1.ITP4 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3322 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3323 a_65333_n39042# a_65505_n33199# a_67309_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3324 a_52828_n16095# CM_n_net_0.IN a_52306_n16095# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3325 a_n7828_n21089# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3326 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3327 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3328 a_2376_n20707# a_n7408_n26036# a_1808_n20707# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X3329 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3330 a_42947_n9787# CM_n_net_1.IN a_42387_n9787# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3331 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3332 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3333 a_108601_n8593# CM_p_net_1.IN a_108033_n8593# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3334 a_45255_n15967# CM_n_net_1.IN a_44733_n15967# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3335 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3336 a_102643_n31143# PRbiased_net_x5_0.IBN5 PRbiased_net_x5_0.ITN5 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3337 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3338 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3339 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3340 a_36377_n32301# a_29999_n40208# PRbiased_net_x5_0.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3341 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3342 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3343 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3344 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3345 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3346 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3347 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3348 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3349 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3350 a_106627_n11308# CM_p_net_1.IN a_106097_n11308# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3351 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3352 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3353 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3354 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3355 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3356 a_51954_n9018# CM_n_net_0.IN a_52828_n7224# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3357 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3358 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3359 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3360 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3361 a_65863_13393# a_65333_10295# a_65333_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3362 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3363 a_63052_n7224# CM_n_net_0.IN a_62492_n7224# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3364 a_56226_n16095# CM_n_net_0.IN a_55704_n16992# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3365 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3366 a_38989_n15967# CM_n_net_1.IN a_38467_n15967# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3367 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3368 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3369 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3370 a_90782_n34225# a_83000_n40208# a_83172_n33199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3371 a_77072_n33067# a_65505_n33199# a_79029_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3372 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3373 a_109439_n10403# CM_p_net_1.IN a_108601_n9498# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3374 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3375 a_108033_n15728# CM_p_net_1.IN a_107465_n15728# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3376 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3377 a_47666_n40208# a_47666_n39042# a_49602_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3378 PRbiased_net_x5_1.ITN5 PRbiased_net_x5_1.IBN5 a_101239_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3379 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3380 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3381 a_65863_11461# a_65333_10295# a_65333_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3382 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3383 a_94942_n10522# CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3384 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3385 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3386 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3387 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3388 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3389 a_90082_n10522# CM_p_net_0.IN a_89244_n10522# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3390 CM_n_net_1.VSS a_41738_4328# a_42260_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3391 a_53388_n19683# CM_n_net_0.IN a_52828_n19683# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3392 a_54044_n33067# a_47666_n40208# PRbiased_net_x5_0.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3393 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3394 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3395 PRbiased_net_x5_1.IBN2 a_47666_11461# a_54044_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3396 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3397 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3398 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3399 a_65333_10295# a_65505_4268# a_67309_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3400 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3401 a_114332_n31143# a_112406_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3402 a_112325_n9498# CM_p_net_1.IN a_111795_n9498# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3403 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3404 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3405 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3406 a_96916_n4187# CM_p_net_0.IN a_96348_n4187# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3407 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3408 a_106627_n15728# CM_p_net_1.IN CM_p_net_1.OUT9 CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3409 a_78998_5486# a_77072_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3410 PRbiased_net_x5_0.VDD a_47666_n39042# a_48196_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3411 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3412 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3413 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3414 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3415 a_37781_n31143# a_29999_n40208# a_30171_n33199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3416 a_33283_n15070# CM_n_net_1.IN a_32723_n14173# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3417 a_114299_n17538# CM_p_net_1.IN a_113731_n17538# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3418 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3419 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3420 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3421 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3422 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3423 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3424 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3425 a_29855_n5302# CM_n_net_1.IN a_29333_n6199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3426 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3427 a_97754_n7807# CM_p_net_0.IN a_97224_n6902# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3428 a_85520_n5092# CM_p_net_0.IN a_84952_n5092# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3429 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3430 a_90782_5486# a_83000_11461# PRbiased_net_x5_1.IBN4 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3431 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3432 a_42387_n6199# CM_n_net_1.IN a_41865_n6199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3433 a_65333_n39042# a_65505_n33199# a_67309_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3434 a_113731_n4973# CM_p_net_1.IN a_113163_n4973# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3435 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3436 a_50520_n21477# CM_n_net_0.IN a_49960_n21477# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3437 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3438 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3439 a_50520_n18786# CM_n_net_0.IN a_49960_n18786# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3440 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3441 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3442 a_94942_n14942# CM_p_net_0.IN a_94412_n18562# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3443 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3444 PRbiased_net_x5_0.VDD a_100667_n40208# a_108449_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3445 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3446 a_90082_n14942# CM_p_net_0.IN a_89244_n14942# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3447 a_103741_n10403# CM_p_net_1.IN a_102903_n9498# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3448 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3449 a_49960_n19683# CM_n_net_0.IN a_49438_n19683# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3450 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3451 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3452 a_51954_n15198# CM_n_net_0.IN a_51394_n14301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3453 a_63926_n9915# CM_n_net_0.IN a_63404_n9915# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3454 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3455 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3456 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3457 a_96696_n39042# PRbiased_net_x5_0.IBP4 PRbiased_net_x5_0.ITP4 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3458 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3459 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3460 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3461 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3462 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3463 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3464 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3465 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3466 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3467 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3468 CM_p_net_1.VDD CM_p_net_1.IN a_114299_n11308# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3469 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3470 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3471 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3472 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3473 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3474 a_89010_10235# PRbiased_net_x5_1.IBP4 a_96696_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3475 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3476 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3477 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3478 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X3479 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3480 a_84936_12227# a_83000_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3481 a_90782_n32301# a_83000_n40208# PRbiased_net_x5_0.IBN4 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3482 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3483 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3484 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3485 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3486 a_83000_n40208# PRbiased_net_x5_0.IBN4 a_84976_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3487 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3488 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3489 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0 ps=0 w=1.2u l=2u
X3490 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3491 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3492 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3493 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3494 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3495 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3496 a_100929_n8593# CM_p_net_1.IN a_100399_n9498# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3497 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3498 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3499 a_114299_n21158# CM_p_net_1.IN a_113731_n21158# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3500 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3501 a_108033_n10403# CM_p_net_1.IN a_107465_n10403# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3502 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3503 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3504 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3505 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3506 a_37555_n3508# CM_n_net_1.IN a_36681_n7096# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3507 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3508 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3509 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3510 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3511 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3512 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3513 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3514 a_54044_n31143# a_47666_n40208# a_53522_n31143# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3515 PRbiased_net_x5_0.IBP2 a_53676_n40268# a_55482_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3516 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3517 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3518 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3519 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3520 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3521 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X3522 a_39549_n4405# CM_n_net_1.IN a_38989_n3508# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3523 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3524 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3525 a_31289_n19555# CM_n_net_1.IN a_30767_n20452# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3526 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3527 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3528 a_65863_n40208# a_65333_n39042# a_65333_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3529 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3530 a_58220_n21477# CM_n_net_0.IN a_57660_n20580# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3531 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3532 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3533 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3534 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3535 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3536 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3537 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3538 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3539 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3540 a_106627_n10403# CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3541 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3542 a_72648_n9756# a_71318_n10715# CM_input_0.IN2 CM_input_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X3543 a_107077_13393# a_106677_10235# PRbiased_net_x5_1.VB PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3544 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3545 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3546 a_115137_n16633# CM_p_net_1.IN a_114299_n15728# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3547 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3548 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3549 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3550 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3551 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3552 CM_n_net_1.VSS a_53676_n40268# a_54076_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3553 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3554 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3555 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X3556 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3557 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3558 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3559 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3560 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3561 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3562 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3563 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3564 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3565 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3566 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3567 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3568 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3569 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3570 a_77623_n37110# a_65505_n33199# a_77072_n33067# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3571 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3572 a_109439_n8593# CM_p_net_1.IN a_108601_n8593# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3573 a_107077_11461# a_106677_10235# PRbiased_net_x5_1.IBP5 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3574 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3575 a_108033_n14823# CM_p_net_1.IN a_107465_n14823# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3576 a_89010_n40268# a_94739_n33067# a_96665_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3577 a_45255_n9787# CM_n_net_1.IN a_44733_n9787# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3578 a_106523_n34225# a_100667_n40208# a_108449_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3579 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3580 PRbiased_net_x5_0.ITN2 a_47838_n33199# a_48238_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3581 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3582 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3583 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3584 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3585 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3586 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3587 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3588 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X3589 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3590 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3591 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3592 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3593 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3594 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3595 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3596 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3597 a_112325_n8593# CM_p_net_1.IN a_111795_n9498# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3598 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3599 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3600 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3601 a_55448_5486# a_47666_11461# PRbiased_net_x5_1.IBN2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3602 a_96916_n3282# CM_p_net_0.IN a_96348_n3282# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3603 a_107465_n5878# CM_p_net_1.IN a_106627_n5878# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3604 a_63926_n15198# CM_n_net_0.IN a_63404_n16095# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3605 a_106627_n14823# CM_p_net_1.IN a_106097_n18443# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3606 a_42289_13393# PRbiased_net_x5_1.IBP1 a_36009_10235# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3607 a_29999_11461# a_29999_10295# a_31935_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3608 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3609 CM_n_net_1.VSS a_53676_10235# a_54076_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3610 a_65360_n7224# CM_n_net_0.IN a_64486_n5430# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3611 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3612 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3613 FC_top_0.VOUT a_n7828_n21089# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3614 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3615 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3616 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3617 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3618 a_50520_n9915# CM_n_net_0.IN a_49960_n9915# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3619 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3620 a_114299_n16633# CM_p_net_1.IN a_113731_n16633# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3621 a_83000_n40208# PRbiased_net_x5_0.IBN4 a_84976_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3622 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3623 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3624 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3625 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3626 a_90816_13393# a_89010_10235# a_88856_4328# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3627 FC_top_0.AVDD FC_top_0.IREF a_n7828_n20082# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3628 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3629 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3630 a_115137_n7688# CM_p_net_1.IN CM_p_net_1.OUT6 CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3631 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3632 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3633 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3634 a_58220_n9018# CM_n_net_0.IN a_57660_n9018# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3635 a_42289_11461# PRbiased_net_x5_1.IBP1 a_36009_10235# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3636 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3637 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3638 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3639 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3640 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3641 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3642 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3643 a_29999_11461# PRbiased_net_x5_1.IBN1 a_31975_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3644 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3645 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3646 a_107077_n38276# a_106677_n40268# PRbiased_net_x5_0.IBP5 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3647 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3648 PRbiased_net_x5_1.ITN5 PRbiased_net_x5_1.IBN5 a_101239_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3649 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3650 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3651 a_90816_11461# a_89010_10235# CM_n_net_1.VSS PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3652 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3653 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3654 a_103741_n8593# CM_p_net_1.IN a_102903_n8593# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3655 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3656 a_43664_4328# a_41738_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3657 a_53676_n40268# PRbiased_net_x5_0.IBP2 a_61362_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3658 CM_n_net_1.VSS a_41738_4328# a_42260_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3659 PRbiased_net_x5_1.VDD a_83000_10295# a_83530_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3660 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3661 a_101767_n22968# CM_p_net_1.IN a_100929_n22968# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3662 a_108601_n11308# CM_p_net_1.IN a_108033_n11308# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3663 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3664 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3665 a_30529_10295# a_29999_10295# a_29999_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3666 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3667 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3668 a_65333_10295# a_65505_4268# a_67309_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3669 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X3670 FC_top_0.AVDD FC_top_0.IREF a_n7828_n21089# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3671 a_71743_n40208# a_71343_n40268# a_71213_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3672 a_2944_n20707# a_n7408_n26036# a_2376_n20707# FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X3673 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3674 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3675 a_58220_n10812# CM_n_net_0.IN a_57660_n10812# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3676 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3677 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3678 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3679 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3680 a_78998_7410# a_77072_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3681 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3682 a_115137_n10403# CM_p_net_1.IN a_114299_n10403# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3683 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3684 a_65360_n14301# CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3685 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3686 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3687 PRbiased_net_x5_1.VDD a_83000_10295# a_83530_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3688 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3689 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3690 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3691 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3692 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3693 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3694 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3695 PRbiased_net_x5_0.ITP2 a_47838_n33199# a_59956_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3696 a_89010_n40268# a_94739_n33067# a_96665_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3697 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3698 a_90782_7410# a_83000_11461# a_83172_4268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3699 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3700 a_61362_10295# PRbiased_net_x5_1.IBP2 PRbiased_net_x5_1.ITP2 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3701 a_102643_4328# PRbiased_net_x5_1.IBN5 PRbiased_net_x5_1.ITN5 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3702 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3703 a_30571_4328# a_30171_4268# a_29999_10295# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3704 a_57660_n21477# CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3705 PRbiased_net_x5_0.ITN2 a_47838_n33199# a_48238_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3706 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3707 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3708 a_114299_n20253# CM_p_net_1.IN a_113731_n20253# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3709 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3710 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3711 a_31849_n8890# CM_n_net_1.IN a_31289_n8890# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3712 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3713 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3714 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3715 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3716 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3717 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3718 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3719 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3720 CM_p_net_0.VDD CM_p_net_0.IN a_96916_n11427# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3721 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3722 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3723 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3724 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3725 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3726 a_56786_n7224# CM_n_net_0.IN a_56226_n7224# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3727 a_59094_n14301# CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3728 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3729 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3730 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3731 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3732 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3733 a_108601_n15728# CM_p_net_1.IN a_108033_n15728# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3734 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X3735 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3736 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3737 a_37815_10295# a_36009_10235# a_35855_7410# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3738 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3739 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X3740 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3741 a_59956_10295# a_47838_4268# a_59405_4328# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3742 a_42947_n15967# CM_n_net_1.IN a_42387_n15070# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3743 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3744 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3745 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X3746 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3747 a_44381_n4405# CM_n_net_1.IN a_43821_n3508# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3748 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3749 PRbiased_net_x5_0.VDD a_83000_n39042# a_83530_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3750 a_92056_n5092# CM_p_net_0.IN a_91218_n4187# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3751 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3752 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3753 PRbiased_net_x5_1.ITP2 PRbiased_net_x5_1.IBP2 a_59956_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3754 a_114607_n18443# CM_p_net_1.IN a_114299_n14823# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3755 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3756 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3757 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3758 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3759 a_114363_n38276# a_100839_n33199# PRbiased_net_x5_0.ITP5 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3760 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3761 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3762 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3763 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3764 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3765 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3766 FC_top_0.VOUT a_n7828_n21089# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3767 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3768 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3769 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3770 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3771 FC_top_0.VOUT a_n7828_n21089# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3772 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3773 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3774 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3775 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3776 a_64486_n16095# CM_n_net_0.IN a_63926_n16095# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3777 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3778 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3779 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3780 PRbiased_net_x5_1.ITP2 PRbiased_net_x5_1.IBP2 a_59956_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3781 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3782 a_97754_n5092# CM_p_net_0.IN a_96916_n5092# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3783 a_106627_n4068# CM_p_net_1.IN CM_p_net_1.OUT3 CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3784 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3785 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3786 PRbiased_net_x5_0.ITP3 a_65505_n33199# a_77623_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3787 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3788 a_97754_n16752# CM_p_net_0.IN a_96916_n15847# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3789 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3790 a_36009_10235# a_41738_4328# a_43664_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3791 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3792 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3793 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3794 a_112957_n38276# PRbiased_net_x5_0.IBP5 a_106677_n40268# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3795 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3796 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3797 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3798 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3799 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3800 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3801 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3802 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3803 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3804 a_62492_n5430# CM_n_net_0.IN a_61970_n6327# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3805 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3806 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3807 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3808 a_107465_n4973# CM_p_net_1.IN a_106627_n4973# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3809 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3810 a_64486_n5430# CM_n_net_0.IN a_63926_n5430# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3811 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3812 a_49642_n34225# a_47838_n33199# PRbiased_net_x5_0.ITN2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3813 CM_n_net_1.VSS a_59405_n33067# a_59927_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3814 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3815 a_55482_10295# a_53676_10235# a_53522_7410# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3816 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3817 a_42387_n21349# CM_n_net_1.IN a_41865_n21349# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3818 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3819 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3820 a_42387_n18658# CM_n_net_1.IN a_41865_n19555# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3821 a_101239_n33067# a_100839_n33199# a_100667_n39042# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3822 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3823 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3824 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3825 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3826 a_100667_11461# PRbiased_net_x5_1.IBN5 a_102643_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3827 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3828 PRbiased_net_x5_1.ITN1 a_30171_4268# a_30571_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3829 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3830 a_37815_n37110# a_36009_n40268# a_35855_n34225# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3831 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3832 a_36681_n21349# CM_n_net_1.IN a_36121_n21349# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3833 a_115137_n7688# CM_p_net_1.IN a_114607_n6783# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3834 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3835 a_36681_n18658# CM_n_net_1.IN a_36121_n18658# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3836 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3837 a_73115_n33067# a_65333_n40208# PRbiased_net_x5_0.IBN3 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3838 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3839 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3840 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3841 a_102603_n39042# a_100667_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3842 a_114332_6252# a_112406_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3843 a_42260_6252# a_41738_4328# a_41738_4328# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3844 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3845 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3846 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3847 PRbiased_net_x5_0.IBP4 a_89010_n40268# a_90816_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3848 a_n7828_n21089# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3849 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3850 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3851 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3852 a_33283_n6199# CM_n_net_1.IN a_32723_n6199# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3853 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3854 a_84952_n4187# CM_p_net_0.IN a_84384_n4187# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3855 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3856 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3857 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3858 a_108601_n10403# CM_p_net_1.IN a_108033_n10403# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3859 a_42387_n10684# CM_n_net_1.IN a_41865_n10684# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3860 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3861 a_42289_n39042# a_30171_n33199# a_41738_n33067# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3862 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3863 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3864 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3865 a_36409_n37110# a_36009_n40268# PRbiased_net_x5_0.VA PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3866 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3867 a_n7828_n21089# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3868 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3869 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3870 a_55448_7410# a_47666_11461# a_47838_4268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3871 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3872 a_36681_n10684# CM_n_net_1.IN a_36121_n10684# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3873 CM_p_net_1.VDD CM_p_net_1.IN a_108601_n11308# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3874 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X3875 PRbiased_net_x5_0.VDD a_65333_n39042# a_65863_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3876 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3877 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3878 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3879 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3880 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3881 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3882 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3883 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3884 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3885 a_56226_n7224# CM_n_net_0.IN CM_n_net_0.OUT4 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3886 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3887 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3888 a_95290_n40208# PRbiased_net_x5_0.IBP4 a_89010_n40268# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3889 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3890 a_86358_n7807# CM_p_net_0.IN CM_p_net_0.OUT2 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3891 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3892 a_38115_n19555# CM_n_net_1.IN a_37555_n19555# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3893 FC_top_0.AVDD FC_top_0.IREF a_n7828_n20082# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3894 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3895 a_86358_n8712# CM_p_net_0.IN a_85520_n5997# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3896 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3897 a_53388_n15198# CM_n_net_0.IN a_52828_n15198# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3898 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3899 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3900 a_102335_n5878# CM_p_net_1.IN a_101767_n5878# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3901 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3902 a_65905_n34225# PRbiased_net_x5_0.IBN3 a_65333_n40208# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3903 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3904 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3905 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3906 a_97754_n10522# CM_p_net_0.IN a_96916_n10522# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3907 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3908 a_36377_n33067# a_29999_n40208# PRbiased_net_x5_0.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3909 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3910 a_32723_n16864# CM_n_net_1.IN a_32201_n18658# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3911 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3912 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3913 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3914 CM_n_net_1.VSS a_112406_4328# a_112928_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3915 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3916 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3917 a_89410_n38276# a_89010_n40268# PRbiased_net_x5_0.IBP4 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3918 FC_top_0.AVDD FC_top_0.IREF a_n7828_n20082# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3919 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3920 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X3921 a_108601_n14823# CM_p_net_1.IN a_108033_n14823# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3922 a_62492_n14301# CM_n_net_0.IN a_61970_n15198# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3923 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3924 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3925 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3926 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3927 a_31935_n40208# a_29999_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3928 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3929 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3930 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3931 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3932 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X3933 CM_n_net_1.VSS a_59405_n33067# a_59927_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3934 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3935 a_49642_n32301# a_47838_n33199# PRbiased_net_x5_0.ITN2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3936 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3937 a_77072_4328# a_77072_4328# a_78998_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3938 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3939 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3940 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3941 a_91526_n6902# CM_p_net_0.IN a_91218_n3282# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3942 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3943 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3944 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3945 a_38989_n9787# CM_n_net_1.IN a_38467_n9787# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3946 a_109439_n16633# CM_p_net_1.IN a_108601_n15728# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3947 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3948 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3949 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3950 a_101239_n31143# a_100839_n33199# a_100667_n39042# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3951 a_72655_n15993# CM_input_0.ISBCS CM_input_0.IP2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X3952 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3953 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3954 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3955 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3956 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3957 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3958 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3959 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X3960 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3961 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3962 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3963 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3964 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3965 a_73115_n31143# a_65333_n40208# a_65505_n33199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3966 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3967 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3968 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3969 a_30529_n40208# a_29999_n39042# a_29999_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3970 a_36121_n16864# CM_n_net_1.IN a_35599_n16864# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3971 PRbiased_net_x5_0.IBP5 a_106677_n40268# a_108483_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3972 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3973 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3974 a_43821_n8890# CM_n_net_1.IN a_43299_n9787# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3975 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3976 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3977 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3978 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3979 a_49960_n15198# CM_n_net_0.IN a_49438_n15198# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3980 a_106627_n3163# CM_p_net_1.IN a_106097_n6783# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3981 a_45815_n8890# CM_n_net_1.IN a_45255_n8890# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3982 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3983 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X3984 a_59094_n7224# CM_n_net_0.IN a_58220_n5430# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3985 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X3986 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3987 CM_p_net_1.VDD CM_p_net_1.IN a_102903_n22968# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3988 a_63926_n5430# CM_n_net_0.IN a_63404_n5430# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3989 a_97224_n18562# CM_p_net_0.IN a_96916_n14942# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3990 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3991 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3992 PRbiased_net_x5_1.ITN3 PRbiased_net_x5_1.IBN3 a_65905_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X3993 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X3994 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X3995 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X3996 a_89244_n19467# CM_p_net_0.IN a_88714_n23087# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X3997 a_49960_n9018# CM_n_net_0.IN a_49438_n9018# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3998 a_73115_4328# a_65333_11461# a_65505_4268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3999 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X4000 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4001 a_30415_n15967# CM_n_net_1.IN a_29855_n15967# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4002 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4003 a_65863_10295# a_65333_10295# a_65333_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4004 a_77594_5486# a_77072_4328# a_71343_10235# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4005 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4006 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4007 CM_n_net_1.VSS a_106677_n40268# a_107077_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4008 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4009 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4010 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4011 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4012 a_29855_n16864# CM_n_net_1.IN a_29333_n16864# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4013 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4014 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4015 a_65920_n6327# CM_n_net_0.IN a_65360_n6327# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4016 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4017 a_48238_4328# a_47838_4268# a_47666_10295# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4018 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4019 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4020 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4021 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4022 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4023 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4024 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4025 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4026 a_65333_n40208# PRbiased_net_x5_0.IBN3 a_67309_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4027 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4028 CM_n_net_1.OUT11 CM_n_net_1.IN a_42387_n14173# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4029 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4030 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4031 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4032 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4033 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4034 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4035 a_65905_n32301# PRbiased_net_x5_0.IBN3 a_65333_n40208# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4036 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4037 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4038 a_31975_5486# a_30171_4268# PRbiased_net_x5_1.ITN1 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4039 a_36377_n31143# a_29999_n40208# a_35855_n31143# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4040 PRbiased_net_x5_0.IBP1 a_36009_n40268# a_37815_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4041 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4042 a_31289_n15070# CM_n_net_1.IN a_30767_n15967# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4043 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4044 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4045 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4046 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4047 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4048 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4049 a_100667_n39042# a_100839_n33199# a_102643_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4050 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X4051 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4052 a_48196_n40208# a_47666_n39042# a_47666_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4053 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4054 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4055 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4056 a_84952_n3282# CM_p_net_0.IN a_84384_n3282# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4057 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4058 CM_n_net_1.VSS CM_input_0.ISBCS a_72655_n16769# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X4059 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4060 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4061 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4062 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4063 PRbiased_net_x5_1.VDD a_100667_10295# a_101197_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4064 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4065 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4066 a_89244_n23087# CM_p_net_0.IN a_88714_n23087# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4067 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4068 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4069 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4070 a_55482_n37110# a_53676_n40268# a_53522_n34225# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4071 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4072 CM_n_net_1.VSS a_36009_n40268# a_36409_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4073 a_109439_n10403# CM_p_net_1.IN a_108601_n10403# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4074 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4075 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4076 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4077 a_90782_n33067# a_83000_n40208# PRbiased_net_x5_0.IBN4 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4078 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4079 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4080 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4081 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4082 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4083 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4084 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4085 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4086 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4087 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4088 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4089 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4090 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4091 a_62492_n4533# CM_n_net_0.IN a_61970_n4533# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4092 a_59956_n37110# a_47838_n33199# a_59405_n33067# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4093 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4094 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4095 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4096 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4097 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4098 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4099 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4100 a_86358_n7807# CM_p_net_0.IN a_85828_n6902# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4101 a_64486_n4533# CM_n_net_0.IN a_63926_n4533# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4102 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4103 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4104 a_58220_n4533# CM_n_net_0.IN a_57660_n3636# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4105 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4106 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4107 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4108 a_112406_n33067# a_100839_n33199# a_114363_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4109 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4110 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4111 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4112 a_107045_n34225# a_100667_n40208# a_106523_n34225# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4113 a_101767_n4068# CM_p_net_1.IN a_100929_n4068# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4114 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4115 a_102335_n4973# CM_p_net_1.IN a_101767_n4973# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4116 a_42387_n20452# CM_n_net_1.IN a_41865_n21349# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4117 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4118 a_42387_n17761# CM_n_net_1.IN CM_n_net_1.OUT12 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4119 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4120 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4121 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4122 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4123 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4124 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4125 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4126 a_36681_n20452# CM_n_net_1.IN a_36121_n20452# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4127 CM_n_net_1.VSS a_n7828_n20082# a_n7828_n20082# CM_n_net_1.VSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X4128 a_36681_n17761# CM_n_net_1.IN a_36121_n17761# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4129 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4130 PRbiased_net_x5_1.IBP5 a_106677_10235# a_108483_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4131 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4132 a_50520_n5430# CM_n_net_0.IN a_49960_n5430# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4133 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4134 a_108909_n18443# CM_p_net_1.IN a_108601_n14823# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4135 FC_top_0.VOUT a_n7828_n21089# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4136 PRbiased_net_x5_0.ITP5 PRbiased_net_x5_0.IBP5 a_112957_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4137 a_2376_n22018# a_n7408_n26036# a_1808_n22018# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X4138 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4139 a_35855_n31143# a_29999_n40208# a_37781_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4140 a_65333_n40208# PRbiased_net_x5_0.IBN3 a_67309_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4141 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4142 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4143 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4144 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4145 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4146 a_45815_n21349# CM_n_net_1.IN a_45255_n21349# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4147 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4148 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4149 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4150 a_45815_n19555# CM_n_net_1.IN a_45255_n18658# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4151 a_36377_4328# a_29999_11461# a_35855_4328# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4152 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4153 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4154 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4155 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4156 a_83572_n34225# PRbiased_net_x5_0.IBN4 a_83000_n40208# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4157 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4158 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4159 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4160 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4161 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4162 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4163 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4164 a_100667_n39042# a_100839_n33199# a_102643_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4165 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4166 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4167 a_106677_10235# a_112406_4328# a_114332_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4168 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4169 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4170 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4171 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4172 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4173 a_36009_n40268# PRbiased_net_x5_0.IBP1 a_43695_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4174 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X4175 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4176 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4177 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4178 a_49602_n38276# a_47666_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4179 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4180 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4181 a_89244_n19467# CM_p_net_0.IN a_88714_n18562# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4182 a_107077_10295# a_106677_10235# a_88880_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4183 CM_n_net_1.VSS a_112406_4328# a_112928_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4184 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4185 a_39549_n21349# CM_n_net_1.IN a_38989_n21349# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4186 a_52828_n9018# CM_n_net_0.IN a_52306_n9915# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4187 a_54076_n40208# a_53676_n40268# a_53546_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4188 a_39549_n19555# CM_n_net_1.IN a_38989_n18658# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4189 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4190 a_45815_n10684# CM_n_net_1.IN a_45255_n10684# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4191 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4192 a_90650_n23087# CM_p_net_0.IN a_90082_n23087# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4193 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4194 a_36009_10235# PRbiased_net_x5_1.IBP1 a_43695_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4195 a_101767_n22063# CM_p_net_1.IN a_100929_n22063# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4196 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4197 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4198 a_90782_n31143# a_83000_n40208# a_83172_n33199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4199 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4200 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4201 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4202 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4203 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4204 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4205 a_113163_n4068# CM_p_net_1.IN a_112325_n4068# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4206 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4207 a_77072_4328# a_77072_4328# a_78998_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4208 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4209 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4210 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4211 a_43821_n15967# CM_n_net_1.IN a_43299_n15967# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4212 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4213 a_31289_n5302# CM_n_net_1.IN a_30767_n5302# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4214 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4215 PRbiased_net_x5_0.ITP1 a_30171_n33199# a_42289_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4216 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4217 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4218 a_79029_n40208# a_65505_n33199# PRbiased_net_x5_0.ITP3 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4219 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4220 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4221 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X4222 FC_top_0.AVDD FC_top_0.IREF a_n7828_n21089# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4223 a_36681_n7993# CM_n_net_1.IN a_36121_n6199# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4224 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4225 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4226 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4227 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4228 a_42947_n5302# CM_n_net_1.IN a_42387_n5302# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4229 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4230 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4231 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4232 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4233 a_95261_n34225# a_94739_n33067# a_89010_n40268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4234 a_39549_n10684# CM_n_net_1.IN a_38989_n10684# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4235 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4236 a_107045_n32301# a_100667_n40208# PRbiased_net_x5_0.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4237 a_103741_n19348# CM_p_net_1.IN CM_p_net_1.OUT8 CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4238 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4239 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4240 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4241 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4242 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4243 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4244 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4245 a_79029_13393# a_65505_4268# PRbiased_net_x5_1.ITP3 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4246 a_96348_n23087# CM_p_net_0.IN a_95780_n23087# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4247 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4248 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4249 a_42289_10295# a_30171_4268# a_41738_4328# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4250 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4251 a_37555_n15967# CM_n_net_1.IN a_37033_n15967# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4252 PRbiased_net_x5_1.ITN3 PRbiased_net_x5_1.IBN3 a_65905_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4253 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4254 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4255 a_n7828_n20082# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4256 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X4257 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4258 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4259 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4260 a_77594_7410# a_77072_4328# a_71343_10235# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4261 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4262 PRbiased_net_x5_0.VDD a_29999_n40208# a_37781_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4263 a_90816_10295# a_89010_10235# a_88856_7410# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4264 a_112406_4328# a_100839_4268# a_114363_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4265 a_45815_n8890# CM_n_net_1.IN a_45255_n7993# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4266 a_89244_n22182# CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4267 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4268 a_79029_11461# a_65505_4268# PRbiased_net_x5_1.ITP3 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4269 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4270 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4271 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4272 a_63926_n4533# CM_n_net_0.IN a_63404_n5430# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4273 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4274 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4275 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4276 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4277 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4278 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4279 a_83572_n32301# PRbiased_net_x5_0.IBN4 a_83000_n40208# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4280 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4281 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4282 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4283 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4284 a_29999_n39042# a_29999_n39042# a_31935_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4285 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4286 a_51954_n19683# CM_n_net_0.IN a_51394_n19683# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4287 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4288 a_49960_n8121# CM_n_net_0.IN a_49438_n9018# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4289 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4290 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4291 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4292 a_112406_4328# a_100839_4268# a_114363_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4293 a_61362_n40208# a_47838_n33199# PRbiased_net_x5_0.ITP2 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4294 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4295 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4296 PRbiased_net_x5_1.VDD a_83000_10295# a_83530_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4297 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4298 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4299 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4300 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4301 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4302 a_31975_7410# a_30171_4268# PRbiased_net_x5_1.ITN1 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4303 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4304 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4305 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4306 a_101767_n3163# CM_p_net_1.IN a_100929_n3163# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4307 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4308 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4309 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4310 a_90082_n4187# CM_p_net_0.IN a_89244_n4187# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4311 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4312 a_89010_10235# a_94739_4328# a_96665_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4313 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4314 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4315 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4316 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4317 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4318 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X4319 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4320 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4321 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4322 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4323 a_96696_13393# a_83172_4268# PRbiased_net_x5_1.ITP4 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4324 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4325 a_37555_n8890# CM_n_net_1.IN a_37033_n9787# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4326 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4327 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4328 a_31289_n14173# CM_n_net_1.IN a_30415_n17761# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4329 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4330 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4331 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4332 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4333 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4334 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4335 a_39549_n8890# CM_n_net_1.IN a_38989_n8890# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4336 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4337 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4338 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4339 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4340 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4341 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4342 a_71343_n40268# PRbiased_net_x5_0.IBP3 a_79029_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4343 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4344 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4345 CM_n_net_0.OUT7 CM_n_net_0.IN a_49960_n14301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4346 a_95261_n32301# a_94739_n33067# a_89010_n40268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4347 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4348 a_96696_11461# a_83172_4268# PRbiased_net_x5_1.ITP4 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4349 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4350 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4351 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4352 PRbiased_net_x5_1.ITN5 a_100839_4268# a_101239_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4353 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4354 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4355 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4356 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4357 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4358 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4359 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4360 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4361 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4362 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4363 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4364 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4365 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4366 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4367 PRbiased_net_x5_1.ITN4 a_83172_4268# a_83572_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4368 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4369 CM_n_net_1.VSS a_41738_4328# a_42260_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4370 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4371 a_47666_n39042# a_47666_n39042# a_49602_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4372 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4373 a_65333_11461# PRbiased_net_x5_1.IBN3 a_67309_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4374 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4375 a_59654_n6327# CM_n_net_0.IN a_59094_n6327# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4376 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4377 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4378 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4379 a_95261_4328# a_94739_4328# a_94739_4328# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4380 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4381 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4382 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4383 CM_n_net_1.VSS a_n7828_n20082# a_n7828_n20082# CM_n_net_1.VSS nfet_03v3 ad=0.9p pd=3.05u as=1.3725p ps=5.72u w=2.25u l=2u
X4384 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4385 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4386 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4387 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4388 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4389 PRbiased_net_x5_1.ITP2 a_47838_4268# a_59956_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4390 a_78998_6252# a_77072_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4391 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4392 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4393 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4394 a_90650_n22182# CM_p_net_0.IN a_90082_n22182# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4395 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4396 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4397 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4398 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4399 a_36121_n6199# CM_n_net_1.IN a_35599_n6199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4400 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4401 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4402 a_52828_n20580# CM_n_net_0.IN a_52306_n20580# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4403 PRbiased_net_x5_0.VDD a_47666_n39042# a_48196_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4404 a_113163_n3163# CM_p_net_1.IN a_112325_n3163# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4405 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4406 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4407 a_52828_n17889# CM_n_net_0.IN a_51954_n16095# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4408 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4409 a_114299_n9498# CM_p_net_1.IN a_113731_n9498# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4410 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4411 a_90782_6252# a_83000_11461# PRbiased_net_x5_1.IBN4 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4412 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4413 a_83172_n33199# a_83000_n40208# a_89378_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4414 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4415 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4416 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4417 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4418 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4419 FC_top_0.AVDD FC_top_0.IREF a_n7828_n20082# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4420 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4421 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4422 a_65920_n16992# CM_n_net_0.IN a_65360_n16095# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4423 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4424 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4425 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4426 a_38115_n15070# CM_n_net_1.IN a_37555_n15070# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4427 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4428 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4429 a_91218_n17657# CM_p_net_0.IN a_90650_n17657# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4430 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4431 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4432 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4433 a_86358_n20372# CM_p_net_0.IN a_85520_n17657# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4434 a_50520_n5430# CM_n_net_0.IN a_49960_n4533# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4435 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4436 a_103741_n19348# CM_p_net_1.IN a_103211_n18443# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4437 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4438 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4439 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4440 a_48238_n34225# PRbiased_net_x5_0.IBN2 a_47666_n40208# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4441 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4442 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4443 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4444 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4445 a_45815_n21349# CM_n_net_1.IN a_45255_n20452# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4446 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4447 a_96348_n22182# CM_p_net_0.IN a_95780_n22182# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4448 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4449 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4450 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4451 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4452 a_86358_n5092# CM_p_net_0.IN a_85520_n5092# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4453 a_44381_n19555# CM_n_net_1.IN a_45255_n17761# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4454 a_56226_n20580# CM_n_net_0.IN a_55704_n21477# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4455 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4456 a_56226_n17889# CM_n_net_0.IN CM_n_net_0.OUT10 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4457 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4458 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4459 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4460 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4461 a_59654_n16992# CM_n_net_0.IN a_59094_n16095# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4462 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4463 a_77623_12227# a_65505_4268# a_77072_4328# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4464 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4465 a_49960_n3636# CM_n_net_0.IN a_49438_n4533# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4466 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4467 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4468 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4469 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4470 a_96696_n40208# a_83172_n33199# PRbiased_net_x5_0.ITP4 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4471 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4472 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4473 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4474 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4475 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4476 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4477 a_84936_n37110# a_83000_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4478 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4479 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4480 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4481 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4482 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4483 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4484 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4485 a_9305_n11560# a_n7828_n21089# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4486 a_45255_n5302# CM_n_net_1.IN a_44733_n5302# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4487 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4488 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4489 a_39549_n21349# CM_n_net_1.IN a_38989_n20452# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4490 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4491 a_65505_n33199# a_65333_n40208# a_71711_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4492 a_38115_n19555# CM_n_net_1.IN a_38989_n17761# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4493 a_52828_n8121# CM_n_net_0.IN a_52306_n8121# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4494 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4495 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4496 a_9305_n11560# a_n7828_n21089# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4497 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4498 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4499 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4500 PRbiased_net_x5_1.VDD a_47666_10295# a_48196_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4501 a_2944_n22018# a_n7408_n26036# a_2376_n22018# FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X4502 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4503 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4504 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4505 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4506 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4507 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4508 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4509 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4510 a_65360_n19683# CM_n_net_0.IN a_64838_n20580# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4511 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4512 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4513 a_65505_4268# a_65333_11461# a_71711_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4514 a_84936_13393# a_83000_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4515 a_91218_n21277# CM_p_net_0.IN a_90650_n21277# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4516 a_85520_n9617# CM_p_net_0.IN a_84952_n9617# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4517 a_35879_n40208# a_53676_n40268# a_55482_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4518 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4519 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4520 a_75637_n15093# CM_input_0.ISBCS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X4521 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4522 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4523 a_86358_n22182# CM_p_net_0.IN a_85520_n21277# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4524 a_33283_n16864# CM_n_net_1.IN a_32723_n15967# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4525 a_103741_n22063# CM_p_net_1.IN a_102903_n22063# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4526 a_90082_n3282# CM_p_net_0.IN a_89244_n3282# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4527 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4528 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4529 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4530 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4531 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4532 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4533 a_49642_n33067# PRbiased_net_x5_0.IBN2 PRbiased_net_x5_0.ITN2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4534 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4535 CM_n_net_1.VSS a_112406_n33067# a_112928_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4536 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4537 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4538 PRbiased_net_x5_0.IBN4 a_83000_n40208# a_89378_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4539 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4540 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4541 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4542 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4543 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4544 a_84936_11461# a_83000_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4545 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4546 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X4547 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4548 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4549 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4550 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4551 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4552 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4553 a_59094_n19683# CM_n_net_0.IN a_58572_n20580# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4554 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4555 a_52828_n10812# CM_n_net_0.IN a_50520_n10812# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4556 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4557 a_53522_n34225# a_53676_n40268# a_54076_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4558 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4559 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4560 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4561 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4562 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4563 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4564 a_59927_4328# a_59405_4328# a_59405_4328# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4565 a_48238_n32301# PRbiased_net_x5_0.IBN2 a_47666_n40208# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4566 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4567 a_44381_n8890# CM_n_net_1.IN a_43821_n8890# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4568 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4569 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4570 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4571 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4572 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4573 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4574 a_29999_10295# a_30171_4268# a_31975_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4575 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4576 a_43664_n34225# a_41738_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4577 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4578 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4579 a_63052_n21477# CM_n_net_0.IN a_62492_n21477# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4580 a_71711_4328# a_65333_11461# a_71189_4328# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4581 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4582 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4583 a_63052_n18786# CM_n_net_0.IN a_62492_n18786# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4584 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4585 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4586 a_43664_5486# a_41738_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4587 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4588 a_55448_6252# a_47666_11461# PRbiased_net_x5_1.IBN2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4589 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4590 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4591 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4592 a_77623_n38276# PRbiased_net_x5_0.IBP3 a_71343_n40268# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4593 a_56226_n10812# CM_n_net_0.IN a_55704_n10812# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4594 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4595 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4596 a_96916_n23087# CM_p_net_0.IN a_96348_n23087# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4597 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4598 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4599 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4600 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4601 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4602 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4603 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4604 a_114299_n8593# CM_p_net_1.IN a_113731_n8593# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4605 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4606 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4607 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4608 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4609 PRbiased_net_x5_0.IBN3 a_65333_n40208# a_71711_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4610 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4611 a_57660_n14301# CM_n_net_0.IN a_56786_n17889# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4612 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4613 a_90816_n37110# a_89010_n40268# a_88856_n34225# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4614 a_56786_n21477# CM_n_net_0.IN a_56226_n21477# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4615 a_31849_n4405# CM_n_net_1.IN a_31289_n4405# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4616 a_56786_n18786# CM_n_net_0.IN a_56226_n18786# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4617 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4618 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4619 a_65905_n33067# a_65505_n33199# a_65333_n39042# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4620 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4621 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4622 a_91218_n16752# CM_p_net_0.IN a_90650_n16752# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4623 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4624 a_102643_5486# a_100839_4268# PRbiased_net_x5_1.ITN5 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4625 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4626 a_30571_5486# PRbiased_net_x5_1.IBN1 a_29999_11461# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4627 a_107077_n39042# a_106677_n40268# PRbiased_net_x5_0.IBP5 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4628 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4629 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4630 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4631 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4632 a_29999_10295# a_29999_10295# a_31935_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4633 a_86358_n16752# CM_p_net_0.IN a_85520_n16752# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4634 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4635 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4636 a_53522_7410# a_53676_10235# a_54076_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4637 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4638 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4639 a_44381_n19555# CM_n_net_1.IN a_43821_n19555# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4640 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4641 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4642 a_39549_n8890# CM_n_net_1.IN a_38989_n7993# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4643 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4644 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4645 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4646 a_112325_n17538# CM_p_net_1.IN a_111795_n17538# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4647 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4648 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4649 a_49642_n31143# PRbiased_net_x5_0.IBN2 PRbiased_net_x5_0.ITN2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4650 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4651 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4652 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4653 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4654 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4655 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4656 CM_n_net_1.VSS a_112406_n33067# a_112928_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4657 a_59405_n33067# a_47838_n33199# a_61362_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4658 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4659 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4660 a_29999_10295# a_29999_10295# a_31935_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4661 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4662 CM_n_net_1.VSS a_53676_10235# a_54076_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4663 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4664 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4665 a_n10081_n11560# a_n7828_n21089# a_9305_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4666 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4667 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4668 a_52828_n3636# CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4669 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4670 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X4671 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4672 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4673 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4674 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4675 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4676 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4677 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4678 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4679 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4680 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4681 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4682 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4683 a_106523_7410# a_100667_11461# a_108449_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4684 a_30171_4268# a_29999_11461# a_36377_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4685 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4686 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4687 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4688 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4689 PRbiased_net_x5_0.ITP2 PRbiased_net_x5_0.IBP2 a_59956_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4690 a_43664_n32301# a_41738_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4691 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4692 a_96916_n5997# CM_p_net_0.IN a_96348_n5997# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4693 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4694 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4695 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4696 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4697 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4698 a_52828_n16992# CM_n_net_0.IN a_52306_n18786# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4699 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4700 a_91218_n20372# CM_p_net_0.IN a_90650_n20372# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4701 a_85520_n8712# CM_p_net_0.IN a_84952_n8712# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4702 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4703 a_86358_n20372# CM_p_net_0.IN a_85520_n20372# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4704 a_38115_n15070# CM_n_net_1.IN a_37555_n14173# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4705 PRbiased_net_x5_0.VDD a_83000_n39042# a_83530_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4706 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4707 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4708 a_83530_12227# a_83000_10295# a_83000_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4709 a_84384_n11427# CM_p_net_0.IN a_83546_n11427# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4710 a_112325_n21158# CM_p_net_1.IN a_111795_n21158# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4711 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4712 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4713 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4714 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4715 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4716 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4717 a_114363_n39042# PRbiased_net_x5_0.IBP5 PRbiased_net_x5_0.ITP5 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4718 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4719 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4720 a_30415_n7096# CM_n_net_1.IN a_29855_n7096# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4721 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4722 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4723 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4724 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4725 a_43695_n37110# PRbiased_net_x5_0.IBP1 PRbiased_net_x5_0.ITP1 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4726 a_107045_4328# a_100667_11461# a_106523_4328# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4727 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4728 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4729 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4730 a_65905_n31143# a_65505_n33199# a_65333_n39042# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4731 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4732 a_62492_n19683# CM_n_net_0.IN a_61970_n19683# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4733 a_56226_n16992# CM_n_net_0.IN a_55704_n16992# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4734 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4735 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X4736 a_75637_n17669# CM_input_0.ISBCS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X4737 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4738 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4739 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4740 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4741 a_100667_n40208# PRbiased_net_x5_0.IBN5 a_102643_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4742 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4743 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4744 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4745 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4746 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4747 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4748 a_29855_n6199# CM_n_net_1.IN a_29333_n6199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4749 PRbiased_net_x5_1.ITP4 a_83172_4268# a_95290_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4750 PRbiased_net_x5_1.IBP3 a_71343_10235# a_73149_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4751 a_112957_n39042# a_100839_n33199# a_112406_n33067# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4752 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4753 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4754 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4755 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4756 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4757 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4758 PRbiased_net_x5_0.ITP3 PRbiased_net_x5_0.IBP3 a_77623_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4759 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4760 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4761 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4762 a_51394_n9018# CM_n_net_0.IN a_50872_n9915# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4763 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4764 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4765 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4766 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4767 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4768 a_53388_n9018# CM_n_net_0.IN a_52828_n9018# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4769 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4770 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4771 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4772 a_84384_n15847# CM_p_net_0.IN a_83546_n15847# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4773 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4774 a_63052_n9915# CM_n_net_0.IN a_62492_n9018# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4775 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4776 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4777 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4778 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4779 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4780 a_114299_n22968# CM_p_net_1.IN a_113731_n22968# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4781 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4782 a_96916_n22182# CM_p_net_0.IN a_96348_n22182# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4783 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4784 a_51954_n15198# CM_n_net_0.IN a_51394_n15198# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4785 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4786 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4787 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4788 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4789 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4790 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4791 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4792 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4793 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4794 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4795 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4796 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4797 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4798 a_107045_n33067# a_100667_n40208# PRbiased_net_x5_0.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4799 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4800 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4801 PRbiased_net_x5_0.IBP4 a_89010_n40268# a_90816_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4802 a_9305_n11560# a_n7828_n21089# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4803 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4804 a_83000_n40208# a_83000_n39042# a_84936_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4805 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4806 a_9305_n11560# a_n7828_n21089# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4807 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4808 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4809 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4810 a_102603_n40208# a_100667_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4811 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4812 a_29999_10295# a_30171_4268# a_31975_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4813 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4814 a_112325_n16633# CM_p_net_1.IN a_111795_n17538# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4815 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4816 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4817 a_102335_n11308# CM_p_net_1.IN a_101767_n11308# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4818 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4819 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4820 a_43664_7410# a_41738_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4821 a_37815_n38276# a_36009_n40268# CM_n_net_1.VSS PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4822 a_38989_n5302# CM_n_net_1.IN a_38467_n5302# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4823 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4824 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4825 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4826 PRbiased_net_x5_0.VDD a_29999_n40208# a_37781_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4827 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4828 a_97754_n10522# CM_p_net_0.IN a_96916_n9617# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4829 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4830 a_42289_n40208# PRbiased_net_x5_0.IBP1 a_36009_n40268# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4831 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4832 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4833 a_64486_n21477# CM_n_net_0.IN a_63926_n20580# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4834 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4835 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4836 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4837 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4838 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4839 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4840 a_83572_n33067# a_83172_n33199# a_83000_n39042# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4841 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4842 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4843 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4844 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4845 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4846 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4847 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4848 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4849 a_94942_n17657# CM_p_net_0.IN a_94412_n17657# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4850 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4851 a_43821_n4405# CM_n_net_1.IN a_43299_n5302# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4852 a_67309_n34225# a_65505_n33199# PRbiased_net_x5_0.ITN3 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4853 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4854 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4855 a_100929_n11308# CM_p_net_1.IN a_100399_n11308# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4856 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4857 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4858 a_90082_n17657# CM_p_net_0.IN a_89244_n17657# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4859 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4860 a_100667_n40208# PRbiased_net_x5_0.IBN5 a_102643_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4861 a_36409_n38276# a_36009_n40268# PRbiased_net_x5_0.IBP1 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4862 a_51394_n21477# CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4863 a_45815_n4405# CM_n_net_1.IN a_45255_n4405# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4864 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4865 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4866 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4867 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4868 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4869 a_79029_10295# PRbiased_net_x5_1.IBP3 PRbiased_net_x5_1.ITP3 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4870 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4871 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4872 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4873 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4874 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4875 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4876 a_102643_7410# a_100839_4268# PRbiased_net_x5_1.ITN5 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4877 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4878 a_30571_7410# PRbiased_net_x5_1.IBN1 a_29999_11461# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4879 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4880 CM_n_net_1.VSS a_112406_4328# a_112928_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4881 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4882 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4883 a_89410_n39042# a_89010_n40268# PRbiased_net_x5_0.IBP4 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4884 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4885 a_102335_n15728# CM_p_net_1.IN a_101767_n15728# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4886 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4887 CM_n_net_1.VSS a_94739_4328# a_95261_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4888 a_102903_n9498# CM_p_net_1.IN a_102335_n9498# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4889 a_106677_10235# PRbiased_net_x5_1.IBP5 a_114363_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4890 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4891 a_73115_5486# a_65333_11461# PRbiased_net_x5_1.IBN3 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4892 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4893 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4894 a_102603_12227# a_100667_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4895 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4896 a_71343_10235# a_77072_4328# a_78998_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4897 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4898 a_84384_n10522# CM_p_net_0.IN a_83546_n10522# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4899 a_71189_n31143# a_71343_n40268# a_71743_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4900 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4901 a_112325_n20253# CM_p_net_1.IN a_111795_n21158# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4902 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4903 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4904 a_88856_n31143# a_83000_n40208# a_90782_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4905 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4906 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4907 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4908 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4909 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4910 a_48238_5486# PRbiased_net_x5_1.IBN2 a_47666_11461# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4911 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X4912 a_95261_n33067# a_94739_n33067# a_94739_n33067# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4913 a_107045_n31143# a_100667_n40208# a_106523_n31143# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4914 a_100929_n15728# CM_p_net_1.IN CM_p_net_1.OUT7 CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4915 PRbiased_net_x5_0.IBP5 a_106677_n40268# a_108483_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4916 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4917 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4918 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4919 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4920 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4921 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4922 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4923 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4924 a_94942_n21277# CM_p_net_0.IN a_94412_n21277# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4925 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4926 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4927 PRbiased_net_x5_1.ITN3 a_65505_4268# a_65905_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4928 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4929 a_61331_4328# a_59405_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4930 a_90082_n21277# CM_p_net_0.IN a_89244_n21277# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4931 FC_top_0.AVDD FC_top_0.IREF a_n7828_n20082# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4932 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4933 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4934 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4935 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4936 FC_top_0.AVDD FC_top_0.IREF a_n7828_n21089# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4937 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4938 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4939 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4940 a_96696_10295# PRbiased_net_x5_1.IBP4 PRbiased_net_x5_1.ITP4 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4941 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4942 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4943 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4944 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4945 a_90650_n4187# CM_p_net_0.IN a_90082_n4187# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4946 a_77594_6252# a_77072_4328# a_77072_4328# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4947 a_35855_n34225# a_29999_n40208# a_37781_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4948 CM_n_net_1.VSS a_106677_n40268# a_107077_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4949 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4950 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4951 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4952 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4953 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4954 a_84384_n14942# CM_p_net_0.IN a_83546_n14942# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4955 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4956 a_83572_n31143# a_83172_n33199# a_83000_n39042# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4957 a_32723_n7096# CM_n_net_1.IN a_31849_n5302# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4958 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4959 a_67269_n37110# a_65333_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4960 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4961 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4962 a_108033_n17538# CM_p_net_1.IN a_107465_n17538# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4963 a_67309_n32301# a_65505_n33199# PRbiased_net_x5_0.ITN3 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4964 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X4965 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4966 a_n10081_n10574# a_n7828_n21089# FC_top_0.VOUT CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4967 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4968 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4969 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4970 a_64486_n10812# CM_n_net_0.IN a_63926_n10812# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4971 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4972 a_n7828_n20082# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4973 a_n10081_n10574# a_n7828_n21089# FC_top_0.VOUT CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4974 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4975 CM_n_net_1.OUT1 CM_n_net_1.IN a_29855_n3508# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4976 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4977 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4978 a_36409_12227# a_36009_10235# PRbiased_net_x5_1.IBP1 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4979 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4980 PRbiased_net_x5_1.VDD a_29999_10295# a_30529_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4981 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4982 a_31975_6252# PRbiased_net_x5_1.IBN1 PRbiased_net_x5_1.ITN1 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4983 a_92056_n7807# CM_p_net_0.IN CM_p_net_0.OUT4 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4984 a_65360_n15198# CM_n_net_0.IN a_64838_n16095# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X4985 a_n7828_n20082# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X4986 a_58220_n10812# CM_n_net_0.IN a_57660_n9915# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X4987 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4988 FC_top_0.VOUT a_n7828_n21089# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X4989 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4990 a_92056_n8712# CM_p_net_0.IN a_91218_n5997# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4991 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X4992 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X4993 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4994 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4995 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4996 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X4997 PRbiased_net_x5_0.VA a_36009_n40268# a_37815_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X4998 a_106627_n17538# CM_p_net_1.IN a_106097_n17538# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X4999 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5000 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5001 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5002 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5003 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5004 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5005 a_102335_n10403# CM_p_net_1.IN a_101767_n10403# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5006 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5007 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5008 a_65360_n9018# CM_n_net_0.IN a_64838_n9915# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5009 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5010 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5011 a_45255_n16864# CM_n_net_1.IN a_44733_n18658# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5012 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5013 PRbiased_net_x5_0.VDD a_83000_n40208# a_90782_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5014 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5015 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5016 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5017 a_97754_n8712# CM_p_net_0.IN a_96916_n8712# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5018 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5019 a_59094_n15198# CM_n_net_0.IN a_58572_n16095# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5020 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5021 a_106627_n5878# CM_p_net_1.IN a_106097_n5878# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5022 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5023 a_95261_n31143# a_94739_n33067# a_94739_n33067# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5024 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5025 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5026 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5027 a_35855_n34225# a_36009_n40268# a_36409_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5028 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5029 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5030 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5031 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5032 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5033 a_94942_n16752# CM_p_net_0.IN a_94412_n17657# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5034 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5035 a_36377_5486# a_29999_11461# PRbiased_net_x5_1.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5036 a_100929_n10403# CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5037 a_84952_n11427# CM_p_net_0.IN a_84384_n11427# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5038 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5039 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5040 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5041 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5042 a_90082_n16752# CM_p_net_0.IN a_89244_n16752# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5043 PRbiased_net_x5_1.IBP1 a_36009_10235# a_37815_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5044 a_53388_n9018# CM_n_net_0.IN a_52828_n8121# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5045 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5046 a_63052_n8121# CM_n_net_0.IN a_62492_n8121# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5047 a_108033_n21158# CM_p_net_1.IN a_107465_n21158# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5048 PRbiased_net_x5_1.VDD a_100667_10295# a_101197_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5049 a_106677_n40268# PRbiased_net_x5_0.IBP5 a_114363_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5050 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5051 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5052 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5053 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5054 a_38989_n16864# CM_n_net_1.IN a_38467_n18658# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5055 a_55482_n38276# a_53676_n40268# CM_n_net_1.VSS PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5056 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5057 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5058 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5059 a_112406_4328# a_112406_4328# a_114332_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5060 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5061 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5062 FC_top_0.AVDD FC_top_0.IREF a_n7828_n21089# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5063 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5064 a_1808_n20707# a_n7408_n26036# a_1278_n21432# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X5065 a_102335_n14823# CM_p_net_1.IN a_101767_n14823# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5066 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5067 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5068 a_102903_n8593# CM_p_net_1.IN a_102335_n8593# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5069 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5070 a_59956_n38276# PRbiased_net_x5_0.IBP2 a_53676_n40268# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5071 a_83546_n11427# CM_p_net_0.IN a_83016_n11427# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5072 PRbiased_net_x5_1.VDD a_100667_10295# a_101197_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5073 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5074 PRbiased_net_x5_0.IBN4 a_83000_n40208# a_89378_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5075 a_106627_n21158# CM_p_net_1.IN a_106097_n21158# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5076 PRbiased_net_x5_0.ITP5 a_100839_n33199# a_112957_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5077 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5078 a_84976_n34225# a_83172_n33199# PRbiased_net_x5_0.ITN4 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5079 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5080 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5081 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5082 a_42947_n15967# CM_n_net_1.IN a_42387_n15967# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5083 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5084 a_n7828_n21089# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5085 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5086 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5087 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5088 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5089 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5090 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5091 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5092 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5093 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5094 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5095 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5096 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5097 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5098 a_73149_n37110# a_71343_n40268# a_71189_n34225# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5099 a_84952_n5997# CM_p_net_0.IN a_84384_n5997# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5100 a_100929_n14823# CM_p_net_1.IN a_100399_n18443# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5101 a_84952_n15847# CM_p_net_0.IN a_84384_n15847# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5102 a_48238_n33067# a_47838_n33199# a_47666_n39042# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5103 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5104 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5105 a_44381_n15070# CM_n_net_1.IN a_43821_n15070# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5106 a_84936_10295# a_83000_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5107 a_88880_13393# a_106677_10235# a_108483_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5108 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5109 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5110 a_56786_n9915# CM_n_net_0.IN a_56226_n9018# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5111 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5112 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5113 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5114 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5115 a_94942_n20372# CM_p_net_0.IN a_94412_n21277# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5116 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5117 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5118 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5119 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5120 a_49602_n39042# a_47666_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5121 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5122 a_42387_n7096# CM_n_net_1.IN CM_n_net_1.OUT6 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5123 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5124 CM_n_net_1.VSS a_41738_n33067# a_42260_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5125 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5126 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5127 a_90082_n20372# CM_p_net_0.IN a_89244_n20372# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5128 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5129 a_2376_n21432# a_n7408_n26036# a_1808_n21432# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X5130 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5131 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5132 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5133 a_115137_n20253# CM_p_net_1.IN a_114299_n17538# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5134 a_90650_n3282# CM_p_net_0.IN a_90082_n3282# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5135 a_50520_n20580# CM_n_net_0.IN a_49960_n19683# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5136 a_41738_n33067# a_30171_n33199# a_43695_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5137 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5138 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5139 a_83546_n15847# CM_p_net_0.IN CM_p_net_0.OUT7 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5140 PRbiased_net_x5_1.IBP5 a_106677_10235# a_108483_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5141 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5142 a_73115_7410# a_65333_11461# a_65505_4268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5143 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5144 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5145 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5146 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5147 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5148 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5149 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5150 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5151 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5152 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5153 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5154 PRbiased_net_x5_0.IBN3 a_65333_n40208# a_71711_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5155 a_102903_n11308# CM_p_net_1.IN a_102335_n11308# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5156 a_91218_n4187# CM_p_net_0.IN a_90650_n4187# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5157 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5158 a_108033_n16633# CM_p_net_1.IN a_107465_n16633# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5159 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5160 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5161 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5162 a_48238_7410# PRbiased_net_x5_1.IBN2 a_47666_11461# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5163 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5164 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5165 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5166 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5167 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5168 PRbiased_net_x5_0.ITP1 PRbiased_net_x5_0.IBP1 a_42289_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5169 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5170 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5171 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.9p pd=3.05u as=0 ps=0 w=2.25u l=2u
X5172 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X5173 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5174 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5175 a_41738_4328# a_30171_4268# a_43695_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5176 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5177 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5178 a_92056_n7807# CM_p_net_0.IN a_91526_n6902# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5179 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5180 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5181 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5182 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5183 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5184 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5185 a_96916_n5092# CM_p_net_0.IN a_96348_n5092# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5186 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5187 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5188 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5189 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5190 a_106627_n16633# CM_p_net_1.IN a_106097_n17538# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5191 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5192 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5193 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5194 CM_n_net_1.VSS a_n7828_n21089# a_n2230_n26552# CM_n_net_1.VSS nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X5195 CM_n_net_1.VSS a_112406_n33067# a_112928_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5196 a_37555_n4405# CM_n_net_1.IN a_37033_n5302# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5197 a_41738_4328# a_30171_4268# a_43695_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5198 a_83172_n33199# a_83000_n40208# a_89378_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5199 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5200 FC_top_0.AVDD FC_top_0.IREF a_n7828_n21089# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5201 a_84976_n32301# a_83172_n33199# PRbiased_net_x5_0.ITN4 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5202 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5203 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5204 CM_input_0.VDD a_71318_n10715# a_72648_n10715# CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X5205 a_94739_4328# a_94739_4328# a_96665_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5206 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5207 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5208 a_51394_n3636# CM_n_net_0.IN a_50520_n7224# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5209 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5210 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5211 CM_p_net_0.VDD CM_p_net_0.IN a_91218_n11427# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5212 a_39549_n4405# CM_n_net_1.IN a_38989_n4405# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5213 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5214 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5215 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5216 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5217 a_115137_n10403# CM_p_net_1.IN a_114299_n9498# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5218 a_53388_n4533# CM_n_net_0.IN a_52828_n3636# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5219 a_115137_n22063# CM_p_net_1.IN a_114299_n21158# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5220 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5221 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5222 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5223 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5224 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5225 a_106627_n4973# CM_p_net_1.IN a_106097_n5878# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5226 a_58220_n21477# CM_n_net_0.IN a_57660_n21477# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5227 CM_n_net_0.OUT5 CM_n_net_0.IN a_62492_n3636# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5228 a_102903_n15728# CM_p_net_1.IN a_102335_n15728# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5229 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5230 a_32723_n3508# CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5231 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5232 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5233 a_62492_n15198# CM_n_net_0.IN a_61970_n15198# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5234 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5235 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5236 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5237 a_100839_4268# a_100667_11461# a_107045_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5238 a_48238_n31143# a_47838_n33199# a_47666_n39042# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5239 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5240 a_29999_11461# a_29999_10295# a_31935_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5241 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5242 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5243 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5244 a_53522_4328# a_53676_10235# a_54076_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5245 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5246 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5247 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5248 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5249 a_84952_n10522# CM_p_net_0.IN a_84384_n10522# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5250 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5251 a_43664_n33067# a_41738_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5252 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5253 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5254 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5255 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5256 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5257 a_108033_n20253# CM_p_net_1.IN a_107465_n20253# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5258 CM_n_net_1.VSS a_41738_n33067# a_42260_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5259 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X5260 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5261 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5262 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5263 PRbiased_net_x5_1.ITN4 PRbiased_net_x5_1.IBN4 a_83572_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5264 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5265 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5266 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5267 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5268 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5269 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5270 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5271 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5272 a_95261_5486# a_94739_4328# a_89010_10235# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5273 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5274 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5275 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5276 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5277 a_95290_12227# a_83172_4268# a_94739_4328# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5278 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5279 a_83546_n10522# CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5280 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5281 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5282 a_92056_n16752# CM_p_net_0.IN a_91218_n15847# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5283 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5284 a_106627_n20253# CM_p_net_1.IN a_106097_n21158# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5285 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5286 a_65505_n33199# a_65333_n40208# a_71711_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5287 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5288 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5289 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5290 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5291 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5292 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5293 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5294 a_56226_n9018# CM_n_net_0.IN a_55704_n9018# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5295 a_114299_n22063# CM_p_net_1.IN a_113731_n22063# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5296 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5297 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5298 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5299 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5300 a_63926_n16095# CM_n_net_0.IN a_63404_n16095# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5301 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5302 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5303 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5304 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5305 a_65360_n8121# CM_n_net_0.IN a_64838_n8121# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5306 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5307 a_49602_12227# a_47666_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5308 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5309 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5310 a_77072_n33067# a_65505_n33199# a_79029_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5311 a_84952_n14942# CM_p_net_0.IN a_84384_n14942# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5312 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5313 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5314 a_36377_7410# a_29999_11461# a_35855_7410# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5315 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5316 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5317 a_32723_n21349# CM_n_net_1.IN a_30415_n21349# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5318 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5319 a_65333_n40208# a_65333_n39042# a_67269_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5320 a_32723_n18658# CM_n_net_1.IN a_32201_n18658# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5321 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5322 a_108601_n17538# CM_p_net_1.IN a_108033_n17538# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5323 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5324 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5325 FC_top_0.AVDD FC_top_0.IREF a_n7828_n20082# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5326 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5327 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5328 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5329 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5330 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5331 CM_n_net_1.VSS a_112406_n33067# a_112928_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5332 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5333 a_112406_4328# a_112406_4328# a_114332_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5334 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5335 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5336 a_115137_n16633# CM_p_net_1.IN a_114299_n16633# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5337 a_47666_n39042# a_47838_n33199# a_49642_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5338 a_108033_n9498# CM_p_net_1.IN a_107465_n9498# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5339 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5340 a_83546_n14942# CM_p_net_0.IN a_83016_n18562# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5341 a_49960_n9915# CM_n_net_0.IN a_49438_n10812# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5342 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5343 a_108601_n4068# CM_p_net_1.IN a_108033_n4068# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5344 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5345 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5346 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5347 a_32723_n10684# CM_n_net_1.IN a_30415_n10684# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5348 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5349 a_36121_n21349# CM_n_net_1.IN a_35599_n21349# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5350 a_102903_n10403# CM_p_net_1.IN a_102335_n10403# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5351 a_91218_n3282# CM_p_net_0.IN a_90650_n3282# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5352 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5353 a_101767_n5878# CM_p_net_1.IN a_100929_n5878# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5354 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5355 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5356 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5357 a_36121_n18658# CM_n_net_1.IN a_35599_n19555# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5358 a_43664_n31143# a_41738_n33067# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5359 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5360 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5361 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5362 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5363 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5364 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5365 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5366 a_97754_n20372# CM_p_net_0.IN a_96916_n17657# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5367 a_59094_n9018# CM_n_net_0.IN a_58572_n9915# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5368 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5369 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5370 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5371 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5372 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5373 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5374 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X5375 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5376 PRbiased_net_x5_1.IBN3 a_65333_11461# a_71711_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5377 a_85520_n11427# CM_p_net_0.IN a_84952_n11427# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5378 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5379 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5380 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5381 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5382 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5383 a_31289_n15967# CM_n_net_1.IN a_30767_n15967# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5384 a_57660_n19683# CM_n_net_0.IN a_57138_n20580# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5385 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5386 a_29855_n21349# CM_n_net_1.IN a_29333_n21349# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5387 a_42387_n3508# CM_n_net_1.IN a_41865_n4405# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5388 a_31849_n10684# CM_n_net_1.IN a_31289_n9787# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5389 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5390 a_95780_n4187# CM_p_net_0.IN a_94942_n4187# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5391 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5392 a_108601_n21158# CM_p_net_1.IN a_108033_n21158# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5393 a_29855_n18658# CM_n_net_1.IN a_29333_n19555# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5394 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5395 a_36121_n10684# CM_n_net_1.IN a_35599_n10684# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5396 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5397 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5398 a_44381_n15070# CM_n_net_1.IN a_43821_n14173# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5399 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5400 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5401 a_92056_n10522# CM_p_net_0.IN a_91218_n10522# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5402 a_56786_n8121# CM_n_net_0.IN a_56226_n8121# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5403 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5404 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5405 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5406 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5407 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5408 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5409 a_115137_n8593# CM_p_net_1.IN a_114299_n8593# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5410 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5411 a_115137_n20253# CM_p_net_1.IN a_114299_n20253# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5412 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5413 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5414 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5415 a_102903_n14823# CM_p_net_1.IN a_102335_n14823# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5416 a_113163_n11308# CM_p_net_1.IN a_112325_n11308# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5417 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5418 a_44381_n4405# CM_n_net_1.IN a_43821_n4405# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5419 a_71343_10235# PRbiased_net_x5_1.IBP3 a_79029_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5420 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5421 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5422 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5423 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5424 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5425 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5426 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5427 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5428 a_59927_5486# a_59405_4328# a_53676_10235# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5429 a_77623_13393# PRbiased_net_x5_1.IBP3 a_71343_10235# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5430 a_29855_n10684# CM_n_net_1.IN a_29333_n10684# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5431 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5432 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5433 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5434 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5435 CM_n_net_0.OUT11 CM_n_net_0.IN a_62492_n14301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5436 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5437 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5438 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5439 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5440 a_71213_n40208# a_71343_n40268# a_73149_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5441 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5442 a_84936_n38276# a_83000_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5443 a_113163_n5878# CM_p_net_1.IN a_112325_n5878# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5444 a_97754_n22182# CM_p_net_0.IN a_96916_n21277# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5445 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5446 a_47666_n39042# a_47838_n33199# a_49642_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5447 a_85520_n15847# CM_p_net_0.IN a_84952_n15847# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5448 a_71711_5486# a_65333_11461# PRbiased_net_x5_1.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5449 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5450 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5451 a_108483_n37110# a_106677_n40268# a_106523_n34225# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5452 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5453 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5454 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5455 a_114363_12227# PRbiased_net_x5_1.IBP5 PRbiased_net_x5_1.ITP5 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5456 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5457 a_77623_11461# PRbiased_net_x5_1.IBP3 a_71343_10235# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5458 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5459 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5460 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5461 a_65920_n21477# CM_n_net_0.IN a_65360_n20580# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5462 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5463 PRbiased_net_x5_1.VDD a_47666_10295# a_48196_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5464 a_64486_n19683# CM_n_net_0.IN a_65360_n17889# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5465 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5466 a_94739_4328# a_94739_4328# a_96665_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5467 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5468 a_91526_n18562# CM_p_net_0.IN a_91218_n14942# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5469 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5470 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5471 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5472 a_65360_n3636# CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5473 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5474 a_2944_n22018# a_n7408_n26036# a_2376_n21432# FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X5475 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5476 CM_n_net_0.OUT9 CM_n_net_0.IN a_56226_n14301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5477 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5478 a_86358_n10522# CM_p_net_0.IN a_85520_n9617# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5479 a_62492_n6327# CM_n_net_0.IN a_61970_n6327# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5480 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5481 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5482 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5483 a_113163_n15728# CM_p_net_1.IN a_112325_n15728# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5484 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5485 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5486 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5487 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5488 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5489 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X5490 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5491 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5492 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5493 a_58220_n5430# CM_n_net_0.IN a_57660_n5430# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5494 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5495 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5496 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5497 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5498 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5499 PRbiased_net_x5_1.VDD a_47666_10295# a_48196_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5500 a_29999_11461# PRbiased_net_x5_1.IBN1 a_31975_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5501 a_59654_n21477# CM_n_net_0.IN a_59094_n20580# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5502 a_42387_n19555# CM_n_net_1.IN a_41865_n19555# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5503 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5504 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5505 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5506 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5507 a_108601_n16633# CM_p_net_1.IN a_108033_n16633# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5508 a_58220_n19683# CM_n_net_0.IN a_59094_n17889# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5509 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5510 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5511 a_84976_4328# PRbiased_net_x5_1.IBN4 PRbiased_net_x5_1.ITN4 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5512 a_43664_6252# a_41738_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5513 PRbiased_net_x5_1.ITN4 PRbiased_net_x5_1.IBN4 a_83572_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5514 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5515 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5516 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5517 a_36681_n20452# CM_n_net_1.IN a_36121_n19555# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5518 a_42947_n7993# CM_n_net_1.IN a_42387_n6199# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5519 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5520 a_100929_n4068# CM_p_net_1.IN CM_p_net_1.OUT1 CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5521 a_92056_n5092# CM_p_net_0.IN a_91218_n5092# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5522 a_77623_n39042# a_65505_n33199# a_77072_n33067# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5523 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5524 a_109439_n20253# CM_p_net_1.IN a_108601_n17538# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5525 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5526 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5527 a_108033_n8593# CM_p_net_1.IN a_107465_n8593# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5528 a_95261_7410# a_94739_4328# a_89010_10235# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5529 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5530 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5531 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5532 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5533 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5534 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5535 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5536 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5537 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5538 a_52828_n9915# CM_n_net_0.IN a_52306_n9915# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5539 a_108601_n3163# CM_p_net_1.IN a_108033_n3163# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5540 a_31849_n8890# CM_n_net_1.IN a_32723_n7096# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5541 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5542 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5543 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5544 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5545 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5546 a_67309_n33067# PRbiased_net_x5_0.IBN3 PRbiased_net_x5_0.ITN3 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5547 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5548 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5549 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5550 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5551 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5552 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5553 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5554 a_101767_n4973# CM_p_net_1.IN a_100929_n4973# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5555 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5556 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5557 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5558 a_n7828_n21089# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5559 a_n10081_n11560# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5560 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5561 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5562 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5563 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5564 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5565 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5566 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5567 a_102643_6252# PRbiased_net_x5_1.IBN5 PRbiased_net_x5_1.ITN5 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5568 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5569 a_30571_6252# a_30171_4268# a_29999_10295# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5570 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5571 PRbiased_net_x5_1.VDD a_100667_11461# a_108449_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5572 PRbiased_net_x5_1.IBN1 a_29999_11461# a_36377_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5573 a_90082_n5997# CM_p_net_0.IN a_89244_n5997# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5574 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5575 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5576 a_97754_n16752# CM_p_net_0.IN a_96916_n16752# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5577 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5578 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5579 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5580 a_88856_n31143# a_89010_n40268# a_89410_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5581 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5582 PRbiased_net_x5_1.IBP4 a_89010_10235# a_90816_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5583 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5584 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X5585 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5586 a_108483_12227# a_106677_10235# CM_n_net_1.VSS PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5587 a_107077_n40208# a_106677_n40268# PRbiased_net_x5_0.VB PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5588 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5589 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5590 a_56226_n8121# CM_n_net_0.IN a_55704_n9018# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5591 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5592 CM_n_net_0.OUT3 CM_n_net_0.IN a_56226_n3636# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5593 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5594 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5595 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5596 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5597 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5598 a_85520_n10522# CM_p_net_0.IN a_84952_n10522# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5599 a_90816_n38276# a_89010_n40268# CM_n_net_1.VSS PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5600 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5601 a_109439_n4973# CM_p_net_1.IN a_108601_n4068# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5602 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5603 a_95780_n3282# CM_p_net_0.IN a_94942_n3282# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5604 a_108601_n20253# CM_p_net_1.IN a_108033_n20253# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5605 PRbiased_net_x5_0.VDD a_83000_n40208# a_90782_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5606 a_53388_n16992# CM_n_net_0.IN a_52828_n16095# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5607 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5608 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5609 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5610 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5611 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5612 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5613 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5614 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5615 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5616 a_32723_n20452# CM_n_net_1.IN a_32201_n20452# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5617 a_32723_n17761# CM_n_net_1.IN a_31849_n15967# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5618 CM_n_net_1.VSS a_89010_10235# a_89410_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5619 a_65333_11461# a_65333_10295# a_67269_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5620 a_65920_n10812# CM_n_net_0.IN a_65360_n10812# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5621 a_2376_n22743# a_n7408_n26036# a_1808_n22743# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.504p ps=2.04u w=1.2u l=2u
X5622 a_109439_n22063# CM_p_net_1.IN a_108601_n21158# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5623 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5624 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5625 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5626 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5627 a_96348_n4187# CM_p_net_0.IN a_95780_n4187# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5628 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5629 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5630 a_107045_5486# a_100667_11461# PRbiased_net_x5_1.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5631 a_112325_n4068# CM_p_net_1.IN CM_p_net_1.OUT5 CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5632 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5633 a_113163_n10403# CM_p_net_1.IN a_112325_n10403# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5634 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5635 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X5636 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5637 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5638 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5639 CM_n_net_1.VSS CM_input_0.ISBCS a_72655_n15093# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X5640 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5641 a_84952_n5092# CM_p_net_0.IN a_84384_n5092# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5642 a_43695_12227# PRbiased_net_x5_1.IBP1 PRbiased_net_x5_1.ITP1 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5643 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5644 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5645 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5646 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5647 a_59654_n10812# CM_n_net_0.IN a_59094_n10812# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5648 a_36121_n20452# CM_n_net_1.IN a_35599_n21349# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5649 a_113163_n4973# CM_p_net_1.IN a_112325_n4973# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5650 a_50520_n16095# CM_n_net_0.IN a_49960_n15198# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5651 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5652 a_97754_n20372# CM_p_net_0.IN a_96916_n20372# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5653 a_n7828_n20082# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5654 a_36121_n17761# CM_n_net_1.IN CM_n_net_1.OUT10 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5655 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5656 a_43821_n9787# CM_n_net_1.IN a_43299_n9787# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5657 a_85520_n14942# CM_p_net_0.IN a_84952_n14942# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5658 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5659 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5660 a_65505_4268# a_65333_11461# a_71711_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5661 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5662 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5663 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5664 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5665 a_n10081_n10574# a_n7828_n21089# FC_top_0.VOUT CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5666 a_95780_n11427# CM_p_net_0.IN a_94942_n11427# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5667 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5668 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5669 a_49960_n16095# CM_n_net_0.IN a_49438_n16992# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5670 a_45815_n10684# CM_n_net_1.IN a_45255_n9787# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5671 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5672 a_59094_n8121# CM_n_net_0.IN a_58572_n8121# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5673 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5674 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5675 a_67309_n31143# PRbiased_net_x5_0.IBN3 PRbiased_net_x5_0.ITN3 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5676 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5677 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5678 PRbiased_net_x5_0.VDD a_83000_n39042# a_83530_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5679 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5680 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5681 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5682 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5683 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5684 PRbiased_net_x5_0.ITN4 PRbiased_net_x5_0.IBN4 a_83572_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5685 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5686 a_103741_n4973# CM_p_net_1.IN a_102903_n4068# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5687 a_47666_11461# PRbiased_net_x5_1.IBN2 a_49642_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5688 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5689 a_89010_n40268# PRbiased_net_x5_0.IBP4 a_96696_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5690 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5691 a_30415_n18658# CM_n_net_1.IN a_29855_n16864# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5692 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5693 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5694 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5695 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5696 a_114363_n40208# a_100839_n33199# PRbiased_net_x5_0.ITP5 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5697 a_86358_n8712# CM_p_net_0.IN a_85520_n8712# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5698 PRbiased_net_x5_1.VDD a_100667_10295# a_101197_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5699 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5700 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5701 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5702 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5703 a_29855_n20452# CM_n_net_1.IN a_29333_n21349# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5704 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5705 a_113163_n14823# CM_p_net_1.IN a_112325_n14823# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5706 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5707 a_29855_n17761# CM_n_net_1.IN CM_n_net_1.OUT8 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5708 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5709 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5710 CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5711 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5712 a_83530_13393# a_83000_10295# a_83000_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5713 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5714 a_64486_n9018# CM_n_net_0.IN a_65360_n7224# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5715 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5716 a_59927_7410# a_59405_4328# a_53676_10235# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5717 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5718 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5719 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5720 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5721 PRbiased_net_x5_0.ITP4 a_83172_n33199# a_95290_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5722 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5723 a_43695_n38276# a_30171_n33199# PRbiased_net_x5_0.ITP1 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5724 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5725 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5726 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5727 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5728 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5729 a_88856_n34225# a_83000_n40208# a_90782_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5730 a_112957_n40208# PRbiased_net_x5_0.IBP5 a_106677_n40268# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5731 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5732 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5733 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5734 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5735 a_100929_n3163# CM_p_net_1.IN a_100399_n6783# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5736 a_109439_n16633# CM_p_net_1.IN a_108601_n16633# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5737 a_71711_7410# a_65333_11461# a_71189_7410# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5738 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5739 a_95780_n15847# CM_p_net_0.IN a_94942_n15847# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5740 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5741 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5742 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5743 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5744 a_83530_11461# a_83000_10295# a_83000_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5745 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5746 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X5747 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5748 a_89244_n4187# CM_p_net_0.IN CM_p_net_0.OUT3 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5749 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5750 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5751 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5752 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5753 PRbiased_net_x5_1.ITP4 PRbiased_net_x5_1.IBP4 a_95290_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5754 a_53546_13393# a_71343_10235# a_73149_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5755 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5756 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5757 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5758 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5759 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5760 a_51394_n14301# CM_n_net_0.IN a_50520_n17889# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5761 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5762 PRbiased_net_x5_1.VB a_106677_10235# a_108483_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5763 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5764 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5765 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5766 a_56226_n3636# CM_n_net_0.IN a_55704_n4533# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5767 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5768 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5769 a_65920_n16992# CM_n_net_0.IN a_65360_n16992# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5770 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5771 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5772 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5773 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5774 a_38115_n15967# CM_n_net_1.IN a_37555_n15967# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5775 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5776 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5777 PRbiased_net_x5_1.ITP4 PRbiased_net_x5_1.IBP4 a_95290_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5778 PRbiased_net_x5_1.IBP3 a_71343_10235# a_73149_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5779 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5780 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5781 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5782 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5783 a_71213_n40208# a_89010_n40268# a_90816_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5784 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5785 a_45255_n6199# CM_n_net_1.IN a_44733_n7993# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5786 a_113731_n11308# CM_p_net_1.IN a_113163_n11308# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5787 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5788 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5789 a_37815_n39042# a_36009_n40268# CM_n_net_1.VSS PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5790 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5791 a_30415_n9787# CM_n_net_1.IN a_29855_n8890# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5792 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5793 a_84976_n33067# PRbiased_net_x5_0.IBN4 PRbiased_net_x5_0.ITN4 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5794 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5795 a_108909_n6783# CM_p_net_1.IN a_108601_n3163# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5796 a_58220_n4533# CM_n_net_0.IN a_57660_n4533# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5797 CM_n_net_1.VSS a_94739_4328# a_95261_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5798 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5799 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5800 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5801 PRbiased_net_x5_0.ITN4 PRbiased_net_x5_0.IBN4 a_83572_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5802 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5803 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5804 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5805 a_83000_n39042# a_83000_n39042# a_84936_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5806 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5807 a_59654_n16992# CM_n_net_0.IN a_59094_n16992# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5808 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5809 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5810 a_109439_n20253# CM_p_net_1.IN a_108601_n20253# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5811 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5812 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5813 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5814 a_33283_n4405# CM_n_net_1.IN a_32723_n3508# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5815 a_35855_7410# a_29999_11461# a_37781_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5816 a_96348_n3282# CM_p_net_0.IN a_95780_n3282# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5817 a_36009_10235# PRbiased_net_x5_1.IBP1 a_43695_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5818 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.48p pd=2u as=0 ps=0 w=1.2u l=2u
X5819 a_112325_n3163# CM_p_net_1.IN a_111795_n6783# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5820 a_31935_12227# a_29999_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5821 a_107465_n11308# CM_p_net_1.IN a_106627_n11308# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5822 a_54076_12227# a_53676_10235# PRbiased_net_x5_1.IBP2 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5823 a_36409_n39042# a_36009_n40268# PRbiased_net_x5_0.IBP1 PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5824 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5825 a_50520_n8121# CM_n_net_0.IN a_49960_n6327# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5826 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5827 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5828 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5829 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5830 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5831 a_106523_4328# a_100667_11461# a_108449_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5832 a_30171_4268# a_29999_11461# a_36377_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5833 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5834 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5835 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5836 CM_n_net_1.VSS a_41738_n33067# a_42260_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5837 CM_input_0.VDD a_71318_n10715# a_72648_n11674# CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X5838 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5839 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5840 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5841 a_45815_n19555# CM_n_net_1.IN a_45255_n19555# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5842 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5843 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5844 a_59094_n3636# CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5845 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5846 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5847 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5848 a_61331_5486# a_59405_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5849 a_113731_n15728# CM_p_net_1.IN a_113163_n15728# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5850 a_73115_6252# a_65333_11461# PRbiased_net_x5_1.IBN3 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5851 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5852 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5853 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5854 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5855 a_49960_n5430# CM_n_net_0.IN a_49438_n6327# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5856 a_89410_n40208# a_89010_n40268# a_88880_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5857 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5858 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5859 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5860 a_95780_n10522# CM_p_net_0.IN a_94942_n10522# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5861 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5862 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5863 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5864 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5865 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5866 a_n1670_n25929# a_n7828_n21089# a_n2230_n25929# CM_n_net_1.VSS nfet_03v3 ad=0.732p pd=3.62u as=0.48p ps=2u w=1.2u l=2u
X5867 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5868 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5869 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5870 a_48238_6252# a_47838_4268# a_47666_10295# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5871 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5872 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5873 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5874 CM_n_net_1.VSS CM_input_0.ISBCS a_72655_n17669# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X5875 a_103211_n6783# CM_p_net_1.IN a_102903_n3163# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5876 a_39549_n19555# CM_n_net_1.IN a_38989_n19555# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5877 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5878 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5879 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5880 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5881 a_107465_n15728# CM_p_net_1.IN a_106627_n15728# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5882 a_107045_7410# a_100667_11461# a_106523_7410# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5883 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5884 a_1808_n22018# a_n7408_n26036# a_1278_n22743# FC_top_0.AVDD pfet_03v3 ad=0.504p pd=2.04u as=0.78p ps=3.7u w=1.2u l=2u
X5885 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5886 a_102603_13393# a_100667_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5887 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5888 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5889 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5890 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5891 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5892 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5893 a_88880_n40208# a_106677_n40268# a_108483_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5894 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5895 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5896 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5897 CM_n_net_1.VSS a_71343_n40268# a_71743_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5898 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5899 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5900 a_n7828_n20082# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X5901 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5902 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5903 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5904 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5905 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5906 a_57660_n15198# CM_n_net_0.IN a_57138_n16095# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5907 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5908 a_36681_n7096# CM_n_net_1.IN a_36121_n7096# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5909 a_84976_n31143# PRbiased_net_x5_0.IBN4 PRbiased_net_x5_0.ITN4 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5910 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5911 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5912 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5913 a_102603_11461# a_100667_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5914 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5915 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5916 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5917 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5918 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5919 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5920 a_95780_n14942# CM_p_net_0.IN a_94942_n14942# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5921 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5922 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5923 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5924 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5925 a_106523_n34225# a_106677_n40268# a_107077_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5926 a_89244_n3282# CM_p_net_0.IN a_88714_n6902# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5927 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5928 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5929 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5930 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5931 CM_n_net_1.VSS CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5932 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5933 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5934 PRbiased_net_x5_0.VDD a_29999_n39042# a_30529_n37110# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5935 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5936 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5937 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5938 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5939 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5940 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5941 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5942 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5943 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5944 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5945 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5946 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5947 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5948 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5949 CM_n_net_1.VSS a_41738_n33067# a_42260_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5950 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5951 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5952 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5953 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5954 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5955 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5956 FC_top_0.AVDD a_n7408_n26036# a_2376_n22743# FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0.504p ps=2.04u w=1.2u l=2u
X5957 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5958 FC_top_0.AVDD FC_top_0.IREF a_n7828_n21089# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5959 a_112325_n22968# CM_p_net_1.IN a_111795_n22968# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5960 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5961 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5962 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5963 a_67269_n38276# a_65333_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5964 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X5965 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5966 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5967 a_113731_n10403# CM_p_net_1.IN a_113163_n10403# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5968 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5969 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5970 CM_n_net_1.VSS a_59405_4328# a_59927_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5971 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5972 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5973 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5974 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5975 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5976 a_36409_13393# a_36009_10235# a_35879_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5977 a_75637_n15993# CM_input_0.ISBCS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X5978 PRbiased_net_x5_1.VDD a_29999_10295# a_30529_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5979 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5980 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X5981 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5982 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X5983 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5984 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5985 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X5986 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5987 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5988 a_n7828_n21089# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5989 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X5990 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5991 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.78p pd=3.7u as=0 ps=0 w=1.2u l=2u
X5992 a_36377_6252# a_29999_11461# PRbiased_net_x5_1.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5993 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X5994 a_29999_n39042# a_30171_n33199# a_31975_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X5995 a_86358_n19467# CM_p_net_0.IN CM_p_net_0.OUT8 CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X5996 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5997 a_36409_11461# a_36009_10235# PRbiased_net_x5_1.IBP1 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5998 PRbiased_net_x5_1.VDD a_29999_10295# a_30529_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X5999 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6000 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6001 a_107465_n10403# CM_p_net_1.IN a_106627_n10403# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6002 a_37555_n9787# CM_n_net_1.IN a_37033_n9787# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6003 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6004 a_42387_n15070# CM_n_net_1.IN a_41865_n15070# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6005 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6006 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6007 a_55482_n39042# a_53676_n40268# CM_n_net_1.VSS PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6008 a_39549_n10684# CM_n_net_1.IN a_38989_n9787# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6009 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6010 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6011 a_106677_10235# a_112406_4328# a_114332_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6012 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6013 a_36681_n15967# CM_n_net_1.IN a_36121_n15070# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6014 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6015 a_112406_n33067# a_100839_n33199# a_114363_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6016 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6017 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6018 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6019 a_47666_n40208# PRbiased_net_x5_0.IBN2 a_49642_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6020 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6021 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6022 a_32723_n8890# CM_n_net_1.IN a_32201_n9787# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6023 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6024 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6025 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6026 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6027 a_83000_11461# PRbiased_net_x5_1.IBN4 a_84976_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6028 a_113731_n14823# CM_p_net_1.IN a_113163_n14823# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6029 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6030 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6031 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6032 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6033 a_59956_n39042# a_47838_n33199# a_59405_n33067# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6034 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6035 a_9305_n11560# a_n7828_n21089# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X6036 a_112928_n34225# a_112406_n33067# a_106677_n40268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6037 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6038 a_52828_n5430# CM_n_net_0.IN a_52306_n5430# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6039 PRbiased_net_x5_1.VA a_36009_10235# a_37815_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6040 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6041 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6042 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6043 a_96665_4328# a_94739_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6044 CM_n_net_1.VSS a_94739_4328# a_95261_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6045 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6046 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6047 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6048 a_84384_n4187# CM_p_net_0.IN a_83546_n4187# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6049 a_58220_n9018# CM_n_net_0.IN a_59094_n7224# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6050 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6051 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6052 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6053 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6054 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6055 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6056 a_72648_n10715# a_71318_n10715# a_71318_n10715# CM_input_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X6057 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6058 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6059 PRbiased_net_x5_0.ITP5 PRbiased_net_x5_0.IBP5 a_112957_n40208# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6060 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6061 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6062 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6063 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6064 a_77623_10295# a_65505_4268# a_77072_4328# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6065 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6066 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6067 a_30415_n7993# CM_n_net_1.IN a_29855_n7993# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6068 PRbiased_net_x5_1.IBP1 a_36009_10235# a_37815_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6069 a_107465_n14823# CM_p_net_1.IN a_106627_n14823# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6070 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6071 a_36121_n7096# CM_n_net_1.IN CM_n_net_1.OUT4 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6072 a_41738_n33067# a_41738_n33067# a_43664_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6073 a_n10081_n11560# a_n7828_n21089# a_9305_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X6074 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6075 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6076 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6077 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6078 a_52828_n21477# CM_n_net_0.IN a_50520_n21477# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6079 a_91218_n23087# CM_p_net_0.IN a_90650_n23087# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6080 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6081 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6082 a_52828_n18786# CM_n_net_0.IN a_52306_n18786# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6083 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6084 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6085 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6086 CM_p_net_0.VDD CM_p_net_0.IN a_85520_n23087# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6087 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6088 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6089 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6090 a_90082_n5092# CM_p_net_0.IN a_89244_n5092# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6091 a_83572_4328# a_83172_4268# a_83000_10295# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6092 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6093 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6094 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6095 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6096 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6097 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6098 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6099 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6100 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6101 PRbiased_net_x5_1.VDD a_47666_10295# a_48196_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6102 a_61331_7410# a_59405_4328# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6103 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6104 a_73149_n38276# a_71343_n40268# CM_n_net_1.VSS PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6105 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6106 a_49602_n40208# a_47666_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6107 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6108 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6109 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6110 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6111 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6112 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X6113 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6114 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6115 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6116 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6117 a_51394_n9915# CM_n_net_0.IN a_50872_n9915# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6118 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6119 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6120 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6121 a_58220_n15198# CM_n_net_0.IN a_57660_n14301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6122 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6123 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6124 a_53388_n10812# CM_n_net_0.IN a_52828_n9915# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6125 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6126 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6127 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6128 a_29999_n39042# a_30171_n33199# a_31975_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6129 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6130 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6131 a_63052_n9915# CM_n_net_0.IN a_62492_n9915# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6132 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6133 a_56226_n21477# CM_n_net_0.IN a_55704_n21477# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6134 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6135 a_56226_n18786# CM_n_net_0.IN a_55704_n19683# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6136 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6137 a_38989_n6199# CM_n_net_1.IN a_38467_n7993# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6138 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6139 PRbiased_net_x5_1.IBN5 a_100667_11461# a_107045_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6140 a_49960_n4533# CM_n_net_0.IN a_49438_n4533# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6141 PRbiased_net_x5_1.ITP5 a_100839_4268# a_112957_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6142 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6143 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6144 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6145 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6146 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6147 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6148 a_47666_n40208# PRbiased_net_x5_0.IBN2 a_49642_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6149 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6150 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6151 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6152 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6153 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6154 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6155 a_112928_n32301# a_112406_n33067# a_106677_n40268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6156 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6157 a_9305_n11560# a_n7828_n21089# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6158 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6159 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6160 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6161 a_89010_10235# a_94739_4328# a_96665_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6162 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6163 a_71189_7410# a_65333_11461# a_73115_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6164 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6165 CM_n_net_1.OUT3 CM_n_net_1.IN a_36121_n3508# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6166 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6167 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6168 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6169 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6170 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6171 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6172 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6173 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6174 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6175 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6176 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6177 a_33283_n16864# CM_n_net_1.IN a_32723_n16864# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6178 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6179 FC_top_0.AVDD FC_top_0.IREF a_n7828_n21089# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6180 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6181 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6182 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6183 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6184 PRbiased_net_x5_1.ITN2 a_47838_4268# a_48238_4328# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6185 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6186 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6187 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6188 a_41738_n33067# a_41738_n33067# a_43664_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6189 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6190 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6191 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6192 a_86358_n19467# CM_p_net_0.IN a_85828_n18562# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6193 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6194 a_42387_n8890# CM_n_net_1.IN a_41865_n8890# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6195 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6196 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6197 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6198 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6199 a_90650_n5997# CM_p_net_0.IN a_90082_n5997# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6200 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6201 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6202 a_31849_n21349# CM_n_net_1.IN a_31289_n21349# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6203 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6204 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6205 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6206 a_112325_n19348# CM_p_net_1.IN a_111795_n22968# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6207 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6208 PRbiased_net_x5_1.ITN4 a_83172_4268# a_83572_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6209 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6210 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6211 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6212 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6213 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6214 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6215 a_95261_6252# a_94739_4328# a_94739_4328# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6216 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6217 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6218 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6219 a_44381_n10684# CM_n_net_1.IN a_43821_n9787# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6220 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6221 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6222 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6223 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6224 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6225 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6226 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6227 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6228 a_77072_n33067# a_77072_n33067# a_78998_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6229 CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD CM_input_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X6230 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6231 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6232 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6233 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6234 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6235 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6236 a_31849_n10684# CM_n_net_1.IN a_31289_n10684# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6237 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6238 a_63052_n20580# CM_n_net_0.IN a_62492_n19683# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6239 a_84384_n3282# CM_p_net_0.IN a_83546_n3282# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6240 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6241 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6242 a_96916_n9617# CM_p_net_0.IN a_96348_n9617# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6243 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6244 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6245 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6246 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6247 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6248 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6249 a_101197_12227# a_100667_10295# a_100667_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6250 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6251 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6252 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6253 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6254 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6255 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6256 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6257 a_95290_13393# PRbiased_net_x5_1.IBP4 a_89010_10235# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6258 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6259 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6260 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6261 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6262 a_91218_n22182# CM_p_net_0.IN a_90650_n22182# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6263 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6264 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6265 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6266 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6267 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6268 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6269 a_86358_n22182# CM_p_net_0.IN a_85520_n22182# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6270 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6271 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6272 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6273 a_31849_n5302# CM_n_net_1.IN a_31289_n5302# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6274 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6275 a_56786_n20580# CM_n_net_0.IN a_56226_n19683# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6276 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6277 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6278 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6279 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6280 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6281 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0 ps=0 w=2.25u l=2u
X6282 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6283 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6284 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6285 a_n10081_n10574# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6286 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6287 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6288 a_95290_11461# PRbiased_net_x5_1.IBP4 a_89010_10235# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6289 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6290 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6291 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6292 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6293 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6294 a_49602_13393# a_47666_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6295 a_42387_n14173# CM_n_net_1.IN a_41865_n15070# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6296 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6297 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6298 a_65333_n39042# a_65333_n39042# a_67269_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6299 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6300 a_108033_n22968# CM_p_net_1.IN a_107465_n22968# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6301 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6302 a_59405_n33067# a_59405_n33067# a_61331_n34225# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6303 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6304 CM_n_net_1.OUT9 CM_n_net_1.IN a_36121_n14173# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6305 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X6306 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6307 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6308 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6309 a_32723_n7993# CM_n_net_1.IN a_32201_n7993# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6310 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6311 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6312 a_83530_10295# a_83000_10295# a_83000_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6313 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6314 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6315 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6316 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6317 a_49602_11461# a_47666_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6318 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6319 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X6320 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6321 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6322 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6323 a_52828_n4533# CM_n_net_0.IN a_52306_n5430# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6324 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6325 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6326 a_45815_n15070# CM_n_net_1.IN a_45255_n15070# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6327 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6328 FC_top_0.AVDD FC_top_0.IREF a_n7828_n21089# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6329 a_36121_n3508# CM_n_net_1.IN a_35599_n4405# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6330 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6331 a_106627_n22968# CM_p_net_1.IN a_106097_n22968# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6332 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6333 PRbiased_net_x5_1.IBN3 a_65333_11461# a_71711_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6334 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6335 a_38115_n4405# CM_n_net_1.IN a_37555_n3508# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6336 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6337 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6338 a_84384_n17657# CM_p_net_0.IN a_83546_n17657# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6339 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6340 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6341 a_77072_n33067# a_77072_n33067# a_78998_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6342 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6343 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6344 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6345 a_71213_13393# a_71343_10235# a_73149_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6346 PRbiased_net_x5_0.ITN4 a_83172_n33199# a_83572_n33067# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6347 PRbiased_net_x5_1.ITP4 a_83172_4268# a_95290_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6348 a_63926_n20580# CM_n_net_0.IN a_63404_n20580# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6349 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6350 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6351 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6352 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6353 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6354 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6355 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6356 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6357 a_65360_n9915# CM_n_net_0.IN a_64838_n9915# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6358 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6359 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6360 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6361 a_39549_n15070# CM_n_net_1.IN a_38989_n15070# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6362 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6363 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6364 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6365 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6366 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.732p pd=3.62u as=0 ps=0 w=1.2u l=2u
X6367 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6368 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6369 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6370 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6371 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6372 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6373 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6374 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6375 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6376 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X6377 a_108449_4328# a_100667_11461# a_100839_4268# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6378 a_59927_6252# a_59405_4328# a_59405_4328# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6379 a_100839_4268# a_100667_11461# a_107045_7410# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6380 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6381 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6382 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6383 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6384 a_112325_n19348# CM_p_net_1.IN a_111795_n18443# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6385 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6386 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6387 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6388 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6389 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6390 a_84936_n39042# a_83000_n39042# PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6391 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6392 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6393 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6394 a_n10081_n10574# a_n7828_n21089# FC_top_0.VOUT CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6395 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6396 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6397 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6398 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6399 a_71711_6252# a_65333_11461# PRbiased_net_x5_1.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6400 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6401 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6402 a_n10081_n11560# FC_top_0.VP a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6403 a_84976_5486# a_83172_4268# PRbiased_net_x5_1.ITN4 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6404 a_45255_n21349# CM_n_net_1.IN a_42947_n21349# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6405 a_91218_n5997# CM_p_net_0.IN a_90650_n5997# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6406 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6407 a_45255_n18658# CM_n_net_1.IN a_44733_n18658# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6408 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6409 a_77072_4328# a_65505_4268# a_79029_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6410 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6411 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6412 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6413 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6414 a_113731_n9498# CM_p_net_1.IN a_113163_n9498# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6415 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6416 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6417 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6418 a_29855_n7096# CM_n_net_1.IN CM_n_net_1.OUT2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6419 a_59405_n33067# a_59405_n33067# a_61331_n32301# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6420 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6421 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6422 a_84384_n21277# CM_p_net_0.IN a_83546_n21277# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6423 a_94942_n19467# CM_p_net_0.IN a_94412_n23087# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6424 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6425 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6426 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6427 a_9305_3068# a_n7408_n26036# a_9305_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6428 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6429 a_96916_n8712# CM_p_net_0.IN a_96348_n8712# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6430 PRbiased_net_x5_0.IBP3 a_71343_n40268# a_73149_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6431 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6432 a_77072_4328# a_65505_4268# a_79029_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6433 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6434 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6435 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6436 a_108483_n38276# a_106677_n40268# CM_n_net_1.VSS PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6437 a_38989_n21349# CM_n_net_1.IN a_36681_n21349# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6438 a_114363_13393# a_100839_4268# PRbiased_net_x5_1.ITP5 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6439 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6440 a_38989_n18658# CM_n_net_1.IN a_38467_n18658# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6441 a_45255_n10684# CM_n_net_1.IN a_42947_n10684# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6442 FC_top_0.VOUT a_n7408_n26036# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6443 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6444 a_51954_n16095# CM_n_net_0.IN a_51394_n16095# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6445 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6446 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6447 a_102335_n17538# CM_p_net_1.IN a_101767_n17538# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6448 a_101197_n37110# a_100667_n39042# a_100667_n39042# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6449 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6450 a_n10081_3068# FC_top_0.VP a_n10081_n11560# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6451 a_44381_n15967# CM_n_net_1.IN a_43821_n15967# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6452 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n11560# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X6453 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6454 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6455 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6456 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6457 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6458 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6459 CM_p_net_1.VDD CM_p_net_1.IN a_114299_n22968# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6460 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6461 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6462 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6463 a_56786_n9915# CM_n_net_0.IN a_56226_n9915# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6464 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6465 PRbiased_net_x5_0.ITN4 a_83172_n33199# a_83572_n31143# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6466 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6467 a_114363_11461# a_100839_4268# PRbiased_net_x5_1.ITP5 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6468 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6469 a_112325_n22063# CM_p_net_1.IN CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6470 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6471 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6472 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6473 a_42387_n7993# CM_n_net_1.IN a_41865_n8890# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6474 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6475 a_55448_n34225# a_47666_n40208# a_47838_n33199# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6476 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6477 a_31849_n21349# CM_n_net_1.IN a_31289_n20452# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6478 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6479 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6480 a_n10081_3068# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6481 CM_n_net_1.IN CM_n_net_1.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6482 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6483 a_77623_n40208# PRbiased_net_x5_0.IBP3 a_71343_n40268# PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6484 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6485 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6486 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6487 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6488 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6489 a_38989_n10684# CM_n_net_1.IN a_36681_n10684# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6490 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6491 a_63926_n10812# CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6492 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6493 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6494 a_100929_n17538# CM_p_net_1.IN a_100399_n17538# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6495 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6496 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6497 a_102603_10295# a_100667_10295# PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6498 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6499 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6500 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6501 PRbiased_net_x5_1.VDD a_100667_11461# a_108449_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6502 PRbiased_net_x5_1.IBN1 a_29999_11461# a_36377_6252# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6503 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6504 a_94942_n23087# CM_p_net_0.IN a_94412_n23087# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6505 a_53676_10235# PRbiased_net_x5_1.IBP2 a_61362_12227# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6506 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6507 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6508 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6509 a_90082_n23087# CM_p_net_0.IN a_89244_n23087# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6510 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6511 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6512 a_64486_n21477# CM_n_net_0.IN a_63926_n21477# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6513 a_89378_4328# a_83000_11461# a_88856_4328# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6514 CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6515 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6516 a_9305_4054# a_n7408_n26036# FC_top_0.VOUT FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6517 a_43821_n5302# CM_n_net_1.IN a_43299_n5302# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6518 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6519 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6520 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6521 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6522 a_90816_n39042# a_89010_n40268# CM_n_net_1.VSS PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6523 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6524 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6525 a_45815_n6199# CM_n_net_1.IN a_45255_n5302# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6526 a_84384_n16752# CM_p_net_0.IN a_83546_n16752# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6527 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6528 a_51394_n19683# CM_n_net_0.IN a_50872_n20580# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6529 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6530 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6531 a_n7828_n20082# FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6532 a_102335_n21158# CM_p_net_1.IN a_101767_n21158# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6533 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6534 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6535 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6536 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6537 a_n7408_n26036# a_n7828_n20082# CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.3725p pd=5.72u as=0.9p ps=3.05u w=2.25u l=2u
X6538 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6539 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6540 CM_p_net_1.VDD CM_p_net_1.IN CM_p_net_1.IN CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6541 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6542 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6543 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6544 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6545 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6546 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6547 CM_n_net_1.VSS a_89010_n40268# a_89410_n38276# PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6548 a_71213_13393# a_89010_10235# a_90816_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6549 a_108483_13393# a_106677_10235# a_106523_4328# PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6550 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6551 a_107045_6252# a_100667_11461# PRbiased_net_x5_1.VDD CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6552 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6553 a_47666_10295# a_47838_4268# a_49642_5486# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6554 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6555 a_92056_n10522# CM_p_net_0.IN a_91218_n9617# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6556 a_n10081_n10574# a_n7828_n21089# FC_top_0.VOUT CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0.8p ps=2.8u w=2u l=2u
X6557 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6558 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6559 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6560 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6561 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6562 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6563 a_100929_n21158# CM_p_net_1.IN a_100399_n21158# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6564 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6565 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6566 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6567 a_106627_n19348# CM_p_net_1.IN a_106097_n22968# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6568 CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6569 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6570 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6571 PRbiased_net_x5_1.IBP4 a_89010_10235# a_90816_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6572 a_9305_3068# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6573 a_108483_11461# a_106677_10235# CM_n_net_1.VSS PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6574 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6575 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6576 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6577 a_88856_7410# a_89010_10235# a_89410_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6578 a_65333_10295# a_65333_10295# a_67269_13393# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6579 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6580 a_108601_n5878# CM_p_net_1.IN a_108033_n5878# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6581 a_114299_n4068# CM_p_net_1.IN a_113731_n4068# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6582 a_36409_10295# a_36009_10235# PRbiased_net_x5_1.VA PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6583 PRbiased_net_x5_1.VDD a_29999_10295# a_30529_10295# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6584 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6585 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6586 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6587 a_33283_n8890# CM_n_net_1.IN a_32723_n8890# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6588 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6589 CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6590 a_55448_n32301# a_47666_n40208# PRbiased_net_x5_0.IBN2 CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6591 a_51394_n5430# CM_n_net_0.IN a_50872_n5430# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6592 a_n10081_3068# FC_top_0.VN a_n10081_n10574# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6593 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6594 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6595 a_106627_n7688# CM_p_net_1.IN a_106097_n11308# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6596 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6597 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6598 a_113731_n8593# CM_p_net_1.IN a_113163_n8593# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6599 a_9305_n11560# a_n7408_n26036# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6600 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6601 a_53388_n6327# CM_n_net_0.IN a_52828_n5430# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6602 FC_top_0.AVDD a_9305_n11560# a_9305_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6603 a_45815_n15070# CM_n_net_1.IN a_45255_n14173# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6604 FC_top_0.AVDD FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6605 CM_n_net_1.VSS a_89010_10235# a_89410_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6606 a_65333_10295# a_65333_10295# a_67269_11461# PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6607 a_63052_n5430# CM_n_net_0.IN a_62492_n5430# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6608 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6609 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6610 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6611 a_84384_n20372# CM_p_net_0.IN a_83546_n20372# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6612 a_94942_n19467# CM_p_net_0.IN a_94412_n18562# CM_p_net_0.VDD pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=2u
X6613 a_43695_13393# a_30171_4268# PRbiased_net_x5_1.ITP1 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6614 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6615 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6616 a_n10081_n10574# FC_top_0.VN a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6617 CM_p_net_0.VDD CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6618 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6619 PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6620 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X6621 a_9305_4054# a_9305_n11560# FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6622 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6623 CM_p_net_0.IN CM_p_net_0.IN CM_p_net_0.VDD CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6624 CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X6625 PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD PRbiased_net_x5_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6626 a_56226_n9915# CM_n_net_0.IN a_55704_n10812# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6627 FC_top_0.AVDD FC_top_0.IREF a_n10081_3068# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6628 CM_n_net_1.VSS a_n7828_n20082# a_n10081_n10574# CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6629 FC_top_0.AVDD a_9305_n11560# a_9305_4054# FC_top_0.AVDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6630 a_95780_n5997# CM_p_net_0.IN a_94942_n5997# CM_p_net_0.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6631 a_108601_n22968# CM_p_net_1.IN a_108033_n22968# CM_p_net_1.VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6632 CM_n_net_1.VSS CM_n_net_0.IN CM_n_net_0.IN CM_n_net_1.VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X6633 a_43695_11461# a_30171_4268# PRbiased_net_x5_1.ITP1 PRbiased_net_x5_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X6634 a_53388_n21477# CM_n_net_0.IN a_52828_n20580# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6635 FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X6636 a_51954_n19683# CM_n_net_0.IN a_52828_n17889# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X6637 FC_top_0.IREF FC_top_0.IREF FC_top_0.AVDD FC_top_0.AVDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6638 a_102335_n16633# CM_p_net_1.IN a_101767_n16633# CM_p_net_1.VDD pfet_03v3 ad=0.84p pd=2.84u as=0.84p ps=2.84u w=2u l=2u
X6639 a_39549_n15070# CM_n_net_1.IN a_38989_n14173# CM_n_net_1.VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
.ends

