* Extracted by KLayout with GF180MCU LVS runset on : 30/04/2024 19:55

.SUBCKT nmos_char VS VG VD1 VD2 VD3
M$1 VS VS VS VS nfet_03v3 L=1U W=5U AS=3.05P AD=2P PS=11.22U PD=5.8U
M$2 VS VS VS VS nfet_03v3 L=1U W=5U AS=2P AD=3.05P PS=5.8U PD=11.22U
M$3 VS VS VS VS nfet_03v3 L=1U W=5U AS=3.05P AD=3.05P PS=11.22U PD=11.22U
M$4 VS VS VS VS nfet_03v3 L=1U W=5U AS=3.05P AD=2P PS=11.22U PD=5.8U
M$5 VS VS VS VS nfet_03v3 L=1U W=5U AS=2P AD=3.05P PS=5.8U PD=11.22U
M$6 VS VS VS VS nfet_03v3 L=1U W=5U AS=3.05P AD=2P PS=11.22U PD=5.8U
M$7 VD1 VG VS VS nfet_03v3 L=0.28U W=5U AS=2P AD=3.05P PS=5.8U PD=11.22U
M$8 VD2 VG VS VS nfet_03v3 L=0.5U W=5U AS=3.05P AD=3.05P PS=11.22U PD=11.22U
M$9 VS VG VD3 VS nfet_03v3 L=1U W=5U AS=3.05P AD=2P PS=11.22U PD=5.8U
M$10 VS VS VS VS nfet_03v3 L=1U W=5U AS=2P AD=3.05P PS=5.8U PD=11.22U
M$11 VS VS VS VS nfet_03v3 L=1U W=5U AS=3.05P AD=2P PS=11.22U PD=5.8U
M$12 VS VS VS VS nfet_03v3 L=1U W=5U AS=2P AD=3.05P PS=5.8U PD=11.22U
M$13 VS VS VS VS nfet_03v3 L=1U W=5U AS=3.05P AD=3.05P PS=11.22U PD=11.22U
M$14 VS VS VS VS nfet_03v3 L=1U W=5U AS=3.05P AD=2P PS=11.22U PD=5.8U
M$15 VS VS VS VS nfet_03v3 L=1U W=5U AS=2P AD=3.05P PS=5.8U PD=11.22U
.ENDS nmos_char
