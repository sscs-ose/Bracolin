* Extracted by KLayout with GF180MCU LVS runset on : 02/05/2024 18:41

.SUBCKT pmos_char VS VG VD1 VD2 VD3
M$1 VS VS VS VS pfet_03v3 L=0.92U W=5U AS=3.25P AD=2.1P PS=11.3U PD=5.84U
M$2 VS VS VS VS pfet_03v3 L=0.92U W=5U AS=2.1P AD=3.25P PS=5.84U PD=11.3U
M$3 VS VS VS VS pfet_03v3 L=0.92U W=5U AS=3.25P AD=3.25P PS=11.3U PD=11.3U
M$4 VS VS VS VS pfet_03v3 L=0.92U W=5U AS=3.25P AD=2.1P PS=11.3U PD=5.84U
M$5 VS VS VS VS pfet_03v3 L=0.92U W=5U AS=2.1P AD=3.25P PS=5.84U PD=11.3U
M$6 VS VS VS VS pfet_03v3 L=1U W=5U AS=3.25P AD=2.1P PS=11.3U PD=5.84U
M$7 VD1 VG VS VS pfet_03v3 L=0.28U W=5U AS=2.1P AD=3.25P PS=5.84U PD=11.3U
M$8 VD2 VG VS VS pfet_03v3 L=0.5U W=5U AS=3.25P AD=3.25P PS=11.3U PD=11.3U
M$9 VS VG VD3 VS pfet_03v3 L=1U W=5U AS=3.25P AD=2.1P PS=11.3U PD=5.84U
M$10 VS VS VS VS pfet_03v3 L=1U W=5U AS=2.1P AD=3.25P PS=5.84U PD=11.3U
M$11 VS VS VS VS pfet_03v3 L=0.92U W=5U AS=3.25P AD=2.1P PS=11.3U PD=5.84U
M$12 VS VS VS VS pfet_03v3 L=0.92U W=5U AS=2.1P AD=3.25P PS=5.84U PD=11.3U
M$13 VS VS VS VS pfet_03v3 L=0.92U W=5U AS=3.25P AD=3.25P PS=11.3U PD=11.3U
M$14 VS VS VS VS pfet_03v3 L=0.92U W=5U AS=3.25P AD=2.1P PS=11.3U PD=5.84U
M$15 VS VS VS VS pfet_03v3 L=0.92U W=5U AS=2.1P AD=3.25P PS=5.84U PD=11.3U
.ENDS pmos_char
