* Extracted by KLayout with GF180MCU LVS runset on : 29/04/2024 18:51

.SUBCKT SAR_logic_dac VSSD VDP VDN vocp D Valid VDDD Set CK_1 clks Reset VCM
M$1 \$8787 \$9466 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$2 \$8818 \$8787 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$3 \$8799 \$8798 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$4 \$8788 \$9472 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$5 \$8819 \$8788 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$6 \$8801 \$8800 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$7 \$8789 \$9478 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$8 \$8820 \$8789 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$9 \$8803 \$8802 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$10 \$8790 \$9484 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$11 \$8821 \$8790 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$12 \$8805 \$8804 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$13 \$8791 \$9490 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$14 \$8822 \$8791 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$15 \$8807 \$8806 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$16 \$8792 \$9496 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$17 \$8823 \$8792 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$18 \$8809 \$8808 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$19 \$8793 \$9502 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$20 \$8824 \$8793 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$21 \$8811 \$8810 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$22 \$8794 \$9508 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$23 \$8825 \$8794 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$24 \$8813 \$8812 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$25 \$8795 \$9514 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$26 \$8826 \$8795 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$27 \$8815 \$8814 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$28 \$8796 \$9520 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$29 \$8827 \$8796 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$30 \$8817 \$8816 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$31 \$1278 \$8818 \$1263 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$32 \$8798 \$8787 \$1263 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$33 \$1278 \$8787 \$8799 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$34 \$1280 \$8819 \$1265 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$35 \$8800 \$8788 \$1265 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$36 \$1280 \$8788 \$8801 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$37 \$1282 \$8820 \$1267 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$38 \$8802 \$8789 \$1267 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$39 \$1282 \$8789 \$8803 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$40 \$2940 \$8821 \$2938 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$41 \$8804 \$8790 \$2938 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$42 \$2940 \$8790 \$8805 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$43 \$5832 \$8822 \$5830 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$44 \$8806 \$8791 \$5830 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$45 \$5832 \$8791 \$8807 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$46 \$1286 \$8823 \$1271 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$47 \$8808 \$8792 \$1271 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$48 \$1286 \$8792 \$8809 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$49 \$1289 \$8824 \$1274 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$50 \$8810 \$8793 \$1274 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$51 \$1289 \$8793 \$8811 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$52 \$1290 \$8825 \$1275 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$53 \$8812 \$8794 \$1275 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$54 \$1290 \$8794 \$8813 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$55 \$2941 \$8826 \$2939 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$56 \$8814 \$8795 \$2939 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$57 \$2941 \$8795 \$8815 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$58 \$5833 \$8827 \$5831 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$59 \$8816 \$8796 \$5831 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$60 \$5833 \$8796 \$8817 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$61 \$9527 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$62 \$9528 \$9527 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$63 \$9461 \$9528 D VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$64 \$10346 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$65 \$9462 \$9461 \$10346 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$66 \$10347 \$9462 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$67 \$9463 clks \$10347 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$68 \$9461 \$9527 \$9463 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$69 \$9465 \$9527 \$9462 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$70 \$10348 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$71 \$9466 \$9465 \$10348 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$72 \$10349 \$9466 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$73 \$9464 Set \$10349 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$74 \$9465 \$9528 \$9464 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$75 \$9529 \$9466 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$76 \$9530 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$77 \$9531 \$9530 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$78 \$9467 \$9531 \$9466 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$79 \$10350 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$80 \$9468 \$9467 \$10350 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$81 \$10351 \$9468 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$82 \$9469 clks \$10351 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$83 \$9467 \$9530 \$9469 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$84 \$9471 \$9530 \$9468 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$85 \$10352 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$86 \$9472 \$9471 \$10352 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$87 \$10353 \$9472 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$88 \$9470 Set \$10353 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$89 \$9471 \$9531 \$9470 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$90 \$9532 \$9472 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$91 \$9533 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$92 \$9534 \$9533 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$93 \$9473 \$9534 \$9472 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$94 \$10354 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$95 \$9474 \$9473 \$10354 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$96 \$10355 \$9474 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$97 \$9475 clks \$10355 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$98 \$9473 \$9533 \$9475 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$99 \$9477 \$9533 \$9474 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$100 \$10356 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$101 \$9478 \$9477 \$10356 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$102 \$10357 \$9478 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$103 \$9476 Set \$10357 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$104 \$9477 \$9534 \$9476 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$105 \$9535 \$9478 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$106 \$9536 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$107 \$9537 \$9536 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$108 \$9479 \$9537 \$9478 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$109 \$10358 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$110 \$9480 \$9479 \$10358 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$111 \$10359 \$9480 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$112 \$9481 clks \$10359 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$113 \$9479 \$9536 \$9481 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$114 \$9483 \$9536 \$9480 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$115 \$10360 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$116 \$9484 \$9483 \$10360 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$117 \$10361 \$9484 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$118 \$9482 Set \$10361 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$119 \$9483 \$9537 \$9482 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$120 \$9538 \$9484 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$121 \$9539 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$122 \$9540 \$9539 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$123 \$9485 \$9540 \$9484 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$124 \$10362 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$125 \$9486 \$9485 \$10362 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$126 \$10363 \$9486 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$127 \$9487 clks \$10363 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$128 \$9485 \$9539 \$9487 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$129 \$9489 \$9539 \$9486 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$130 \$10364 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$131 \$9490 \$9489 \$10364 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$132 \$10365 \$9490 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$133 \$9488 Set \$10365 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$134 \$9489 \$9540 \$9488 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$135 \$9541 \$9490 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$136 \$9542 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$137 \$9543 \$9542 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$138 \$9491 \$9543 \$9490 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$139 \$10366 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$140 \$9492 \$9491 \$10366 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$141 \$10367 \$9492 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$142 \$9493 clks \$10367 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$143 \$9491 \$9542 \$9493 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$144 \$9495 \$9542 \$9492 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$145 \$10368 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$146 \$9496 \$9495 \$10368 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$147 \$10369 \$9496 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$148 \$9494 Set \$10369 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$149 \$9495 \$9543 \$9494 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$150 \$9544 \$9496 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$151 \$9545 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$152 \$9546 \$9545 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$153 \$9497 \$9546 \$9496 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$154 \$10370 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$155 \$9498 \$9497 \$10370 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$156 \$10371 \$9498 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$157 \$9499 clks \$10371 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$158 \$9497 \$9545 \$9499 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$159 \$9501 \$9545 \$9498 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$160 \$10372 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$161 \$9502 \$9501 \$10372 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$162 \$10373 \$9502 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$163 \$9500 Set \$10373 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$164 \$9501 \$9546 \$9500 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$165 \$9547 \$9502 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$166 \$9548 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$167 \$9549 \$9548 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$168 \$9503 \$9549 \$9502 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$169 \$10374 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$170 \$9504 \$9503 \$10374 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$171 \$10375 \$9504 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$172 \$9505 clks \$10375 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$173 \$9503 \$9548 \$9505 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$174 \$9507 \$9548 \$9504 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$175 \$10376 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$176 \$9508 \$9507 \$10376 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$177 \$10377 \$9508 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$178 \$9506 Set \$10377 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$179 \$9507 \$9549 \$9506 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$180 \$9550 \$9508 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$181 \$9551 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$182 \$9552 \$9551 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$183 \$9509 \$9552 \$9508 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$184 \$10378 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$185 \$9510 \$9509 \$10378 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$186 \$10379 \$9510 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$187 \$9511 clks \$10379 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$188 \$9509 \$9551 \$9511 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$189 \$9513 \$9551 \$9510 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$190 \$10380 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$191 \$9514 \$9513 \$10380 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$192 \$10381 \$9514 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$193 \$9512 Set \$10381 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$194 \$9513 \$9552 \$9512 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$195 \$9553 \$9514 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$196 \$9554 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$197 \$9555 \$9554 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$198 \$9515 \$9555 \$9514 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$199 \$10382 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$200 \$9516 \$9515 \$10382 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$201 \$10383 \$9516 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$202 \$9517 clks \$10383 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$203 \$9515 \$9554 \$9517 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$204 \$9519 \$9554 \$9516 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$205 \$10384 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$206 \$9520 \$9519 \$10384 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$207 \$10385 \$9520 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$208 \$9518 Set \$10385 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$209 \$9519 \$9555 \$9518 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$210 \$9556 \$9520 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$211 \$9557 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$212 \$9558 \$9557 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$213 \$9521 \$9558 \$9520 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$214 \$10386 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$215 \$9522 \$9521 \$10386 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$216 \$10387 \$9522 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$217 \$9523 clks \$10387 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$218 \$9521 \$9557 \$9523 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$219 \$9526 \$9557 \$9522 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$220 \$10388 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$221 CK_1 \$9526 \$10388 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$222 \$10389 CK_1 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$223 \$9525 Set \$10389 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$224 \$9526 \$9558 \$9525 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$225 \$9559 CK_1 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$226 \$10972 \$11176 \$10973 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$227 VDDD \$10973 \$11809 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$228 \$11016 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$229 \$11017 \$11016 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$230 \$11792 \$11811 \$11747 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$231 \$12323 Set \$11792 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$232 \$10974 \$11017 \$10973 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$233 VDDD \$10973 \$12323 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$234 \$11392 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$235 \$10975 \$10974 \$11392 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$236 \$12324 \$11747 \$10973 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$237 VDDD Reset \$12324 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$238 \$11393 \$10975 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$239 \$10976 Reset \$11393 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$240 \$11793 \$11810 \$11747 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$241 \$10974 \$11016 \$10976 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$242 \$11794 \$11810 \$11782 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$243 \$10979 \$11016 \$10975 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$244 \$12325 Reset \$11794 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$245 VDDD \$11793 \$12325 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$246 \$11394 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$247 \$10977 \$10979 \$11394 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$248 \$12326 \$11782 \$11793 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$249 VDDD Set \$12326 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$250 \$11395 \$10977 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$251 vocp \$11811 \$11782 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$252 \$10978 Set \$11395 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$253 \$10979 \$11017 \$10978 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$254 VDDD \$11810 \$11811 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$255 VDDD \$11015 \$11810 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$256 \$11018 \$10977 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$257 VDDD \$11176 \$11015 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$258 VDDD CK_1 \$11176 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$259 \$10970 \$11190 \$10980 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$260 VDDD \$10980 \$11813 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$261 \$11020 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$262 \$11021 \$11020 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$263 \$11795 \$11815 \$11748 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$264 \$12327 Set \$11795 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$265 \$10981 \$11021 \$10980 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$266 VDDD \$10980 \$12327 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$267 \$11396 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$268 \$10982 \$10981 \$11396 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$269 \$12328 \$11748 \$10980 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$270 VDDD Reset \$12328 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$271 \$11397 \$10982 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$272 \$10983 Reset \$11397 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$273 \$11796 \$11814 \$11748 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$274 \$10981 \$11020 \$10983 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$275 \$11797 \$11814 \$11783 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$276 \$10986 \$11020 \$10982 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$277 \$12329 Reset \$11797 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$278 VDDD \$11796 \$12329 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$279 \$11398 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$280 \$10984 \$10986 \$11398 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$281 \$12330 \$11783 \$11796 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$282 VDDD Set \$12330 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$283 \$11399 \$10984 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$284 vocp \$11815 \$11783 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$285 \$10985 Set \$11399 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$286 \$10986 \$11021 \$10985 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$287 VDDD \$11814 \$11815 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$288 VDDD \$11019 \$11814 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$289 \$11022 \$10984 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$290 VDDD \$11190 \$11019 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$291 VDDD \$9520 \$11190 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$292 \$10987 \$11203 \$10988 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$293 VDDD \$10988 \$11817 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$294 \$11024 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$295 \$11025 \$11024 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$296 \$11798 \$11819 \$11749 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$297 \$12331 Set \$11798 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$298 \$10989 \$11025 \$10988 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$299 VDDD \$10988 \$12331 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$300 \$11400 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$301 \$10990 \$10989 \$11400 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$302 \$12332 \$11749 \$10988 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$303 VDDD Reset \$12332 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$304 \$11401 \$10990 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$305 \$10991 Reset \$11401 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$306 \$11799 \$11818 \$11749 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$307 \$10989 \$11024 \$10991 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$308 \$11800 \$11818 \$11784 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$309 \$10994 \$11024 \$10990 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$310 \$12333 Reset \$11800 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$311 VDDD \$11799 \$12333 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$312 \$11402 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$313 \$10992 \$10994 \$11402 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$314 \$12334 \$11784 \$11799 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$315 VDDD Set \$12334 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$316 \$11403 \$10992 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$317 vocp \$11819 \$11784 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$318 \$10993 Set \$11403 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$319 \$10994 \$11025 \$10993 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$320 VDDD \$11818 \$11819 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$321 VDDD \$11023 \$11818 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$322 \$11026 \$10992 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$323 VDDD \$11203 \$11023 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$324 VDDD \$9514 \$11203 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$325 \$10971 \$11216 \$10995 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$326 VDDD \$10995 \$11821 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$327 \$11028 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$328 \$11029 \$11028 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$329 \$11801 \$11823 \$11750 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$330 \$12335 Set \$11801 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$331 \$10996 \$11029 \$10995 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$332 VDDD \$10995 \$12335 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$333 \$11404 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$334 \$10997 \$10996 \$11404 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$335 \$12336 \$11750 \$10995 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$336 VDDD Reset \$12336 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$337 \$11405 \$10997 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$338 \$10998 Reset \$11405 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$339 \$11802 \$11822 \$11750 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$340 \$10996 \$11028 \$10998 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$341 \$11803 \$11822 \$11785 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$342 \$11001 \$11028 \$10997 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$343 \$12337 Reset \$11803 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$344 VDDD \$11802 \$12337 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$345 \$11406 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$346 \$10999 \$11001 \$11406 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$347 \$12338 \$11785 \$11802 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$348 VDDD Set \$12338 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$349 \$11407 \$10999 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$350 vocp \$11823 \$11785 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$351 \$11000 Set \$11407 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$352 \$11001 \$11029 \$11000 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$353 VDDD \$11822 \$11823 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$354 VDDD \$11027 \$11822 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$355 \$11030 \$10999 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$356 VDDD \$11216 \$11027 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$357 VDDD \$9508 \$11216 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$358 \$11002 \$11229 \$11003 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$359 VDDD \$11003 \$11825 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$360 \$11032 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$361 \$11033 \$11032 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$362 \$11804 \$11827 \$11751 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$363 \$12339 Set \$11804 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$364 \$11004 \$11033 \$11003 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$365 VDDD \$11003 \$12339 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$366 \$11408 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$367 \$11005 \$11004 \$11408 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$368 \$12340 \$11751 \$11003 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$369 VDDD Reset \$12340 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$370 \$11409 \$11005 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$371 \$11006 Reset \$11409 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$372 \$11805 \$11826 \$11751 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$373 \$11004 \$11032 \$11006 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$374 \$11806 \$11826 \$11786 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$375 \$11009 \$11032 \$11005 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$376 \$12341 Reset \$11806 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$377 VDDD \$11805 \$12341 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$378 \$11410 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$379 \$11007 \$11009 \$11410 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$380 \$12342 \$11786 \$11805 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$381 VDDD Set \$12342 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$382 \$11411 \$11007 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$383 vocp \$11827 \$11786 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$384 \$11008 Set \$11411 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$385 \$11009 \$11033 \$11008 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$386 VDDD \$11826 \$11827 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$387 VDDD \$11031 \$11826 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$388 \$11034 \$11007 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$389 VDDD \$11229 \$11031 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$390 VDDD \$9502 \$11229 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$391 VDDD \$12776 \$12774 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$392 \$12743 \$12968 \$12698 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$393 \$13225 Set \$12743 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$394 VDDD \$12776 \$13225 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$395 \$13226 \$12698 \$12776 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$396 VDDD Reset \$13226 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$397 \$12744 \$12775 \$12698 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$398 \$12745 \$12775 \$12732 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$399 \$13227 Reset \$12745 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$400 VDDD \$12744 \$13227 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$401 \$13228 \$12732 \$12744 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$402 VDDD Set \$13228 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$403 \$12746 \$12968 \$12732 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$404 VDDD \$12775 \$12968 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$405 VDDD clks \$12775 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$406 \$12746 \$12777 \$12733 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$407 \$9382 \$11015 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$408 VDDD \$11808 \$9382 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$409 \$11808 \$11176 \$10973 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$410 VDDD \$12780 \$12778 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$411 VDDD \$11015 \$11808 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$412 \$12747 \$12982 \$12699 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$413 \$13229 Set \$12747 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$414 VDDD \$12780 \$13229 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$415 \$13230 \$12699 \$12780 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$416 VDDD Reset \$13230 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$417 \$12748 \$12779 \$12699 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$418 \$12749 \$12779 \$12734 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$419 \$13231 Reset \$12749 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$420 VDDD \$12748 \$13231 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$421 \$13232 \$12734 \$12748 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$422 VDDD Set \$13232 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$423 \$12750 \$12982 \$12734 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$424 VDDD \$12779 \$12982 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$425 VDDD clks \$12779 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$426 \$12750 \$12781 \$12735 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$427 \$5831 \$11019 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$428 VDDD \$11812 \$5831 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$429 \$11812 \$11190 \$10980 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$430 VDDD \$12784 \$12782 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$431 VDDD \$11019 \$11812 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$432 \$12751 \$13004 \$12700 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$433 \$13233 Set \$12751 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$434 VDDD \$12784 \$13233 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$435 \$13234 \$12700 \$12784 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$436 VDDD Reset \$13234 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$437 \$12752 \$12783 \$12700 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$438 \$12753 \$12783 \$12736 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$439 \$13235 Reset \$12753 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$440 VDDD \$12752 \$13235 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$441 \$13236 \$12736 \$12752 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$442 VDDD Set \$13236 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$443 \$12754 \$13004 \$12736 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$444 VDDD \$12783 \$13004 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$445 VDDD clks \$12783 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$446 \$12754 \$12785 \$12755 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$447 \$2939 \$11023 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$448 VDDD \$11816 \$2939 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$449 \$11816 \$11203 \$10988 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$450 VDDD \$12788 \$12786 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$451 VDDD \$11023 \$11816 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$452 \$12756 \$13010 \$12701 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$453 \$13237 Set \$12756 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$454 VDDD \$12788 \$13237 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$455 \$13238 \$12701 \$12788 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$456 VDDD Reset \$13238 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$457 \$12757 \$12787 \$12701 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$458 \$12758 \$12787 \$12737 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$459 \$13239 Reset \$12758 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$460 VDDD \$12757 \$13239 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$461 \$13240 \$12737 \$12757 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$462 VDDD Set \$13240 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$463 \$12759 \$13010 \$12737 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$464 VDDD \$12787 \$13010 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$465 VDDD clks \$12787 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$466 \$12759 \$12789 \$12738 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$467 \$1275 \$11027 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$468 VDDD \$11820 \$1275 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$469 \$11820 \$11216 \$10995 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$470 VDDD \$12792 \$12790 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$471 VDDD \$11027 \$11820 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$472 \$12760 \$13024 \$12702 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$473 \$13241 Set \$12760 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$474 VDDD \$12792 \$13241 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$475 \$13242 \$12702 \$12792 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$476 VDDD Reset \$13242 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$477 \$12761 \$12791 \$12702 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$478 \$12762 \$12791 \$12739 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$479 \$13243 Reset \$12762 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$480 VDDD \$12761 \$13243 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$481 \$13244 \$12739 \$12761 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$482 VDDD Set \$13244 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$483 \$12763 \$13024 \$12739 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$484 VDDD \$12791 \$13024 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$485 VDDD clks \$12791 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$486 \$12763 \$12793 \$12740 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$487 \$1274 \$11031 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$488 VDDD \$11824 \$1274 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$489 \$11824 \$11229 \$11003 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$490 VDDD \$12796 \$12794 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$491 VDDD \$11031 \$11824 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$492 \$12764 \$13046 \$12703 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$493 \$13245 Set \$12764 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$494 VDDD \$12796 \$13245 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$495 \$13246 \$12703 \$12796 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$496 VDDD Reset \$13246 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$497 \$12765 \$12795 \$12703 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$498 \$12766 \$12795 \$12741 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$499 \$13247 Reset \$12766 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$500 VDDD \$12765 \$13247 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$501 \$13248 \$12741 \$12765 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$502 VDDD Set \$13248 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$503 \$12767 \$13046 \$12741 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$504 VDDD \$12795 \$13046 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$505 VDDD clks \$12795 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$506 \$12767 \$12797 \$12742 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$507 \$12777 \$9466 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$508 \$12977 \$12777 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$509 \$13735 \$12977 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$510 \$13879 \$13735 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$511 \$13705 \$13879 vocp VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$512 \$14359 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$513 \$13706 \$13705 \$14359 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$514 \$14360 \$13706 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$515 \$13707 Reset \$14360 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$516 \$13705 \$13735 \$13707 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$517 \$13709 \$13735 \$13706 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$518 \$14361 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$519 \$12746 \$13709 \$14361 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$520 \$14362 \$12746 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$521 \$13708 Set \$14362 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$522 \$13709 \$13879 \$13708 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$523 \$13736 \$12746 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$524 \$12781 \$9472 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$525 \$12991 \$12781 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$526 \$13738 \$12991 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$527 \$13880 \$13738 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$528 \$13710 \$13880 vocp VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$529 \$14363 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$530 \$13711 \$13710 \$14363 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$531 \$14364 \$13711 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$532 \$13712 Reset \$14364 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$533 \$13710 \$13738 \$13712 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$534 \$13714 \$13738 \$13711 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$535 \$14365 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$536 \$12750 \$13714 \$14365 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$537 \$14366 \$12750 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$538 \$13713 Set \$14366 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$539 \$13714 \$13880 \$13713 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$540 \$13739 \$12750 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$541 \$12785 \$9478 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$542 \$13005 \$12785 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$543 \$13741 \$13005 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$544 \$13881 \$13741 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$545 \$13715 \$13881 vocp VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$546 \$14367 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$547 \$13716 \$13715 \$14367 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$548 \$14368 \$13716 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$549 \$13717 Reset \$14368 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$550 \$13715 \$13741 \$13717 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$551 \$13719 \$13741 \$13716 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$552 \$14369 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$553 \$12754 \$13719 \$14369 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$554 \$14370 \$12754 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$555 \$13718 Set \$14370 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$556 \$13719 \$13881 \$13718 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$557 \$13742 \$12754 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$558 \$12789 \$9484 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$559 \$13019 \$12789 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$560 \$13744 \$13019 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$561 \$13882 \$13744 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$562 \$13720 \$13882 vocp VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$563 \$14371 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$564 \$13721 \$13720 \$14371 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$565 \$14372 \$13721 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$566 \$13722 Reset \$14372 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$567 \$13720 \$13744 \$13722 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$568 \$13724 \$13744 \$13721 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$569 \$14373 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$570 \$12759 \$13724 \$14373 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$571 \$14374 \$12759 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$572 \$13723 Set \$14374 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$573 \$13724 \$13882 \$13723 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$574 \$13745 \$12759 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$575 \$12793 \$9490 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$576 \$13033 \$12793 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$577 \$13747 \$13033 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$578 \$13883 \$13747 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$579 \$13725 \$13883 vocp VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$580 \$14375 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$581 \$13726 \$13725 \$14375 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$582 \$14376 \$13726 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$583 \$13727 Reset \$14376 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$584 \$13725 \$13747 \$13727 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$585 \$13729 \$13747 \$13726 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$586 \$14377 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$587 \$12763 \$13729 \$14377 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$588 \$14378 \$12763 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$589 \$13728 Set \$14378 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$590 \$13729 \$13883 \$13728 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$591 \$13748 \$12763 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$592 \$12797 \$9496 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$593 \$13047 \$12797 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$594 \$13750 \$13047 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$595 \$13884 \$13750 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$596 \$13730 \$13884 vocp VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$597 \$14379 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$598 \$13731 \$13730 \$14379 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$599 \$14380 \$13731 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$600 \$13732 Reset \$14380 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$601 \$13730 \$13750 \$13732 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$602 \$13734 \$13750 \$13731 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$603 \$14381 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$604 \$12767 \$13734 \$14381 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$605 \$14382 \$12767 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$606 \$13733 Set \$14382 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$607 \$13734 \$13884 \$13733 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$608 \$13751 \$12767 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$609 \$13737 \$12977 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$610 \$12746 \$12777 \$13737 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$611 \$1263 \$13737 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$612 VCM \$12977 \$1263 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$613 \$13740 \$12991 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$614 \$12750 \$12781 \$13740 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$615 \$1265 \$13740 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$616 VCM \$12991 \$1265 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$617 \$13743 \$13005 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$618 \$12754 \$12785 \$13743 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$619 \$1267 \$13743 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$620 VCM \$13005 \$1267 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$621 \$13746 \$13019 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$622 \$12759 \$12789 \$13746 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$623 \$2938 \$13746 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$624 VCM \$13019 \$2938 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$625 \$13749 \$13033 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$626 \$12763 \$12793 \$13749 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$627 \$5830 \$13749 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$628 VCM \$13033 \$5830 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$629 \$13752 \$13047 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$630 \$12767 \$12797 \$13752 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$631 \$1271 \$13752 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$632 VCM \$13047 \$1271 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$633 \$1278 \$8787 \$1263 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$634 \$8798 \$8818 \$1263 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$635 \$1278 \$8818 \$8799 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$636 \$1280 \$8788 \$1265 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$637 \$8800 \$8819 \$1265 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$638 \$1280 \$8819 \$8801 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$639 \$1282 \$8789 \$1267 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$640 \$8802 \$8820 \$1267 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$641 \$1282 \$8820 \$8803 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$642 \$2940 \$8790 \$2938 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$643 \$8804 \$8821 \$2938 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$644 \$2940 \$8821 \$8805 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$645 \$5832 \$8791 \$5830 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$646 \$8806 \$8822 \$5830 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$647 \$5832 \$8822 \$8807 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$648 \$1286 \$8792 \$1271 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$649 \$8808 \$8823 \$1271 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$650 \$1286 \$8823 \$8809 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$651 \$1289 \$8793 \$1274 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$652 \$8810 \$8824 \$1274 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$653 \$1289 \$8824 \$8811 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$654 \$1290 \$8794 \$1275 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$655 \$8812 \$8825 \$1275 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$656 \$1290 \$8825 \$8813 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$657 \$2941 \$8795 \$2939 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$658 \$8814 \$8826 \$2939 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$659 \$2941 \$8826 \$8815 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$660 \$5833 \$8796 \$5831 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$661 \$8816 \$8827 \$5831 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$662 \$5833 \$8827 \$8817 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$663 \$8787 \$9466 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$664 \$8818 \$8787 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$665 \$8799 \$8798 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$666 \$8788 \$9472 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$667 \$8819 \$8788 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$668 \$8801 \$8800 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$669 \$8789 \$9478 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$670 \$8820 \$8789 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$671 \$8803 \$8802 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$672 \$8790 \$9484 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$673 \$8821 \$8790 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$674 \$8805 \$8804 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$675 \$8791 \$9490 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$676 \$8822 \$8791 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$677 \$8807 \$8806 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$678 \$8792 \$9496 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$679 \$8823 \$8792 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$680 \$8809 \$8808 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$681 \$8793 \$9502 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$682 \$8824 \$8793 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$683 \$8811 \$8810 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$684 \$8794 \$9508 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$685 \$8825 \$8794 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$686 \$8813 \$8812 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$687 \$8795 \$9514 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$688 \$8826 \$8795 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$689 \$8815 \$8814 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$690 \$8796 \$9520 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$691 \$8827 \$8796 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$692 \$8817 \$8816 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$693 \$9461 \$9527 D VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$694 \$9462 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$695 VSSD \$9461 \$9462 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$696 \$9463 \$9462 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$697 VSSD clks \$9463 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$698 \$9461 \$9528 \$9463 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$699 \$9465 \$9528 \$9462 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$700 \$9466 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$701 VSSD \$9465 \$9466 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$702 \$9464 \$9466 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$703 VSSD Set \$9464 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$704 \$9465 \$9527 \$9464 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$705 \$9467 \$9530 \$9466 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$706 \$9468 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$707 VSSD \$9467 \$9468 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$708 \$9469 \$9468 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$709 VSSD clks \$9469 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$710 \$9467 \$9531 \$9469 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$711 \$9471 \$9531 \$9468 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$712 \$9472 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$713 VSSD \$9471 \$9472 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$714 \$9470 \$9472 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$715 VSSD Set \$9470 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$716 \$9471 \$9530 \$9470 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$717 \$9473 \$9533 \$9472 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$718 \$9474 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$719 VSSD \$9473 \$9474 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$720 \$9475 \$9474 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$721 VSSD clks \$9475 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$722 \$9473 \$9534 \$9475 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$723 \$9477 \$9534 \$9474 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$724 \$9478 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$725 VSSD \$9477 \$9478 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$726 \$9476 \$9478 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$727 VSSD Set \$9476 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$728 \$9477 \$9533 \$9476 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$729 \$9479 \$9536 \$9478 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$730 \$9480 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$731 VSSD \$9479 \$9480 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$732 \$9481 \$9480 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$733 VSSD clks \$9481 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$734 \$9479 \$9537 \$9481 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$735 \$9483 \$9537 \$9480 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$736 \$9484 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$737 VSSD \$9483 \$9484 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$738 \$9482 \$9484 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$739 VSSD Set \$9482 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$740 \$9483 \$9536 \$9482 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$741 \$9485 \$9539 \$9484 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$742 \$9486 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$743 VSSD \$9485 \$9486 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$744 \$9487 \$9486 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$745 VSSD clks \$9487 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$746 \$9485 \$9540 \$9487 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$747 \$9489 \$9540 \$9486 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$748 \$9490 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$749 VSSD \$9489 \$9490 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$750 \$9488 \$9490 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$751 VSSD Set \$9488 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$752 \$9489 \$9539 \$9488 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$753 \$9491 \$9542 \$9490 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$754 \$9492 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$755 VSSD \$9491 \$9492 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$756 \$9493 \$9492 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$757 VSSD clks \$9493 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$758 \$9491 \$9543 \$9493 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$759 \$9495 \$9543 \$9492 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$760 \$9496 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$761 VSSD \$9495 \$9496 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$762 \$9494 \$9496 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$763 VSSD Set \$9494 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$764 \$9495 \$9542 \$9494 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$765 \$9497 \$9545 \$9496 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$766 \$9498 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$767 VSSD \$9497 \$9498 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$768 \$9499 \$9498 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$769 VSSD clks \$9499 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$770 \$9497 \$9546 \$9499 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$771 \$9501 \$9546 \$9498 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$772 \$9502 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$773 VSSD \$9501 \$9502 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$774 \$9500 \$9502 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$775 VSSD Set \$9500 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$776 \$9501 \$9545 \$9500 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$777 \$9503 \$9548 \$9502 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$778 \$9504 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$779 VSSD \$9503 \$9504 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$780 \$9505 \$9504 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$781 VSSD clks \$9505 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$782 \$9503 \$9549 \$9505 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$783 \$9507 \$9549 \$9504 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$784 \$9508 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$785 VSSD \$9507 \$9508 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$786 \$9506 \$9508 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$787 VSSD Set \$9506 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$788 \$9507 \$9548 \$9506 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$789 \$9509 \$9551 \$9508 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$790 \$9510 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$791 VSSD \$9509 \$9510 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$792 \$9511 \$9510 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$793 VSSD clks \$9511 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$794 \$9509 \$9552 \$9511 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$795 \$9513 \$9552 \$9510 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$796 \$9514 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$797 VSSD \$9513 \$9514 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$798 \$9512 \$9514 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$799 VSSD Set \$9512 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$800 \$9513 \$9551 \$9512 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$801 \$9515 \$9554 \$9514 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$802 \$9516 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$803 VSSD \$9515 \$9516 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$804 \$9517 \$9516 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$805 VSSD clks \$9517 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$806 \$9515 \$9555 \$9517 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$807 \$9519 \$9555 \$9516 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$808 \$9520 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$809 VSSD \$9519 \$9520 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$810 \$9518 \$9520 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$811 VSSD Set \$9518 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$812 \$9519 \$9554 \$9518 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$813 \$9521 \$9557 \$9520 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$814 \$9522 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$815 VSSD \$9521 \$9522 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$816 \$9523 \$9522 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$817 VSSD clks \$9523 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$818 \$9521 \$9558 \$9523 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$819 \$9526 \$9558 \$9522 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$820 CK_1 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$821 VSSD \$9526 CK_1 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$822 \$9525 CK_1 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$823 VSSD Set \$9525 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$824 \$9526 \$9557 \$9525 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$825 \$9527 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$826 \$9528 \$9527 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$827 \$9529 \$9466 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$828 \$9530 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$829 \$9531 \$9530 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$830 \$9382 \$10972 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$831 \$10972 \$11015 \$10973 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$832 VSSD \$11176 \$10972 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$833 \$11016 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$834 \$11017 \$11016 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$835 \$11792 \$11810 \$11747 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$836 \$9532 \$9472 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$837 \$11792 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$838 \$10974 \$11016 \$10973 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$839 \$9533 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$840 VSSD \$10973 \$11792 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$841 \$10975 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$842 \$9534 \$9533 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$843 VSSD \$10974 \$10975 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$844 \$10973 \$11747 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$845 VSSD Reset \$10973 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$846 \$10976 \$10975 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$847 VSSD Reset \$10976 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$848 \$11793 \$11811 \$11747 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$849 \$10974 \$11017 \$10976 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$850 \$11794 \$11811 \$11782 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$851 \$10979 \$11017 \$10975 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$852 \$11794 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$853 VSSD \$11793 \$11794 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$854 \$10977 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$855 VSSD \$10979 \$10977 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$856 \$11793 \$11782 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$857 VSSD Set \$11793 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$858 \$10978 \$10977 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$859 vocp \$11810 \$11782 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$860 VSSD Set \$10978 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$861 \$10979 \$11016 \$10978 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$862 \$11018 \$10977 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$863 \$9535 \$9478 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$864 \$9536 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$865 \$9537 \$9536 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$866 \$5831 \$10970 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$867 \$10970 \$11019 \$10980 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$868 VSSD \$11190 \$10970 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$869 \$9538 \$9484 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$870 \$11020 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$871 \$9539 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$872 \$11021 \$11020 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$873 \$11795 \$11814 \$11748 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$874 \$9540 \$9539 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$875 \$11795 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$876 \$10981 \$11020 \$10980 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$877 VSSD \$10980 \$11795 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$878 \$10982 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$879 VSSD \$10981 \$10982 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$880 \$10980 \$11748 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$881 VSSD Reset \$10980 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$882 \$10983 \$10982 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$883 VSSD Reset \$10983 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$884 \$11796 \$11815 \$11748 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$885 \$10981 \$11021 \$10983 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$886 \$11797 \$11815 \$11783 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$887 \$10986 \$11021 \$10982 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$888 \$11797 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$889 VSSD \$11796 \$11797 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$890 \$10984 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$891 VSSD \$10986 \$10984 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$892 \$11796 \$11783 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$893 VSSD Set \$11796 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$894 \$10985 \$10984 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$895 vocp \$11814 \$11783 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$896 VSSD Set \$10985 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$897 \$10986 \$11020 \$10985 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$898 \$11022 \$10984 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$899 \$9541 \$9490 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$900 \$9542 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$901 \$9543 \$9542 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$902 \$2939 \$10987 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$903 \$9544 \$9496 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$904 \$10987 \$11023 \$10988 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$905 VSSD \$11203 \$10987 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$906 \$9545 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$907 \$9546 \$9545 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$908 \$11024 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$909 \$11025 \$11024 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$910 \$11798 \$11818 \$11749 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$911 \$11798 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$912 \$10989 \$11024 \$10988 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$913 VSSD \$10988 \$11798 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$914 \$10990 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$915 VSSD \$10989 \$10990 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$916 \$10988 \$11749 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$917 VSSD Reset \$10988 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$918 \$10991 \$10990 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$919 VSSD Reset \$10991 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$920 \$11799 \$11819 \$11749 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$921 \$10989 \$11025 \$10991 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$922 \$11800 \$11819 \$11784 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$923 \$10994 \$11025 \$10990 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$924 \$11800 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$925 VSSD \$11799 \$11800 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$926 \$10992 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$927 VSSD \$10994 \$10992 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$928 \$11799 \$11784 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$929 VSSD Set \$11799 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$930 \$10993 \$10992 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$931 vocp \$11818 \$11784 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$932 VSSD Set \$10993 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$933 \$9547 \$9502 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$934 \$10994 \$11024 \$10993 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$935 \$9548 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$936 \$11026 \$10992 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$937 \$9549 \$9548 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$938 \$9550 \$9508 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$939 \$1275 \$10971 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$940 \$9551 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$941 \$9552 \$9551 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$942 \$10971 \$11027 \$10995 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$943 VSSD \$11216 \$10971 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$944 \$11028 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$945 \$11029 \$11028 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$946 \$11801 \$11822 \$11750 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$947 \$11801 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$948 \$10996 \$11028 \$10995 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$949 VSSD \$10995 \$11801 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$950 \$10997 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$951 VSSD \$10996 \$10997 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$952 \$10995 \$11750 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$953 VSSD Reset \$10995 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$954 \$10998 \$10997 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$955 VSSD Reset \$10998 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$956 \$11802 \$11823 \$11750 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$957 \$10996 \$11029 \$10998 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$958 \$11803 \$11823 \$11785 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$959 \$11001 \$11029 \$10997 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$960 \$11803 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$961 VSSD \$11802 \$11803 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$962 \$10999 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$963 VSSD \$11001 \$10999 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$964 \$11802 \$11785 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$965 \$9553 \$9514 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$966 VSSD Set \$11802 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$967 \$11000 \$10999 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$968 vocp \$11822 \$11785 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$969 VSSD Set \$11000 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$970 \$9554 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$971 \$9555 \$9554 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$972 \$11001 \$11028 \$11000 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$973 \$11030 \$10999 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$974 \$9556 \$9520 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$975 \$9557 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$976 \$9558 \$9557 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$977 \$1274 \$11002 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$978 \$11002 \$11031 \$11003 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$979 VSSD \$11229 \$11002 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$980 \$11032 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$981 \$11033 \$11032 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$982 \$11804 \$11826 \$11751 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$983 \$11804 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$984 \$11004 \$11032 \$11003 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$985 VSSD \$11003 \$11804 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$986 \$11005 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$987 VSSD \$11004 \$11005 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$988 \$11003 \$11751 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$989 VSSD Reset \$11003 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$990 \$11006 \$11005 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$991 VSSD Reset \$11006 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$992 \$11805 \$11827 \$11751 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$993 \$11004 \$11033 \$11006 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$994 \$11806 \$11827 \$11786 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$995 \$11009 \$11033 \$11005 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$996 \$9559 CK_1 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$997 \$11806 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$998 VSSD \$11805 \$11806 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$999 \$11007 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1000 VSSD \$11009 \$11007 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1001 \$11805 \$11786 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1002 VSSD Set \$11805 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1003 \$11008 \$11007 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1004 vocp \$11826 \$11786 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1005 VSSD Set \$11008 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1006 \$11009 \$11032 \$11008 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1007 \$11034 \$11007 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1008 \$12743 \$12775 \$12698 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1009 \$12743 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1010 VSSD \$12776 \$12743 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1011 \$12776 \$12698 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1012 VSSD Reset \$12776 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1013 \$12744 \$12968 \$12698 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1014 \$12745 \$12968 \$12732 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1015 \$12745 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1016 VSSD \$12744 \$12745 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1017 \$12744 \$12732 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1018 VSSD Set \$12744 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1019 \$12746 \$12775 \$12732 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1020 \$12733 \$12777 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1021 \$12746 \$12977 \$12733 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1022 VSSD \$12733 \$1263 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1023 \$9382 \$11176 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1024 \$11808 \$11015 \$10973 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1025 \$12747 \$12779 \$12699 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1026 VSSD \$10973 \$11809 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1027 \$12747 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1028 VSSD \$12780 \$12747 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1029 \$12780 \$12699 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1030 VSSD Reset \$12780 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1031 \$12748 \$12982 \$12699 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1032 \$12749 \$12982 \$12734 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1033 \$12749 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1034 VSSD \$12748 \$12749 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1035 \$12748 \$12734 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1036 VSSD Set \$12748 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1037 \$12750 \$12779 \$12734 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1038 VSSD \$11810 \$11811 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1039 \$12735 \$12781 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1040 VSSD \$11015 \$11810 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1041 \$12750 \$12991 \$12735 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1042 VSSD \$11176 \$11015 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1043 VSSD \$12735 \$1265 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1044 VSSD CK_1 \$11176 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1045 \$5831 \$11190 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1046 \$11812 \$11019 \$10980 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1047 \$12751 \$12783 \$12700 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1048 VSSD \$10980 \$11813 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1049 \$12751 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1050 VSSD \$12784 \$12751 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1051 \$12784 \$12700 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1052 VSSD Reset \$12784 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1053 \$12752 \$13004 \$12700 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1054 \$12753 \$13004 \$12736 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1055 \$12753 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1056 VSSD \$12752 \$12753 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1057 \$12752 \$12736 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1058 VSSD Set \$12752 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1059 \$12754 \$12783 \$12736 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1060 VSSD \$11814 \$11815 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1061 \$12755 \$12785 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1062 VSSD \$11019 \$11814 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1063 \$12754 \$13005 \$12755 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1064 VSSD \$11190 \$11019 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1065 VSSD \$12755 \$1267 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1066 VSSD \$9520 \$11190 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1067 \$2939 \$11203 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1068 \$11816 \$11023 \$10988 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1069 \$12756 \$12787 \$12701 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1070 VSSD \$10988 \$11817 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1071 \$12756 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1072 VSSD \$12788 \$12756 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1073 \$12788 \$12701 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1074 VSSD Reset \$12788 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1075 \$12757 \$13010 \$12701 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1076 \$12758 \$13010 \$12737 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1077 \$12758 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1078 VSSD \$12757 \$12758 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1079 \$12757 \$12737 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1080 VSSD Set \$12757 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1081 \$12759 \$12787 \$12737 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1082 VSSD \$11818 \$11819 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1083 \$12738 \$12789 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1084 VSSD \$11023 \$11818 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1085 \$12759 \$13019 \$12738 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1086 VSSD \$11203 \$11023 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1087 VSSD \$12738 \$2938 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1088 VSSD \$9514 \$11203 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1089 \$1275 \$11216 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1090 \$11820 \$11027 \$10995 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1091 \$12760 \$12791 \$12702 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1092 VSSD \$10995 \$11821 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1093 \$12760 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1094 VSSD \$12792 \$12760 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1095 \$12792 \$12702 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1096 VSSD Reset \$12792 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1097 \$12761 \$13024 \$12702 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1098 \$12762 \$13024 \$12739 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1099 \$12762 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1100 VSSD \$12761 \$12762 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1101 \$12761 \$12739 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1102 VSSD Set \$12761 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1103 \$12763 \$12791 \$12739 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1104 VSSD \$11822 \$11823 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1105 \$12740 \$12793 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1106 VSSD \$11027 \$11822 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1107 \$12763 \$13033 \$12740 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1108 VSSD \$11216 \$11027 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1109 VSSD \$12740 \$5830 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1110 VSSD \$9508 \$11216 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1111 \$1274 \$11229 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1112 \$11824 \$11031 \$11003 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1113 \$12764 \$12795 \$12703 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1114 VSSD \$11003 \$11825 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1115 \$12764 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1116 VSSD \$12796 \$12764 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1117 \$12796 \$12703 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1118 VSSD Reset \$12796 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1119 \$12765 \$13046 \$12703 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1120 \$12766 \$13046 \$12741 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1121 \$12766 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1122 VSSD \$12765 \$12766 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1123 \$12765 \$12741 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1124 VSSD Set \$12765 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1125 \$12767 \$12795 \$12741 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1126 VSSD \$11826 \$11827 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1127 \$12742 \$12797 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1128 VSSD \$11031 \$11826 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1129 \$12767 \$13047 \$12742 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1130 VSSD \$11229 \$11031 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1131 VSSD \$12742 \$1271 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1132 VSSD \$9502 \$11229 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1133 VSSD \$12776 \$12774 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1134 \$13705 \$13735 vocp VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1135 \$13706 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1136 VSSD \$13705 \$13706 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1137 \$13707 \$13706 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1138 VSSD Reset \$13707 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1139 \$13705 \$13879 \$13707 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1140 \$13709 \$13879 \$13706 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1141 \$12746 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1142 VSSD \$13709 \$12746 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1143 \$13708 \$12746 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1144 VSSD Set \$13708 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1145 \$13709 \$13735 \$13708 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1146 VSSD \$12775 \$12968 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1147 VSSD clks \$12775 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1148 VSSD \$12780 \$12778 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1149 \$13710 \$13738 vocp VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1150 \$13711 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1151 VSSD \$13710 \$13711 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1152 \$13712 \$13711 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1153 VSSD Reset \$13712 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1154 \$13710 \$13880 \$13712 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1155 \$13714 \$13880 \$13711 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1156 \$12750 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1157 VSSD \$13714 \$12750 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1158 \$13713 \$12750 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1159 VSSD Set \$13713 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1160 \$13714 \$13738 \$13713 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1161 VSSD \$12779 \$12982 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1162 VSSD clks \$12779 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1163 VSSD \$12784 \$12782 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1164 \$13715 \$13741 vocp VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1165 \$13716 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1166 VSSD \$13715 \$13716 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1167 \$13717 \$13716 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1168 VSSD Reset \$13717 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1169 \$13715 \$13881 \$13717 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1170 \$13719 \$13881 \$13716 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1171 \$12754 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1172 VSSD \$13719 \$12754 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1173 \$13718 \$12754 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1174 VSSD Set \$13718 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1175 \$13719 \$13741 \$13718 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1176 VSSD \$12783 \$13004 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1177 VSSD clks \$12783 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1178 VSSD \$12788 \$12786 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1179 \$13720 \$13744 vocp VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1180 \$13721 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1181 VSSD \$13720 \$13721 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1182 \$13722 \$13721 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1183 VSSD Reset \$13722 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1184 \$13720 \$13882 \$13722 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1185 \$13724 \$13882 \$13721 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1186 \$12759 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1187 VSSD \$13724 \$12759 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1188 \$13723 \$12759 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1189 VSSD Set \$13723 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1190 \$13724 \$13744 \$13723 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1191 VSSD \$12787 \$13010 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1192 VSSD clks \$12787 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1193 VSSD \$12792 \$12790 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1194 \$13725 \$13747 vocp VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1195 \$13726 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1196 VSSD \$13725 \$13726 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1197 \$13727 \$13726 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1198 VSSD Reset \$13727 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1199 \$13725 \$13883 \$13727 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1200 \$13729 \$13883 \$13726 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1201 \$12763 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1202 VSSD \$13729 \$12763 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1203 \$13728 \$12763 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1204 VSSD Set \$13728 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1205 \$13729 \$13747 \$13728 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1206 VSSD \$12791 \$13024 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1207 VSSD clks \$12791 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1208 VSSD \$12796 \$12794 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1209 \$13730 \$13750 vocp VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1210 \$13731 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1211 VSSD \$13730 \$13731 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1212 \$13732 \$13731 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1213 VSSD Reset \$13732 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1214 \$13730 \$13884 \$13732 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1215 \$13734 \$13884 \$13731 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1216 \$12767 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1217 VSSD \$13734 \$12767 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1218 \$13733 \$12767 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1219 VSSD Set \$13733 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1220 \$13734 \$13750 \$13733 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1221 VSSD \$12795 \$13046 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1222 VSSD clks \$12795 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1223 \$12777 \$9466 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1224 \$12977 \$12777 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1225 \$13735 \$12977 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1226 \$13879 \$13735 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1227 \$13736 \$12746 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1228 \$12746 \$12977 \$13737 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1229 VCM \$12777 \$1263 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1230 \$12781 \$9472 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1231 \$12991 \$12781 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1232 \$13738 \$12991 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1233 \$13880 \$13738 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1234 \$13739 \$12750 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1235 \$12750 \$12991 \$13740 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1236 VCM \$12781 \$1265 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1237 \$12785 \$9478 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1238 \$13005 \$12785 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1239 \$13741 \$13005 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1240 \$13881 \$13741 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1241 \$13742 \$12754 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1242 \$12754 \$13005 \$13743 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1243 VCM \$12785 \$1267 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1244 \$12789 \$9484 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1245 \$13019 \$12789 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1246 \$13744 \$13019 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1247 \$13882 \$13744 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1248 \$13745 \$12759 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1249 \$12759 \$13019 \$13746 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1250 VCM \$12789 \$2938 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1251 \$12793 \$9490 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1252 \$13033 \$12793 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1253 \$13747 \$13033 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1254 \$13883 \$13747 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1255 \$13748 \$12763 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1256 \$12763 \$13033 \$13749 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1257 VCM \$12793 \$5830 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1258 \$12797 \$9496 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1259 \$13047 \$12797 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1260 \$13750 \$13047 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1261 \$13884 \$13750 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1262 \$13751 \$12767 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1263 \$12767 \$13047 \$13752 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1264 VCM \$12797 \$1271 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
C$1265 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1266 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1267 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1268 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1269 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1270 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1271 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1272 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1273 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1274 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1275 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1276 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1277 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1278 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1279 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1280 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1281 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1282 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1283 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1284 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1285 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1286 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1287 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1288 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1289 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1290 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1291 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1292 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1293 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1294 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1295 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1296 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1297 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1298 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1299 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1300 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1301 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1302 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1303 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1304 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1305 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1306 \$1265 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1307 \$1267 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1308 \$1265 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1309 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1310 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1311 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1312 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1313 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1314 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1315 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1316 \$1274 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1317 \$1275 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1318 \$1274 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1319 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1320 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1321 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1322 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1323 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1324 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1325 \$1280 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1326 \$1282 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1327 \$1280 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1328 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1329 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1330 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1331 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1332 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1333 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1334 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1335 \$1289 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1336 \$1290 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1337 \$1289 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1338 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1339 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1340 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1341 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1342 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1343 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1344 \$1265 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1345 \$1267 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1346 \$1265 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1347 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1348 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1349 \$2938 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1350 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1351 \$2939 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1352 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1353 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1354 \$1274 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1355 \$1275 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1356 \$1274 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1357 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1358 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1359 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1360 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1361 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1362 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1363 \$1280 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1364 \$1282 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1365 \$1280 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1366 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1367 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1368 \$2940 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1369 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1370 \$2941 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1371 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1372 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1373 \$1289 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1374 \$1290 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1375 \$1289 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1376 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1377 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1378 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1379 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1380 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1381 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1382 \$1265 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1383 \$1267 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1384 \$1265 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1385 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1386 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1387 \$2938 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1388 \$1272 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1389 \$2939 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1390 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1391 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1392 \$1274 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1393 \$1275 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1394 \$1274 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1395 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1396 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1397 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1398 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1399 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1400 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1401 \$1280 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1402 \$1282 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1403 \$1280 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1404 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1405 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1406 \$2940 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1407 \$1287 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1408 \$2941 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1409 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1410 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1411 \$1289 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1412 \$1290 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1413 \$1289 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1414 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1415 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1416 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1417 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1418 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1419 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1420 \$1265 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1421 \$1267 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1422 \$1265 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1423 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1424 \$1263 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1425 \$5830 VDP 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1426 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1427 \$5831 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1428 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1429 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1430 \$1274 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1431 \$1275 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1432 \$1274 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1433 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1434 \$1271 \$1272 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1435 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1436 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1437 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1438 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1439 \$1280 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1440 \$1282 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1441 \$1280 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1442 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1443 \$1278 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1444 \$5832 VDN 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1445 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1446 \$5833 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1447 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1448 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1449 \$1289 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1450 \$1290 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1451 \$1289 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1452 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1453 \$1286 \$1287 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1454 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1455 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1456 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1457 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1458 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1459 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1460 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1461 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1462 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1463 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1464 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1465 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1466 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1467 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1468 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1469 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1470 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1471 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1472 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1473 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1474 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1475 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1476 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1477 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1478 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1479 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1480 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1481 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1482 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1483 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1484 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1485 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1486 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1487 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1488 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1489 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1490 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1491 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1492 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
.ENDS SAR_logic_dac
