** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/Folded/FC_bias_pfets.sch
.subckt FC_bias_pfets IREF VDD VB1 VB2 VB3
*.PININFO IREF:B VDD:B VB1:B VB2:B VB3:B
M13[1] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[2] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[3] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[4] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[5] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[6] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[7] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[8] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[9] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[10] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[11] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[12] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[13] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[14] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[15] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[16] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[17] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[18] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[19] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[20] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[21] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M13[22] IREF VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[1] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[2] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[3] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[4] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[5] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[6] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[7] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[8] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[9] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[10] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[11] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[12] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[13] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[14] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[15] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[16] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[17] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[18] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[19] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[20] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[21] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M14[22] VB3 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[1] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[2] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[3] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[4] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[5] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[6] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[7] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[8] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[9] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[10] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[11] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[12] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[13] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[14] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[15] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[16] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[17] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[18] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[19] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[20] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[21] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M15[22] VB2 VB1 VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[1] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[2] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[3] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[4] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[5] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[6] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[7] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[8] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[9] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[10] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[11] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[12] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[13] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[14] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[15] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[16] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[17] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[18] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[19] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[20] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[21] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[22] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[23] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[24] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[25] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[26] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[27] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[28] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[29] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[30] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[31] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[32] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[33] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[34] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[35] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[36] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[37] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
M1[38] VDD VDD VDD VDD pfet_03v3 L=2u W=2u nf=1 m=1
.ends
.end
