* Extracted by KLayout with GF180MCU LVS runset on : 30/04/2024 12:06

.SUBCKT SAR_top clks Vinp Vinn C B A D VDDA VSSD Vcom Valid VDDD Set Reset VCM
M$1 \$69 clks VDDA VDDA pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$2 \$70 \$69 VDDA VDDA pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$3 VDDA \$1087 \$4104 \$4104 pfet_03v3 L=0.28U W=4U AS=2.6P AD=2.6P PS=9.3U
+ PD=9.3U
M$4 \$1087 \$67 \$4104 \$4104 pfet_03v3 L=0.28U W=4U AS=2.6P AD=2.6P PS=9.3U
+ PD=9.3U
M$5 \$4106 \$75 \$73 \$4106 pfet_03v3 L=0.28U W=4U AS=2.6P AD=2.6P PS=9.3U
+ PD=9.3U
M$6 \$4106 \$73 VDDA \$4106 pfet_03v3 L=0.28U W=4U AS=2.6P AD=2.6P PS=9.3U
+ PD=9.3U
M$7 \$8656 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$8 \$8657 \$10778 \$8656 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$9 \$7400 Valid \$8657 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$10 \$8126 \$7400 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$11 \$67 \$70 VDDA VDDA pfet_03v3 L=0.28U W=4U AS=2.6P AD=2.6P PS=9.3U PD=9.3U
M$12 VDDA \$70 \$75 VDDA pfet_03v3 L=0.28U W=4U AS=2.6P AD=2.6P PS=9.3U PD=9.3U
M$13 \$7891 \$8126 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$14 \$8395 \$7891 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$15 \$8398 \$8396 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$16 \$8399 \$8371 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$17 \$9906 \$9904 \$8396 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$18 \$8396 \$9904 \$9906 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$19 \$9906 \$9904 \$8396 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$20 \$8396 \$9904 \$9906 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$21 \$9909 \$8385 \$8371 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$22 \$8371 \$8385 \$9909 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$23 \$9909 \$8385 \$8371 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$24 \$8371 \$8385 \$9909 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$25 \$10042 \$10720 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$26 \$10072 \$10042 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$27 \$10053 \$10052 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$28 \$10043 \$10726 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$29 \$10073 \$10043 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$30 \$10055 \$10054 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$31 \$10044 \$10732 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$32 \$10074 \$10044 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$33 \$10057 \$10056 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$34 \$10045 \$10738 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$35 \$10075 \$10045 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$36 \$10059 \$10058 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$37 \$10046 \$10744 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$38 \$10076 \$10046 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$39 \$10061 \$10060 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$40 \$9904 \$7891 VDDD VDDD pfet_03v3 L=0.28U W=2.35U AS=1.5275P AD=1.5275P
+ PS=6U PD=6U
M$41 VDDD \$7891 \$9904 VDDD pfet_03v3 L=0.28U W=2.35U AS=1.5275P AD=1.5275P
+ PS=6U PD=6U
M$42 \$8385 \$7891 VDDD VDDD pfet_03v3 L=0.28U W=2.35U AS=1.5275P AD=1.5275P
+ PS=6U PD=6U
M$43 VDDD \$7891 \$8385 VDDD pfet_03v3 L=0.28U W=2.35U AS=1.5275P AD=1.5275P
+ PS=6U PD=6U
M$44 \$10047 \$10750 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$45 \$10077 \$10047 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$46 VDDD \$8371 \$9906 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$47 \$9906 \$8371 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$48 VDDD \$8371 \$9906 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$49 \$9906 \$8371 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$50 VDDD \$8396 \$9909 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$51 \$9909 \$8396 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$52 \$10063 \$10062 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$53 VDDD \$8396 \$9909 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$54 \$9909 \$8396 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$55 Valid \$8399 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$56 VDDD \$8398 Valid VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$57 \$10048 \$10756 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$58 \$10078 \$10048 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$59 \$10065 \$10064 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$60 \$10049 \$10762 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$61 \$10079 \$10049 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$62 \$10067 \$10066 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$63 \$10050 \$10768 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$64 \$10080 \$10050 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$65 \$10069 \$10068 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$66 \$10051 \$10774 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$67 \$10081 \$10051 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$68 \$10071 \$10070 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$69 \$1630 \$10072 \$1624 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$70 \$10052 \$10042 \$1624 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$71 \$1630 \$10042 \$10053 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$72 \$1631 \$10073 \$1625 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$73 \$10054 \$10043 \$1625 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$74 \$1631 \$10043 \$10055 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$75 \$1632 \$10074 \$1626 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$76 \$10056 \$10044 \$1626 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$77 \$1632 \$10044 \$10057 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$78 \$3104 \$10075 \$3102 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$79 \$10058 \$10045 \$3102 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$80 \$3104 \$10045 \$10059 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$81 \$6827 \$10076 \$6823 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$82 \$10060 \$10046 \$6823 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$83 \$6827 \$10046 \$10061 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$84 \$1633 \$10077 \$1627 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$85 \$10062 \$10047 \$1627 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$86 \$1633 \$10047 \$10063 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$87 \$1634 \$10078 \$1628 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$88 \$10064 \$10048 \$1628 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$89 \$1634 \$10048 \$10065 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$90 \$1635 \$10079 \$1629 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$91 \$10066 \$10049 \$1629 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$92 \$1635 \$10049 \$10067 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$93 \$3105 \$10080 \$3103 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$94 \$10068 \$10050 \$3103 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$95 \$3105 \$10050 \$10069 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$96 \$6828 \$10081 \$6824 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$97 \$10070 \$10051 \$6824 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$98 \$6828 \$10051 \$10071 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$99 \$10781 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$100 \$10782 \$10781 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$101 \$10715 \$10782 D VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$102 \$11599 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$103 \$10716 \$10715 \$11599 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$104 \$11600 \$10716 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$105 \$10717 clks \$11600 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$106 \$10715 \$10781 \$10717 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$107 \$10719 \$10781 \$10716 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$108 \$11601 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$109 \$10720 \$10719 \$11601 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$110 \$11602 \$10720 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$111 \$10718 Set \$11602 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$112 \$10719 \$10782 \$10718 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$113 \$10783 \$10720 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$114 \$10784 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$115 \$10785 \$10784 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$116 \$10721 \$10785 \$10720 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$117 \$11603 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$118 \$10722 \$10721 \$11603 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$119 \$11604 \$10722 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$120 \$10723 clks \$11604 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$121 \$10721 \$10784 \$10723 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$122 \$10725 \$10784 \$10722 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$123 \$11605 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$124 \$10726 \$10725 \$11605 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$125 \$11606 \$10726 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$126 \$10724 Set \$11606 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$127 \$10725 \$10785 \$10724 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$128 \$10786 \$10726 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$129 \$10787 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$130 \$10788 \$10787 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$131 \$10727 \$10788 \$10726 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$132 \$11607 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$133 \$10728 \$10727 \$11607 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$134 \$11608 \$10728 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$135 \$10729 clks \$11608 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$136 \$10727 \$10787 \$10729 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$137 \$10731 \$10787 \$10728 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$138 \$11609 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$139 \$10732 \$10731 \$11609 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$140 \$11610 \$10732 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$141 \$10730 Set \$11610 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$142 \$10731 \$10788 \$10730 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$143 \$10789 \$10732 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$144 \$10790 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$145 \$10791 \$10790 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$146 \$10733 \$10791 \$10732 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$147 \$11611 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$148 \$10734 \$10733 \$11611 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$149 \$11612 \$10734 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$150 \$10735 clks \$11612 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$151 \$10733 \$10790 \$10735 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$152 \$10737 \$10790 \$10734 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$153 \$11613 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$154 \$10738 \$10737 \$11613 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$155 \$11614 \$10738 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$156 \$10736 Set \$11614 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$157 \$10737 \$10791 \$10736 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$158 \$10792 \$10738 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$159 \$10793 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$160 \$10794 \$10793 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$161 \$10739 \$10794 \$10738 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$162 \$11615 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$163 \$10740 \$10739 \$11615 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$164 \$11616 \$10740 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$165 \$10741 clks \$11616 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$166 \$10739 \$10793 \$10741 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$167 \$10743 \$10793 \$10740 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$168 \$11617 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$169 \$10744 \$10743 \$11617 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$170 \$11618 \$10744 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$171 \$10742 Set \$11618 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$172 \$10743 \$10794 \$10742 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$173 \$10795 \$10744 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$174 \$10796 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$175 \$10797 \$10796 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$176 \$10745 \$10797 \$10744 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$177 \$11619 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$178 \$10746 \$10745 \$11619 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$179 \$11620 \$10746 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$180 \$10747 clks \$11620 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$181 \$10745 \$10796 \$10747 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$182 \$10749 \$10796 \$10746 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$183 \$11621 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$184 \$10750 \$10749 \$11621 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$185 \$11622 \$10750 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$186 \$10748 Set \$11622 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$187 \$10749 \$10797 \$10748 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$188 \$10798 \$10750 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$189 \$10799 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$190 \$10800 \$10799 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$191 \$10751 \$10800 \$10750 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$192 \$11623 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$193 \$10752 \$10751 \$11623 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$194 \$11624 \$10752 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$195 \$10753 clks \$11624 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$196 \$10751 \$10799 \$10753 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$197 \$10755 \$10799 \$10752 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$198 \$11625 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$199 \$10756 \$10755 \$11625 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$200 \$11626 \$10756 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$201 \$10754 Set \$11626 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$202 \$10755 \$10800 \$10754 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$203 \$10801 \$10756 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$204 \$10802 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$205 \$10803 \$10802 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$206 \$10757 \$10803 \$10756 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$207 \$11627 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$208 \$10758 \$10757 \$11627 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$209 \$11628 \$10758 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$210 \$10759 clks \$11628 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$211 \$10757 \$10802 \$10759 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$212 \$10761 \$10802 \$10758 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$213 \$11629 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$214 \$10762 \$10761 \$11629 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$215 \$11630 \$10762 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$216 \$10760 Set \$11630 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$217 \$10761 \$10803 \$10760 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$218 \$10804 \$10762 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$219 \$10805 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$220 \$10806 \$10805 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$221 \$10763 \$10806 \$10762 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$222 \$11631 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$223 \$10764 \$10763 \$11631 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$224 \$11632 \$10764 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$225 \$10765 clks \$11632 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$226 \$10763 \$10805 \$10765 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$227 \$10767 \$10805 \$10764 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$228 \$11633 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$229 \$10768 \$10767 \$11633 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$230 \$11634 \$10768 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$231 \$10766 Set \$11634 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$232 \$10767 \$10806 \$10766 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$233 \$10807 \$10768 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$234 \$10808 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$235 \$10809 \$10808 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$236 \$10769 \$10809 \$10768 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$237 \$11635 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$238 \$10770 \$10769 \$11635 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$239 \$11636 \$10770 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$240 \$10771 clks \$11636 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$241 \$10769 \$10808 \$10771 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$242 \$10773 \$10808 \$10770 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$243 \$11637 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$244 \$10774 \$10773 \$11637 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$245 \$11638 \$10774 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$246 \$10772 Set \$11638 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$247 \$10773 \$10809 \$10772 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$248 \$10810 \$10774 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$249 \$10811 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$250 \$10812 \$10811 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$251 \$10775 \$10812 \$10774 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$252 \$11639 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$253 \$10776 \$10775 \$11639 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$254 \$11640 \$10776 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$255 \$10777 clks \$11640 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$256 \$10775 \$10811 \$10777 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$257 \$10780 \$10811 \$10776 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$258 \$11641 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$259 \$10778 \$10780 \$11641 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$260 \$11642 \$10778 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$261 \$10779 Set \$11642 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$262 \$10780 \$10812 \$10779 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$263 \$10813 \$10778 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$264 \$12222 \$12428 \$12227 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$265 VDDD \$12227 \$13062 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$266 \$12268 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$267 \$12269 \$12268 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$268 \$13045 \$13064 \$13000 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$269 \$13576 Set \$13045 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$270 \$12228 \$12269 \$12227 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$271 VDDD \$12227 \$13576 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$272 \$12645 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$273 \$12229 \$12228 \$12645 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$274 \$13577 \$13000 \$12227 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$275 VDDD Reset \$13577 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$276 \$12646 \$12229 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$277 \$12230 Reset \$12646 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$278 \$13046 \$13063 \$13000 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$279 \$12228 \$12268 \$12230 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$280 \$13047 \$13063 \$13035 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$281 \$12233 \$12268 \$12229 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$282 \$13578 Reset \$13047 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$283 VDDD \$13046 \$13578 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$284 \$12647 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$285 \$12231 \$12233 \$12647 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$286 \$13579 \$13035 \$13046 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$287 VDDD Set \$13579 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$288 \$12648 \$12231 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$289 \$8399 \$13064 \$13035 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$290 \$12232 Set \$12648 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$291 \$12233 \$12269 \$12232 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$292 VDDD \$13063 \$13064 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$293 VDDD \$12267 \$13063 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$294 \$12270 \$12231 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$295 VDDD \$12428 \$12267 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$296 VDDD \$10778 \$12428 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$297 \$12223 \$12442 \$12234 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$298 VDDD \$12234 \$13066 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$299 \$12272 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$300 \$12273 \$12272 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$301 \$13048 \$13068 \$13001 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$302 \$13580 Set \$13048 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$303 \$12235 \$12273 \$12234 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$304 VDDD \$12234 \$13580 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$305 \$12649 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$306 \$12236 \$12235 \$12649 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$307 \$13581 \$13001 \$12234 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$308 VDDD Reset \$13581 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$309 \$12650 \$12236 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$310 \$12237 Reset \$12650 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$311 \$13049 \$13067 \$13001 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$312 \$12235 \$12272 \$12237 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$313 \$13050 \$13067 \$13036 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$314 \$12240 \$12272 \$12236 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$315 \$13582 Reset \$13050 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$316 VDDD \$13049 \$13582 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$317 \$12651 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$318 \$12238 \$12240 \$12651 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$319 \$13583 \$13036 \$13049 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$320 VDDD Set \$13583 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$321 \$12652 \$12238 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$322 \$8399 \$13068 \$13036 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$323 \$12239 Set \$12652 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$324 \$12240 \$12273 \$12239 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$325 VDDD \$13067 \$13068 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$326 VDDD \$12271 \$13067 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$327 \$12274 \$12238 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$328 VDDD \$12442 \$12271 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$329 VDDD \$10774 \$12442 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$330 \$12224 \$12455 \$12241 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$331 VDDD \$12241 \$13070 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$332 \$12276 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$333 \$12277 \$12276 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$334 \$13051 \$13072 \$13002 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$335 \$13584 Set \$13051 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$336 \$12242 \$12277 \$12241 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$337 VDDD \$12241 \$13584 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$338 \$12653 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$339 \$12243 \$12242 \$12653 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$340 \$13585 \$13002 \$12241 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$341 VDDD Reset \$13585 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$342 \$12654 \$12243 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$343 \$12244 Reset \$12654 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$344 \$13052 \$13071 \$13002 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$345 \$12242 \$12276 \$12244 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$346 \$13053 \$13071 \$13037 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$347 \$12247 \$12276 \$12243 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$348 \$13586 Reset \$13053 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$349 VDDD \$13052 \$13586 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$350 \$12655 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$351 \$12245 \$12247 \$12655 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$352 \$13587 \$13037 \$13052 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$353 VDDD Set \$13587 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$354 \$12656 \$12245 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$355 \$8399 \$13072 \$13037 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$356 \$12246 Set \$12656 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$357 \$12247 \$12277 \$12246 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$358 VDDD \$13071 \$13072 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$359 VDDD \$12275 \$13071 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$360 \$12278 \$12245 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$361 VDDD \$12455 \$12275 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$362 VDDD \$10768 \$12455 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$363 \$12225 \$12468 \$12248 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$364 VDDD \$12248 \$13074 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$365 \$12280 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$366 \$12281 \$12280 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$367 \$13054 \$13076 \$13003 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$368 \$13588 Set \$13054 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$369 \$12249 \$12281 \$12248 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$370 VDDD \$12248 \$13588 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$371 \$12657 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$372 \$12250 \$12249 \$12657 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$373 \$13589 \$13003 \$12248 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$374 VDDD Reset \$13589 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$375 \$12658 \$12250 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$376 \$12251 Reset \$12658 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$377 \$13055 \$13075 \$13003 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$378 \$12249 \$12280 \$12251 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$379 \$13056 \$13075 \$13038 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$380 \$12254 \$12280 \$12250 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$381 \$13590 Reset \$13056 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$382 VDDD \$13055 \$13590 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$383 \$12659 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$384 \$12252 \$12254 \$12659 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$385 \$13591 \$13038 \$13055 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$386 VDDD Set \$13591 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$387 \$12660 \$12252 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$388 \$8399 \$13076 \$13038 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$389 \$12253 Set \$12660 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$390 \$12254 \$12281 \$12253 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$391 VDDD \$13075 \$13076 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$392 VDDD \$12279 \$13075 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$393 \$12282 \$12252 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$394 VDDD \$12468 \$12279 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$395 VDDD \$10762 \$12468 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$396 \$12226 \$12481 \$12255 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$397 VDDD \$12255 \$13078 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$398 \$12284 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$399 \$12285 \$12284 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$400 \$13057 \$13080 \$13004 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$401 \$13592 Set \$13057 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$402 \$12256 \$12285 \$12255 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$403 VDDD \$12255 \$13592 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$404 \$12661 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$405 \$12257 \$12256 \$12661 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$406 \$13593 \$13004 \$12255 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$407 VDDD Reset \$13593 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$408 \$12662 \$12257 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$409 \$12258 Reset \$12662 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$410 \$13058 \$13079 \$13004 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$411 \$12256 \$12284 \$12258 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$412 \$13059 \$13079 \$13039 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$413 \$12261 \$12284 \$12257 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$414 \$13594 Reset \$13059 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$415 VDDD \$13058 \$13594 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$416 \$12663 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$417 \$12259 \$12261 \$12663 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$418 \$13595 \$13039 \$13058 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$419 VDDD Set \$13595 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$420 \$12664 \$12259 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$421 \$8399 \$13080 \$13039 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$422 \$12260 Set \$12664 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$423 \$12261 \$12285 \$12260 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$424 VDDD \$13079 \$13080 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$425 VDDD \$12283 \$13079 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$426 \$12286 \$12259 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$427 VDDD \$12481 \$12283 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$428 VDDD \$10756 \$12481 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$429 VDDD \$14029 \$14027 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$430 \$13997 \$14221 \$13951 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$431 \$14478 Set \$13997 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$432 VDDD \$14029 \$14478 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$433 \$14479 \$13951 \$14029 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$434 VDDD Reset \$14479 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$435 \$13998 \$14028 \$13951 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$436 \$13999 \$14028 \$13985 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$437 \$14480 Reset \$13999 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$438 VDDD \$13998 \$14480 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$439 \$14481 \$13985 \$13998 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$440 VDDD Set \$14481 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$441 \$14000 \$14221 \$13985 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$442 VDDD \$14028 \$14221 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$443 VDDD clks \$14028 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$444 \$14000 \$14030 \$13986 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$445 \$10635 \$12267 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$446 VDDD \$13061 \$10635 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$447 \$13061 \$12428 \$12227 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$448 VDDD \$14033 \$14031 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$449 VDDD \$12267 \$13061 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$450 \$14001 \$14235 \$13952 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$451 \$14482 Set \$14001 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$452 VDDD \$14033 \$14482 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$453 \$14483 \$13952 \$14033 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$454 VDDD Reset \$14483 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$455 \$14002 \$14032 \$13952 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$456 \$14003 \$14032 \$13987 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$457 \$14484 Reset \$14003 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$458 VDDD \$14002 \$14484 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$459 \$14485 \$13987 \$14002 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$460 VDDD Set \$14485 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$461 \$14004 \$14235 \$13987 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$462 VDDD \$14032 \$14235 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$463 VDDD clks \$14032 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$464 \$14004 \$14034 \$13988 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$465 \$6824 \$12271 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$466 VDDD \$13065 \$6824 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$467 \$13065 \$12442 \$12234 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$468 VDDD \$14037 \$14035 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$469 VDDD \$12271 \$13065 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$470 \$14005 \$14257 \$13953 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$471 \$14486 Set \$14005 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$472 VDDD \$14037 \$14486 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$473 \$14487 \$13953 \$14037 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$474 VDDD Reset \$14487 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$475 \$14006 \$14036 \$13953 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$476 \$14007 \$14036 \$13989 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$477 \$14488 Reset \$14007 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$478 VDDD \$14006 \$14488 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$479 \$14489 \$13989 \$14006 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$480 VDDD Set \$14489 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$481 \$14008 \$14257 \$13989 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$482 VDDD \$14036 \$14257 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$483 VDDD clks \$14036 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$484 \$14008 \$14038 \$13990 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$485 \$3103 \$12275 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$486 VDDD \$13069 \$3103 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$487 \$13069 \$12455 \$12241 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$488 VDDD \$14041 \$14039 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$489 VDDD \$12275 \$13069 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$490 \$14009 \$14263 \$13954 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$491 \$14490 Set \$14009 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$492 VDDD \$14041 \$14490 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$493 \$14491 \$13954 \$14041 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$494 VDDD Reset \$14491 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$495 \$14010 \$14040 \$13954 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$496 \$14011 \$14040 \$13991 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$497 \$14492 Reset \$14011 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$498 VDDD \$14010 \$14492 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$499 \$14493 \$13991 \$14010 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$500 VDDD Set \$14493 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$501 \$14012 \$14263 \$13991 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$502 VDDD \$14040 \$14263 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$503 VDDD clks \$14040 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$504 \$14012 \$14042 \$13992 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$505 \$1629 \$12279 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$506 VDDD \$13073 \$1629 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$507 \$13073 \$12468 \$12248 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$508 VDDD \$14045 \$14043 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$509 VDDD \$12279 \$13073 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$510 \$14013 \$14277 \$13955 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$511 \$14494 Set \$14013 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$512 VDDD \$14045 \$14494 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$513 \$14495 \$13955 \$14045 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$514 VDDD Reset \$14495 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$515 \$14014 \$14044 \$13955 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$516 \$14015 \$14044 \$13993 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$517 \$14496 Reset \$14015 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$518 VDDD \$14014 \$14496 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$519 \$14497 \$13993 \$14014 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$520 VDDD Set \$14497 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$521 \$14016 \$14277 \$13993 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$522 VDDD \$14044 \$14277 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$523 VDDD clks \$14044 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$524 \$14016 \$14046 \$13994 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$525 \$1628 \$12283 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$526 VDDD \$13077 \$1628 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$527 \$13077 \$12481 \$12255 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$528 VDDD \$14049 \$14047 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$529 VDDD \$12283 \$13077 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$530 \$14017 \$14291 \$13956 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$531 \$14498 Set \$14017 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$532 VDDD \$14049 \$14498 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$533 \$14499 \$13956 \$14049 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$534 VDDD Reset \$14499 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$535 \$14018 \$14048 \$13956 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$536 \$14019 \$14048 \$13995 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$537 \$14500 Reset \$14019 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$538 VDDD \$14018 \$14500 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$539 \$14501 \$13995 \$14018 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$540 VDDD Set \$14501 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$541 \$14020 \$14291 \$13995 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$542 VDDD \$14048 \$14291 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$543 VDDD clks \$14048 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$544 \$14020 \$14050 \$13996 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$545 \$14030 \$10720 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$546 \$14230 \$14030 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$547 \$14988 \$14230 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$548 \$15132 \$14988 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$549 \$14958 \$15132 \$8399 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$550 \$15612 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$551 \$14959 \$14958 \$15612 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$552 \$15613 \$14959 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$553 \$14960 Reset \$15613 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$554 \$14958 \$14988 \$14960 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$555 \$14962 \$14988 \$14959 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$556 \$15614 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$557 \$14000 \$14962 \$15614 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$558 \$15615 \$14000 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$559 \$14961 Set \$15615 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$560 \$14962 \$15132 \$14961 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$561 \$14989 \$14000 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$562 \$14034 \$10726 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$563 \$14244 \$14034 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$564 \$14991 \$14244 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$565 \$15133 \$14991 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$566 \$14963 \$15133 \$8399 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$567 \$15616 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$568 \$14964 \$14963 \$15616 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$569 \$15617 \$14964 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$570 \$14965 Reset \$15617 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$571 \$14963 \$14991 \$14965 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$572 \$14967 \$14991 \$14964 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$573 \$15618 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$574 \$14004 \$14967 \$15618 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$575 \$15619 \$14004 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$576 \$14966 Set \$15619 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$577 \$14967 \$15133 \$14966 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$578 \$14992 \$14004 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$579 \$14038 \$10732 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$580 \$14258 \$14038 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$581 \$14994 \$14258 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$582 \$15134 \$14994 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$583 \$14968 \$15134 \$8399 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$584 \$15620 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$585 \$14969 \$14968 \$15620 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$586 \$15621 \$14969 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$587 \$14970 Reset \$15621 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$588 \$14968 \$14994 \$14970 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$589 \$14972 \$14994 \$14969 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$590 \$15622 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$591 \$14008 \$14972 \$15622 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$592 \$15623 \$14008 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$593 \$14971 Set \$15623 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$594 \$14972 \$15134 \$14971 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$595 \$14995 \$14008 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$596 \$14042 \$10738 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$597 \$14272 \$14042 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$598 \$14997 \$14272 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$599 \$15135 \$14997 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$600 \$14973 \$15135 \$8399 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$601 \$15624 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$602 \$14974 \$14973 \$15624 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$603 \$15625 \$14974 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$604 \$14975 Reset \$15625 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$605 \$14973 \$14997 \$14975 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$606 \$14977 \$14997 \$14974 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$607 \$15626 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$608 \$14012 \$14977 \$15626 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$609 \$15627 \$14012 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$610 \$14976 Set \$15627 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$611 \$14977 \$15135 \$14976 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$612 \$14998 \$14012 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$613 \$14046 \$10744 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$614 \$14286 \$14046 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$615 \$15000 \$14286 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$616 \$15136 \$15000 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$617 \$14978 \$15136 \$8399 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$618 \$15628 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$619 \$14979 \$14978 \$15628 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$620 \$15629 \$14979 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$621 \$14980 Reset \$15629 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$622 \$14978 \$15000 \$14980 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$623 \$14982 \$15000 \$14979 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$624 \$15630 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$625 \$14016 \$14982 \$15630 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$626 \$15631 \$14016 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$627 \$14981 Set \$15631 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$628 \$14982 \$15136 \$14981 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$629 \$15001 \$14016 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$630 \$14050 \$10750 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$631 \$14300 \$14050 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$632 \$15003 \$14300 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$633 \$15137 \$15003 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$634 \$14983 \$15137 \$8399 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$635 \$15632 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$636 \$14984 \$14983 \$15632 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$637 \$15633 \$14984 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$638 \$14985 Reset \$15633 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$639 \$14983 \$15003 \$14985 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$640 \$14987 \$15003 \$14984 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$641 \$15634 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$642 \$14020 \$14987 \$15634 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$643 \$15635 \$14020 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$644 \$14986 Set \$15635 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$645 \$14987 \$15137 \$14986 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$646 \$15004 \$14020 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$647 \$14990 \$14230 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$648 \$14000 \$14030 \$14990 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$649 \$1624 \$14990 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$650 VCM \$14230 \$1624 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$651 \$14993 \$14244 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$652 \$14004 \$14034 \$14993 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$653 \$1625 \$14993 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$654 VCM \$14244 \$1625 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$655 \$14996 \$14258 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$656 \$14008 \$14038 \$14996 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$657 \$1626 \$14996 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$658 VCM \$14258 \$1626 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$659 \$14999 \$14272 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$660 \$14012 \$14042 \$14999 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$661 \$3102 \$14999 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$662 VCM \$14272 \$3102 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$663 \$15002 \$14286 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$664 \$14016 \$14046 \$15002 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$665 \$6823 \$15002 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$666 VCM \$14286 \$6823 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$667 \$15005 \$14300 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$668 \$14020 \$14050 \$15005 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$669 \$1627 \$15005 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$670 VCM \$14300 \$1627 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$671 \$69 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$672 \$70 \$69 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$673 \$1647 VSSD Vcom VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$674 \$1647 \$1087 Vinp VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P
+ PS=13.22U PD=13.22U
M$675 \$1647 VSSD Vcom VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$676 \$1647 \$1087 Vinp VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P
+ PS=13.22U PD=13.22U
M$677 \$1647 VSSD Vcom VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$678 \$1647 \$1087 Vinp VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P
+ PS=13.22U PD=13.22U
M$679 \$1647 VSSD Vcom VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$680 \$1647 \$1087 Vinp VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P
+ PS=13.22U PD=13.22U
M$681 \$1647 VSSD Vcom VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$682 \$1647 \$1087 Vinp VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P
+ PS=13.22U PD=13.22U
M$683 \$67 \$70 \$66 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$684 \$67 \$1087 \$66 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$685 VSSD \$69 \$66 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$686 Vinp \$1087 \$66 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$687 \$68 VDDA \$1087 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$688 VSSD \$69 \$68 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$689 \$72 \$69 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$690 \$73 VDDA \$72 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$691 \$74 \$73 Vinn VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$692 \$74 \$69 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$693 \$74 \$73 \$75 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$694 \$74 \$70 \$75 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$695 Vinn \$73 \$1651 VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$696 Vcom VSSD \$1651 VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$697 Vinn \$73 \$1651 VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$698 Vcom VSSD \$1651 VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$699 Vinn \$73 \$1651 VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$700 Vcom VSSD \$1651 VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$701 Vinn \$73 \$1651 VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$702 Vcom VSSD \$1651 VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$703 Vinn \$73 \$1651 VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$704 Vcom VSSD \$1651 VSSD nfet_03v3 L=0.28U W=6U AS=3.66P AD=3.66P PS=13.22U
+ PD=13.22U
M$705 \$7400 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$706 VSSD \$10778 \$7400 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$707 VSSD Valid \$7400 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$708 \$7890 \$7400 VSSD VSSD nfet_03v3 L=35U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$709 \$7890 \$7400 \$8126 VSSD nfet_03v3 L=35U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$710 \$8382 \$7400 \$8911 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$711 \$8382 \$7400 VSSD VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$712 \$8126 A \$8911 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$713 \$8383 \$7400 VSSD VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$714 \$8126 B \$8912 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$715 \$8383 \$7400 \$8912 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$716 \$8384 \$7400 VSSD VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$717 \$8126 C \$8913 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$718 \$8384 \$7400 \$8913 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$719 \$7891 \$8126 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$720 \$8394 \$1647 \$8385 VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$721 \$8394 \$1651 \$9904 VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$722 \$9904 \$1651 \$8394 VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$723 \$8385 \$1647 \$8394 VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$724 \$8394 \$7891 VSSD VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$725 \$8394 \$1647 \$8385 VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$726 \$8394 \$1651 \$9904 VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$727 VSSD \$7891 \$8394 VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$728 \$9904 \$1651 \$8394 VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$729 \$8385 \$1647 \$8394 VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$730 \$8394 \$7891 VSSD VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$731 \$8394 \$1647 \$8385 VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$732 \$8394 \$1651 \$9904 VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$733 \$8385 \$1647 \$8394 VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$734 \$9904 \$1651 \$8394 VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$735 \$8395 \$7891 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$736 \$8396 \$8395 VSSD VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$737 VSSD \$8396 \$8371 VSSD nfet_03v3 L=0.28U W=6.3U AS=3.843P AD=2.52P
+ PS=13.82U PD=7.1U
M$738 \$8396 \$8371 VSSD VSSD nfet_03v3 L=0.28U W=6.3U AS=2.52P AD=3.843P
+ PS=7.1U PD=13.82U
M$739 \$8371 \$8395 VSSD VSSD nfet_03v3 L=0.28U W=3.1U AS=1.891P AD=1.891P
+ PS=7.42U PD=7.42U
M$740 \$8398 \$8396 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$741 \$8399 \$8371 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$742 \$8372 \$8399 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$743 Valid \$8398 \$8372 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$744 \$1630 \$10042 \$1624 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$745 \$10052 \$10072 \$1624 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$746 \$1630 \$10072 \$10053 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$747 \$1631 \$10043 \$1625 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$748 \$10054 \$10073 \$1625 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$749 \$1631 \$10073 \$10055 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$750 \$1632 \$10044 \$1626 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$751 \$10056 \$10074 \$1626 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$752 \$1632 \$10074 \$10057 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$753 \$3104 \$10045 \$3102 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$754 \$10058 \$10075 \$3102 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$755 \$3104 \$10075 \$10059 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$756 \$6827 \$10046 \$6823 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$757 \$10060 \$10076 \$6823 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$758 \$6827 \$10076 \$10061 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$759 \$1633 \$10047 \$1627 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$760 \$10062 \$10077 \$1627 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$761 \$1633 \$10077 \$10063 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$762 \$1634 \$10048 \$1628 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$763 \$10064 \$10078 \$1628 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$764 \$1634 \$10078 \$10065 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$765 \$1635 \$10049 \$1629 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$766 \$10066 \$10079 \$1629 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$767 \$1635 \$10079 \$10067 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$768 \$3105 \$10050 \$3103 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$769 \$10068 \$10080 \$3103 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$770 \$3105 \$10080 \$10069 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$771 \$6828 \$10051 \$6824 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$772 \$10070 \$10081 \$6824 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$773 \$6828 \$10081 \$10071 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$774 \$10042 \$10720 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$775 \$10072 \$10042 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$776 \$10053 \$10052 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$777 \$10043 \$10726 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$778 \$10073 \$10043 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$779 \$10055 \$10054 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$780 \$10044 \$10732 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$781 \$10074 \$10044 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$782 \$10057 \$10056 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$783 \$10045 \$10738 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$784 \$10075 \$10045 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$785 \$10059 \$10058 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$786 \$10046 \$10744 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$787 \$10076 \$10046 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$788 \$10061 \$10060 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$789 \$10047 \$10750 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$790 \$10077 \$10047 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$791 \$10063 \$10062 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$792 \$10048 \$10756 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$793 \$10078 \$10048 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$794 \$10065 \$10064 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$795 \$10049 \$10762 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$796 \$10079 \$10049 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$797 \$10067 \$10066 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$798 \$10050 \$10768 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$799 \$10080 \$10050 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$800 \$10069 \$10068 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$801 \$10051 \$10774 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$802 \$10081 \$10051 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$803 \$10071 \$10070 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$804 \$10715 \$10781 D VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$805 \$10716 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$806 VSSD \$10715 \$10716 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$807 \$10717 \$10716 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$808 VSSD clks \$10717 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$809 \$10715 \$10782 \$10717 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$810 \$10719 \$10782 \$10716 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$811 \$10720 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$812 VSSD \$10719 \$10720 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$813 \$10718 \$10720 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$814 VSSD Set \$10718 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$815 \$10719 \$10781 \$10718 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$816 \$10721 \$10784 \$10720 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$817 \$10722 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$818 VSSD \$10721 \$10722 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$819 \$10723 \$10722 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$820 VSSD clks \$10723 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$821 \$10721 \$10785 \$10723 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$822 \$10725 \$10785 \$10722 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$823 \$10726 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$824 VSSD \$10725 \$10726 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$825 \$10724 \$10726 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$826 VSSD Set \$10724 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$827 \$10725 \$10784 \$10724 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$828 \$10727 \$10787 \$10726 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$829 \$10728 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$830 VSSD \$10727 \$10728 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$831 \$10729 \$10728 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$832 VSSD clks \$10729 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$833 \$10727 \$10788 \$10729 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$834 \$10731 \$10788 \$10728 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$835 \$10732 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$836 VSSD \$10731 \$10732 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$837 \$10730 \$10732 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$838 VSSD Set \$10730 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$839 \$10731 \$10787 \$10730 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$840 \$10733 \$10790 \$10732 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$841 \$10734 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$842 VSSD \$10733 \$10734 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$843 \$10735 \$10734 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$844 VSSD clks \$10735 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$845 \$10733 \$10791 \$10735 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$846 \$10737 \$10791 \$10734 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$847 \$10738 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$848 VSSD \$10737 \$10738 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$849 \$10736 \$10738 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$850 VSSD Set \$10736 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$851 \$10737 \$10790 \$10736 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$852 \$10739 \$10793 \$10738 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$853 \$10740 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$854 VSSD \$10739 \$10740 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$855 \$10741 \$10740 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$856 VSSD clks \$10741 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$857 \$10739 \$10794 \$10741 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$858 \$10743 \$10794 \$10740 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$859 \$10744 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$860 VSSD \$10743 \$10744 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$861 \$10742 \$10744 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$862 VSSD Set \$10742 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$863 \$10743 \$10793 \$10742 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$864 \$10745 \$10796 \$10744 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$865 \$10746 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$866 VSSD \$10745 \$10746 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$867 \$10747 \$10746 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$868 VSSD clks \$10747 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$869 \$10745 \$10797 \$10747 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$870 \$10749 \$10797 \$10746 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$871 \$10750 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$872 VSSD \$10749 \$10750 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$873 \$10748 \$10750 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$874 VSSD Set \$10748 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$875 \$10749 \$10796 \$10748 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$876 \$10751 \$10799 \$10750 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$877 \$10752 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$878 VSSD \$10751 \$10752 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$879 \$10753 \$10752 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$880 VSSD clks \$10753 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$881 \$10751 \$10800 \$10753 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$882 \$10755 \$10800 \$10752 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$883 \$10756 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$884 VSSD \$10755 \$10756 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$885 \$10754 \$10756 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$886 VSSD Set \$10754 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$887 \$10755 \$10799 \$10754 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$888 \$10757 \$10802 \$10756 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$889 \$10758 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$890 VSSD \$10757 \$10758 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$891 \$10759 \$10758 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$892 VSSD clks \$10759 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$893 \$10757 \$10803 \$10759 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$894 \$10761 \$10803 \$10758 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$895 \$10762 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$896 VSSD \$10761 \$10762 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$897 \$10760 \$10762 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$898 VSSD Set \$10760 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$899 \$10761 \$10802 \$10760 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$900 \$10763 \$10805 \$10762 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$901 \$10764 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$902 VSSD \$10763 \$10764 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$903 \$10765 \$10764 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$904 VSSD clks \$10765 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$905 \$10763 \$10806 \$10765 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$906 \$10767 \$10806 \$10764 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$907 \$10768 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$908 VSSD \$10767 \$10768 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$909 \$10766 \$10768 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$910 VSSD Set \$10766 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$911 \$10767 \$10805 \$10766 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$912 \$10769 \$10808 \$10768 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$913 \$10770 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$914 VSSD \$10769 \$10770 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$915 \$10771 \$10770 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$916 VSSD clks \$10771 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$917 \$10769 \$10809 \$10771 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$918 \$10773 \$10809 \$10770 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$919 \$10774 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$920 VSSD \$10773 \$10774 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$921 \$10772 \$10774 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$922 VSSD Set \$10772 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$923 \$10773 \$10808 \$10772 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$924 \$10775 \$10811 \$10774 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$925 \$10776 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$926 VSSD \$10775 \$10776 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$927 \$10777 \$10776 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$928 VSSD clks \$10777 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$929 \$10775 \$10812 \$10777 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$930 \$10780 \$10812 \$10776 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$931 \$10778 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$932 VSSD \$10780 \$10778 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$933 \$10779 \$10778 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$934 VSSD Set \$10779 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$935 \$10780 \$10811 \$10779 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$936 \$10781 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$937 \$10782 \$10781 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$938 \$10783 \$10720 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$939 \$10784 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$940 \$10785 \$10784 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$941 \$10635 \$12222 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$942 \$12222 \$12267 \$12227 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$943 VSSD \$12428 \$12222 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$944 \$12268 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$945 \$12269 \$12268 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$946 \$13045 \$13063 \$13000 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$947 \$10786 \$10726 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$948 \$13045 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$949 \$12228 \$12268 \$12227 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$950 \$10787 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$951 VSSD \$12227 \$13045 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$952 \$12229 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$953 \$10788 \$10787 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$954 VSSD \$12228 \$12229 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$955 \$12227 \$13000 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$956 VSSD Reset \$12227 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$957 \$12230 \$12229 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$958 VSSD Reset \$12230 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$959 \$13046 \$13064 \$13000 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$960 \$12228 \$12269 \$12230 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$961 \$13047 \$13064 \$13035 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$962 \$12233 \$12269 \$12229 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$963 \$13047 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$964 VSSD \$13046 \$13047 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$965 \$12231 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$966 VSSD \$12233 \$12231 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$967 \$13046 \$13035 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$968 VSSD Set \$13046 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$969 \$12232 \$12231 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$970 \$8399 \$13063 \$13035 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$971 VSSD Set \$12232 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$972 \$12233 \$12268 \$12232 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$973 \$12270 \$12231 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$974 \$10789 \$10732 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$975 \$10790 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$976 \$10791 \$10790 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$977 \$6824 \$12223 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$978 \$12223 \$12271 \$12234 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$979 VSSD \$12442 \$12223 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$980 \$10792 \$10738 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$981 \$12272 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$982 \$10793 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$983 \$12273 \$12272 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$984 \$13048 \$13067 \$13001 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$985 \$10794 \$10793 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$986 \$13048 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$987 \$12235 \$12272 \$12234 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$988 VSSD \$12234 \$13048 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$989 \$12236 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$990 VSSD \$12235 \$12236 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$991 \$12234 \$13001 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$992 VSSD Reset \$12234 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$993 \$12237 \$12236 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$994 VSSD Reset \$12237 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$995 \$13049 \$13068 \$13001 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$996 \$12235 \$12273 \$12237 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$997 \$13050 \$13068 \$13036 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$998 \$12240 \$12273 \$12236 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$999 \$13050 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1000 VSSD \$13049 \$13050 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1001 \$12238 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1002 VSSD \$12240 \$12238 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1003 \$13049 \$13036 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1004 VSSD Set \$13049 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1005 \$12239 \$12238 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1006 \$8399 \$13067 \$13036 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1007 VSSD Set \$12239 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1008 \$12240 \$12272 \$12239 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1009 \$12274 \$12238 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1010 \$10795 \$10744 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1011 \$10796 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1012 \$10797 \$10796 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1013 \$3103 \$12224 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1014 \$10798 \$10750 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1015 \$12224 \$12275 \$12241 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1016 VSSD \$12455 \$12224 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1017 \$10799 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1018 \$10800 \$10799 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1019 \$12276 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1020 \$12277 \$12276 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1021 \$13051 \$13071 \$13002 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1022 \$13051 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1023 \$12242 \$12276 \$12241 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1024 VSSD \$12241 \$13051 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1025 \$12243 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1026 VSSD \$12242 \$12243 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1027 \$12241 \$13002 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1028 VSSD Reset \$12241 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1029 \$12244 \$12243 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1030 VSSD Reset \$12244 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1031 \$13052 \$13072 \$13002 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1032 \$12242 \$12277 \$12244 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1033 \$13053 \$13072 \$13037 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1034 \$12247 \$12277 \$12243 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1035 \$13053 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1036 VSSD \$13052 \$13053 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1037 \$12245 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1038 VSSD \$12247 \$12245 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1039 \$13052 \$13037 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1040 VSSD Set \$13052 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1041 \$12246 \$12245 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1042 \$8399 \$13071 \$13037 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1043 VSSD Set \$12246 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1044 \$10801 \$10756 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1045 \$12247 \$12276 \$12246 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1046 \$10802 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1047 \$12278 \$12245 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1048 \$10803 \$10802 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1049 \$10804 \$10762 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1050 \$1629 \$12225 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1051 \$10805 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1052 \$12225 \$12279 \$12248 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1053 \$10806 \$10805 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1054 VSSD \$12468 \$12225 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1055 \$12280 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1056 \$12281 \$12280 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1057 \$13054 \$13075 \$13003 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1058 \$13054 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1059 \$12249 \$12280 \$12248 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1060 VSSD \$12248 \$13054 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1061 \$12250 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1062 VSSD \$12249 \$12250 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1063 \$12248 \$13003 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1064 VSSD Reset \$12248 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1065 \$12251 \$12250 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1066 VSSD Reset \$12251 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1067 \$13055 \$13076 \$13003 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1068 \$12249 \$12281 \$12251 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1069 \$13056 \$13076 \$13038 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1070 \$12254 \$12281 \$12250 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1071 \$13056 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1072 VSSD \$13055 \$13056 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1073 \$12252 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1074 VSSD \$12254 \$12252 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1075 \$13055 \$13038 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1076 \$10807 \$10768 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1077 VSSD Set \$13055 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1078 \$12253 \$12252 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1079 \$8399 \$13075 \$13038 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1080 VSSD Set \$12253 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1081 \$10808 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1082 \$10809 \$10808 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1083 \$12254 \$12280 \$12253 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1084 \$12282 \$12252 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1085 \$10810 \$10774 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1086 \$10811 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1087 \$10812 \$10811 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1088 \$1628 \$12226 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1089 \$12226 \$12283 \$12255 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1090 VSSD \$12481 \$12226 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1091 \$12284 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1092 \$12285 \$12284 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1093 \$13057 \$13079 \$13004 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1094 \$13057 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1095 \$12256 \$12284 \$12255 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1096 VSSD \$12255 \$13057 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1097 \$12257 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1098 VSSD \$12256 \$12257 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1099 \$12255 \$13004 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1100 VSSD Reset \$12255 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1101 \$12258 \$12257 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1102 VSSD Reset \$12258 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1103 \$13058 \$13080 \$13004 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1104 \$12256 \$12285 \$12258 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1105 \$13059 \$13080 \$13039 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1106 \$12261 \$12285 \$12257 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1107 \$10813 \$10778 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1108 \$13059 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1109 VSSD \$13058 \$13059 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1110 \$12259 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1111 VSSD \$12261 \$12259 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1112 \$13058 \$13039 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1113 VSSD Set \$13058 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1114 \$12260 \$12259 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1115 \$8399 \$13079 \$13039 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1116 VSSD Set \$12260 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1117 \$12261 \$12284 \$12260 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1118 \$12286 \$12259 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1119 \$13997 \$14028 \$13951 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1120 \$13997 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1121 VSSD \$14029 \$13997 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1122 \$14029 \$13951 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1123 VSSD Reset \$14029 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1124 \$13998 \$14221 \$13951 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1125 \$13999 \$14221 \$13985 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1126 \$13999 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1127 VSSD \$13998 \$13999 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1128 \$13998 \$13985 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1129 VSSD Set \$13998 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1130 \$14000 \$14028 \$13985 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1131 \$13986 \$14030 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1132 \$14000 \$14230 \$13986 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1133 VSSD \$13986 \$1624 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1134 \$10635 \$12428 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1135 \$13061 \$12267 \$12227 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1136 \$14001 \$14032 \$13952 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1137 VSSD \$12227 \$13062 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1138 \$14001 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1139 VSSD \$14033 \$14001 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1140 \$14033 \$13952 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1141 VSSD Reset \$14033 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1142 \$14002 \$14235 \$13952 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1143 \$14003 \$14235 \$13987 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1144 \$14003 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1145 VSSD \$14002 \$14003 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1146 \$14002 \$13987 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1147 VSSD Set \$14002 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1148 \$14004 \$14032 \$13987 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1149 VSSD \$13063 \$13064 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1150 \$13988 \$14034 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1151 VSSD \$12267 \$13063 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1152 \$14004 \$14244 \$13988 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1153 VSSD \$12428 \$12267 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1154 VSSD \$13988 \$1625 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1155 VSSD \$10778 \$12428 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1156 \$6824 \$12442 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1157 \$13065 \$12271 \$12234 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1158 \$14005 \$14036 \$13953 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1159 VSSD \$12234 \$13066 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1160 \$14005 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1161 VSSD \$14037 \$14005 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1162 \$14037 \$13953 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1163 VSSD Reset \$14037 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1164 \$14006 \$14257 \$13953 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1165 \$14007 \$14257 \$13989 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1166 \$14007 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1167 VSSD \$14006 \$14007 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1168 \$14006 \$13989 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1169 VSSD Set \$14006 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1170 \$14008 \$14036 \$13989 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1171 VSSD \$13067 \$13068 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1172 \$13990 \$14038 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1173 VSSD \$12271 \$13067 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1174 \$14008 \$14258 \$13990 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1175 VSSD \$12442 \$12271 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1176 VSSD \$13990 \$1626 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1177 VSSD \$10774 \$12442 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1178 \$3103 \$12455 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1179 \$13069 \$12275 \$12241 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1180 \$14009 \$14040 \$13954 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1181 VSSD \$12241 \$13070 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1182 \$14009 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1183 VSSD \$14041 \$14009 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1184 \$14041 \$13954 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1185 VSSD Reset \$14041 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1186 \$14010 \$14263 \$13954 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1187 \$14011 \$14263 \$13991 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1188 \$14011 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1189 VSSD \$14010 \$14011 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1190 \$14010 \$13991 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1191 VSSD Set \$14010 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1192 \$14012 \$14040 \$13991 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1193 VSSD \$13071 \$13072 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1194 \$13992 \$14042 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1195 VSSD \$12275 \$13071 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1196 \$14012 \$14272 \$13992 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1197 VSSD \$12455 \$12275 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1198 VSSD \$13992 \$3102 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1199 VSSD \$10768 \$12455 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1200 \$1629 \$12468 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1201 \$13073 \$12279 \$12248 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1202 \$14013 \$14044 \$13955 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1203 VSSD \$12248 \$13074 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1204 \$14013 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1205 VSSD \$14045 \$14013 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1206 \$14045 \$13955 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1207 VSSD Reset \$14045 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1208 \$14014 \$14277 \$13955 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1209 \$14015 \$14277 \$13993 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1210 \$14015 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1211 VSSD \$14014 \$14015 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1212 \$14014 \$13993 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1213 VSSD Set \$14014 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1214 \$14016 \$14044 \$13993 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1215 VSSD \$13075 \$13076 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1216 \$13994 \$14046 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1217 VSSD \$12279 \$13075 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1218 \$14016 \$14286 \$13994 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1219 VSSD \$12468 \$12279 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1220 VSSD \$13994 \$6823 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1221 VSSD \$10762 \$12468 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1222 \$1628 \$12481 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1223 \$13077 \$12283 \$12255 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1224 \$14017 \$14048 \$13956 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1225 VSSD \$12255 \$13078 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1226 \$14017 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1227 VSSD \$14049 \$14017 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1228 \$14049 \$13956 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1229 VSSD Reset \$14049 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1230 \$14018 \$14291 \$13956 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1231 \$14019 \$14291 \$13995 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1232 \$14019 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1233 VSSD \$14018 \$14019 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1234 \$14018 \$13995 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1235 VSSD Set \$14018 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1236 \$14020 \$14048 \$13995 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1237 VSSD \$13079 \$13080 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1238 \$13996 \$14050 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1239 VSSD \$12283 \$13079 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1240 \$14020 \$14300 \$13996 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1241 VSSD \$12481 \$12283 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1242 VSSD \$13996 \$1627 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1243 VSSD \$10756 \$12481 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1244 VSSD \$14029 \$14027 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1245 \$14958 \$14988 \$8399 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1246 \$14959 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1247 VSSD \$14958 \$14959 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1248 \$14960 \$14959 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1249 VSSD Reset \$14960 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1250 \$14958 \$15132 \$14960 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1251 \$14962 \$15132 \$14959 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1252 \$14000 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1253 VSSD \$14962 \$14000 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1254 \$14961 \$14000 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1255 VSSD Set \$14961 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1256 \$14962 \$14988 \$14961 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1257 VSSD \$14028 \$14221 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1258 VSSD clks \$14028 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1259 VSSD \$14033 \$14031 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1260 \$14963 \$14991 \$8399 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1261 \$14964 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1262 VSSD \$14963 \$14964 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1263 \$14965 \$14964 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1264 VSSD Reset \$14965 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1265 \$14963 \$15133 \$14965 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1266 \$14967 \$15133 \$14964 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1267 \$14004 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1268 VSSD \$14967 \$14004 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1269 \$14966 \$14004 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1270 VSSD Set \$14966 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1271 \$14967 \$14991 \$14966 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1272 VSSD \$14032 \$14235 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1273 VSSD clks \$14032 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1274 VSSD \$14037 \$14035 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1275 \$14968 \$14994 \$8399 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1276 \$14969 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1277 VSSD \$14968 \$14969 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1278 \$14970 \$14969 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1279 VSSD Reset \$14970 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1280 \$14968 \$15134 \$14970 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1281 \$14972 \$15134 \$14969 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1282 \$14008 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1283 VSSD \$14972 \$14008 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1284 \$14971 \$14008 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1285 VSSD Set \$14971 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1286 \$14972 \$14994 \$14971 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1287 VSSD \$14036 \$14257 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1288 VSSD clks \$14036 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1289 VSSD \$14041 \$14039 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1290 \$14973 \$14997 \$8399 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1291 \$14974 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1292 VSSD \$14973 \$14974 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1293 \$14975 \$14974 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1294 VSSD Reset \$14975 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1295 \$14973 \$15135 \$14975 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1296 \$14977 \$15135 \$14974 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1297 \$14012 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1298 VSSD \$14977 \$14012 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1299 \$14976 \$14012 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1300 VSSD Set \$14976 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1301 \$14977 \$14997 \$14976 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1302 VSSD \$14040 \$14263 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1303 VSSD clks \$14040 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1304 VSSD \$14045 \$14043 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1305 \$14978 \$15000 \$8399 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1306 \$14979 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1307 VSSD \$14978 \$14979 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1308 \$14980 \$14979 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1309 VSSD Reset \$14980 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1310 \$14978 \$15136 \$14980 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1311 \$14982 \$15136 \$14979 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1312 \$14016 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1313 VSSD \$14982 \$14016 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1314 \$14981 \$14016 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1315 VSSD Set \$14981 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1316 \$14982 \$15000 \$14981 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1317 VSSD \$14044 \$14277 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1318 VSSD clks \$14044 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1319 VSSD \$14049 \$14047 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1320 \$14983 \$15003 \$8399 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1321 \$14984 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1322 VSSD \$14983 \$14984 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1323 \$14985 \$14984 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1324 VSSD Reset \$14985 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1325 \$14983 \$15137 \$14985 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1326 \$14987 \$15137 \$14984 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1327 \$14020 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1328 VSSD \$14987 \$14020 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1329 \$14986 \$14020 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1330 VSSD Set \$14986 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1331 \$14987 \$15003 \$14986 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1332 VSSD \$14048 \$14291 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1333 VSSD clks \$14048 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1334 \$14030 \$10720 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1335 \$14230 \$14030 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1336 \$14988 \$14230 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1337 \$15132 \$14988 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1338 \$14989 \$14000 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1339 \$14000 \$14230 \$14990 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1340 VCM \$14030 \$1624 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1341 \$14034 \$10726 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1342 \$14244 \$14034 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1343 \$14991 \$14244 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1344 \$15133 \$14991 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1345 \$14992 \$14004 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1346 \$14004 \$14244 \$14993 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1347 VCM \$14034 \$1625 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1348 \$14038 \$10732 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1349 \$14258 \$14038 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1350 \$14994 \$14258 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1351 \$15134 \$14994 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1352 \$14995 \$14008 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1353 \$14008 \$14258 \$14996 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1354 VCM \$14038 \$1626 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1355 \$14042 \$10738 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1356 \$14272 \$14042 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1357 \$14997 \$14272 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1358 \$15135 \$14997 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1359 \$14998 \$14012 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1360 \$14012 \$14272 \$14999 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1361 VCM \$14042 \$3102 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1362 \$14046 \$10744 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1363 \$14286 \$14046 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1364 \$15000 \$14286 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1365 \$15136 \$15000 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1366 \$15001 \$14016 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1367 \$14016 \$14286 \$15002 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1368 VCM \$14046 \$6823 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1369 \$14050 \$10750 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1370 \$14300 \$14050 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1371 \$15003 \$14300 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1372 \$15137 \$15003 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1373 \$15004 \$14020 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1374 \$14020 \$14300 \$15005 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1375 VCM \$14050 \$1627 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
C$1376 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1377 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1378 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1379 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1380 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1381 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1382 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1383 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1384 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1385 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1386 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1387 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1388 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1389 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1390 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1391 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1392 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1393 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1394 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1395 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1396 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1397 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1398 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1399 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1400 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1401 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1402 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1403 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1404 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1405 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1406 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1407 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1408 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1409 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1410 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1411 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1412 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1413 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1414 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1415 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1416 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1417 \$1625 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1418 \$1626 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1419 \$1625 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1420 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1421 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1422 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1423 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1424 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1425 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1426 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1427 \$1628 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1428 \$1629 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1429 \$1628 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1430 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1431 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1432 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1433 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1434 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1435 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1436 \$1631 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1437 \$1632 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1438 \$1631 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1439 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1440 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1441 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1442 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1443 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1444 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1445 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1446 \$1634 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1447 \$1635 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1448 \$1634 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1449 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1450 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1451 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1452 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1453 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1454 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1455 \$1625 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1456 \$1626 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1457 \$1625 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1458 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1459 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1460 \$3102 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1461 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1462 \$3103 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1463 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1464 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1465 \$1628 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1466 \$1629 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1467 \$1628 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1468 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1469 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1470 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1471 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1472 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1473 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1474 \$1631 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1475 \$1632 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1476 \$1631 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1477 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1478 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1479 \$3104 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1480 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1481 \$3105 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1482 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1483 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1484 \$1634 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1485 \$1635 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1486 \$1634 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1487 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1488 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1489 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1490 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1491 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1492 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1493 \$1625 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1494 \$1626 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1495 \$1625 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1496 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1497 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1498 \$3102 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1499 \$1649 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1500 \$3103 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1501 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1502 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1503 \$1628 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1504 \$1629 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1505 \$1628 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1506 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1507 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1508 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1509 \$66 \$4104 2e-13 cap_mim_2f0_m4m5_noshield A=100P P=40U
C$1510 \$66 \$4104 2e-13 cap_mim_2f0_m4m5_noshield A=100P P=40U
C$1511 \$66 \$4104 2e-13 cap_mim_2f0_m4m5_noshield A=100P P=40U
C$1512 \$74 \$4106 2e-13 cap_mim_2f0_m4m5_noshield A=100P P=40U
C$1513 \$74 \$4106 2e-13 cap_mim_2f0_m4m5_noshield A=100P P=40U
C$1514 \$74 \$4106 2e-13 cap_mim_2f0_m4m5_noshield A=100P P=40U
C$1515 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1516 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1517 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1518 \$1631 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1519 \$1632 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1520 \$1631 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1521 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1522 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1523 \$3104 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1524 \$1653 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1525 \$3105 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1526 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1527 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1528 \$1634 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1529 \$1635 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1530 \$1634 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1531 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1532 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1533 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1534 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1535 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1536 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1537 \$1625 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1538 \$1626 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1539 \$1625 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1540 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1541 \$1624 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1542 \$6823 \$1647 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1543 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1544 \$6824 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1545 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1546 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1547 \$1628 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1548 \$1629 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1549 \$1628 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1550 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1551 \$1627 \$1649 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1552 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1553 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1554 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1555 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1556 \$1631 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1557 \$1632 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1558 \$1631 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1559 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1560 \$1630 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1561 \$6827 \$1651 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1562 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1563 \$6828 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1564 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1565 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1566 \$1634 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1567 \$1635 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1568 \$1634 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1569 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1570 \$1633 \$1653 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1571 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1572 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1573 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1574 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1575 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1576 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1577 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1578 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1579 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1580 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1581 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1582 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1583 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1584 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1585 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1586 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1587 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1588 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1589 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1590 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1591 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1592 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1593 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1594 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1595 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1596 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1597 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1598 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1599 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1600 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1601 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1602 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1603 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1604 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1605 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1606 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1607 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1608 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
C$1609 VSSD VSSD 5e-14 cap_mim_2f0_m4m5_noshield A=25P P=20U
.ENDS SAR_top
