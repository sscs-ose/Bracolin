* Extracted by KLayout with GF180MCU LVS runset on : 15/04/2024 20:03

.SUBCKT clock_generator_delay_cell IN OUT VDDD VSSD A B C
M$1 OUT IN VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$2 \$2 IN VSSD VSSD nfet_03v3 L=35U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$3 \$2 IN OUT VSSD nfet_03v3 L=35U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$4 \$10 IN VSSD VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$5 \$11 IN VSSD VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$6 \$12 IN VSSD VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$7 \$10 IN \$17 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$8 \$11 IN \$18 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$9 \$12 IN \$19 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$10 OUT A \$17 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$11 OUT B \$18 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
M$12 OUT C \$19 VSSD nfet_03v3 L=2U W=1.56U AS=0.9516P AD=0.9516P PS=4.34U
+ PD=4.34U
.ENDS clock_generator_delay_cell
