** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/Folded/FC_net.sch
.subckt FC_net AVDD AVSS VOUT VP VN VB1 VB2 VB3 VB4
*.PININFO AVDD:B AVSS:B VOUT:B VP:B VN:B VB1:B VB2:B VB3:B VB4:B
x1 net1 net1 net2 net3 VP VN AVDD FC_pfets_x4
x2 AVDD AVDD net1 net1 VB1 VB1 AVDD FC_pfets_x4
x3 AVDD AVDD net4 net5 M3_D M3_D AVDD FC_pfets_x4
x4 net4 net5 M3_D VOUT VB4 VB4 AVDD FC_pfets_x4
x5 net2 net3 M3_D VOUT VB3 VB3 AVSS FC_nfets
x6 AVSS AVSS net2 net3 VB2 VB2 AVSS FC_nfets_x2
.ends

* expanding   symbol:  /home/gmaranhao/Desktop/Bracolin/TIA_Filter/Folded/FC_pfets_x4.sym # of
*+ pins=7
** sym_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/Folded/FC_pfets_x4.sym
** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/Folded/FC_pfets_x4.sch
.subckt FC_pfets_x4 S1 S2 D1 D2 G1 G2 B
*.PININFO S1:B S2:B D1:B D2:B G1:B G2:B B:B
x1[1] S1 S2 D1 D2 G1 G2 B FC_pfets
x1[2] S1 S2 D1 D2 G1 G2 B FC_pfets
x1[3] S1 S2 D1 D2 G1 G2 B FC_pfets
x1[4] S1 S2 D1 D2 G1 G2 B FC_pfets
.ends


* expanding   symbol:  /home/gmaranhao/Desktop/Bracolin/TIA_Filter/Folded/FC_nfets.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/Folded/FC_nfets.sym
** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/Folded/FC_nfets.sch
.subckt FC_nfets S1 S2 D1 D2 G1 G2 B
*.PININFO S1:B S2:B D1:B D2:B G1:B G2:B B:B
M1[1] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[2] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[3] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[4] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[5] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[6] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[7] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[8] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[9] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[10] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[11] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[12] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[13] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[14] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[15] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[16] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[17] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M1[18] D1 G1 S1 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[1] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[2] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[3] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[4] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[5] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[6] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[7] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[8] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[9] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[10] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[11] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[12] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[13] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[14] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[15] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[16] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[17] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M2[18] D2 G2 S2 B nfet_03v3 L=2u W=2u nf=1 m=1
M3[1] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[2] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[3] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[4] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[5] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[6] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[7] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[8] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[9] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[10] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[11] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[12] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[13] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[14] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[15] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[16] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[17] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[18] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[19] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[20] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[21] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[22] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[23] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[24] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[25] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[26] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[27] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[28] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[29] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
M3[30] B B B B nfet_03v3 L=2u W=2u nf=1 m=1
.ends


* expanding   symbol:  /home/gmaranhao/Desktop/Bracolin/TIA_Filter/Folded/FC_nfets_x2.sym # of
*+ pins=7
** sym_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/Folded/FC_nfets_x2.sym
** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/Folded/FC_nfets_x2.sch
.subckt FC_nfets_x2 S1 S2 D1 D2 G1 G2 B
*.PININFO S1:B S2:B D1:B D2:B G1:B G2:B B:B
x1[1] S1 S2 D1 D2 G1 G2 B FC_nfets
x1[2] S1 S2 D1 D2 G1 G2 B FC_nfets
.ends


* expanding   symbol:  /home/gmaranhao/Desktop/Bracolin/TIA_Filter/Folded/FC_pfets.sym # of pins=7
** sym_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/Folded/FC_pfets.sym
** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/Folded/FC_pfets.sch
.subckt FC_pfets S1 S2 D1 D2 G1 G2 B
*.PININFO S1:B S2:B D1:B D2:B G1:B G2:B B:B
M1[1] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[2] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[3] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[4] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[5] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[6] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[7] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[8] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[9] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[10] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[11] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[12] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[13] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[14] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[15] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[16] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[17] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[18] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[19] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[20] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[21] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M1[22] D1 G1 S1 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[1] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[2] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[3] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[4] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[5] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[6] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[7] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[8] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[9] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[10] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[11] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[12] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[13] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[14] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[15] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[16] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[17] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[18] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[19] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[20] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[21] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M2[22] D2 G2 S2 B pfet_03v3 L=2u W=2u nf=1 m=1
M3[1] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[2] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[3] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[4] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[5] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[6] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[7] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[8] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[9] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[10] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[11] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[12] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[13] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[14] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[15] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[16] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[17] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[18] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[19] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[20] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[21] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[22] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[23] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[24] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[25] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[26] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[27] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[28] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[29] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[30] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[31] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[32] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[33] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
M3[34] B B B B pfet_03v3 L=2u W=2u nf=1 m=1
.ends

.end
