* NGSPICE file created from CM_input.ext - technology: gf180mcuD

.subckt CM_input ISBCS INP INP2 INN INN2 VDD VSS
X0 a_3930_2285# ISBCS.t4 VSS.t57 VSS.t48 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X1 a_948_n291# ISBCS.t2 ISBCS.t3 VSS.t47 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X2 INN.t0 a_n389_6663.t0 a_3947_7622# VDD.t9 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3 a_3930_609# ISBCS.t5 VSS.t56 VSS.t48 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X4 INN2.t0 a_n389_6663.t0 a_3947_5704# VDD.t9 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X5 VSS.t45 VSS.t44 VSS.t45 VSS.t10 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X6 VSS.t43 VSS.t42 VSS.t43 VSS.t7 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X7 VSS.t41 VSS.t40 VSS.t41 VSS.t24 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X8 a_n389_6663.t0 ISBCS.t6 a_3930_609# VSS.t46 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X9 VDD.t47 VDD.t46 VDD.t47 VDD.t9 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X10 VSS.t55 ISBCS.t7 a_948_1385# VSS.t50 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X11 a_n389_6663.t1 a_n389_6663.t0 a_3947_6663# VDD.t9 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X12 a_3930_n291# ISBCS.t8 VSS.t54 VSS.t48 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X13 VDD.t45 VDD.t44 VDD.t45 VDD.t9 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X14 VSS.t53 ISBCS.t9 a_948_609# VSS.t50 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X15 VSS.t39 VSS.t38 VSS.t39 VSS.t10 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X16 VSS.t37 VSS.t36 VSS.t37 VSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X17 VSS.t35 VSS.t34 VSS.t35 VSS.t7 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X18 a_3947_7622# a_n389_6663.t0 VDD.t8 VDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X19 VDD.t43 VDD.t42 VDD.t43 VDD.t30 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X20 VSS.t33 VSS.t32 VSS.t33 VSS.t10 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X21 VSS.t31 VSS.t30 VSS.t31 VSS.t7 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X22 a_3947_5704# a_n389_6663.t0 VDD.t7 VDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X23 VSS.t29 VSS.t28 VSS.t29 VSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X24 VSS.t52 ISBCS.t10 a_948_2285# VSS.t50 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X25 VDD.t41 VDD.t40 VDD.t41 VDD.t30 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X26 a_948_609# ISBCS.t11 INP2.t1 VSS.t47 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X27 VSS.t27 VSS.t26 VSS.t27 VSS.t1 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X28 a_941_7622# a_n389_6663.t0 INN2.t1 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X29 VDD.t39 VDD.t38 VDD.t39 VDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X30 a_n389_6663.t0 ISBCS.t12 a_3930_1385# VSS.t46 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X31 a_3947_6663# a_n389_6663.t0 VDD.t6 VDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X32 VDD.t37 VDD.t36 VDD.t37 VDD.t30 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X33 VDD.t35 VDD.t34 VDD.t35 VDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X34 VDD.t33 VDD.t32 VDD.t33 VDD.t30 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X35 a_941_5704# a_n389_6663.t0 INN.t1 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X36 VDD.t31 VDD.t29 VDD.t31 VDD.t30 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X37 a_948_1385# ISBCS.t13 INP2.t0 VSS.t47 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X38 VDD.t4 a_n389_6663.t0 a_941_7622# VDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X39 VDD.t28 VDD.t27 VDD.t28 VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X40 VSS.t25 VSS.t23 VSS.t25 VSS.t24 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X41 VSS.t51 ISBCS.t14 a_948_n291# VSS.t50 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X42 VDD.t26 VDD.t25 VDD.t26 VDD.t13 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X43 a_941_6663# a_n389_6663.t0 a_n389_6663.t0 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X44 VSS.t22 VSS.t21 VSS.t22 VSS.t7 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X45 VDD.t24 VDD.t23 VDD.t24 VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X46 VDD.t22 VDD.t21 VDD.t22 VDD.t13 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X47 VDD.t2 a_n389_6663.t0 a_941_5704# VDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X48 VSS.t20 VSS.t19 VSS.t20 VSS.t10 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X49 VDD.t20 VDD.t19 VDD.t20 VDD.t13 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X50 VDD.t18 VDD.t17 VDD.t18 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X51 VDD.t16 VDD.t15 VDD.t16 VDD.t13 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X52 VDD.t1 a_n389_6663.t0 a_941_6663# VDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X53 ISBCS.t1 ISBCS.t0 a_3930_2285# VSS.t46 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X54 a_3930_1385# ISBCS.t15 VSS.t49 VSS.t48 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X55 VSS.t18 VSS.t17 VSS.t18 VSS.t7 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X56 VSS.t16 VSS.t15 VSS.t16 VSS.t10 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X57 VDD.t14 VDD.t12 VDD.t14 VDD.t13 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X58 VDD.t11 VDD.t10 VDD.t11 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X59 VSS.t14 VSS.t12 VSS.t14 VSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X60 a_948_2285# ISBCS.t16 INP.t1 VSS.t47 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X61 VSS.t11 VSS.t9 VSS.t11 VSS.t10 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X62 VSS.t8 VSS.t6 VSS.t8 VSS.t7 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X63 INP.t0 ISBCS.t17 a_3930_n291# VSS.t46 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X64 VSS.t5 VSS.t3 VSS.t5 VSS.t4 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X65 VSS.t2 VSS.t0 VSS.t2 VSS.t1 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
R0 ISBCS.n8 ISBCS.t1 10.2879
R1 ISBCS ISBCS.n31 6.52263
R2 ISBCS.t0 ISBCS.n9 4.39661
R3 ISBCS.n7 ISBCS.t12 4.39661
R4 ISBCS.t6 ISBCS.n1 4.39661
R5 ISBCS.t17 ISBCS.n25 4.39661
R6 ISBCS.n10 ISBCS.t0 4.39661
R7 ISBCS.n26 ISBCS.t17 4.39661
R8 ISBCS.n13 ISBCS.t16 4.39651
R9 ISBCS.n12 ISBCS.t16 4.39651
R10 ISBCS.n21 ISBCS.t11 4.39651
R11 ISBCS.n19 ISBCS.t13 4.39651
R12 ISBCS.n29 ISBCS.t2 4.39651
R13 ISBCS.n28 ISBCS.t2 4.39651
R14 ISBCS ISBCS.t3 3.79155
R15 ISBCS.n13 ISBCS.t10 2.96638
R16 ISBCS.t10 ISBCS.n12 2.96638
R17 ISBCS.t4 ISBCS.n9 2.96638
R18 ISBCS.n10 ISBCS.t4 2.96638
R19 ISBCS.t5 ISBCS.n1 2.96638
R20 ISBCS.n7 ISBCS.t15 2.96638
R21 ISBCS.n21 ISBCS.t9 2.96638
R22 ISBCS.n29 ISBCS.t14 2.96638
R23 ISBCS.t14 ISBCS.n28 2.96638
R24 ISBCS.t8 ISBCS.n25 2.96638
R25 ISBCS.n26 ISBCS.t8 2.96638
R26 ISBCS.t7 ISBCS.n19 2.96638
R27 ISBCS.n6 ISBCS.t5 2.52844
R28 ISBCS.n18 ISBCS.t11 2.52844
R29 ISBCS.t13 ISBCS.n18 2.52844
R30 ISBCS.t15 ISBCS.n6 2.52844
R31 ISBCS.n3 ISBCS.t12 2.52844
R32 ISBCS.n20 ISBCS.t7 2.52844
R33 ISBCS.t9 ISBCS.n20 2.52844
R34 ISBCS.n3 ISBCS.t6 2.52844
R35 ISBCS.n31 ISBCS.n30 1.5005
R36 ISBCS.n27 ISBCS.n24 1.5005
R37 ISBCS.n23 ISBCS.n22 1.5005
R38 ISBCS.n4 ISBCS.n0 1.5005
R39 ISBCS.n17 ISBCS.n16 1.5005
R40 ISBCS.n15 ISBCS.n14 1.5005
R41 ISBCS.n11 ISBCS.n8 1.5005
R42 ISBCS.n5 ISBCS.n4 1.19221
R43 ISBCS.n4 ISBCS.n2 1.16411
R44 ISBCS.n11 ISBCS.n10 0.88285
R45 ISBCS.n14 ISBCS.n9 0.88285
R46 ISBCS.n17 ISBCS.n7 0.88285
R47 ISBCS.n22 ISBCS.n1 0.88285
R48 ISBCS.n27 ISBCS.n26 0.88285
R49 ISBCS.n30 ISBCS.n25 0.88285
R50 ISBCS.n12 ISBCS.n11 0.858643
R51 ISBCS.n14 ISBCS.n13 0.858643
R52 ISBCS.n19 ISBCS.n17 0.858643
R53 ISBCS.n22 ISBCS.n21 0.858643
R54 ISBCS.n28 ISBCS.n27 0.858643
R55 ISBCS.n30 ISBCS.n29 0.858643
R56 ISBCS.n18 ISBCS.n2 0.367144
R57 ISBCS.n5 ISBCS.n3 0.365787
R58 ISBCS.n16 ISBCS.n0 0.210297
R59 ISBCS.n23 ISBCS.n0 0.207257
R60 ISBCS.n31 ISBCS.n24 0.1805
R61 ISBCS.n15 ISBCS.n8 0.179588
R62 ISBCS.n16 ISBCS.n15 0.0935405
R63 ISBCS.n24 ISBCS.n23 0.0935405
R64 ISBCS.n6 ISBCS.n5 0.0804816
R65 ISBCS.n20 ISBCS.n2 0.0795377
R66 VSS.t47 VSS.t10 997.681
R67 VSS.t4 VSS.t7 977.011
R68 VSS.t1 VSS.t46 727.312
R69 VSS.t50 VSS.t13 727.312
R70 VSS.n64 VSS.n4 697.422
R71 VSS.n66 VSS.n5 693.922
R72 VSS.n64 VSS.n5 693.645
R73 VSS.n66 VSS.n4 688.856
R74 VSS.t7 VSS.n4 484.967
R75 VSS.t10 VSS.n5 484.966
R76 VSS.n65 VSS.t48 445.214
R77 VSS.n65 VSS.t24 428.455
R78 VSS.t46 VSS.t4 32.3999
R79 VSS.t48 VSS.t1 32.3999
R80 VSS.t24 VSS.t50 32.3999
R81 VSS.t13 VSS.t47 32.3999
R82 VSS.n57 VSS.t14 3.3605
R83 VSS.n61 VSS.t25 3.3605
R84 VSS.n26 VSS.t2 3.3605
R85 VSS.n22 VSS.t29 3.3605
R86 VSS.n30 VSS.t52 3.3605
R87 VSS.n30 VSS.t57 3.3605
R88 VSS.n29 VSS.t55 3.3605
R89 VSS.n29 VSS.t49 3.3605
R90 VSS.n28 VSS.t53 3.3605
R91 VSS.n28 VSS.t56 3.3605
R92 VSS.n27 VSS.t51 3.3605
R93 VSS.n27 VSS.t54 3.3605
R94 VSS.n42 VSS.t37 3.3605
R95 VSS.n38 VSS.t41 3.3605
R96 VSS.n68 VSS.t27 3.3605
R97 VSS.n72 VSS.t5 3.3605
R98 VSS.t34 VSS.n73 2.53859
R99 VSS.t15 VSS.n43 2.53859
R100 VSS.n21 VSS.t30 2.53837
R101 VSS.n56 VSS.t32 2.53837
R102 VSS.n19 VSS.t30 2.52844
R103 VSS.t6 VSS.n17 2.52844
R104 VSS.n18 VSS.t6 2.52844
R105 VSS.t21 VSS.n15 2.52844
R106 VSS.n16 VSS.t21 2.52844
R107 VSS.t17 VSS.n12 2.52844
R108 VSS.n13 VSS.t17 2.52844
R109 VSS.t42 VSS.n0 2.52844
R110 VSS.n11 VSS.t42 2.52844
R111 VSS.n74 VSS.t34 2.52844
R112 VSS.n54 VSS.t32 2.52844
R113 VSS.t9 VSS.n52 2.52844
R114 VSS.n53 VSS.t9 2.52844
R115 VSS.t19 VSS.n50 2.52844
R116 VSS.n51 VSS.t19 2.52844
R117 VSS.t38 VSS.n47 2.52844
R118 VSS.n48 VSS.t38 2.52844
R119 VSS.t44 VSS.n45 2.52844
R120 VSS.n46 VSS.t44 2.52844
R121 VSS.n44 VSS.t15 2.52844
R122 VSS.n71 VSS.n70 2.1005
R123 VSS.n41 VSS.n40 2.1005
R124 VSS.n25 VSS.n24 2.1005
R125 VSS.n60 VSS.n59 2.1005
R126 VSS.n20 VSS.t31 1.6805
R127 VSS.n7 VSS.t8 1.6805
R128 VSS.n8 VSS.t22 1.6805
R129 VSS.n9 VSS.t18 1.6805
R130 VSS.n10 VSS.t43 1.6805
R131 VSS.n1 VSS.t35 1.6805
R132 VSS.n55 VSS.t33 1.6805
R133 VSS.n32 VSS.t11 1.6805
R134 VSS.n33 VSS.t20 1.6805
R135 VSS.n34 VSS.t39 1.6805
R136 VSS.n35 VSS.t45 1.6805
R137 VSS.n36 VSS.t16 1.6805
R138 VSS.n2 VSS.t3 1.26547
R139 VSS.n69 VSS.t26 1.26547
R140 VSS.n39 VSS.t40 1.26547
R141 VSS.n37 VSS.t36 1.26547
R142 VSS.n23 VSS.t28 1.26547
R143 VSS.n6 VSS.t0 1.26547
R144 VSS.n31 VSS.t23 1.26547
R145 VSS.n58 VSS.t12 1.26547
R146 VSS.t25 VSS.n60 1.2605
R147 VSS.n60 VSS.t14 1.2605
R148 VSS.n25 VSS.t29 1.2605
R149 VSS.t2 VSS.n25 1.2605
R150 VSS.n41 VSS.t41 1.2605
R151 VSS.t37 VSS.n41 1.2605
R152 VSS.t5 VSS.n71 1.2605
R153 VSS.n71 VSS.t27 1.2605
R154 VSS.n30 VSS.n29 0.240145
R155 VSS.n28 VSS.n27 0.240145
R156 VSS.n29 VSS.n28 0.207127
R157 VSS.n62 VSS.n30 0.160263
R158 VSS.n27 VSS.n3 0.160263
R159 VSS.n14 VSS.n4 0.0933571
R160 VSS.n49 VSS.n5 0.0917281
R161 VSS.n72 VSS.n2 0.069264
R162 VSS.n70 VSS.n2 0.069264
R163 VSS.n70 VSS.n69 0.069264
R164 VSS.n69 VSS.n68 0.069264
R165 VSS.n39 VSS.n38 0.069264
R166 VSS.n40 VSS.n39 0.069264
R167 VSS.n40 VSS.n37 0.069264
R168 VSS.n42 VSS.n37 0.069264
R169 VSS.n23 VSS.n22 0.0685756
R170 VSS.n24 VSS.n23 0.0685756
R171 VSS.n24 VSS.n6 0.0685756
R172 VSS.n26 VSS.n6 0.0685756
R173 VSS.n61 VSS.n31 0.0685756
R174 VSS.n59 VSS.n31 0.0685756
R175 VSS.n59 VSS.n58 0.0685756
R176 VSS.n58 VSS.n57 0.0685756
R177 VSS.n67 VSS.n66 0.0519852
R178 VSS.n66 VSS.n65 0.0519852
R179 VSS.n64 VSS.n63 0.0519852
R180 VSS.n65 VSS.n64 0.0519852
R181 VSS.n43 VSS.n42 0.0456011
R182 VSS.n57 VSS.n56 0.0451496
R183 VSS.n73 VSS.n72 0.0359944
R184 VSS.n22 VSS.n21 0.035639
R185 VSS.n19 VSS.n18 0.0192683
R186 VSS.n54 VSS.n53 0.0192569
R187 VSS.n45 VSS.n44 0.0192569
R188 VSS.n68 VSS.n67 0.0181966
R189 VSS.n63 VSS.n26 0.0180195
R190 VSS.n17 VSS.n16 0.0174024
R191 VSS.n12 VSS.n11 0.0174024
R192 VSS.n52 VSS.n51 0.0173921
R193 VSS.n47 VSS.n46 0.0173921
R194 VSS.n20 VSS.n19 0.0167439
R195 VSS.n18 VSS.n7 0.0167439
R196 VSS.n17 VSS.n7 0.0167439
R197 VSS.n16 VSS.n8 0.0167439
R198 VSS.n15 VSS.n8 0.0167439
R199 VSS.n13 VSS.n9 0.0167439
R200 VSS.n12 VSS.n9 0.0167439
R201 VSS.n11 VSS.n10 0.0167439
R202 VSS.n10 VSS.n0 0.0167439
R203 VSS.n74 VSS.n1 0.0167439
R204 VSS.n55 VSS.n54 0.016734
R205 VSS.n53 VSS.n32 0.016734
R206 VSS.n52 VSS.n32 0.016734
R207 VSS.n51 VSS.n33 0.016734
R208 VSS.n50 VSS.n33 0.016734
R209 VSS.n48 VSS.n34 0.016734
R210 VSS.n47 VSS.n34 0.016734
R211 VSS.n46 VSS.n35 0.016734
R212 VSS.n45 VSS.n35 0.016734
R213 VSS.n44 VSS.n36 0.016734
R214 VSS VSS.n0 0.0105976
R215 VSS VSS.n74 0.00917073
R216 VSS.n38 VSS.n3 0.00788202
R217 VSS.n62 VSS.n61 0.00780812
R218 VSS.n15 VSS.n14 0.00779878
R219 VSS.n21 VSS.n20 0.00681098
R220 VSS.n56 VSS.n55 0.00680713
R221 VSS.n73 VSS.n1 0.00659146
R222 VSS.n43 VSS.n36 0.00658775
R223 VSS.n49 VSS.n48 0.00592962
R224 VSS.n50 VSS.n49 0.00516179
R225 VSS.n14 VSS.n13 0.00329878
R226 VSS.n67 VSS.n3 0.00191573
R227 VSS.n63 VSS.n62 0.00190156
R228 a_n389_6663.t1 a_n389_6663.t0 9.72448
R229 INN INN.t0 17.8765
R230 INN INN.t1 3.47857
R231 VDD.n52 VDD.n23 614.001
R232 VDD.n52 VDD.n51 613.338
R233 VDD.n54 VDD.n23 607.537
R234 VDD.n54 VDD.n51 606.872
R235 VDD.t9 VDD.t30 338.731
R236 VDD.t3 VDD.t13 338.731
R237 VDD.t5 VDD.t9 260.622
R238 VDD.t0 VDD.t3 260.622
R239 VDD.t30 VDD.n23 167.008
R240 VDD.t13 VDD.n51 167.008
R241 VDD.n53 VDD.t5 156.792
R242 VDD.n53 VDD.t0 155.268
R243 VDD.n30 VDD.t24 3.20383
R244 VDD.t11 VDD.n5 3.20383
R245 VDD.t35 VDD.n4 3.20383
R246 VDD.n12 VDD.t45 3.20383
R247 VDD.n57 VDD.t4 3.20383
R248 VDD.n57 VDD.t8 3.20383
R249 VDD.n58 VDD.t1 3.20383
R250 VDD.n58 VDD.t6 3.20383
R251 VDD.n59 VDD.t2 3.20383
R252 VDD.n59 VDD.t7 3.20383
R253 VDD.n43 VDD.t28 3.20383
R254 VDD.n39 VDD.t18 3.20383
R255 VDD.n61 VDD.t39 3.20383
R256 VDD.n65 VDD.t47 3.20383
R257 VDD.t29 VDD.n13 2.55028
R258 VDD.t12 VDD.n31 2.55028
R259 VDD.t36 VDD.n66 2.55022
R260 VDD.t19 VDD.n44 2.55022
R261 VDD.n14 VDD.t29 2.54061
R262 VDD.n16 VDD.t42 2.54061
R263 VDD.t42 VDD.n15 2.54061
R264 VDD.n20 VDD.t32 2.54061
R265 VDD.t32 VDD.n17 2.54061
R266 VDD.t40 VDD.n0 2.54061
R267 VDD.n19 VDD.t40 2.54061
R268 VDD.n67 VDD.t36 2.54061
R269 VDD.n32 VDD.t12 2.54061
R270 VDD.n34 VDD.t25 2.54061
R271 VDD.t25 VDD.n33 2.54061
R272 VDD.n48 VDD.t15 2.54061
R273 VDD.t15 VDD.n35 2.54061
R274 VDD.t21 VDD.n46 2.54061
R275 VDD.n47 VDD.t21 2.54061
R276 VDD.n45 VDD.t19 2.54061
R277 VDD.n64 VDD.n63 1.73383
R278 VDD.n42 VDD.n41 1.73383
R279 VDD.n11 VDD.n10 1.73383
R280 VDD.n29 VDD.n28 1.73383
R281 VDD.n7 VDD.t31 1.60217
R282 VDD.n6 VDD.t43 1.60217
R283 VDD.n21 VDD.t33 1.60217
R284 VDD.n18 VDD.t41 1.60217
R285 VDD.n1 VDD.t37 1.60217
R286 VDD.n25 VDD.t14 1.60217
R287 VDD.n24 VDD.t26 1.60217
R288 VDD.n49 VDD.t16 1.60217
R289 VDD.n36 VDD.t22 1.60217
R290 VDD.n37 VDD.t20 1.60217
R291 VDD.n29 VDD.t11 1.4705
R292 VDD.t24 VDD.n29 1.4705
R293 VDD.t45 VDD.n11 1.4705
R294 VDD.n11 VDD.t35 1.4705
R295 VDD.n42 VDD.t18 1.4705
R296 VDD.t28 VDD.n42 1.4705
R297 VDD.t47 VDD.n64 1.4705
R298 VDD.n64 VDD.t39 1.4705
R299 VDD.n2 VDD.t46 1.27155
R300 VDD.n62 VDD.t38 1.27155
R301 VDD.n40 VDD.t17 1.27155
R302 VDD.n38 VDD.t27 1.27155
R303 VDD.n8 VDD.t44 1.27155
R304 VDD.n9 VDD.t34 1.27155
R305 VDD.n27 VDD.t10 1.27155
R306 VDD.n26 VDD.t23 1.27155
R307 VDD.n58 VDD.n57 0.249951
R308 VDD.n59 VDD.n58 0.249951
R309 VDD.n57 VDD.n56 0.192465
R310 VDD.n60 VDD.n59 0.192465
R311 VDD.n51 VDD.n50 0.119368
R312 VDD.n23 VDD.n22 0.119368
R313 VDD.n65 VDD.n2 0.0677787
R314 VDD.n63 VDD.n2 0.0677787
R315 VDD.n63 VDD.n62 0.0677787
R316 VDD.n62 VDD.n61 0.0677787
R317 VDD.n40 VDD.n39 0.0677787
R318 VDD.n41 VDD.n40 0.0677787
R319 VDD.n41 VDD.n38 0.0677787
R320 VDD.n43 VDD.n38 0.0677787
R321 VDD.n12 VDD.n8 0.0677787
R322 VDD.n10 VDD.n8 0.0677787
R323 VDD.n10 VDD.n9 0.0677787
R324 VDD.n9 VDD.n4 0.0677787
R325 VDD.n27 VDD.n5 0.0677787
R326 VDD.n28 VDD.n27 0.0677787
R327 VDD.n28 VDD.n26 0.0677787
R328 VDD.n30 VDD.n26 0.0677787
R329 VDD.n55 VDD.n54 0.0628762
R330 VDD.n54 VDD.n53 0.0628762
R331 VDD.n52 VDD.n3 0.061665
R332 VDD.n53 VDD.n52 0.061665
R333 VDD.n66 VDD.n65 0.0370902
R334 VDD.n44 VDD.n43 0.0370902
R335 VDD.n13 VDD.n12 0.0370902
R336 VDD.n31 VDD.n30 0.0370902
R337 VDD.n33 VDD.n32 0.0266202
R338 VDD.n46 VDD.n45 0.0266202
R339 VDD.n15 VDD.n14 0.0266202
R340 VDD.n35 VDD.n34 0.0203361
R341 VDD.n48 VDD.n47 0.0203361
R342 VDD.n17 VDD.n16 0.0203361
R343 VDD.n20 VDD.n19 0.0203361
R344 VDD.n32 VDD.n25 0.0167842
R345 VDD.n33 VDD.n24 0.0167842
R346 VDD.n34 VDD.n24 0.0167842
R347 VDD.n49 VDD.n48 0.0167842
R348 VDD.n47 VDD.n36 0.0167842
R349 VDD.n46 VDD.n36 0.0167842
R350 VDD.n45 VDD.n37 0.0167842
R351 VDD.n14 VDD.n7 0.0167842
R352 VDD.n15 VDD.n6 0.0167842
R353 VDD.n16 VDD.n6 0.0167842
R354 VDD.n21 VDD.n20 0.0167842
R355 VDD.n19 VDD.n18 0.0167842
R356 VDD.n18 VDD.n0 0.0167842
R357 VDD.n67 VDD.n1 0.0167842
R358 VDD VDD.n0 0.0160738
R359 VDD.n50 VDD.n35 0.014653
R360 VDD.n22 VDD.n17 0.014653
R361 VDD.n61 VDD.n60 0.0137787
R362 VDD.n56 VDD.n4 0.0137787
R363 VDD.n39 VDD.n3 0.0133852
R364 VDD.n55 VDD.n5 0.0133852
R365 VDD VDD.n67 0.0110464
R366 VDD.n44 VDD.n37 0.00716667
R367 VDD.n66 VDD.n1 0.00716667
R368 VDD.n31 VDD.n25 0.00711202
R369 VDD.n13 VDD.n7 0.00711202
R370 VDD.n50 VDD.n49 0.00263115
R371 VDD.n22 VDD.n21 0.00263115
R372 VDD.n60 VDD.n3 0.000893443
R373 VDD.n56 VDD.n55 0.000893443
R374 INN2 INN2.t1 18.1027
R375 INN2 INN2.t0 3.43357
R376 INP2 INP2.t0 3.81472
R377 INP2 INP2.t1 3.67076
R378 INP INP.t1 17.3056
R379 INP INP.t0 3.66129
C0 INP2 VDD 0.004028f
C1 a_941_6663# a_941_7622# 0.005385f
C2 INP2 ISBCS 1.14676f
C3 a_3947_6663# VDD 0.027393f
C4 a_3930_n291# ISBCS 0.134577f
C5 a_3947_7622# INN2 3.94e-19
C6 INN a_3947_7622# 0.010547f
C7 a_948_609# INP 0.029925f
C8 a_3947_6663# a_3947_5704# 0.005385f
C9 INP a_948_1385# 0.03013f
C10 a_3947_5704# VDD 0.03531f
C11 INP a_948_2285# 0.01763f
C12 ISBCS VDD 0.030253f
C13 a_948_1385# a_948_2285# 0.005955f
C14 a_948_n291# INP 0.007229f
C15 a_3930_609# a_3930_n291# 0.005955f
C16 ISBCS a_3930_1385# 0.159888f
C17 a_941_5704# VDD 0.03531f
C18 a_948_609# a_948_n291# 0.005955f
C19 VDD INN2 4.29151f
C20 INN VDD 2.65405f
C21 INP2 INP 0.32406f
C22 a_3947_5704# INN2 0.010168f
C23 INN a_3947_5704# 7.79e-19
C24 a_3930_n291# INP 0.010567f
C25 a_948_609# INP2 0.009765f
C26 INP2 a_948_1385# 0.009765f
C27 a_941_6663# VDD 0.027393f
C28 a_3930_609# ISBCS 0.159921f
C29 a_3930_2285# a_3930_1385# 0.005955f
C30 ISBCS a_3930_2285# 0.144473f
C31 INP2 a_948_2285# 0.00209f
C32 a_941_5704# INN2 0.032393f
C33 INN a_941_5704# 0.01055f
C34 a_941_7622# VDD 0.03531f
C35 INN INN2 4.90563f
C36 a_948_n291# INP2 0.001895f
C37 INP a_3930_1385# 8.06e-19
C38 INP ISBCS 10.9255f
C39 a_941_6663# a_941_5704# 0.005385f
C40 a_948_609# ISBCS 0.158537f
C41 ISBCS a_948_1385# 0.158318f
C42 a_941_6663# INN2 0.032392f
C43 a_3947_6663# a_3947_7622# 0.005385f
C44 ISBCS a_948_2285# 0.134725f
C45 a_3947_7622# VDD 0.03531f
C46 a_3930_609# INP 8.1e-19
C47 a_941_7622# INN2 0.042203f
C48 a_941_7622# INN 7.75e-19
C49 INP a_3930_2285# 8.06e-19
C50 a_948_n291# ISBCS 0.14436f
C51 INP2 VSS 1.59743f
C52 INP VSS 7.18598f
C53 ISBCS VSS 46.01309f
C54 INN VSS 9.654295f
C55 INN2 VSS 6.649196f
C56 VDD VSS 0.172401p
C57 a_3930_n291# VSS 0.036472f
C58 a_948_n291# VSS 0.036472f
C59 a_3930_609# VSS 0.02091f
C60 a_948_609# VSS 0.02091f
C61 a_3930_1385# VSS 0.020886f
C62 a_948_1385# VSS 0.02091f
C63 a_3930_2285# VSS 0.036472f
C64 a_948_2285# VSS 0.036472f
C65 INP.t1 VSS 5.06175f
C66 INP.t0 VSS 0.250813f
C67 INN2.t0 VSS 0.198984f
C68 INN2.t1 VSS 5.41973f
C69 VDD.n0 VSS 0.22353f
C70 VDD.t37 VSS 0.02503f
C71 VDD.n1 VSS 0.132032f
C72 VDD.t46 VSS 0.169724f
C73 VDD.n2 VSS 0.330319f
C74 VDD.t39 VSS 0.018381f
C75 VDD.n3 VSS 0.021563f
C76 VDD.n4 VSS 0.136455f
C77 VDD.n5 VSS 0.135816f
C78 VDD.t43 VSS 0.02503f
C79 VDD.n6 VSS 0.182634f
C80 VDD.t31 VSS 0.02503f
C81 VDD.n7 VSS 0.131745f
C82 VDD.t44 VSS 0.169724f
C83 VDD.n8 VSS 0.330319f
C84 VDD.t35 VSS 0.018381f
C85 VDD.t34 VSS 0.169724f
C86 VDD.n9 VSS 0.330319f
C87 VDD.n10 VSS 0.218506f
C88 VDD.n11 VSS 0.011731f
C89 VDD.t45 VSS 0.018381f
C90 VDD.n12 VSS 0.174311f
C91 VDD.n13 VSS 0.412458f
C92 VDD.t29 VSS 0.170729f
C93 VDD.n14 VSS 0.279019f
C94 VDD.n15 VSS 0.279019f
C95 VDD.t42 VSS 0.169711f
C96 VDD.n16 VSS 0.245956f
C97 VDD.n17 VSS 0.234743f
C98 VDD.t33 VSS 0.02503f
C99 VDD.t41 VSS 0.02503f
C100 VDD.n18 VSS 0.182634f
C101 VDD.t40 VSS 0.169711f
C102 VDD.n19 VSS 0.245956f
C103 VDD.t32 VSS 0.169711f
C104 VDD.n20 VSS 0.245956f
C105 VDD.n21 VSS 0.108169f
C106 VDD.n22 VSS 0.085677f
C107 VDD.n23 VSS 1.1143f
C108 VDD.t26 VSS 0.02503f
C109 VDD.n24 VSS 0.182634f
C110 VDD.t14 VSS 0.02503f
C111 VDD.n25 VSS 0.131745f
C112 VDD.t23 VSS 0.169724f
C113 VDD.n26 VSS 0.330319f
C114 VDD.t11 VSS 0.018381f
C115 VDD.t10 VSS 0.169724f
C116 VDD.n27 VSS 0.330319f
C117 VDD.n28 VSS 0.218506f
C118 VDD.n29 VSS 0.011731f
C119 VDD.t24 VSS 0.018381f
C120 VDD.n30 VSS 0.174311f
C121 VDD.n31 VSS 0.412458f
C122 VDD.t12 VSS 0.170729f
C123 VDD.n32 VSS 0.279019f
C124 VDD.n33 VSS 0.279019f
C125 VDD.t25 VSS 0.169711f
C126 VDD.n34 VSS 0.245956f
C127 VDD.n35 VSS 0.234743f
C128 VDD.t16 VSS 0.02503f
C129 VDD.t22 VSS 0.02503f
C130 VDD.n36 VSS 0.182634f
C131 VDD.t20 VSS 0.02503f
C132 VDD.n37 VSS 0.132032f
C133 VDD.t27 VSS 0.169724f
C134 VDD.n38 VSS 0.330319f
C135 VDD.t18 VSS 0.018381f
C136 VDD.n39 VSS 0.135816f
C137 VDD.t17 VSS 0.169724f
C138 VDD.n40 VSS 0.330319f
C139 VDD.n41 VSS 0.218506f
C140 VDD.n42 VSS 0.011731f
C141 VDD.t28 VSS 0.018381f
C142 VDD.n43 VSS 0.174311f
C143 VDD.n44 VSS 0.412178f
C144 VDD.t19 VSS 0.170722f
C145 VDD.n45 VSS 0.279019f
C146 VDD.n46 VSS 0.279019f
C147 VDD.t21 VSS 0.169711f
C148 VDD.n47 VSS 0.245956f
C149 VDD.t15 VSS 0.169711f
C150 VDD.n48 VSS 0.245956f
C151 VDD.n49 VSS 0.108169f
C152 VDD.n50 VSS 0.085677f
C153 VDD.n51 VSS 1.11408f
C154 VDD.t30 VSS 2.43248f
C155 VDD.t9 VSS 2.88265f
C156 VDD.t5 VSS 2.00759f
C157 VDD.n52 VSS 0.197128f
C158 VDD.t13 VSS 2.43248f
C159 VDD.t3 VSS 2.88265f
C160 VDD.t0 VSS 2.00026f
C161 VDD.n53 VSS 1.50088f
C162 VDD.n54 VSS 0.195044f
C163 VDD.n55 VSS 0.021563f
C164 VDD.n56 VSS 0.066776f
C165 VDD.t8 VSS 0.012515f
C166 VDD.t4 VSS 0.012515f
C167 VDD.n57 VSS 0.113777f
C168 VDD.t6 VSS 0.012515f
C169 VDD.t1 VSS 0.012515f
C170 VDD.n58 VSS 0.127125f
C171 VDD.t7 VSS 0.012515f
C172 VDD.t2 VSS 0.012515f
C173 VDD.n59 VSS 0.113777f
C174 VDD.n60 VSS 0.066776f
C175 VDD.n61 VSS 0.136455f
C176 VDD.t38 VSS 0.169724f
C177 VDD.n62 VSS 0.330319f
C178 VDD.n63 VSS 0.218506f
C179 VDD.n64 VSS 0.011731f
C180 VDD.t47 VSS 0.018381f
C181 VDD.n65 VSS 0.174311f
C182 VDD.n66 VSS 0.412178f
C183 VDD.t36 VSS 0.170722f
C184 VDD.n67 VSS 0.197079f
C185 INN.t1 VSS 0.23606f
C186 INN.t0 VSS 3.70135f
C187 a_n389_6663.t0 VSS 19.538f
C188 a_n389_6663.t1 VSS 16.362f
C189 ISBCS.t3 VSS 0.020838f
C190 ISBCS.n0 VSS 0.103861f
C191 ISBCS.n1 VSS 0.256662f
C192 ISBCS.t11 VSS 0.31814f
C193 ISBCS.n2 VSS 0.072615f
C194 ISBCS.t12 VSS 0.317363f
C195 ISBCS.t6 VSS 0.317363f
C196 ISBCS.n3 VSS 0.346678f
C197 ISBCS.n4 VSS 0.052027f
C198 ISBCS.n5 VSS 0.072917f
C199 ISBCS.t5 VSS 0.264098f
C200 ISBCS.n6 VSS 0.290443f
C201 ISBCS.t15 VSS 0.264098f
C202 ISBCS.n7 VSS 0.256662f
C203 ISBCS.t1 VSS 0.101213f
C204 ISBCS.n8 VSS 0.272154f
C205 ISBCS.n9 VSS 0.256662f
C206 ISBCS.t16 VSS 0.389255f
C207 ISBCS.t0 VSS 0.387701f
C208 ISBCS.t4 VSS 0.28117f
C209 ISBCS.n10 VSS 0.256662f
C210 ISBCS.n11 VSS 0.036537f
C211 ISBCS.n12 VSS 0.257861f
C212 ISBCS.t10 VSS 0.28117f
C213 ISBCS.n13 VSS 0.257861f
C214 ISBCS.n14 VSS 0.036537f
C215 ISBCS.n15 VSS 0.067851f
C216 ISBCS.n16 VSS 0.075508f
C217 ISBCS.n17 VSS 0.036537f
C218 ISBCS.n18 VSS 0.346416f
C219 ISBCS.t13 VSS 0.31814f
C220 ISBCS.n19 VSS 0.257861f
C221 ISBCS.t7 VSS 0.264098f
C222 ISBCS.n20 VSS 0.29042f
C223 ISBCS.t9 VSS 0.264098f
C224 ISBCS.n21 VSS 0.257861f
C225 ISBCS.n22 VSS 0.036537f
C226 ISBCS.n23 VSS 0.07475f
C227 ISBCS.n24 VSS 0.068079f
C228 ISBCS.n25 VSS 0.256662f
C229 ISBCS.t2 VSS 0.38531f
C230 ISBCS.t17 VSS 0.384486f
C231 ISBCS.t8 VSS 0.28117f
C232 ISBCS.n26 VSS 0.249989f
C233 ISBCS.n27 VSS 0.036537f
C234 ISBCS.n28 VSS 0.257861f
C235 ISBCS.t14 VSS 0.28117f
C236 ISBCS.n29 VSS 0.249661f
C237 ISBCS.n30 VSS 0.036537f
C238 ISBCS.n31 VSS 0.22612f
.ends

