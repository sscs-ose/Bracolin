* Extracted by KLayout with GF180MCU LVS runset on : 05/04/2024 12:28

.SUBCKT CM_block GND iref_un ibias iref iref_diff
M$1 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$2 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$3 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$7 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$8 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$9 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$10 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$11 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$12 iref_un ibias GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$13 GND ibias iref_un GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$14 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$15 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$16 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$17 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$18 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$19 iref ibias GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$20 iref_diff ibias GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$21 GND ibias iref_diff GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$22 GND ibias iref GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$23 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$24 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$25 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$26 iref_un ibias GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$27 GND ibias iref_diff GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$28 iref_diff ibias GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$29 GND ibias iref_diff GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$30 iref_diff ibias GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$31 GND ibias iref_un GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$32 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$33 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$34 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$35 iref ibias GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$36 iref_diff ibias GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$37 GND ibias iref_diff GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$38 GND ibias iref GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$39 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$40 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$41 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$42 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$43 ibias ibias GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$44 iref_un ibias GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$45 GND ibias iref_un GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$46 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$47 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$48 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$49 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$50 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$51 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$52 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$53 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$54 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$55 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$56 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
.ENDS CM_block
