** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/CurrentMirrors/CM_n_net.sch
.subckt CM_n_net IN OUT1 OUT2 VSS OUT3 OUT4 OUT5 OUT6 OUT7 OUT8 OUT9 OUT10 OUT11 OUT12
*.PININFO IN:B OUT1:B OUT2:B VSS:B OUT3:B OUT4:B OUT5:B OUT6:B OUT7:B OUT8:B OUT9:B OUT10:B OUT11:B
*+ OUT12:B
x1 IN OUT1 OUT2 VSS CM_nfets
x2 IN OUT3 OUT4 VSS CM_nfets
x4 IN OUT9 OUT10 VSS CM_nfets
x5 IN OUT7 OUT8 VSS CM_nfets
x3 IN OUT5 OUT6 VSS CM_nfets
x7 IN OUT11 OUT12 VSS CM_nfets
.ends

* expanding   symbol:  CurrentMirrors/CM_nfets.sym # of pins=4
** sym_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/CurrentMirrors/CM_nfets.sym
** sch_path: /home/gmaranhao/Desktop/Bracolin/TIA_Filter/CurrentMirrors/CM_nfets.sch
.subckt CM_nfets IN OUT1 OUT2 VSS
*.PININFO IN:B OUT1:B OUT2:B VSS:B
M2[1] IN IN VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M2[2] IN IN VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M2[3] IN IN VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M2[4] IN IN VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M2[5] IN IN VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M2[6] IN IN VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M2 OUT1 IN net3 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M11 net4 IN net6 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M12 net6 IN net7 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M13 net7 IN net8 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M14 net8 IN net9 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M15 net9 IN net10 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M16 net10 IN net11 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M17 net11 IN net12 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M18 net12 IN net13 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M19 net13 IN net14 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M20 net14 IN net1 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M21 net1 IN net15 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M22 net15 IN net16 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M23 net16 IN net17 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M24 net17 IN net18 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M25 net18 IN net19 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M26 net19 IN net20 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M27 net20 IN net21 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M28 net21 IN net22 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M29 net22 IN net23 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M30 net23 IN net2 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M31 net2 IN net24 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M32 net24 IN net25 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M33 net25 IN net26 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M34 net26 IN net27 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M35 net27 IN net28 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M36 net28 IN net29 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1 net29 IN net30 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M37 net30 IN net31 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M38 net31 IN net32 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M9 net32 IN VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M5 net3 IN net4 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M8 net5 IN net33 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M10 net33 IN net34 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M39 net34 IN net35 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M40 net35 IN net36 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M41 net36 IN net37 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M42 net37 IN net38 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M43 net38 IN net39 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M44 net39 IN net40 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M45 net40 IN net41 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M46 net41 IN VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M47 OUT2 IN net42 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M48 net42 IN net43 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M49 net43 IN net44 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M50 net44 IN net45 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M51 net45 IN net46 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M52 net46 IN net5 VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[1] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[2] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[3] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[4] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[5] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[6] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[7] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[8] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[9] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[10] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[11] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[12] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[13] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[14] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[15] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[16] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[17] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[18] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[19] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[20] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[21] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[22] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[23] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[24] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[25] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[26] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[27] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[28] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[29] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[30] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[31] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[32] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[33] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
M1[34] VSS VSS VSS VSS nfet_03v3 L=2u W=2u nf=1 m=1
.ends

.end
