* NGSPICE file created from CM_input.ext - technology: gf180mcuD

.subckt CM_input_pex IN IN2 IP2 IP ISBCS VDD VSS
X0 a_3930_2285# ISBCS.t4 VSS.t11 VSS.t2 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X1 a_948_n291# ISBCS.t0 ISBCS.t1 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X2 IN.t0 a_n389_6663.t0 a_3947_7622# VDD.t9 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X3 a_3930_609# ISBCS.t5 VSS.t10 VSS.t2 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X4 IN2.t0 a_n389_6663.t0 a_3947_5704# VDD.t9 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X5 VSS.t57 VSS.t56 VSS.t57 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X6 VSS.t55 VSS.t54 VSS.t55 VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X7 VSS.t53 VSS.t52 VSS.t53 VSS.t36 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X8 a_n389_6663.t0 ISBCS.t6 a_3930_609# VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X9 VDD.t55 VDD.t54 VDD.t55 VDD.t9 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X10 VSS.t9 ISBCS.t7 a_948_1385# VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X11 a_n389_6663.t2 a_n389_6663.t0 a_3947_6663# VDD.t9 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X12 a_3930_n291# ISBCS.t8 VSS.t8 VSS.t2 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X13 VDD.t53 VDD.t52 VDD.t53 VDD.t9 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X14 VSS.t7 ISBCS.t9 a_948_609# VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X15 VSS.t51 VSS.t50 VSS.t51 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X16 VSS.t49 VSS.t48 VSS.t49 VSS.t25 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X17 VSS.t47 VSS.t46 VSS.t47 VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X18 a_3947_7622# a_n389_6663.t0 VDD.t8 VDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X19 VDD.t51 VDD.t49 VDD.t51 VDD.t50 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X20 VSS.t45 VSS.t44 VSS.t45 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X21 VSS.t43 VSS.t42 VSS.t43 VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X22 a_3947_5704# a_n389_6663.t0 VDD.t7 VDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X23 VSS.t41 VSS.t40 VSS.t41 VSS.t16 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X24 VSS.t6 ISBCS.t10 a_948_2285# VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X25 VDD.t48 VDD.t46 VDD.t48 VDD.t47 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X26 a_948_609# ISBCS.t11 IP2.t0 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X27 VSS.t39 VSS.t38 VSS.t39 VSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X28 a_941_7622# a_n389_6663.t0 IN2.t1 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X29 VDD.t45 VDD.t44 VDD.t45 VDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X30 a_n389_6663.t0 ISBCS.t12 a_3930_1385# VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X31 a_3947_6663# a_n389_6663.t0 VDD.t6 VDD.t5 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X32 VDD.t43 VDD.t41 VDD.t43 VDD.t42 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X33 VDD.t40 VDD.t39 VDD.t40 VDD.t5 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X34 VDD.t38 VDD.t36 VDD.t38 VDD.t37 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X35 a_941_5704# a_n389_6663.t0 IN.t1 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X36 VDD.t35 VDD.t33 VDD.t35 VDD.t34 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X37 a_948_1385# ISBCS.t13 IP2.t1 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X38 VDD.t4 a_n389_6663.t0 a_941_7622# VDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X39 VDD.t32 VDD.t31 VDD.t32 VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X40 VSS.t37 VSS.t35 VSS.t37 VSS.t36 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X41 VSS.t5 ISBCS.t14 a_948_n291# VSS.t4 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X42 VDD.t30 VDD.t28 VDD.t30 VDD.t29 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X43 a_941_6663# a_n389_6663.t0 a_n389_6663.t0 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=6u
X44 VSS.t34 VSS.t33 VSS.t34 VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X45 VDD.t27 VDD.t26 VDD.t27 VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X46 VDD.t25 VDD.t23 VDD.t25 VDD.t24 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X47 VDD.t2 a_n389_6663.t0 a_941_5704# VDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X48 VSS.t32 VSS.t31 VSS.t32 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X49 VDD.t22 VDD.t20 VDD.t22 VDD.t21 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X50 VDD.t19 VDD.t18 VDD.t19 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X51 VDD.t17 VDD.t15 VDD.t17 VDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X52 VDD.t1 a_n389_6663.t0 a_941_6663# VDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=6u
X53 ISBCS.t3 ISBCS.t2 a_3930_2285# VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X54 a_3930_1385# ISBCS.t15 VSS.t3 VSS.t2 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X55 VSS.t30 VSS.t29 VSS.t30 VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X56 VSS.t28 VSS.t27 VSS.t28 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X57 VDD.t14 VDD.t12 VDD.t14 VDD.t13 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=6u
X58 VDD.t11 VDD.t10 VDD.t11 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=6u
X59 VSS.t26 VSS.t24 VSS.t26 VSS.t25 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X60 a_948_2285# ISBCS.t16 IP.t1 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=6u
X61 VSS.t23 VSS.t21 VSS.t23 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X62 VSS.t20 VSS.t18 VSS.t20 VSS.t19 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
X63 IP.t0 ISBCS.t17 a_3930_n291# VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=6u
X64 VSS.t17 VSS.t15 VSS.t17 VSS.t16 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=6u
X65 VSS.t14 VSS.t12 VSS.t14 VSS.t13 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=6u
R0 ISBCS.n8 ISBCS.t3 10.2879
R1 ISBCS ISBCS.n31 6.52263
R2 ISBCS.t2 ISBCS.n9 4.39661
R3 ISBCS.n7 ISBCS.t12 4.39661
R4 ISBCS.t6 ISBCS.n1 4.39661
R5 ISBCS.t17 ISBCS.n25 4.39661
R6 ISBCS.n10 ISBCS.t2 4.39661
R7 ISBCS.n26 ISBCS.t17 4.39661
R8 ISBCS.n13 ISBCS.t16 4.39651
R9 ISBCS.n12 ISBCS.t16 4.39651
R10 ISBCS.n21 ISBCS.t11 4.39651
R11 ISBCS.n19 ISBCS.t13 4.39651
R12 ISBCS.n29 ISBCS.t0 4.39651
R13 ISBCS.n28 ISBCS.t0 4.39651
R14 ISBCS ISBCS.t1 3.79155
R15 ISBCS.n13 ISBCS.t10 2.96638
R16 ISBCS.t10 ISBCS.n12 2.96638
R17 ISBCS.t4 ISBCS.n9 2.96638
R18 ISBCS.n10 ISBCS.t4 2.96638
R19 ISBCS.t5 ISBCS.n1 2.96638
R20 ISBCS.n7 ISBCS.t15 2.96638
R21 ISBCS.n21 ISBCS.t9 2.96638
R22 ISBCS.n29 ISBCS.t14 2.96638
R23 ISBCS.t14 ISBCS.n28 2.96638
R24 ISBCS.t8 ISBCS.n25 2.96638
R25 ISBCS.n26 ISBCS.t8 2.96638
R26 ISBCS.t7 ISBCS.n19 2.96638
R27 ISBCS.n6 ISBCS.t5 2.52844
R28 ISBCS.n18 ISBCS.t11 2.52844
R29 ISBCS.t13 ISBCS.n18 2.52844
R30 ISBCS.t15 ISBCS.n6 2.52844
R31 ISBCS.n3 ISBCS.t12 2.52844
R32 ISBCS.n20 ISBCS.t7 2.52844
R33 ISBCS.t9 ISBCS.n20 2.52844
R34 ISBCS.n3 ISBCS.t6 2.52844
R35 ISBCS.n31 ISBCS.n30 1.5005
R36 ISBCS.n27 ISBCS.n24 1.5005
R37 ISBCS.n23 ISBCS.n22 1.5005
R38 ISBCS.n4 ISBCS.n0 1.5005
R39 ISBCS.n17 ISBCS.n16 1.5005
R40 ISBCS.n15 ISBCS.n14 1.5005
R41 ISBCS.n11 ISBCS.n8 1.5005
R42 ISBCS.n5 ISBCS.n4 1.19221
R43 ISBCS.n4 ISBCS.n2 1.16411
R44 ISBCS.n11 ISBCS.n10 0.88285
R45 ISBCS.n14 ISBCS.n9 0.88285
R46 ISBCS.n17 ISBCS.n7 0.88285
R47 ISBCS.n22 ISBCS.n1 0.88285
R48 ISBCS.n27 ISBCS.n26 0.88285
R49 ISBCS.n30 ISBCS.n25 0.88285
R50 ISBCS.n12 ISBCS.n11 0.858643
R51 ISBCS.n14 ISBCS.n13 0.858643
R52 ISBCS.n19 ISBCS.n17 0.858643
R53 ISBCS.n22 ISBCS.n21 0.858643
R54 ISBCS.n28 ISBCS.n27 0.858643
R55 ISBCS.n30 ISBCS.n29 0.858643
R56 ISBCS.n18 ISBCS.n2 0.367144
R57 ISBCS.n5 ISBCS.n3 0.365787
R58 ISBCS.n16 ISBCS.n0 0.210297
R59 ISBCS.n23 ISBCS.n0 0.207257
R60 ISBCS.n31 ISBCS.n24 0.1805
R61 ISBCS.n15 ISBCS.n8 0.179588
R62 ISBCS.n16 ISBCS.n15 0.0935405
R63 ISBCS.n24 ISBCS.n23 0.0935405
R64 ISBCS.n6 ISBCS.n5 0.0804816
R65 ISBCS.n20 ISBCS.n2 0.0795377
R66 VSS.t1 VSS.t22 992.053
R67 VSS.t16 VSS.t19 971.501
R68 VSS.t13 VSS.t0 723.211
R69 VSS.t4 VSS.t25 723.211
R70 VSS.n64 VSS.n4 697.422
R71 VSS.n66 VSS.n5 693.922
R72 VSS.n64 VSS.n5 693.645
R73 VSS.n66 VSS.n4 688.856
R74 VSS.t19 VSS.n4 482.233
R75 VSS.t22 VSS.n5 482.231
R76 VSS.n65 VSS.t2 442.702
R77 VSS.n65 VSS.t36 426.038
R78 VSS.t0 VSS.t16 32.2172
R79 VSS.t2 VSS.t13 32.2172
R80 VSS.t36 VSS.t4 32.2172
R81 VSS.t25 VSS.t1 32.2172
R82 VSS.n57 VSS.t26 3.3605
R83 VSS.n61 VSS.t37 3.3605
R84 VSS.n26 VSS.t14 3.3605
R85 VSS.n22 VSS.t41 3.3605
R86 VSS.n30 VSS.t6 3.3605
R87 VSS.n30 VSS.t11 3.3605
R88 VSS.n29 VSS.t9 3.3605
R89 VSS.n29 VSS.t3 3.3605
R90 VSS.n28 VSS.t7 3.3605
R91 VSS.n28 VSS.t10 3.3605
R92 VSS.n27 VSS.t5 3.3605
R93 VSS.n27 VSS.t8 3.3605
R94 VSS.n42 VSS.t49 3.3605
R95 VSS.n38 VSS.t53 3.3605
R96 VSS.n68 VSS.t39 3.3605
R97 VSS.n72 VSS.t17 3.3605
R98 VSS.t46 VSS.n73 2.53859
R99 VSS.t27 VSS.n43 2.53859
R100 VSS.n21 VSS.t42 2.53837
R101 VSS.n56 VSS.t44 2.53837
R102 VSS.n19 VSS.t42 2.52844
R103 VSS.t18 VSS.n17 2.52844
R104 VSS.n18 VSS.t18 2.52844
R105 VSS.t33 VSS.n15 2.52844
R106 VSS.n16 VSS.t33 2.52844
R107 VSS.t29 VSS.n12 2.52844
R108 VSS.n13 VSS.t29 2.52844
R109 VSS.t54 VSS.n0 2.52844
R110 VSS.n11 VSS.t54 2.52844
R111 VSS.n74 VSS.t46 2.52844
R112 VSS.n54 VSS.t44 2.52844
R113 VSS.t21 VSS.n52 2.52844
R114 VSS.n53 VSS.t21 2.52844
R115 VSS.t31 VSS.n50 2.52844
R116 VSS.n51 VSS.t31 2.52844
R117 VSS.t50 VSS.n47 2.52844
R118 VSS.n48 VSS.t50 2.52844
R119 VSS.t56 VSS.n45 2.52844
R120 VSS.n46 VSS.t56 2.52844
R121 VSS.n44 VSS.t27 2.52844
R122 VSS.n71 VSS.n70 2.1005
R123 VSS.n41 VSS.n40 2.1005
R124 VSS.n25 VSS.n24 2.1005
R125 VSS.n60 VSS.n59 2.1005
R126 VSS.n20 VSS.t43 1.6805
R127 VSS.n7 VSS.t20 1.6805
R128 VSS.n8 VSS.t34 1.6805
R129 VSS.n9 VSS.t30 1.6805
R130 VSS.n10 VSS.t55 1.6805
R131 VSS.n1 VSS.t47 1.6805
R132 VSS.n55 VSS.t45 1.6805
R133 VSS.n32 VSS.t23 1.6805
R134 VSS.n33 VSS.t32 1.6805
R135 VSS.n34 VSS.t51 1.6805
R136 VSS.n35 VSS.t57 1.6805
R137 VSS.n36 VSS.t28 1.6805
R138 VSS.n2 VSS.t15 1.26547
R139 VSS.n69 VSS.t38 1.26547
R140 VSS.n39 VSS.t52 1.26547
R141 VSS.n37 VSS.t48 1.26547
R142 VSS.n23 VSS.t40 1.26547
R143 VSS.n6 VSS.t12 1.26547
R144 VSS.n31 VSS.t35 1.26547
R145 VSS.n58 VSS.t24 1.26547
R146 VSS.t37 VSS.n60 1.2605
R147 VSS.n60 VSS.t26 1.2605
R148 VSS.n25 VSS.t41 1.2605
R149 VSS.t14 VSS.n25 1.2605
R150 VSS.n41 VSS.t53 1.2605
R151 VSS.t49 VSS.n41 1.2605
R152 VSS.t17 VSS.n71 1.2605
R153 VSS.n71 VSS.t39 1.2605
R154 VSS.n30 VSS.n29 0.240145
R155 VSS.n28 VSS.n27 0.240145
R156 VSS.n29 VSS.n28 0.207127
R157 VSS.n62 VSS.n30 0.160263
R158 VSS.n27 VSS.n3 0.160263
R159 VSS.n14 VSS.n4 0.0933571
R160 VSS.n49 VSS.n5 0.0917281
R161 VSS.n72 VSS.n2 0.069264
R162 VSS.n70 VSS.n2 0.069264
R163 VSS.n70 VSS.n69 0.069264
R164 VSS.n69 VSS.n68 0.069264
R165 VSS.n39 VSS.n38 0.069264
R166 VSS.n40 VSS.n39 0.069264
R167 VSS.n40 VSS.n37 0.069264
R168 VSS.n42 VSS.n37 0.069264
R169 VSS.n23 VSS.n22 0.0685756
R170 VSS.n24 VSS.n23 0.0685756
R171 VSS.n24 VSS.n6 0.0685756
R172 VSS.n26 VSS.n6 0.0685756
R173 VSS.n61 VSS.n31 0.0685756
R174 VSS.n59 VSS.n31 0.0685756
R175 VSS.n59 VSS.n58 0.0685756
R176 VSS.n58 VSS.n57 0.0685756
R177 VSS.n67 VSS.n66 0.0519852
R178 VSS.n66 VSS.n65 0.0519852
R179 VSS.n64 VSS.n63 0.0519852
R180 VSS.n65 VSS.n64 0.0519852
R181 VSS.n43 VSS.n42 0.0456011
R182 VSS.n57 VSS.n56 0.0451496
R183 VSS.n73 VSS.n72 0.0359944
R184 VSS.n22 VSS.n21 0.035639
R185 VSS.n19 VSS.n18 0.0192683
R186 VSS.n54 VSS.n53 0.0192569
R187 VSS.n45 VSS.n44 0.0192569
R188 VSS.n68 VSS.n67 0.0181966
R189 VSS.n63 VSS.n26 0.0180195
R190 VSS.n17 VSS.n16 0.0174024
R191 VSS.n12 VSS.n11 0.0174024
R192 VSS.n52 VSS.n51 0.0173921
R193 VSS.n47 VSS.n46 0.0173921
R194 VSS.n20 VSS.n19 0.0167439
R195 VSS.n18 VSS.n7 0.0167439
R196 VSS.n17 VSS.n7 0.0167439
R197 VSS.n16 VSS.n8 0.0167439
R198 VSS.n15 VSS.n8 0.0167439
R199 VSS.n13 VSS.n9 0.0167439
R200 VSS.n12 VSS.n9 0.0167439
R201 VSS.n11 VSS.n10 0.0167439
R202 VSS.n10 VSS.n0 0.0167439
R203 VSS.n74 VSS.n1 0.0167439
R204 VSS.n55 VSS.n54 0.016734
R205 VSS.n53 VSS.n32 0.016734
R206 VSS.n52 VSS.n32 0.016734
R207 VSS.n51 VSS.n33 0.016734
R208 VSS.n50 VSS.n33 0.016734
R209 VSS.n48 VSS.n34 0.016734
R210 VSS.n47 VSS.n34 0.016734
R211 VSS.n46 VSS.n35 0.016734
R212 VSS.n45 VSS.n35 0.016734
R213 VSS.n44 VSS.n36 0.016734
R214 VSS VSS.n0 0.0105976
R215 VSS VSS.n74 0.00917073
R216 VSS.n38 VSS.n3 0.00788202
R217 VSS.n62 VSS.n61 0.00780812
R218 VSS.n15 VSS.n14 0.00779878
R219 VSS.n21 VSS.n20 0.00681098
R220 VSS.n56 VSS.n55 0.00680713
R221 VSS.n73 VSS.n1 0.00659146
R222 VSS.n43 VSS.n36 0.00658775
R223 VSS.n49 VSS.n48 0.00592962
R224 VSS.n50 VSS.n49 0.00516179
R225 VSS.n14 VSS.n13 0.00329878
R226 VSS.n67 VSS.n3 0.00191573
R227 VSS.n63 VSS.n62 0.00190156
R228 a_n389_6663.t2 a_n389_6663.t0 9.72448
R229 IN IN.t0 17.8765
R230 IN IN.t1 3.47857
R231 VDD.n54 VDD.n23 614.001
R232 VDD.n54 VDD.n51 613.338
R233 VDD.n58 VDD.n23 607.537
R234 VDD.n58 VDD.n51 606.872
R235 VDD.t50 VDD.t34 575.871
R236 VDD.t47 VDD.t42 575.871
R237 VDD.t29 VDD.t13 575.871
R238 VDD.t24 VDD.t21 575.871
R239 VDD.n53 VDD.t47 513.138
R240 VDD.n56 VDD.t24 513.138
R241 VDD.n52 VDD.t50 493.298
R242 VDD.n55 VDD.t29 493.298
R243 VDD.t5 VDD.t9 230.343
R244 VDD.t0 VDD.t3 230.343
R245 VDD.t9 VDD.n53 143.458
R246 VDD.t3 VDD.n56 143.458
R247 VDD.n57 VDD.t5 138.577
R248 VDD.n57 VDD.t0 137.228
R249 VDD.t37 VDD.n52 20.912
R250 VDD.t16 VDD.n55 20.912
R251 VDD.n30 VDD.t27 3.20383
R252 VDD.t11 VDD.n5 3.20383
R253 VDD.t40 VDD.n4 3.20383
R254 VDD.n12 VDD.t53 3.20383
R255 VDD.n61 VDD.t4 3.20383
R256 VDD.n61 VDD.t8 3.20383
R257 VDD.n62 VDD.t1 3.20383
R258 VDD.n62 VDD.t6 3.20383
R259 VDD.n63 VDD.t2 3.20383
R260 VDD.n63 VDD.t7 3.20383
R261 VDD.n43 VDD.t32 3.20383
R262 VDD.n39 VDD.t19 3.20383
R263 VDD.n65 VDD.t45 3.20383
R264 VDD.n69 VDD.t55 3.20383
R265 VDD.t33 VDD.n13 2.55028
R266 VDD.t12 VDD.n31 2.55028
R267 VDD.t41 VDD.n70 2.55022
R268 VDD.t20 VDD.n44 2.55022
R269 VDD.n14 VDD.t33 2.54061
R270 VDD.n16 VDD.t49 2.54061
R271 VDD.t49 VDD.n15 2.54061
R272 VDD.n20 VDD.t36 2.54061
R273 VDD.t36 VDD.n17 2.54061
R274 VDD.t46 VDD.n0 2.54061
R275 VDD.n19 VDD.t46 2.54061
R276 VDD.n71 VDD.t41 2.54061
R277 VDD.n32 VDD.t12 2.54061
R278 VDD.n34 VDD.t28 2.54061
R279 VDD.t28 VDD.n33 2.54061
R280 VDD.n48 VDD.t15 2.54061
R281 VDD.t15 VDD.n35 2.54061
R282 VDD.t23 VDD.n46 2.54061
R283 VDD.n47 VDD.t23 2.54061
R284 VDD.n45 VDD.t20 2.54061
R285 VDD.n68 VDD.n67 1.73383
R286 VDD.n42 VDD.n41 1.73383
R287 VDD.n11 VDD.n10 1.73383
R288 VDD.n29 VDD.n28 1.73383
R289 VDD.n7 VDD.t35 1.60217
R290 VDD.n6 VDD.t51 1.60217
R291 VDD.n21 VDD.t38 1.60217
R292 VDD.n18 VDD.t48 1.60217
R293 VDD.n1 VDD.t43 1.60217
R294 VDD.n25 VDD.t14 1.60217
R295 VDD.n24 VDD.t30 1.60217
R296 VDD.n49 VDD.t17 1.60217
R297 VDD.n36 VDD.t25 1.60217
R298 VDD.n37 VDD.t22 1.60217
R299 VDD.n29 VDD.t11 1.4705
R300 VDD.t27 VDD.n29 1.4705
R301 VDD.t53 VDD.n11 1.4705
R302 VDD.n11 VDD.t40 1.4705
R303 VDD.n42 VDD.t19 1.4705
R304 VDD.t32 VDD.n42 1.4705
R305 VDD.t55 VDD.n68 1.4705
R306 VDD.n68 VDD.t45 1.4705
R307 VDD.n2 VDD.t54 1.27155
R308 VDD.n66 VDD.t44 1.27155
R309 VDD.n40 VDD.t18 1.27155
R310 VDD.n38 VDD.t31 1.27155
R311 VDD.n8 VDD.t52 1.27155
R312 VDD.n9 VDD.t39 1.27155
R313 VDD.n27 VDD.t10 1.27155
R314 VDD.n26 VDD.t26 1.27155
R315 VDD.n53 VDD.t37 1.07289
R316 VDD.n56 VDD.t16 1.07289
R317 VDD.n62 VDD.n61 0.249951
R318 VDD.n63 VDD.n62 0.249951
R319 VDD.n61 VDD.n60 0.192465
R320 VDD.n64 VDD.n63 0.192465
R321 VDD.n51 VDD.n50 0.119368
R322 VDD.n55 VDD.n51 0.119368
R323 VDD.n23 VDD.n22 0.119368
R324 VDD.n52 VDD.n23 0.119368
R325 VDD.n69 VDD.n2 0.0677787
R326 VDD.n67 VDD.n2 0.0677787
R327 VDD.n67 VDD.n66 0.0677787
R328 VDD.n66 VDD.n65 0.0677787
R329 VDD.n40 VDD.n39 0.0677787
R330 VDD.n41 VDD.n40 0.0677787
R331 VDD.n41 VDD.n38 0.0677787
R332 VDD.n43 VDD.n38 0.0677787
R333 VDD.n12 VDD.n8 0.0677787
R334 VDD.n10 VDD.n8 0.0677787
R335 VDD.n10 VDD.n9 0.0677787
R336 VDD.n9 VDD.n4 0.0677787
R337 VDD.n27 VDD.n5 0.0677787
R338 VDD.n28 VDD.n27 0.0677787
R339 VDD.n28 VDD.n26 0.0677787
R340 VDD.n30 VDD.n26 0.0677787
R341 VDD.n59 VDD.n58 0.0628762
R342 VDD.n58 VDD.n57 0.0628762
R343 VDD.n54 VDD.n3 0.061665
R344 VDD.n57 VDD.n54 0.061665
R345 VDD.n70 VDD.n69 0.0370902
R346 VDD.n44 VDD.n43 0.0370902
R347 VDD.n13 VDD.n12 0.0370902
R348 VDD.n31 VDD.n30 0.0370902
R349 VDD.n33 VDD.n32 0.0266202
R350 VDD.n46 VDD.n45 0.0266202
R351 VDD.n15 VDD.n14 0.0266202
R352 VDD.n35 VDD.n34 0.0203361
R353 VDD.n48 VDD.n47 0.0203361
R354 VDD.n17 VDD.n16 0.0203361
R355 VDD.n20 VDD.n19 0.0203361
R356 VDD.n32 VDD.n25 0.0167842
R357 VDD.n33 VDD.n24 0.0167842
R358 VDD.n34 VDD.n24 0.0167842
R359 VDD.n49 VDD.n48 0.0167842
R360 VDD.n47 VDD.n36 0.0167842
R361 VDD.n46 VDD.n36 0.0167842
R362 VDD.n45 VDD.n37 0.0167842
R363 VDD.n14 VDD.n7 0.0167842
R364 VDD.n15 VDD.n6 0.0167842
R365 VDD.n16 VDD.n6 0.0167842
R366 VDD.n21 VDD.n20 0.0167842
R367 VDD.n19 VDD.n18 0.0167842
R368 VDD.n18 VDD.n0 0.0167842
R369 VDD.n71 VDD.n1 0.0167842
R370 VDD VDD.n0 0.0160738
R371 VDD.n50 VDD.n35 0.014653
R372 VDD.n22 VDD.n17 0.014653
R373 VDD.n65 VDD.n64 0.0137787
R374 VDD.n60 VDD.n4 0.0137787
R375 VDD.n39 VDD.n3 0.0133852
R376 VDD.n59 VDD.n5 0.0133852
R377 VDD VDD.n71 0.0110464
R378 VDD.n44 VDD.n37 0.00716667
R379 VDD.n70 VDD.n1 0.00716667
R380 VDD.n31 VDD.n25 0.00711202
R381 VDD.n13 VDD.n7 0.00711202
R382 VDD.n50 VDD.n49 0.00263115
R383 VDD.n22 VDD.n21 0.00263115
R384 VDD.n64 VDD.n3 0.000893443
R385 VDD.n60 VDD.n59 0.000893443
R386 IN2 IN2.t1 18.1027
R387 IN2 IN2.t0 3.43357
R388 IP2 IP2.t1 3.81472
R389 IP2 IP2.t0 3.67076
R390 IP IP.t1 17.3056
R391 IP IP.t0 3.66129
C0 ISBCS IP2 1.14676f
C1 IN IN2 4.90563f
C2 IP ISBCS 10.9255f
C3 VDD IN2 4.41958f
C4 IN VDD 2.66124f
C5 IP2 VSS 1.59743f
C6 IP VSS 7.18598f
C7 ISBCS VSS 46.01309f
C8 IN VSS 9.647114f
C9 IN2 VSS 6.571406f
C10 VDD VSS 0.190456p
C11 IP.t1 VSS 5.06175f
C12 IN2.t1 VSS 5.46769f
C13 VDD.n53 VSS 1.17735f
C14 VDD.t9 VSS 2.26658f
C15 VDD.t5 VSS 2.23697f
C16 VDD.n56 VSS 1.17735f
C17 VDD.t3 VSS 2.26658f
C18 VDD.t0 VSS 2.22881f
C19 VDD.n57 VSS 1.67237f
C20 IN.t0 VSS 3.70135f
C21 a_n389_6663.t0 VSS 19.538f
C22 a_n389_6663.t2 VSS 16.362f
.ends

