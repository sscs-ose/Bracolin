magic
tech gf180mcuC
magscale 1 5
timestamp 1698433737
<< checkpaint >>
rect 650 8796 3100 8826
rect 650 1814 3520 8796
rect 650 1784 3940 1814
rect 650 1678 4360 1784
rect -1030 -730 4360 1678
rect -1000 -880 4360 -730
rect -1000 -2600 1100 -880
rect 1490 -910 4360 -880
rect 1910 -940 4360 -910
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
rect 0 -1200 100 -1100
rect 0 -1400 100 -1300
rect 0 -1600 100 -1500
use nfet_03v3_QVD5W3  M1
timestamp 0
transform 1 0 195 0 1 474
box -225 -204 225 204
use nfet_03v3_QVD5W3  M2
timestamp 0
transform 1 0 1035 0 1 414
box -225 -204 225 204
use pfet_03v3_ANSKCD  M3
timestamp 0
transform 1 0 615 0 1 444
box -225 -204 225 204
use pfet_03v3_ANSKCD  M4
timestamp 0
transform 1 0 1455 0 1 384
box -225 -204 225 204
use nfet_03v3_V3AFXU  M5
timestamp 0
transform 1 0 1875 0 1 3988
box -225 -3838 225 3838
use pfet_03v3_5MBUKS  M6
timestamp 0
transform 1 0 2295 0 1 3958
box -225 -3838 225 3838
use nfet_03v3_QVDB54  M7
timestamp 0
transform 1 0 2715 0 1 452
box -225 -362 225 362
use pfet_03v3_ANSKZB  M8
timestamp 0
transform 1 0 3135 0 1 422
box -225 -362 225 362
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 640 0 0 0 VA
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 640 0 0 0 VB
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 640 0 0 0 VG_N
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 640 0 0 0 VG_P
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 640 0 0 0 IB_N
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 640 0 0 0 IB_P
port 5 nsew
flabel metal1 0 -1200 100 -1100 0 FreeSans 640 0 0 0 VDD
port 6 nsew
flabel metal1 0 -1400 100 -1300 0 FreeSans 640 0 0 0 VSS
port 7 nsew
flabel metal1 0 -1600 100 -1500 0 FreeSans 640 0 0 0 VC
port 8 nsew
<< end >>
