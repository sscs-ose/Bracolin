* NGSPICE file created from DiffN_net.ext - technology: gf180mcuD

.subckt DiffN_net VSS VDD VN IT OUT VP
X0 VDD.t71 VDD.t70 VDD.t71 VDD.t7 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X1 VDD.t69 VDD.t68 VDD.t69 VDD.t4 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X2 a_438_9747# a_n92_682.t12 OUT.t1 VDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X3 a_1844_8581# a_n92_682.t13 VDD.t75 VDD.t41 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X4 a_438_7815# a_n92_682.t14 OUT.t3 VDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X5 OUT a_n92_682.t15 a_1844_6649# VDD.t46 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X6 VDD.t67 VDD.t66 VDD.t67 VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X7 OUT VN.t0 a_1834_682# VSS.t2 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X8 VSS.t71 VSS.t70 VSS.t71 VSS.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X9 a_1834_682# VN.t1 IT.t2 VSS.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X10 a_438_6649# a_n92_682.t4 a_n92_682.t5 VDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X11 VDD.t65 VDD.t64 VDD.t65 VDD.t41 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X12 VSS.t69 VSS.t68 VSS.t69 VSS.t15 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X13 VSS.t67 VSS.t66 VSS.t67 VSS.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X14 VSS.t65 VSS.t64 VSS.t65 VSS.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X15 VDD.t63 VDD.t62 VDD.t63 VDD.t46 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X16 VSS.t63 VSS.t62 VSS.t63 VSS.t8 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X17 VSS.t61 VSS.t60 VSS.t61 VSS.t15 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X18 VSS.t59 VSS.t58 VSS.t59 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X19 VSS.t57 VSS.t56 VSS.t57 VSS.t15 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X20 VSS.t55 VSS.t54 VSS.t55 VSS.t8 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X21 VSS.t53 VSS.t52 VSS.t53 VSS.t8 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X22 VSS.t51 VSS.t50 VSS.t51 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X23 VDD a_n92_682.t16 a_438_9747# VDD.t15 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X24 VDD.t61 VDD.t60 VDD.t61 VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X25 VDD a_n92_682.t17 a_438_7815# VDD.t15 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X26 VDD.t59 VDD.t58 VDD.t59 VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X27 VDD.t57 VDD.t56 VDD.t57 VDD.t7 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X28 VDD.t55 VDD.t54 VDD.t55 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X29 OUT a_n92_682.t18 a_1844_8581# VDD.t46 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X30 VDD.t53 VDD.t52 VDD.t53 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X31 VDD.t51 VDD.t50 VDD.t51 VDD.t36 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X32 VSS.t49 VSS.t48 VSS.t49 VSS.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X33 a_1834_2606# VN.t2 IT.t3 VSS.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X34 OUT VN.t3 a_1834_2606# VSS.t2 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X35 a_438_8581# a_n92_682.t8 a_n92_682.t9 VDD.t36 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X36 VDD a_n92_682.t19 a_438_6649# VDD.t15 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X37 VDD.t49 VDD.t48 VDD.t49 VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X38 VDD.t47 VDD.t45 VDD.t47 VDD.t46 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X39 VSS.t47 VSS.t46 VSS.t47 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X40 VSS.t45 VSS.t44 VSS.t45 VSS.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X41 VDD.t44 VDD.t43 VDD.t44 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X42 IT VP.t0 a_430_682# VSS.t1 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X43 VDD.t42 VDD.t40 VDD.t42 VDD.t41 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X44 VDD.t39 VDD.t38 VDD.t39 VDD.t4 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X45 VDD.t37 VDD.t35 VDD.t37 VDD.t36 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X46 a_1834_3764# VP.t1 IT.t6 VSS.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X47 a_430_2606# VP.t3 a_n92_682.t1 VSS.t0 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X48 VSS.t43 VSS.t42 VSS.t43 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X49 VDD.t34 VDD.t33 VDD.t34 VDD.t7 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X50 VDD.t32 VDD.t31 VDD.t32 VDD.t7 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X51 VDD.t30 VDD.t29 VDD.t30 VDD.t4 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X52 VSS.t41 VSS.t40 VSS.t41 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X53 a_1834_1840# VP.t5 IT.t5 VSS.t3 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X54 VSS.t39 VSS.t38 VSS.t39 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X55 VDD.t28 VDD.t27 VDD.t28 VDD.t4 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X56 VDD.t26 VDD.t25 VDD.t26 VDD.t4 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X57 VDD.t24 VDD.t23 VDD.t24 VDD.t7 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X58 a_430_3764# VN.t4 OUT.t5 VSS.t0 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X59 a_1844_9747# a_n92_682.t20 VDD.t74 VDD.t41 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X60 a_1844_7815# a_n92_682.t21 VDD.t80 VDD.t41 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X61 a_430_1840# VN.t5 OUT.t0 VSS.t0 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X62 VDD a_n92_682.t22 a_438_8581# VDD.t15 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X63 VDD.t22 VDD.t21 VDD.t22 VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X64 VSS.t37 VSS.t36 VSS.t37 VSS.t15 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X65 VDD.t20 VDD.t19 VDD.t20 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X66 a_1844_6649# a_n92_682.t23 VDD.t83 VDD.t41 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X67 VSS.t35 VSS.t34 VSS.t35 VSS.t2 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X68 VDD.t18 VDD.t17 VDD.t18 VDD.t15 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X69 VDD.t16 VDD.t14 VDD.t16 VDD.t15 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X70 VDD.t13 VDD.t11 VDD.t13 VDD.t12 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X71 VSS.t33 VSS.t32 VSS.t33 VSS.t3 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X72 VSS.t31 VSS.t30 VSS.t31 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X73 VSS.t29 VSS.t28 VSS.t29 VSS.t8 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X74 VSS.t27 VSS.t26 VSS.t27 VSS.t2 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X75 VDD.t10 VDD.t9 VDD.t10 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X76 IT VP.t6 a_430_2606# VSS.t1 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X77 VSS.t25 VSS.t24 VSS.t25 VSS.t3 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X78 VSS.t23 VSS.t21 VSS.t23 VSS.t22 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X79 a_430_682# VP.t7 a_n92_682.t0 VSS.t0 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X80 VSS.t20 VSS.t19 VSS.t20 VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X81 VSS.t18 VSS.t17 VSS.t18 VSS.t15 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X82 VSS.t16 VSS.t14 VSS.t16 VSS.t15 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X83 VDD.t8 VDD.t6 VDD.t8 VDD.t7 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X84 VDD.t5 VDD.t3 VDD.t5 VDD.t4 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X85 VSS.t13 VSS.t12 VSS.t13 VSS.t8 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X86 VSS.t11 VSS.t10 VSS.t11 VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X87 IT VN.t6 a_430_3764# VSS.t1 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X88 VSS.t9 VSS.t7 VSS.t9 VSS.t8 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X89 VDD.t2 VDD.t0 VDD.t2 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X90 VSS.t6 VSS.t4 VSS.t6 VSS.t5 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X91 IT VN.t7 a_430_1840# VSS.t1 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
R0 VDD.n79 VDD.n5 477.971
R1 VDD.n76 VDD.n6 470.842
R2 VDD.n79 VDD.n6 470.842
R3 VDD.n76 VDD.n5 469.683
R4 VDD.t46 VDD.t12 142.93
R5 VDD.t36 VDD.t4 142.93
R6 VDD.t12 VDD.t1 96.8792
R7 VDD.t41 VDD.t46 96.8792
R8 VDD.t15 VDD.t36 96.8792
R9 VDD.t4 VDD.t7 96.8792
R10 VDD.t1 VDD.n5 81.1238
R11 VDD.t7 VDD.n6 81.1238
R12 VDD.n77 VDD.t41 70.2717
R13 VDD.n78 VDD.t15 64.1315
R14 VDD.n78 VDD.n77 8.52856
R15 VDD.n18 VDD.t66 8.10567
R16 VDD.n18 VDD.t0 8.10567
R17 VDD.n16 VDD.t60 8.10567
R18 VDD.n16 VDD.t54 8.10567
R19 VDD.n15 VDD.t21 8.10567
R20 VDD.n15 VDD.t19 8.10567
R21 VDD.n0 VDD.t58 8.10567
R22 VDD.n0 VDD.t52 8.10567
R23 VDD.n89 VDD.t48 8.10567
R24 VDD.n89 VDD.t43 8.10567
R25 VDD.n87 VDD.t11 8.10567
R26 VDD.n87 VDD.t9 8.10567
R27 VDD.n71 VDD.t50 8.10567
R28 VDD.n25 VDD.t17 8.10567
R29 VDD.n7 VDD.t40 8.10567
R30 VDD.n21 VDD.t62 8.10567
R31 VDD.n48 VDD.t56 8.10567
R32 VDD.n48 VDD.t27 8.10567
R33 VDD.n46 VDD.t33 8.10567
R34 VDD.n46 VDD.t38 8.10567
R35 VDD.n45 VDD.t6 8.10567
R36 VDD.n45 VDD.t3 8.10567
R37 VDD.n41 VDD.t31 8.10567
R38 VDD.n41 VDD.t29 8.10567
R39 VDD.n40 VDD.t23 8.10567
R40 VDD.n40 VDD.t25 8.10567
R41 VDD.n38 VDD.t70 8.10567
R42 VDD.n38 VDD.t68 8.10567
R43 VDD.n32 VDD.t35 8.10567
R44 VDD.n33 VDD.t14 8.10567
R45 VDD.n82 VDD.t64 8.10567
R46 VDD.n3 VDD.t45 8.10567
R47 VDD.n68 VDD.n67 4.61205
R48 VDD.n57 VDD.n56 4.61205
R49 VDD.n61 VDD.n59 4.5005
R50 VDD.n54 VDD.n52 4.5005
R51 VDD.n51 VDD.t83 4.00848
R52 VDD.n56 VDD.n55 4.00554
R53 VDD.n70 VDD.n69 3.87081
R54 VDD.n51 VDD.t80 3.78097
R55 VDD.n62 VDD.t74 3.78097
R56 VDD.n61 VDD.n60 3.77818
R57 VDD.n54 VDD.n53 3.77818
R58 VDD.n58 VDD.n57 3.61296
R59 VDD.n64 VDD.n58 3.34333
R60 VDD.n69 VDD.n68 3.26458
R61 VDD.n50 VDD.t51 3.20383
R62 VDD.n74 VDD.t18 3.20383
R63 VDD.n24 VDD.t42 3.20383
R64 VDD.n20 VDD.t63 3.20383
R65 VDD.n63 VDD.t75 3.20383
R66 VDD.n66 VDD.n65 3.20383
R67 VDD.n36 VDD.t37 3.20383
R68 VDD.t16 VDD.n4 3.20383
R69 VDD.n81 VDD.t65 3.20383
R70 VDD.n85 VDD.t47 3.20383
R71 VDD.n64 VDD.n63 3.1154
R72 VDD.n62 VDD.n59 2.65924
R73 VDD.n52 VDD.n51 2.65924
R74 VDD.n66 VDD.n64 2.61766
R75 VDD.n84 VDD.n83 1.73383
R76 VDD.n35 VDD.n34 1.73383
R77 VDD.n23 VDD.n22 1.73383
R78 VDD.n73 VDD.n72 1.73383
R79 VDD.t18 VDD.n73 1.4705
R80 VDD.n73 VDD.t51 1.4705
R81 VDD.n23 VDD.t63 1.4705
R82 VDD.t42 VDD.n23 1.4705
R83 VDD.n35 VDD.t16 1.4705
R84 VDD.t37 VDD.n35 1.4705
R85 VDD.t47 VDD.n84 1.4705
R86 VDD.n84 VDD.t65 1.4705
R87 VDD.n8 VDD.t2 1.00929
R88 VDD.n9 VDD.t55 1.00929
R89 VDD.n10 VDD.t20 1.00929
R90 VDD.n11 VDD.t53 1.00929
R91 VDD.n1 VDD.t44 1.00929
R92 VDD.n2 VDD.t10 1.00929
R93 VDD.n26 VDD.t28 1.00929
R94 VDD.n27 VDD.t39 1.00929
R95 VDD.n28 VDD.t5 1.00929
R96 VDD.n29 VDD.t30 1.00929
R97 VDD.n30 VDD.t26 1.00929
R98 VDD.n31 VDD.t69 1.00929
R99 VDD.n8 VDD.t67 1.00871
R100 VDD.n9 VDD.t61 1.00871
R101 VDD.n10 VDD.t22 1.00871
R102 VDD.n11 VDD.t59 1.00871
R103 VDD.n1 VDD.t49 1.00871
R104 VDD.n2 VDD.t13 1.00871
R105 VDD.n26 VDD.t57 1.00871
R106 VDD.n27 VDD.t34 1.00871
R107 VDD.n28 VDD.t8 1.00871
R108 VDD.n29 VDD.t32 1.00871
R109 VDD.n30 VDD.t24 1.00871
R110 VDD.n31 VDD.t71 1.00871
R111 VDD.n63 VDD.n62 0.805146
R112 VDD.n67 VDD.n66 0.80221
R113 VDD.n37 VDD.n31 0.468749
R114 VDD.n39 VDD.n30 0.468749
R115 VDD.n42 VDD.n29 0.468749
R116 VDD.n44 VDD.n28 0.468749
R117 VDD.n47 VDD.n27 0.468749
R118 VDD.n49 VDD.n26 0.468749
R119 VDD.n86 VDD.n2 0.468749
R120 VDD.n88 VDD.n1 0.468749
R121 VDD.n12 VDD.n11 0.468749
R122 VDD.n14 VDD.n10 0.468749
R123 VDD.n17 VDD.n9 0.468749
R124 VDD.n19 VDD.n8 0.468749
R125 VDD.n69 VDD.n58 0.3755
R126 VDD.n68 VDD.n59 0.157683
R127 VDD.n57 VDD.n52 0.157683
R128 VDD.n43 VDD.n6 0.10728
R129 VDD.n76 VDD.n75 0.10728
R130 VDD.n77 VDD.n76 0.10728
R131 VDD.n13 VDD.n5 0.10728
R132 VDD.n80 VDD.n79 0.1055
R133 VDD.n79 VDD.n78 0.1055
R134 VDD.n48 VDD.n47 0.0382419
R135 VDD.n39 VDD.n38 0.0382419
R136 VDD.n18 VDD.n17 0.0382419
R137 VDD.n88 VDD.n87 0.0382419
R138 VDD.n46 VDD.n45 0.0364748
R139 VDD.n41 VDD.n40 0.0364748
R140 VDD.n16 VDD.n15 0.0364748
R141 VDD.n21 VDD.n20 0.0346711
R142 VDD.n22 VDD.n21 0.0346711
R143 VDD.n22 VDD.n7 0.0346711
R144 VDD.n24 VDD.n7 0.0346711
R145 VDD.n74 VDD.n25 0.0346711
R146 VDD.n72 VDD.n25 0.0346711
R147 VDD.n72 VDD.n71 0.0346711
R148 VDD.n86 VDD.n85 0.0308563
R149 VDD.n37 VDD.n36 0.0308563
R150 VDD.n50 VDD.n49 0.0308128
R151 VDD.n20 VDD.n19 0.0308128
R152 VDD.n85 VDD.n3 0.0293162
R153 VDD.n83 VDD.n3 0.0293162
R154 VDD.n83 VDD.n82 0.0293162
R155 VDD.n82 VDD.n81 0.0293162
R156 VDD.n33 VDD.n4 0.0293162
R157 VDD.n34 VDD.n33 0.0293162
R158 VDD.n34 VDD.n32 0.0293162
R159 VDD.n36 VDD.n32 0.0293162
R160 VDD.n70 VDD.n50 0.0272991
R161 VDD.n44 VDD.n43 0.0270708
R162 VDD.n14 VDD.n13 0.0270708
R163 VDD.n43 VDD.n42 0.0222742
R164 VDD.n13 VDD.n12 0.0222742
R165 VDD.n49 VDD.n48 0.0193079
R166 VDD.n47 VDD.n46 0.0193079
R167 VDD.n45 VDD.n44 0.0193079
R168 VDD.n42 VDD.n41 0.0193079
R169 VDD.n40 VDD.n39 0.0193079
R170 VDD.n38 VDD.n37 0.0193079
R171 VDD.n19 VDD.n18 0.0193079
R172 VDD.n17 VDD.n16 0.0193079
R173 VDD.n15 VDD.n14 0.0193079
R174 VDD.n12 VDD.n0 0.0193079
R175 VDD.n89 VDD.n88 0.0193079
R176 VDD.n87 VDD.n86 0.0193079
R177 VDD VDD.n0 0.0188661
R178 VDD.n81 VDD.n80 0.0185609
R179 VDD VDD.n89 0.0181087
R180 VDD.n75 VDD.n74 0.0175856
R181 VDD.n75 VDD.n24 0.0159011
R182 VDD.n71 VDD.n70 0.0108166
R183 VDD.n80 VDD.n4 0.00983484
R184 VDD.n67 VDD.n61 0.00523684
R185 VDD.n56 VDD.n54 0.00523684
R186 a_n92_682.t1 a_n92_682.t9 12.6502
R187 a_n92_682.t1 a_n92_682.t6 10.2828
R188 a_n92_682.t1 a_n92_682.t10 10.2828
R189 a_n92_682.t1 a_n92_682.t18 10.2828
R190 a_n92_682.t1 a_n92_682.t15 10.2828
R191 a_n92_682.t1 a_n92_682.t12 10.1333
R192 a_n92_682.t1 a_n92_682.t14 10.1333
R193 a_n92_682.t1 a_n92_682.t8 10.1333
R194 a_n92_682.t1 a_n92_682.t4 10.1333
R195 a_n92_682.t1 a_n92_682.t0 9.7247
R196 a_n92_682.t1 a_n92_682.t23 9.57156
R197 a_n92_682.t1 a_n92_682.t20 9.57156
R198 a_n92_682.t1 a_n92_682.t21 9.57156
R199 a_n92_682.t1 a_n92_682.t13 9.57156
R200 a_n92_682.t1 a_n92_682.t19 9.57156
R201 a_n92_682.t1 a_n92_682.t16 9.57156
R202 a_n92_682.t1 a_n92_682.t17 9.57156
R203 a_n92_682.t1 a_n92_682.t22 9.57156
R204 a_n92_682.t1 a_n92_682.n2 8.03774
R205 a_n92_682.t0 a_n92_682.n1 8.03774
R206 a_n92_682.t1 a_n92_682.n0 7.97167
R207 a_n92_682.t1 a_n92_682.n3 7.97167
R208 a_n92_682.t5 a_n92_682.t1 7.35438
R209 OUT.n3 OUT.t1 10.6384
R210 OUT.n6 OUT.t5 10.1588
R211 OUT.n5 OUT.n4 9.34003
R212 OUT.n8 OUT.t0 7.9312
R213 OUT.n2 OUT.t3 7.66186
R214 OUT.n2 OUT.n1 7.2428
R215 OUT.n8 OUT.n7 7.23802
R216 OUT OUT.n9 6.76897
R217 OUT OUT.n0 3.63761
R218 OUT.n9 OUT.n8 2.2505
R219 OUT.n3 OUT.n2 2.2505
R220 OUT.n6 OUT.n5 0.79175
R221 OUT.n9 OUT.n6 0.726875
R222 OUT.n5 OUT.n3 0.67625
R223 VN.n1 VN.t1 8.41259
R224 VN.n4 VN.t2 8.41259
R225 VN.n1 VN.t0 8.3889
R226 VN.n4 VN.t3 8.3889
R227 VN.n21 VN.t5 8.06917
R228 VN.n16 VN.t7 8.06917
R229 VN.n6 VN.t6 8.06917
R230 VN.n5 VN.t4 8.06917
R231 VN.n16 VN.n0 4.64616
R232 VN.n7 VN.n6 4.64616
R233 VN.n19 VN.n15 4.64379
R234 VN.n10 VN.n3 4.64379
R235 VN.n9 VN.n8 4.5005
R236 VN.n18 VN.n17 4.5005
R237 VN.n13 VN.n3 3.48816
R238 VN.n15 VN.n14 3.43191
R239 VN.n2 VN.n1 2.78312
R240 VN.n12 VN.n4 2.78312
R241 VN.n20 VN.n19 2.35902
R242 VN.n11 VN.n10 2.35902
R243 VN.n14 VN.n2 2.30675
R244 VN.n21 VN.n20 2.28769
R245 VN.n11 VN.n5 2.28769
R246 VN.n13 VN.n12 2.2505
R247 VN.n7 VN.n5 2.01635
R248 VN.n22 VN.n0 1.96437
R249 VN.n20 VN.n2 1.34566
R250 VN.n12 VN.n11 1.34566
R251 VN.n14 VN.n13 0.666125
R252 VN.n8 VN.n3 0.157683
R253 VN.n8 VN.n7 0.157683
R254 VN.n17 VN.n15 0.157683
R255 VN.n17 VN.n0 0.157683
R256 VN VN.n22 0.137512
R257 VN.n22 VN.n21 0.0521211
R258 VN.n19 VN.n18 0.00405263
R259 VN.n10 VN.n9 0.00405263
R260 VN.n18 VN.n16 0.00168421
R261 VN.n9 VN.n6 0.00168421
R262 VSS.n58 VSS.n6 523.342
R263 VSS.n61 VSS.n5 521.869
R264 VSS.n58 VSS.n5 519.659
R265 VSS.n61 VSS.n6 516.342
R266 VSS.t2 VSS.t22 442.449
R267 VSS.t0 VSS.t5 442.449
R268 VSS.t22 VSS.t15 301.425
R269 VSS.t3 VSS.t2 301.425
R270 VSS.t1 VSS.t0 301.425
R271 VSS.t5 VSS.t8 301.425
R272 VSS.t15 VSS.n5 251.454
R273 VSS.t8 VSS.n6 251.454
R274 VSS.n59 VSS.t3 216.381
R275 VSS.n60 VSS.t1 210.998
R276 VSS.n60 VSS.n59 26.9134
R277 VSS.n20 VSS.t30 8.06917
R278 VSS.n20 VSS.t68 8.06917
R279 VSS.n18 VSS.t40 8.06917
R280 VSS.n18 VSS.t17 8.06917
R281 VSS.n17 VSS.t46 8.06917
R282 VSS.n17 VSS.t36 8.06917
R283 VSS.n13 VSS.t38 8.06917
R284 VSS.n13 VSS.t14 8.06917
R285 VSS.n12 VSS.t42 8.06917
R286 VSS.n12 VSS.t56 8.06917
R287 VSS.n69 VSS.t21 8.06917
R288 VSS.n69 VSS.t60 8.06917
R289 VSS.n53 VSS.t19 8.06917
R290 VSS.n27 VSS.t58 8.06917
R291 VSS.n7 VSS.t32 8.06917
R292 VSS.n23 VSS.t34 8.06917
R293 VSS.n50 VSS.t62 8.06917
R294 VSS.n50 VSS.t48 8.06917
R295 VSS.n48 VSS.t12 8.06917
R296 VSS.n48 VSS.t66 8.06917
R297 VSS.n47 VSS.t28 8.06917
R298 VSS.n47 VSS.t4 8.06917
R299 VSS.n43 VSS.t7 8.06917
R300 VSS.n43 VSS.t64 8.06917
R301 VSS.n42 VSS.t52 8.06917
R302 VSS.n42 VSS.t70 8.06917
R303 VSS.n40 VSS.t54 8.06917
R304 VSS.n40 VSS.t44 8.06917
R305 VSS.n34 VSS.t10 8.06917
R306 VSS.n35 VSS.t50 8.06917
R307 VSS.n64 VSS.t24 8.06917
R308 VSS.n3 VSS.t26 8.06917
R309 VSS.n52 VSS.t20 3.3605
R310 VSS.n56 VSS.t59 3.3605
R311 VSS.n26 VSS.t33 3.3605
R312 VSS.n22 VSS.t35 3.3605
R313 VSS.n38 VSS.t11 3.3605
R314 VSS.t51 VSS.n4 3.3605
R315 VSS.n63 VSS.t25 3.3605
R316 VSS.n67 VSS.t27 3.3605
R317 VSS.n66 VSS.n65 2.1005
R318 VSS.n37 VSS.n36 2.1005
R319 VSS.n25 VSS.n24 2.1005
R320 VSS.n55 VSS.n54 2.1005
R321 VSS.t59 VSS.n55 1.2605
R322 VSS.n55 VSS.t20 1.2605
R323 VSS.n25 VSS.t35 1.2605
R324 VSS.t33 VSS.n25 1.2605
R325 VSS.n37 VSS.t51 1.2605
R326 VSS.t11 VSS.n37 1.2605
R327 VSS.t27 VSS.n66 1.2605
R328 VSS.n66 VSS.t25 1.2605
R329 VSS.n8 VSS.t69 0.918039
R330 VSS.n9 VSS.t18 0.918039
R331 VSS.n10 VSS.t37 0.918039
R332 VSS.n11 VSS.t16 0.918039
R333 VSS.n0 VSS.t57 0.918039
R334 VSS.n2 VSS.t61 0.918039
R335 VSS.n28 VSS.t49 0.918039
R336 VSS.n29 VSS.t67 0.918039
R337 VSS.n30 VSS.t6 0.918039
R338 VSS.n31 VSS.t65 0.918039
R339 VSS.n32 VSS.t71 0.918039
R340 VSS.n33 VSS.t45 0.918039
R341 VSS.n8 VSS.t31 0.91749
R342 VSS.n9 VSS.t41 0.91749
R343 VSS.n10 VSS.t47 0.91749
R344 VSS.n11 VSS.t39 0.91749
R345 VSS.n0 VSS.t43 0.91749
R346 VSS.n2 VSS.t23 0.91749
R347 VSS.n28 VSS.t63 0.91749
R348 VSS.n29 VSS.t13 0.91749
R349 VSS.n30 VSS.t29 0.91749
R350 VSS.n31 VSS.t9 0.91749
R351 VSS.n32 VSS.t53 0.91749
R352 VSS.n33 VSS.t55 0.91749
R353 VSS.n39 VSS.n33 0.582999
R354 VSS.n41 VSS.n32 0.582999
R355 VSS.n44 VSS.n31 0.582999
R356 VSS.n46 VSS.n30 0.582999
R357 VSS.n49 VSS.n29 0.582999
R358 VSS.n51 VSS.n28 0.582999
R359 VSS.n68 VSS.n2 0.582999
R360 VSS.n1 VSS.n0 0.582999
R361 VSS.n14 VSS.n11 0.582999
R362 VSS.n16 VSS.n10 0.582999
R363 VSS.n19 VSS.n9 0.582999
R364 VSS.n21 VSS.n8 0.582999
R365 VSS.n45 VSS.n6 0.0886356
R366 VSS.n58 VSS.n57 0.0886356
R367 VSS.n59 VSS.n58 0.0886356
R368 VSS.n15 VSS.n5 0.0886356
R369 VSS.n62 VSS.n61 0.0871667
R370 VSS.n61 VSS.n60 0.0871667
R371 VSS.n50 VSS.n49 0.0390622
R372 VSS.n41 VSS.n40 0.0390622
R373 VSS.n20 VSS.n19 0.0385696
R374 VSS.n48 VSS.n47 0.0371211
R375 VSS.n43 VSS.n42 0.0371211
R376 VSS.n18 VSS.n17 0.0366533
R377 VSS.n13 VSS.n12 0.0366533
R378 VSS.n23 VSS.n22 0.0341
R379 VSS.n24 VSS.n23 0.0341
R380 VSS.n24 VSS.n7 0.0341
R381 VSS.n26 VSS.n7 0.0341
R382 VSS.n56 VSS.n27 0.0341
R383 VSS.n54 VSS.n27 0.0341
R384 VSS.n54 VSS.n53 0.0341
R385 VSS.n53 VSS.n52 0.0341
R386 VSS.n39 VSS.n38 0.0302339
R387 VSS.n46 VSS.n45 0.0301981
R388 VSS.n68 VSS.n67 0.0301505
R389 VSS.n52 VSS.n51 0.0300328
R390 VSS.n22 VSS.n21 0.0299989
R391 VSS.n16 VSS.n15 0.0298187
R392 VSS VSS.n1 0.0297548
R393 VSS.n67 VSS.n3 0.0294988
R394 VSS.n65 VSS.n3 0.0294988
R395 VSS.n65 VSS.n64 0.0294988
R396 VSS.n64 VSS.n63 0.0294988
R397 VSS.n35 VSS.n4 0.0294988
R398 VSS.n36 VSS.n35 0.0294988
R399 VSS.n36 VSS.n34 0.0294988
R400 VSS.n38 VSS.n34 0.0294988
R401 VSS.n45 VSS.n44 0.0203634
R402 VSS.n15 VSS.n14 0.0201097
R403 VSS.n57 VSS.n56 0.01994
R404 VSS.n51 VSS.n50 0.0196517
R405 VSS.n49 VSS.n48 0.0196517
R406 VSS.n47 VSS.n46 0.0196517
R407 VSS.n44 VSS.n43 0.0196517
R408 VSS.n42 VSS.n41 0.0196517
R409 VSS.n40 VSS.n39 0.0196517
R410 VSS.n21 VSS.n20 0.019407
R411 VSS.n19 VSS.n18 0.019407
R412 VSS.n17 VSS.n16 0.019407
R413 VSS.n14 VSS.n13 0.019407
R414 VSS.n12 VSS.n1 0.019407
R415 VSS.n69 VSS.n68 0.019407
R416 VSS.n63 VSS.n62 0.0183136
R417 VSS.n57 VSS.n26 0.01514
R418 VSS.n62 VSS.n4 0.0120995
R419 VSS VSS.n69 0.00931476
R420 IT.n9 IT.t2 6.55856
R421 IT.n2 IT.t6 6.51441
R422 IT.n2 IT.n1 5.98782
R423 IT.n8 IT.n2 4.04004
R424 IT.n9 IT.n8 3.979
R425 IT.n6 IT.n4 3.89695
R426 IT.n3 IT.t3 3.89695
R427 IT.n6 IT.n5 3.73116
R428 IT.n3 IT.t5 3.73116
R429 IT IT.n0 3.55589
R430 IT.n8 IT.n7 3.39813
R431 IT.n7 IT.n3 2.58466
R432 IT IT.n9 2.44554
R433 IT.n7 IT.n6 2.22759
R434 VP.n5 VP.t2 11.4656
R435 VP.n1 VP.t4 11.4656
R436 VP.n5 VP.t1 10.736
R437 VP.n1 VP.t5 10.736
R438 VP.n17 VP.t0 8.06917
R439 VP.n9 VP.t6 8.06917
R440 VP.n8 VP.t3 8.06917
R441 VP.n15 VP.t7 8.06917
R442 VP VP.n0 4.73347
R443 VP.n10 VP.n9 4.64616
R444 VP.n17 VP.n16 4.64616
R445 VP.n18 VP.n0 4.5005
R446 VP.n11 VP.n7 2.43517
R447 VP.n7 VP.n6 2.38451
R448 VP.n19 VP.n2 2.38035
R449 VP.n12 VP.n4 2.31238
R450 VP.n13 VP.n3 2.31238
R451 VP.n12 VP.n11 2.2505
R452 VP.n14 VP.n13 2.2505
R453 VP.n8 VP.n4 2.20398
R454 VP.n15 VP.n14 2.20398
R455 VP.n10 VP.n8 2.01137
R456 VP.n16 VP.n15 2.01137
R457 VP.n6 VP.n5 1.05605
R458 VP.n2 VP.n1 1.05605
R459 VP.n13 VP.n12 0.65975
R460 VP.n6 VP.n4 0.118858
R461 VP.n14 VP.n2 0.118858
R462 VP.n3 VP.n0 0.114585
R463 VP VP.n19 0.0644474
R464 VP.n11 VP.n10 0.0435986
R465 VP.n16 VP.n3 0.0435986
R466 VP.n19 VP.n18 0.00760526
R467 VP.n9 VP.n7 0.00562075
R468 VP.n18 VP.n17 0.00168421
C0 VN VP 3.20803f
C1 VDD a_438_6649# 0.071285f
C2 OUT a_430_1840# 0.029214f
C3 a_430_1840# VP 0.018108f
C4 IT a_430_682# 0.055103f
C5 OUT a_438_7815# 0.042859f
C6 IT a_430_2606# 0.042833f
C7 VDD a_438_9747# 0.071615f
C8 VN a_1834_3764# 0.063013f
C9 VN a_1834_682# 0.146345f
C10 VDD a_1844_9747# 0.05845f
C11 OUT a_1844_6649# 0.05266f
C12 a_430_682# VP 0.111688f
C13 IT a_1834_1840# 0.042422f
C14 VN a_430_1840# 0.094098f
C15 VDD a_438_7815# 0.060056f
C16 OUT a_430_2606# 0.013188f
C17 a_430_2606# VP 0.111688f
C18 VDD a_1844_6649# 0.05812f
C19 IT a_430_3764# 0.055502f
C20 a_1834_1840# VP 0.078551f
C21 OUT a_1844_7815# 0.024944f
C22 IT a_1834_2606# 0.029143f
C23 VDD a_438_8581# 0.074277f
C24 OUT a_430_3764# 0.029162f
C25 a_430_3764# VP 0.018108f
C26 OUT IT 4.3178f
C27 IT VP 2.22362f
C28 VN a_1834_1840# 0.064867f
C29 VDD a_1844_7815# 0.046892f
C30 OUT a_1834_2606# 0.044666f
C31 a_1834_2606# VP 0.01303f
C32 OUT a_1844_8581# 0.039403f
C33 IT a_1834_3764# 0.041812f
C34 IT a_1834_682# 0.041413f
C35 OUT VP 0.902686f
C36 VN a_430_3764# 0.094098f
C37 OUT a_438_6649# 0.013996f
C38 VN IT 1.6819f
C39 IT a_430_1840# 0.056112f
C40 VN a_1834_2606# 0.148004f
C41 VDD a_1844_8581# 0.061113f
C42 OUT a_1834_682# 0.032229f
C43 a_1834_3764# VP 0.078551f
C44 a_1834_682# VP 0.01303f
C45 OUT VDD 4.54076f
C46 OUT a_438_9747# 0.042379f
C47 OUT a_1844_9747# 0.024463f
C48 VN OUT 2.05197f
.ends

