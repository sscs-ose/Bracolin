* Extracted by KLayout with GF180MCU LVS runset on : 29/04/2024 18:36

.SUBCKT SAR_Asynchronous_top_neg_logic vocp D Valid VSSD Bit_10 Bit_10_n Bit_9
+ Bit_9_n Bit_8 Bit_8_n Bit_7 Bit_7_n Bit_6 Bit_5 Bit_4 Bit_3 Bit_2 Bit_2_n
+ Bit_1 Bit_1_n VDDD Set CK_1 clks Reset VCM
M$1 \$9 \$707 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$2 \$59 \$9 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$3 \$22 \$21 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$4 \$10 \$713 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$5 \$60 \$10 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$6 \$26 \$25 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$7 \$11 \$719 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$8 \$61 \$11 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$9 \$30 \$29 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$10 \$12 \$725 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$11 \$62 \$12 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$12 \$34 \$33 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$13 \$13 \$731 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$14 \$63 \$13 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$15 \$38 \$37 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$16 \$14 \$737 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$17 \$64 \$14 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$18 \$42 \$41 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$19 \$15 \$743 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$20 \$65 \$15 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$21 \$46 \$45 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$22 \$16 \$749 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$23 \$66 \$16 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$24 \$50 \$49 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$25 \$17 \$755 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$26 \$67 \$17 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$27 \$54 \$53 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$28 \$18 \$761 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$29 \$68 \$18 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$30 \$58 \$57 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$31 Bit_10_n \$59 Bit_10 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$32 \$21 \$9 Bit_10 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$33 Bit_10_n \$9 \$22 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$34 Bit_9_n \$60 Bit_9 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$35 \$25 \$10 Bit_9 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$36 Bit_9_n \$10 \$26 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$37 Bit_8_n \$61 Bit_8 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$38 \$29 \$11 Bit_8 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$39 Bit_8_n \$11 \$30 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$40 Bit_7_n \$62 Bit_7 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$41 \$33 \$12 Bit_7 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$42 Bit_7_n \$12 \$34 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$43 \$36 \$63 Bit_6 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$44 \$37 \$13 Bit_6 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$45 \$36 \$13 \$38 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$46 \$40 \$64 Bit_5 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$47 \$41 \$14 Bit_5 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$48 \$40 \$14 \$42 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$49 \$44 \$65 Bit_4 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$50 \$45 \$15 Bit_4 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$51 \$44 \$15 \$46 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$52 \$48 \$66 Bit_3 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$53 \$49 \$16 Bit_3 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$54 \$48 \$16 \$50 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$55 Bit_2_n \$67 Bit_2 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$56 \$53 \$17 Bit_2 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$57 Bit_2_n \$17 \$54 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$58 Bit_1_n \$68 Bit_1 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$59 \$57 \$18 Bit_1 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$60 Bit_1_n \$18 \$58 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$61 \$768 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$62 \$769 \$768 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$63 \$702 \$769 D VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$64 \$1587 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$65 \$703 \$702 \$1587 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$66 \$1588 \$703 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$67 \$704 clks \$1588 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$68 \$702 \$768 \$704 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$69 \$706 \$768 \$703 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$70 \$1589 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$71 \$707 \$706 \$1589 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$72 \$1590 \$707 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$73 \$705 Set \$1590 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$74 \$706 \$769 \$705 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$75 \$770 \$707 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$76 \$771 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$77 \$772 \$771 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$78 \$708 \$772 \$707 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$79 \$1591 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$80 \$709 \$708 \$1591 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$81 \$1592 \$709 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$82 \$710 clks \$1592 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$83 \$708 \$771 \$710 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$84 \$712 \$771 \$709 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$85 \$1593 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$86 \$713 \$712 \$1593 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$87 \$1594 \$713 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$88 \$711 Set \$1594 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$89 \$712 \$772 \$711 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$90 \$773 \$713 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$91 \$774 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$92 \$775 \$774 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$93 \$714 \$775 \$713 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$94 \$1595 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$95 \$715 \$714 \$1595 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$96 \$1596 \$715 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$97 \$716 clks \$1596 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$98 \$714 \$774 \$716 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$99 \$718 \$774 \$715 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$100 \$1597 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$101 \$719 \$718 \$1597 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$102 \$1598 \$719 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$103 \$717 Set \$1598 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$104 \$718 \$775 \$717 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$105 \$776 \$719 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$106 \$777 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$107 \$778 \$777 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$108 \$720 \$778 \$719 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$109 \$1599 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$110 \$721 \$720 \$1599 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$111 \$1600 \$721 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$112 \$722 clks \$1600 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$113 \$720 \$777 \$722 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$114 \$724 \$777 \$721 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$115 \$1601 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$116 \$725 \$724 \$1601 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$117 \$1602 \$725 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$118 \$723 Set \$1602 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$119 \$724 \$778 \$723 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$120 \$779 \$725 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$121 \$780 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$122 \$781 \$780 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$123 \$726 \$781 \$725 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$124 \$1603 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$125 \$727 \$726 \$1603 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$126 \$1604 \$727 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$127 \$728 clks \$1604 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$128 \$726 \$780 \$728 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$129 \$730 \$780 \$727 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$130 \$1605 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$131 \$731 \$730 \$1605 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$132 \$1606 \$731 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$133 \$729 Set \$1606 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$134 \$730 \$781 \$729 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$135 \$782 \$731 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$136 \$783 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$137 \$784 \$783 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$138 \$732 \$784 \$731 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$139 \$1607 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$140 \$733 \$732 \$1607 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$141 \$1608 \$733 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$142 \$734 clks \$1608 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$143 \$732 \$783 \$734 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$144 \$736 \$783 \$733 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$145 \$1609 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$146 \$737 \$736 \$1609 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$147 \$1610 \$737 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$148 \$735 Set \$1610 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$149 \$736 \$784 \$735 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$150 \$785 \$737 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$151 \$786 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$152 \$787 \$786 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$153 \$738 \$787 \$737 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$154 \$1611 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$155 \$739 \$738 \$1611 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$156 \$1612 \$739 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$157 \$740 clks \$1612 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$158 \$738 \$786 \$740 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$159 \$742 \$786 \$739 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$160 \$1613 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$161 \$743 \$742 \$1613 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$162 \$1614 \$743 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$163 \$741 Set \$1614 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$164 \$742 \$787 \$741 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$165 \$788 \$743 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$166 \$789 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$167 \$790 \$789 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$168 \$744 \$790 \$743 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$169 \$1615 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$170 \$745 \$744 \$1615 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$171 \$1616 \$745 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$172 \$746 clks \$1616 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$173 \$744 \$789 \$746 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$174 \$748 \$789 \$745 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$175 \$1617 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$176 \$749 \$748 \$1617 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$177 \$1618 \$749 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$178 \$747 Set \$1618 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$179 \$748 \$790 \$747 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$180 \$791 \$749 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$181 \$792 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$182 \$793 \$792 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$183 \$750 \$793 \$749 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$184 \$1619 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$185 \$751 \$750 \$1619 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$186 \$1620 \$751 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$187 \$752 clks \$1620 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$188 \$750 \$792 \$752 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$189 \$754 \$792 \$751 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$190 \$1621 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$191 \$755 \$754 \$1621 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$192 \$1622 \$755 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$193 \$753 Set \$1622 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$194 \$754 \$793 \$753 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$195 \$794 \$755 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$196 \$795 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$197 \$796 \$795 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$198 \$756 \$796 \$755 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$199 \$1623 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$200 \$757 \$756 \$1623 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$201 \$1624 \$757 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$202 \$758 clks \$1624 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$203 \$756 \$795 \$758 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$204 \$760 \$795 \$757 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$205 \$1625 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$206 \$761 \$760 \$1625 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$207 \$1626 \$761 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$208 \$759 Set \$1626 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$209 \$760 \$796 \$759 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$210 \$797 \$761 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$211 \$798 Valid VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$212 \$799 \$798 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$213 \$762 \$799 \$761 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$214 \$1627 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$215 \$763 \$762 \$1627 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$216 \$1628 \$763 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$217 \$764 clks \$1628 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$218 \$762 \$798 \$764 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$219 \$767 \$798 \$763 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$220 \$1629 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$221 CK_1 \$767 \$1629 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$222 \$1630 CK_1 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$223 \$766 Set \$1630 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$224 \$767 \$799 \$766 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$225 \$800 CK_1 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$226 \$2211 \$2417 \$2215 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$227 VDDD \$2215 \$3049 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$228 \$2257 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$229 \$2258 \$2257 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$230 \$3032 \$3051 \$2987 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$231 \$3563 Set \$3032 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$232 \$2216 \$2258 \$2215 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$233 VDDD \$2215 \$3563 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$234 \$2632 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$235 \$2217 \$2216 \$2632 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$236 \$3564 \$2987 \$2215 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$237 VDDD Reset \$3564 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$238 \$2633 \$2217 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$239 \$2218 Reset \$2633 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$240 \$3033 \$3050 \$2987 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$241 \$2216 \$2257 \$2218 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$242 \$3034 \$3050 \$3022 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$243 \$2221 \$2257 \$2217 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$244 \$3565 Reset \$3034 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$245 VDDD \$3033 \$3565 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$246 \$2634 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$247 \$2219 \$2221 \$2634 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$248 \$3566 \$3022 \$3033 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$249 VDDD Set \$3566 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$250 \$2635 \$2219 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$251 vocp \$3051 \$3022 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$252 \$2220 Set \$2635 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$253 \$2221 \$2258 \$2220 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$254 VDDD \$3050 \$3051 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$255 VDDD \$2256 \$3050 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$256 \$2259 \$2219 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$257 VDDD \$2417 \$2256 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$258 VDDD CK_1 \$2417 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$259 \$2222 \$2431 \$2223 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$260 VDDD \$2223 \$3053 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$261 \$2261 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$262 \$2262 \$2261 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$263 \$3035 \$3055 \$2988 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$264 \$3567 Set \$3035 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$265 \$2224 \$2262 \$2223 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$266 VDDD \$2223 \$3567 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$267 \$2636 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$268 \$2225 \$2224 \$2636 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$269 \$3568 \$2988 \$2223 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$270 VDDD Reset \$3568 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$271 \$2637 \$2225 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$272 \$2226 Reset \$2637 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$273 \$3036 \$3054 \$2988 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$274 \$2224 \$2261 \$2226 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$275 \$3037 \$3054 \$3023 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$276 \$2229 \$2261 \$2225 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$277 \$3569 Reset \$3037 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$278 VDDD \$3036 \$3569 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$279 \$2638 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$280 \$2227 \$2229 \$2638 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$281 \$3570 \$3023 \$3036 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$282 VDDD Set \$3570 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$283 \$2639 \$2227 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$284 vocp \$3055 \$3023 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$285 \$2228 Set \$2639 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$286 \$2229 \$2262 \$2228 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$287 VDDD \$3054 \$3055 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$288 VDDD \$2260 \$3054 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$289 \$2263 \$2227 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$290 VDDD \$2431 \$2260 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$291 VDDD \$761 \$2431 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$292 \$2212 \$2444 \$2230 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$293 VDDD \$2230 \$3057 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$294 \$2265 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$295 \$2266 \$2265 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$296 \$3038 \$3059 \$2989 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$297 \$3571 Set \$3038 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$298 \$2231 \$2266 \$2230 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$299 VDDD \$2230 \$3571 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$300 \$2640 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$301 \$2232 \$2231 \$2640 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$302 \$3572 \$2989 \$2230 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$303 VDDD Reset \$3572 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$304 \$2641 \$2232 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$305 \$2233 Reset \$2641 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$306 \$3039 \$3058 \$2989 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$307 \$2231 \$2265 \$2233 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$308 \$3040 \$3058 \$3024 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$309 \$2236 \$2265 \$2232 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$310 \$3573 Reset \$3040 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$311 VDDD \$3039 \$3573 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$312 \$2642 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$313 \$2234 \$2236 \$2642 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$314 \$3574 \$3024 \$3039 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$315 VDDD Set \$3574 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$316 \$2643 \$2234 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$317 vocp \$3059 \$3024 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$318 \$2235 Set \$2643 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$319 \$2236 \$2266 \$2235 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$320 VDDD \$3058 \$3059 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$321 VDDD \$2264 \$3058 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$322 \$2267 \$2234 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$323 VDDD \$2444 \$2264 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$324 VDDD \$755 \$2444 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$325 \$2213 \$2457 \$2237 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$326 VDDD \$2237 \$3061 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$327 \$2269 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$328 \$2270 \$2269 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$329 \$3041 \$3063 \$2990 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$330 \$3575 Set \$3041 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$331 \$2238 \$2270 \$2237 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$332 VDDD \$2237 \$3575 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$333 \$2644 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$334 \$2239 \$2238 \$2644 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$335 \$3576 \$2990 \$2237 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$336 VDDD Reset \$3576 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$337 \$2645 \$2239 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$338 \$2240 Reset \$2645 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$339 \$3042 \$3062 \$2990 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$340 \$2238 \$2269 \$2240 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$341 \$3043 \$3062 \$3025 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$342 \$2243 \$2269 \$2239 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$343 \$3577 Reset \$3043 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$344 VDDD \$3042 \$3577 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$345 \$2646 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$346 \$2241 \$2243 \$2646 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$347 \$3578 \$3025 \$3042 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$348 VDDD Set \$3578 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$349 \$2647 \$2241 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$350 vocp \$3063 \$3025 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$351 \$2242 Set \$2647 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$352 \$2243 \$2270 \$2242 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$353 VDDD \$3062 \$3063 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$354 VDDD \$2268 \$3062 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$355 \$2271 \$2241 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$356 VDDD \$2457 \$2268 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$357 VDDD \$749 \$2457 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$358 \$2214 \$2470 \$2244 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$359 VDDD \$2244 \$3065 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$360 \$2273 clks VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$361 \$2274 \$2273 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$362 \$3044 \$3067 \$2991 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$363 \$3579 Set \$3044 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$364 \$2245 \$2274 \$2244 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$365 VDDD \$2244 \$3579 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$366 \$2648 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$367 \$2246 \$2245 \$2648 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$368 \$3580 \$2991 \$2244 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$369 VDDD Reset \$3580 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$370 \$2649 \$2246 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$371 \$2247 Reset \$2649 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$372 \$3045 \$3066 \$2991 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$373 \$2245 \$2273 \$2247 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$374 \$3046 \$3066 \$3026 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$375 \$2250 \$2273 \$2246 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$376 \$3581 Reset \$3046 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$377 VDDD \$3045 \$3581 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$378 \$2650 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$379 \$2248 \$2250 \$2650 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$380 \$3582 \$3026 \$3045 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$381 VDDD Set \$3582 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$382 \$2651 \$2248 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$383 vocp \$3067 \$3026 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$384 \$2249 Set \$2651 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$385 \$2250 \$2274 \$2249 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$386 VDDD \$3066 \$3067 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$387 VDDD \$2272 \$3066 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$388 \$2275 \$2248 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$389 VDDD \$2470 \$2272 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$390 VDDD \$743 \$2470 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$391 VDDD \$4016 \$4014 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$392 \$3983 \$4208 \$3938 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$393 \$4464 Set \$3983 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$394 VDDD \$4016 \$4464 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$395 \$4465 \$3938 \$4016 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$396 VDDD Reset \$4465 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$397 \$3984 \$4015 \$3938 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$398 \$3985 \$4015 \$3972 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$399 \$4466 Reset \$3985 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$400 VDDD \$3984 \$4466 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$401 \$4467 \$3972 \$3984 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$402 VDDD Set \$4467 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$403 \$3986 \$4208 \$3972 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$404 VDDD \$4015 \$4208 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$405 VDDD clks \$4015 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$406 \$3986 \$4017 \$3987 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$407 \$620 \$2256 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$408 VDDD \$3048 \$620 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$409 \$3048 \$2417 \$2215 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$410 VDDD \$4020 \$4018 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$411 VDDD \$2256 \$3048 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$412 \$3988 \$4230 \$3939 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$413 \$4468 Set \$3988 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$414 VDDD \$4020 \$4468 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$415 \$4469 \$3939 \$4020 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$416 VDDD Reset \$4469 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$417 \$3989 \$4019 \$3939 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$418 \$3990 \$4019 \$3973 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$419 \$4470 Reset \$3990 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$420 VDDD \$3989 \$4470 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$421 \$4471 \$3973 \$3989 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$422 VDDD Set \$4471 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$423 \$3991 \$4230 \$3973 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$424 VDDD \$4019 \$4230 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$425 VDDD clks \$4019 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$426 \$3991 \$4021 \$3974 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$427 Bit_1 \$2260 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$428 VDDD \$3052 Bit_1 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$429 \$3052 \$2431 \$2223 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$430 VDDD \$4024 \$4022 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$431 VDDD \$2260 \$3052 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$432 \$3992 \$4236 \$3940 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$433 \$4472 Set \$3992 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$434 VDDD \$4024 \$4472 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$435 \$4473 \$3940 \$4024 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$436 VDDD Reset \$4473 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$437 \$3993 \$4023 \$3940 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$438 \$3994 \$4023 \$3975 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$439 \$4474 Reset \$3994 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$440 VDDD \$3993 \$4474 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$441 \$4475 \$3975 \$3993 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$442 VDDD Set \$4475 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$443 \$3995 \$4236 \$3975 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$444 VDDD \$4023 \$4236 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$445 VDDD clks \$4023 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$446 \$3995 \$4025 \$3976 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$447 Bit_2 \$2264 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$448 VDDD \$3056 Bit_2 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$449 \$3056 \$2444 \$2230 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$450 VDDD \$4028 \$4026 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$451 VDDD \$2264 \$3056 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$452 \$3996 \$4258 \$3941 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$453 \$4476 Set \$3996 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$454 VDDD \$4028 \$4476 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$455 \$4477 \$3941 \$4028 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$456 VDDD Reset \$4477 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$457 \$3997 \$4027 \$3941 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$458 \$3998 \$4027 \$3977 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$459 \$4478 Reset \$3998 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$460 VDDD \$3997 \$4478 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$461 \$4479 \$3977 \$3997 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$462 VDDD Set \$4479 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$463 \$3999 \$4258 \$3977 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$464 VDDD \$4027 \$4258 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$465 VDDD clks \$4027 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$466 \$3999 \$4029 \$3978 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$467 Bit_3 \$2268 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$468 VDDD \$3060 Bit_3 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$469 \$3060 \$2457 \$2237 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$470 VDDD \$4032 \$4030 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$471 VDDD \$2268 \$3060 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$472 \$4000 \$4264 \$3942 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$473 \$4480 Set \$4000 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$474 VDDD \$4032 \$4480 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$475 \$4481 \$3942 \$4032 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$476 VDDD Reset \$4481 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$477 \$4001 \$4031 \$3942 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$478 \$4002 \$4031 \$3979 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$479 \$4482 Reset \$4002 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$480 VDDD \$4001 \$4482 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$481 \$4483 \$3979 \$4001 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$482 VDDD Set \$4483 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$483 \$4003 \$4264 \$3979 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$484 VDDD \$4031 \$4264 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$485 VDDD clks \$4031 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$486 \$4003 \$4033 \$3980 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$487 Bit_4 \$2272 VCM VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$488 VDDD \$3064 Bit_4 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$489 \$3064 \$2470 \$2244 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$490 VDDD \$4036 \$4034 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$491 VDDD \$2272 \$3064 VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$492 \$4004 \$4278 \$3943 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$493 \$4484 Set \$4004 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$494 VDDD \$4036 \$4484 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$495 \$4485 \$3943 \$4036 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$496 VDDD Reset \$4485 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$497 \$4005 \$4035 \$3943 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$498 \$4006 \$4035 \$3981 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$499 \$4486 Reset \$4006 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$500 VDDD \$4005 \$4486 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$501 \$4487 \$3981 \$4005 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$502 VDDD Set \$4487 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$503 \$4007 \$4278 \$3981 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$504 VDDD \$4035 \$4278 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$505 VDDD clks \$4035 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$506 \$4007 \$4037 \$3982 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$507 \$4017 \$707 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$508 \$4217 \$4017 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$509 \$4974 \$4217 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$510 \$5118 \$4974 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$511 \$4944 \$5118 vocp VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$512 \$5598 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$513 \$4945 \$4944 \$5598 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$514 \$5599 \$4945 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$515 \$4946 Reset \$5599 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$516 \$4944 \$4974 \$4946 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$517 \$4948 \$4974 \$4945 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$518 \$5600 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$519 \$3986 \$4948 \$5600 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$520 \$5601 \$3986 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$521 \$4947 Set \$5601 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$522 \$4948 \$5118 \$4947 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$523 \$4975 \$3986 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$524 \$4021 \$713 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$525 \$4231 \$4021 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$526 \$4977 \$4231 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$527 \$5119 \$4977 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$528 \$4949 \$5119 vocp VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$529 \$5602 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$530 \$4950 \$4949 \$5602 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$531 \$5603 \$4950 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$532 \$4951 Reset \$5603 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$533 \$4949 \$4977 \$4951 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$534 \$4953 \$4977 \$4950 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$535 \$5604 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$536 \$3991 \$4953 \$5604 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$537 \$5605 \$3991 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$538 \$4952 Set \$5605 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$539 \$4953 \$5119 \$4952 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$540 \$4978 \$3991 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$541 \$4025 \$719 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$542 \$4245 \$4025 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$543 \$4980 \$4245 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$544 \$5120 \$4980 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$545 \$4954 \$5120 vocp VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$546 \$5606 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$547 \$4955 \$4954 \$5606 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$548 \$5607 \$4955 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$549 \$4956 Reset \$5607 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$550 \$4954 \$4980 \$4956 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$551 \$4958 \$4980 \$4955 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$552 \$5608 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$553 \$3995 \$4958 \$5608 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$554 \$5609 \$3995 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$555 \$4957 Set \$5609 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$556 \$4958 \$5120 \$4957 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$557 \$4981 \$3995 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$558 \$4029 \$725 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$559 \$4259 \$4029 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$560 \$4983 \$4259 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$561 \$5121 \$4983 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$562 \$4959 \$5121 vocp VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$563 \$5610 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$564 \$4960 \$4959 \$5610 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$565 \$5611 \$4960 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$566 \$4961 Reset \$5611 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$567 \$4959 \$4983 \$4961 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$568 \$4963 \$4983 \$4960 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$569 \$5612 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$570 \$3999 \$4963 \$5612 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$571 \$5613 \$3999 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$572 \$4962 Set \$5613 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$573 \$4963 \$5121 \$4962 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$574 \$4984 \$3999 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$575 \$4033 \$731 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$576 \$4273 \$4033 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$577 \$4986 \$4273 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$578 \$5122 \$4986 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$579 \$4964 \$5122 vocp VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$580 \$5614 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$581 \$4965 \$4964 \$5614 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$582 \$5615 \$4965 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$583 \$4966 Reset \$5615 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$584 \$4964 \$4986 \$4966 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$585 \$4968 \$4986 \$4965 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$586 \$5616 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$587 \$4003 \$4968 \$5616 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$588 \$5617 \$4003 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$589 \$4967 Set \$5617 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$590 \$4968 \$5122 \$4967 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$591 \$4987 \$4003 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$592 \$4037 \$737 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$593 \$4287 \$4037 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$594 \$4989 \$4287 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$595 \$5123 \$4989 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$596 \$4969 \$5123 vocp VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$597 \$5618 Set VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P PS=9.1U
+ PD=9.1U
M$598 \$4970 \$4969 \$5618 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$599 \$5619 \$4970 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$600 \$4971 Reset \$5619 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$601 \$4969 \$4989 \$4971 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$602 \$4973 \$4989 \$4970 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$603 \$5620 Reset VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$604 \$4007 \$4973 \$5620 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$605 \$5621 \$4007 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$606 \$4972 Set \$5621 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$607 \$4973 \$5123 \$4972 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$608 \$4990 \$4007 VDDD VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$609 \$4976 \$4217 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$610 \$3986 \$4017 \$4976 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$611 Bit_10 \$4976 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$612 VCM \$4217 Bit_10 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$613 \$4979 \$4231 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$614 \$3991 \$4021 \$4979 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$615 Bit_9 \$4979 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$616 VCM \$4231 Bit_9 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$617 \$4982 \$4245 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$618 \$3995 \$4025 \$4982 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$619 Bit_8 \$4982 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$620 VCM \$4245 Bit_8 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$621 \$4985 \$4259 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$622 \$3999 \$4029 \$4985 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$623 Bit_7 \$4985 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$624 VCM \$4259 Bit_7 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$625 \$4988 \$4273 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$626 \$4003 \$4033 \$4988 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$627 Bit_6 \$4988 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$628 VCM \$4273 Bit_6 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$629 \$4991 \$4287 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$630 \$4007 \$4037 \$4991 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$631 Bit_5 \$4991 VDDD VDDD pfet_03v3 L=1.1U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$632 VCM \$4287 Bit_5 VDDD pfet_03v3 L=0.28U W=3.9U AS=2.535P AD=2.535P
+ PS=9.1U PD=9.1U
M$633 Bit_10_n \$9 Bit_10 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$634 \$21 \$59 Bit_10 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$635 Bit_10_n \$59 \$22 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$636 Bit_9_n \$10 Bit_9 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$637 \$25 \$60 Bit_9 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$638 Bit_9_n \$60 \$26 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$639 Bit_8_n \$11 Bit_8 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$640 \$29 \$61 Bit_8 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$641 Bit_8_n \$61 \$30 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$642 Bit_7_n \$12 Bit_7 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$643 \$33 \$62 Bit_7 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$644 Bit_7_n \$62 \$34 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$645 \$36 \$13 Bit_6 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$646 \$37 \$63 Bit_6 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$647 \$36 \$63 \$38 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$648 \$40 \$14 Bit_5 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$649 \$41 \$64 Bit_5 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$650 \$40 \$64 \$42 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$651 \$44 \$15 Bit_4 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$652 \$45 \$65 Bit_4 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$653 \$44 \$65 \$46 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$654 \$48 \$16 Bit_3 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$655 \$49 \$66 Bit_3 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$656 \$48 \$66 \$50 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$657 Bit_2_n \$17 Bit_2 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$658 \$53 \$67 Bit_2 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$659 Bit_2_n \$67 \$54 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$660 Bit_1_n \$18 Bit_1 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$661 \$57 \$68 Bit_1 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$662 Bit_1_n \$68 \$58 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$663 \$9 \$707 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$664 \$59 \$9 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$665 \$22 \$21 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$666 \$10 \$713 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$667 \$60 \$10 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$668 \$26 \$25 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$669 \$11 \$719 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$670 \$61 \$11 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$671 \$30 \$29 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$672 \$12 \$725 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$673 \$62 \$12 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$674 \$34 \$33 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$675 \$13 \$731 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$676 \$63 \$13 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$677 \$38 \$37 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$678 \$14 \$737 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$679 \$64 \$14 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$680 \$42 \$41 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$681 \$15 \$743 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$682 \$65 \$15 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$683 \$46 \$45 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$684 \$16 \$749 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$685 \$66 \$16 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$686 \$50 \$49 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$687 \$17 \$755 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$688 \$67 \$17 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$689 \$54 \$53 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$690 \$18 \$761 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$691 \$68 \$18 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$692 \$58 \$57 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$693 \$702 \$768 D VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$694 \$703 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$695 VSSD \$702 \$703 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$696 \$704 \$703 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$697 VSSD clks \$704 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$698 \$702 \$769 \$704 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$699 \$706 \$769 \$703 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$700 \$707 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$701 VSSD \$706 \$707 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$702 \$705 \$707 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$703 VSSD Set \$705 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$704 \$706 \$768 \$705 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$705 \$708 \$771 \$707 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$706 \$709 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$707 VSSD \$708 \$709 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$708 \$710 \$709 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$709 VSSD clks \$710 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$710 \$708 \$772 \$710 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$711 \$712 \$772 \$709 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$712 \$713 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$713 VSSD \$712 \$713 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$714 \$711 \$713 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$715 VSSD Set \$711 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$716 \$712 \$771 \$711 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$717 \$714 \$774 \$713 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$718 \$715 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$719 VSSD \$714 \$715 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$720 \$716 \$715 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$721 VSSD clks \$716 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$722 \$714 \$775 \$716 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$723 \$718 \$775 \$715 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$724 \$719 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$725 VSSD \$718 \$719 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$726 \$717 \$719 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$727 VSSD Set \$717 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$728 \$718 \$774 \$717 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$729 \$720 \$777 \$719 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$730 \$721 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$731 VSSD \$720 \$721 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$732 \$722 \$721 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$733 VSSD clks \$722 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$734 \$720 \$778 \$722 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$735 \$724 \$778 \$721 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$736 \$725 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$737 VSSD \$724 \$725 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$738 \$723 \$725 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$739 VSSD Set \$723 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$740 \$724 \$777 \$723 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$741 \$726 \$780 \$725 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$742 \$727 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$743 VSSD \$726 \$727 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$744 \$728 \$727 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$745 VSSD clks \$728 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$746 \$726 \$781 \$728 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$747 \$730 \$781 \$727 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$748 \$731 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$749 VSSD \$730 \$731 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$750 \$729 \$731 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$751 VSSD Set \$729 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$752 \$730 \$780 \$729 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$753 \$732 \$783 \$731 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$754 \$733 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$755 VSSD \$732 \$733 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$756 \$734 \$733 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$757 VSSD clks \$734 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$758 \$732 \$784 \$734 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$759 \$736 \$784 \$733 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$760 \$737 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$761 VSSD \$736 \$737 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$762 \$735 \$737 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$763 VSSD Set \$735 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$764 \$736 \$783 \$735 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$765 \$738 \$786 \$737 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$766 \$739 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$767 VSSD \$738 \$739 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$768 \$740 \$739 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$769 VSSD clks \$740 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$770 \$738 \$787 \$740 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$771 \$742 \$787 \$739 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$772 \$743 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$773 VSSD \$742 \$743 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$774 \$741 \$743 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$775 VSSD Set \$741 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$776 \$742 \$786 \$741 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$777 \$744 \$789 \$743 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$778 \$745 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$779 VSSD \$744 \$745 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$780 \$746 \$745 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$781 VSSD clks \$746 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$782 \$744 \$790 \$746 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$783 \$748 \$790 \$745 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$784 \$749 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$785 VSSD \$748 \$749 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$786 \$747 \$749 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$787 VSSD Set \$747 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$788 \$748 \$789 \$747 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$789 \$750 \$792 \$749 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$790 \$751 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$791 VSSD \$750 \$751 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$792 \$752 \$751 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$793 VSSD clks \$752 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$794 \$750 \$793 \$752 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$795 \$754 \$793 \$751 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$796 \$755 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$797 VSSD \$754 \$755 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$798 \$753 \$755 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$799 VSSD Set \$753 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$800 \$754 \$792 \$753 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$801 \$756 \$795 \$755 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$802 \$757 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$803 VSSD \$756 \$757 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$804 \$758 \$757 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$805 VSSD clks \$758 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$806 \$756 \$796 \$758 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$807 \$760 \$796 \$757 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$808 \$761 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$809 VSSD \$760 \$761 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$810 \$759 \$761 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$811 VSSD Set \$759 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$812 \$760 \$795 \$759 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$813 \$762 \$798 \$761 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$814 \$763 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$815 VSSD \$762 \$763 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$816 \$764 \$763 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$817 VSSD clks \$764 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$818 \$762 \$799 \$764 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$819 \$767 \$799 \$763 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$820 CK_1 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$821 VSSD \$767 CK_1 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$822 \$766 CK_1 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$823 VSSD Set \$766 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$824 \$767 \$798 \$766 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$825 \$768 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$826 \$769 \$768 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$827 \$770 \$707 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$828 \$771 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$829 \$772 \$771 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$830 \$620 \$2211 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$831 \$2211 \$2256 \$2215 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$832 VSSD \$2417 \$2211 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$833 \$2257 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$834 \$2258 \$2257 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$835 \$3032 \$3050 \$2987 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$836 \$773 \$713 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$837 \$3032 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$838 \$2216 \$2257 \$2215 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$839 \$774 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$840 VSSD \$2215 \$3032 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$841 \$2217 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$842 \$775 \$774 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$843 VSSD \$2216 \$2217 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$844 \$2215 \$2987 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$845 VSSD Reset \$2215 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$846 \$2218 \$2217 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$847 VSSD Reset \$2218 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$848 \$3033 \$3051 \$2987 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$849 \$2216 \$2258 \$2218 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$850 \$3034 \$3051 \$3022 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$851 \$2221 \$2258 \$2217 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$852 \$3034 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$853 VSSD \$3033 \$3034 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$854 \$2219 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$855 VSSD \$2221 \$2219 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$856 \$3033 \$3022 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$857 VSSD Set \$3033 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$858 \$2220 \$2219 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$859 vocp \$3050 \$3022 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$860 VSSD Set \$2220 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$861 \$2221 \$2257 \$2220 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$862 \$2259 \$2219 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$863 \$776 \$719 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$864 \$777 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$865 \$778 \$777 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$866 Bit_1 \$2222 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$867 \$2222 \$2260 \$2223 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$868 VSSD \$2431 \$2222 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$869 \$779 \$725 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$870 \$2261 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$871 \$780 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$872 \$2262 \$2261 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$873 \$3035 \$3054 \$2988 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$874 \$781 \$780 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$875 \$3035 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$876 \$2224 \$2261 \$2223 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$877 VSSD \$2223 \$3035 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$878 \$2225 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$879 VSSD \$2224 \$2225 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$880 \$2223 \$2988 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$881 VSSD Reset \$2223 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$882 \$2226 \$2225 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$883 VSSD Reset \$2226 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$884 \$3036 \$3055 \$2988 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$885 \$2224 \$2262 \$2226 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$886 \$3037 \$3055 \$3023 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$887 \$2229 \$2262 \$2225 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$888 \$3037 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$889 VSSD \$3036 \$3037 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$890 \$2227 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$891 VSSD \$2229 \$2227 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$892 \$3036 \$3023 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$893 VSSD Set \$3036 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$894 \$2228 \$2227 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$895 vocp \$3054 \$3023 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$896 VSSD Set \$2228 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$897 \$2229 \$2261 \$2228 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$898 \$2263 \$2227 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$899 \$782 \$731 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$900 \$783 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$901 \$784 \$783 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$902 Bit_2 \$2212 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$903 \$785 \$737 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$904 \$2212 \$2264 \$2230 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$905 VSSD \$2444 \$2212 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$906 \$786 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$907 \$787 \$786 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$908 \$2265 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$909 \$2266 \$2265 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$910 \$3038 \$3058 \$2989 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$911 \$3038 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$912 \$2231 \$2265 \$2230 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$913 VSSD \$2230 \$3038 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$914 \$2232 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$915 VSSD \$2231 \$2232 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$916 \$2230 \$2989 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$917 VSSD Reset \$2230 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$918 \$2233 \$2232 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$919 VSSD Reset \$2233 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$920 \$3039 \$3059 \$2989 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$921 \$2231 \$2266 \$2233 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$922 \$3040 \$3059 \$3024 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$923 \$2236 \$2266 \$2232 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$924 \$3040 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$925 VSSD \$3039 \$3040 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$926 \$2234 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$927 VSSD \$2236 \$2234 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$928 \$3039 \$3024 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$929 VSSD Set \$3039 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$930 \$2235 \$2234 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$931 vocp \$3058 \$3024 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$932 VSSD Set \$2235 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$933 \$788 \$743 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$934 \$2236 \$2265 \$2235 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$935 \$789 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$936 \$2267 \$2234 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$937 \$790 \$789 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$938 \$791 \$749 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$939 Bit_3 \$2213 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$940 \$792 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$941 \$793 \$792 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$942 \$2213 \$2268 \$2237 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$943 VSSD \$2457 \$2213 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$944 \$2269 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$945 \$2270 \$2269 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$946 \$3041 \$3062 \$2990 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$947 \$3041 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$948 \$2238 \$2269 \$2237 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$949 VSSD \$2237 \$3041 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$950 \$2239 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$951 VSSD \$2238 \$2239 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$952 \$2237 \$2990 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$953 VSSD Reset \$2237 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$954 \$2240 \$2239 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$955 VSSD Reset \$2240 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$956 \$3042 \$3063 \$2990 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$957 \$2238 \$2270 \$2240 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$958 \$3043 \$3063 \$3025 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$959 \$2243 \$2270 \$2239 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$960 \$3043 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$961 VSSD \$3042 \$3043 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$962 \$2241 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$963 VSSD \$2243 \$2241 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$964 \$3042 \$3025 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$965 \$794 \$755 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$966 VSSD Set \$3042 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$967 \$2242 \$2241 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$968 vocp \$3062 \$3025 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$969 VSSD Set \$2242 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$970 \$795 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$971 \$796 \$795 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$972 \$2243 \$2269 \$2242 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$973 \$2271 \$2241 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$974 \$797 \$761 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$975 \$798 Valid VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$976 \$799 \$798 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$977 Bit_4 \$2214 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$978 \$2214 \$2272 \$2244 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$979 VSSD \$2470 \$2214 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$980 \$2273 clks VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$981 \$2274 \$2273 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$982 \$3044 \$3066 \$2991 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$983 \$3044 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$984 \$2245 \$2273 \$2244 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$985 VSSD \$2244 \$3044 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$986 \$2246 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$987 VSSD \$2245 \$2246 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$988 \$2244 \$2991 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$989 VSSD Reset \$2244 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$990 \$2247 \$2246 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$991 VSSD Reset \$2247 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$992 \$3045 \$3067 \$2991 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$993 \$2245 \$2274 \$2247 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$994 \$3046 \$3067 \$3026 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$995 \$2250 \$2274 \$2246 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$996 \$800 CK_1 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$997 \$3046 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$998 VSSD \$3045 \$3046 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$999 \$2248 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1000 VSSD \$2250 \$2248 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1001 \$3045 \$3026 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1002 VSSD Set \$3045 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1003 \$2249 \$2248 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1004 vocp \$3066 \$3026 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1005 VSSD Set \$2249 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1006 \$2250 \$2273 \$2249 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1007 \$2275 \$2248 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1008 \$3983 \$4015 \$3938 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1009 \$3983 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1010 VSSD \$4016 \$3983 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1011 \$4016 \$3938 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1012 VSSD Reset \$4016 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1013 \$3984 \$4208 \$3938 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1014 \$3985 \$4208 \$3972 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1015 \$3985 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1016 VSSD \$3984 \$3985 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1017 \$3984 \$3972 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1018 VSSD Set \$3984 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1019 \$3986 \$4015 \$3972 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1020 \$3987 \$4017 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1021 \$3986 \$4217 \$3987 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1022 VSSD \$3987 Bit_10 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1023 \$620 \$2417 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1024 \$3048 \$2256 \$2215 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1025 \$3988 \$4019 \$3939 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1026 VSSD \$2215 \$3049 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1027 \$3988 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1028 VSSD \$4020 \$3988 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1029 \$4020 \$3939 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1030 VSSD Reset \$4020 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1031 \$3989 \$4230 \$3939 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1032 \$3990 \$4230 \$3973 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1033 \$3990 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1034 VSSD \$3989 \$3990 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1035 \$3989 \$3973 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1036 VSSD Set \$3989 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1037 \$3991 \$4019 \$3973 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1038 VSSD \$3050 \$3051 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1039 \$3974 \$4021 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1040 VSSD \$2256 \$3050 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1041 \$3991 \$4231 \$3974 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1042 VSSD \$2417 \$2256 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1043 VSSD \$3974 Bit_9 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1044 VSSD CK_1 \$2417 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1045 Bit_1 \$2431 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1046 \$3052 \$2260 \$2223 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1047 \$3992 \$4023 \$3940 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1048 VSSD \$2223 \$3053 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1049 \$3992 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1050 VSSD \$4024 \$3992 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1051 \$4024 \$3940 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1052 VSSD Reset \$4024 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1053 \$3993 \$4236 \$3940 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1054 \$3994 \$4236 \$3975 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1055 \$3994 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1056 VSSD \$3993 \$3994 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1057 \$3993 \$3975 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1058 VSSD Set \$3993 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1059 \$3995 \$4023 \$3975 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1060 VSSD \$3054 \$3055 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1061 \$3976 \$4025 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1062 VSSD \$2260 \$3054 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1063 \$3995 \$4245 \$3976 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1064 VSSD \$2431 \$2260 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1065 VSSD \$3976 Bit_8 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1066 VSSD \$761 \$2431 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1067 Bit_2 \$2444 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1068 \$3056 \$2264 \$2230 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1069 \$3996 \$4027 \$3941 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1070 VSSD \$2230 \$3057 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1071 \$3996 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1072 VSSD \$4028 \$3996 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1073 \$4028 \$3941 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1074 VSSD Reset \$4028 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1075 \$3997 \$4258 \$3941 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1076 \$3998 \$4258 \$3977 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1077 \$3998 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1078 VSSD \$3997 \$3998 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1079 \$3997 \$3977 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1080 VSSD Set \$3997 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1081 \$3999 \$4027 \$3977 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1082 VSSD \$3058 \$3059 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1083 \$3978 \$4029 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1084 VSSD \$2264 \$3058 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1085 \$3999 \$4259 \$3978 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1086 VSSD \$2444 \$2264 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1087 VSSD \$3978 Bit_7 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1088 VSSD \$755 \$2444 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1089 Bit_3 \$2457 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1090 \$3060 \$2268 \$2237 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1091 \$4000 \$4031 \$3942 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1092 VSSD \$2237 \$3061 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1093 \$4000 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1094 VSSD \$4032 \$4000 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1095 \$4032 \$3942 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1096 VSSD Reset \$4032 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1097 \$4001 \$4264 \$3942 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1098 \$4002 \$4264 \$3979 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1099 \$4002 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1100 VSSD \$4001 \$4002 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1101 \$4001 \$3979 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1102 VSSD Set \$4001 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1103 \$4003 \$4031 \$3979 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1104 VSSD \$3062 \$3063 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1105 \$3980 \$4033 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1106 VSSD \$2268 \$3062 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1107 \$4003 \$4273 \$3980 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1108 VSSD \$2457 \$2268 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1109 VSSD \$3980 Bit_6 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1110 VSSD \$749 \$2457 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1111 Bit_4 \$2470 VCM VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1112 \$3064 \$2272 \$2244 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1113 \$4004 \$4035 \$3943 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1114 VSSD \$2244 \$3065 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1115 \$4004 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1116 VSSD \$4036 \$4004 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1117 \$4036 \$3943 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1118 VSSD Reset \$4036 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1119 \$4005 \$4278 \$3943 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1120 \$4006 \$4278 \$3981 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1121 \$4006 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1122 VSSD \$4005 \$4006 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1123 \$4005 \$3981 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1124 VSSD Set \$4005 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1125 \$4007 \$4035 \$3981 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1126 VSSD \$3066 \$3067 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1127 \$3982 \$4037 VSSD VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1128 VSSD \$2272 \$3066 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1129 \$4007 \$4287 \$3982 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1130 VSSD \$2470 \$2272 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1131 VSSD \$3982 Bit_5 VSSD nfet_03v3 L=1.1U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1132 VSSD \$743 \$2470 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1133 VSSD \$4016 \$4014 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1134 \$4944 \$4974 vocp VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1135 \$4945 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1136 VSSD \$4944 \$4945 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1137 \$4946 \$4945 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1138 VSSD Reset \$4946 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1139 \$4944 \$5118 \$4946 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1140 \$4948 \$5118 \$4945 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1141 \$3986 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1142 VSSD \$4948 \$3986 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1143 \$4947 \$3986 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1144 VSSD Set \$4947 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1145 \$4948 \$4974 \$4947 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1146 VSSD \$4015 \$4208 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1147 VSSD clks \$4015 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1148 VSSD \$4020 \$4018 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1149 \$4949 \$4977 vocp VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1150 \$4950 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1151 VSSD \$4949 \$4950 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1152 \$4951 \$4950 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1153 VSSD Reset \$4951 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1154 \$4949 \$5119 \$4951 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1155 \$4953 \$5119 \$4950 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1156 \$3991 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1157 VSSD \$4953 \$3991 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1158 \$4952 \$3991 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1159 VSSD Set \$4952 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1160 \$4953 \$4977 \$4952 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1161 VSSD \$4019 \$4230 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1162 VSSD clks \$4019 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1163 VSSD \$4024 \$4022 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1164 \$4954 \$4980 vocp VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1165 \$4955 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1166 VSSD \$4954 \$4955 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1167 \$4956 \$4955 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1168 VSSD Reset \$4956 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1169 \$4954 \$5120 \$4956 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1170 \$4958 \$5120 \$4955 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1171 \$3995 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1172 VSSD \$4958 \$3995 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1173 \$4957 \$3995 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1174 VSSD Set \$4957 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1175 \$4958 \$4980 \$4957 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1176 VSSD \$4023 \$4236 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1177 VSSD clks \$4023 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1178 VSSD \$4028 \$4026 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1179 \$4959 \$4983 vocp VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1180 \$4960 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1181 VSSD \$4959 \$4960 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1182 \$4961 \$4960 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1183 VSSD Reset \$4961 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1184 \$4959 \$5121 \$4961 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1185 \$4963 \$5121 \$4960 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1186 \$3999 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1187 VSSD \$4963 \$3999 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1188 \$4962 \$3999 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1189 VSSD Set \$4962 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1190 \$4963 \$4983 \$4962 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1191 VSSD \$4027 \$4258 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1192 VSSD clks \$4027 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1193 VSSD \$4032 \$4030 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1194 \$4964 \$4986 vocp VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1195 \$4965 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1196 VSSD \$4964 \$4965 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1197 \$4966 \$4965 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1198 VSSD Reset \$4966 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1199 \$4964 \$5122 \$4966 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1200 \$4968 \$5122 \$4965 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1201 \$4003 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1202 VSSD \$4968 \$4003 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1203 \$4967 \$4003 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1204 VSSD Set \$4967 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1205 \$4968 \$4986 \$4967 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1206 VSSD \$4031 \$4264 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1207 VSSD clks \$4031 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1208 VSSD \$4036 \$4034 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1209 \$4969 \$4989 vocp VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1210 \$4970 Set VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1211 VSSD \$4969 \$4970 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1212 \$4971 \$4970 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1213 VSSD Reset \$4971 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1214 \$4969 \$5123 \$4971 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1215 \$4973 \$5123 \$4970 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1216 \$4007 Reset VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1217 VSSD \$4973 \$4007 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1218 \$4972 \$4007 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1219 VSSD Set \$4972 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1220 \$4973 \$4989 \$4972 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1221 VSSD \$4035 \$4278 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1222 VSSD clks \$4035 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1223 \$4017 \$707 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1224 \$4217 \$4017 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1225 \$4974 \$4217 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1226 \$5118 \$4974 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1227 \$4975 \$3986 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1228 \$3986 \$4217 \$4976 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1229 VCM \$4017 Bit_10 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1230 \$4021 \$713 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1231 \$4231 \$4021 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1232 \$4977 \$4231 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1233 \$5119 \$4977 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1234 \$4978 \$3991 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1235 \$3991 \$4231 \$4979 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1236 VCM \$4021 Bit_9 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1237 \$4025 \$719 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1238 \$4245 \$4025 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1239 \$4980 \$4245 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1240 \$5120 \$4980 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1241 \$4981 \$3995 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1242 \$3995 \$4245 \$4982 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1243 VCM \$4025 Bit_8 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1244 \$4029 \$725 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1245 \$4259 \$4029 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1246 \$4983 \$4259 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1247 \$5121 \$4983 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1248 \$4984 \$3999 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1249 \$3999 \$4259 \$4985 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1250 VCM \$4029 Bit_7 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1251 \$4033 \$731 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1252 \$4273 \$4033 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1253 \$4986 \$4273 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1254 \$5122 \$4986 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1255 \$4987 \$4003 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1256 \$4003 \$4273 \$4988 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1257 VCM \$4033 Bit_6 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1258 \$4037 \$737 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1259 \$4287 \$4037 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1260 \$4989 \$4287 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1261 \$5123 \$4989 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1262 \$4990 \$4007 VSSD VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
M$1263 \$4007 \$4287 \$4991 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P
+ AD=0.9516P PS=4.34U PD=4.34U
M$1264 VCM \$4037 Bit_5 VSSD nfet_03v3 L=0.28U W=1.56U AS=0.9516P AD=0.9516P
+ PS=4.34U PD=4.34U
.ENDS SAR_Asynchronous_top_neg_logic
