* NGSPICE file created from DiffP_net.ext - technology: gf180mcuD

.subckt DiffP_net IT VN VDD VP VSS OUT
X0 VSS.t75 VSS.t74 VSS.t75 VSS.t1 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X1 VSS.t73 VSS.t72 VSS.t73 VSS.t35 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2 a_1771_2657# a_n179_6700.t11 VSS.t76 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X3 VSS.t71 VSS.t70 VSS.t71 VSS.t20 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X4 a_367_1891# a_n179_6700.t12 OUT.t0 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X5 VDD.t71 VDD.t70 VDD.t71 VDD.t2 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X6 VSS a_n179_6700.t13 a_367_733# VSS.t2 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X7 VSS.t69 VSS.t68 VSS.t69 VSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X8 VSS.t67 VSS.t66 VSS.t67 VSS.t2 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X9 VSS a_n179_6700.t14 a_367_1891# VSS.t2 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X10 VSS.t65 VSS.t64 VSS.t65 VSS.t17 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X11 VSS.t63 VSS.t62 VSS.t63 VSS.t52 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X12 VSS.t61 VSS.t60 VSS.t61 VSS.t20 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X13 VSS.t59 VSS.t58 VSS.t59 VSS.t35 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X14 VSS.t57 VSS.t56 VSS.t57 VSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X15 VSS.t55 VSS.t54 VSS.t55 VSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X16 VDD.t69 VDD.t68 VDD.t69 VDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X17 VDD.t67 VDD.t66 VDD.t67 VDD.t39 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X18 VDD.t65 VDD.t64 VDD.t65 VDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X19 VDD.t63 VDD.t62 VDD.t63 VDD.t39 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X20 VSS.t53 VSS.t51 VSS.t53 VSS.t52 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X21 VSS.t50 VSS.t49 VSS.t50 VSS.t20 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X22 a_1771_1891# a_n179_6700.t15 VSS.t83 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X23 VSS.t48 VSS.t47 VSS.t48 VSS.t20 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X24 VSS.t46 VSS.t45 VSS.t46 VSS.t35 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X25 VDD.t61 VDD.t60 VDD.t61 VDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X26 VDD.t59 VDD.t58 VDD.t59 VDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X27 VSS.t44 VSS.t43 VSS.t44 VSS.t35 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X28 VSS.t42 VSS.t41 VSS.t42 VSS.t35 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X29 IT VN.t0 a_351_9798# VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X30 VDD.t57 VDD.t56 VDD.t57 VDD.t39 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X31 IT VN.t1 a_351_7866# VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X32 VDD.t55 VDD.t54 VDD.t55 VDD.t39 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X33 a_367_733# a_n179_6700.t9 a_n179_6700.t10 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X34 VDD.t53 VDD.t52 VDD.t53 VDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X35 VDD.t51 VDD.t50 VDD.t51 VDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X36 VDD.t49 VDD.t48 VDD.t49 VDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X37 VDD.t47 VDD.t46 VDD.t47 VDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X38 VDD.t45 VDD.t43 VDD.t45 VDD.t44 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X39 VDD.t42 VDD.t41 VDD.t42 VDD.t39 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X40 a_1771_733# a_n179_6700.t16 VSS.t79 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X41 VDD.t40 VDD.t38 VDD.t40 VDD.t39 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X42 IT VP.t0 a_351_8632# VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X43 VDD.t37 VDD.t36 VDD.t37 VDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X44 IT VP.t1 a_351_6700# VDD.t3 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X45 VDD.t35 VDD.t34 VDD.t35 VDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X46 VDD.t33 VDD.t32 VDD.t33 VDD.t11 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X47 VDD.t31 VDD.t30 VDD.t31 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X48 VDD.t29 VDD.t28 VDD.t29 VDD.t3 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X49 VDD.t27 VDD.t26 VDD.t27 VDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X50 a_351_9798# VN.t2 OUT.t5 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X51 VDD.t25 VDD.t24 VDD.t25 VDD.t11 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X52 a_351_7866# VN.t3 OUT.t6 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X53 VDD.t23 VDD.t22 VDD.t23 VDD.t11 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X54 a_1757_9798# VP.t4 IT.t0 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X55 a_1757_7866# VP.t5 IT.t6 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X56 OUT a_n179_6700.t18 a_1771_733# VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X57 VSS.t40 VSS.t39 VSS.t40 VSS.t17 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X58 OUT a_n179_6700.t19 a_1771_2657# VSS.t0 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X59 a_351_8632# VP.t6 a_n179_6700.t0 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X60 OUT VN.t4 a_1757_8632# VDD.t2 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X61 VDD.t21 VDD.t20 VDD.t21 VDD.t11 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X62 a_351_6700# VP.t7 a_n179_6700.t0 VDD.t1 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X63 OUT VN.t5 a_1757_6700# VDD.t2 pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X64 VDD.t19 VDD.t18 VDD.t19 VDD.t11 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X65 a_367_3815# a_n179_6700.t20 OUT.t1 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X66 a_1757_8632# VN.t6 IT.t3 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X67 a_1757_6700# VN.t7 IT.t2 VDD.t0 pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X68 VSS.t38 VSS.t37 VSS.t38 VSS.t17 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X69 VSS.t36 VSS.t34 VSS.t36 VSS.t35 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X70 VSS.t33 VSS.t32 VSS.t33 VSS.t0 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X71 VDD.t17 VDD.t15 VDD.t17 VDD.t16 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X72 VDD.t14 VDD.t13 VDD.t14 VDD.t2 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X73 VDD.t12 VDD.t10 VDD.t12 VDD.t11 pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X74 VSS a_n179_6700.t21 a_367_3815# VSS.t2 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X75 VSS.t31 VSS.t30 VSS.t31 VSS.t20 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X76 VSS.t29 VSS.t28 VSS.t29 VSS.t17 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X77 VDD.t9 VDD.t8 VDD.t9 VDD.t1 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X78 VDD.t7 VDD.t6 VDD.t7 VDD.t1 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X79 a_367_2657# a_n179_6700.t7 a_n179_6700.t8 VSS.t1 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X80 VDD.t5 VDD.t4 VDD.t5 VDD.t0 pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X81 VSS.t27 VSS.t26 VSS.t27 VSS.t0 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X82 VSS.t25 VSS.t24 VSS.t25 VSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X83 a_1771_3815# a_n179_6700.t22 VSS.t80 VSS.t52 nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X84 VSS.t23 VSS.t22 VSS.t23 VSS.t17 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X85 VSS.t21 VSS.t19 VSS.t21 VSS.t20 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X86 VSS.t18 VSS.t16 VSS.t18 VSS.t17 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X87 VSS.t15 VSS.t14 VSS.t15 VSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X88 VSS.t13 VSS.t12 VSS.t13 VSS.t1 nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X89 VSS a_n179_6700.t24 a_367_2657# VSS.t2 nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X90 VSS.t11 VSS.t9 VSS.t11 VSS.t10 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X91 VSS.t8 VSS.t7 VSS.t8 VSS.t2 nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
R0 VSS.n72 VSS.n6 523.342
R1 VSS.n75 VSS.n5 521.869
R2 VSS.n72 VSS.n5 519.659
R3 VSS.n75 VSS.n6 516.342
R4 VSS.t0 VSS.t20 442.449
R5 VSS.t1 VSS.t10 442.449
R6 VSS.t20 VSS.t35 301.425
R7 VSS.t52 VSS.t0 301.425
R8 VSS.t2 VSS.t1 301.425
R9 VSS.t10 VSS.t17 301.425
R10 VSS.t35 VSS.n5 251.454
R11 VSS.t17 VSS.n6 251.454
R12 VSS.n73 VSS.t52 216.381
R13 VSS.n74 VSS.t2 210.998
R14 VSS.n74 VSS.n73 26.9134
R15 VSS.n18 VSS.t49 8.06917
R16 VSS.n18 VSS.t43 8.06917
R17 VSS.n16 VSS.t19 8.06917
R18 VSS.n16 VSS.t72 8.06917
R19 VSS.n15 VSS.t70 8.06917
R20 VSS.n15 VSS.t58 8.06917
R21 VSS.n0 VSS.t47 8.06917
R22 VSS.n0 VSS.t41 8.06917
R23 VSS.n85 VSS.t30 8.06917
R24 VSS.n85 VSS.t34 8.06917
R25 VSS.n83 VSS.t60 8.06917
R26 VSS.n83 VSS.t45 8.06917
R27 VSS.n67 VSS.t74 8.06917
R28 VSS.n25 VSS.t66 8.06917
R29 VSS.n7 VSS.t51 8.06917
R30 VSS.n21 VSS.t26 8.06917
R31 VSS.n64 VSS.t22 8.06917
R32 VSS.n64 VSS.t56 8.06917
R33 VSS.n62 VSS.t39 8.06917
R34 VSS.n62 VSS.t24 8.06917
R35 VSS.n61 VSS.t37 8.06917
R36 VSS.n61 VSS.t9 8.06917
R37 VSS.n57 VSS.t16 8.06917
R38 VSS.n57 VSS.t54 8.06917
R39 VSS.n56 VSS.t64 8.06917
R40 VSS.n56 VSS.t14 8.06917
R41 VSS.n54 VSS.t28 8.06917
R42 VSS.n54 VSS.t68 8.06917
R43 VSS.n49 VSS.t12 8.06917
R44 VSS.n48 VSS.t7 8.06917
R45 VSS.n78 VSS.t62 8.06917
R46 VSS.n3 VSS.t32 8.06917
R47 VSS.n38 VSS.n37 4.61205
R48 VSS.n45 VSS.n44 4.61205
R49 VSS.n35 VSS.n33 4.5005
R50 VSS.n42 VSS.n40 4.5005
R51 VSS.n32 VSS.t76 4.16278
R52 VSS.n39 VSS.t79 4.16278
R53 VSS.n37 VSS.n36 4.15984
R54 VSS.n44 VSS.n43 4.15984
R55 VSS.n46 VSS.n38 3.98482
R56 VSS.n47 VSS.n46 3.97971
R57 VSS.n32 VSS.t80 3.93054
R58 VSS.n39 VSS.t83 3.93054
R59 VSS.n35 VSS.n34 3.92774
R60 VSS.n42 VSS.n41 3.92774
R61 VSS.n66 VSS.t75 3.3605
R62 VSS.n70 VSS.t67 3.3605
R63 VSS.n24 VSS.t53 3.3605
R64 VSS.n20 VSS.t27 3.3605
R65 VSS.n52 VSS.t13 3.3605
R66 VSS.t8 VSS.n4 3.3605
R67 VSS.n77 VSS.t63 3.3605
R68 VSS.n81 VSS.t33 3.3605
R69 VSS.n46 VSS.n45 3.27473
R70 VSS.n33 VSS.n32 2.68012
R71 VSS.n40 VSS.n39 2.68012
R72 VSS.n80 VSS.n79 2.1005
R73 VSS.n51 VSS.n50 2.1005
R74 VSS.n23 VSS.n22 2.1005
R75 VSS.n69 VSS.n68 2.1005
R76 VSS.t67 VSS.n69 1.2605
R77 VSS.n69 VSS.t75 1.2605
R78 VSS.n23 VSS.t27 1.2605
R79 VSS.t53 VSS.n23 1.2605
R80 VSS.n51 VSS.t8 1.2605
R81 VSS.t13 VSS.n51 1.2605
R82 VSS.t33 VSS.n80 1.2605
R83 VSS.n80 VSS.t63 1.2605
R84 VSS.n8 VSS.t44 0.918039
R85 VSS.n9 VSS.t73 0.918039
R86 VSS.n10 VSS.t59 0.918039
R87 VSS.n11 VSS.t42 0.918039
R88 VSS.n1 VSS.t36 0.918039
R89 VSS.n2 VSS.t46 0.918039
R90 VSS.n26 VSS.t57 0.918039
R91 VSS.n27 VSS.t25 0.918039
R92 VSS.n28 VSS.t11 0.918039
R93 VSS.n29 VSS.t55 0.918039
R94 VSS.n30 VSS.t15 0.918039
R95 VSS.n31 VSS.t69 0.918039
R96 VSS.n8 VSS.t50 0.91749
R97 VSS.n9 VSS.t21 0.91749
R98 VSS.n10 VSS.t71 0.91749
R99 VSS.n11 VSS.t48 0.91749
R100 VSS.n1 VSS.t31 0.91749
R101 VSS.n2 VSS.t61 0.91749
R102 VSS.n26 VSS.t23 0.91749
R103 VSS.n27 VSS.t40 0.91749
R104 VSS.n28 VSS.t38 0.91749
R105 VSS.n29 VSS.t18 0.91749
R106 VSS.n30 VSS.t65 0.91749
R107 VSS.n31 VSS.t29 0.91749
R108 VSS.n53 VSS.n31 0.582999
R109 VSS.n55 VSS.n30 0.582999
R110 VSS.n58 VSS.n29 0.582999
R111 VSS.n60 VSS.n28 0.582999
R112 VSS.n63 VSS.n27 0.582999
R113 VSS.n65 VSS.n26 0.582999
R114 VSS.n82 VSS.n2 0.582999
R115 VSS.n84 VSS.n1 0.582999
R116 VSS.n12 VSS.n11 0.582999
R117 VSS.n14 VSS.n10 0.582999
R118 VSS.n17 VSS.n9 0.582999
R119 VSS.n19 VSS.n8 0.582999
R120 VSS.n38 VSS.n33 0.157683
R121 VSS.n45 VSS.n40 0.157683
R122 VSS.n59 VSS.n6 0.0886356
R123 VSS.n72 VSS.n71 0.0886356
R124 VSS.n73 VSS.n72 0.0886356
R125 VSS.n13 VSS.n5 0.0886356
R126 VSS.n76 VSS.n75 0.0871667
R127 VSS.n75 VSS.n74 0.0871667
R128 VSS.n64 VSS.n63 0.0390622
R129 VSS.n55 VSS.n54 0.0390622
R130 VSS.n18 VSS.n17 0.0385696
R131 VSS.n84 VSS.n83 0.0385696
R132 VSS.n62 VSS.n61 0.0371211
R133 VSS.n57 VSS.n56 0.0371211
R134 VSS.n16 VSS.n15 0.0366533
R135 VSS.n21 VSS.n20 0.0341
R136 VSS.n22 VSS.n21 0.0341
R137 VSS.n22 VSS.n7 0.0341
R138 VSS.n24 VSS.n7 0.0341
R139 VSS.n70 VSS.n25 0.0341
R140 VSS.n68 VSS.n25 0.0341
R141 VSS.n68 VSS.n67 0.0341
R142 VSS.n67 VSS.n66 0.0341
R143 VSS.n53 VSS.n52 0.0302339
R144 VSS.n60 VSS.n59 0.0301981
R145 VSS.n82 VSS.n81 0.0301505
R146 VSS.n66 VSS.n65 0.0300328
R147 VSS.n20 VSS.n19 0.0299989
R148 VSS.n14 VSS.n13 0.0298187
R149 VSS.n81 VSS.n3 0.0294988
R150 VSS.n79 VSS.n3 0.0294988
R151 VSS.n79 VSS.n78 0.0294988
R152 VSS.n78 VSS.n77 0.0294988
R153 VSS.n48 VSS.n4 0.0294988
R154 VSS.n50 VSS.n48 0.0294988
R155 VSS.n50 VSS.n49 0.0294988
R156 VSS.n52 VSS.n47 0.0221222
R157 VSS VSS.n0 0.0217704
R158 VSS.n59 VSS.n58 0.0203634
R159 VSS.n13 VSS.n12 0.0201097
R160 VSS.n71 VSS.n70 0.01994
R161 VSS.n65 VSS.n64 0.0196517
R162 VSS.n63 VSS.n62 0.0196517
R163 VSS.n61 VSS.n60 0.0196517
R164 VSS.n58 VSS.n57 0.0196517
R165 VSS.n56 VSS.n55 0.0196517
R166 VSS.n54 VSS.n53 0.0196517
R167 VSS.n19 VSS.n18 0.019407
R168 VSS.n17 VSS.n16 0.019407
R169 VSS.n15 VSS.n14 0.019407
R170 VSS.n12 VSS.n0 0.019407
R171 VSS.n85 VSS.n84 0.019407
R172 VSS.n83 VSS.n82 0.019407
R173 VSS.n77 VSS.n76 0.0183136
R174 VSS VSS.n85 0.0153829
R175 VSS.n71 VSS.n24 0.01514
R176 VSS.n76 VSS.n4 0.0120995
R177 VSS.n49 VSS.n47 0.0108347
R178 VSS.n37 VSS.n35 0.00523684
R179 VSS.n44 VSS.n42 0.00523684
R180 a_n179_6700.n1 a_n179_6700.t3 10.2515
R181 a_n179_6700.n1 a_n179_6700.t5 10.2515
R182 a_n179_6700.n1 a_n179_6700.t19 10.2515
R183 a_n179_6700.n1 a_n179_6700.t18 10.2515
R184 a_n179_6700.n1 a_n179_6700.t9 10.096
R185 a_n179_6700.n1 a_n179_6700.t12 10.0935
R186 a_n179_6700.n1 a_n179_6700.t7 10.0859
R187 a_n179_6700.n1 a_n179_6700.t20 10.0808
R188 a_n179_6700.n1 a_n179_6700.t13 9.53981
R189 a_n179_6700.n1 a_n179_6700.t21 9.53981
R190 a_n179_6700.n1 a_n179_6700.t14 9.53981
R191 a_n179_6700.n1 a_n179_6700.t24 9.53981
R192 a_n179_6700.n1 a_n179_6700.t16 9.53744
R193 a_n179_6700.n1 a_n179_6700.t22 9.53744
R194 a_n179_6700.n1 a_n179_6700.t15 9.53744
R195 a_n179_6700.n1 a_n179_6700.t11 9.53744
R196 a_n179_6700.n1 a_n179_6700.n0 8.41434
R197 a_n179_6700.n1 a_n179_6700.n3 8.14082
R198 a_n179_6700.n0 a_n179_6700.n4 8.13828
R199 a_n179_6700.t0 a_n179_6700.n5 7.91099
R200 a_n179_6700.t0 a_n179_6700.n2 7.91099
R201 a_n179_6700.t0 a_n179_6700.n1 7.50545
R202 a_n179_6700.n0 a_n179_6700.t10 7.48586
R203 a_n179_6700.n1 a_n179_6700.t8 7.48333
R204 OUT.n3 OUT.t5 10.5425
R205 OUT.n6 OUT.t1 9.99909
R206 OUT.n5 OUT.n4 9.47655
R207 OUT.n2 OUT.t6 7.77927
R208 OUT.n8 OUT.t0 7.74799
R209 OUT.n8 OUT.n7 7.46478
R210 OUT.n2 OUT.n1 7.08235
R211 OUT OUT.n9 6.58315
R212 OUT OUT.n0 3.62813
R213 OUT.n9 OUT.n8 2.2505
R214 OUT.n3 OUT.n2 2.2505
R215 OUT.n6 OUT.n5 0.797
R216 OUT.n5 OUT.n3 0.7685
R217 OUT.n9 OUT.n6 0.723125
R218 VDD.n59 VDD.n5 477.971
R219 VDD.n56 VDD.n6 470.842
R220 VDD.n59 VDD.n6 470.842
R221 VDD.n56 VDD.n5 469.683
R222 VDD.t2 VDD.t16 142.93
R223 VDD.t1 VDD.t39 142.93
R224 VDD.t16 VDD.t11 96.8792
R225 VDD.t0 VDD.t2 96.8792
R226 VDD.t3 VDD.t1 96.8792
R227 VDD.t39 VDD.t44 96.8792
R228 VDD.t11 VDD.n5 81.1238
R229 VDD.t44 VDD.n6 81.1238
R230 VDD.n57 VDD.t0 70.2717
R231 VDD.n58 VDD.t3 64.1315
R232 VDD.n58 VDD.n57 8.52856
R233 VDD.n18 VDD.t15 8.10567
R234 VDD.n18 VDD.t32 8.10567
R235 VDD.n16 VDD.t52 8.10567
R236 VDD.n16 VDD.t24 8.10567
R237 VDD.n15 VDD.t36 8.10567
R238 VDD.n15 VDD.t20 8.10567
R239 VDD.n0 VDD.t48 8.10567
R240 VDD.n0 VDD.t22 8.10567
R241 VDD.n69 VDD.t34 8.10567
R242 VDD.n69 VDD.t18 8.10567
R243 VDD.n67 VDD.t26 8.10567
R244 VDD.n67 VDD.t10 8.10567
R245 VDD.n51 VDD.t8 8.10567
R246 VDD.n25 VDD.t30 8.10567
R247 VDD.n7 VDD.t58 8.10567
R248 VDD.n21 VDD.t70 8.10567
R249 VDD.n48 VDD.t60 8.10567
R250 VDD.n48 VDD.t38 8.10567
R251 VDD.n46 VDD.t68 8.10567
R252 VDD.n46 VDD.t66 8.10567
R253 VDD.n45 VDD.t50 8.10567
R254 VDD.n45 VDD.t56 8.10567
R255 VDD.n41 VDD.t64 8.10567
R256 VDD.n41 VDD.t62 8.10567
R257 VDD.n40 VDD.t46 8.10567
R258 VDD.n40 VDD.t54 8.10567
R259 VDD.n38 VDD.t43 8.10567
R260 VDD.n38 VDD.t41 8.10567
R261 VDD.n32 VDD.t6 8.10567
R262 VDD.n33 VDD.t28 8.10567
R263 VDD.n62 VDD.t4 8.10567
R264 VDD.n3 VDD.t13 8.10567
R265 VDD.n50 VDD.t9 3.20383
R266 VDD.n54 VDD.t31 3.20383
R267 VDD.n24 VDD.t59 3.20383
R268 VDD.n20 VDD.t71 3.20383
R269 VDD.n36 VDD.t7 3.20383
R270 VDD.t29 VDD.n4 3.20383
R271 VDD.n61 VDD.t5 3.20383
R272 VDD.n65 VDD.t14 3.20383
R273 VDD.n64 VDD.n63 1.73383
R274 VDD.n35 VDD.n34 1.73383
R275 VDD.n23 VDD.n22 1.73383
R276 VDD.n53 VDD.n52 1.73383
R277 VDD.t31 VDD.n53 1.4705
R278 VDD.n53 VDD.t9 1.4705
R279 VDD.n23 VDD.t71 1.4705
R280 VDD.t59 VDD.n23 1.4705
R281 VDD.n35 VDD.t29 1.4705
R282 VDD.t7 VDD.n35 1.4705
R283 VDD.t14 VDD.n64 1.4705
R284 VDD.n64 VDD.t5 1.4705
R285 VDD.n8 VDD.t33 1.00929
R286 VDD.n9 VDD.t25 1.00929
R287 VDD.n10 VDD.t21 1.00929
R288 VDD.n11 VDD.t23 1.00929
R289 VDD.n1 VDD.t19 1.00929
R290 VDD.n2 VDD.t12 1.00929
R291 VDD.n26 VDD.t40 1.00929
R292 VDD.n27 VDD.t67 1.00929
R293 VDD.n28 VDD.t57 1.00929
R294 VDD.n29 VDD.t63 1.00929
R295 VDD.n30 VDD.t55 1.00929
R296 VDD.n31 VDD.t42 1.00929
R297 VDD.n8 VDD.t17 1.00871
R298 VDD.n9 VDD.t53 1.00871
R299 VDD.n10 VDD.t37 1.00871
R300 VDD.n11 VDD.t49 1.00871
R301 VDD.n1 VDD.t35 1.00871
R302 VDD.n2 VDD.t27 1.00871
R303 VDD.n26 VDD.t61 1.00871
R304 VDD.n27 VDD.t69 1.00871
R305 VDD.n28 VDD.t51 1.00871
R306 VDD.n29 VDD.t65 1.00871
R307 VDD.n30 VDD.t47 1.00871
R308 VDD.n31 VDD.t45 1.00871
R309 VDD.n37 VDD.n31 0.468749
R310 VDD.n39 VDD.n30 0.468749
R311 VDD.n42 VDD.n29 0.468749
R312 VDD.n44 VDD.n28 0.468749
R313 VDD.n47 VDD.n27 0.468749
R314 VDD.n49 VDD.n26 0.468749
R315 VDD.n66 VDD.n2 0.468749
R316 VDD.n68 VDD.n1 0.468749
R317 VDD.n12 VDD.n11 0.468749
R318 VDD.n14 VDD.n10 0.468749
R319 VDD.n17 VDD.n9 0.468749
R320 VDD.n19 VDD.n8 0.468749
R321 VDD.n43 VDD.n6 0.10728
R322 VDD.n56 VDD.n55 0.10728
R323 VDD.n57 VDD.n56 0.10728
R324 VDD.n13 VDD.n5 0.10728
R325 VDD.n60 VDD.n59 0.1055
R326 VDD.n59 VDD.n58 0.1055
R327 VDD.n48 VDD.n47 0.0382419
R328 VDD.n39 VDD.n38 0.0382419
R329 VDD.n18 VDD.n17 0.0382419
R330 VDD.n68 VDD.n67 0.0382419
R331 VDD.n46 VDD.n45 0.0364748
R332 VDD.n41 VDD.n40 0.0364748
R333 VDD.n16 VDD.n15 0.0364748
R334 VDD.n21 VDD.n20 0.0346711
R335 VDD.n22 VDD.n21 0.0346711
R336 VDD.n22 VDD.n7 0.0346711
R337 VDD.n24 VDD.n7 0.0346711
R338 VDD.n54 VDD.n25 0.0346711
R339 VDD.n52 VDD.n25 0.0346711
R340 VDD.n52 VDD.n51 0.0346711
R341 VDD.n51 VDD.n50 0.0346711
R342 VDD.n66 VDD.n65 0.0308563
R343 VDD.n37 VDD.n36 0.0308563
R344 VDD.n50 VDD.n49 0.0308128
R345 VDD.n20 VDD.n19 0.0308128
R346 VDD.n65 VDD.n3 0.0293162
R347 VDD.n63 VDD.n3 0.0293162
R348 VDD.n63 VDD.n62 0.0293162
R349 VDD.n62 VDD.n61 0.0293162
R350 VDD.n33 VDD.n4 0.0293162
R351 VDD.n34 VDD.n33 0.0293162
R352 VDD.n34 VDD.n32 0.0293162
R353 VDD.n36 VDD.n32 0.0293162
R354 VDD.n44 VDD.n43 0.0270708
R355 VDD.n14 VDD.n13 0.0270708
R356 VDD VDD.n0 0.0247356
R357 VDD.n43 VDD.n42 0.0222742
R358 VDD.n13 VDD.n12 0.0222742
R359 VDD.n49 VDD.n48 0.0193079
R360 VDD.n47 VDD.n46 0.0193079
R361 VDD.n45 VDD.n44 0.0193079
R362 VDD.n42 VDD.n41 0.0193079
R363 VDD.n40 VDD.n39 0.0193079
R364 VDD.n38 VDD.n37 0.0193079
R365 VDD.n19 VDD.n18 0.0193079
R366 VDD.n17 VDD.n16 0.0193079
R367 VDD.n15 VDD.n14 0.0193079
R368 VDD.n12 VDD.n0 0.0193079
R369 VDD.n69 VDD.n68 0.0193079
R370 VDD.n67 VDD.n66 0.0193079
R371 VDD.n61 VDD.n60 0.0185609
R372 VDD.n55 VDD.n54 0.0175856
R373 VDD.n55 VDD.n24 0.0159011
R374 VDD VDD.n69 0.0122391
R375 VDD.n60 VDD.n4 0.00983484
R376 VN.n3 VN.t7 8.44198
R377 VN.n3 VN.t5 8.44198
R378 VN.n5 VN.t6 8.44198
R379 VN.n5 VN.t4 8.44198
R380 VN.n6 VN.t2 8.10925
R381 VN.n18 VN.t3 8.10567
R382 VN.n2 VN.t1 8.10567
R383 VN.n7 VN.t0 8.10567
R384 VN VN.n20 4.74531
R385 VN.n19 VN.n18 4.64261
R386 VN.n2 VN.n1 4.63432
R387 VN.n7 VN.n4 4.63432
R388 VN.n20 VN.n0 4.5005
R389 VN.n12 VN.n4 3.48966
R390 VN.n13 VN.n1 3.43191
R391 VN.n14 VN.n3 2.78312
R392 VN.n11 VN.n5 2.78312
R393 VN.n16 VN.n15 2.36376
R394 VN.n10 VN.n9 2.36376
R395 VN.n14 VN.n13 2.30825
R396 VN.n10 VN.n6 2.29458
R397 VN.n15 VN.n0 2.29243
R398 VN.n17 VN.n16 2.25205
R399 VN.n9 VN.n8 2.25205
R400 VN.n12 VN.n11 2.2505
R401 VN.n8 VN.n6 2.09285
R402 VN.n15 VN.n14 1.34566
R403 VN.n11 VN.n10 1.34566
R404 VN.n13 VN.n12 0.66725
R405 VN.n19 VN.n17 0.476265
R406 VN.n8 VN.n4 0.234207
R407 VN.n17 VN.n1 0.234207
R408 VN.n20 VN.n19 0.157683
R409 VN VN.n0 0.0597105
R410 VN.n16 VN.n2 0.00997368
R411 VN.n9 VN.n7 0.00997368
R412 VN.n18 VN.n0 0.00523684
R413 IT.n2 IT.t0 6.52632
R414 IT.n9 IT.t2 6.39955
R415 IT.n2 IT.n1 5.96327
R416 IT.n8 IT.n2 4.07346
R417 IT.n9 IT.n8 3.98123
R418 IT.n6 IT.n4 3.73554
R419 IT.n3 IT.t3 3.73554
R420 IT.n6 IT.n5 3.57923
R421 IT.n3 IT.t6 3.57923
R422 IT IT.n0 3.47265
R423 IT.n8 IT.n7 3.39848
R424 IT.n7 IT.n3 2.58435
R425 IT IT.n9 2.3644
R426 IT.n7 IT.n6 2.22754
R427 VP.n7 VP.t2 11.5068
R428 VP.n2 VP.t3 11.5068
R429 VP.n7 VP.t4 10.7772
R430 VP.n2 VP.t5 10.7772
R431 VP.n6 VP.t6 8.10766
R432 VP.n1 VP.t7 8.10567
R433 VP.n16 VP.t1 8.10567
R434 VP.n9 VP.t0 8.10567
R435 VP.n24 VP.n23 4.79742
R436 VP.n9 VP.n5 4.7915
R437 VP.n16 VP.n15 4.7915
R438 VP.n12 VP.n11 4.64734
R439 VP.n19 VP.n18 4.64734
R440 VP VP.n0 4.57511
R441 VP.n11 VP.n5 4.5005
R442 VP.n18 VP.n15 4.5005
R443 VP.n25 VP.n24 4.5005
R444 VP.n17 VP.n3 2.38035
R445 VP.n10 VP.n8 2.38035
R446 VP.n14 VP.n4 2.31238
R447 VP.n21 VP.n20 2.31238
R448 VP.n14 VP.n13 2.2505
R449 VP.n22 VP.n21 2.2505
R450 VP.n6 VP.n4 2.20772
R451 VP.n23 VP.n22 2.20362
R452 VP.n12 VP.n6 2.00763
R453 VP.n8 VP.n7 1.05605
R454 VP.n3 VP.n2 1.05605
R455 VP.n21 VP.n14 0.663125
R456 VP.n19 VP.n0 0.389655
R457 VP.n24 VP.n0 0.157683
R458 VP.n8 VP.n4 0.118858
R459 VP.n22 VP.n3 0.118858
R460 VP.n13 VP.n5 0.114585
R461 VP.n20 VP.n15 0.114585
R462 VP VP.n25 0.0727368
R463 VP.n13 VP.n12 0.0435986
R464 VP.n20 VP.n19 0.0435986
R465 VP.n11 VP.n10 0.00760526
R466 VP.n18 VP.n17 0.00760526
R467 VP.n10 VP.n9 0.00642105
R468 VP.n17 VP.n16 0.00642105
R469 VP.n23 VP.n1 0.00523684
R470 VP.n25 VP.n1 0.00286842
C0 IT a_351_7866# 0.055781f
C1 a_1771_3815# OUT 0.023318f
C2 a_1771_733# OUT 0.05062f
C3 VN VDD 5.66978f
C4 VP a_1757_8632# 0.013454f
C5 VN a_1757_9798# 0.06302f
C6 VDD OUT 2.47667f
C7 a_1757_9798# OUT 0.017032f
C8 VP VN 3.21018f
C9 VP OUT 0.999978f
C10 VDD a_351_6700# 0.029536f
C11 IT a_1757_6700# 0.042056f
C12 a_367_1891# OUT 0.042182f
C13 VP a_351_6700# 0.112267f
C14 VN a_351_7866# 0.093125f
C15 a_351_7866# OUT 0.029087f
C16 VDD a_1757_9798# 0.024759f
C17 VP VDD 5.58399f
C18 VN a_1757_6700# 0.144764f
C19 IT a_351_8632# 0.042212f
C20 VP a_1757_9798# 0.077197f
C21 a_1757_6700# OUT 0.031959f
C22 a_367_733# OUT 0.012591f
C23 VDD a_351_7866# 0.017204f
C24 IT a_1757_7866# 0.042616f
C25 VP a_351_7866# 0.019637f
C26 a_351_8632# OUT 0.013857f
C27 VDD a_1757_6700# 0.021515f
C28 a_1771_1891# OUT 0.023412f
C29 VP a_1757_6700# 0.013454f
C30 IT a_351_9798# 0.04226f
C31 VN a_1757_7866# 0.065048f
C32 VDD a_351_8632# 0.017204f
C33 IT a_1757_8632# 0.029048f
C34 a_367_3815# OUT 0.042089f
C35 VP a_351_8632# 0.112267f
C36 VN IT 1.39374f
C37 VN a_351_9798# 0.093125f
C38 IT OUT 4.41873f
C39 a_351_9798# OUT 0.042426f
C40 VDD a_1757_7866# 0.012306f
C41 IT a_351_6700# 0.055221f
C42 a_1771_2657# OUT 0.038791f
C43 VP a_1757_7866# 0.077197f
C44 VN a_1757_8632# 0.14651f
C45 a_1757_8632# OUT 0.045043f
C46 VN OUT 2.3496f
C47 VDD IT 2.51055f
C48 VDD a_351_9798# 0.029536f
C49 IT a_1757_9798# 0.029095f
C50 VP IT 2.11529f
C51 VP a_351_9798# 0.019637f
.ends

