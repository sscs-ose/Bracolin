* Extracted by KLayout with GF180MCU LVS runset on : 24/12/2023 18:44

.SUBCKT CM_input ISBCS IP IP2 VDD IN IN2 VSS
M$1 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$3 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$4 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$5 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$6 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$7 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$8 \$63 \$58 IN VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$9 VDD \$58 \$63 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$10 \$64 \$58 VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$11 IN2 \$58 \$64 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$12 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$13 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$14 \$71 \$58 \$58 VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$15 VDD \$58 \$71 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$16 \$72 \$58 VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$17 \$58 \$58 \$72 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$18 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$19 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$20 \$80 \$58 IN2 VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$21 VDD \$58 \$80 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$22 \$81 \$58 VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$23 IN \$58 \$81 VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$24 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$25 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$26 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$27 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$28 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=0.84P PS=5.3U PD=2.84U
M$29 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=0.84P AD=1.3P PS=2.84U PD=5.3U
M$30 VDD VDD VDD VDD pfet_03v3 L=6U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$31 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$32 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$33 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$34 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$35 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$36 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$37 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$38 \$9 ISBCS ISBCS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$39 VSS ISBCS \$9 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$40 \$10 ISBCS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$41 IP ISBCS \$10 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$42 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$43 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$44 \$20 ISBCS IP2 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$45 VSS ISBCS \$20 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$46 \$21 ISBCS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$47 \$58 ISBCS \$21 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$48 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$49 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$50 \$28 ISBCS IP2 VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$51 VSS ISBCS \$28 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$52 \$29 ISBCS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$53 \$58 ISBCS \$29 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$54 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$55 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$56 \$38 ISBCS IP VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$57 VSS ISBCS \$38 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$58 \$39 ISBCS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$59 ISBCS ISBCS \$39 VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$60 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$61 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$62 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$63 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$64 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$65 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$66 VSS VSS VSS VSS nfet_03v3 L=6U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
.ENDS CM_input
