* Extracted by KLayout with GF180MCU LVS runset on : 03/04/2024 17:11

.SUBCKT clockGeneratorLayout GND VDD IBIAS OUT
M$1 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$2 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$3 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$4 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$5 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$6 \$54 \$54 \$57 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$7 \$28 \$54 \$58 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$8 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$9 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$10 \$58 \$54 VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$11 \$57 \$54 VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$12 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$13 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$14 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$15 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$16 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$17 \$189 \$191 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.52P PS=5.3U PD=2.52U
M$18 VDD \$191 \$189 VDD pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$19 \$189 \$191 VDD VDD pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$20 VDD \$191 \$189 VDD pfet_03v3 L=2U W=2U AS=0.52P AD=1.3P PS=2.52U PD=5.3U
M$21 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$22 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$23 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$24 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$25 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$26 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$27 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$28 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$29 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$30 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$31 \$189 \$191 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.52P PS=5.3U PD=2.52U
M$32 VDD \$191 \$189 VDD pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$33 \$189 \$191 VDD VDD pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$34 VDD \$191 \$189 VDD pfet_03v3 L=2U W=2U AS=0.52P AD=1.3P PS=2.52U PD=5.3U
M$35 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$36 \$47 \$299 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$37 \$48 \$298 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$38 \$48 \$298 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$39 \$47 \$299 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$40 \$47 \$299 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$41 \$48 \$298 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$42 \$48 \$298 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$43 \$47 \$299 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$44 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$45 \$189 \$191 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.52P PS=5.3U PD=2.52U
M$46 VDD \$191 \$189 VDD pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$47 \$189 \$191 VDD VDD pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$48 VDD \$191 \$189 VDD pfet_03v3 L=2U W=2U AS=0.52P AD=1.3P PS=2.52U PD=5.3U
M$49 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$50 \$48 \$298 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$51 \$47 \$299 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$52 \$47 \$299 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$53 \$48 \$298 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$54 \$48 \$298 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$55 \$47 \$299 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$56 \$47 \$299 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$57 \$48 \$298 \$189 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$58 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$59 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$60 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$61 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$62 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$63 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$64 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$65 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$66 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$67 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$68 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$69 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$70 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$71 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$72 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$73 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$74 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$75 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$76 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$77 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$78 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$79 \$391 \$191 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.52P PS=5.3U PD=2.52U
M$80 VDD \$191 \$391 VDD pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$81 \$391 \$191 VDD VDD pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$82 VDD \$191 \$391 VDD pfet_03v3 L=2U W=2U AS=0.52P AD=1.3P PS=2.52U PD=5.3U
M$83 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$84 \$438 \$299 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$85 \$427 \$505 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$86 \$427 \$505 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$87 \$438 \$299 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$88 \$438 \$299 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$89 \$427 \$505 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$90 \$427 \$505 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$91 \$438 \$299 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$92 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$93 \$391 \$191 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.52P PS=5.3U PD=2.52U
M$94 VDD \$191 \$391 VDD pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$95 \$391 \$191 VDD VDD pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U PD=2.52U
M$96 VDD \$191 \$391 VDD pfet_03v3 L=2U W=2U AS=0.52P AD=1.3P PS=2.52U PD=5.3U
M$97 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$98 \$427 \$505 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$99 \$438 \$299 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$100 \$438 \$299 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P
+ PS=3.52U PD=3.52U
M$101 \$427 \$505 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P
+ PS=3.52U PD=3.52U
M$102 \$427 \$505 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P
+ PS=3.52U PD=3.52U
M$103 \$438 \$299 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P
+ PS=3.52U PD=3.52U
M$104 \$438 \$299 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P
+ PS=3.52U PD=3.52U
M$105 \$427 \$505 \$391 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P
+ PS=3.52U PD=3.52U
M$106 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$107 \$391 \$191 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=0.52P PS=5.3U PD=2.52U
M$108 VDD \$191 \$391 VDD pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U
+ PD=2.52U
M$109 \$391 \$191 VDD VDD pfet_03v3 L=2U W=2U AS=0.52P AD=0.52P PS=2.52U
+ PD=2.52U
M$110 VDD \$191 \$391 VDD pfet_03v3 L=2U W=2U AS=0.52P AD=1.3P PS=2.52U PD=5.3U
M$111 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$112 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$113 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$114 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$115 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$116 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$117 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$118 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$119 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$120 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$121 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$122 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$123 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$124 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$125 OUT \$659 \$642 VDD pfet_03v3 L=0.6U W=0.6U AS=0.39P AD=0.39P PS=2.5U
+ PD=2.5U
M$126 \$642 \$654 VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.39P AD=0.39P PS=2.5U
+ PD=2.5U
M$127 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$128 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$129 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$130 \$645 \$618 VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$131 \$646 \$618 VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$132 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$133 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$134 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$135 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$136 \$618 \$618 \$646 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P
+ PS=3.52U PD=3.52U
M$137 \$654 \$618 \$645 VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P
+ PS=3.52U PD=3.52U
M$138 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$139 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$140 \$724 \$724 \$725 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$141 \$299 \$724 \$726 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$142 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$143 \$709 OUT \$659 VDD pfet_03v3 L=0.6U W=0.6U AS=0.39P AD=0.39P PS=2.5U
+ PD=2.5U
M$144 VDD \$28 \$709 VDD pfet_03v3 L=0.6U W=0.6U AS=0.39P AD=0.39P PS=2.5U
+ PD=2.5U
M$145 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$146 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$147 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$148 VDD VDD VDD VDD pfet_03v3 L=0.6U W=0.6U AS=0.696P AD=0.696P PS=3.52U
+ PD=3.52U
M$149 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$150 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$151 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$152 \$299 \$724 \$726 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$153 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$154 \$724 \$724 \$725 VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$155 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$156 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$157 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$158 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$159 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$160 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$161 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$162 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$163 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$164 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$165 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$166 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$167 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$168 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$169 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$170 \$726 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$171 \$725 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$172 \$726 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$173 \$725 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$174 \$726 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$175 \$725 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$176 \$726 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$177 \$725 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$178 \$726 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$179 \$725 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$180 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$181 \$505 \$505 VDD VDD pfet_03v3 L=4U W=5U AS=3.25P AD=3.25P PS=11.3U
+ PD=11.3U
M$182 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$183 \$725 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$184 \$726 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$185 \$725 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$186 \$726 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$187 \$725 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$188 \$726 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$189 \$725 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$190 \$726 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$191 \$725 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$192 \$726 \$725 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$193 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$194 \$191 \$191 VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$195 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$196 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$197 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$198 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$199 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$200 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$201 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$202 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$203 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$204 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$205 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$206 VDD VDD VDD VDD pfet_03v3 L=2U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$207 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$208 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$209 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$210 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$211 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$212 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$213 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$214 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$215 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$216 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$217 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$218 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$219 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$220 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$221 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$222 \$47 \$47 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$223 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$224 \$47 \$48 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$225 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$226 \$48 \$47 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$227 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$228 \$48 \$48 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$229 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$230 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$231 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$232 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$233 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$234 \$28 \$48 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$235 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$236 \$54 \$47 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$237 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$238 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$239 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$240 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$241 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$242 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$243 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$244 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$245 \$46 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$246 \$46 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$247 \$46 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$248 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$249 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$250 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$251 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$252 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$253 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$254 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$255 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$256 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$257 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$258 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$259 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$260 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$261 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$262 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$263 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$264 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$265 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$266 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$267 \$48 \$48 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$268 \$48 \$47 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$269 \$47 \$48 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$270 \$47 \$47 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$271 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$272 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$273 \$54 \$47 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$274 \$28 \$48 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$275 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$276 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$277 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$278 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$279 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$280 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$281 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$282 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$283 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$284 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$285 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$286 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$287 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$288 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$289 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$290 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$291 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$292 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$293 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$294 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$295 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$296 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$297 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$298 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$299 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$300 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$301 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$302 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$303 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$304 \$240 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$305 \$240 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$306 \$240 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$307 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$308 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$309 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$310 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$311 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$312 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$313 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$314 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$315 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$316 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$317 \$240 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$318 \$240 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$319 \$240 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$320 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$321 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$322 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$323 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$324 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$325 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$326 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$327 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$328 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$329 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$330 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$331 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$332 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$333 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$334 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$335 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$336 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$337 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$338 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$339 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$340 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$341 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$342 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$343 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$344 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$345 \$187 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$346 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$347 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$348 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$349 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$350 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$351 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$352 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$353 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$354 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$355 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$356 \$46 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$357 \$46 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$358 \$46 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$359 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$360 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$361 \$56 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$362 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$363 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$364 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$365 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$366 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$367 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$368 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$369 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$370 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$371 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$372 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$373 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$374 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$375 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$376 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$377 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$378 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$379 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$380 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$381 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$382 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$383 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$384 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$385 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$386 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$387 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$388 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$389 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$390 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$391 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$392 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$393 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$394 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$395 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$396 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$397 \$708 IBIAS \$56 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$398 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$399 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$400 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$401 OUT \$654 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.366P AD=0.366P PS=2.42U
+ PD=2.42U
M$402 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$403 \$438 \$438 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$404 \$438 \$427 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$405 \$427 \$438 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$406 \$427 \$427 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$407 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$408 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$409 \$618 \$427 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$410 \$654 \$438 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$411 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$412 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$413 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$414 \$708 IBIAS \$56 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$415 \$724 IBIAS \$187 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$416 \$708 IBIAS \$56 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$417 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$418 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$419 GND \$659 OUT GND nfet_03v3 L=0.6U W=0.6U AS=0.366P AD=0.366P PS=2.42U
+ PD=2.42U
M$420 \$659 OUT GND GND nfet_03v3 L=0.6U W=0.6U AS=0.366P AD=0.366P PS=2.42U
+ PD=2.42U
M$421 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$422 \$427 \$427 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$423 \$427 \$438 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$424 \$438 \$427 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$425 \$438 \$438 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$426 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$427 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$428 \$654 \$438 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$429 \$618 \$427 GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$430 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$431 GND \$28 \$659 GND nfet_03v3 L=0.6U W=0.6U AS=0.366P AD=0.366P PS=2.42U
+ PD=2.42U
M$432 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$433 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$434 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$435 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$436 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$437 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$438 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$439 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$440 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$441 GND GND GND GND nfet_03v3 L=0.6U W=0.6U AS=0.672P AD=0.672P PS=3.44U
+ PD=3.44U
M$442 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$443 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$444 \$708 IBIAS \$56 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$445 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$446 \$724 IBIAS \$187 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$447 \$708 IBIAS \$56 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$448 \$724 IBIAS \$187 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$449 \$298 IBIAS \$240 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$450 \$708 IBIAS \$56 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$451 \$724 IBIAS \$187 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$452 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$453 \$708 IBIAS \$56 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$454 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$455 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$456 VDD OUT \$708 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$457 \$299 \$659 \$708 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$458 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$459 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$460 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$461 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$462 IBIAS IBIAS \$46 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$463 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$464 \$708 IBIAS \$56 GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$465 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$466 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$467 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$468 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$469 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$470 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$471 GND GND GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$472 \$191 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$473 GND \$46 \$191 GND nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$474 \$191 \$46 GND GND nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
M$475 \$191 \$46 GND GND nfet_03v3 L=2U W=2U AS=1.22P AD=0.8P PS=5.22U PD=2.8U
M$476 GND \$46 \$191 GND nfet_03v3 L=2U W=2U AS=0.8P AD=0.8P PS=2.8U PD=2.8U
M$477 \$191 \$46 GND GND nfet_03v3 L=2U W=2U AS=0.8P AD=1.22P PS=2.8U PD=5.22U
R$478 \$2281 \$505 GND 98000 ppolyf_u_1k L=98U W=1U
R$479 \$298 \$1737 GND 98000 ppolyf_u_1k L=98U W=1U
R$480 \$1955 \$1737 GND 98000 ppolyf_u_1k L=98U W=1U
R$481 GND GND GND 98000 ppolyf_u_1k L=98U W=1U
R$482 \$1955 \$2172 GND 98000 ppolyf_u_1k L=98U W=1U
R$483 \$2281 \$2172 GND 98000 ppolyf_u_1k L=98U W=1U
R$484 GND GND GND 98000 ppolyf_u_1k L=98U W=1U
C$485 GND \$299 8.4e-13 cap_mim_2f0_m4m5_noshield A=420P P=104U
C$486 GND \$299 8.4e-13 cap_mim_2f0_m4m5_noshield A=420P P=104U
C$487 GND \$299 8.4e-13 cap_mim_2f0_m4m5_noshield A=420P P=104U
C$488 GND \$299 8.4e-13 cap_mim_2f0_m4m5_noshield A=420P P=104U
.ENDS clockGeneratorLayout
