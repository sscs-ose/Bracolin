** sch_path: /home/gmaranhao/Desktop/Juan_bracolin/PICO_contest/CDAC/Differential_capacitive_DAC/xschem/Differential_capacitive_DAC_array.sch
.subckt Differential_capacitive_DAC_array VD Bit_3 Bit_8 Bit_5 Bit_6 Bit_7 Bit_4 Bit_9 Bit_10 Bit_2 Bit_1
*.PININFO Bit_1:B Bit_2:B Bit_3:B Bit_4:B Bit_5:B Bit_6:B Bit_7:B Bit_8:B Bit_9:B Bit_10:B VD:B
C1 net1 Bit_1 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C2[1] net1 Bit_2 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C2[2] net1 Bit_2 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C3[1] net1 Bit_3 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C3[2] net1 Bit_3 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C3[3] net1 Bit_3 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C3[4] net1 Bit_3 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C4[1] net1 Bit_4 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C4[2] net1 Bit_4 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C4[3] net1 Bit_4 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C4[4] net1 Bit_4 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C4[5] net1 Bit_4 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C4[6] net1 Bit_4 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C4[7] net1 Bit_4 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C4[8] net1 Bit_4 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[1] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[2] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[3] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[4] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[5] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[6] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[7] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[8] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[9] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[10] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[11] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[12] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[13] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[14] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[15] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C5[16] net1 Bit_5 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C6 VD Bit_6 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C7[1] VD Bit_7 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C7[2] VD Bit_7 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C8[1] VD Bit_8 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C8[2] VD Bit_8 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C8[3] VD Bit_8 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C8[4] VD Bit_8 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C9[1] VD Bit_9 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C9[2] VD Bit_9 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C9[3] VD Bit_9 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C9[4] VD Bit_9 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C9[5] VD Bit_9 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C9[6] VD Bit_9 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C9[7] VD Bit_9 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C9[8] VD Bit_9 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[1] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[2] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[3] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[4] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[5] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[6] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[7] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[8] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[9] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[10] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[11] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[12] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[13] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[14] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[15] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C10[16] VD Bit_10 cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C11 net1 VD cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[1] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[2] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[3] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[4] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[5] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[6] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[7] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[8] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[9] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[10] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[11] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[12] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[13] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[14] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[15] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[16] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[17] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[18] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[19] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[20] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[21] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[22] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[23] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[24] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[25] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[26] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[27] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[28] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[29] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[30] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[31] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[32] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[33] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[34] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[35] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[36] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[37] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[38] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[39] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[40] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[41] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[42] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[43] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[44] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[45] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[46] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[47] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[48] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[49] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[50] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
C12[51] GND GND cap_mim_2f0_m4m5_noshield W=5e-6 L=5e-6 m=1
.ends
.GLOBAL GND
.end
