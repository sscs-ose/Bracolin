* NGSPICE file created from PR_net.ext - technology: gf180mcuD

.subckt PR_net VSS VC VG_N IB_N VDD VB VA IB_P VG_P
X0 a_387_2075# VG_N VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X1 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X2 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X3 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X4 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X5 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X6 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X7 VC VG_N a_387_151# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X8 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X9 a_375_8672# VG_P IB_P VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X10 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X11 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X12 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X13 a_375_6740# VG_P VA VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X14 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X15 a_1781_8672# VG_P VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X16 a_1781_6740# VG_P a_n135_3233# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X17 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X18 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X19 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X20 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X21 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X22 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X23 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X24 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X25 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X26 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X27 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X28 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X29 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X30 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X31 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X32 VDD VG_N a_1791_1309# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X33 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X34 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X35 a_387_151# VG_N a_n135_151# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X36 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X37 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X38 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X39 a_1791_151# VG_N VC VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X40 a_n135_3233# VG_P a_375_9838# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X41 VSS VG_P a_375_7906# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X42 VA VG_P a_1781_9838# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X43 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X44 IB_P VG_P a_1781_7906# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X45 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X46 IB_N VG_N a_387_1309# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X47 a_1791_1309# VG_N IB_N VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X48 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X49 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X50 a_n135_151# VG_N a_1791_3233# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X51 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X52 a_387_1309# VG_N VDD VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X53 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X54 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X55 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X56 a_n135_3233# VG_N a_1791_151# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X57 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X58 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X59 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X60 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X61 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X62 VDD VG_N a_1791_2075# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X63 a_375_9838# VG_P VB VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X64 a_375_7906# VG_P IB_P VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X65 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X66 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X67 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X68 VC VG_N a_387_3233# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X69 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X70 a_1781_9838# VG_P a_n135_151# VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X71 a_1781_7906# VG_P VSS VDD pfet_03v3 ad=0.84p pd=2.84u as=1.3p ps=5.3u w=2u l=2u
X72 VDD VDD VDD VDD pfet_03v3 ad=1.3p pd=5.3u as=0 ps=0 w=2u l=2u
X73 VSS VG_P a_375_8672# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X74 a_n135_151# VG_P a_375_6740# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X75 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X76 a_1791_3233# VG_N VC VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X77 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X78 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X79 IB_P VG_P a_1781_8672# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X80 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X81 VB VG_P a_1781_6740# VDD pfet_03v3 ad=1.3p pd=5.3u as=0.84p ps=2.84u w=2u l=2u
X82 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X83 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X84 IB_N VG_N a_387_2075# VSS nfet_03v3 ad=1.22p pd=5.22u as=0.8p ps=2.8u w=2u l=2u
X85 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X86 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X87 a_387_3233# VG_N a_n135_3233# VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X88 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X89 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X90 a_1791_2075# VG_N IB_N VSS nfet_03v3 ad=0.8p pd=2.8u as=1.22p ps=5.22u w=2u l=2u
X91 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
X92 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X93 VDD VDD VDD VDD pfet_03v3 ad=0.84p pd=2.84u as=0 ps=0 w=2u l=2u
X94 VSS VSS VSS VSS nfet_03v3 ad=1.22p pd=5.22u as=0 ps=0 w=2u l=2u
X95 VSS VSS VSS VSS nfet_03v3 ad=0.8p pd=2.8u as=0 ps=0 w=2u l=2u
.ends

